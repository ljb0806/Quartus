��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`����<�V0`Q��ťɊ#�MwU�P�X���s��j8C��eZH�4�L���M��-oi佴���y�w��KX2���M��f�� rF���O`)���3������Ў��T����.���FN�Oݯ�����U��&~��Ōı�r�j���'���6��`bFM,��g:8���?<p�U+�k|YwIj�F�C�&�5�v�0��c���8�N枫?K���|څ�m�!�����8z���|[�pz�<�����ާ\�[s���J�0���S��f`$�z�>$��>H�{`��s �=Os��a��73ݯ5���N�sx�� &��n��z������t���������n��#/r���y����~�>K��3fď�k��c@�pS�i�D���� @�biMYl@2��ӅfznDO/v���K}�dq&�K@�BK�|��I�dP�?CcRB�ewⱰ�1�,2I�n��	����U�I�	P��YaLr�q�U�$Q���@�b�cA@�v�ԫH8��,y�J�3c7� Dh���?�3Q�����˛He� t���s� �Z��0�*��R���h���JyǱU\\�RR��ڨ<=��Կ�Od�|�@�~W���!��i��H�������+����ꤺ!��+�M&i�yB먪�0�a�{��m. ��Z2l�]�c;eۢ8e��� ~�[��Μ N^av�A�0ׂK(#�gr�,t�`;�X6�{���>���� G�j�_w=lQ������V�R���՝��,�Y�dfv��O�r�݄�9�[�_�u����bD�ij�TM�c�D~�0�,Yӂ:]3���W�W�����|�E�2�lY�>���
�U�HkV��Y������
� ��E0��!�{��N�Nl?b"�lK&jS'�E�<m@Ծ6w�1�z���,,{�DM���O��	��Wϕ^._4�uLL�{�;<B�S�|]S�iC�:7zٓx�����v;�C�s޾?yc�s��ٰ]��.��軷n�+ޤ�IH��ږ�w����P4�q˜�-�c�ɋ�T�$ڴ`�n�P�;a�~�M�پ�m��p�iO��Ť����k\/b�e�=Ǉ��Ir	��W�h�Tk54i?� �{)"!���t���Ő����0R��W�����_03�~��#�AƄ)��"�ap��L��0{c,]ATDĨL/�/�hPι�J�)fc#�4(�<�u�-�Ų��� 1rm�6�Lԣk�2�\$?^O��q��&�HE���6�뤿{Cܥp�=Υ'$��� 1|�D���X�ۣwN�8�����*K�#��%0R�������A.���Z<�y��#�0���x5���!�ELH�͝�[�d8�z���D�iǕ�R�c����TjM�輼,T�m֢5�y���=��cI�C���n�qۯ�`�b��h��ĭ�! �?��'s�:�#@ �,�`^'����q�	�l/��KGv��T
#��Ot�п��4��*�SL����f�i����KL5�aF�4)����pr-����ם�g�h䪠2Q��i�C���1�$�5$�*{����/�w��ap!A��*��@'���l�کiz��o�Aa�+=�	׆IQ� !{[C���ڱ)ٷIl�`�8��f����9��&�X��6���s'�x�i�.Y\�1��z-�$ԥe����f��:9j#���B
W���)�(�*��qO	�����e��L?SFGP2���(VUd8\�����.mx�rը��r߀^��l	��^�4z����M���{7& ���(�h_1��bV����OBA��~'�h�)�8n�{���[	�l��(@���00�
�R��g4�k��Aȣ�0o��g����,
���f��Z��F����mwc:�w�c����>�N9�F)�o��Z���A��u��R��=}�e|�b��Lh��H�#��]��p��N8��j1���Ğ�-���� E���o�1[S��`)���Ôl�>R> ��dJ4���Ѳ��E��p�}�X�On��3i�p�aM�u׻�#��n�Bn�4��>B��f��uu�p˱(���A���`r����-�I���/���>B� ������:�b��/�B���p(o�J�Y�����;:"�8����6� ?�t=j.��D����2�!)!q:M������Au������i¶��D�����p����;�46T��T����Yb#�҆@�䰭������D��$m��g�����	�}LB���s�]Lս\�l�!؏w�c�C�����3��[��R���iF���[}��ι�l�;�l�W�	U�*��q�� �GS�11��e,�i�Q�p�#�ƤG�]ab{���hn��e ku"_�{�$s(�Q%��`I0�>'��AZq�9��c[�|���t�H\�2�Y�NB��rMrSZBȚ�r�=�A۵����+8[����Sd��uO��P�`;��x�p�D�(^��>|#�  �ܙ�4.HW��+R��O,\��:t\i@
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
U0Cxj/qh3WJ0XqiaKbrHqO5prYe5jn1r+xbvD+oPufkxSFNETvuInzlSg/GPq7b+pdjlBsiT0qBt
r270umIrJzuFq19oNJrijNIc4LS+cmWp9CFxmfV85EPJYZRY7cWjFjUUysiOVjUUXILNbQJB8Cuq
O6GgkYGWIrcpk+/1Kb0JqD3vCdxrgxp42/KTYIwW4UINoaqXow7S+prDNr3Hrh5U8uQeeiOv23D/
dSwLY0qCw5MMATxI04eOs/aD2AsC5JQ02CgSsGSfsy+ZHo5KdVjTduRElWgRrQ3UW23sc9xDJZzS
XaTyrI7X5fNK8h2UD1MdYC9jebtCEFfb6SPlUw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6784)
`protect data_block
soPOf68o7/noxlWY9CwCluw/icMLkhZDw84t17TgTNyocTz8ThTJ38jgNdw5Jh3WprSz1mhrvQHS
LJQzhssh1vjDcxjK2rGnBq+jdnwqfeEFnzbjaAiCxXwQhhmPjoOUKqWauZur+FP985o+/tsEU5Ep
BGquYaKZ5gD7x71BA5LAmDOzXg7YhJv29+40R+sTygOvUG2/nRCWt/rcyFGGtlIHJSUVNf9Rj/i0
fr2VT7rel5rCp+RsL4c+h5gGFIukru2KmMCd/8+5h3o3Omx50fstOYBYc/rM8ECir4/1Lw5ZA8Bz
f7UQlJE8Tb/EwIKarGdAUnpUCNPkds8ICeEjLDeoq1RvyFORa2xYdvzpM1SC0RV5qKOfDdtbLF4e
tccTaj0G0/s8EvpfSyT3M7qX4yaWv2HN3CMeQxZ/YXkE8CjyrVwEkCwdIsUvUMIFEwR2y+C+0bWH
1oZre21/mVoOmFq3icH/fj6wf6DMi954llYwBJ4b+5NUmakYpI0F0yN9BmrXCix5T8L+rwxSke1W
5CzlMZm7yL6VjHqSnpkMNglhkKmED6huI7dxpP7umUNn3pD1Sq8Dz5SeYjJSGs/tI8KN2TvNaxkn
gsKKd39f3xqBjr1VdDMlPm3eqDeI0zBDiOEDDmaowV4dm5pMQNzHfvHsE0MVlv2TNYs7Yl9QQZRB
6g7RfO7RYu2GnPcxzbs5m3+DUqmSOCXdakyjKIkH/Xkzpw1MvBqY9LZJvb1R8TwDYk9CUGzNKQCX
czLKumQP3Ywy0xytCa5epamb1LNkEfRdjmIA1lNMHG58K4Y8CS2PDZkEYYmK2yU9/RQ8YvVQ0Dhl
Z3Wa+xxsoMrOrvypE8YrX3pow0q/n0yg7qdUzBk/AY0le0TAoXUwUwlnu5Tvs98LuI9TEsdGLwOe
3fK6QnqHcv4OVB13c/tYVIpBkDuSfE4AnAiPsKvgz+K6fEqf7+8Vzhm5QzkcJb6L9I8mSZaFdizL
cLccIHSigOqvYeVaNp07/fPxJot3zyFgYnKD8jM9iWI7Ikwb+M+iwSmxY1qcSqVk0hvYwUOOIAUy
4elqNYGqi1n1h6ytaYzP0wv8M7UCnXi/ixWV/zcJADJ6JmdE0CoKBwRrWm8NfbhLHtj3QxFsRlX0
xuwlYOBa3uV1Q9KRHlEWiuRXDawPMi5hk7AAptTPNxr6aiWF0lp1sZ/R1tAbGMwN3ufaV5hNwia3
8SJTLkMLFK/nbkcIjdHYwz7VOT/Jk4+0XVugkgUn4rq/dopwzYB4n5R+v/snlvRYSa9/G1f4ZS3O
J2lwWhjGZQ/rftroHp+cZspsYUrQPFpqa6ksxYAs71Zmzd+KHgyyZvi9vDtylkpS95wnjn0F/TZd
v9W5U9kumurljdYO5CiEWzudOaHUQumspI5DBV5A1iQ7LuzvjKM4A3T0jEs8FMrujAlLQJNM4ge9
G62svVVdz7durn3XjEucmm9uOWGPbKeFYFhEgMtmeScNj33GuUay50hkrRwHaLAG6iPB7pbqKtgF
DyDVZSWUrzRlUtdeHVveev9bD73yIaRPp0SwQ6nVYIx3I8bUPmHvS/FDEWL+SSA9lkrrHl5KdaA+
mpsQBmFlwMnf9+VmLJO80u09EE2+stYyP5aEZHPeS+YCUkt8ZyCKxct6wdCQixtee28j/1vKQa0e
aaicoWU6IzTFvQDKEEKucGs8yOUkT3nkhz+CuovWFIjG3WoayJQQrEd61LhC1aarfhbazKuwoP5G
6k008LcKCYCq16/k/t48wTzaOWhMlq0+xdmGto9pY66QvM0dsZK2TZ7wnfsbVkLvSUjxaZlKY2MH
RxivSkaDx90aj6NDImPq/ZnEByi6fiJPczNY0vaJTEdaMVy19ndJedE5YGTrnDnuZIxGeiMGMK/i
lwkzKAkcpK663TuAyFjTUxPNkO9wezY2JUbNf7FT4hpXsDg3J+S1N/+9JXNlOKHeRL17j9UoPrhN
rZPr9kEDn5Wj2WpqanGzJB6NCxBjIOGVGsWbKBdm8mJC4Lgg9z9K6jEBW7SDCm1J7iFvqUDuQFO1
6rOGQD6xZA7pk0b5gbDy1Dwi96abqrH+ymE34jvOFemGs6Nnw0wotC1rZ2yHGlrr0ym2/jVvoi9g
6YN/tlQkUIvEPy/qhTmfj9LYb3npVxHYLCnyOZjKk6GWt7P+jVUdEJupKzmGLDnz6GrXz2i8c206
KBTw3xk0XGCl7zue9iO+99X61Uu39wI8tiwr/uRG1Mkh73a9R9SKf3g3Fgl9nDO68FbX+veel7Ey
EXPj3toubxqE8DNX3HpfmXGrfJAwFN+QGv25ad+nPTJQW+UFdwrH9WWK2TYDt894VDE8gqNnvc9D
QRSyQldhh44W2KHSEAIclmHM0aoKftOYVxpDTaKqWOExG4ZgU63yGaHoCfYO+SoKtxvDyvaRtIIl
u6ZubND2Ds/SRW9gXAmubrls8H+wH8g2SPbXe7nvcUUDlwqJ5U1G//HHlPk+JNY8mw8xUaZKNeeO
5Rq6L1RkX38VZ3UXSEjk0cLmKiL4Ol34J/hia2X7dOUJLDiNNvxdhyJf7FhDmjoJ46pc4cAMXUWy
isGBR71qLLFd0PvM0Swq27f75wVP1bkZsTJrFDQW/sNhvhWeRcBwMa6WA2dTEi6tc1OF+zlJErlR
bBD8SYwDFjHLvU7QbHpNMr80f5RtfbVy/Ps6/zzyuRaZKVD+6qtswQhtrjn8Kaq3qS1YopIqyGr9
8dc4Rv426qJD/vfs44lgLBCjR+SEJzgV7zEG9Y67MoiXSZK13tCnHoc8i2TtjOQGxUmgNwkc7/Uk
JOevam/vuO2nLOx7RxvSH/IUUsxAQ0H7ikyl4HAZH6G2CKetN/dYS8mJ/5ovLb76uV2d2qYL7bKv
5LKCWlYx+KN83vwXNlrwtE0V6f1Li/nA8eyHTlEPJyoqZgYxb+Xh2Ac4tzBnrzHMYv7Olcox5TJl
BvQYueohl0tCmmrAm2ABpfELh/fExRoRjCxNxpmqaQlKQ+2LniAqXh1SAStaAWL4Y7OLuuGXP72A
6VdGOhM0lfTunjP7c2RicT/mBYESNpDtuNUvHPnopJeuRadYUvPOb+Vq0mdeq1u0zUUNSWHQh5tk
Ekmz++DRWj5lYXPZcdinMV+eDnRabqz4AxhTZp2NaNjwI3Omuftze3BUIr5OrWtReDEeLjTPpKKN
r+o3ASQtWNG0qw1EVjNwvjhmS/lBoCUEXeNx8PFMK+svszJJBApRrInI9nmSsjbT8pRUm3tmJQTo
4QMzgEyx6cQwL23eVbaG4dovCRsjvt+7mCf9ltxFqUjRkZs+cXlMdBi6yHVpRzlx3K8FfhQdB9+K
yJUImXHwp1GGuUq/JByAjXtfu0juFuWglsa8CKqhpVjeRb6fd+chLB6WMz/5kN22KryIBMnAojkb
MWF0BmdPqJYU8uoKMzaOkb3p5BomZYjB/BT5QKYfuKT7DS0EA/CW0GG/LAJkdeSnSrBER2gheSiC
8QfjzBVzXgrXWfiGPkiWxa3vZjSBykFpynerf2p4o7wJVEGQdGa2fqScv7FBui3Iiw5CLgDQKxff
QJvfbVP5isZ/aL2jbSIwdIvgCbsow49+qnZ4A0oUQ1TNOleftHdBxapk0GIYPBKIIJLuv0vmgwjx
JFEtDGfv/o8/OokY2jpjyanxEc+drxvF2UUFEU3zWfbJkUSMg1rsJxbFx3r70lw8CbY2a3mr66tj
ysI2ltCTe8H2IpG7ZKA7daYbhvD7pZ5+OKAX3AHeUNVckLfDn1J4EL5UPgfbfTRQfGHq4Rw0ON0Q
gRBzlmH5TBxdrJPj1dZv9i6/kd/4kOTaZdthVsAPnmvbs0hRqpgF3wiYazv7i2NIQz4uKIDhGw4C
NOyiwc4/TxNwPv6Q94wZwHzxIEyQPDct3VxOyYhbmLDvxciXWnj18ToUr7GOftpAX96wBPmkKJ9k
RQJzwRUJTjlYrpsovSDK/btanXBp4g2bnhH8xffDDltJAHzAY4xYzDSwq9vVHEOu8G3gHqhpi+ft
26tTx8l0HJJUKvjIRPYTObc26qn6MEEtsjvRyunwB4+62huWz3+j6XYFW+eb7Z7oltoIEqtnF6F5
CHN43QlgObyF5Sjzf4FYnqRMy8N3eL/jyhaYSbCjIuJDHsxBfcjy9vrfoeZ49hU8FT6kQF2NP50t
9c0P6opZr9nAZPyCe3ev41PQdbB1Ep1w9moGjW5RjD1UUQS9hBSFEy8EGpKasL9G1qEDEUeEv3K6
u2jMQaLnZz3FprpgEphlZQBsOqsU5O8/RKeYtqspp1g1pOyGgrt7mWanlQl9bp37biMGkYp2fVX7
SdN80/CG8TUTNu4ad2Vxp17sgsiCo9xwUTJvRqsKIVe7Zbuyazis7GLxVDwQ3evZF5rCAsNsfDjD
ZetolBxOO6KxJ/wkNADxg+RGSGxnQPrAOuj9eOUmgeWYI14d1hZYEmNsJEFcEt9ULyO8WBkbdgnO
BmeSRwyv0CMspj8C2NJnhTpDjEHstr1fS7hzP8JLlxqO01Trg4RaOUhP4eoZ5OzqbdtrfAjZ9yQ2
8PZtmLwMntio9FkHE75D8FTTDn+2GSg6ftTGadWn2WmV2xxuqeOSjWYviuRCuOtjS+jomCUkpReN
muDOTtqlcmMAVu/9Z0qGIJM9DH/+bFiHaHbEBlPeKX5C/SEGK/Q6uAr8N3fPN0Zpb/2JCRAQ7IbH
SU/BTEDakTidyQh3wYona/JaqU9vmQ+k3CM/1OILkL1RUQFQzlv4l/+oUcVAUvVOCcWnO0GjTYaX
mLz5dSqDF0LPJrXOWAl2FpOfp6Bf+59ubv8gkxetplf9FFhW9M1BnF7VK0tk4IkCi7Kx4e2PXVp1
m6w3bnTazhzyvV8QIt2dN8sscp1HpIs1clrXTtAVA+aqDV5wO9qlAdS5yVnF7FGYxG8Qw28SokGz
KJEWJe1J33afHXk2L3GDo0Z68FmQopZ24X2qhlj/yPAhx5IA80iRkO6NJUtyc3KKQ9u3fjNCZsD9
0/lJ9kB+ORJLwW4FK0gDlcEXVJQZ/VUcdDEbtVchQrAfzFfcwSj13y4kNSvKUElFHc0RbEpP/EMP
mEQ/QnQ/EH3hcYghIvvoLCsN4Z+s3xbMqMsqYYYbOxEB6agwMUPbbgfHz1VS78BEa6U+tG5bNT8r
1cj5KAdPA72K3+NPgHfBf0SwNwF+dWo1/RVdrbFUmfm6OspA5kl7Y5iXOHYoid+axdBN511cfDpv
ioMLe+h5X19PmnHq3UbFKQ6vbHYv50GB4Mfjk5KSEvH7IyNW/74+D2JtfQdKJnCB4eRYYvrAru9D
IPH6KO/cgi30wYRCtDE3SY1UxXp/4wzRmyvwV/kE6so+G/VEQecFHuQRXJzgcB+NnypawL2lAMR5
/Sh11cvT8ZQCbPjyjSsk2rMzDpJTC2tgpzkEB9Mz3ZKhCKsS1FrbofkwN6AmiI1BR5yfkbpulB/C
efIvymsyongGg7kmTDguvnkOKu1Qm3zFB+tlcYlKtA16lc+x/WKt1uZo3sFYCH7BChzpFWwh0tJa
0TNmXcp/PJzcdqPpW3XB2fgQKdekSATJ0IEzHDucCiy0yWCu+NA/urcNc+whs596I2+56G83q+gz
Z6YmGE/we+ren94SvPm8WjBUt0+WbtAHYN3OU+w1Q/7lJAwQKB/0RDKwZxGtbTj83AlfNUpLhuli
XN2zq+drt/2OVIdTG28aP0MYlNhzxdPAcsXFc/Bsc2TQbuqnymJ8y/guOXTmpJBT1t5g6xw2eVyO
/8ZL5j8Z8ZRpQ1EyON9Z19Qj/ImIyKTI2dM+1bxcXz+jdrcC6EyBRoNdGRws0vi65GuT1bQvdzkn
CptTx3DUFhpxwjphNm0Y9rJN/cRWfOYB+FciicCuwZslQ3wFAukijUqCWcPWLo4J0GGuq5ovbQxh
5qapBlr99eHlHlw4xaJnwr9QfYHpp8f51aSrqpEl7cx55GxaC/4+xu1EsUxKrK8BQBRFiL4OstQ+
ouVUNxM8VQJBgToLmok8caWLTmn0HtJdL2CSJLehxWcZk6iQlltCmH0FuyhTDH8atxiNEkeqGOi+
MDbZVkIqq8GVM+XlkIOXBN8lMMaf3b4aIbYJPNiLIaBG66fh45miTmfIo2QtaDnDLtgqpALNy5Pm
49HH8WAtBgQC1sRIvJj4wkPRUpcCrwN/SRDKizHZs80KCbOCaZN5CFkvve5W3celZ3/YiaoKQuoL
87r+xPDLT5mvAiSx5vtcN6Rn60Dbz8CEJqjqBRgehmJvXa3bTCr3oWAp3iNgjamH9L9dNZ8f8x+k
LQz6op87W+LKUJugkN/pjhSkqfFE3yfavJJkWSpdEl4m+LBJS4xBac8knqqJ4lcCweNN8yFcRIdT
SxcLQ+4VfcOb/YMHvpH2s0zMpNrqIPI9723DR+2gCkZTFmTawNl2Kt7OzWFSUvFal2e5lc+K6M6k
qGMjHrgSlc+S5Bi14CzqGwjWzshlQN7h4L3upKxEb+bAJjDQWxb1PKuVbuEuu3xBWUJEGr4lBSr1
5b2b47Rxw5jvg443lYSOMsvXQ9RCLeGScstavdF0wmqZPrGwZ0/HcJZeKmIA13xyle1UNrIH4X/U
P17kIXBGcZ1kSeUY0U7Gy56GQQA8game0b6miFqylNnKk2abbI01BfQxAYEfBywc7f7jg0cxQf+r
Dp6WiBDqMA9KEY/sCkKr8iQ9g2Ya8LZBX06zEABa1Ylq8rlGSq7XBQvWRd/9PvvwylF5jdJ2byB3
ICoiL9GS0EDNNpq0ADJF2g04iHfbf47mLYXjWEYzTLRz5HwAFnyQ20J6/EysbsSX2I33ddRmyY1J
WVuhRNwnveU+qIAHMepyVoWrVBQjTQQoMm5GOVzfsap8ADFSQHHNCUpZh8MmEnkITsrPaN+peyIL
uAaBgIxH0+K92Bruew0Mn+QGRSoyflK+Usi9h3eYXrh0xJY2FR3qNLOLVeVOcSTVZO/WmJGHcprA
d/p6lZoc3ccZd+0J7Se/EnPOae8MptJudCYLrDg0cXnMxcGoE5zeaq/uo1yuoYy+1ZR5SAtfqkv1
HNW4V2SF+HmLIcY7kDkp582N909m6wJ+PCfptDKUriFDwdj65pyxETg8xaXF4N7arklvhuCBi0mq
R+48ikd0WzrEOJoEfzWz9HOpzi8+ktgRTBIA0d3y2fkR2iyQhU87b4NTBjdcCfidEeKAL9EVclTA
5xxoNGiQI0tjiZo7bYPpPx5aiMksNSenFdEZF2Bkv/T3IeDgfdnbjf7kEjbMv4kD24Zmut6uhl/c
QY6KfsWUDwozMiw1BRu3XRuzqXx1IYBGmURZBlN0pwZVFNR3yGOlScNDpTeEgSt2NN1IQvNd9jQp
QSpLQSWmry65UhFNKO1+dHjVrx9WHkjMvEGtfRuz+2i1fD89vnV7OGywheurXJX7io8Ishmz3jSH
g4FIZ65/95scNWPyLTTt9OP3qB9iP8B6ZZq/y3lqcMH3jyKUSevR0haUyJxqh6y2rmMYvqOpbzj+
GYea0S+ax5KPErhN9/FqLzRm/kPzSKF9aie3ppLO2V1m0Ds/iS/BsUHb/uGqM13UxnGNoDJxiaxB
zn4rECelBcpJXNmgEop69QG101yTj4/BrAECgb9V8UNQ4ywgaat1FNTeVx0Raag+f1oNuPMHIhUQ
10TCIch6rqciWFzJKnMqC++GZQKOyvTkay5vNbYcKlUK+ndR0Dm6KaVWUx39cDkzxk2y14Xd1Z+l
dXmGBYP30elRfyjRDOn8p9n+ykNJ+9nKCuGRYkLxtEvtyDrAI+hLymkenq/wuHon3Wx5cyS6GI2l
Go5wJuxMozqsZgLyp6xh4iIlepm7QtooG63PzfFr36GNBcAG5eRLutfkj7sE/JS/22xeAKqsTFcO
BDI2WyjT6WcsdGp1tBFUg9oA1QVnZlvTyv2tUDGFSy3hjL+zI9Covw1sJEeFcEetnvbBr7bBIhFc
fIqo6QPJSnslAVqlOfQvEgK5VPNLwFVlAtuudBLqRLKODD9P51RKgmPiRzMQP5ByENM3npdDmS+D
TSfCGWXqikYyUbQF1dznOo5/FyQDsHN4xBp5aHazLHR1555HXRjUJMq+KKsqBiLJOOa25O9XXGVy
AbTrIqJNbcXG5D+sl4Fr96x7JhzIbbH0+CN+2BHR2r/31nz+NABrfm4GBYjaMDI+f26DuNQRnpLH
DxylmfX8b5Q82/3Y3WlAlNiDIWZeppVWQUDiSIruJf9VzYdgCw7KfzMW53AmhXtipesr0eCBQe2/
55SvHi/4Db7sctKzcXp43KWirF1TEZmUUvjoU8PYouy0KvKAIImRrqy/LrZ3CK67gh9reqLtomgz
xkcx+hrQT+3XQ9uE0oJhXBCe2fSG9J7HLPC1NCt+LsFTt8mOaBTr/aKdX+iACeHLL5hIskuXIxTB
ygx3x8MFXstAOiVxtjVhgXqlIjyR/QG6vnTdNRuiS0ntS9f5rgY2LPmTmwnNrvG0ll3lELnG+2ef
SP9tR4a9MaLsAMbxV8Tpkee2SLpGegbc2BfFuiChTSX4uZlGdjPGsmIhJ9En6K9Wi6lEM5eMHXpb
R6TFDdLpguO5cuyhFos9TNCbcnwArlTh4RUr8QXAj2mOnYRNAt2FnSQkEgKeFPvBMuo258OImPsO
2M4G9Ev7abWnBuoFUmAyhnjE65EqVqefFGq7YB8jKme0LvHvIjAP78J18EkDcJu/gFgy7BycKuvT
9VxeQp68HmUNfG8BM+ThwtS9XNfJcyuUVNBAcwoMqIwxav/KhdVK1bazIe9tpE5jF/QfhWe4Sdxn
BBjyvhyx/lBnHBSWeLJEalKOFwo0T+TKywfScAr0jcI9xlZ+lun0+skbkQUiYoqYTXJ8nX4PP2KT
f2fE03eTu9HDOZWTc+wacX168u+zCFJc3Da3P3TjDahgDHmLxg60AvdSRH5cWDe+TauHGn9aqPzp
WYDwEESRBJeqlGfKV5tUN0MQZ8yDj//EKKabtyYywR2oG4xId9FbpT9/mW80ncQ4Npu3BNvAjK1F
Og==
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�C2��~[�X"Hl3G�z���'�K���6qַ}Y��.� N�v<�]�-��������l&ʛn��������?�y��C�'� ���,BY������B�6�i��z"{���j�M5��^�̺ �K�5W���\��x�1���Ė��	�@0u�0Ry �1Y8�������"�*��M�~�ft O�"w�xՄ��ب_?��.�A��0���0_�%<j�T)_xݑ�������M���S�l��ڿ�!AX�j�N�yov�u��>��2gi5Mlft"b ʪ+���Y��t�&��H�y�GEm��* ]VRg[����"�e@AF�U��˘l��cߎW&�(��қ3흽�.w�����zX�k����l��ez�m�K̅���qܱ�j-�H�^i������,JK�����ZZ�	@�o��չ�G���4%5��9���
��q)5�F��ga�A�_z�,t?��JB#H,�qJ�'L�ɱ�P4T��3������Y���=��7s��位%c�����qCӸ���S��SY���e��V-�!�N�ZD?�`������[���#t�b$����g�*�u���&�G��� Z?�!3c�Z�3��>��Dak/Bzc	n�%](wB8ߢ�]��f�ő9�z'����t.O:���5a�*}F����_�e��g�L��bS~0�Y������W���i���5�9�����8n}֟G���=[4>n(hnU7�=o!3U�j��wR�j�n����բ���!8�;mw�:G��e���H�z;�D�gӖ��J����_}��R��NB��ջ�>FC��1k�4�,���Lt��F�@a�9����k���&�)=��I�<��D�A���Z���(��?1<����h���С(?��&[ V�L�3 :۪�j����粬�&���/�s�����������r�%�1܃��g�%�x"�[�7�M�
À���laj�A
��J�����ADdw(`l��bHkN�nAI{��{R���͞��s�8�;r�ӈæ��'�H���\i��:��^��\��ե�̒�(D!^�T_M�ed���`}k2/�&���荜�7$#ޛ���a6�),���,5G�.�BO:w(�����*�F,/����xuw;��8 ��P"-M��7Y�侧�bl��b �ո���w,�4~�iY/�4m[$;�:X�p�ie�P�[��;Ȅϯ�q�V��[:O̙/+�ZP��m_]�ۍy0� �y�%OZ�������h����.�rr��Yg�0�o����E��T��R��9������?�ը6=O�9޾2�2eaz,�����/�=�C
���m�)͡��YL.7N��뿆fU�ՊPKk�Q��._�M�}������F"��k.�"��1?w�ae�w�p�w�mm������"Q�6���᡽�.���C1�h�G ,	�i�:�F�
lV���:kН篒E��~�9׼�>p/܉�R���'s��տz��*%��""��~��7< 9��{T�SlZ�{��!����7�CU������ �C���]���|X�ߔp^h�9^���{S�EJ���V�%�����Yw�;����^Iɒ�˶���6#��_)Q�<�Pٰ���Ǣt�p_���k�4u�,P�G�z|Bd}X��.�4�pa�D� �v�*(TyC
z��6G������{�ʊ5�C��I�r3ݞ��L6+5�+��I�d�H�:ԝ\?�����C���:�)��W��x���TB�	Db>�7��BU/.k���ĳ�|�����h��)��ō"�M$U5<2��";�X.�����ecI�j�_�U�5_�P<{�R,ZD ���pI�x�<�~c���u��{p��� ����LNi��+Z )��FN�lئ�%��ԧP���q��-S�n�!9�,WÎ���93�x�c�A���k�7�+�T�bK����,lW.3jV�fb�0�q�so�ǒS�\/.Z6��ÔE��#�O����q����m(�CۃUd��3��Fn�~�@�r�9��N3�p���yru{�t�D!`qߝ��(xW�8����]Z��x��k �/r�t�)�?�M�	�#l�������l�O�������kɖ��n��xݒ؄4w���zk�P#?X�A���rX;��щ����o��boc�A�G���VG��B-�A.q�3�<���s����@7bF�^���/���hf��;֬�Q��Z1g�q�k��(�B����� v=u��	���`���M�޻f�Ui��z�o����1�F�t{e�}Q5��]�q� ��i��3� �З%&��ݷ���%Mq��b��tO��#�ⱈ���'}(��7!&9 �f���-�I�{�[�K'}f�1��;|�[�cwյ!�:�?�똌��n
1�����_�Dx�(����q�ܰ��:,��'�F�7j]%:��X[2"lꬥ��w�j<�R�A�x�G|%=ۂ�M��i�Ϯvۂ�?(�l@O����-�l(3��*i<��^Fʓ�ުh):̇pĶOx��|M��lѡSM����B�Srծz6L�7y�iOU؛�O��/��ߓ�6� ��K	���V?_�Ж;���!�Ӧq�5�Gf���t��ٹ�H�� }��.����Mn����z�"�y�B\2�Q����
��yL�\�T��?�H�qD���w��HN�^]�K���{ѦD��b�c��X��J����K��� ��R*jZ�*5�JplE�������y5���,��H)%d���YiJe�SQd���|�6���ج��@�ZM�{�?��w\(k����ҵ8��)�����Yo,i�e����~3Sq�G�w+���u�D
�V��g��H����i&\��c&�Z]:� ��a���O��)a�A����g�~7�쟇����H�~�`�Y�@�s��:�"f�=�Ț�"FP?�Y�k�O)����s��2�+m�@}4��0��B&uj�&��T�'����5�CZ��I@���<Ѧk}f�Lw�WA��;s]�?$�}E1��J�+pB��J�L4���(�@����.���?(���J)��l�OUJ�*IS�;bq{�A	�u�3`3T�r<F�jp킃�e?=�~����ŭ���2t®�[)�#�dh�j�vHoW@/�b��`�`�(��Y ���7�vzs��ꡞ[N-e�)����'?�1��C1�䐃9��c,��5��������U��p��!�94/�8���x-a�m��RM�~��ِ~��Ze�(��q�)���ӕ�]H㕦�n�þF�u}/��j� ��*g�
��Yg� �^n)�.�����wpLH��|z��
��V���i�[���$�)3طÝj~60��fzu�9޸�@+w�\V�b��~����1ğ`�j=]CD&�AP�)�Ȩ�7��t��~��_�6�舣�����l�������X�nY�����䅌��}/3��n��r2Iz��%��aˢ�^��˪�X�P쨍��D:�8�.w
8���EN�?R���q �[��8�����l}3���N.�!D���P���5�p�SZ�n�.�GL@��̒��ށ��n��5y���ǒ��@}w.A��-�P�/4U[����<>yxa>���\��U~K0��c	���=����Kܤ���6�c����o6
�M���A�;��̸�@���;�ԗʀPR���(l|��Z���s���	&ڪ��rDH�l��T"�cY��f�2�nF�$�L�䮥	��/�= z6��i/7.˗Ωc4�V�������末���ӬH�{���+o���ضY��
1��塂��w��ȫ��!U�Wb�R��R<fl��:`4�r�0�h�[�!m/�.l�/"];����9> ���,�Key��p@�یP�~��XqgtG�;q��O�6���"�Fʨ�#f����4a@ `!������b� �wZ�U>�ŀ9�.�Nj���g/C�v_����Q�����B����B]��n�>=p\��9�t�~�=�4��<���� ӳ���{��7wOF�E��C7��H���Yi���K��Ơ�Mm"R��T�z{��V�:�`8�j��пH����ɑ�|��O&AT`��>ya�˳B��U��v�M�	��]�M�|��\+FW7�"��ALQ��[��a�xK0�������/�7���v��^�El��"j�<�UlO��N�~�Ejf�ة/��'i;�k���쿝l,��p�hN���i�E%d�
���E���C OO.Ia\��hG5�ͯ�4�t���j�?�kgZ<�'x{A�y�u\�U!�m�L���}��ᐊ�d	�Ru�*����S��u1�t��dC
�{)���x�w��ۯ̰�}�8a$ք�l��C�v
RTc�!��D�������=Ȧ%+Y�!RF�G`�P{���Ǽ��X�-o����{X�X��$�	��I(�Z1��0E��g�r�4��#�fY�@��YP��"�+ٴ!�� �O�i*#�>=�Q�bl�l��_(qS�Vz9ǳBH��- �b��Ir����	�U|x=G"O���Ӈ�a��`�yV"3���4�	��חO�K��[M��7��6ܵ��8�Go+ҿ/G�/E��_��� ���>�㓎"�9�oh��}�
��/�B��&��:*���)��0DӲ6��|�r���ʠ�"� �a��x:oW�)�,�&Kද�*���4)h%�f�M�#���M$���ռT�� �G�ꔳ��Va���%������@y��SDK�&D[/���[��.���;��i+���G,��Ҥ��1�qM�A,����&C���s��"���<ʹ���+��N��A�s2pL!<��^������~��2v�.�'��N�@�"N���0��2̰�0aA��Y�]�����1mY���Qy��p��hn)��S#vB������c�ŜS�r���y?6I1��[��J�d�j]����r���}�G-��I�������w)�G��-1�+a��!p�v���k�<Zބ믟S۱>������-�WS�`(!c��p�Yo��˷�M֢���+`�o)0L��z����%h+��)�xش�5ڋK�[I�W�ٴ��ݓ{=�c��,-�Vi���������-l1U�4��ЯZ�=�
���w�*�}I�U��I:���n�1�إ�b�����
q>��3.ŉ\;���P���O�?v�p�`����^���R-��B}b��6O�K�8���Ǻ˞��N�}���ؙh�yND�3@0�z[��-�k��槊'A��3�����(M	���=XAob:��N��MU,G�mZ�:Xat��rRg�+��F��jVaޚ;�$3hB������=\E��xM�g'B�?vO�Px��<ݞ{��|W���H��w�fg��[z�����ӎн��z���G�W���a`
�%'(�ꅢ��l��V��},	�*<8}ݕ�o1��v0^�8|����S#�pSh73��tR3��j	Q��x��*c��9z>�2�WU��C��z��V�X�t}^b��X��8��_	dL�;FH\t`"Y,r�	Z)e;k#!�됂)�
�*$���cV�%[2FztV��El��яB3�g��c2!͵pS%I|�(�{a��u�۽��"��|��BԚ#���#9��_�y	���}��`��x*	��wk�(�ʳ�$�������N�y&�Um,��(����?u��� l��ܖ:
�1�e,
�瘝G�7U�iQ�>�g�y[@�NP-���G��XeA+v�$@į��4���n��i�8c[��ޱHI�7H����S���D^d��KV�AYc܋<�� Jq�eVdJJTf�?>kf���jJ8���ɶ����O�I�oxEԿ�U��f*��$ޘ4����Tw��Ȣ�)牽'Z��V
��x���B������F���N錎��c�R�jQ��'�׽L�ӯ���IQ��]�"f{%g�N.u�y�$�Ȳ��2�-�@x�������P%�[�����4�E���s�(0~����mB�֩�G�����	A�0e�c�*oD���(噀�,���:�{},>����I��}]��T�w]W�����1ƒ�X��vF�XDϟ6�١�_7E�������C��l� L57�5�W���U]��xL/TR ����d=�R��O�ś
F���'^c���<d�b�®���wˬJA�b�+b�>#v
%��ie��#�_���߸����t:�Rg^>�<�*�z�ղ��?�B�Q�rq�;������ H���dj��8��bR��1fuSN!l��Lx���r�K%l��d�X��40Rρ��$�:������&�TF�|ì�~%�(��'���vQ��Ŀ����jk��+��yEٝ�@�ڋ��+�3o?-�0߾(��R��O��r�<+7C�������X������Oh���Z�H����Hb�)�-̏��i|�C��=$9���њ���l,o���v'��ݧqg:�ةr�f����Sm�� �A�
5c�E��mW�q�oڡ�I���ӪօN�P^4>x��':~<+��7��߁�7������W����u󤎄�.U6Em8�)TЗ�\ۡbH�QZ�?������-'�)���N���:xEQL�F�}��!{Q�kY����S�9�sł����d�a��V��0t
H;-�l|�S�ᇽڧpS������ ����m�i) ����l�Y��������)5� �����U��U�����d)QBc��U2�|Sw ����e��;�������y�D��L�1M*}U��fK�T���E��i�D[�_)�4��g�X���a�!�F���*&R���t
<�oF�p f�C��M���W�踙�R�%*bAp�si�c1�5&��h�z;���-�t�+�2��E�����7^�%Z�¼�D��+XO�����2�*����{p �Qm.ݐ��J�{��9ѭ[�Ӎ͔�Q����KA�mv�`sl���2X��2��W�O��[�
L\I�3DB0�:�ph|����oQ%	�̣���rD�zM���
�{e�]����"G��ʘ�f^>@����h�1UQ��g�6��9����u�i%���I5$�Wɶ��:�s*;`�a��bj���*-]�&�U�%�=����Y��>��^�S� ���b'2��?fl:<�1*��9T^fя$u0��q�_�=4��ncY$׾�u>0���	���0�P�*�d��AWڶCy.U��`
te��
�A"Pp��#_x^��U�5}{�zF�م����*5�&�ߟ��1�^ŀ����I{$j7�c״��$̕ښ8'���a,�Jq:MR���el0V�4%̏��-��6�r>3eZQ�%�t�'?P���'���߷�LREK�������LǴA�
)i2D�uJg���&,;I�6�_j8��l)�WO��"��<2���:��x�o*i�Y��r<�S��_D��b�7̆l5U�1Ngƕ�a�Ю�
��u�v��mUi�ZN`5�_�`��V������/	�e�𩇁�u.a�Qe�ܸ��X�j������B�p�kY0_���������ˆ��������v����_�ģ2�ȓ�"����oA���ƽ�6���hC)=  A-"��(�A>�e��I��f&��s��L��{�8�ݢF"W��l���k�.P�)�:i�8�8�͒�lj��������zꔑ^�������0��Li?�%N��#y[�j����ּ3����������-\1�1TX�`�.c�N�Oڒ��Gpn�_.�^ywo���$N����K��+&��n؅\�y�ǵ���3E�;C儱1d8"�^8P&����J��R�m�7Z��$����s~�����`/��7Ά�/����;4�ܦjl��il�J�h��Lg����	��i���zP�>i+��i��N�<i���3�	�&�c1�C>�a��0��"��x,���;�\8�hG��	�3�1BV��ɰ����ƌ�qpCx��y�0�m繱��i
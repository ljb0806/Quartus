��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X�D�(lQ9e-.?������������!F���O�ZU"�������Bu>�sa��Ҁ� ��uɸ���p}0�~]��è>Aܝ��i��|D"����1<l4�3	V�-(#���%��;=��p��;�BJ���W�8^/Z�0�8�#��9���QSK^oh0�x�$���\�1�E�J��H+Ds5n��:�bW:����:FNd^B����{df/O�����zcs���e�v�Nݮ`��\2xf�A�{��H�~ZѮ�ُ�,q���4'h����:�f�J�I���iC�]��P��`�4YG���̊�aYw�2����x�k��0���m���=|:��3���2|�y@�U��Q��/����eoԌ����v��3�����#��<Qa����A����'��\�(�Վ_����h�� O�Ծ;/��`��Gn���>��&��`�bA���8��rߡ��,`���������J��M�gk*�Z�e�L��>�*�R� ���l�t"�O�&��Ɓ!K�t��C�6�́ZA���^}���Gd4	|��4g
Ԣ/M����SF��VE�"�U��h������[F�� i[Ka�cE7f�gD��Ъ�<�i���ud�k���1rW���L��1��F�G���z)�]1�+�I&�*2��~�f_lev%�I�uO(iH�CL1=w�A�Ke���"�"D3�=�$et'G�D� ��/8�O�Α�L�SmU�	&����w�0���ZE?yqA����ا��Hl��4#V�;##�/�QӶ�#e�;�-�6��ϢG��]���/�3��	�s�H�%4]��7�Yd�����ؽ(�e!��&���8��^���$�"��ƅq�>CZ͎'���Z'����Ј[�R{;|��P5��R3�,���~�X���������ª���zcI9{�u�>6�e���mp�u��q�oB9���sS�uS��`�q�P*9�;�A����ï�q�~K hR.$��ޫ����ݖ���Q�]���O	k�ꘃ}��H|��;�������������X;7�4�=�Gf�����EKwR�G'��b���$bHm�B��Wd	�90w�
؈���%�A��3yx�F H�Q��߿������@��:-��Q�����ڌ7���[�Cc��.w�z�jd��$���싻�h1�o�F.N�]�%�^-*�cC��=��W�~]���4�� �	��\,�4c�c/�`�j#��rbܩu���}���]Yړ9�oe��fq�ӳ^�B�c��55.
����7��D3ب">��c�����]f�Zʉ�	�q�#S�i_�	�e�U�.����º�`�J��8�s��ͨ9�.Cra�>�(���l��He��S�T��~A���g�#�c��*Bꄡ�U�����H�/a��V�S����D0��֫T�a&�X�k�:h�9��
���'�3pxғI�P�j봞@$H��]�n��߈Y�N����a.Nɺ��d�A$�,%Fk�NޙO���Ds�U �#�M��y�9��և��T�dwTNGz$��f����6����c��O�Uj܊n�j9 �i&�Pͭqa�t&����2&���f��|ȺcN���E$��&'�k�ZF�ݖ���F�|�����xu9�+���<}��s����û�uc�t(��R�6M+���E��PX�B���)n��[���vAó�<�ɹ���,ط�ˡ���T!?�J�mZ8���fE���y������=˥�, �ZV�W?ۺ,*�|�#������Z�r��)�iUm�/7�N��I�g��Ov��e�HU�䣙��F�M��~i#�T'Lc|q���^��J�����s�w�L�N?��?=�ㇰ�j��Y_�2 �w-ak�5�=����7	�d����ۙQ� ��CPTʛ�#.T%�wP2��-���A�X�C^�G&���ठ8��¤@�@�;���p�i��Τ|��#��Y��G����PG���+iM���@)��5�& ��f*`IÁmzM�v��jO4VL�+iq8� j�<i<���Hg�!R�?y�鰈)�,��mBR{.�4nE��G�n�0���U?[�
UߺE��hc4L��%P�*埛\��\��ҍ|8Tz,��H=�n�3��MuS��=�7��A��j�oea¨=�n�9J�m*��M����n�ּ��W@��ϳ�B������(�rt��_-N��k�\�]^�KC2e��'(��~!���t�̯=�Q8����O��ىvR+�^�M���&������X_��A^������h=0K�I@(��2I�xI�ۀ��/�ݡj!�'�	�^L�N/r�B� P*�-t�d&ͷ ~hLi䫍����+VT.�[#�Z22��o	�~�ߔ)7r���]"�D���l5�!)��3[�爙��E���ƸA����CBYc�2E/�Om�#_U#����aQ�ø���Xyqc��{&�u��=�N�ڢ1���_�O�K�yBl��e\�h������t/�s%9S�"���x�������	�����}��*ky|���S��1���$ NY{#<潿��=ח⳶�Zj�T�(�=�=%����!��d^X2�]�Dt������ƹ��L.a�~� I}��;�Y��uu���R��'N	�����,xq�������2u����:L�
��_��~�3]�d�sʧci�'73�?1�P	�e��\(�\��ׯ���7P�{�k�]"��̖�U��%�bJ�Ȓ�Hڏ�ra����R�@2��D��������RB"�o�}�y�����2����w�l�(�3BV�	�rԾ��"����`�l|����:��
��|�4f���te�]������V}��0ȆBW�Z,Vj�n(��`�T�H�e��\�0:k�r�[�C���Y��ڇ��� �$|՟f:�.u*�2�<>#�z&N5f��o!Fl�*z�u�6���;T=w�Q*0T��u�m܁�X���o4$Bz���d��Y�g����&�S
��)C�m�4�Q��D�.���dj��:�+fet�-�6G����C�,6N�M�Zu��t jW&Gϰ/!2�����ߖ0#t�� ��k
�i]A�Ɇ��P�
5/K��#ǴDB��0Y$��pftxC�9�T�%g�o0B��YN�'n͘;��6�䧿��k�u���]�n�Ƚ[�%���Y�l��R�{�X�3Z�-$L��A7ЯA~Lk��b�q )���Ⱦ�՞����#������j�13-�H�[z��p�l0����	3����$�a+�����,ǩ�� �Ĳϗ��<R��")Y7�ɒ�1��9򲠏��d�]���E��hL9AO��%[<�C!G͇DN�VC���M+<_#f�����`���_�ѓ?F�����ʬ��VL�c�堗��g|�����9�8�0&A|�ݵ��3�]Ҩ-�r���zN�@}����&�ٶ}��f"�6��抄��`.��R��;��(��1�x�r���b���',T(��9)�����
b����.�&7���~�=��<�����B����Y>����]B���R_�sb6Pnݽb�(?�����1g�<*Cf���k�m(  XC]���C�׶Q]A�Vr�^���l�SH��`C4��L�j�x^D���G�'y˘�7�$�m�(��iHP�,Y��/�g qE��	{���<���%I�՘��Y��n�r�&Q��(�tYC�u�����%�`�3�mdloy%�c��g#��z
��/�/�Ri��V(ʹ&$�㭔��v��1I�ѩ�X�ި���
�A'�N�f �\�5��)�j����~�CE$.=W�ԨM�=�]�oa�X�`�v��	b�ĉ��o͊��wFX84���S���i��U�f��	�c���p�u?.Ҟ]}a�b��c?P�G|{|#�T�H���[�k͘+Y�&:/��,�Cd��ԉ���s91�n+rOt��ߗ��lT}�	��lK�dvr~�ځ�c/'����7t��?�	(�⯪ڑN �9�4;x�����b�� NК����`�P]Bj�TU⟕�Dm�����6�Y2V宧��W�Tz���ḞxŗCۼ�	����q����>��=��*K�Hjl|�&Fi�����U��ɉ��\Z�c0A�P�޷X=�ޭ��AkX�ې��Z���e������֜�*Ia�H�&Xe']l��$���9�����mɘ0�I�����	u��@��
��W�wR�-Wv��ei�jYׂ�٤�t���6�䬗P����A�����f�_�	�v����CA�j�Eedt��ľ᠚�$з����,pD�,�s\��������rN�r�DՃ��=}�l�M/=nS������G�܀B��`��=9���,�>(~�kЛs���AB��J�x<��G�b<lB�c\�0p�L�x�x��l�%)��q��[��`J��a�D{��K�V���ߑQ\��	�	N@�B1���wÕ7�+�mu�z�F������V��<�>�ݫ�
�I#���t��!>�*�?����@A����_��NBCT�m'/-���A���	�l�8��2����,������5��m��W[*���ɻ������W���t��gVA�8H�2���\�I���T���r˴�� l�JqQK,��_8*S�b�O���| B�O�ݠ`*7�J�q:@��x���61��ܨ�9���a�i�h������=��]j��1O;�l�?o���Q�%��<�@��8��O���R�ͤw�Z���m��ZQ�`���s���2Y�!tI�0�:"�奫�}�!��㸧�*���#�c��}&�.x��h|N�ᄲ'��/���٠��8�@"Hf��D!�_+ܶ 6�F	��qK�iWP��'/�"U̶�f��I���?¤�W��^�5�5��Ccyn"��gʋ��D��b���Q�6�{�_!�i<��N$
��m�	f{�e��.2��Y/��#1�@UtZdBWm�jǉu��V��)x|�)q�٬�Ȍ��eВ�r�6a	���jvL��mD�Q��ñٜ5:c��H�����kw͂�Qo_A�W��b$h"zɵY�_]�qvi1{Ҽ)7�^�>b��X���+"/.���E���n��^��L����ժ�����C%�m&(r}��^���
�ƭK%rD�BzI��B�7�����8Wy��f� �
��ԅ}6v��@�%��B��]��1��:sY�SM�0S8^�z�J�gsr;܍<��E9��rm��F���u�w;�H�o5�3��~#
����,v�S3A�T`�(q�(
pqW��¯B���.8S��" �P��T|ۉ����E�[;�V?��7��K��qg>/���]L,�8� ݩb/F���oэ1�ŏ0D�k�����U�J���-&�T�θ|���y�D
ClL��j�6]Ϝ��8�$q��@)���w/���6����{�j"��� ��
�V�ǙuR Ѷ� �n���5,LG�n�����Ϻ�BJj84���0�x^1�c|x���,��0��?��Ws�X���oܙ-��~+��e�^/`�Bg1�$@����F
&�a�5>��jY&�U0?�&��d�w�6�������ꖥ��iX:�(rxE�D��m|����~���G�w^�@���U厪RN�PՇ��Y7�ڛ�|�<u��)
V����p�>Q�z��������Mz���Rn��V)�;y`zO�hf�����Q����
*�p)����'R��ӵ\2vJ!=f���� l��G����!��7,����|�p�U.u�d�c4���q�y���.ԬD/�ׯ�e�zY��b[���3=$,��{��W���X�_�ת8k$�O���m<g���Y&����T�NBM���Ip) TY�EIM�����.gkb#Ye>"�)s�P�.�n��qFJ���b��\�f�Vqk�����a_�ʟ'Uw�S���3♣z�ٸ �`�,��n��v�0Eۯja.���%�`q�c�ɵ�j������Uz�H/)A�0�fȽaJ��M!����
E?ֆ� Q_�$�O�$�I6'Zo��4=s�UiUP��.:H��oy����n?G�ɶ�tr��^6W�
K�A3�sS\@�|X}�ǃUi��7��m������cW>L�щMJ���J��zH�}�zt��6rr��:��D�ڍZ�Z�dnGOf�s����n��2�I��9Z����)�Q|�*ş�*�:����,�^��;0o�hG;���Dd ������f'�Ȍ�f��M��q�h6a�FB��r݁�'&��h��ve2�vR'�>j1w����!�'=�*�`�Џ"F��K�f��l�"B{p���da�TA}<��k�mrQ?8�2�!Ș�J��@����29"�ܛO���ᰠ��wk�v��~�+����s���D7����j�r���jV2qדs"��,���}^)�I���p�Ձ��l���,IY��g{x�)w� c`	]h��+���������c�4n��X�?`> ۟��Z����c4�g���#\^2Z;���1Lj�ͧ���҅��5��}\��?�J�{6{q�ж��Ŕǒ��|�0A��V\�3�E�#p����^����{��lf ;΄���e�s��	6��1KG����7�W�N��o�q1����A����A���a�e��E�~���8���{��a3;�A��hVBˣ�����O��Zi���5��|�q�d�1�,� �a}�҅!�2b2�*3*�3��wS?��̴z�U�N�=���y�2���}pr�49�AV��VM%��;���������Oi��x"�ȧ7D�'sV���4��I��xb�TU��� 1�zʲ,-_P(w͠f��p�U !x[����%���H��Tֱ���GXb��-�;[2*:��9�h\ۃMձ����ȃQ��i�c�Pjs=�P=ze-̶� �o*n]�}�����'�Tc4��L^�h1��u^-��Z�/hq��q��h/4�)��<e({�0:.5H/Y2و���-硧ԓU�PA����<��BV1�G�)�9[�@�F��� Cvn��|�KW��0�I��:Q�œFWO�Oz�a�������@eeyLS4S��yͤ�n@p� ���w��t����,����Ş��]'&�j�?�9�pV_�I����&x3t���ҮvK�f$����׽/aoϭ$�o/��h��ڔ �
�fN�rb�3ޣ*+�FϷ�t'f��-�;yŝ#V�|�Qv�YZ�F��A�w�����c���+�ݷL>wj���M�k�[�'�&Z����L�P���hw&�ת�:�������
�A�Z���1�Z^��1(�[�`.�?��忀Lk&�=�e7��\�ڑH�u�g)����1e�yo���:#gT	і��R��x
���-���`�� �O"Z�I��ѿq,�����-���r�J�\��D!�NO~bd��Ϙ�(�w{ϺAa�˟�p�MQ�b?>��V�L�
[��f���"�<i��w�~]ĭ�c�'qĘR��4vٍ3a����|��=�B�h> �o&O��l����b{�K�sҢ����$e�~q۷_0dR��.4r3Ԩ/����u�Ć�1j�\̙�� O<�0�	~�>���@l%%@��n5^t@�G����ܳ�� �s������^/�Wz=��yO����K�	��	���
ūP)5�(�<�,*{m#`�e=筚n�/#���F��}��B푨�Ze}�p%�U��tFO`�4/�n���;��3�D��rM��<�k����"��J(X�@d��`k)�:�&C_��;fĴ�d�bҪ�9Ǧ��j��թҲ�#�#�9��.�ITdd�zm]feuq���Sdb_Sp&�{����$�
�}�*/�#������!�m-N%^�R�f�ϭN�P���*Hd>GQ����\��ؼR�Z	�r�J�;77��j��V?�� (S���5V<IЌ����]��L,�ԙ��w���0�^�My#C��vn;�릵b#:����w�~��9*V��7WY7x���$ʄbu�O�4����G���A�'ky~��^�k���^�����(��D��O���6�8cZ[?w��h��B¯b_>؄*[f#��SҖ���o��B�깙2�8	�95��}y����C'=M3�lL�t�ec�y��MB�a�"A�;�T�ɱM��~80�
����� �'P�RA�#rF��[^�3������H��&%fm�&�1�&sQ����i�c����_ӧ�F��]��M%�3��z�����|��SQ�A�E9�-�Dz�F�C�ꨒ)f;<��<BJMѬ��/ng���d��9Ԍ$�X���SGQ�U�%��kP��uқ���z����:sO�����2��,��u*j�<���t����WgG�;��f�Vq�����N�g�bt����sDƻM�����)c�)�j��z�5����k�X�謻"/�m����)-�Yb���g��.kk�x_�G��t��Jb�n�^����r�@]��ݥJZ�t�ɩFH�#+F��L����p����A0@��9�D`����;���*\ۂ���ra��=Iw�oS�&���qū�#q���g~h���e��)�뙌�.A]���AZO6�SZ���퉪ZjW�Y��zG.u;�� �J9��"��ʆ��VА�sj�C.M�j����$�6��TP�C���%����}�x^��&��/z�w�n`�t�7vE$�&X�-�qǹ����z�N)4g���~��
2�{��\��Gu��x��Cpr�'kRA����$�.���n�V>Z�=�N~
&�Td��s��"Y��]���!!�V=}��IR�S1��4��D�L��.{��%�&^��@�QL(��,9�s�T�=h�
�wj@��ǴQ���� p�J1ϫ@^N��a�n�8� ���ɋ��0�tQo&�Nˢmo5EZ�XU��;7�|j�u�r�F�{���dGF?p�(�+���
�����<�@��^
F�%�q�AB��ݺ˱��H�ʆ��쇗�i���Ȼ��������x��n����K5g�c-�ݤi�O!�՞U�ski�C��\kQ3��Ė���X/��� �	�t.�a<��JC�]����	��~�+p�v�<urf���6m{)�TY�_���S��n�2/&^K��G��HK}���]O=8bl[�Ϫjj�:�[#��0h��}���l �s�%��A�lJ$Jrx����jKA����X'�@���a18�r������'����C�`�>T��R`D�4�&#���Y�t1��[m ո�0r�o?�Ѵba�X);�A��$C��U�^Vq���T���2���Q�	�.�3�K)@T�Ef/jOZ/�Δ���P|]֘�]η��>�K?o�s/bg�dL��$r�f�wr2ws�+Fn����O�O�w��J6��i��B+��w:6�����u$�����qR'�e�B�hf@��[��7�����hKd ��ZPt%��%�Dd�@ި]T���o���_��Z|6IAOgt��8��|_�fؓ�-�	�L��QE���-��ʜ743�(�����#�N/�5�a�tcx����(�z��PX�pk��������������d��/넫�2r�c�(��<�9�ڳu�
l䖀��&[��)r:�g�F���B3q3OJ3�����u��#i|�&�l�)�l��؉��݆��+\ںVF|N��w1aą�{m� g��-L{���T��9~S������D#/?|�<���4d����L�O��׉�<�[��J�p#�G��I�k�noX�7��Y��$��tv
��_>5w�泯�=1��g�nAJ[�]����T2�5��a�����
ۡ舒�6E ��g�������V���o]�Sd��I�lM�x0�
OdŘesʿ�w��<F'T��(�9�sK~���2�34!l�+�&��c�3��@��o��˕3��D����#�uO	�϶�����$K�5xak/���9�3b��C{��
����?�L���*Rp����j	��!��f��!�3RD����!_>���(w�ʚ^��4��j%�0(����
��OVVL-���y7Sw�Z��'l@c�I1SW�5������ɓ�튴^]��=��i��b���y�v AدRr�ץ���lf(����>�92�R�&n���*#���
ƨ��#ы)g��G]v]z�ކF,v���zP���	�|˞X� %�vF�b{N2�!�k/ɬƓp�Yy��,�]u�<~)��ϑ0�i�����]��:����B<8��*�`��p6�.:�^u�g�`�8QI�*�Rt#��+NҾU~@�����������>^���s�`'A��ۭ����a�PG!;Og"{��&�d*%���}��}?.�r�'�#���)��I�8��hu6 ��}#�i��0qw�&si9���Z5�2S�+�p����w�ʃ�@C������'6��'����[��s���&���"�����V�<kT~/�R<��_Tn7����(r;�pY�/���,�<pR���@v��Ȥ$ޭ��|ߍ�����0����01�1���+�終�V<�[��=�y�Lb�k�77������ˉ������~��Zd�c��r�������	T��lOU��Y���@��C��^�ING���
���M(��QP����>�'4���J�OL-��pE=:�ŞMe,|^c�u�
.gt>d�=���5_�����O�?Qz����+���'�w���+�JU��Pm��ڼ>h=%�A��#�H2���Z��C�������B�˫���]�W��]��� ��Zp�m)�)�/e�p�aQ�t����К��H�Ӽģ'�w(�A-q -�[����^���C��>�~�i��m��L]�m��N�n)��J"X�`��"�pR̦�ɠ�E�������_��"�*��-�h��6�z�@�Zl����B�!���ݑZPq�H
�릾O�ԇL,;��}×~I�E�}kI�{��si��$�.������_J���e�ͻ�_ς��z��ف���eU���V�������qwn� �����B�~�>����:��-��h�Rf_V��:�7��١��h��Ft�rh�T�I�`��JZ��C+0"}`� ӱQ�2�E�� �K�|e3�;6s�+����n����ƛ�w����U-�
̟���Z���g��Zr��{$,q �OS�T ���z^1uJ	����l�B��A�+:��6;)b��yՑ�x�2g�q�c�4O�dC�	��s}�kV���?U�[
w�3��.�Aa����W�Y=�;E�ƈ����)�BN+�m�᭦m"D����Bd�ݸ"_")���¼�(���޾0�%��+/�:�[ �=�D&��0	��ћ�|䋏���Ŋ��Safcrl�מ������c<ԏj�;���>xԽ�b�-��xG�j��热�8F)�-����3[��Άc\��K(Uߔ�+�/�N���h��	�X��0(=�iz��"z�5�m��X]'3������Ro:�n��!��  ~���`^���q6��)剳�˗0#A����z5���)��a��v�Vg]�! ��CgָĢ&� {����Z�MN�ɽ�˞�A���
��}�{���7Q��X2s���@��I�_t��d���E.�j�DBT��?%����F�H��8�y>j��Q��@ɥ2�(GN�45t�U�-o���840g:�C��4�Œ	�f�}��80�F���_ ��P޷���A�ҬՆ����ehy~�N�����)��e����B/��s���B���uE�G{�H�Q���,wwCub�
��|ݯ�Oo�<f���{����-�I7S
ܢ��TbX�Y+�!�j��w O(�Ͳy����H(�o�X�4D`ڞ��
�nN3�n�hJN�PB�Z'���qk}������@������mf�0�lb�V���Y�!a�U+3��j�BM[����ś;�oE���7�"C��Ӵ�8ѫM�bN�h����׺M������kzm�
:�w�9]�)���(�r]�Z��Mˀ����:֣^&=���t��p��㊡2�/ڃ�qI�d��׉Cb�3n��(tf�6(�^���Ci����W��>��J?��H|�O?�mA�ۥ�(�E�=��ؤ�u.Y��$�?��C��̯N`�r�����˂Z�X���T��#�p̘�<��4��pk>�^��u.:���@���2�s�g�t�t"\1P�ߠ�(��}�?���8ഌSc��K0z��,�cL>��#+
J����� �Ŧ*S��v���vE��d���iEk�����{Ŷ	�6�����)rK��'V��
�]f�
_ �����
������"h�O4q�U�!���e���a�?��D���.�ی[<gf��RC?���]l�I,�K7$�ԁ6G�M ���Hh3(�-`Z�9���+��^���n��Y�g�����H9��s�C�����$Y�h�t�W��'��F❗�ӕ�rߜ6rq8W�**�G�[��/o�5���8K��JX'k�V��v5>�Q(��汘���G}��u��#����>�g}?��8�uύ��CO�4w��o�R�W�f��cd�d���rB�"���������ϡ<���0t�	�,�秝�j�K�N��	��ze+{�� �u������ϋ��#y+ e�q�����p�7���:P;E��X;���>�j���I@��.*n��\�l~A3Y�;���ɼ$σ�T;Q��,~��ф/��6Mb�y���C�"q����flv+�5�:N�F�ڏiC���a�X�E�l��0{��+�Y�
�/q�����\�zd�捠%��)w=d�7�O�F�N[S&�g�F��
	�j�ސ]��"u�"����/g~F���{�&�~�� �7������Pr&��?���M"}�����"���Z��*P+��r�f�6G�(๜f	\�0��k�sD;w���|����5���ڡ�?�#���P����ǌ\v�w�+`�7�q�V���/����N�XV���X�̄�:�U�6����-#a3p���l.a�מaZ�e�F�$_eSsx{��)5?Z�,{+���h��A֙�7�����?�Y�޵����WRG�-�U�ܺy`uΈ�	�<���l[3�Ih�޾�@��v:�3�6�R�n�[���������fA��;�Uo��{�VZ�7�rI�2G�Qk��(Y��x���q�w�����)Θu�ݼ�����d���KLc�4�
��a9�T;����51"��-��	-W�@�%�RYX3r��:EVᰀ���B\Z5�?�T��{9�f/�2rȔ�msV~	����xeD'�L����3�'<Їp�ԛ:r���-{�[�Ux�3�'��؄�QZ��4�Μy�����?�U�Zg�?#��3�f��,�m����2$¢�����j��ٲ`2�j����|U��]�5#D}�A�*v��0�Crp}-�z��`���`��1���{e� մ�΀�W遣d���\|*�k:�`ɥ!�Boiʘt*�gl������&0�0��/��n��p���N���Ѥ⟈ⱀ���֪�F���@�O-W�)ܢ;IM���C�I�m�V��O{r<pz���-*3|��O���^5����9�U����O&�JE<$f1Ia\�&�3��̼w�˭["��M٣�h��]EO�0�s���\��?�B�j�R+.��T�齢c�X���>mӎN6M���J& (QE���l��Ҩ�,��݀P�Ȧs�a!��L�P��8�,��ۂoB�ɗQ��*��׀��sКЖg��M���B�|Yo�8<V�����4�U�ڨ�M�%MM����Y�Q�ӄ���ᚐ1Dū)�,? �O|�91�5=&&���S���	�߳�q��� �B�k������@/�����q�xZG!|�R����<Nu��� ����5��7���USI�ޖQ׌J� ������O��!D��g���
k�f��_�6��\��P��9q��L�+�ʤ��1�Tn��L���z3������;�SN�:�U�Q�)sԨ>y��V�u�r�A Hna�����}�Vz�B�����S�[P�V?�}͝���ؕ��Qd�~���;��TQY=Ӫ-�FJ!,��gdK7�� �T�F��+�@��N0���~�!6�m�F�U�����tF`N��8֓��1	$�ͷ�<�.hµ^a��i���u���aD��v�j�[�T�~rr�P3O��]�􄩰�3�w5X2�pa9����X���(�bj�۾�F�C�p�}d�Uh���J���㌌����%+�{���I̳�� ������Ab�h��Ή�����'�gn;�9�����B`�ſr4��W�2v}��rO%�Uj�-�� +pt�S=B�F<�9�c
��+уGu��H��<u�(B!��W�J�B��H����7ge�*�.7x(6����E�oA3�y}a��L$���P$j��7) ����d�B�r���]�/�^�|s�y��Y.Xl��P���to8T���>;@"ir�P�`G����)�G[5
���1��d������+��מ��ǯIכJz�rQ���0��z���Yڎ�P�=�6���k��t��K�(� �4�g��M���m~���Fմ��@�ֹXp�u�nJ��˺����\T�3�V���{U�M\��ԯ���I�xI��˺73n}"*��W@C(Y��~}]z��
��`�%�h	�3 ��0呩 N��]-o��/0M��aA�D��>@�A�Bn/�y�"	�|�4���:]J�������[���?R�
@��i$�C�ѢN�j��Ƹ�x���ptn�:nŴ�P���"ɶ��-uM4��"P�VyW��$E�5b�O	�/�;.߄����5��'����j�q�-ʩ��x;�=/ϊ*�sÕ��w3�yy^��P�[�jФ�Q�`��xn����Ai2��j�Ԕ=�+4n�]����!q#*�^p��ࠃ�A+[��%�J�b�1����|=���#"���Qg���C���I��af^�3J�/��7l�d�R����Z�п(���d��Ԋ����s�?�8B �,�����7�K�n@�a��G��z4�\�8[��P����j�9�H%l�C���5!0f+�?�HL/�#�P�Y��y�!(ě�`�Y,M�0��� �+�]��S��XnL:b�ޚi�ُ������j���L�үn�3���4�L�z?
��!�'~M����a��E(Z*X�n�,����1Dr�ֳwܯ�|����B_����&n���fL�f�,hV�-��%�@I����mg��5��J�S�>{����m;~��w�ކZ<x�Hqڅ����B�)��(aȺ���E�7�8�vi���-�=~��@�ZN�/�df�n��>����PB+����l
��D��[����H�5oH8Q�D�S��mx���"��ib����g��$0���퐤��=D!;�g����yض�#�O�)�0��cR�e	�?�Rh�'�N�}��tÔ�wu�Wg�WD;�c��3;�Y�,�)��&���������S�(�|>&P|/�`[T������6ر�^�Bq�p�xE���	q��]gq�L����y���`Dg��)�w���I4»��e'�W��Q����'zD��"W�j��7J���n�+p�fH�띘n��
���B+r�V�������k�8��b����+���C���k�����ǈ?�V
`R:	��E� �wZ�����	~��s�g}x"��?>�c�#�z�����+o�5	>���NMO-���Er1f�/y�S].F)�����4M�%���&I����?}	i�/��_��:cd�8U�h���q�AR���TS�������3�Ej#���,vܫ*y/�ǥ*�qI��դxD����JIyɪ��1ܱ3ep�a�&�`�^Id�����]��@A�С���Z���9�\�R*?d�=����3�A'۩��b˩�4h�9����XU!����_YtyP�_&e�!�6Zg�)�.��㈃EۢpSQb~*Sk3�z��Z����!Ԥ= |K��D�rS_^����9zd	{���[HF�r[-�4�V��w��4��K���'!�ao-@���?�fV�K�������Ѭ��F�1;Y��
��u�DT������V6!��#B�u3�K�JK;ZLƬ�Xh���D� H�{��\�%�Y'S�}��{҃�j+�US�`����w�AY�`u�o3�=�
�;E�t�Ν ǰ?���݅��JD�ȼ'�4�7V 4!΁I�¢[g���%`md����������)&*���%٣fID�'��uO��ݞA�ɶ-L��)�/�Rx���8�uH!�3S��y,+��&�r�z��1hB6ɚ<2rp��]���F��5v�{h�����xs���Ɋ&/�p��Iگ)N���=+�`%HRƶ�$��r�� `!�Pu���@����.�3�3���÷���"鿲t���r��	�y$R���d̔�.<�v���I&6K˒��:������}�Uc��x�4n|�U��Zv0��$W~��D׌���A]#���P���
1�Q�H�Ϋ��t��N����0N]�K�	����74
$�����N�3�h�6ۺ�)�C-&7���,g�C�f��?��O�~ j"�h�x�	��]�I��P$�h��t�)��-� B�%X��݊��Ep3��j��(� (��(Ǥ���d2nLce��U�/���C�w��9�|iH�{����l~q�R-!�N������;�FP��oc��L<���[���j��4����L6~�}��	غ�I�ۙ�d�08�p��o�@����
�i(��jM����D�>����'��ώ ��C�;��X;�f�`���JFtqq�Bڜs�/���-
��暪�@PR��Ü4+]�,�ee�ˣn	WR�5��+6�;\�&U^��](Ҩ�px�լ?�:b}M6ED�B�ګ�=�6�F�����9�����<���!�Fm�y����d��[]i��԰P봭k̈hY-X
��t�X�+�?rđ�s8Y�XrC��Y�����T�+a�ky�)I�~��� ��.��=�L�"��`%�ەM������0�$��htY]���Ё������FI���$�\�n[��oƔ���a�S㔬�w���g=;�ī�<R/���W�w)l:��=6a�c"�K�Y��T4�!�.N�����JaL1��b�#�aD8���hS����S�L�P(U3����T؅ q��'�V��S�ܺ.�����ßB�f�!��X�;+֭��|	@yI'��H�s�#����7���z3� ��u"4(��u�D~S�T�7�Lw�l��w��#?��G�rc�a�E��.oYS�/k!`в���X��6�� ߇�$���\@�iWӁ^�<���#�n��l0�'B�AY"����iuA<�����]0�\Zj�*(��п���T�HՓ�j��;}�NS���ݍ�	���9�����j��5���3���R�sn@%�KFGW2�ja=}n��-[���{ ����F:󣀘d�=��X?DJ���:�\��}n�USkj
CR�b���e��ӎ�k*	a9�����UG����/�X�_�Mf�Grșy��a5M�֜o
�W��d$j�W��m�H=Ǝ�����szm	`�����á���"��Б��q2}'��͋�?+T$��o�E��������=��D䷌m� �sf�y]�yc|����>��	}N����V�b3Bl�U)"CQ<��Ps���%��'F
�I�Hޟd��V!�{������
���y�ˍW�{�*r�>��mB�'{.�f,*��_�N����at�e4 �wrD�'�E���k2��>�2w`���h�������2�o1�ɣ�<�g��ǳ���e
ʲx/���A�&�Q�4M<�+��@�Ss3�n��D�Bf�E ���k\��4Ęȍ��fe�!U�+���d��WJUn�\D�@f�}����^~ )x{1�W>�*���1�(j�s�T���‐��G-ܓ����2�ˇ �݈��XA*	&���`pL&ʄ���\��o���l�c�r&(\��/RzA��)�p������Hc".ة���Z�? k:�-p�������`�G���$�'�k+��]�"��M�F��$�-r���C��K�6������m�GD%�4��P-
U����i՟������D�[ WJ�t�,�eBA�k��=vh��IM(բ�p�~��y�G�޸�4�\H����{�B�����CvI�.��q��jG�����96�'@�r])�C�2"չ���jQ�u�4zs~xgȞ��^w�3��.O� �bl�
�q�*����̺C��>���3��NQ96 ��(q���vo�Z:f�:z��s�Y��q�鋌Hy��X9:s��|R���B-(  ��t�f�����F�c5�H� 	ﰹ�3LJ���b�۶��˝��x��,#�'S*��I9�Օt7����F��l֫�<l�T9��74^�Q���k��Sݭ�+���<����|�٧��tPi�ۨ��2CD��6���~����Z��;���A�R=]���2MP������hsd�y��^�_�r��~��z>I�W������6��dDr0��r	5 ��`!į
.O#�j�-�8��h�� �1R�ݭ�@����g$���n�)��e�)hÎ����XMK�nb�����4U��,=R؉׬��U}ǆ�h\k�>f���]���M0�VI�:��*u�����;�+n���t�[�
>@��/l�)
�VF��tʨu���*��U�ʫ�T�� ��������c��mjjF�9'�.^t��17��fj��bR����G��N��I�2f���x�?�.���O�A1��Ǹ6B����y�o�1���t�d�ŦY�vP��i�S;�4R�<j����`� ��8��6�G6������n���{uX��|�Q��g�~��#�� �"K����'�D������x��������q�Т���o��^�!��#ؘvPGv�~@�]��b� ���}�F�0?=���|��D�G�e�_j�"�_������Ư�3a�M�����
�N�'�/��͑8-O�@I�n8mɌ�-O�=i"�{���IC��h;o��o�7;�M �@�=Y�): �3�)ZS�6�V�,�[���rwT�z�X Fu�WZ���MweV�	���нEݮ\����b׊��Ҁ[��(�{��#ܛ8a�z�j=Ŧ!}��@oƵ�Ya.�,.8���	3�+������^��8�����vS��C��L'��X+�2:��v���v�}goylD4�)��8����:����7�Q����p�����C�(��7C�`8��ω�"�v�`��rt�_.��,L���C�T�ȫz�k�,����
�T=Va��#I;�1���=���}�^o�ńu�E|��١��C�?IKpn�&�]�+.Ӳ�t��-3iQ֔&�{��/�5^��?�Pf�n��R�j��B�K/��^s����~��)x�x<.��FAB&�>5Ѫ�L�,2��3�����$�
T���;'��wh��L��Pԫ>B��!���>�џ��Ι�?�P����Fo�@���Z��W�P�R5*e;gȇ�p��
��1|B ��^�U��5R<�7��Β���7G��׬^���q�|j�!���������g{�>`v��
���/=b`�q����<gSm��y��Mp�[ikTE��t�	��-�{[̄�	��[-�t�k4uen�CzK���e�$Aƃ��٥� t �x�vc�9���� ��r�o4@҂�1=Zn���6����Q�:�hP�iy��c�)��߬P0��S���I�08ih����%���\�҉P�Xȟj�	�b�A��l�/5bBB��㤎&O)��/Nn�e#�zN�)gk<��\5��������=�VY�<��?�}D }�"XP���wY-��h���u�]_;�X�SmbE��{��M2_��9[�]z�ג3�#����;�v]/���l���G�+��ك���<��ch�{#p�^V��*�����w�Ьڎ=�@�n�<j�`P9��˖WdEv�Z�Ԝ5�4/v!��ǳ]�C���k���x~�oLf�R�$Y��Z@�8W�JXq��R�Q٧�/�!��v������wg߷} �,�UvƯ������ն��D�B�t�Yz��FsY�H���Y�`�3�i}u��1h���� g�:��m�),��'�̱|T9Ret��m�1I P#����OE��-�Z9�*�w|y�?�C��r௢��ef���Ug�,�.���1I�v���.9�6��18�4����Y-�Y��tUH%��t��.p��Umd:πJ���,#ǘ�����ʌ��̐�Dw:~r�<&��vj�:[6dɢ����ԃ(���1�@�m.��x�|`7�	O�7�ռ5�V�mL_�@���P%�;�<*c;m�jRHH��-�0����NA�>���_ԁ��$����ǵ�Ĭ،N5�]�B}xa˟�3luh,�8M�c�R`?$����y߫����X����I)A}�K��"f<��
Ue��Zp�}����k*�p{?3��7L�� ���%�[qܵ�,3��e���)�E�c�tV]"]H[�������� ;D���wn�O^��r��2V�i�'���YF��+<�P����g�]�d��;��GW.��]6Nyf�R����˚�oL\S}�0�%5��~m4�h��(���ܑ�-��2�X�"�YHE`��S튉�+�c��֧4��^H=��ѱ�>y|,"c�/�5պ4�@��u2����� ���v�
4g��[�`u�Z �O��(}ܠ~�.$�z�����Ċ�^	-�u�5�;6��'��޼��9��4͍P���1��n�w&M�[bf�'�*��O��<N#_�ax�Ț�����>\G�{�P뫇�<�Z��&cUԠ���	��/r�[�%��`���u�p����T�x?	�KMC	��&��o�����^��0�CS�����DfC̈;�I�d�b�zϩc�΋�Y�� O��#?Z���P��t�n|�w��AL�pv�miN�R��M�w�`�+�1
������*b��^���;�c�b{�,���Q�]i������2o9�2��\���ζg �Y�����HWs�υ�c�pP��$g�����Ņc�!��/"�z�5� ���P��|�x׆�6l{q��g�@����R�!��}�Y�Ss;g�$l�I+k���쪘�9�9�]�ݦ�z}V�^>hiWGzcg���B4�7Y!䀦Fּ��JLI'���e/r�`W/�#�s0�(vm)W��"N�:�֝�Ce�����) �S�t����	��Y������m=�A��x��!�7�ś��\������SS�4���wRw���y����j`ɿ��Hk-���h�?J�` �����<g���F*~E.j�0�Q-��l�%��N쫴NI���&���r�74�"��!WH/ܻM雃�1sq�򯜥��|���$�w��'%��$%h�#q�M�����A������(�]*��V��J�[k#��]1>���֮o�5&�+@$���W��|a�= ����8��]��c�閴8$�H�����Qx�7��zJ{<K��xe��:�t 03�)t�b�OV�#Ǜί���Q���N��v�P�@��gY� ��B;s>'рg���ȶ��d^	�'V�	6*8	�J;_i��(�lW�����؝S�M�[b�C���T��_F��ws6�(����EN�q�N�Zj
r�~��:8�b��fezk��"z+a�85�ǜ�:쥷Z ������=�(�.�HeY�2z�WX;:���VO� k�����՗��}嘒�����P6�M���
:jg�7����NP$䣰�`�^VqX�5����f�$��e�	�ze�w��� �3I�y^�[���~MWd
_�&�|5��#-�ߞ���Z�~Sz����O�����`��4���]�f�V�������9�4�P����\OӋ��[�\�@zL�58[����F-�13H}���Ph r!�����Ě����������\���X8T�t��۸��	᱾�W�4;7bq�<j�3�,�w��V���5j :*��Y���W�5����\��Z���r����ZD��O�X��Qtw���}<�X��Zt*VM������]�I:~=���:�S�	��^���p]��M�����7@s�%{��"e��1�&��ݒ�w��;�9��[_��L��o�0K(l�26��m�3�c1,�X$e����v{ؕH'P_S1����O}�jO���/�U@{X���0J);tv�c����j'�yLޙHK��ٿhe��-�ݲ����b�wU&�Ns�ykuqɁr�ģ8��T��� &;�Vx!S���ŻW;���\9:��H���;��g��H�P�
R<�U���[{�*�S@�lr��t�#�2:1�%�3�-`w�J���+�dE����~@A�v oL��E�0�ݗVlr;�h��	�(�:=��'l��y��Mn���/ˆ	)��mbiI�
�9v�S�9�}�	^��b~�|;R��0���7a��\J�Z6n���%Zx�
`D8g��$��='`؇9_/��%N�e�tw��=N;승/�h�9�y��i[�/z/�!i�n�D�M@��E�%�d�4�gW<�{�i@���B}"��۵���߷) ���3w5��"��D��0Ѵ�Itp9���2���-���U���'t]����=*ƿ٭���h��B╹���?CO�|v�4f�CI{(]�=�PT��@`�Y��M�zr3v�o�2ߓ�AF``���)R��-����ݱ�B�����cm)�ͤ���� �۸B��yA�<%�7
9	�RVUl������,2�X�Om)e��=6�N��`�)��>���{�J�K���g����I�[}̂0������.D�-�E�=�0&X��J�/p�Y�@C�u�}oYOg-��Q2�Oc�N�i�̷7A�6�u�E���Y#@2�r� �4K��<c�n���L �(@W���p��l�D1v焑�Y	-Y	 �d]���5�`��=��L�%���.
˪7������nE��t�a���d��V�C��ѫH�����{��[�7�f�i�"���L\U�/t��O4';��
������U��;5�zn�
�1.(2auTq��1���I_�_R�o�Ұ��S��NvEX���,vJ@�����Kk;D����`�G�l�{����v�r�JZI�[���N8BL�� ��.�b|��r? �f>uV��C��J�M���Cl��)� ܱ�������س嬍�=ͪ���Mm��K[9s���
Ώ ���Ûl�!;�]gKH4V���\_�v,;���ۤ�
�l'�^��y��5��䫙޻6� $k�B��d|�	�Fk,��c>��6
�T�؆Y}\^B�9�W������⾧ne���r�����|"���=_ҩ�+ɶ�?�r�W;֣ꟲ0�"���L�n�)�he��Omϼ�{~@���P0� U޺)A�^�"��<v�'�e�o��ZG����S�+���3E�r�.�a��R��������2h��+)�|��Y���I-��Js�Z���kZb� }"3y �&�V/�8e4z\r�Z�$@�|�XM2�KW:P_�*�g�����6/
���0���:d
��@�0pm���e�oq���wӻ���ێg�6乨y`h%Fgt����l۵��?��+�+��J2C������4���[��+�P�;W�(򆿹�8�;��&��٦���N�J���4<a��"煻?��D�ʊFΎ���QSX�<����5��O��,���!����4�	U�����N8��1�$��&��z���d�(��=�����L��&��`B����m:Ǻ�!԰�-_�nD��Æ�I�'�����ط7�m�
�I���v!���ڣ @�%���g��.�0-R�dx�:h�e0T��`C�+%GS'v-�q�{i8�w��
D��:�U�Aly�oY������}��8��A�[�M��w��8�o�z�+�OaD�b.:�~+�1!4�%Gw6ܓ9畴�**��J7���.��2.ě�N�c��3��)���C�Ѐ�
�j�0?�`�c��಍�6�5�%��il�V��U&AG0���DheJ�1�~qp-\��e�n�(�*��d�!a_Ѽ2�4O�$ =�,����*dm�o�zm�n��X�R�d��5��N���'a�ߌ��B�,�Y���$-��o��e�/y�K��E! Nd�u�yI(�^��x#�KuܞO;OIR� ��l�|�d�����������K�n1�hܖ�Xk{�
�Z����V7�(fr�~�^b�I!j�c#f�d�eͿK��0�N��	�H`d����{PK�s�t���)��6�=y��q��Y� \k�U�`5e �>�R�`�K�7��E�� /�~f�r-�{<�v�|�a]�%�ò�q���M�#o.�*���U��4��T�X���#Q7�S�@�Xb4��I�&�����5��Kj*��,��`��X�CF|�=�r6j��;o#�b��	��5�8-�#n�;�zG����-� �;;���.ߴLR^��$ʷ6�@�5P���&T��뻱�Q�l��mU��V�rsz��l�k�ct�.0F��w5��a����PLS���J�#�j{e����"�ҳد�*gy��tcX�X29W42@�6�c�5�ʾy�F�x�)_� ��F3�-��!@��z'�����9���gҢH�v�w�r��\!4~	BWX)��n(W.�D�Vy����s�n��rýZ�����gA3�"�Hw�^�Ĥ�c&�sN8���}�T����TA��9����rZѿ#��D��g�B{U�u��L5)�|*.m�fW��-��+jS߶�����s�4-&�׳4���pו�U>@o�c:�(7U��1�]�z���	f7�i(�1vD_̻�����b�P��3g��Q&��OZ�V䳘r�����}���cZ��_fٳe�$�0�bcs�⤽XQ��<"�\�<���c���h,x$e����=���x͖Q������Y�����b�pF#�f�xa�ʼ�wOo�"t�Ӓ�H�@\����K�ɠ��B��9��M�Ԇ�X՛���L��ϻ�$c�p�s0��K�3H8�#��Xsw��Dg�ް�O�e/���N���n�_Oئ�I]db�Ռ��i-9{�ᗪU8/�z3_��R�D�!�4]'4r�� o!:�U���h��+{�t�̰lX�Ϛp�=�L)_4�m���JpڂP�E��7:,k�M��Z�df�����_�t��?A���f[����@O5k�$)���w���Oz{�3q�#l��N<Ȃ)�f��3`;ٚg{�Â��d1w�D��.E���GO����N�%!��\�\S��I�7������(��g> ��I�ΆҩkFS��s�m5+���=��)�G6�z��g5}�儂t�}Z�Cm?^�.�͠u�E���4p�Xj���M�.���8��e�X2�G��茧g� ���k�A}Ŵ(!J̕�d�i�8\y��ʳ���;�����&RȎ>�����E1Gn��n#S�����8Id�~��f��눨�T.�D�^�9�u:�
��;��2�<e�n=�k9�O�.��.ڛe� �^M�����=k�~�B��!Ee��h٬�jܬ��=�ht��¶���h8+��NP��q4Ű]����-��@� K.�N��R˰�8��<�1�p�(�wѭ% 7h��i?U>:?�.H6lq`��;��j��H�^Fq�v吃�+��ى"�~ي��1i�7�K���������a��R�{(��:�1As���^�M=9�"�|ky:��;��m����+�i�j+�<O����Y�G����-�%�į-��� �7��@O���Qa�d��
���<},�yկ}p���ͣ�5-�����eKqN"ƿk�M���6���n�î����T6�b�k��	&�`�e_��>%�.�7�"���{�e�fBY4qI����w7 �����`:Zn%��&m���9��5�7=��Zf�lO��+l��SU۸F�����Gv^��;	�]��t�>�Z�##��7��h�m��#�j�2��JdW��ٮ���F;pv/�S�֋�`���9���P~�B3�}��ٚ�ʥ��.�3��)��V>*qƐ�V�ձ����=&h�6Rg�cAn��<��D�z���n��A����7�B*�BXo\6���$�kHΧr���2]�W�������."c�@����P\�4�#��|+�~8��X�����o�g:ö�=6P�g����\�\�o�X;����SIa2�݋���U3��wdr��tF����;��k&�^8!�R��VSZ�~�Zi��jt	O�$v�uL/�5�VpYF�?��e����ŋ�u����\����p��V�=���(�G��I�ݯ��Nh�7��%ׅ�O@�}��[��Je�N:�g�q��$MqL�q;�j�տ��y����'{���a��{���DKzQ�z/Q�7���lӆ�/�����8�-z��sǢ���cI㰖#Y�4XTAB���F��Y�,������d+c�p'����L��!i����֢��}���ZW��K���A�ś���7�2G�
ju~�e[��e���wo��+b(�0��x�HsD(�h��|�'Ni�2�Xc��
�Eo�����']��$&�� oF��}���@	B9`�d��&LAR{Ӿ#�؏�P�q���)6�_�&����%�'��J.���H'vP���Yl���?�|�W���<����=�m�����,�u[8�ol��i1�~pr|���f��%D|��&����ś��)|!�;��kif��j;�5�e�$��\M�dL�%XYs �B��f���	��7+�a�i[;�қ�X�x���A���%i֒�%�1��e�ƕ�zR�%ɔ���[Sn��Þ�n�?�b���]
~��8���B�XxWы]0t����'_ �W��j�;E�y<�X�����Y��@~L�v���9�ٔVn���rF��0��+[E��ր;a��~�Ze܁E:����8�WP�4��VB���or}+d�|O�2{b�g��%2�y��J_��O5k�W��l��H�|�n��)�t�eQ�7b�0L�4�9�D�Zu�{4k�ݾ���7��f�,N�<;�o�C�vz������;g*a)g���hg�S��΍�2�Sò;��#�'���_U�G��~��Q��t �2�,P�B��9g<3�
e��t�Ss	8���%�$�x���N(�"�)���FmY�ء��(�ZHZr�5����	�e���2��'ؽ\k����!�<I�ށ����.���O���.�ɭ���%�ÁZ����Z6b���������&��
��ʾT�ff���%�ǜ�H����ϯ��!cp UK][�\�ڌ��h��!�@��3Bj��TEz�K	�����N���9���uQO-������eS�`a,��_��.�F���_I������p<�~��v�+r���	f�����A1�W�*T�9�*��:Α��	W�2��P_>�*�C�L������BC�{��`�=�ߵ>��k��J8O$�
��9�0���B��TZ`%��q�&���Xʹ���e�^5onhz7��Ɨ�xr�l-kwpkYƳtqã���~�A4 ���4�&�J�5R���~1:�;ă�HWLK��ǿpl����`k>�
_�oT��	F��+��h�1& uf�����ՑWą��Pc�N�^YpXD
u�zk<�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��YN��C({rϴD�9��Q���7u]��-��Z�s���)�S�2�ڔ�$mJ�����y�N�!���zGc�����e�6~�A��R�y*�ϐ)���K��Qr�gٶ��V���ٱ	*�&[1��3����80�o\
�*��3�<�B1���Ix�F��e��a��:Xr�v��݇3�j~T's���w�f������!S>Ų!-&4Yw�+P�B@� �n���������g����lC(�.�3[�������9�+���a5S�[v�i��Fԥ=�1���(�q\��&*�Z��E��mLL
�80F́�Rh=��J��F����	�0:�2����<^|L��Tf��I�@��z(8@x��}+��ӄ�<U�J����*S%Y�$j=�L�~�i��`�^׺6�o�����\Ԍ/�
�*�8��;9[`޽��MEe�٪Q��L������y��{�����wLKt���XE`������C�[R�x�@�/�P����=@�^K�~�t}�=��*�]������\���K�p��ڵ'^�ϱ�^�����N�@f�����kV�,:�|?�� �w#����	�ڦ��򙤃����T�GL*(%gu��	�b?�ч��4�.6�]Pme:88Ħ�
)EX+r��D�r�� �̢��X;���)�y�t�rr7����/�Nx	E94�3�;*!���#��$�?w�Eki�WK�>��z�C��t�]X���w��M{��崥��sծC�a�����vy�X�XM#
<o�h^��K��Q���S�^-�2}#��� J��=%�%SV�1D�B>l�*�V�|��b����۠�d�����͂�J���"����m�A����$��`��j���@�E�6�q9��J,aLj�g��/w�꯺�\�f��	V1� o+���Θ���	�[����qo������ �A��^�94+Ot6����nΜ�!��'�:H���r���Fy��]�hi���Q=!���C��m��<C<�X1UA�_�=NK���B���~��Iҧ�,7�Q�
�x&���w��@��a<�)�����Cec9�pS<S�74$�GM���e��}�ó��5��j";PGX�u�C���n�s^���8�̀�{��:r��}���R�O�`z��&}�3�BѺ��x��"*O���s]�/T֔ǌ���9~�sձ��ͼ'�֦�}�)���=���&��͏�#rʌ���m���S*�Y�@s�����֔�NA�q�.zK��&0k���۔I�����Jw-(ܣU�6X%|��d�M�����Z3���_���9�6���S���7n2�ݨAI�@���I��EU��k�v&��b8q�ny"�J��m4][YÕc,^�}�Wc�fF��+F�F1%
NT�BR����deA_����%!cF�6g�����Tk�e������C��S�3��<.b�LVT
w붧�
n� 4g�� �����rG�h$~�-��=�ׂd �oN�������a�6d{VڢJ�L��j|�U��A��jC`{
h�'����	�'�L=������lVĽ���B����>���kw���x���KՄjׇ<<�$���hߠ����V*�[v�28$l\^n�6��]G%]|SFWr�
N��RL�{䨩��`��_���_�G���K��'�:���ځ��6�����������J2$�[�H4��[�brn�ڲJ����PS`"�#?
PG&�f�b���)��ư.�2�߮'|�0����hW�A�Ύ@����p=ˠ*���o��Hs2rr���He"�,�v|Ӣ_�Ø���I�	"�y��oR�\E�uE�L��޴D��r�Ƭ&R�Vk�=:Y���l�W7H���i-x4f�{,�AWf��o(�f�<^�>#�jPeoD}�!�(Q$��c��+ �;�$u_�iu���M���9������n���X��}�*%��T�	W����n��Ԧ�&�{�a�~�P$d��Cin�Aq��۝u���K7E�v��\��CT7��y=��骠�PXL,VW)�w؀�u���B��'V�}�&!OO���M�ό����%5����ЮN�:�:�Z�)�^{�z�2м���7�KRF34�j�{���b��x�|܂��3��r��9�Ωn�Y������'z���h� ���$ķ�M﹛��@ۍ�q�p��s-��i� Q�BɃ\�ԛ���,����빊�X4N���)��h嘙B�&r���ʹy�=\�
����C �M� �qԶ≼>����YD�	�$�Q)F����M���W@<�{I��I�j-��a�ֱ�9-ܩ`�T�Wǽ�DCK���~�>psnWh�����U��_G!���}X~��ݜb\�3|\�o��]/[ўq����9����`R�^w����"�g�B���>�.3���8����I3L�nDQi�xt������'v|��<����fm�)��7C�&�[Y�_y���l�h�l��m�jc��y�g�sey�]'�VZE�����Z;��^ ��V�AX�?��7�50������Ӌ/M���x�X,�c*��;�X�QN)��Ȝ���h����Q �y�.g������,����	�a:~��5? W����6��t��_��<��"�6(5�!֎������HzF~�<-��zT�kw	)�Ck�Q)&h�9�xu��T������%3�Z���&�Q�����`c2�b@�&74���A�A���G0�1��)*�t_�r}2�.ە[��i �ƾ����(@�%�SSKƥ t�<0��ui�Cm˷�r�"͸&��/��I�]��{�u�b2���4T�+���%�ӧi&d�9c�K�J\�^R�y#�]�e~a��\c���7Q���K9o���(%����E�	H�^����IDer�x�_��4!��W]�pd��@�!�m��Y�OM��Q�����OFyO��3�Y�����/�P n��O�����EQ�$��6Ϡ齒�%���;RS���:e�����Pۦ�#t[�T2{~�G�xb̙�l܆�nR�-�-�%�|5���D��<���g0aV�f�`��C���=���f�����}�S"�/!+'H|j0cE�h���o���%ĭ�f���i3;4�=N�;��MO�@�R�yi�����	�~��#�(�s �g�<d,�ǯ�L�B��m�����T���E�'�v W��V)�3V����E@��?%?�c�~=$�@��Ү߂�MD��t�%�:��-֙���!^�f_�K,��vJ��i��#}2��Z|>J�����S�s�U�.�M$s���M��b��q`��k1Ȇr�������St,�N�����m���L9�Y'x9��*I���v�����b�� y��+�Y�Ez�+��R���q��˘��I��#�(o��Nme�f}x�X��X	d9|"���S� 朆������"�{ukP%{��+lM7�:^̀�ĉ�$2�?��?h�IU0�>~�ǽ�j��oI _�:��7�eE�"�s�OXn���
doʓ��8��#��0r�kS���60ʓ����m�����X񣃊&2�6�@�5�kC�����%��e|$���}pQ�=�.��e��P��IL���I�~i_6$�a���{����%��bP����M8@WvT��d�q��|81:��Z��{���)i��������j�MP;�x\'C�Ȋ�����p��mO��Tȓ	�ȏ�ȸ�A���|���k���`�"�M�pg�a�"��\إ����1#ױ"�WG��ʁS	q!���" >�e�/��܀8]�֑rgb{KE+�HpgK"��ȥh	�)`+q��]��/Wkr>ؔ0p%;c7�XMV���[��H�7@�mk��ʇ�/A�{�`��X[˷����_Cο6>�,c}�hdh��j���VtW���J�f����%�hL�ɈG�+��7��iK͓�t]5c$��vҗ<������cH�3G"��`��`aB�0�ݺx���Ir!X"˕�	��P��� ad�KhFvN#�{�ѵ"\'X���P�VO���!5���
���[.9�F�Ԯ@4�t��U�՝SAzR?���2j;��wy�Q}cSM�!S����_��$,3Yk1��Ū�l�KF���\�$=C�1Թ�R����vD(B�N0A��x�ń��Y�S�'�B�4����Z(�C7EŠ�>��%A_^KM��o"%N]8F��/@��6�}? �$��Cn��a��}$͞Xb��J�����dJ�B��@���|!���BQ2��*��@A /�Q'a��V�|�ISϸY�z�T35����i#���>�(
@8���;�w��ô���A@\F�H]�l�R�U��!Բ�9���)Qsu|����
�Y̓D�p-��׫j����iI�t��&D`̞3]�e(̢��1PP&���qwK��h4������v@��%�V}{Q뱕lѕ~�vo��aM�3��#���{k�ɨA�)������\h�&[�|�~_0�{���c��͝Lo��	�q-`D�0oc�u�I��I�#�8�� �*�%����?� -��U�%t�:�*c��HːV��׷�
�qz��	�G����@ߤ*���-�YCv9�?OS�1�d� ���Y7�O��6#��:;Pf����u(��wy�@!u�dg���л�����a�-�~��oW��
�nwmf@2Ӆp����ī1ʷ�i���3N��F�|��5��}.٘UZ�z���ՖN���'�i�|;g����Y+O�W����H��ڕ��}����J]�y�����Gf�Z����+Kו��1�q��Ɗ����7U6�3c��.&�v!���j��(�9�U�1�I�e�Rq�/}�S��7%)�DI6��{�J��b���)}Nd��]��Q�^w�FFy�&�}ڒ�L��O|�,G ]v>Q���?�R�-87�T��M���nkޮ0٣�߁��)�R:�W��g� ~mA�Ўf��V�ϗJ��d�Sg;�w��bFw�fY�����=�8��PMVA�=��x��՝� q�kЩ� Q
�cu����4�y6�X��ۅj�9�I����Z1نY�i���I�R� 
����.®��*NA�jQ*T�rj�W�<P�@o֟[��w�[7N�@s��O.m�fm����!S���7efj��t�Po=�ҺNeB�I����J���$��$P�"��h���|�y�l�N�v�1������^#��Hҝ|�~,��ٍ���b��� ��qfo�r:߯}�b跺�0�	w�yG	N�?�����ߜ�q�S4��gŇ!�]�NY��3�Z�8��;($>��E]��+E�rĕ�A��0{RX\�r��."g�wӻ�j[���\�_�����F ��f�tgCE1�:ंܨ�-�=Gɏe��ڏ�9�;�!�v ��m2Z�n�>�t*��I$�������3�lll+ ���2ӹ8�,�N�D�,~a����>�5�6>4�{�h�PL�P;��,WǠ}�W���x���@ݻ�CH;��1 �4���t����	
�EL����۔�P�|�K�n��J<��W�9���� ��*�ӾbD�ј��8��$������ST�yVڱ�����~�Z<ֻ�(��~�O�L�/!y��w�P	(����h��{xH� ��'^>��TK0�8Ԏ�(���K�l��+О�ja�^����vX�9Ի���@!�W52|W�+x�s,���O�^4�c����:�'sר �*GNX��w7~�
�B�����<s*v���f�p/ߝ9X�6<q@@T(E�h�n?P��wA�<���n٩z
�k���Ō�P6�<�_�'�B�놪�_6��|�3LB^�|P�qq�R2 <����,���8���;�F��]�;,mQK?_�S9��PB�iϼf~����ML�B�_� bl�;�� ������U��Իrs��aɰ��H�|�c66����s���Uل�/�Ѡ�T?�*�:�&��fF��-`Ek	P2���S�P�:���l�}�����k����a�\�^7������$���NF b>od6|�c�ނ:��k�����"6�N����ı�|�����˔"��l;��"�o]��7Y�e*l !�S"#d�h	�Y�l�`q����D�0Ԓ�L�x�w����w!�Ʒ�3�2�]8 �Al�����d��'�[�7��~8&{|�{m�oWV:L�N��zI�Oi�O���q����Sy�Or�R�Q�h����^c�&��ƾt�zAQ�R�����K%-1e���'�j�_�Ÿ�`%�Émaݑ�M��g�ʋ(���6Z��L��D=͎๦�/8S�>��bi��I�%<�����	n�#�,��cdݱ������Bh����I�I��=�ޣ*�̑� 0�fV֗'=HD�}p�[É��|�d,ҥUTYUg��	�Ee-��E��}Z�S�j�9�J3�Z���O�6g�3��� ��rfX��0��_V1~�Ym�P�AD}����%#ְE�v�+Q���8��A0��A�%�|h���
�U�2���{���*I�5�G�3A�����-L-�~�WN��Z�D�$�p_"9����	�	m:��u׉�����l��˻���^������(^hVn������lU�K�9E4"�ą/���q�a!Q K*l;ؿ8^��n�8�Z8t�f�����>fE!ע��`&s�����ͩt��r�L[�8��B��gϽ�t���	�����R[#NJ��-h�~��ü�ai�����'�"[�0�}�(|������!�Z���i� ���zGY��\��l�3���B��M"&��a]U	�b/�I���qz��\!���8�K��iY�z +��/�Yi��S��?�#���^��t�vI�12��:��P��g��f���V>�4�SU�;p�tG	{�7�h�>��{_k
t�������������ڌ	�
���v�:V�`���C%O�>5���f�xa�ΓGP}XWg��6�a�$\=�@����/��q�ޖ�M�&��?[S�`aLm�M!�������Y��*,g��7R��9����e�Z�?�&��TrRw�*��!j%�˰�'������ʄ���᯴t۱�GY�`��_��Q��k��>���	q
_9����@�Iڒ�+Θ�<o�Q:/�>���R�Eʩ ����P��?���rͱ=�����h^�s�B�_}F�w;l��̐���$�n���s�k*O����������̓/yx��L��i4�S`;�_
�S�_�(��ס�+��	P�@�Qρ��LQw+���M�PE�R��~1�����4`6�sA_3U��۷�q[�$��#֋"��I:�i�'�/[w��;@�Kb

����k\�T0<lX��l�\�/�rKJ��a|
s��徧%���9	�0�s0�╄��uJ��s�x��#�U�5����Z��L�iQ �?iGu���Jo\M��sOp9px.�b�C�L��˃��م:���u_���fD �vl��s{��s{_N�u尠[� \��%]8����e�>�jos��6�V�~{9L�G|��Q��%�o3��R�,��. ���[�aƋ������Ii1����C��6=�f���f>�5�Ѐ�����TK�ѳf�Ng��1�l�0�T���);����T|� �|K�V,'i�ǹ���`�+~L�W"z�Р*"������o����Eӯ� 9Mt0�=ϤEc�O�2��)y����y�i+�����f?�Mdij���_(`]��y%�N��
ߕUJ���㚟\/��R{3�O�Hj����L��DVm�2��])�%�'����WN� 5~�&�N�$-Ld��E*'��!��Q���n"���q�8`>��I����&Vp������ÍXqf�h����'|ue��5�`�W���JJU��g�J�9�1dj,�9�>�y�+(T5����AR�j\}��[A �~"�b�R�b�������A�z�8���O. �Y��O�b8�k>�=���/��P�?��p���86� ��)�s�<\���u~��q���Uo
�b�HEǜ�2)�2$L�%������J׷�C^���n��DI�q�M�+���3�Tɳ+����h:���d�K�'��qLA���x�%,*֧�0�yfw/� �՜�N��,�#>�g�i��E��u��ک3�C���JH��M��bzt=�݁/�?����^���Q��+��V�i��N�� �I�]�NBp���b*���*|aл�p�-���^�S��Iu{�B��Q����#"�r�h(J&�5��Ôtc='xr�(���I3��[}�AU׌�Q�m�"�[�x!wP:a�,����Ov����4�d�4=P�f5�	���U'iu�帙b��^U;~�t��$\J ���ݾ��1�[��$���1*L������W<�5����ȃ�/��~�S=�E�\=�TI��tlc��K���ޛ-�)"~q���M���[\��ݣ;�F��d-��7���� Bf�J�ʙ���T$)I��{��Oٳ�F��m~�C���w������	\'M"�nC<ċ�ތ�����tv{	n�H�Z
>."d�4i
����̿��L�~�~1)��L��2�Zu�u<p�A�=(�Zg	���9���81L�����e��Î�k��gU�����x}�� u�CH���"�g����rjШ���L��܏S[Ƿ��.W��-��9;�v*V���b��Ŗ���r0a��[=+�?P ��ƮFe��;���c�ŉDy���W�S>���\���S�,��>�\��(���&����et,'�ûr�{� d��Z7����0����9�L� *���o��e ��5�����C>�m�$RY�rʷ�/���j~��[��7���_4�k�]�z��k%��OUE����b:��7��ϩ�A��utT�b�e�VIk��x]�ǁ�0����<�Z��L�Ap쨔D_[!�-h���V����mJ�ՑG�"�[P�f������EG���`9D	�Nq�ԀL�G�K���J󸂍�P��Ƞ	w=�w���Cyl�ޖ����g1���y���_[�ē�1��#7�+�u�t�%�:�Y�r}��/��`a+�mw�p��µ�J���|��h]o�`�,ڵ^k��Q�b�9:�,�[cX��;ks�&���g��tt�*tJ�)o��	��_*'����v}��Oq�m�yD��G����.EH���O�����"{�����=�(�ϥF�yw$��/�fr�fa���"��|Ɯ���gs�	#�Z�Z��Z��똮pʽx�E��WC'��7����S[�?�ރXY�(V�ո����n�v��&V���jSi��Db��3�טˤ��ݫ9����
*F�E��w�A���a�@�+�,/8�p�z���%5����q(W^���!֖���/u�W�Aʉ��U7C�<I������ĵa��{�n��	=zfX�s�)g��Wn���Qe�1%��k�3�ߡI��ӽ���!��'lyxƥ]��E�{\I�
rY�������Iw�Q-��d�$ǉ���'^���$�(-b����J|(���4-8ڴs:�W�"vG&$��� #-6�&Q���gQԷ�>�6�F����E�%���U�����$
	�����Q���s�M���$9TcX�2e�� ^�R�zj�琮�v#��E��H���������� /'�)c�����u�DO+�)��I����*ʐ��e�G�HX�D�M��	�	ZdNwf���ՒCp�kw�`��`�.�4�N���|�v��Lt@�ۢ��ٻsu s�U�ۤ�>$/,RςA� &���sw�S�^b�3��J�$�XR�7��e����m�������)��7��Wa��g�ڥc�#c�4�s�!f������2uٌ4�y75飶�	���F�������6|��0���WI�D�y~�C�cv��P*�М`���E��X��A�uNԾ�l� �O7Վ-k�Q��"{l,x���vd��>��.�P�$��B�~���挽���s}<���>��ȱ
g��ދN<�n�vL�a���J�za=�?��z�[G"��'�9��{[�eAǟ�S ��x�@��~���[�si���Ч�T>�ݠ��@�W~�?�2�GN���)RJ�Z����	&�xZf�Ǿ�u�����/L*�%��8�3�Y��s�S7vh�3+�]������|��"��2I�v�S��N� /�3�����\9m�He3"eX��Q ��/��4�q1�ZPo��f�B�]�	 �R� o9��=�S�:J�4Ŀ ��G�@�;�^�U�
(>4ҧ�p���aE���������.ۨ��\��H&�2��W�W��_��^��V�7���`�����I�Nd��ӗ=oɜ���TC[�[`W�i]iKbzp"nQ�/�+9q���uӝ������o+8���j��O�x�J�l���F+�˼��^��٘�������#T��t7�'s��-�K�JAhE���.����YZS��DI�l�4+e;�QVڄ=�C��Y�$i��a�!�.F����z��W�Ғ.R,u	!����^c�r�|@��dVc��m��A\x���Җ��$:�ew��@���_d�?or�5@	9�R=�s�z
_@�D�?�7���	Zo4�$>r��L�^���)$@��~ ^&X��U���le���fK���ڤ��&1h�7�H�d�XU�Ĭ V��a�c���L�,�N�Ȕ���9!-���x��V��z�J�fm�AЇ�
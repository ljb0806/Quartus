-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZpeEopvISJKx1+NRyeAWX96jR8MejYSG5GV+Qy/d9iOj7vftTqPC1yqV+O7nYDqWn7NzGSNcSBjM
ybTcJVMeVShv88VGYlF8CHb1wJTN2qdtlIaoJhcVHV+b/UMSiYEetrJk7EKRRYl6LkdpiMV5bOw7
pJfIEpHqVYwzehahXMzgAARFimEnG0SBIlIvPHZxYMVaouk5EEUfbN29R1jR0N5HytHHnv6TiWNL
vIyiDjqJ15xlxWU9Hz7bsdyU4hLeXBfEk5TpGDPu485hyHevLO0lqIo5ovecdOLtfGWrH5uOdYnT
JIGH2Mko/eY2Vsn9XLpaVZM5PckY9e333UF4nQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 86768)
`protect data_block
bc+ktTbJoJnZRVuGWPLDdQi+wOaIy3SzEvwztXV5fwlCmVm6DbF3ApwNVZTyYeEzYDiwJauq2+nE
wcEgjKOqr5R74bFOi1JuZEBkg0fQUAkwgadUEsCcpr6sdWnzFebTAccVAN/+jwxYVpU2+e09RBZH
j0gocs32mnuixyrsyU8E6/51AYyF58P8Tr52teLNE0mMHoON9FbtHdiMjpGeLIxSQdW+4Kr4Uq5V
P6Nc4xe6tpuI1Hc6DcY9/74iiGLbIrHnlXsMcK2s/c7hN5hD1McMe984vvxyxTGSylFoA+2C5iDd
4OdhEGTn7+uF2X3sR4FH3nJf+VF2YScDBH7iBjPvDoNWFrJrVxHlyzq3Gg0BhBvJk7tsbSX1Quzh
a1/8kq8nwIQ/xZJwqOGITUQ97wC8QB+983Y2/Hpq7YFNW9DCm2I/Sve2+JZ4sYjbbZjNycrLi/qQ
pIjxemmZuZBl5XFUZu+ZPSbtNTldfnU+pVFYL5g5LL4lyc34JDL2JwmX+WltcbHIT6j6nlGmac8N
4LUozXcuhrySPwzL133Q/c2Kdn1cpPNSrIg2AUFYtb9mZzpYIKNX1/FWpLEcnj21q+FwJn6j2Hl5
q4cvdrvGSmbFws3xh7Zp/PKvvon9Qu7m4D4vrgH5bSoHhtVZHoOjhSzvaoK92mTu2o3pMySVcz+F
iaLXVzl1IMD9AfqNCvZVlRSjSC7ec6QYYoXwLBrjExZmubX+9tEZr0lyVo9rBHb07ltRtxHRb6N9
efLORGshVXZVRV0LgFRwxX89ho0nD3rGnTDW9teOVgY9NqTVjA9gZN1QLG+dqcvBIdM56/VKeuC0
PoLEKDhJNs1n+TWz9QRbpfE65omp4CMiDt6k7zcR6FHbMKjOlrFzcRnXC47Q6WNdq39ccJbONwD+
ua10wsz8jofOJatpppqlzsYKKPTwNPk94fMOtg0WkExIuuQPsXxD6aoELE+BZGd3oMhnMVGa3/56
j7QxGadV4BoaLr5y7xlGmzrT5bAowpO/xYrv/fLYLDUOQTe2p6YyDHjnMkoclh/qQ2s6lnBWg/Rp
PXFozY5qSCNit4W6vvdJdgNUN/3lnn9A9kr6W15zgdpCgE6aGJrykbCVsimv/HuLoYA8SfwSXzWe
lGZp5R+hEtQ93/MG5iCZaPDB4W0fCZCuZptoc9W3fuOIsUK45VIAd8hBVvBuo2sndiQDp5EkFkYa
uVCQD5qrY6+ykCCuMcgsn0ZeW+d8WSn2Ev+Dutv/eBmBCGeCesrlGi+nWaq2yPbfadAeesG6KM7V
Gqp3aaozgj01lrSw41W2AdL4JwWdMj/D4QxhqCPxBWhjALxkf/lgzGfazncCP3tctLVWfxHuKlqz
N4TL5XUstbVJS9ojIVSaZBVZ71mnZU9kgVaIl7lb2ap/2uO6GeX+lmNkvq8lOOjdVPkgIkVwJjcf
Idv9NAzGMKXvayquYWO05JLovusno1lJ7IvDwXJHNqyk9AhcdyFM/V2PgXubb4NY1M3tEBZ7l6rD
ntMCDcMlOa8ODuoCSqSv5/toXJ30Z7hfh14qMsw+/yUAqE4k0D1Fj+D3vxo6WfMJHDKaXbaXaWWO
ZOX6u4md/livOcxBKf2hpfWeJdN+m+9xLQ6ydtT1H9cFO/pi8OYpzgxwsUMK95feFUDbFF0at3X7
uXpFktv1M6NZD41NZd3/N74MGaqpElWwEqcNBHyBzx3LW+0vrwry/JYOdYibqW6DnSXYKFWJYgK2
Z+hScBPrp8vgj10lZrv9Jx/nicQ6ooz+QqSfa76QCH+y4HLCakuToZXSjhFCulYTLuwV3n3iclL5
u3w1XVYL1ZgE6gEfpYmKw1VWLfD+U7yKA8FEvqWJrkShLJVEA02qnhW9YDaXUM0awjh9prOjNV3f
9m+zLKumtynLoYpLkD22MasoeDE2xYojaETKznGSHc0uP7QpOu/98rfRM/SNLr5BifOkjOXjx5WZ
8pSaP67ODjXnGFh/u39PUDDQoqPway+qvVAkcm+o/RgaQOFYaf+xUvsbqhi6ndKfZE9LCeAGgaqh
rrivdHVFwg1k2pFIsekHmCybBvAeRvbgXJXjVtOcG4EdmckbKufRba+5R3A9QXR4da0NmYvEtDsd
T8Z/nDansf5AziwjCr07fIUG6zF3c8A7r9bKXwwBK+5BCRshNr4hIrbhhkj39z6B7oz60w3Uq8hN
gPt8fv9U3DNA+kjnfG4ryeQIG+jXYBZq8ymeL/IMJttc2FBe+yTs59lQLJJQpUB/TTIstbebxVsa
hedkLXtJnHKnvkK0uym7h9h/tc29NocI0Td7bDiL/oMllEKaeCrjkqi9zBHmFg0PIg0+b/rbeHTv
J1LwBA63ieStsTB2g985msdJ3iyGLFgHTCHV8EzB0YXfY5IBioD63f8ENM/14QwbHa9QISRX5L8Z
gRkQH9ahBjHq2c7RrFzglUCCtlHT+Mx9r3hdt477FqG3joj1GLVnOyguKNYDtMcNj1/HqfC8LqIu
oFGvwwVPaCSFj3IhdifgqoMupoNAOsOhByTEyOwWRjtOcqRPgWVkI8uvv9uLfsLBmYprex1WX9+K
GYivrLazM5Jvtad9aW09tO7gzV1Vnjhnr04iUaMUfEFcckajBHsT6V8pIiMaWFO0txIsuQBboLRI
vDIC2hRrCHgc2I+uPdXcrE0SktGvGQS67TbuF+IhbBHqF5JXLDY0gC/NmeGjFjknWdmyVss1wV8s
UyrywJb/IZo7512khIJC2+rEP49HSgEMErsNk62XlVoMTCoIvubzFiG2P+nXAuoxXtg/umW180FQ
Wsf7R1g+JN1dHSXfNH8nAHJNgs7ckhCE83KdOOaO2lNfP87se0wTJk0fnkaOkZhrFjKs6Td46LKe
OTkZEpOTJtk1mNVkkscz7gaw763Y0zxyFzePSy+NYPFjVSbQWAQhACCZhjE8RddCPGh6serzfjTW
iFfjbH56a/dZe8ASHFpccWIwCavIUvF6Zv1Jt4VQY+o+kdNEz7p1zxz4Li57wSuILUgg8gQ8aHLb
zFCgEZzQECnuVaV3lt3qmBgJQX3OiT5tKBPynkNl379wEXwoQG/X1fE8VqmYgEe02G3SujHalHbg
hLamHMYAIgmUV3YBa3MXCcRJ3YYdp8EPgo14a7BT5Im4fzZ7eiPHGcbAFKvy8UJIYCerC5/0UWR9
CC/4avEprw6gmY/rJY8tnSVfnFxoAg0we9CB6p7GShWtOhfXyGRcRLRPTo71SaDBFJjdC20XhMnI
v62wi781xMbMyaYSkrmPFi3wY0ynYMPx3g8V4gxq4vG39QuT3+CKCqh2O8LoaSrS1S+kkh7X2lp5
qFrNvuAMhjaSmJitm/HtZpRTqxQOz8trJ2bM2eEhTZg0uDRK9zA8GCYm/3skfyLaxyda7rdkhYX1
GJgPduyRvpYh0W06CtPOTniYILUOaD1K/a0xKVSx123/6gB6iENAsR59HTyJjnVFzW+Ibe/YjiLZ
l6dxn/k98lTsRlfyIqtifKTF/hkp9VnPZb4vr8QI+PJnEjjGZjS9tBtmhd6u6i8QuvfnuvYfuSpG
5+YXCWMT07Ksngcg1s7ZVHwjcD+4UhU3sCfgU/KwQ6rptHLoKEfuOzIhHhrMTLgYFBU/kF9jYhk0
ZHWy4Cx6YFAgRFfR0wCok7fDmZ4uItkfcheJrVhc3wfH31CJ9CzRFTNZlzib0LABWEqDO0NHld8+
bmweAvGfh0y+oH8g8GRHYOCuwMaRh3jjcaBzYGImstqw7dPu+V/5Blv9EhCr2+e5cHdMJOhJt/za
G5AMY7AboVTBFigZdaGNcAYZ61Jd5XDT10bPhUlK7hQbhgrxxdJBKP7jplW43GXQ9WsZqBYqc+lZ
8lyxDl2ZI0oN73AwP4T1vziFmyODxjHIpbyG30GmLiHRzR+XdrpfYi8gy0Ss2zAK+j6vo8O0BoaK
RwoTomQw0VmiRLBQp/rnurUmNIu17owMn82u8LL74CkwEXK2SFEp8sHy2dmjaRWBysoaZWxRzLYb
5xyPOp8Qo4bEr0dPfpkrdBM8lssoGsDuwqegJqeURKdUgz80eY2q4S7wRKW3En8IuMG34DcWlvij
USy+KVHnoELeYPlYKKg7neoAoZMFXmPirXQEMUx/WiFYNC5+Ee75vtzCNcqschVLkDUsRMDHOOuQ
uwQxyyW+nyy0p+mIjn+nIfeaydPZmx0Z7W/FHjxIuwr9l/+QZb3ag9YM64CRNuQSuRobb6kWUvQc
eCLqe376Klse4+HoLa5PO2vGGAU8I4eDaahGyqWDpFaikUeZjED16x24PzOrOQ/KuIE7Y29RVgf6
l1+Vzy4EdrBn6sfuyLHnYZt8DnRT0pCj/b/e1yKaHVjrBgzp1hufS8LCTT5cPW5lL/nr5aMZ6gXe
Uoorrq9vKnG2nDSDv6opRnSTvb4f0xx6nFvwmHnEEyMRjSYbzEu4nEACnt5h/DMR/wbDX7tZo2Rg
ff9jGN0V9Ls+8aaeSKpcc5QAxyr0bOLkHHFfYcpFfIQ4EoS0J31icvCV17fXFAXX2FVxjbv84Ybh
yWMSncvegLwcgyT5Axu3Dq9YB/sgcUPUy4KVSvdjxj+rCcA48zHMBLLmkM14NKHLSMcLRScQlL7v
Z6UpxHtVn95efbLlt7ricpQtj86zw5meXAkIpilutWX9/NDFu9W6D4N3Fgnba/2lXd9o26FS4Yni
SAJC762V4XoELhK316X9XPifuVBumROS/Q1kCKK8OynhRyaYX+ihkcqNmamazQl0AIO1NavcT8ba
g2XtI6Xf7PryWVAZ7v1FJdXaV3Riu0Fn19V//e4CySO2GMGrkpDXfdlLR1NFgnz7Ts2Qn2lQilxK
l0Fx3OA4wfiLpPNLoNv7W/GbY864NuHhPNuD4SBJjBuw6Gww06LHlYV9bN6Ea3taP9Cy6fDvdiJp
wpeXwywE6s9m7R/MlqVDVx6U/MMz6UpdekXnoDmwTF6Zf6CfA6cGwE7t0cLLUTTpQzR1kfH2AZvN
YrkfMFcprhJrWD64D7vSVhHEzQ+iuqt13opt9Lr4L2UmWqPMkPbsASfGlTVqow0/YmfOT0uvYE3+
D3Vh3qEuBdZ4fK6wbQNvmg+4XENrZ69xLfMmGbymDwFUevEOhmeQ3UdfnH5vgnnxZ91y4hY9mhYV
c0RUuPpNPWaa2XtSxHZuz/LxMDnKEQt7j1SUloJZkYS6jvC2xqtY+g7j9c8T+Cc1jUxYuGrJ+p5e
qe5eTXgRGdf/3E5s9UDwO2lY/lshFDGZUDc6yX0jSLDlpJ8n0IcpaXRCWWS8+u2cQE1wcBTvoY0R
0EAz4B4MfqK6kScGOa/FCv6qRYnSen/D7Yqhyidz7v8HWQ8in4SwjxnzJ+WYYlTYEu+isBe/pzfG
RjrJdlMg1Qn7UPnfTuAFrmmzoLf7ZQoBuZCqE77fUy73a0XVKrD4ereXjXWV18+EHOdSQL/KbFxF
puSGR/aoiqWxsEWD0qSDPKh01/L9QVJB4buSaEbO0k0QM68nj6aVjZYwG0W/yoTtNBXQWZbedk45
9+rUDMRd8OEsghVgOWqsYnyRjWFqV8DHtyObMliZc54SrLJTGbkMmIjc+0XdzOWtZkmxqtUimKIe
+Vr+WLOcQ2ntpb1w0Do4IXY5mhVVHjYsyTzTpJr8WtW5LnO2OepBlnIc4nqzDgYgl0fnMoVzgCCF
QWm2aEn+fH27zT2Rb7/ca9xtS3nMCGQtec9OrgtZ+mZqTxwxG8NtDZFji0zEtrj2DLuP/xbEwIWS
7ddml2ldoq6GGFvB8fI11ZfrhYi1DSvEffWfAaRjRip+4qc8pIu28akX8QZNUUNy+J8RIKsn2O/K
vjy368ilb3wVL1zmOERM8D2FMT71xuthhgenisdJAxiZGS5LeeQ7XprlLTW+j1Dfe7/aJvBxGkuW
/Oc7MdO2vAw8z7VUtWwgb360n4BRR+3FTNtvNIfnB/EPxwtg3G2HrBkWltLOBrQjikeSKroz+251
M1KsFERJAsjgcTPGVLW29kuvlp9o7j7yDfqQJmELJKEsdUVJTwev1xqfTjfFQAYB/ClLSKSCa0BV
fiFvGksdbwmKGETQwRG68uN/6rDTdCUBH+j1aJbur8hZ2iHYPU64Kuy7Q7PGngu/8pucB/lQs38u
QC7Wd7x8eNi5CiDZ1msWcn16u/kZ6QpeTHkZH8jFAnHrrZw+9LeOWp115gds0oll8ktSXiC3jyLL
7hz47Lc90Sgol6QJwgoGkbxrrjJuVM/wszFrLuStsndnyJ2r4TN0oTBuqGOXLLqFeLWOTlnspv41
TRjm/0bsd1fEgGlLVTZ3hS4Rqyl1gLoIbQFicYItaKBe7yx/hTzw749IkqfTB5XWlNGPCEBTuKGR
o6pLzphK4H6S8v+ANmd8vcWdLSa9eQWHjwVna29ZK7U4TDuugKWl3+T/OQVCpMYcIWqqeg+MlbgZ
glfp5upCv4gjzqL0gzFg1qkLP8Lfa8rzklvXhMxXOropJ2bk47+TNkB+VrLSyWh3EsLIe7EaaQBD
MurYp8ZbBTgZ5Nvb8oETd5zUxPSuynsnyQpYXxVBwIy40N6x6lu7RwDVFo1B5uFvveyZqO7X8Dqg
HmvGMOOaKbQJgTlHjLESkXkUScXXGoqEs/0LSq7w6F3zaJfJOYvhe+8JlTInuDtuNw5RUaqp6Q6x
bB5zRQWkZ0gxQU2Zx6bOUHs4BzJtBfxKRIT6Xmn1VRUxGRXiu5wm+sigZmxhsHGzdA1xuoJCUSwB
K2nz79+vxnni4/WtcHWhlxRQnvDRW2gDpq4a14qoUbeYuhRhVfwIsO7Jay4eT8j3IN+JWKHP6aF1
uabRe7n7nnb+5+jbuMPrkSQXv1KQcUzZsj0eoj7wKGw4MPBTBFU4IhJA56x4cJy89EsAPnt8D7yw
9QEA3diP7d1oH7vu8p7iXTVSzmVOOrOqaTJIgMWzF5uxkU5cc8w2DHXguO3HXSILAluvjO9BcOvZ
svlYPSCXKPaPXeIvj0o7DITpvjWjhbWUPeGYwojKVATV5FaD1kbwFi1FPvRAd9x0dh4Pwo3BJnJj
VKn/YvpycNd+eaG+EJ7I/LFjKDdDKpsT+YhIn4FELb8mtMy5eeVFj5wnk78NEulpBxpUttQ1FtGT
q+fMUpoepnwBYMf/W86dqgcf1trcOpBRgRpdP8Sj6jYNbzRslIvV6tUjQKnr3aYkfISZsSsOv+tG
jYzqks8anz3Rx44EdJLqL9WTehGaqazNYCIm9RCeTspBqAijsLV1VJhCjjSYW7zkzCFJnSJljcdn
DplOqKsmzP+mizuzTeW71KWph2NCs9RF5t8aXiOlR013XORLxgMw9FnaGV9jouRr175AZc0uiZKD
qnT3zVyDIVjxBfP9hlNgGr/uqgjOpRmCdMIRoHl202w7s+QvrXNxO4xglw3JNagv5L6x4dhU5bPU
el7cD7Mj9+Q9Gp4W9GdKiwxuc3r3n15NzgJokS5/94ot9TGxY53Dv7qzBycY3T1JlsDa9AcrACrV
yLVXfBT5jROW0oU/PU3YBRKHr/byeZ+q5wNXNNp1MN63/QKXVQ6FEnALAPpZFT72OxMKpwrdtlSx
kc6WAEVVyRZkl+w4sb+sJX6D3S6m8gUSXhcoyu+3+YMrI9e9lxaPty8HlwcJYJz5ZZprimzN6DXQ
k9UBQerW/hJdhcQ9Vm74I6RiWDJHiZlZiB0aHQWYbrZUgAz6ZdlxxbRgU+idOIy0Fbi4opCeLcnI
wkzc2hmP4rGpXXTudQPDPdyyCkhaijpSsoEC934z6wiZ8U8U2o2jMjMT7g4LUFYWhjiJj3dzCqdS
03Nekl0CVXRRq+quodYBwjecE+zvk39T+8D+/ME4K8sVA8RJc2UGESHMNswMi8btyGgeTWXnSxl0
RarCjebFOUOdbqeBtv/Q3hyW8z6lfoebAWkTon3Jq01SADiK5UQpskUg6ZAN4n6B4xFnLQ8EA1Cp
/9veosmw4Y7AJx3sh93czp/9PVmYB/OGU/T1u+ipRaNZZ+nslr9t4h7pkni4ubkYCoy0gZE4xUvT
431djWRtfRjvMkq8RlSmSyZHcDsvvNem1WBNvlFt6yC5NZby0MZ0oNAAawTCcu5WL6Nk3A6wYx9t
WXIWkOmPOwbOxIDCHgqKTxmXDYOOZT0Fk/J+tRDUliWOsU+kG9d75HhoTMG4RGYGR215p0HoPTs0
o6w9AZNfqphGIidF8u2oS7frLXCoVv7Av6bhtbneivJ442hlZ743u0/UaaNI8Q0hdGXxDUDp2+43
KwnjP6nKE0TkxUkueKdTYTDN21R9Ev5wAIj7w6RZ0CddiKzzmfERuo28KJTWbBW3WMGYjTzb4798
K/V8mkosxGkdU196WrMnJsoJfdJynd8oxMrnTnDqzVZ4RWfKu2AEyreVzkPKMm7vYCMUfEnNEQN9
lDfYbMwyb2BGz0wD04y6Whg+ljK/Z5RWr1603bad+3U40cYbhRhiZHGaxk94GEer//+zo36ZDe5r
7gJE3tcKIqoUvOI8P0VRDGr0i6U/ffx1KbtdnwN/ESfkwflqgpugouKg9zI/aSG2mUEjKkRu728w
4vhA7kUb/Of0ccnoLsT/WrKpdQNGxW3v+Dnrui5L4Vmfs3E39sQ3FbNS2wc++6RFgfaRoygIe1P6
r60AOt+Jnt9xYlL/dSWVCkuRq63IGpECTPlf1+lev4iBj/ksXEHyLgbFMCEzeuV4b09DP4N8JKkG
yOqtHn3tLf5OnDV1XeZo70oEEjnei129yJ+f9lPVSgrhZ3KOjvdxpzLqSzgOozWFJWMMZcjFxF5J
FKH5u5Twj4RxF2JpO9n8BTm+CcsgOVWGfho+6WWaRz4umq8f7GKu1IUYnxq0kNM3+u4vmrDkKe8c
Qr391e/tfs0s9/T5o+YXuMvVlKykzqwiCO7RCDhZageBjPcctvxZexmJ7ikAi2acCPtgYs9BnmGd
gp+Cm9Lt5kS8ngN91Jz+Hdk6NoHvSLvsvh5Vlefzkz/ixYhkwIw130uuapr0rKn3wz9SfeT8ss2s
XbI6XnsvtgBcCjomgPwl0UqQl6ZcGsZ8TbghjZJAX2HsSTnBMtdkiCXk7DUpHgYZVB0NWXBKZMhz
GcrpwRZujr4X71yXH6arK0nrZtWYiEWnQuebLEzB/g1KjOKxfQq48fI/bj1Twq/k9nCCx9DbnCgL
IAzuLePLl1wMvYTGhFTh+NMiP8fHWF1bhXE6YTaoOS/DPn2dTnGaO64pvgEa5047iaI7uW9JLl/M
Be870jSD/dMkpIWWv+ROFs50QD7w2n4kTYrJyfu1e+ouo+YxZpesQZprpaWWYOH9mN83RmE2U2mz
cPcB9+skw/+f36yLGNQXdkA19hLSmvwzJO2XeP7ykgOWqbbJZrhUt+T2ilbHsZK44T65EMiKIwwW
AcqBY8s4YytLdg/dHcnugSwQGly3j4jXOjdYmQ9dsr5gli0go9Cu6fWBkIJuP0guKNGbIX4pIyEm
dXUmHgpxoqeMH67/gw/k0lGnDiPgzFcNnNeWBoSVKtdG0ezE1pGqLrzkLNn2oPraAGxd4YsAPnQc
ij/VeWn/qufDCrxI1u2li8QcbIvgIIjFiorysCpK4xu900G/jZcXE3j50McL+W9fgOFyyw2IXfFp
rpQofkazzb2jNJi/IK0tydonCyKgmwF6ZMEOFJYlKxfrnUeNqkwBtY6Jn08xBazNn6Z2hnleHo1l
Y2Y0H6lwvYHcovmX1FmuZtGllOJpSN4xU4LXBE/J8ItUKv1o9jPF6Ta0/xf+TsuZtPgDKzZd1gNe
h0azrRLHjF1hesSlgZmIAosfnVMHAIc+LDm8ajyrrUJcktTxYub6SqLVGs7EP4MICq6bZCenh51J
WPVlzRm43w9xembDm3bD4/JK9gBjXuky/Nm09D3vJLOzaHZIWyPgR5NP2Fb86yDcCLtfcqpdllPO
ikqxz3iOnQIlA2Xv4PN7/Zsz68Y9p9WHoH01kgMB4pA/C8wxAtrQZi5jtb1d/torm/MLvQ6x+n7S
Ueh5X6clMzkpdEc357ACRzdTRLDtAcYbxhWpnXPJO4GWUdLCekaoPtWcweM/NnPaqRKKNfPPsrhV
sel1jQQF4FZjCl/FfPlGK8wWndVpG1K4qVLJxvY+j9bFeOLMysqkutEJUPytNNKEHEYIgt55D98z
LEpSNAQKlTAFGpIxMQOmugcCh7Qi8Bjog3qpw5r64XURbFNLGIJJfoKBJuB8MwT61jNvFJZqMxLy
MkUF9ALtR0sNNYg4H9X8T2zguwTUMJxugkO20N6454zYrbEsqo7brhX00Gw2VdSvuIjZs1OIX9Ey
0HbSrFDcCCc14IOXxwfebeh3xOSTS+mvHV/BgufRHbsA0QHQUZl4UbWNFnS7LkZorcdWZzke9qZN
alfbyKHImMRTjCgzQF+774Y2W8Uz5nbyCJFsfSi7Ih9MCol00C9KpTfPKTIdg7jIOHX5fz29nlc/
Bae5PfYdr+ufzrkrnX8J2knO83WC+C5fk6sQfHhv1+GX+hc9WOX3oqA/iShyFClMBLKFP5LEQ3iJ
tOux6NfSkAvpQAhoeMf2NiS+pn8b4h4IzFL2C3ChpRo9fYWpfp/lEns1fBm+K++YgiJrXJHmJXjt
alxfAJjG05kYII+DK+E3ibkpkzgQCM5g3LDLFk9GMR2JZ/vS1zPELR8CwqTvTOtrTNLD0IUdI12g
OHKsvFkDpd5wH1rlTXaV6IdUZWJIZRotbkL2+3wlTbKK9edbBKXBHSJD1xmsdl4YtG5Z2MHbyG2O
9WTT+dvLAimaUELWpMnsDe2DEblB6a4lw2A9bCNR9lR+uaJzybepZyNKi+th+ERPUdeZrNA/pJ7l
MPhQXXS84bWteEJ9DQjSRgeC0B36UFCZJla/PdMAPCQjW5DmW+La2+hfuyct3eyiWsxOor7ngirp
47Wq30pazzoMVy8KoB5a3Cv8UokzzoC/g7ZpPcIOmlpheENrsNi17EUuwXp1U7bgISSKK+3w1lDD
0yRCItnq9QQf4A+D2rhs9d1JkrXzj2OlGOoIUXY3690rqtbYrqF9QO1pV6CLOTlfW2jX/HgNV7f7
QMlpvZSkvockoRPa1R6tCjKFlt1L4GxDFXP+WKRUOJZJkClTL0rUy0El59eBZTbq/SZNiH7ibn9I
zbxchDwqiCnAxnvpSRctD7KNsXQ5mOwpzjHjrB+oSAI+Or/NY3rB5LSYpAFhfS7HK07KjSc2HmF8
dR57buGsRum+qLLwgHuyxmvo6TPm+uYM2Cz4ha5tAWlxCEa6sjXPSUHCPbdubKfta4il+owl1PxM
IQnBQnyBdW6LcBsBZoACrXGee9zDWs9ntJk+jzl9kzvgNjI28t2JAWCCoYkLhKgAgIle5EAwsaSw
T8ywBE5h/AH9AOx3pfOFlvN3LIqTFdLJYL7mjDOneAFM+D1fHB0/MRNaf96rHF2tHy5uUBawg9dn
voc00+VuaOMyVgoWmx6yAvUx7vvVT8CQ3Mun1nSOe77qXAEeSFSQvHRyMPG6ziR+di9Vcm3UIqFe
NjLd0donj7N/13vdR24kGmzFhlGI88qCDej3+2VTvaYkQbOREqCTBbGmh4aol5xi+LnfQgmL8yiK
tQYHu/LQ/4d4vnUMNjd5QJ/MejDrvBM9XKL4pHn/h0jPBrYoqYU54pu2d20SRmBDFKNaO9wp7VVz
vcVBtDSU0EEQ0I+3rA/frAzP7e1OPKYXy/onPIQF0nXq5dgULcs8jxHLIb2EH7jI1nl60/X7X/1V
sNrhmxhy6Wr6DEpWQ32jm7hbSA5H7/S06gVNhMdroVipz6ymZdS5MhUmV/ip2OGUCLEjT4NP4YdQ
59d4mbLoN1qpYUKIzSvuKCUfSc+fmvYB1PMJRFLiDhccH0dFFkE322ve3XXuuBZ+SiTyhSpgO96P
PEJNkjvo7tTe9S9wIuepyfOZ23tOvtgbYD17OBZ5R4cHOYI+bca+4XMDuBFal9UboiDjVtfJjoRu
06OuWHYtprcymLSj6kMvncABCAWqX1sOj3EDxWm+Sp2u5Yii4KQg6O6HvPIN2SiIHkwuIh9nTaNx
BW0cOtYoxOy9OloUGUFQkIkPLMRqlahcupUMoKwXDjnkRrfaSlHvRCW0tvLWVCDmjbT8Fd4/teyy
UodQRcxCxQ9myoshPIfM2ERMXB8l6pMZVi5Zs6ZTr6HABuJjRnpimz6AALGO2ZjPgyM5bQTXsfKl
51oapyrh8LRSMxLtbsCtVoNmvnpxXWbq2IwtaQ0ZDs0d1utNvq5EqHYs9Wt74kHy+PEB5oPdz2dA
/cTf1CuVL3naSEsxPkqnH/BlsAP/LVaPoS4PLXZB6NEjQ7ki3Yx8xukgIzDQVv0/2H5lmeBadm3Q
ylwlZxDpu6dj6TJNjFv3Ch+1Nus7tshNZ6/X19EWHFhYlGuA6UnFYLEoxK9UUiv9UthTuoR93Wgn
7ymtbuWNebUTG68VQOWEmckJjgMTPROrERwuEtYXtwu00ExhZIT5OeWwk40zvuaTAnlpRGMzalQZ
uvbNQ0HfKnrJlUsnlTsluQ2/WHa8LZKnmDF4jJEVTLynGaVKhFoxCbv9rI+11JMN1aJt5F5mh2RV
QIU19SCMiiFcfym5C8BzI7EE0x+weyxSSk6gPc4eavWgAGT04p/2oPJD9AnrARGmQhIBzphlycBm
FmLwhmusQEQnYXCRBFsQ5PBs4xmiSk4OEQ82iCrzvRI+J4+MDmnK4upPptJQ+SZBxv0aSzP7Cz2l
HRsSPVGmdHqSfDBzSrFkNud4spLL/yCMHEY4AJv+MF6bppsLqNF66jfmyGuCodTHaumVnP3WknRi
B1+YbfbL0/ljg7jRy5jGzNmzN2IwdD3RPtVzW6rrRjVC9SyzPkrtntYmCIrJ/NmRnTlFUnQm6a/h
BvJSgbairvjk8SDOJLFZkEh19sYd5/F+3xpOIIqgSADm5KmxjMvxzaEEC1A+0w+dO7blMWcNPKfm
V9H4A4402xr7GYmoN4AN1UC5aViro9cRgDlq4kImApFNpOxAmkAtOZFaeZjvLvNKN/izM2NVRxZV
xBj+rii0HT9vgjAHjrPhn617RKi/yJf384HBglHL/IWPxHDDZMx3lXEJvoRAMuvIW3ff+EABJ9oE
lQIqZfanUwc7dVUkZtoY054rmaU/Nn1fONwHvGAkPuONOJQYNkuazPoAyOy22auwJKwQSuKOSoW7
OBmN0Sure48c54tKWKAsNFY73vNFZ/iJQghXOPd5AKNXEcn6e1ev3myxLg2fiDjENP6h9m+R8tn3
BnxOWprChBclBDXh1U/juXxvvaXaNiUKJ+fz08jMQ7hOA4y2Zlw5GXDY7Mk+Ibs27ANg6k89sX5d
qoyGUiaMtZSMQ+jC6yDak7AT1dLtEYDy3sek31IB5qKgpgumvIMCHYK2GqrMe2E3SmznW1ZZLTtt
7xVcxyACy23tS/v7wNYZKlLLoSs8aPZXVjeDn4y7j8Gj0PnAkVQ18+rDWVbE5Q7C+kaNkqKBzyyy
xiw8viXBxJiRwX650xiw57cVfYD3oknOH++YYGMEzOm2+w0x+FXZtgwsFrfUuh1BCbT03bun/cCL
hzRjMmsAkeg35bw3+bdZf+IuWEZq2dJy/mD3XRtIC2GZqWDiitNnkgkSPfiRGEayVG/ciqY0UUH9
k8ZJfa7gwkyiCXR9jh9+dvgnDZGYHPV3uA1u/NA4pwVR0y4tSzHLmDJl+rzBCoW3BcMooguNZx1u
rbaGpyTobljmf3F4nWM4hplzwgrD7GWH3o0E6shHJUkJik03fX3gEHGE4dlhfmYvg1hW/fnJNndw
gN7QL+p/+be6nx0O+iGTPTE7loqxC7eAx1DeBsn4/eY1oHdvAhR97k3focY74CncdObrAPElAZEl
9lNs+P+8ymtYL2ofcVWqqFW45ik1CmU1U/VcthpxoNH27O0LMBk1jLbZZ5qgsytZtrWC8HgaDKnc
X3hGduMg7oUx8AlV0qLRDra7w1YFhSz9VgQxNsAUzQ40Km3IJ+cAouR41Ozqm417/O4OYhnKQlqJ
Y0q/V8ba4SJgd8Opz2JEd8Nb2zqW9UXKLi0KD6RTkb+MNdvR64KOtl0ys68w4RDvG6pZiUnmOOma
jEcrFKbGzMnYMjKgWQuITlr9e5oz9e/QDhbta5a8ESHmjz2xygC7apr5aJ+7Kj+lnYFz5kyNYU7a
bZrwIveKi9QbgmrvkEaNF30Of6RQl365krZW7mFDw5OHUSQ0bUtaaov0EMmJlAmuNoC0NMszP9yt
m9Carb9+4msnOSBR6C3Z4RzAxkWatfgenVV/8GSkS1pnCcrEiXA+/yaC+vOL5fCJmenH9kehEjfp
uXxY3wLK4UEJXocnRZ5VDGZ+hXreCKYi8tSmNST+te7IAjjC/qH911GXut45bfSfGcp3RfkBZEbh
4lMHCl6LWNxKNn0lRCWG/7HmiI3PVpeb6J+lgCW5A3OEIpQ7ncfh9U5qbHSVtUf69aSZ0uM7oE3m
o6uHy111hDGIKkmC8Ghp8A/LqC8imHLvUyrZqS4kTovyGW/asy4POM0kg6YKfrvn0PhiIr06yccE
uJUwDuC6SE6MglG9eos9KtUac/Erz3hmnCG2hMgKWXrhXR80q0hqCziHuLL4FY66AaHLp1hhjwbQ
VVo0UXD4sF4l8uXs2chCiQjHJ7AxhuxVr7nAaNMpKn95sFvVIxBOOprJDKVCVPJBDUo/AWDUDXKL
2yTwrXWAdGMgttw5jnPiBp2EZgR3DQGcwbkbUJdenHQ63/D2mKb6GO/7GezfiuYnwBoktYVrLqNB
s3A3k102VbvVnuGkfw7k1xjUVRcRv6dJZKHRRsk/BeK5CheAQ44KL7T8CwEHQflIYS6qts7HdY/2
fGkE60247yoE6ZZKHr/ZMWEkJi4m5oA1vSvCOBSRDGUjM35jaPOVKQ8F6WaK/w1/mPDIQYDa2W/g
Oj9a/b7K1eMXlv4h9ZYTBRP44+FI12e1BQ1h+xE3UshXBYv8pfJnmhAoW7AD3jzJM6cdRM/YCcnK
CQ/YGKzihx8AqrwctvY9/A/BAXsQGVTwwKa/9kM4HmYy+X5CxSmkHMW0d4xqbE8kTpSAyuQwCoEG
p7NMuLpjkaGMZuNt+xZ+KHKJIcm19nWDKK+gbAsZJUr9LhBPOfca+dyEz+3pmbuRxlMx2cTAC6ya
V0GB59d5Zsbwq2kjkGhdyigir38mpI8zj0hZmfYZDOPYv+1XldUK7jQQe5zWwuG5DnCAnlRjKmPI
Ems5miCglLAmp0ybsUQxT7X9c2KcKhaTtzJq/ec3i5UkxliRR/FT02juuFNkOnA4V0BxJ0PFxQl6
4/+E77CYpvq6scOlGUDR56XKNcW0a3dmJmZ47V3RQe161vNhRhuDUuzfv0cVvy6e9YsnZJSxhT43
GYBZUmxIu5KxeUSSPli3MO2zr+fxiQLHkKYOsUeoeFj+rOTYuyWyoVwqQLlwcmwUrLQ8puaHGjl+
37L6qlSKmpmHSr+4fpHlT/dj6fCYWSKk54OJ7qkrQk7fcuffLGy7aHrgmtqqMubCAASsYlfqvi+r
jORNS/stePHs4SSjHHNguclDTTbZhuLFuTeHFlQwK4RYkxCP4RCZNmntXBvV4o51XCHP20zvIW1o
S9YWdnG6MK8TQlR4UPDq2dR63UncCitjivWF5xRY7/LUmMaf5YM3wq/QqqkCCvCIwmFjZXh459TR
WUJNlewiJMFVMF3DBR9GQJ4dwH6u5HSiAoMekeRLqFnv7j9x63wNHYPFqrewiXKPZWioDr3foccs
rTEof20uD0piDXy7+BcYyub4FMfRGKJvxR0Gb2TUP5UAV5Jz3k6dHo7cNdjCwWzEIDtMJ8xxDFve
r0blv58lG4ksDatrCXM+kLJMQQM/bzqF8TreuaFjN4oM11J2r/0sXPZ4dMua1oc43Ic6oqL5Nd8F
cw4UD8vqWfF5iJ+2dkZde+zj2wWFMPezRbrLrif2sEMnCtVe0uQTsbZeBU/dvEP0D0n2jq+ytJjI
hqRaDABalu7HWfw0NvC0y7LbgwIF7szqPFWZMhqRjhhVrC613VkJ1BjNQf5A4XQi566oyafagyEF
XLx2pocKn+hJUNE482YHUtmGTXdE8fNO2l9iJsOoapwIEBXQ0LlaDmxyisaF0GwRWkbzSRHeEdX+
jViZP4yhJAqFYNn15xMCSabcZleZbobaIXNKC4SMweSBNHN3tlVIXgJYbh9whCFbtZx7LkCAQfaJ
FtFvhJ08A8Bn5yOLtvm5lZoA1cZdlYuhNCK8LVdSWkoVlyipA7UA7W/Cm/7ZRYvG2bGTyOspmWQw
WOCmR4X1qX3XJ6roaIy/qBUhlz9lXHUqNPhtzS5hBHz68HkSmSJGvWXKTLxBr78RCc1BCK5bwL12
c7EeSlh6VTC6cSgShQ9GdugpI1SRr0lHEnbeoe9e8QiS308tmv+NWYbaZA8n69uI3qU5OK1pJ0lP
Vy/JEKIYhX1uzKBtjaDKeQ4HeIU55Y55PpBG+cORUyMvsq8tzTpOfuf1AQqRYMIT5shicUbeO3eZ
bo9JXTadIBa5viAuCmAb3kKz0eNTGp9k4Dqrb8kOTZLdokd3jYlzJWx95PRW6cTze9aUOVgwqbw8
1sHp0KckX1y+8C1k1yyXbaKfcfhGsN8jw+jC31ykwhgR+aNi+QVTb8I4vPH5n0bCWW2mLooSCjf7
GOXk88WZbsbaPpdergp5GGyzZ4xZfeb7Xpw/27Pa6cg2hBdcCHFzQheS6MZh/heT3c1OsFv/yb0h
TiBwaL3A3B/EbXXusKHpbjQxcN110VnSj/fvBDzhBz4JXCbtylMqupZqJ7xRCsZfTvLVCtyt6hro
x3yNnlaDYe/VozkpE2YFHlLvV3+rsS133u7l+UUUfPSxhgRCmBgXON6YS3sGkL6qJytfLuCtVW1f
5Qtf+Tq3JA9udtW8gws1E/o/lhuoulzLWVkiDqF9OaUs6tB96PCUua6ABUVv+6spVBWSdL/DaAjq
PTEXZJR47Rgs5cQVWOYIL4Nn2Am8VrRivSwAekE5T08ABGjxvztvSdmhjjYZmSRtcmxqP5wHduZh
YLwLTXiiy1Ey0qvmhgqTIQPoepwUX9LABGKkbk+pk4HtZtejUdTVT1uC9OB/Wlebk9Fr1/zWXxGJ
3UQrnj+PpOssz3PovVE3RpQzhzYIBhIWMQjfN4U8LnGJX9QTq6FHmy2WTUSz0qEGB/w24jpWO7nv
3J6dBV0VxCD/0i5EzkZErWr00nDaulrQwEsdJMmXCgjKfTeGsEaxGEvpCXTbxZX01MiIemxPArON
IeLhLjE/+AVt8PPsoma7pBkx15RZK8dagOxohSB8zZpxlBSk0FfDlPdWRX72pkzwzkolpRJQFxLV
klxQlggpx+c3bdIDmRL9LJJdYNzIjUIbhjv5TR4vYA+s3pb5Vgpur9uNR2OToCgafrNY21m6EFCg
xhyUvuRXaxrMJRwptuT3BpPRLnudkW/Ok7ZwQssafsuhzzYhARg8n2Neg3ASxFZorPVT2T0F4DG7
mSfgI5dgeok52J+siesqHfjHDlIT/q+J8kQB0ZbP7aYCmK/b6thfKarOE49Fulafr12zVP1zoDN/
c0aReO+P0nL8Bsn6cQxvqhAV2A9FcM7jF5B4wvBmrQtAqXAVuaFPe9UbXu6E2PAATL5JwcwJeBIq
fwiKxh2li4b7q0zWkRkt4v7hDQcAQlKyisdFuRXstjvkN8XnTPWlxOTYHSq6X703gNUBiwZtRcS9
pW7DRCcn0cAd7E3gjULmQLHNz/nQPIewIbpRe31QUj52iIizyDHPUEo9P9XCU1Sfzlaqm2WXdX96
2+AJQCJWZPyfW6R7+RY9my2eJFVICwTTtQhJnbsfA0HjkxAxzI+VQCvtaHi1SmYDTzJ/bcqXh4AZ
HxcnNn6UIWXxXk0BqPQf0hFCUMOhK9CpduyDcM0+EnqOvJzmOb0gGZ57l2XMYD1tyxNK/LqkX5iQ
UWXJATxAF5JfbpfrINLfMLtxLe3Q/wo0M7R2sj/MCpeRPBV4lzKc/d+E5h+D4vr3455vHVgUa/Kh
FVmoUcVANzAl50UC4K9v+Iwb/xQ7OZVHG3dgFYlH8L+1Dc3N81/US9oyw4fTARVIHwcv9EqWJE2U
FkrOwBb8KW74JocRf4+hgpHiwu3V38wzq1p/fhKs7woPdDgPou1a43XVDDNX2iNvOyaFXhBoXue/
4rpO33yOvUJuWFHAkd35jJqC6mqdDgmY/yWdWUKVCsO2AeNHN7qCw4oKRRD0z07ko/3U+Gfdp+nc
lqd30TegcP0HgvlSUQ0kekpuDrtydjlOG91Sv64u9fTup/8APtXHJmzLHA+pvCtcZdWTcM2jQzKc
bM2qG0ssFdAmrbIJLFm/zIPK+azfdbRkcmBt/MdHFyTjvA9GDtl0V7satSviPfya7bvS1shwHnI5
Hg/0VBsP1olAvX35H2dfRgXQF3VgeyD5GHdtpUrDZfIS1pxS8k7Ic6iGEHh9o9ugt52CARXT+AEs
TkBnye8S8xfzkfEE6e4Cbd36RdmLiQAjU3DxT/xxRoulAO5+IcX2E15AsuPfGTk90HaZndbFBwgA
3YoZ2iB00DmHMOHc3XDdO5PbliptkvUCHnNfnk78/dRpvv6jB2v4ZdI1p4uDqrEQCsRoWyNkMB05
w5ekEFEImgnLXS0PVcP+KB99okssOwUEGv8BKIwC3Qb0MKVpink9qtKXuNuxNnn6U1HBWHT3WDMN
a1/Ugf6kXJOWiOj5nmZ5JaDpsp1De1AmsfnqGaTqzGnsHeovtQCGD+5m6GPSZdaZ2aMyjO8GWNi+
4KSnawVQir98c0rhnVXYXpyLsO9C5oOm27H9CeOexd3ciSeSmU98fFQqcWuRleIsPwIx07rcYFSp
IHtCTMiKdrKsj70+XADh74HUgm2iObeF1I+x5tvek0JU4QBbInr5uawxzMakUGK7aAxjaE+oTwjV
IWJ5QHH1Xwovc+d7MRhUhLAku1aGKUiCkTxp7Q0sU9imOdc/Btrg4PE5Ek0Kg1jlQXbFRAEgrAJT
IC4+teg6qmCHExq+ru1rDy3+iMVKRIhYdrWx+kvOmDgHorqWJbLnbmRy4bytWbVmNUCBWr01DFoW
3Hd2WcCLO1GYz0F/L5JtHM9f/wd+bHwthyEX1GRkzwh0FSY0sTlBF/P5q22qmE+iSVPChOQtqz7v
riekjg1VuKkOPIxeuRmoZ6GkJGEkmLXOdYJSd5Y3mVdWmihlQ2H1KnZg+LpuVYem4Jt2w5e9QRQ5
X7mcTXUZQeKyOCCGOfwNziKJXFUmLNnBm5Ign27h1jXHqLSoBK1wDidD9fYvHsJam9iB4yEQ9Cv9
pmgG82mY0Zu8DvfDQNroGQGAZcD8E56kAKKy2LLoI4A9dpIyOEkPMqOKnIUbGl7RPF9tLGtxM1vf
s4l+ykC92Cc7lVOpRmLMMug/QxeWt8OWw7oQ5+qfsWl99xZgKDQ9CgSBYOFnkwkcPX4ckMh/FblJ
wd2nuxv4Y3C2mtDEu2E0ZWmib6RzUHkzBoqOSIVdsBRrGTlM7msv07XPpKBnUYFT6q4gAmZrKJ/A
FCMF3oFtkkA7Km1mkeDIM147gTlnPDmvxh68PfBDyFCzly0Nam0BjsB0m9TBd3Ts1qlwTPfMgxqn
ohXN7462yK0Wk4s4jl6T2Jg1zqzX7SIc8Z/EtJfT1olxeUpAAPRtLOIOLdBFNThkyVDbcZFKpMQj
PS8v7gbHmg9vcYZ9VM/eiRzDp9R4UjtYpmOjS0CML4Kast+NMJcJW+PM12kxJebPltOmpU1HnJGH
R5Dl7tKI5ZO3A8nBIJAi3p46enO6WhIVYd49z31zO05cbUrCRlzKaMb+P0T8rJ/IOI0Qhh6B6oon
lZiPioHEFpOHum4B7WCrMre3Zdwe6zokeDbT3xOZ9ajD79wM+MKdlNZoUJhK/R0UaOYcMxttZO2z
zNR72xnC18UV7J1xbdHqY6h5lyBF8xIH97z33/f8Jy8K8WTwBqM1+6gTIeRjlPfzwmMWviIC3NSB
AzYa9gOBiXotX8ZxqVYiGHrIAFeypD3N3wotgLkaQ1xEQEds7wWc50TKn3fGJDFuacIwE51A29nI
nvFZRvFD+7LNhDPhRZ2eeRlgGRfP23gPRILMU4bihOt9VyNzx3WspusUOZWH2cajhjN7eaNtg/8Y
cELw2WTrkpapLMNbLG65gkxXs3bYjE23MX7CGTGNadCxDDAaGhlYwAatrlBkL70J4/3/hM9NVPC1
lZ8pkXXwzNYzdbUsWbPijt+d6nwz894WMA400iSk0YOIlYbkhchua/uJKdk5VleJKtXU744+1yX5
ctcwMUhPfTv5PlJM7JDixwD/HgjcY7dSLCicEC0Z8KX2UvGRD7dGOUutLliMy/+pMQcuhl1jP1VI
oFavHo1VmrASPkxn/qEzTwkYjU3iXzkQnCqr56huhJzZx9KdC5ebyuTOVp+B9ass9u9cZQJtoM2I
wpd17AiyiqceL+Tlr99eA21NMAvHhwDEbomVlshjmGBeKJUIcOSHo7m/m5RK3Q1XOTuW8C1pvsBk
tgdDQDS50J9PfGiby2GYoLfWlTjTQkQdFlLi0Fg28sXY8V6qNg0m6yEyc/ZmWWUVRETL1Di7nbcL
+9eRc2RX+PZVBAKPc5iJkRl9xexJ+AuyWmPUquh21Csws9hBMM90CFccywNrtHYONUwaZTcYimKU
gRBRA1O+Z4RfKpro9iCIehJLVDX3F81vi1YACrNzblAsr3i0u2WMf1+vRjnJxY2n2MzEKheDVN+/
Ayclt7G/3iYkyfpQ3NSFJE2yQ3idr6z8TRS+xwj/+2z5Yvkt45XsxzpggQ6080y/Rdu098a4RFNY
vcV/K/xUUNxwwnav6Qsz8TNE+qvwhwL3VglFNtGLf879YjKgL9kyCb5jRYF/RImvQxBLNkefgCST
PRdX0FwDgjnGoQqrQcNkhvXbeP2LmeX7wJ/A9BbE/RZvjvkmvhsgumq+qAu5qkCLSkbjF850EgMt
AkTZLsS6npdu5hsc9CoLoq2XjwSWJV+6JuTvlc6zcU+cRhEnJ8VoRX5DmXf3fvd0wlIYWJq5hGYp
EXnKqx/XD+a7dJ87oRvZrgEgXjDSQTFZN+jMewosZCSq2kAipTv8GWm66otGTwNpP92FS+xKMHep
IyevoeapCJhtYCl+tImkktS/iqWFPmHMVg7Cj2/aWflMYlAMx7bzspYXbzJpZkCcoZyzqeLvPvbL
qzGgnWQMuAx8XkBAgJJ6ZThFwF4njsJlAZg9LTJp2MhaRSG/rK0RVmg5QHhgRJt8iO2gunYkJINd
Ddqq9RjolRmlArILO8g7nfg42qUnbJzEeJZtFp5x+emY1gCaOZb69b1Ne1T7Yz8agUGOsxunq0MK
lOWHrO8noR4/NG/+sflko0dpWkL3dHoWKmaiftFQojdP4zZq/t58elKI9vgqOOxuh67g575V0Gg2
x2jyHhcP2fnMWYaMSGX4+YHYhUP2sDqjL57MPHFlz7LFa8/TD52Gzn7Q0HJ3wh48Sxlt89M21eil
/X9wkwAJWrB7ZrW8tF5Sni1jdN0fydZ/H8m6utd+Weys4GA+XmCNLGfktcx07SGzi56K9G5Mba01
CRthKr3vB5/UBwoTd2QLotq2T6EhsHakuta1LgEzm3TNON+FeNHnFBq3CLA6IBBp/7qyDpQrfPg9
jm2L3vod5lWz0wcQb39v9t5IgP0kxlutkyp0yqSAl8zlVosCPnU7CYvIWJG+5Wj+AJ4E4ZZcK3j8
06ejjVW6wUrkWBaBWazLEe2VAZ/TUmN5R6uUU36DRiWVyaNYyJI/JMKy4US9u3z5UfOAnvjshNX9
m13IVAQjCKqhV6AuSmOTEtWLEKZEJ3IWFzQ51keDezPptfEL2Vb7QHueepTL7ytZ45nDBw1FrQvA
P8o2gG/0xIHm0lrhqtYkg2S2yCqeFZUGn9YJlwl4A7DCHq8ZHU22W3yS94aQJuqTzWPHIfPIGC/x
4XPSE0KrCpFuB6F30VpL6qlmMHa3qpkI2tY0yux9E4ZXclgbuVeySD+7u+X5N4a/hh+s5GeYLo99
HQ46afZsbz9BNbjStjJPDB4MVVaMLKTM2MiohnDoyWxhIMLgTtVFg9xDMvOW/Wa8OHLQppWqwcRy
Nh9FmY7Xyobs56GZnzLE0VG3eHtm+1XGSmEthjvcQ0ZQcH/xbinB9DlWCiqbeSg++xJXcg83rvJC
fVV9A4RCs8jkX5RtRMT0j42WVt0LyrcGs4dxVyHbcMeRPPxSDc1OLcO4gmfAGwD6wIfYAWucRJnw
TtDodbpXsk0l3VeK6vfOy6tp40ImGJ8CXTQiMpUmF1u99PdSzshSF2b/N2mnCHE+dC+vzJd6S6QR
YCxagQUc1FJLypMNglMsUSeLwiNk8vxUvUtpI15ExCggzWCDSYOVwr/ArvddACV+malYCtHIZKwb
M5/OI3cMGUmc4NqvdJlNI6QlFTshZCD1C5D6skMt7VV0Bji1m+oK6Ag6/istT/w2SAMzgzeNPuYz
ZcwgB+zPiAlj6AN14q8R5DTMwYUTGN2tvJGBtJzHg4bsfefKgrOoMuMVMk4l2tt2uOJ6d0z1Bd/o
hoT8j0oM5rtIsM7G6Ztv3BSrUI0h9uagBmiiLWqkhmM2hH2ZZFZkww+bfPsLLA+AAV12DUYEyuVz
lxu3e/lBceqt4jPNnED3B9OtRaA7yhO81LJI+p4I1EtLARo93hgbavC9IFsYMuClaG55RFgDhvw9
/bIk/gxoTBw8f0mcKcPcgk6wJHycOGw6UL4te4o1upOr2rmlePCoHClfAvd31zPqotlF/xVe3aLw
qxM+Uf0hDuEga9mo0d2hdkkJdiXKjPczXju4EvmQ+xe+E2dnQbZmEt9jR/CsGopck4Uu8we6FI3c
R7LG/I6krtE8twjHF18WQ7ZNlEx1r7tMKdl/VktmGG7XIn4jRNyXGj1RXFF41RHvrjxk8WAhqqBh
YRS5uK7a8bm955g2jkyqxdCnLj0ELn0YOjfeSEBcUdB3GH3gSAbCnxs401Fcq4LeXbUoXzMf1Yjm
qHncAt/5ge8yUiQF40xIGdlnAv/7ZcOZNb9Up4y6X/pLmXCu9wyzE2w0FvTDcb7WaD6xhz1+wIMP
+Q1kc/bMWnpWNxXHtxanZVFYNkwKa55fp2QV8dGSZmOZagYuqY4fSZjv9wWeWj/BZDogYFb7rRLp
Oa9tRORY1ZiuFDKdOXs/UUuY8wbuqyo26iK3wfRgl9J4sXUQY+JQY0/0jAyBz5LIyPGGAYM20ijn
Ddd3M9PR4YOEycbboKEyC9qMKWcGvJIZbd55NolJWwj073e6DhdpVTgWGXCxX2BfKQ6ZBa8/joyD
DSjh3xL7SUTGMD6duOUfVzIspV46kujp9omBvT2l2OMdQt4pJw8eqgZ3OIkDuV52mjpP6IBvoV9L
PQhx/8cD+veszH2etiKSBq3dbqK1lp1QyDx8J1oe1PqCxTGV6sFGPi7HS2lqg1IbGRZSGEK1iJh6
GI6Nd5SRvK95GQpVzQWTCuIKapD3A23bKEetOJBquZIEpUU7/xdD03MhavDyMnoWJsYX0/Z4e1GK
+4KERdN1q/B/9g/JE+5ffFIEQd8FmZH5iYiW0Wb4pGOcCE97ipUxltVZWicJqKppCCs4JAE+hkwX
jMHTBOPAVZxqurtzdZVoPDUk+vghXfzNS0nZI7mr2EalNYlisi9Yi84OaokpOB+TfY5aVBCnY3lC
8b+Kr63uVKcq6BHSyucn0jzcOSbkxs7HPuNBMM1yXpnplAUjfvm7Oz+gY/HD8WFCV3I+thGqdTpc
Tup723YyODCsixf73Q7vWuuutQYntsROCM8h9c2JfYk8IsiE0vsv6GvjBBhWRMu7RkZI3Bf966el
9uwq4XRrdWlYiwn+Dz/QdhmiIjtBWKzK+PJe9r2cskioKcP2L/pEC59vXs/KpVOSYzsZvtm10Ufk
EB1cQEQReCmR0hFrd4LNKKHD5BIonqW/XOxm2R2QEWpGojfS/22UA0Ncw7kb9QOmZvTHmG5sJCFC
nc5h1+HXoTRuFSKFrqKj+e+k38gUoipPz1FwJpevRKmoIT06sAmigYOH/3oNDoI82DT0cu6tfqIN
ot2CYCSWbMVg0HO7ar4S5lSJXVeoBg8511ieeELTm2dPlv0wFdSqvOQvmiEzwW2cz4MtvjdZ2Qu0
mdp3v0Uc7A9BD78udanVyVziF8lWLkPHncDexBJrL13C1KL3OhK5zzfuEAElEf9lplrA8KoShE1c
pEaM7glHfjINJFOr4e1HsVknGC4DRu8AeT5iNOAr/JJqPyoWRcWMQVHHLMkPaJQRZwWds+4qjOtm
O+sTsubAskdJr9Bt2ufWGZIjfQsvo4LPgC7u7ADxo6Zlnn0Uonuy14IKT7T6NOQmmmbNXsBCfGyq
KQb3WcPfIJK1PM/ACvV7zLrrX2sbX8M458cP6orksntCR0rWDUKAWON3fLu1RfLkolWDJMUoqGY6
ynTtACWVkYdhrlKrgn3/dOQcpRLdq5vgwF9RuroeuweaAaKxoQi19Y2gs4u6uLBordu0ldS63n5O
hwKZkAbDYbCcc/F17ejQUa3zH6QthYHEPqH8xblD6wjNp3f8U1YLpSJdYm9pfDBHehzOU0vS7v9b
v/Ieyw2S/luwd5juozYKKm0ARdLDlulJsOgQT6IQvxP06640YpSA9mA59w1DbMrHNuGMq4GuyHfq
zXvPhTcXQd2zHoICfqAzh/szk3gqQA5AUolJAqMlfo4nhQmLfvmjcRn1j35sLlAbecn1ela21A1i
JoXdTzD0ixAYpbhHU+3e+ul9/Eeh+Arr7kdGdbW/rhQdRX8xZ+ZzgIBCXtDeo/eoMNUv0gt2vh5Q
+7zWDP/EJcMYetOPlHk+RVSnbf11KSpjRp6+RmjQE16E/OIJf7ktcipgT3sSsSda1X3Cfv/SnNni
N9CJfSHMtiRpGjwkelwy9o3HdIf9N9sbBlwJ43MheWmpJeickhOsbnIOojLr4r7dyvSCWQRtoB4B
3N27RWS/jHBfSmhlfw2GRugKZIEM3tO5CyX88WurMAAEdmqQHhAk8BeeAIubT0vUHJIUnhoP1Nvb
g1zBB+EO5CroAqz5CLlHPRRayFdUmFcQXjqCjFygtVeBCoDXGNIpMvk42itK7Oh0v4WduadCXG2U
yP75ejyOFJVRDP0ZRdoO8P/b+BZC0PQrLi7d4D2hX1AMiSRYIRwEAuRO0KlfxiIa7QT+JSa0jF6O
n5fAHOUd4oMsue3OiJUERfLtcIQ7uWWFoWsTUJ6V1VMaeh6PJouZ3OkO28rQNdZUBzo8xMiLQCT5
GHbc67nebQ0rbhThwEeYgBG6byFKPLSB6v2Yn/1H0LJ+oN0PjYscMP4xrWlzhoiVGnncznmwzyUV
Ry1+BZTcQE02fgS6/OdAT6DYeZdHg9uBdmZKfnJtHKt2bgB95qSgB5Yl2pNAyjh4gxFTcsyHay9r
ITqCCYAsdtYfTza4ctrvk5Pn4avNO3Hd5s8J79pUvmwrZ2fV6ANvmnpM1rWj5IQouOYjLm5E8gjg
/cpoMZrIK2E5c1Gi6+QnIQlqW9guJcmUeGv5+9MkXLq2wQwJtT54iSxU+rEquLdQJ2SutdnfGiUr
UtdScdPHFFh86LhezHjBnk3zaQQXhxM0mZ9atrQrDgi7XEw6WgZXgFmyt2FtH2fheU+KtrC03Klr
cVgmlYl6n1M3b5oPVWoXdmZwRHDFW5cs+dyyls6aSCORM+4iSM4DqiThqzXGeY1wdaMaM/Q4c/oy
aJrtd3qHsu5EUevWA6X3avFgRnF7UiioU033TPo2JhI6qyi0XNM+GepbcKBjFCV+fRsIIYIuISkm
nB2zYrTRQuwiaObFfPZ1t6Hd+YqTUZmzY+3/rKkBmYNfNEbU2d/qUjOumYiKPMFNr+2VVh3bliRr
XDwTkQ9pI2m6IDlhJSbI1jFM2ZdB+miC4kDcN2bP7S4BVrRogUMBOHPhPkJ3EOCqHaGBHeTrf+IC
uj0eZ/RPHydn0J8uujuXdAFebbKE4ZThK+wdySeCiXjLRNf4woAiQiiY495cpXpQ+1Su5UjC4Hkq
cZ5yPTinZ3r9UXjbfD2khIPpKxfktQr5MEWSKWNGMRh9wYDdHphZBBtdszmVn1pYN4GtcQcmXVpK
7K4PMeW7TSR/Tuqcs4nap7Q/HSikFzPn4m2ajV8Obh+DzcuYVykTZ7bgZJ6THOQ0IwgTXCwsd4uB
in9VKJ2Tjng+b8cRWeM6VKPAu6VYkrIt76SxGb4RsUUUw7DwUZzmtktTQBTTrZtnrmRSuo3NY2D9
CchiadF3ovXR50jDECgXdFwVme/vlecgOkCnlG44Q27tgHRf1TDN94ljDmTtXnwHVrFiqn6lm56t
1NBmu/R0jHjxLbTkoi+dsbggHsFMoRhRgi1YCA67uE1fNrpZ4ipf0G24dYoKWVZnSbvms9ENGK8g
eDBk5uDtw3xxtWF7YJSYWaHu7d46cecHzcDhC8S8Ym5ErASqvNogk4eRutEdglnA+W4no8Kk5szI
y03sX6UqljwUUsYb0DQUtwgKlikEcqpNhy9z7ifqSsF7SZUpqT4Co7ud3Surfq8OVZ5H9tYgcCOR
Gky+kgFalVoRlSs4vuJdxqX3k9NfgVJ7apJLEgznGkhsTWXq1uaxtLw81/rk/+MaLx9Jp1hC072x
JsBJIGH9+jT6pwa+QLTGV14XubHxqic5H8RDleytLVxeXI7qqJuZyRV7dhb2uxJcWKsVbfbMDu6/
4DxBeJBJ07yAKLrIR1nT/9OD8JSgV3koDv5oNYQIhKU9qEbcg9O7toJAv/HjSrQMGbtvhdt2YYkk
HcTPrI07CtCejDPwQbSfuxZQ81f8sRlFjlKGp4gbEtsXYD7a9Nqn+NfRcs5qbUjPq/sFKhiCdOg9
5+4Vqe3d5SeKuYMyikpKes+cpVV6e0NuwslVE07UTfPffwzkUIDF3e2vjJGgcn53CX05Nb86b4au
abc2ELzQqak+Y2M1xrHcgwCsVqfsbaWXxtvVm0p2h65NZOwxPWTWIjs99Df6tM59IkP84PhJnuLE
iHpjDZr8Iwo9js17jxH+09likZm7C4Sa+uAvvd097e1+9UuE4Zuhn0Ylg95rz/XM4NzNtDtwIzG/
vwCEcVPdCwG8Vv7gcFtHs9/kIf7YBHii2hdvZOZH6uj8RnmscyeW2kjwFJtFNuCiGHiyK/jscr90
3gH0zfoA+4v7iYrgQO3n+zKhEVsTT+8q3msYl8O0S6qY6K5Uvtl803O0tXAYs5kKV+wEL2EnnQZo
+nWK9EqT4ZghsZxrXzssC6lLTfK0VG2s9T7GcLozza2yEkhijWacmakXHuqy9MFdizEfj6dj3xm3
pWWfxUADS3M9oWx1scLbwYB0Yaom5MnooadxR/gguvNEpVFA4uOhRp5WYIPPp30Ew8J1u6Um51al
tXIQS/LQpELtBWMlaSENYTAFcey7KRpet6M9WiUuXKR82VN8G2kZYM9qmbuw/kfn/pw/WFaMBk/S
ud3/Z8p766TLakuDx+RRkayAvVoi9wvjEwdDevEE0HwDa7murLMncqfUEWC5BfneWz3zQ5WMcl/m
QJ/Fs9JTOEMznvvbKhW06db7NQ1k4rA7OeS3VW8VNFSUlOm5PVwAbFuRikR9i0/wPKMiaD4noc5d
wkJWal4F83WnN/GELz/ojeC92azm7nXeiy0okty71aDY1NXQ5Fho4SaYIHBiLMdJC71ZPgygLNdX
BwiCFdctYQhPL5MyVOgoXCBKC0lgziypbmt89CBEYIXjg88/NEFes7YeXLDltK5sIawoDmTg3dVc
hMzl+qd0MZ8MT+b5mlYfWDRq/WZQxievgHmxkjGxYpogMyI8QJVimO7NG2xqY4TxYSX5k5OLVHav
8e73qF1WPTk/4LZ5+3VsWrTi7faZrpQYrOLgvStqK8bM32qfH9aA+CkEDDwAN94emVT0j6zvic+E
SoH6VwKxJuS2CJjor9pzBva/r4wcPybIzP9zoNt0PLBdndt3JddXnpt7xqusotth+YbNo7tuxWzB
D6K8EtgMhUsetY3lrdAZ8PWOaY6OqL3cTJEAyUbwVPtr4YivQDNbhi3Mcr7Y3sJocD1K8dpB0N6Z
IuH67svdhMVFx69N2ZhFaJVD1ySyVEXNbU2LGOA9AnRYrG8RPoNI6ODzpGag6i+UuMelvBZ0xHUa
otTHbW4Iw2DUGzlvQ4KZXTM7SIwXOCviF0ikTWxqpcznOLJiDW74CI+ZABPR55WpVSp2pPAT1WOi
Cw4qZsTavnScPA9pU2RUIq7b73PZc+lW2MwdJf2zwpDPil/wuV9AQ1VJkvvDInJI8AWXCsXCZdlq
10kDfdFwbMkj0l5SKlPLCCeOlPnvQENkpP/ndH9nimm6YtrFlkqRHBormcjssbVveDqK68bTnAH0
cuRJkus8jn5rfCMP0zRTi64zXw8FCv39en9RuovTwEKlAjaVFgkv+TPdKzD/+S2LM/X4y7gn5AG/
XNjGC1M1QA05lCd7uEaD11uAf7KfLxw6Dj4H+y5w8MC87pxfLj9EmoVnY8rtwrNdWFuZfirGsuMn
MfqKC4eQuJEXqWCXlMVwpCf4NaCk9/1E1w4kabuV5KbeEB21j9VZjTmPODPVfX5y0jNIF0kqQS5y
jexCfKMIUgfpECnbQL8jbiRol4zELt7ZwTmbUKvOFod2l5sBFQZA4NlQyzO+fjuzlXWyjBKNNRhT
dQcnMLP82QF/V6nMdS34nhX3s/6JPoLsl+7bV138eyeDlwkUkyFVeRjqYOexXBBxbF3U+zfCQSlx
qKMt74rY6okrn2wEfnZDpALRT9EcyfBvsPeKw5zG3G8IlqObvwUH+y3bhZST0Rg6zO9lHllYM79E
6evGPrPm8flzICzcbOqflC0U11s2TFvGSKlgB+NQkaZUSOEfzLRwEVAToXszelJhlfF8uk55SsJq
QFaL730XoVL6XzvWfflg3i3+CZMo/vNDGzeQ06aJyBSJRrs1uwMYOPNVZD4RAGrK4MQabo8QmiW/
Jc4t1h3M58FZ2m/lQfKM06YS5IW5eWZrysMyZ9lWAuDhmGpGMJVJNjgVw422tBueLGeffGAauSTa
eAWRR8RJtiA7iQbHuUJvW9Ze7IZXbqOKw4E9uqZETl4rG9SEwaAxKHNL73XBW1r/ubFGF1CYR7Rj
pz7nF/XApzY9XJNIOfYSlBxoE+XBxDAgiVQiKfaqRjUGwsqXxzjVeuEW4VMjYX8yqvgBlGYgt/co
N+SBfZz8J/yghDNfxqBJK3zfnce9Ecd+ZYFfEqrJRfpQsJH3fJQ5Y+gUV/3i4MwnVR8ZzmZJ0Boa
SPTdviGkkdwB0icT8kshg0RHVQSUeILnljuwmLOporj7PM5yUyA/bif7zT4RrTvMDMR7b/CmB4w/
aiz1ZR+TCRphE2On39muHXwQEAW+uENtbwY9TjIiSP/PTA6bYJ6JX32A+F/JHRWAWOToUErt0CR5
KrY76OEDZ3RxCk7gBlozvi1UD518c+r67TulBB23R0WWZIY6aKvqKTUyfllPy9C67PrImxhlBCX6
ZHAgNws5S4F2R2co29AO/7t2Zf2oiDJVIpdE4hXMFLR95/lKoE5E4ppJOA/4/pSPd21GY9WkCfRf
Pb89xvbGhbc4MQG/hF3pqbyK+HXHB8SBaMgz+zD2T+Fn3Qww4tnRAniP1+6CFmb1t3vuSC5GRADm
SoJw3nv1cdIWq1VXDc7htXP544FcJYl4VJcgLxM1bBCAcJ24EPdoCpeDTk/0Xcd4C945TBzQXoGE
8wpJuS2HeuFPFKRxh9uv7qfmt62dXj2uCh/0sCT4n1CUv0l3PKRtSj+Svj+1qG3/WbOMzvQyY01z
gDXB+WLQKcCckXDuFzvLspGJepyn/JrvTjbhACmvfEjMnlfzZtlYo99K0wYR8ORNCWWSz1wq14W7
ky/xpSVhNNjBsZlo/tBuMGAkebqo+466baoaw9Mv2iMg7WGuWIFGTRRExWesQPAUwTv0JWsKFoDJ
SQiU1xBhEquBb5CHS/Jf1OiPZO9Tz96rbobVFET26sFDY1OHzurLVJviuG4G0JidAhgFeS3g7cYF
xK8HzZL7XvyJURrlQcW/OosaolPkU1z/xmeanqSgQwSRHMgORzy74NDlGPpDpA6MYgTbMo+lnTl7
aulRI/0N3uHmgXiE0aDOaiqFc6S4+tJDXA0uRq/+El7oNeUbK3PbUNzTwqOptzAmJRbEjFrOwvhD
pjUkXXA0zfiWafYan3JxK/ywXnN2nlz7PYAo/riSnefGHpFF8oZ8JqMy9A4FhNCZBZa+Qyog8jG3
/oWqYHQEQNKW5nzK38lgMvaaMTzIpklPupLuiKRJctPws1JhPJY7QbcvORJ7Cw67UJXoD0QJ74xs
RuaGX4CyMcnylh1IDS+moRaKeJsH6d2pzqg/VZA6uCNXIX69rNIQPACrvVpygg4WRv5SMrxsIah7
qxndqkweVMxQxduUeRda2zW1uoSAcatnvFVjnFzxxPc8/HvvC+hxgE0Eg1dMIMtT/32JKOo/wde7
bmoP+1jhaLoNQqPAoo+2fryWnI/1Tw5+pwgiWNjEh47X9bkl0iNs1jAIbQ2S9ruboloIZlRkKv2P
oAsgf4009OlIxvbLC1rrmmWUVqO7whlekJPa3VBFSde7UJNHm6i6V433lr6VlqH4cugGA7NsDCBu
9BGSBUXifffuY0rrrWHXX+abipD2WDyJrI21yHTMTiE3wr70AjIzLtYb3dP3lR8FHhU9/Y63Tnn8
soA/ySo+fTCcXV+a8CptDRVtFzYbQMsw6CpxKSP50xA21sYxOs7LcihRbh/EaehxRWgDZT+gdtn7
sFX39ACJBeB24pZupPQ9e3Roh9lLSN0lMQHDsM3AQLaX7+rfEDn/Plpov6tUEdayFSH1RKTG3zL5
g8QQuIJKgjI8J4iKEM4y7u8rHFNwvKT9/sb+bynYCSPFJrSrH0u8ljnXL8TzKiuriyi2DZ+HWras
2mUJDeJYvlAQGHz4I05enFP0B658eA6/fu9Ys8PNqbbdX25Lj0uN34TPewpm5t3nlEEGUG3efOFU
UCXSplrrg8PXUEEDqrbGXhVit0fyw/tDVpNLBHfDogAtJgoH0zF3Ts95EbIposeJtuis/3sHEJHs
m4kgzQ/dy50ccnWnuI9e3ELhhclu0VORXaedAsYnTgBkSDYYcfyRDueo/adKXLaUpKpNEd0dA4aO
eLhmubcb++Xv0h7bHZrlVXiRVn84YYErO7DsnRHgEMBe6GCrL9ENWWewKeuoI8pMxMgm+d45DUuI
iWS2JAkEoeVgOvlh34X6OOyGxZhi4NRbBRuOzjyrcXtvOrA60BGd9EPoDG6cJ5BkNy+ELvfx/d22
1h5d17eAFW6yTDs+3QfxC9tsrIJjNYD3lurnsscY5/MnOh3KNKxVKyHw6aWxhtTURnJShQpXadLx
utojxOk4/4XdRPFRxxZhXD4MbWeTrslvyIXi7zpS1d9ZDZQYYUs8XirSV6BzYeFfx1RIVqkl0ioN
DnUNUKLUiIo17kPAWVlL811CZpty9rZbbwi1TXiqaSiModCxMNOY7WNUD7aGUO6LmMpF95LYH2Od
QNbtzaldkFVnU9/2eXalQ80sGUY3J+4dDA3+0y+IOz9mlkTKqvR4Y2f6Cv8O+gtd5JUM6j9D68ku
Lt5nBsmUf3c/kAL5ltDgeuD2PM3oeKzbqjcev/KWrzbw7OzMvJbweWOiS13/8CN3oPlKFq7lYC1q
3U8NLt0Vnr7nS692nGg0agwHfJkj1qAYrU0lyS5zPlp0qSj4UWhKi9EOuWycjtks5XHumHziYZNG
8u7jUOJuKlUyrJ+NfgYbw0EX3oGkUNMmTfu8xQSmT+g18kjZkje93igzJkf17+Ji1ESiCSAjnk0+
JgKr8U1U8AkHB9QrccF2nZoeiP1rh3ZqhuJhvMk9LJlyP9ef06g4CDDUdiCs04Ssxnot6dmG0ZMp
YlAQvNqVaT/pWyCZ+UlobDtGJDksM1Bcm7zfZ35nCr799mW69FjTMc6VU+jFrxLM6X3LjKy9L+3M
FiApJZIo92d90VYiOHfl1ef+DsrdUsrsycQ0NIRCDaRAKYrP6mTxVz/7HTXOmW/1rUYrOzkWhLKp
OxHDP8Uk311hbvmKtq+J08PNdXnPtsLUyE61GRE7h2WKMcYQjy+iG6ShVjunx7d95PcRfSoKf8ni
hwESz5QqkuWTgIbhjvCQUfoOIk+iUZMTB7r35528Mu1EIg2+xWKrIV8PWHm5KYE86WTG+wQ7wVO5
kRq172sDMyBxROAnrQMf4XXwGt49hvloZzh5lgXlncWbQ9JXRTPkFGBSaaWS6Q8cN16tbT+51ZDD
AGAYKcyec15fA/xMBLMNn+8DsU9Hqt00+dT/GgUWC4wmnc6jrw95VAuN6lu0ncxZ2clSk+XzAn8U
acnB86SsPKl3wgmXxKxgwdwhpM0k+pKEcG2KAeamJjGv59F2LtrVDymgIrgp+9zNeZGUSdL6U0La
U75EgfFPFvel5k0ygzZNURUdwYzqqGPoGLUW8cY+mTauuAou4apIrBkLecULhTU+P2OoVUwRtMPn
y7XtLpTGEco4FGPHmAWmuq9rFJ+WI/2FJG9EBWflbMCvQOr1QfmEc4ClDsi9oixv/nUW/cc3Vd37
TgcbON/j+9pvIhAHEJj1/F+UmuWtvoo5ZJROowatNBTODHlfyMs6uFWh+GYi3erPiRwHtH8jzafQ
QgZ+ksnrrYPIG7q1bSaajUr8zqikKwa4xCR7ZP8gzBFOq1WXy8QPB2LFkXJtxx7mo72QVEFHwrgc
NOqCySRuJj+5x7BA7Gd8eo+AI3fQpOuAd3hRvCMgwy6mgcNTeZtogWtcyev7YB8olGOn6h/XGGqQ
PWPn9jOuwaNWDpquBG/yMADCnKupoA/hL83+vAfwxKsUXKtLzsn4VRHWdCAWJDrjfP2Zxng98VCp
FUI77prWr7UOSG4zpVDvm14+MypVrxFa2SGp2oijI1wiPMDB3DXeU38EYuvOrKQdzGlSYMAzkXwm
VV1ySR42aArQ6mxNFP7jbtpasAnQte0ZZ3Mk4YbpGNvaHBsLCr0KHfGz1d2RfbOxmzZ8OHwmG2bq
nbtAjs0ge4p3BYnir4DCFP3JnZKryPofNFUP1XtNrbH4smFuBQpVAUV6OGPFPsCf9qEatBR5J8qi
6Gl+VDFrwfB5tEVK7KRj2M5c+sU4IAkIPwx4dmjTf+ra5JxeVJKz5QGUT3dngk0dyBFfLStUibUg
mP8Wyx/v1goTGE3KlDCsi0Kikq3Ae18fmZB7Gb94vzvaZuZ0GLRK5JtoZ8oKpVZnvVXV08+xPKnl
pqQhBhS+MJTlC1dw/o3OgrTdzR3V8TNMb57MQ9Qyw1Pxr8nwuA6MsePyvBdFumN9B8jS9c6g/1ob
Yzh4wYIkr5JME6Z59nU5uptL7FOAeExslrqyAK/6bTBte1oPtndeu4Uy686vzyIs5nNj2qezFZap
SFfgO9knaWYa1Z2/31ia1lZeWf5zQmTg0+UYH+dUu7wyUkFz+4har9iKp0HiKppHKaquLXW7DVt9
Eyo4SoNjI+lZjmTs8nESIr8sI8wNIWAbsFKW8XteuuROdydvz6IFPzkyezjyEzpc0yPXYzPBU0h8
6hqiCSNXdwuVeXfHGbfvB+DApuK+dHiYCcM4mXEcFlYkiTIq54stzdO5WumavwPIctEfG58aPbE6
88vK6H+K2hp6bcHW3LO3xuZWgDg1TbZ82chjiRgqilWkTZHXp8OOd2dAZBF492KLFWfUd0fUnlng
fK4GD7ed7f5FbWv1AzfLYVVgPzgBe8GbvuNZPxKGMx9UV9wbq58cmm4OOZbira15CjZC0/4QzfDn
fH0C76k7oFT8zYftjoegnf47d5NBHZ8ftaSkhDdxcuQNUCTgxW7J5OebChEmc3FpggrcpP54myKc
81Y4Z15AoCTq233luEgGrgXpImD+DJzJOOkl+DAH1iKsG2fuixoRfLD/tB4rb1FKwk1gfpR0iKic
su99SXhZTqIO4j2MWBNs3t+HLxeOtJWoxsww/CZNuGFkTe0JmDLQ4DaUQuX+DZgjtzE6j8wllmf6
bJ4fSmiFPES1bCdsYEwTO1cyqJ/1QnL20A/ykGP1SLYTow10nLLAn0BC/+/0ODzqKNQaKmkq0CW9
28JUVi7kaTxL5q3sUZImKQiH+3BMR4aUt5m1FCOr7bJOGYXzoCpSBAR9THw2duMdElyRihPviSmo
VjimO7Vz9oy+MpfPQqOihHYr21K3GUlV2HhkiUc+IVT8VgrqHAk/I0O9MkGvzOqGhmlYtHPYWuEu
WXhDkUlBm226LhSsLy/vPRfmqW38yra3IHFBPN9EjO3n1MgqOO+pVWkOF4b11eKql9whV+IjsJ/G
blCOXmBcrpWpPiWqBoJiEXjWCnB642+C+DxyaDpj5oNBzWk+louHRfMX0okOgZMOlwxSpFgt9U1n
l97/9e7uphSCPwugJlCfMFipqRNUQnweYYbpFiQiPh8iy2Ufi7KpC8d+BkpLMYowwEXqpdT/gr8p
VACIh95HVkOFk1UIrUo4h/jRvLYpThxTAOmXv2C6Klxhj6AtHY/0RoxQCDsw+0C72ppM3u9v0LLB
q1xe09EzhHGl+Zd8iz0Ej4twlYYzOhuSch6ZDrFKctH+Pepx5lyLgo71n6sSgb8eZC0LJRbgVzVn
iUU34jNPx6w7tUIDEINlFBv1xc2bJ+0MkLQ/TDcOglB/tcjSVuYJuBW7iAMGFgjlo3J1uNwa7tjH
U+1LLzvTyVDGZgum2/iK31vIs2LUK2XdXfVaJSS9lYyOe6ZDzabwGovoR9rv686IAFz1wKOGhrmZ
2g2aAwi3izwi9H18Y/IPSnidePXJnd4/eWGbEVL0QvJuzqupusNXf/8IhVeDSFXT3szqy6tyvWTh
m0cU8BTC1UYhi0h08OwV7IlnTmaBr5MPXOeLAJTh3j/fCPJs84U1YLACeg2ZlAJu3HOVESh68fAF
zXlzj5yaWj4Gm+E5PqEGWcx/p63o/t9H479hUrytYZpmllcKgwoaGtfs+vBJLeU1QSHCA/4py60Z
kq4+B887fqU2yxoxtVLW5yKACg2P0Hxra63sbwjttbX/DbJ+xXVSXK0i05KKCDYur7pmqU5ZyPT2
3ANEotPg3wQs9jKwVPVdTNYzTUuxR5kGthKBbJAZxezQHutwW98PtPHcUqrvqa4spB5Ye4ZqNpEN
VoNLBqpM2wqyHfqHTnutpJQSGkUOoKSqqXVEOsSXxxp7cyETYR1m4dxv5V+FMaqp/Mk1oTchVKAB
N0Y0b7RVyHC0ny/c5Mp9c0dML4NweuFhBVXM7zSZ5/56N6XiutLJpgMhxCxOfP5wLUY34t5/RPW1
z0U0id3WtyuaXNMpE76RAKHCWRteDiOvSa+YiXRCEMyAw2Uorz8zV08F+1EViHALovClEus+BXld
w6ASBHVp1ow3GBroAUKTtjZBTs5jCZ2O4dxLCg95dsR7RVekuvwdAZhT9FO6QoJWSrL4unY24xqY
k82fSdzoFK3KxNu3BEgHub81ZUY25Avs6Qs+Yc4hJMMMpAA/ysaWCRuf7dVjnA2onT9QNjy44K9U
CVm2PBePvJDfadvyLRMs/2S7bycJJ9Ux6F6u7G4kaN75++UDdmcFzVXUa29linqEXVgNl4eMEehG
UlBzYmeDyhi2x7HAcx3DZlO7yqwAJ3RfIZ8YoUAGf9B/C0qDbrPTsUNE7eFozH9GlXQ/XyQWFdW6
2z50/002qg3DTyTspvBAwpmCQ5FEryeHUzz61JqD9TDFNQQ0CGEQC4PTFQThb1HfhCaWyHiIjRht
mMopgbABiqfD76lxoPGT+nY2fwqldhMk6mHWO0VI9AbdCagOb8peTOnm+CrTQPu7q/4iKoAuxMHL
HU2/lE0yHbOUz7H/cVFlD7wCDKU/WCeGxqLOxjBc8dB1czvQ/WrCHxNsHC+gUibiGQAqMT/eXc9c
HxS7qX5gQ34e8/QTOu/J1oirzW1isMuyds1/kL4fk/+GJc/Rka7fqA+/8+Utpx2iMB2Py66vMCkl
OS8DCNKOLfAeW3uMoPYKTdTlhlixv1uhFBHvZbpeOuP2higlRpo4RWqELxSwEtH3oeMDo3u+cT9B
oEYesFIqk24msnnyP3PFpXpsLPStU/P5NuEvtwey5ZZK+jzeVTk4LOlRPweP95NttngNmpupAh62
qt6emqhbHYSM1H+XcJNdSBGnrqLhmp/WcdaHSYPqWmh770krnEZomyJrDkWjlsg3NxtGce9prv2T
XH8zYZu9BXA/2J0IgQ/Sg4ECgKNWM/2CvUEpbWOJ33fnJKaAqSMV0FlSq+aAM0ThJexV4DoxWyjo
MN8QJSguFUbbEb/+EEbQUmmJk2hbOW5KBDL0oex60sfZB3QhB0c2F2FjGtnpRCIvsY4gVPAqUHDf
qwS3qmRIT0PaeN5l80x0dndMtYchgogWB3uep+Ob4c5Y0jGl3zqlUv8YJ3ZedB4DKEUxUr7OB7sX
GHs8iAiVngQXTLgjDxW1u3LGG84awLHNYuNIEj9K/wcgYII78wDJ5anEmLW6WtWNlW29aRKk4C8r
4LXYg+p9YPIWivk0Yiio+4SAQy+N8nrsfx4rvy2Sh7JBS7mj/03JrhCPnyxl8tigQdAOEgYgPHAn
FaJDnng6B4O95+XsunrS+yxoBb7jE2ewJSwZ9fZ5sXFD3M3YAmIRhSWgJ9Myi+orxvhgJQjpo7Qu
bR6xCAATwofUpa4vFajhU0RwRLRhnyxfqpmvNCVZuLqd0qjDLAwl2HQ2uqxvSDTpA/aSGvJCJwXL
zrvgk0x3knJrGg00PMd7E9w2KdbffZryDEdcgnynpuWVHKPvXgCRZZ0D8koY171mVZ7T0X4AyzgI
AKUxZhNdRJZp8TqqvAcf9cvCgF51awrc3m2/kXRK2TC3bFHvKBUhIXBlDpttDWe9N+UkytRwGx5H
qjrF7j4uwuzoiyj3arKOn8r5P5MemHs108itFu3C86qNFB5pAu3BCfFx7muM6XEMC8XabD9+p3Ll
zXR8xMCN/YQ7EWvsNuUxgnXoYEpaCBMEAUfBcUu4AcBxFSvORwsiaThr6Naw9BUhrCJLE8pgI04q
eminxOu2q3hpBWUGwNefgcUBgQm9V0hZF3iYdTsiUIsj66cgkXJ21vr7FbWKY1P/B2F/8uH3j4Le
lX7OlHrpxAZb2avznvsc9eTODmH3M6OWvl+qwjo8JprQjvKlBFIoapdqb3XXfoekCw6k3k3JupCA
QGd03CybGoehqNhxzOoRbx+u37ZnXSPZeMJg5iIgA5l3a5KyEhjgDeHza+CJRwnOes/gwD48nYUn
xZMtSleCY3xBHVs9BhfZqWsRRgve8JvTHX3MFPsIMZyuo3UtKDVSVuvzVBuC+5JcXq3syjfa/jgk
H8tl/r2m3riVLjmON747OZhMRB8l05sw3Ju3ti5VlWeFZ8rS1m3DARqz05t5HjtmD5qxWc4THFI0
RQW64s0sdN1yYM071B28uPHpLdTZfcckXtvl1YW+UfxXfWjllWarIcUFAx7h4rvwqf1rnfHh2Im2
e/YYWjHNyJjfvHj1cmsyCREYwoVS2qNsZKy2dDsRFENL5XYTV/XFAmfdFOqrleor0J4EWO63BEM9
odUQfQkLsmZwppI7lGus5dZyDvy61KhQ4upBn0ayseRPfk1LWaf9wxUDySWqnpR+G57NinR5QvnO
gRVqBn13DvkgiDm2/wNAMavzm8Gms+EFIdaCx30agrXRrTiz+PG0NvZoDlFjjBMRHDYL6H+9kJUy
mECO+qKm2JN1geaFaHI9VJ6MVfzRD2tMyLnW3AZRsTnICJR0W/r8WXDRrnJTTwRjKladehnUkLaC
5pTA8h/e3b0EdDsguD/gERXES0c0b3VlmdW8n1Q+MlNmQyC8yr6jBuvI5p99aB494ZUZWcWNSMb3
2oMoSQoUQ6hUTtBsDK0Rbmf/5oDFZ+uiIkWlceQE1Fp2N/HvSpD1cuSkKzoIsdYX5T6aGksYNhTw
+t7/9sA5r1nyMCaotvChBYuxtCh8fx3Kej64J3kZd7ffDryun8SrG6dxnyWe7fWG2Y5uKe8Xbo/m
ad4zx6M5tnr1yfLxsQldBi3kF6UZ+Mlnoqbom+iiHmcMNx//IJ7rmvWYx50yYY0XndGfV/MrLgF9
16yDVOkaIvSYJsfW6ZROuvsSUSIlBebuj+Jok8Jh86CHVrEFhmZZY1ouyRuViOvA+xuXQCBHmwWu
Gvo5kjyXNsLrAmEeZGM22RmpCCb1vNfo+4c2dSJbHk+2Enh3ZVvWE8a4K1VbTpoQ6Vm1/BzlVLv7
eQxBsl1/wFyGoGTYAe/G89AVFMOs2cO+gtbn1uLXIGZtqKYavu0zlDRM/GoxI0o74TbXlXty9Lv6
RG7kJyjdlU3nAWaPk1sqlPwvN/bNFpw+4ZfLYSRdMeclPvl8oyUyrLD3Wd+wWt4ZVJvVF63HuBuM
gsAmBEEV7wNReerCsLf7bGxt1cXfCA7Wul1aUsa0ntRAQXoVUQ+GsdnvANMu+Kq+MCyaO5mZ/fYK
UZzUdOe0JlUzsROJT1rA2CKIJ/vIILESHSYDj6ZdsWmNLclzLkpd9PmQ4oCPq1GwTPK8EyYEC/W/
CJDA2XcU1x0lVdC8KMzB7IZ5/CT5RFLmDhHjhqWR632/mjj08mBbUH9Diu2LVJ5nBjGLOBJKhLhW
BQQ42Hhilxmn6RR6S31bMxup2eLBx3l+WfrXmSH6475YS3ClK1eIvew9fNE6mhBoMLFUbA7TaGsI
HhJoMcM2lk+FtXx7Kq4DWMDQH/6oMcZU/3o3qN/u5KWChH8pj44Pr0DBy3aUUPHY2ayWmGV+jnA0
cLxCv7hE3RoTjIWizdZOwPoeumCALO7BoggwdsN1DkD+NXZRL7KrQ8eKdzexbTsJ7Ef9LDe1FFn0
abkSM+u2DtIqlTMTO356OmUb6h+E2oKjPfC29e+sQk7Fgi+JhDEXml9JHmpX8I/TDaxJKBjBoEzE
fmcCuMOCST9aKYpxsqFr2P1ncyAxRQGBFGND10VFzztKCT0OOHqd/3sqF9yEcAIFMkFhf5drtjW9
nF836Lr/L0NMQdEABij2AUbgN1swMXita7+xEasvDYCx5mZsnNv44LFrPCYP6PlTnxpfpJI0Bw0f
NNl65uxjbbyxanzALWNMnFFIwmAaAU+9kb48zw9ui8YBmhHCDYALvwac1upBaxEtSuTYS5+F747/
f0FjXfBpoVaJHBHVGzmEQH05fiqSm7IKvOS6eiJs3+UlBRphbQsuCtMmFzRiFiKfqvnBP6F9/Rv7
Ezw64tL1wNk4UXv9uH7tRah0hYWQd41oQyZjc5/kCpFwP/bcSj9Dx2oz+Sw4wBjibesTw7+SJKC7
ZGJZtURmqQW6jqNxtbWv9HSoh8Dvkc/JkKKEDE7w2bsUlzXaN6uZE0D4N+K6e20XbV3Vvi72m0OT
Dd6PZHFRT/Rso27NOfWu5F6hixFe7JDj91vTsg2iwH6WCfMlinrslFqNcmNs59FdiWURfzDHGCK8
pXMlNrmeXePZRWcmaWdtPmLeVGhgEmWtqSxYxvYpMUqVKpjxbvofi5cWeRadsg1zQ8tiA60S/wa1
FMbyk+DIRFex2AjLqTiLRjof2TS0RVM3oUFdLhteDoN0zpJqGOA7S1gY0+gH7tRb2fF/xB5RYNEW
zW769NrpKs/C9ztH2AtTU6ARs3BuNKZ+OTHtEFOmcvlnFYt6dvZL16cNe1h7NpLNF2lMcrpxdjMy
+yRreVd8s+4hQtGXC3FTgYNrU5sYbNR54M/eJY1+t1/FpI9u/0hhnorOYBNcYEJToFQx+nqVTLsn
/ycGebqEc/W1RbzzbQ9Pnkd5WXPzT7SDFM8EKDtMX7rytk2EBo4c/C+r5NaGc7XXofib9ahhEnMS
YgNtURHKoKSFA7cKKqFwuIMbsr64atU+PinIQXvCpvLvyz8+7xLVWi/GsSWK87ogmw2v/GY56u9T
18d9LG0nji4SyxAgUa7oLFpfr30qpmnjuZhKlA0cMWOfnUJt5Jiz1T+9DpELPOv9gPl1SO6ICQ7j
Tnr3CRYwsTwrnDQk4OZgYxODM7cVnlEXoK/M+tlGTV2Z7HLHax+yAZcsY6tonaF5WNdFLVRcpu5F
lHBalwxkB48XOsxtHkQUqKaUU6kO9IbP1tdhA1qtByNQtYDaR1NXpM2K8FRo1mz0+l0gnDtShrRR
0CzIca/Vd3i9/aS6zfWYS3XH5fnFh6uxr+6h4PaIgeYeIpCsup6kBE9pX4p8TjM2S0TnglI5RI2x
V+i9EPMKurmskQh0g7d8Zhgvv4gKWizLBlmXRiGz54YXSKqE9QgEnvXblIIabwIlFZMbfRTqm9t9
OTFDL3cH2KkJ+EBaBDPWeHGtEDWL5nYmC4d/oXVfUkglQKFHch7+aLQwcilGLyaxGrEa0eGLwlwR
mRNV97BfV5diwkqrQxaYdcZtgfLtsYKOkpAxuSsp2r4rZxRp3Zx2VTz4ppCEbVFu37RmZKsnpHCQ
y+1BftKnGl5wSA34LeZV3CEskQZ7A1/tI/3xqXWQWeUrEIJ0UsZ86S3wxw5YSka8UqCfvK/z6hWg
OlaXdlIX+HXY8rZD3LtI/9fAinvoEK3GF4Q+6VuxH000qXHGVRmj1ZBWzE+dUFp/SRxOuxWMuJhT
zAGHRIAO7/e/TpkUFteYMCjQK0/AM9UTBDbGTektAsXSMmx4qwaM2c/9KxfnnWPibniR8jy6SNA/
kJ/N+CHgz8nNDQv4pZrY1aWeU1vSW8cwTbzZ4k5ql96oDdxNWSnTuIslvfC1a1+GvfQey+lEm2JU
xrWBjSIs3eJM/gy7mMC3341p5fsFNSJ2RsewMv8V/oiqJ/4uY02oMw/rw9/m7JmEhNs+p36fvFjc
gxpj6V/QglWD6wFbjXFaPOsUwIBm3KQ1l1MYlLzau08bzdNJ5NjWs0qHICUus29HJs10cipZPASl
/iqEokTroZ/gHi1knY1bpPtX/Ng3u+YwN1rBklatC165iPZgx7mru9OET96anIlhxgAkFL/V1x0D
I0Ajac9v+FiqZc34NgURr+HQXhVzaytyZJ3KxdYyznbVoqShS19c2lLXPwg4G5i1SDtMrEMPyOwc
WKxBuJOaV23oHvz8BQybc+TECwhP89bUqKjbYLWt/j6LnX5jSNxjNBdus01aBYL0KqdN4tjHPQsN
m35UpNTkdIXTBdpORhk1SRu2/hc00ea/2/E9xdiahiIEy5FY13nvNkdQiWNqNokrff8uMj8porEe
z9lT15qcoRWR1qXX2KnXxaGUWUQ4egmo+f47CRc/I932B58xNpIyfDqlXY4RNmfWO8VUcZZb7ec5
cbmkoSH1BzE3LW4hwBc3daXbKp5i3jO+UKZ0raAXPwDRy83OrVjQlglR8qR1uAd60vs3H3JHqepb
FG5QME1H9/zm50xtyPFHanOA5WeNeHL2c1ZI4X4DzIB3DY0IxrDYE7MHoNKGOufMrycR0HlM5sTA
H/WoLaineLQ/zq7wW4qdXPYZmdUh6mWpS7BAk1c0z6Sp8xB9POxUeAzNlr0K6Sp/VKrFB0rreYzQ
8NFXNqBM/emY2SedDjoxXMtqMXgGzFyzT6SWXNrrRUTKHjF9LDa166GzfgV1rusGTzlgKFMTmqen
hRi8I5ElWLR2Hx+xRZ/RvOja599z3BL3syc7AA3kvfgm7I2aPA8pdUL62UPuvttQ8GtJzMA5cN3u
JSc0F+j7xbMy9g0QO1ArOKF7gjCesmEIInqYCBlNqeIo7WWmExwuNQehwaqJ7ez0xbsFoCCw/X0o
bOx7yVVOHxiRvDfZZxfVZQ5ZEy/IdSJKdKje1LqxjTTxGadh1fOX+4w1e5Hc8YAKvgu8ojKtLB0H
m5pPnjA5T5BnLWr6hlTpdJg8semAIxjKB8AWRomigSdazLz0mHmxK0hqTRTq4V3FE2glU8ByAVxI
C45HPMrpoZ3N0a9xpCfu4Cxw7FKsggT2MFBUt5wRxMjmDyETWjbU/bS6137fqAMNDHpPaNTUKDbf
0hnTQgjgFUxhWNOvX0UIw/Upx771HOSvi9t2DVk7dIR8CXXFEJDQfR0Q4Cgi4kl3kogWhAdOjyix
8WD07x/OU34iPjcQwP/K19hnLVuVdM6oh7QbhSpJsHv3mADA+ORIiFzvnyqqRGyrrkrm2No6+aZz
al+IVh5X1DKNyVbbwRZhWSReK08+K61wXiP0SvVDnsFR59ZOYDpCWAYSYTnCAqm9lCGWIKQiXYGK
4dwZHPaj0Mlm0bMEGmZCF5thZdsZezD4TnKFcRbQibmGAFIun/IOv7zSZ52w4Sg4Ugyl/qw2NVeK
TffRqtgWdTPf7XYXhszKyS7EBtxPX4QkgxgGivkKw9pkTEa8FR4loNm23S2sepaoL+tKioiR4Jvu
e8GkOpY8qySU/mKQXRKYsfsr6xe7WoHxmzcKw1Qs6EwWqbTi+9d4NnG9U6K0AB/eronxInv8wN7t
GmAMKyTtRzYykDudmtMFOxZUIYD/7zbifObBjmSTB7UrMS4VdMh4mPXxnN3QrwFavIRicur00oJN
xaFTgB0GSbrkTh0iF62kRa5tme1zrqVHDrWYH3ouHFj7ghcxGyZPEgMByN3CY0lqrfnN87YoeEQB
wDOWF92ijbPwopdJjiAeBJ2lsPoycX+6ifu1SMdRTwa3frhSkX5/BZZnzh5ZO2I2uUAGjiq+lxLC
Euk8HjLxkBQ5ROM15L/xdhSmlkT+9NGEkNcjUivaf10pHMuvtFfYK0oJgr+hsHtGdrpQOHJr1gvI
c9LEN7FwsOZoXdrxIaoK+7zlEKQ6kwfS820WviWFJncNJkeM2DbNwg6poWYQghI4hLm3NDo5OzFM
vCx64EYwC47EV7+D/0HkdVo9V/zSZYVkIGELiYQddsCUEShYkQ6sznRKxMtzZNwcc31eg4BB1Lfi
pFh6yc97EAKApGeShdpce3wD3NGtNBuIAMMMKKpv7295VtRzw6c0VkaT2WZnrf+r6+1RPlgfvvk0
2npEHFLezKuY9CQdEM7oyK/b/E38hDbKX0QfI+WrGTXVYTINo30zfkcvV9MO5yHfxO9CYyLlAU1w
Ir7ZAhAJCal2rs/+zmY/pwOGH/Y+E7+hXLA13FssbtXnq3cukw7sRRlnj8E5jM11lvbgM0xa9J68
VwBwpf2Tr+HSZ2/+9TL6hsFzO3xWn8T6BVtRUP1NqzxJpJjyrb2LDmO8pt5y8pcrFuhqFqPrecRe
WRdPrfBfevAX0HUSjhcTQnLLFhc4CEZL4Yni5wv4d0AzP1qWYkviU1HAVIvA69pUsjiT78/3uWX+
rBEUhTvP2GtN66aD8jq6XGZxzYq7ZU9zuu9jkEcCG3MQ302GfynW5MFJnuOyo+4e3FnReBxmzWHz
sbkWIjBSwlsVYpgxWpQ/Nt3FQZQFPjADayd4omqSTvhN6j1Thp3kNyuEMh0AIl1iOS4qMwbwilnv
/mdE7lAKfM6Vzg3zwGgrgPwu3QVFEV9dyFtLIiHMRGkHRjmSpzzT3aoby7WH+UasMsefUG6B+/sK
CkJhyz7uvExHRPCaOiE/MPWmfoVpz7oH+PfRvq02hOq7pyKoFYgHkPePwaGCTmTR8UmeUFEN3Vei
q4InSVnbPyXx2Gh4L2aO9t1PMBkdUWKS0hV0s8i+7WDAZ1twrk1+DU0tjIUHHHSy5Y1DGtm+mdS6
8UDbtMy6vEFUPtSt6s6GDr8tF6YK06hk0mNXaI42aT+pFP5mpDkiuVaBHGKxuOMaQs59Je5QM6hG
mGAtQr5YmOHuoKrQBFrFP1f2nRQ89szUXeQNv/38Kxo4+ozOHLucvPMfCd0ORhg6AJOU0v/g73vR
zwaw9DM5SfhjLHxML0bF7lW4u+RZtRYSxE07fTROitEndTNDe2ZCAqG27xKScue89mJ+x4WX/Guk
hRz73LeaBNU1dqazr6bjHf7yuZBil/FJ1eulUr+3f6IDaWrjQlRyzR3JS4u8wzLuqi43sA0VIPt5
9Xj/kSVGyh8WwmHvU4QZ9vyIUsyBSwdh8m/B0CxN0Vf1mbazQ9Qt+tGovR93TjATwCcuAQHBu2wj
T7nPgPA3ZGohNCNFuYxWQWsxp+oteDQBiq0D3tbgWJtNIqk3uTNUysxTar5tatdoYZjPiaFLNNjt
k4T/vpqlYbhfKIHWtOe3qwVT6AfLiEQRA2ipmqlriz3Qe/KRUwOvTt2eyBhsfc5YUhIK6+rZq7kL
vcDtfJ4UbCwj2nXol7xGEpsOdm7Io8UaMjFkT8D92f77eWZhfjlQQioexQn+zv7XDtcNArFhGrvc
5lqYk/rkutbyj+Yn3jtD/XSHzIqUkH5S2QhbqUTWzJsB+fB2fw20cOJ4cpOzfl9sqidaIf3yFJdl
IIdQ8U5zvi260m5mIe/ziTxSKqJCpKlueMSBZ0oPD+adX+yTaJSkpf9r6mmsNilx4p43OkvjkIi1
INRUA/Z+3Azt6Iv1ab9L+EBAqa4SCBD8VVHwTVxqs1fdtotFEoPbY7ELzzhIS6SRa1Oflf3Yd2+s
t0Od2ChLjef4ArdtjIPbUD3TV1JhMY5gW50lq50aVXUOglGQUdNXky4xmVbBLcLcv0qG9Qv4MsJa
P2ZDr1S9/toDT5LHZjKaTAC8P33qxJlSS3apgnyvR3mNcDZpWqdVhT+QZZSSYdVCVnK1cHWVVpX2
3FwJy9ztUnmcJqmxkZFk+CxDRY0/80/JL6coVYYfIIaJD8kZg3yGjpp5HKOSedxPxq3nXse8893m
3v9q9WCgxsJz1jBHNnB4mLuDoOV1nQSv4mMtZ+Gyy+z7/BZgzuP85y8E/CvPtBQbNsTuNeGEJh/D
W1uNhG9WxIRBHgAqVG8n51IRzxFfNg+itmOcysNH9Px+9UQY+tIu5huIkftjOgjXe22Joy69uRSK
utezc6HOWWkrQdf3tfRmoS0kjR2CZDoyY7/tWYTrVB6cuzJzWb6rT7dz6eLutGQKEsym3pcpazcw
5jsCaLo5dnDV0FMDbiYZsNbYAi2bDbHKog8vCRqI7HIMdiCI3Nf/8fb1RTMICwy7UsgPIiUEqzQ/
kFFck3/o02oQC2DJZe7dKkssTN0tWvj1Hqn9pTtma8PSMU/i7oAh4zzUzRgV5GwdT+5mPePgl3qN
c/OBzHEjrDaqJza37qBc84QJnXZ/FTjgrd0JOZYeu11sqi0yOsjSV821n2sqgFOr/8vFcyPmMJf4
2ghiaGGoIBe2U8tCI1YV9DezXTZEDo6t8fzcTeylAZx0qpHULKWXPW+EM6jEaz/ZUewY+Q6g45Lz
bBUJZ73aGiVXebcwJ8p/bP/BNXn1f/uT+GAqiLIpELfqq9dytkRLOP+hwqyOh+qWz3tgrHjRmfNa
Xmrr5LVBoXArZd2z7aPWBvgavhmKgbRhG8m6cYd1yAmMEYXXf523xoYiHCFtZcn01O/asG100u06
YmRbiYasqBIkgzAK+B22EsHkGYx/lxeeqQfzE8ImvQnaTrxh5pjP1L7/888ZhEBknhSyJNF93/M6
bz5lDqNphQPuc2+2XMDz0cPwLK8w3HHgbDt2X1S/bn4ZzDGib7DcAR2nQa3D/2HzZ6PgHYtH++rR
Z47qY6MHqS5V6abgOJLZ2aBz5RgR8/aw7OaTn5KrP8H0FFOrr8Aj+x2x96hvPZ1SzMzdrxOeBHNs
EQFSrrQX9K2P+rAB8qMCzhsl9/lFx2d+7VTb04KcUhLShmvWnd3G9AeVJlb/cn4gHHIQt1GYELBP
ma9hZG/kdBfglkYuVJ4x8f2edksMYohC8vru6FbddAYFB0NHCpNY5KNVLgVT0EBAhNOT+yX4cQeQ
1ciExl4tpsfp3p48L3oHbBWZY1gWXmF3mz6y8WkFQTf/0fy+Yjds9kd7Xt+sI0R0zdKQUtb001bS
64FIWwBCuoKqJ3Z9I5QWp2vVhpha8aynXeGRGP3q47kfuR3CMhHER/OwOxPIgpJMck45kcicghMB
PGPBbE5B0KpuOCF0LaS6DTpKFr/hinQdP6AEE8kVcWcfAEDCgG0Q7VsMbBfiVQDy2i3xlBxot/C4
Ssi/DCXMKoMdbaysOxx/hOsVqRCwzv1sTQ0mOKMrpvFSM/PUy/UhvYqSs2yqGs6CCTzxy+sc096P
qFjzN0TM2FSs+maMSkKKmpXOe4v4ATmYeM9ep/1zn5OpW2GPAa6HbgFqcOHrgYSA+befmAZZG1HM
Os6t6F7fgQv/+omWuIReNVic6H/teQcbhFydkkhyGGgVhwGOPcMwDKCdsArbGh9Sv83vluiIEGoW
7g8DfN7Y/ZnNpIYxj6s56xbJUnsYkHupW+Vca3msQD2RfmQ5CW6SXWO6g/qmfO2RRhtAAApyyQa0
sayZYwFzuE6N/0ywOhxM0bzqoKnLRmBn6DadbrlqpiYQOSAc56TE8iyLAGp1AxsNu23U6HaoX9q9
XOqtacQntrSSw2Ok5+1CEGJuEpVkGBT+DeC2Xh864I9FKra4vMAcQPjP9XLshXXDZRi2Vsh4o3vr
j/PxXTjN/KxMzxxONjbIN7AQ00xmMgG9remDDiMA7+ReesMgj8kEh6hKqRcnsC7OufFm51goagWz
hAvVrkL0VfbMWm6v8OqjK4njduN5+9d6vGq+icpiTWvmgjV/p8LXK11ZWM48n7kYY3179cUH3NYC
bqreRRgiNJroVFLbjaT/znp2kvnz2+4hNr3SwIa7RHXtwnrejn5yyrFim0CzQJyC9N0uOIf7ESII
3uHdsQOIvj+Tf45nE+QL79fORnaXn64Ld1JA73UnhgInNMpexV5jN4Yhc0p8nYgT55YaCfFw+vOs
cUegVtukcyr4vC7AobUJzfxl5FsWXhq2ae/DTCTnKJ38v4xAc8S9zJ8U8hnSi72WZMVaYgy9xsgB
6k04VtQeAGwDFMbYim596S7FYwb3wqXby1M5d95xOTtC5NbCUL3coAZRWCBg4Lj9fDYekmoWrWd0
hen7dDpmYw+gW6TEvBF7uqC7pCYcQhL304EkCR17nNUt6L4y3k75oni+aBkxDEXsRLRNNhzNP/cm
B62jZCsUsQQE9rKFlz9gWgMquvTER5wxtZATFE0lK6mxHoz+ZefsSSNScVd24bIygGtWSnqQ92jO
Q5SyT5ptAPi+25umd99hpDCxkQJMz0tEKcClaA64IvZ9oUmW0ysjWC0zX9mY66F/n1F5Wo6U5Bcm
svmmPFlhOhEx2W+Z7QFE6TqG7mshQ8nTTCrRkWJbbaTDMtT21NYctVw/GpUjZ0ihPP0ELBqTK4Nq
ntAYMRdRA74TAKyfOMYgX+E55mOWiQl2IT+8tYAMasR6qIPUt3tsULsEArixsJaD6u4xgBtTsc1d
jF0yVhBYxcLqjn5RibB18yEMHWKX0mlsDCo1Q1AXWc/FF8qFU2wlLPZUWsvR8iUNojbgJqzX7Br0
Wo7xWm2lt72AqjxarTBXP1eeF84kTr0RQDO/CwT0cdvJpJFOzfbcTJiL9Db8EZGEPW1jMcxhSbbH
vZ+u8ZbCdlyVDjQHjXf3koKKTwKoiIZIcGQGvnFlpUWKnNGo5VS/Vrbx66KsfxRFh/B2D+16Cn40
EvlfBdtxOJsuFMChaLzjasLj9o7mOWO5GnLxk1VIGBVoyWrN+LURQgNNzt3+Y5IxhX3Mo8t7bXU2
jsArpuiY5ZnkvHb8Pusi2OUQtgoGxtARoPWhaBc2XYKNF3KVg2w4mUAijzqj7w7Ar5gHScwLY8Jh
1CbDTvR1yNUWQZ7PEQA850oZmD+luzMEDLDl+AeGU0ih8Q+cqJu55e0Aslz1qYy+FN3mlyieY9p+
VtAulcTCk0owmpfjnC6M0lbmOQeJe8E/7JyJexqZ0+O8IvMMSLb9/HxfkwC89AbCMHAR1jt+xuxs
5pLBJTzKeCZtQRVP92uPZL2fJdNhPbQJAKLEM2sLNR9XawSmqfyq4LwOTcX1qY7UL8oFeRPP2ET+
4tw178BF0bc6FxA6evickSIA8SEiOhiBr5xAL7eWBD1EMNmPRy+4q0M38BnQMAt1GEiiZNgoGQ2t
8jVg5abUDWyGlO0DT8Zs+tX/OEM2hFsN1TqUAmi6sg+zNfJh8o2TsYcOrJ9okwZfeXeeiQOM3ezk
UvUR52n9N7y2CFREi9BMwlOc2hF5Pxh7LgBhrX8rmvuTbjuHL3Ezb5Avwf8No9mN9SEb625CW9/M
YC/ZoHD2Wh8MKJKC2BkB58q5YYICL1DXMees8WKPIEtSevkqiBxp+PgHmkPrWwK4ifi4ZrJSR694
xB3jTL0NRChLqKXfdvQQpcOQqYaWSin9bFwzC4QeW+Lk2wjYTA1CLMgsKSVn1XpLqkaSEKId3S6N
Db1wn9Ragg1tcTRVHQ+AYdFB+FG5UPI+J23mfzrPB3cekYR7ql2pyNVuvDZX2F3WBHmP/89dc8zA
JQ4CvOnRqno6yKaMQ5hgKRtIvBqauDCoLegeS3b+mUTHPrbXcqxiC7DNPJ9euz2Ric69dIe1e3XT
IVOtkvStG87CCVu9UIkXaqHUFlgyNvB3B2mYPaA2gsobnLfmsCMG1yNGYcnejrX76ukfFQjFqkws
CG4teiDHrznaL3eA60Z4PPSIPYG9HT0VKkNoo10GquHMcHUZ18pPr0BhDJlkoEb9pq2yiy/FZCAi
uA91VTDp5As0eNhuDB9kLHkABqJCzFMWCgBrk++OgLSkRWfrD7gPfpwfyyejwuZ5dvNYB+Xz1foX
DJxISrKGnUbDnN4Te372qkEx4Zg46RnU0lheweFYEkzOIGch7IPXvtoJPW4DmdmWYvGh/QLnzUpj
SWAFuni7SUcJ2iCwB8GAdEWu/e6rxL5n3Bsll9F0zall8jOaBoVRETyJIoDjJakhX3B9knmZGe2w
6XiVV19svj1J05owtyoBRTc72FF2IpnkkvPnyrQ2XM8XBc7M9AotPsIo5BQ8+bul9bMDKcK49YjY
Mh2K+iPLzSPvZewhif2FDM6plOY5VS+IsBE3cDEktKbEG1QUTQlB6RsrtCAtE77wOYjQWc4z20mT
YZrpHYBXke5uVz+ObKVJLFr1z1OchVl+aPpiK5RcR5wJVXKU3XfBK27ky5B0XluC2ypbneN28XL4
0KHQWf4PJK/nGBDJvgbSrkBx72Q21FcaDhfHVQUyrfU50PoRL5MpmmQNKaOipekEKg1rIIqUPK8H
Bg5DLjy7O5SqbMfd0wbWAggmEfVyKKt7W+wxnggtp07NwvaC+g+9qAnoTRwwCzJCx+18Z7zPdPk0
q5We8PJaAQnHeUNbusLFKDp3D+2WGQXXNKry5WEog2RodwyLXrbZ5WOGUPRC7utOonCyYkkiwnpi
T1itdh8DaS8ZVy3j0Me3MGxh1OM7QLpof40WvObjRwwZezhrfTmXgPIeduT37zAYRNe1/yIpI1Vh
iji4FDOgIBJOpqJi8A6rUt+nmAQadmReMXISEROpK4wVdTLOGJ8FkcjyFUoXGrQORJdyiLiO05o2
dG+aMOtqE0hqtvS65mAKf0Rcuf0a6zUcm5PXDEIFOU3leY9cP2LQf50l1mzPLgObbmd0eEVXup0V
lVcBihIAC9U9ngVfr4JYM2jHte2x/vFqTtLi5JfFS0nglY49tHTU45iA2LvrmjC8/Lpdw2E8/zeP
cyT/u/f5pBmYM1dbooy01bV3sbHjoOljNn2Dmx8iJDbY4aFYUwuPZMNyOxRTyywRTHAs8Viy4r7C
CkIM1RKKoLT3Ug1H6fMZ6VnH8+WWQZrB17JXLtgj3KCB+31tzf+Mn0VFeobUYgKDGg7jQXQqlIea
9sfWeo7O9gQFHQGtU3ePomD8Amrd1B9ye7hDLSkbCUA1SQfEJzDjCqh9q5DQE1hTuWFoIAeuiGay
OnUc3fs7EnkrHkGrF/usq4HvGrkyndHzMfndynykicsNkS78CsrsYa68FvNIll248s3XgVDjCrlN
CLGA5vqkS68Ynpy/BCo2nXc/4qQyMIc3iLFDK8EDjzHdjvFovgoUeh5rNdNrShqnCM4zl0K31DSr
AxYVUzC6wftwzLtyHr5elL65zk5GZlAAmsIY6VENXnQxF3y6HDTo2PibX7GhaXmPirJwIvommISl
pciLmCUYQi9MjO/gwWxWJFawo6/v4s6M/QT8MCOhPKJ5MdBwxg8D9jMXSi8zxJaD1PCqju5bAY2Q
EKZ8b/KTKoJrUcGkiCnF99oQp5IdUCs3/wlhBQsvXgOCXRKPsrEArSWXQQseEdWWT8aeuaWBWVVt
3D7DAIyAQL5eLCz5Rf1vhs95pTdltbDXpSSsAqDgIqdYGTdhgmfQ3rEc/5n1ASj6s2Eqh84PksJt
BLqtZA5ADVEiM+e8QaobRd9HbwWFLkLah4TIxzXuEkgQT6NREWWt7b89G1Nk3OxDIGe/TxmUb5EJ
hnrO39QztIGW+FGC1scrjPgWaheM12jjmtpiY4QZsFICn8x+a7HMN3OVNIF/lUGRO3pg5tmhkHog
McPf3kjJYowXBO1AeNnEP8YA0vVefz0Ud162RUCnzD+heOVpHTEX3ByV3dUPfTMep9hy0YOMiT4/
fV2QlU8fLKTZEtrQUrIaZN3Ut6ZSjsa2zAAbw14lQLdM7J10aHdEFEUp20Zv0Xs2R5aOAIFXaKT3
5bGePqEJ7xkJIZP9y0QGY3Fhb5/FRizZDUWLKBgWygtJh5KR4eov0wrKZYEjxdQG1DTG/1qntero
aMmL62swpq3uKzREEZh0X2fS3Ng7IeM37jAlgCHH8aeSwP1fDJzHUFkMNPhHGsqEGHNA9KWBkLkL
fUWY6Da2ZEsia0IyroUpaOBJEkxh51QhqqKNGTeadq7NnKdiyOoRhtl72ZpRtBCyBSPcmSqDYH9f
rTNQrQTeqFkBUj8rXyCra0vGJl2uTwAAvoDbWkVjwp1NHfLCdRq0FET/wilCRceVKF85MZkLKA6E
qN7yLneyJJ1oOnenZ7ORlB6oY1+uMrY9YvaAK7Htz5f7ngcwhFhp29MkeD1NeeAvbfv8hscEC54e
+AbxIQAxio8EFljDopuM/XECpCPBz3QpVmDnXxmY64ynI79iPPWx4bEvuLMnlKGen5ucl0wpMIYL
EvtxMM06QPrhh0MYTz3pON1MbIHxiQjyqsgdoivQO7tg25NUZIZX5nPX7EMSd0qvBZ0tiPvdYNPN
unKqxtvfjacc0HnDIlOV8O9YeBBZdlOMIikIX4oXwUL+t93YYuR4SFLXFbfeg3+23O+dREvZS/ww
ug9BxEdUgIPAi7fwAUB2eWsKvXroF+C4ejKLLbHiRjdByQpBPnGXN1LwpRV2i3P8BEDysUCdne6I
Nf/iD/KriaUQBr0nnDhcU/CeXhIxXcyHbO5nc4ePkqznbzhIuBkmb1UBS+mCOyONEtWa1aIu9reI
nQdF+fLnxD/4nyQyCDuckwTBlQinIqXBznkG249nOoRPUR686du6NrLhg+16lTR4f3iFziL4/Qao
ppnkb15Uc6x9KQhggZ1TJBFyczPkeF1x+IzSX5QjMRZtvTn/mIdRlrq6KDgtQu5YEWLZkYvum8zg
TyJYm/ZMfb8gMeZMUors+N67k2+GfrsogJmpOjwGBv04lec/PwAL+Hag6Lbnhji4hz9l0aEcSWu/
Yvia5VFCnxofBeskvE8NNw9fOtL/RoPT0muXdlCR0sLUHr2QXpyjvjYKfX8yo4EmRpUNc9qNdom/
h9K8Le87dsJgl8Tr43cRfVIuB0IiJVxgYMqHW9KGX5Vi836iBUOm2s1yujhzQUTaAX9OLBT1Tu8p
oAH8sgxSD/BgABoWvu2cj1LKmF2lzbnJkoRYWppabpwWIniY6mTb0fnMMPAf7GZl0ef/5vzlge1e
hMXBEOkArjC6arTaoywnvYDARY5vFtRbEFo6UyZCx9aCr7XiTHqVEQj0uMJbewOCQl1XCFjUSDVV
Z5IYzIm/8vyBKxz28ylE0AfkSifRzbDmMnCUnSRhucLMGmdS8tyONtHYMk1Jmw+9LZ2r6scy3Q01
Q94zKS8Df9emPn613bQqGVUVgP53yfLEuPGPJxdd0rHPBYyA/iPjmUNzqiVsOma9Fa76b1tu5ezl
FUprmTfAMgD31MJg9nX7InkVogOe+HEIqa5tHHrB1GRgk07SyJKtMdORpSNnE4nSrQisTNi7/zsq
1TG/rRz8GrZBIx1iW23LUqPMgH6/LvS07lXNRgiiQAZ5SD1n56ouoLO9ivRG1tkk4CGrkYOMfD+p
lR6CkoIUkvhsxnhEc0gAwLCPI9hPjCv0j3UU0OUQ+VI4YBplnSCtFuHzMkMqf/IcM0wRD7oIvo4O
7uAmqPaOK5aAUkwy/LbT0zt0wN5/1hBaVcQ5pdYuyz+KJuWydaMFUvOxq64Szspf1diH7SokBUUV
TBBx/9OTB/niX+IUFGAMViEXkfDhUKyN5DJSOFNU4p7XIpYVOf/3Oq7RysdK4tPudDaonEerHjrl
8SqNqOWI8cLBS76djU8x4SwP5od2dSVXVisk/afvBVpRtMOAzV3OsmF9zRjoiE7slNyGCsIUISPP
1N3drmk4Int58DkoufvecPrb3mfZ76sOLUaZZnLqbv3VyFzTTb+kf+GE+hwB5rg3LvTobeQcKwYl
TpnB0AvjJ7K0OMJ4e72aulrLMpZ5tG8uQ2ZJHz2Gr2VmsuIqka1WSCWS9tWLhc/A1UL69vvXn0tr
T0zAGD6/hUmL5Wn/E/HiXKuSKJYIxSGqQUbwjTbf76BcCk1AmEC51ah+HowN5JYfCuzEA4kc7JMK
BPLafEtydOp4+ZibDzVfOhx2kP65pRyCk55V4hdyzxPsX2XNNbnVCEaBHLC0b+xY3NBhHmskrYt1
d42J9atFipVAqNmQPCh+e6i4uowP+Jr5ctgiutQReM2toD/5SvT9NAcWuRIJ7W3cfp7C0shgrS56
4OchSruHmynkkOa+AQ6Tib3kcqidGGuoRTRFS6NSWh8fp2BMgP4BBznaEO1LWycKXHejAzYn0/bP
bNPb11tFle3/L1BiJZp9Jkg9b+WVyrGRD39Yx9aa92WQVuUa0FQ/xzC+3gAvs214pyn+VmDFw+Oq
6uVG+YAn+0CzML+t53Js1me1TRhrOZbGI4e4POW3ldRU4fNe3hw8RGktxv1VUyBj2M2FY2Wtpfpo
ELU5Wxqo0LTlcdxRj7pqiD4V0/0w8I9wwk2rnUPrjgI86iu2/SkG1ILx0C9QFFDM0yFh7bODVZg0
IHvXrOyeNVUqn563qt0G/swc5bhs+7VrZG3gBbd2fUcsuAuYAbYg9UKG1t38F0GIpckHtpnYTz5i
1DkbI+FzLi+qTilcJhSJMMcvfCH8kDdHqNQBIE+47626/yLKCu/O0yDkhZtvqMbzGaFu9KuwitzO
itdCqcn69Vj40MrSr/nxIXDBIVZPXO7slSWx63oX0wOUbfz29Gx/TLnTUz9l5d7iUuTI6Tzw4HxC
7Ty540nDrhtKZ32nnP3vYiozJAxQjEYUGwyFAu3oT3Eodwbivuqyt7VMx+PUdNBoF42SGYLiBqWO
5UxV4kNelcsJmT2Bu19VCMdFz1XTR+oOLwaw3noxq0YsTu1T0D/9G2auxNI/Uuj/yVxXPdCGClr1
Tm8hKtjf+vvduL4o/lNRLjPIetqFdsmqtJWpIjZM/eg4Dse3UsgtH18FJilpPN2hIFZT88GIudm5
tJhQ6om5E6SNSNKCAx0VRnqsysE3wSt7l6l92biqTIJTCyToDQgRIQVrEeEUpGafShuUj7/sjM4W
g/DPs1YzIfPHx59V09K643vZTflDhXhmc/iCG/AnyeAzqKmkwk+X11g2fbiInq89Lv0MLXR0DmWJ
HCR3r0EPfUrRfVLL2Pi1U4ZFbBmVaT+FhWU4UziPbslUlBRLdOY5Ejjt+YPMfIz4PhUYrAr99+Pv
Ssy1K1C3yyCC7Y3RRmGFs6AH+tC/z1LJ+jvW+71Kp1EkK9tbklKyXQrgop77EtXM+ttd+pYats2b
FPPYreeLEvhu8npGHMdb8n03fdWI8IVho9butt9Kwxpmn2WDNmehGoVmpdLTBxvfN/s/vU71VOud
xpTwh4eH4jayuY1zrDZ6tqxY8d1tfvFK8fZ1vHqaentJbvy/2EJiXQ4lfMKwtr81abxvnWPJyMcA
kxhC2rluMXoQV/XBG6WpOy4CbnY8ONl+MVYmQhN5EwErdwM9zIlTul4BSamw/nbXykpjxtOg8242
SE/gnevy0sAslbDl5rg8qfMeqXTYPu6ku3egCqg0zKOQ/aN9xhlLAYs2SNAmzHD5e8zz8zXqA1KM
PTpWvIkXYS8E9nHiNU9/w+s2Fklet9IDczjAHi0vRvoL5qlw+uIKVjKHurLFZutHGryk9CPkXNsf
7P25OGsZ7+jvjmI60a2LoGlH57sbh5cdJZErdHB9x62Ely5hS7nwLoedFu+q5aTha5ScmjCuvZFz
Qsg+3/QjasLqHB2/1ldjGeviHag2lvBCVGi1jkibK4BOCj1S4rGtR/HoTesPF/HU8QFXMRp87u/3
dIKUgZ6UiuZWL5WU6688tIRcANPNKOMLa37uL/SNQpj94s9k1Vz2tCIZMSn5NVw4UPZrIp7JZpbL
VSTWB/869lOzHRNDBgglZXe9QJUiQI8HkuJPGRtpRN+x+Gmt032wJGjvA7wQ0xxWwms1lILbDXp9
yYNFTPZIFnKJ15aPzkco63nnJs4bQubMXjBBH89PTfJRkLoAsqJyEERwijunFKlgn1dsgJ9NjCeb
wQMTWcOy035iireJthHDreGCCGqRXwmBZ+5LPIghG4gCtb/jBCpxv+6JB6IhVYa33NhR6rbHGY+Z
Ez2jdyOgPQ4RgtPLsHpiFrZodwBPx3VR3e4xomQ4c48p9xc4dG9iPf7s1do9rIT4sojkqSDGGYZ8
vp6oD8phuKNnPL7vGpod3peKD5TL9s4P1gn8YHWY3PkstWHdUjGVcUWo/pKGK6PuVpnPmt76UVoy
+Ibdrk66glTdIvN2lB1UHZEKSbF+0BGI/oUgLKWWuaXuNLhc/akl33TSkiMKm7DclMbT1W+t/IX1
1vS1a98fvaOcd7ttaUgOlmDcElqkm7zfvk5SSFb4c0+PwVlU3dUNaNuxTfbrZwt6qiUcW9NoQhYN
6cIhQv3VJZfDDcol3puEfsKGIepLP665HblNBQmHC4YRjCd8QBfoCHeweMEWvyrxP/yYr6CRtIGi
HMs+TrVWKxbAFWCxG7lWNauCbOrsp3qG5+XbffO77nuvzPcgI0FX6HioKey8QkZbl1CUnY5RnC+S
lWORG/5hvOkovNk3LR4Kw/4RZ4vrejxO14tb1yHulciWZGBRSAK/jCFvxqjQXyvQEmPiMJF3PZ+d
RKz6GrUddqRHh+7fdXDrJxPJoO7acmygLnhMLgSfv+EbhzceSO08eb8bPZgOXx5/1W4NXcceDF1b
rGS4U6CD302nDvXFjCPHTPWd+A77w5yhPcSrcRb5I0TkdzSRB7nE7qFQ438lYsO8fPRtaHY8vhYN
9MfhWtXPe2qFGYYSII5B2DMnQGjjLXOEk7wR7QotX5cHM88T3YqDmr1VnwoBtKsf+pSMcf3BY710
+b5NtY0dtWCMQFQBAuBFakmm5AjvT9Xw+9/VtD7TM+BZPNj5Y56MbaCTkuFJ8NOcfvZzn7CNtA7H
rb0ltcL+Iddc9ERjepd0LnLjFKxnxWu89PtM7E/y5DJBQCxRNzbwyc5Eva6ZC9b5JB+/900ff1Oj
xWjxpJQA4Z06HnGCdKKcar/3SgswEix19mclE8Z5OaWEvogpQefhwX1v7ktzKV3HmQjSWBpSX33p
5z9iS5k2te9HfKywxGeGZsh7G0ALGFvAo72Zzsu5XrXh3rlGCUP8LuSd+9VKPqK+HOGihZXjUQwo
bEWO4f2lPcozvpbZizpcgaGc1ZhczwgZ0sswaS6uAs26AUpJ/pe8Uj/zgxdWP5KTwb8mWr3e7dMQ
6N6jNYlcciGldB/gw+3RaPOpjK9KUIeSFB3WvXxFRGAW88uTnjJ8f1gHpAhgKTKly0zSoalBlqAi
34yAr7TPjmmjn1AHPzAxLo2KKvuT2K+BJmrJ5351yVF23pKyIGLcIt7kpBdLwQmnbIahcyqjt2oj
frlPaT15cnlxBpr2o7wxLAKrB2nCFTzecijJCkJ6c4fKtBJ7mKtfg8FZOovhWghKcp0EKVmMtV6C
iaxcKK3zX7iujqYH0GvTzraRqT64OgfXPO087CvCQDnBoVBbJKarP6RhZh/9q9ol6kUFnDLiGFvr
t5A7R4S5N2+ehnbm9hPkZqxW3ByBK0MWqmcS/prlPfuJuysYrYooeXDYBC3sD7rlwgjpUT6m/8Uo
igNG+HxHkvlYzGZzD7/Z0tZnYJqWUm13ktyb9RAnFfk7xoLdNA06cBS+SnjGmttJMecS/48uRrey
w2+76lQs7uNTLi5jLXKh2zs0c7qcR5WT0pBPjNjkKzL/CoBY9tH8iYqsxqQMkNpgrfZpI8OcMBiT
pJadWcnxC1qgirfNCKGCOhKv/FFO2c3yS4NvbysdVJRWNbEUzFXtcuXZ5ahVWkF7LGeKXp/BFYxZ
JiyYFAcFapu2YNmh1Fbih+/U5hmwjSqHnwKR05IMVJkd9BFsRT4b1CQ8oz9UnXvJ1wWvegSG10Bb
p4tIow2wH5PfDIyOlCpDsEgGzcf2CEcqjPv0zkNLxBiUnc27VahUW6VsBQXe5C1fdIMccVuk3Lrz
B5TNSmoepktYnBc+bkfLDsVGCyZEwIzVhdVZXKnKmqzH7Aguf0MUl/X2mG4CxHXOu4lxTzmpqZ4I
BLKmtBSOW4Xt41pKsKnvpNZeETbdWA7EUepMvUoY91CcTOQ3sCnrWj7sYkUvIOggy57C06Kkhczt
aSUFgGv6iyuEfNkFJXXfbxZq1WL+C81ElIZypurWFz3DHFDcayiBwNIlk2N5JbcoQC+OZg4Gjlso
zq+RpWtnukPbth+rGFoUF7fspT5Nd2xgHoYRK9wWgQ5ZBjY6Z4Nlja2fsBed/RSFbzyXKY0R68Go
WxSdx7ULRKiCeyX13xkSMeosGxgpli4r3jEVws6lxdcu84GTm0KfOkTYSLouiqY1VsrA54lrel7i
7mcSw60udB5COwZBK3mrYPT/jpZ6hMePWl41ohC1qF8pXr8TkoqdeDtWxL6KVbG5WYGllwXaTdXc
DvJT/6Y/O0TqWDZk3Ls4IeSQ/Be9K84bqIZ6Y7MZbQgH5niW5rcSnQqvgVw6oo4bwrk1fyJTckIO
X9hNYYLAGaK0vrJHLQRha4dJnK844BdSgLYChP1KRWodvNLoSGVQISs6tR/lfejJ34yp3w2H9nXR
x3NQ+s8J0FClx9XpdjGzrks/qcnpxyH7tQJraK8AVMkyHJafHBIcc3jRF7n+KjjQ5Yxyrd2EaVBX
TJpDw6qCH8Bp3Prb6jCZZ/tnragoJQE2ZbH/HHYE1NS+gw4ObP5wTWPn6tvV/f/1dyoalSvNR0t5
CK+EqLLDCKHa9jWu1+Be7HEzcX8zO9UfHJWlwi9+fSLpFDIU7eVg8lx9hb/fMBfuhLcWx2koOrR7
QV51940wsWSrIffzOD1Fx0YNMTfH1LTHvmYoUKBTomUH2KmUyWx2PmqxLcdNPjac8TqNqa9JmxSk
KdLJQS46CnRoenbi7WSrBMzcdCRe9SM6zyyMjcTIXZ8NyRn0HzYUkds4gPW8QWxxUe2mEuis3q4M
824Ao9lnuXNrDKy5NTZSZO8XMDJdjSYrbs6PUzaNjji9HGmhF/HiRZ3pcvxqLdzeFU2et3nga9yI
tGO2/ua06bMgY/uKY7i/5vaATne6c+USiPvQPc/G6cdhJqBFJmyJEFJE7UBrpoLv/n2FSDRjRbgM
mOxwJbgGTEp/9W3+9pJ6GXlLuAFaIph6kWNDEhcXaG1gLnxT1LS+ExSz0qS+ab9ff/N2iD/hIb/o
8BesYmzpPPSLg/lORunflMHKaxdTujCuj7BrsB0MSWLkcRnS6pVj8OpOt4XdW//5MQTuvw0oRzOp
DQBR07hxI95cAIm62zHq5kJ6FfuFSCyhrrS7UiBZdoSavXkusdy/kpiGFrwV27MQTjxVKTaQ3J2A
HABgN8ifT4YYHY2UgwcVNwBWHAWu9LkGxbCD2a+ivY/hk+brGdqtmpWVmpln/7hZBTOQQ3//OatO
4gCrakZxNi3lrngUm/MZLUslMMGbv9wWQOy1EkrZ55Il3rkYnoTeZPrDGwCs7EpVujBHhYvp3EJz
LC9hNFnmt5mx+A8ff7ql+tD9TWWnLAFFhSg31CwzKNwDIEJEMb8DV4Q91woqoon8vJG3B3VKuexy
ylthIzUrKqgkWKhZlNSqLaPD3Cwp+XfwV1Yep9tSBOfdb3uF5m1SzLNoN+7SCXMds9qJicAiAnwv
9YtsKff1gjUAdIwAGiNOK8OFHsh9yC/V4Ynq9qgyk06BpbZwt0dpXPzN0fqSoURuLYgQKUqUH6zc
yYNX1EWyJTVvnwVjqamQFLKX5XPcwxJvfUfcPE5XTMEvjmu+r3SdqQNUiXp5NYfqi/pSAdOZ3CMY
RKReYvMxFonuOLKOi4d1FXx+t+M3x0y4a2/sp0JlNFUuL9MDjO9fQaOb6kutqnQXxgzJvclC2cUr
5J4wxZrftbMmlUWSvPjp2V7s3L02mSLA4IWvKoo1ta8rX2h8wrgkGqpsTTDfVknXaGxxau9RaM9z
Y2bKGF005ZXMwFr683Yf18uEsgzX9mv+LxhIYm1igHNETFRKMezYaAjdTm3ZOETLhHsFp8b/a7tc
L7+qgaD9XsQ5sR+/KWGHO7zN2w0tv82ine6cCO9PML67jpuErCe2T5eC2bGbPIpz9uB8rXuLlj1v
VcIp8m4j2qepAGxpQI5N9HOkXBEkRV8KK06hZGuBTkp3dvJAW+jOHyuge9Y8Qp2OawkqGKZgZeCi
YrA3Q1VAXGw3JCD/Ne3rLT/Qz3fVZ0Ublh1wIUAWZkvtceMO0TagbCQsUlSAxWeB00IGDzKYKHe9
hWl5qfI+MK43nAozSA1qcfR8CZ8NFLUvvWZ4IjyOqhvrVFLIn4eagIGug/0nhqkcnAjxhjw2xNQQ
00LwE8ARpiQN3P2xgLgsTlPZcimjhSt17pqSMAQ/5stDk13YogaJ+zoRRza6gI/aeY0WdqPzG7+P
KiAWyGO/6bjY+ti+nH4gge0cRBbWw07mxNLVHsxofTejnllIwUgFWQH5T33rVEqXxKkRdVqR9tN7
cr83MSGwi2gq0zdamFi+KTWHzkf+VCZHkCUxQ5c+sZQFLcF65/W5KCAbzNF0FuUKF8yAmuxifmNe
w8wuy4vPvHwtAzq6qVJpa6x/kJI9slPVZyixyOa533v1I2YA4aDh+TJJdk/dgRAMsVw09WkYt4nL
aMtH3TYwA86OA4ycJBOgo++At1MitmmAExdkTMwCzOywhCsEq/lEmbyiK4dhQnNLcWZXBGAV64SE
DgMBDQQ8eFFK3Jga+PNxGgi3U/aD9Ho4ijMwm1IR9ZyCt+sVHwsR+oS6k4jPOR2WpECPnYy79Kan
Sx+aa0fJCgEFnOV3wOQEgzRA2yXR4jg0n6sdKYzqwdHh4UV6Aszp07sxxCPS2ehoWG6ItlYbW/3b
AbGMlyWoFE+6Ht7Yta513PYIuwcR+vtn9t5HuA3HwWCl40O4yvnBamEdBDEi41aHakTYB3J6Qbrp
sch1Pri08cY1rJ+f+eLm3BfJHGs8ihmckTUo2VZasKIwkGAsyc0H73Ilq5kBzGL0so2D00TF3SQp
mzCST0zvQvhoHtQv7ATo5tBo6NDyqRFsVOkmqevqGZUBgCJCnD6cwsRadmqhXhys2Ah3tvkYevv9
C6N4k9gt4H5T0MWyD8994IE1ZgJ7GsrN4F9wsJyQIOK8SYdcdgUGddXWB+kCNHfKFqgC2rq5vvaH
u8t7aMRH3ZR5tIowC46wcDjA/m3qGBDtJx6bB44F1kLcpX8sBaz/W86Ed0ChdNEtSRVT/LOXKpdD
pj/tfDxC0BaxGoslJoD7sHloyaYBYgmlioCykDEuNL4jlzWRciYN/6L4f6rXvNCXq7ghksT4lg8f
5Y7gc102Ai0g1tS4Yq9vUdqEtzpTE7zbDU9/dclx1aaGjDJFRu7ya1Xe0lmoFUbIOcfrZ/YGRHzU
fSyeXaXU65P1Y1HTffmyvIeLOJUhOQN8YuH38MgfJX+gtUnrUDezdB6P48CU37x68k5zOuIJq+mK
L1Pa90HJTR5Bm6hMoEfhcq7CzumQP5UyjNc6OUCFn92kkcd7wluRs4QU5PfmHSWRX7T5xv8Ul7Ml
kcW5Ik0Clx5SpDYu77IvipqgoMTv7dyINjzdrCmPJvpRqAa9V6TXle79hCQqbPEMHAKIMLORlr55
dM9VlllYdGF9xR+mwjuZDLza9w4K3Iz6qZesz83/6sCIVjgXoZerSMvhmh+Sq0I/ta29zckZfM4F
YkkxO3479e75OGQagS0RoVJBzmkxYms4sCFWMoiKk/1ldI2JxhSrvTmfePNVp4jf8tHqn2FhvfcF
c2xBgHEBxNmXtrIP8mCAyvDORrFH2RgnzIDBITH5hl1s+OA4kKPlYa1SeKSpRIJ2RRVh3mdwQcIU
KYrC8fwgiGo9sEhFAMAWTr5jwwlkBoZrRiZufXNxEX9Gl2XUv+HFxaCQeIqeu8mzBpemCKHURHxf
JGUziV1fgn+zWu0oZHxB4W7TmM8GK6Q/U7vrKAYec6BVnPMY4VQVfi/pEaDhduKkvqJuu95IhjC9
+j4vME3JJ2MEAikjHVOsr1D3jhangWpI2C1gb+BLlCDMXFuMHAygdrs3aoRwpFczoQ9hY9V1p7YJ
h6Xi9eYg4wVs3R7Lnivf8HY75D3Cu0o1PWzjgIMZJs1EUiLUdVhj8DeCqysWn7n/GtDQR+/pF7Cs
OqiK3lTnqvKMJd2fN/Jz2w2vHTSjAx8wX5j5pfHD0isWmXRDo0wB2jfnxcaaqWezwJYSb7ar1IMj
7745rfqf5VWALdpQmweiNiF+26ynOfcAhn/RHU5TbhJ5ynMHSBgp+gvJ/65f4EihmnHgUA+U4imQ
0VH8ULMp8cPi+vzIDMNXTlohVydS62gqjwBGvZA9DMpQEGkq0TaFjJ0LK0sCSZRt49aul/uMq2L1
rbiAUe/kPZmdogJodta8O1KKM+HdrAoMXFhB8/19LsNKkPWiuqKQBzXgZ7YbnUs9+BZf0+Yx+umf
/85O82olp40Qsv3WBV6fr6b74rRkzrcOs0HOVgwkILlHnqyJr4h88ZGoajdT55Dh5kVPfIJWYi6P
ivjWpgMWBWcVhVF070zsG/OuuQODKtAziQo6UyC2io4oh9EMKqDX2r7SHbd/PcyzbBnXxdphs78S
Ys5/WPhobt9NcTUOhbeVjMvmUW8/S66JXqOCn9bCXEtVsVPs0pY4YrUD4Ct1XXG3C4XWNiP7Bclf
ZulBGLHpsqm+HbHyQs10vtv8GzAeP8lKS+niTsgGJtEzef6il+ZzhS7M18wFos05S6sesoUTrScC
cY3Ax78iiyKQDuWrJoHa0ewy2BFIT+q8kbUFwHLdCnjsC0Q1gcX73qF+0PVdsetONUgRkN1lETxf
G4FmUedysVHLruln4y0V+uo5X0UWrKrvFnTMBMQinjF4MRz+/KV6R3GRqXWFba4uztCBuwvYO4Xb
xfXFsmy7FVg574T0SBioEo9mxKrYm7oF0OBmZjAJqHESUPztMSHyc+ym+SuusYnn93u2TwxN/vl9
1nZdecPFObD5ojZ612Fz22jxfvP8lJehCbdP/q2os47/sb0LebCLlGwkg39Baf2rLfQDdMOXdhgD
nGG+Otsv2fa7XLFCVysSBBgrF+IBhrABvEI1b3CIRCAGV27JC2QUgxaBiCWpQu9d634QguSKays3
HhKQPUQlj+l4BeneOrVJpgUZY+CVlxWX2zLV7LB2oBQEl78o4GkIdir4RQlv0aCIEQlgYHyoNXUz
kpto3EqUvwf/Vpke06vpDtB0nyv/HElOxTIRK/9oi+TAa4gYobIAONzE0lIb27zalyEkSDbYTjJe
QEWriEjuHxtLpCt/mcBbp5+d0sBHvGCCghlUrVkbB8yxd/VnHl4n/gNKB8mF1V33TkYLsfdBpZ7O
UhhF2gEs7ourgi26Mp69HEDzfWFN39ySkfw5t/522n+J6QFW4f0xD3fvFX4isJl7FR+0ukztuZnG
9MBt011lyzQacOMIVCgWForfJNXYT7N7NYnmQWWMihX7cptnBfKhSliiYWKmiGoCEGX3ZM1/dkin
jssovDCwwF3qr7Wi82iA2Dw6jByaMNEeth66NPUQpUJdxVpAwwpVX1iG2qCW9LloPjMtPNkvTBrJ
YZM40N6ZF1RI92UJhLki2h5+bK9s+h1UZcbWj1l6EHRmj51I9nX0TyswSm+wiMV8qUfzkipelZYK
+/tWj2csFH5yqBoyjNLOhv2MCQq2zQIjZgZege4Heh4LHhCgazYBUzl/cVXJWGUt38KTmppdRrZJ
C2HvmCV6RAhYvkXVU4gmty4RDn9NNHxFCRHCL8EafLYhy6VLg7v3FkISkTD9INNF/7YKSAyyr+V7
uauhVx53pKz+A0ZA6b5HyvdkikFPH2PEoEmOJCh4fZx8X1p+uPdYXCdtjT77FVSpb2+mY7UGrQaD
FJOVw9SlO4sqwuW6UcWee+tICLjV0BE1FLeFMaTDXxYPLAnrZBpZEIcr4+V0ij5zZ1miGz62x5B+
PRWIBMRUIAKECwTgRVoP7UiiLuwRW7B8NpCrpInVGGWNTc6FL7+BKJhb/7Os2+qGUquIRMn6aRzy
YLewJ9ZVDptSXPpk3WM577OK6/LCmYCDonj9ckEsEaM+cCHwEpBDTi+fjIh8w6BqAvBN11FTR9+m
OuCA6vfCtAtoBnoCYFeEC+sMiR1/k99Zgjaxigm4J6rv3ZVOPN5Pcn8eqDvTbHxdWxKpcsqo1hSJ
/HYkApdGUoEK3mr5tUNAl/7KvPLcvVnRu2QRtDHKRuTDFnlshMVDSJR2kh+DtgXDl7Wm5ZMEZOwp
2I/gjXgaSmsGdWGIWy786y4sIIlm3zT+byyTW4BFCJMbDAWOAl0+pWvrF0jsPqjEIL3yAHscK2p6
aqdoAhdp5u/s/8ShqhVjnPmG8mntK5LgM3izyXcXibMTkDLCHH8sSSWnM2nrU/AbKcSOX+qu3mnv
MifjYUsHKRAUmZLWYzFLsGtHUqHvhwf7pvdC/2br39eChWhU0aoS+djgbWzfYv/ZJ27fgpDQlygf
iDbXSNA4kcRH97vjWpEcvDrsAoxlP7nQpIjd92HtlsVHVWd9a0WymwyjmiuMwEOtLN1gnCh0V8rZ
P3ZyfL/JucxeMTb9+0+sP7UM2PLJrKxafJi0JLrPik/hMpEGY7lVZI76XQFLtAfMEf2DbqhN49CK
la9gQHeemF6eIXxSK01iw+AYt1ZhysuOfC86SeYohYLy2jy01ul5Jahw5uT8UVhjYmZO6qpf7zAv
MIcOVWTgo+nY0wnNzIvrR7+WfEeGWVijuzVrZJrIHMjLLuw6pqV19DeV6gahD8x5zB8G2WER9Ayy
ysW1ox8iJ7QqO+jWGo3R7+ACIcIkfq55i5aNnEirBRXT2f6FXtwu/2RaaCHP1iT+CSXPaIRpyQOe
ZIx3R5uot9tqSZ+qr9xe9ZqpPDDkhLRTpFxXYcvuf+60DWrKttFp77FwISamgBdReFjgbYawFTYK
YqOI62uS1BrFa/G2ZvgEMWbIxRCiZKWW3e2ckjVSs0Bk+0mHz4KHTs7feY6jF8Y4BtSmt7n7KREw
qsYbV58hm+1kNjKRRqHn9OGOSCgGAsZuFvH0G2JU+zFKOzUg07b4fo0uhL3MbEQV6z+mIbLjhLfU
TTj6QgN8g3adOvYfOLfmSdQ7K9S2RzG0eMaJyAyrY5rtSSYS/L7YlAumIREtSgywE95Yahbp3s37
fw4849K3datgH2WVoDmzLuJkBjKaAKolAAkRjtLbPEzdVD9aqPiIaWsmwSMGSzvK8rLUwU+1sN93
DP0jzqfbSJV4so1p1eqkDkw5Yq8HAFKn0BIBsiCtnf/WKJaffXGzcfoP/118HLN1wouEKhRt1Ldo
RhhIhtEo7w0X1b9xXWVY/CDeciSE4smVSbpyQRV7rRIdmGztlBw8/P9YbkISjTDNpV95KnxUC1hX
kIMyZJ/YCcGw6hKIXAvdpzEkbbXhrx2lO2WaGSh1E41DHS/fkZf32LcJ7IXgbKn/BhEM6CoWO8gc
o5B1XFGSbdlziJGISmzuOenlQ9m5Y67vIVNoF5+ef+1mLzfSB6tKfKJCvRcGctVA/yyA2DC607E6
GNR1XD+AsytTXeArKp4edeXqeuu+cdWEQ3OrY2aKN3ehVkFnFFAP9K1Aazaufs33xNsvg2GOhuS3
PqB1KqearqW1kKNiFESlqfZAYkjk3/HAJC2yCKhSzLB7ZYUs89lUe0QYCGHXiCDRGoWTYLOO0PL8
WrD+0nC3yHcqpM9urbjnN44DYqHgcKPm8IpT7PnRpX6Co8BffmqsrkO4yk1G+BXZjq60DyIQluM5
2/24GcZT4u+2lCLkS6/Ei33uebFy+wOXKsu24CsujFfDPxHDq4VeYK6+/K53vBKLQfMpT/51guEM
ZMx2B4hOzfkG8Nv3Epn1Nhp61zE1mPet+9A7f//3etw9+8HWeyqcSZ1YM3smSUecyxe5HdN3gCwp
YemEfTK34gKqzzfpWpe6wsomA7VSkfqjbxPe0BeeEPb9Sx2K0tAFOuFvvnHxcBsg5C+T+TMa8fzx
Wmy+gj+/TDA/X6zIS/i7OCq9FVxuijp5TSYgxjhMa3uWZBrlv/UXiEmAZ6AAUwWlW38+DretF+++
3k0tHS9CG0dxGLiT3TkDHnzDtBl4rk492JxrV3I1BZqasmWgYDM1vC4Ogtv6f40ib2OOXlv6UUOW
O0E3qY/7pxIf1SmrSwiZ7NJbmToXayHyFnGVolKGxAm4lcvHbgeNpHcGkFnZbNKZdlv8DynFqWup
kGVoIOPtg0ONIpFiF7C1vhMqLzw4WDopqz7+XAMM84BhgxBkdml/+Ef4DB4xYzOz+D5zdEzrV1BV
Ufm0orIwXg55KeMJPKWC7IdOT/DMrQDNNvLU5ji48A0cSn0kSeBY065vl7Swnvk9K9Azn1JRpg0Z
8x5OQLFVJeV7UBw21868PURz22KcvLxhHjqvD1fe/AGuo9zWOhbxt2NWTNH0ZMx5018NqemypiHa
/W2LgYXf/T70kdU89B8qo0DERcusRFtYdH9lkcUDezMXX3PQjjWbfiLPRMaJ1vh+0M5OG/rTdLdN
VJLFjgugmVIckGFtc8bx6CxqZeh+NSc7EqHobV06CcmrFE3nrsULJ1KIna8q20iXIXXmNFEW9c/7
EHo3R+PjAHsocShyatxLYbGTJN86wni4BDvPjCzaxh0lN1z61tmtELJZCZXFYYS4NWcuI14ff3Eg
LhCR/MuxamruH64lHA4HZ0T91ys7ffXZFoGWFfjNFiIvOzcEmddd6WgFpAH2a6hii8LrEx+HbqWm
cCuhgbooPwpPq33q75C/SoNtihT8kjinyU9hAPO2lSo1mlWg7xZyBSZ6iye2mD/JG12YTlI38s9p
1LpvWiogCfjrESaCYVaxxj7TQmECVEpUYaxhTFotP6lvy6crHGNlQuhcl5b3+Rdd1gDiCd2vNFiF
gfBSZeFdfbf8tKBB7JqjC8XqGO8P9Isb+chbay+tQZC6hfrBRGkWpZGsNFYHA8jK99cL9XZ44by6
O94TbaIT/wTPcqfi4ts+9NTbXNv/UeF2sqiyzLLw5SzghN03pWZymE0ZN2Ih0GwKotLidOvl/T8a
9TpobXWB1f+BLpemx+14dXvwNimY6PItaAcBB3d2uojR3KzsMS19I5w6XGTpm5jcq+QPfUnBmYev
HDDKOEOwp4iFROho8Pm4YpOXIm+j065st1tQuke7MLMYWLhtOe/aTxI6ovxExU9mA5aSJyec5jo3
1f59iobHTBHSyzXYLy9YtEGpgjCuIX2rAPzWC2RTvI/rxNwan14saOXpjWV73ExbjIWD4z8yZLLL
XPmHJFXZSGzhiz9o3oqKHfN31/xs5zZAOMF1aNLavy4UOakKzVhFz5pbgloG4etq/eQ6lFY2TlTS
f+1sLcSlyd0q+j5usSN2QJCXXHlRkLJWw9QdlLI9Fq3W4tokMAhwAlkiSS6DtKTJv3GYlLdk8HQZ
DPaVNSv/UPntjrbwrkRBSUDyqk8Ocz4jtSxOMPvOeLNEayj9LsY3yQ5+IwlwL3Hk+NYs01v6oGXU
SsN3vK/7xK+CB7rCSKNF7D1Iz3Dok7xYs47RZR9AIAJLY6HCOlnIVYEOLgQJC5Bm5WDMiCgdLH75
Lw/zmu0CzzYOmxyX6ZW0NBJVyZLGTji5nwY9ZGj9RK6g/WyDlg72mlkXHLBZMf4vQxAzTLpYZ9Dq
rjy4gz56iHrlrrqwNwSac8NTtj+LFD4nd8CZdt2nbmCw9K7uDs3oC7aLnVgT36Pjc1Tjq3JDt4ob
dq/l3eZwzlrYBCdJQk0tR5xJEiV3YbAhx/hmwFm0lbh93+aTZqxe+h069NbIEWdobFnIqAdIJg2Q
YoQntaTw8iujzTgzufq0fAzGLN1YqJq62MgQoZfmBtUD8Ohx/TGd0lwRCxdVVFXKlyhGFyZvxCOx
dgxdtqkEKoN/w6mHzwv0Xg3qhVqF5zHSgP+bsiNEw4LyndXdXYWt4KqVQHLeCNNgtDDG0HUlGa8H
amYxLg4GHejk7u3B7IPsSUR7fGCQgE/5uHnQ1I+30YjjW2NLtxtscyRfq5d+nZRrmsZAVfTyWTtC
Goh8EA6+uCvHEy9WEWfgC0w2x2hN3jXE9jt2B3eKEs4qiP090nwHCrAJXA6I1pJygvz0tGzEwM1L
fy80RXbsNuPyg2guE1D9cv5upAfKW7GUB+yujuRDf7DDWoIpXvgvUmM3O3g+dyb6QW0v72qNveXQ
avtDF78PPsj/8hm44fkdsb2BgJrREMe7yTJehB6/nIdMIvBHTrj5Xj7JYVN5usCrs1dxG1SAUQd3
T7t7oy0k+ivWinwp+hF5Mb/UzHU7LqoGLfUMZbCJ4+M/B5GKX6bFOgWw+L/cqlvJKkTQ9g9oRNZA
4w9akIC+pXrwlmXYqTucRR2g64X/IlGA5wdqmTLHlfpKiRwdYBCajeDS/vJRLYjV6e4iX8aiijha
uHVihURimbW2UhC7yC4iJgmgU+G/xlCBP7O4DrLhEnrFJ1FapqlxvYJCEo2aXR/ixRaoAEZuhCa1
yTmGSEbWTOuBWWV0XNIXVi7Le40kb63vFCRDqSUmB/hoKQQEHNTWiserHc36uwBXB61afJZimFco
0kE7gY8wvTylB2OiPDaClEJ6/Yq3eBO47fMDClRNF0NOArsHBDNaYO0Ogw2q5Z8s5P2iMhp7mOOd
wW875+2bVDhGlXlvPAUmsTyd+0stDHyEVzf08mD5fpjudzTwFmbgUak1XCshXdoeut/gKO5W6SoD
uGBU157DWvO4bSYo872rZ+XyZpEb2a2AdQ2aeb+rqVgfYZcArgjYzrc8km2h6M5Nci60Ys29QI6+
9oGoGJMLFojJLALf+RDfSURTIbkbULpFCzMD5x4Yjm+YyfW8qAKEz8RGSjxTND0A/Q4N0vEf1gox
C0Ky4hz5ygE/1GEarOGN29zEH9toS3+l3mMQKVHPBObo04kq+XuiajssOLaScq4jAm7KXG4vBOBE
DORbYqKMm5/5z6wzOVQpEHE0DlFeeml7wUZNSKOyy208oOhzO+g/u0xZxJklKp4+RRbDymZBekTq
9G+TbhZf8k6p3UOZaGG1T8WZOWV9ZWjjy9oReSuJKaF3cQi66kMzDv/159+QBd1HrJP85m6y2Pdv
23Ylyf/E+3AbbOs/Ttw44S0u0umugkkf6uGf1d1Fv9fTlKbkefUMPxYhqiYb82iHOx/b2LGdJWsi
8BQrobiGz5BdGHcekHNhUk9xbjakQafU7zFeeivyDlxPZlAiUWucB7nR73uuCrvaHnqyklVB67KX
sSUXCMo1mHHkMLxZlLDMb2qMwbL8EoHG+j54qV0wGy8HiOP+USq1ucNHEln5q3DmFSZYjAS62oYT
zUv2chJM/n8sd4xh7jBg6x1w7KI/mI6hVstWcaaKmEJJuqcsbBsiVt2Z4kFcirUIeY2kIZuX6TVF
FOuFHvLuetH0O+SBllTBzoKo7oehIyj7YNSNYT7SJ+7ueBv81rqSnL8bQ7z2kyHCjSXclb9LGptd
WK6YK+WNWs/h/2CCNSPf4DW97bSV/XAnZGS7SSej4f3vV3HRvnwe6lR2ssTCBqaEzjKhlYdmMJLe
H+fl8F9zMy4yuE53zvqWDg11+/30V057r2Qq68udBSTCTA9fWpm3UTDCORnbq+vN/yqYHqPRH5L9
KEpzwbTsAo4uifWhv/0BfzVXWOpIjHlDkiL3MGAmFsW3iN3nM8xXFY0Nn5d2zaiVGshKXrDH9QoL
dXts+WaLo264lVgqy5SLVfNnupZuVU9H9DKUwA8yxVGrZaLu7KOUOJ1ugG8G2VxtQgcjUfsl0zEe
jNR7SbohXTcrtkF7Uq9JZaqHhytbWv64nYYxvWAmpIb9wIK3cF5UeT6ENiRg0c/CFEQer1FK0dYx
TbUKUWeXWdscXMyStek5ia9pDAe6BX8hGNNY4vbaHdf+zqoEgx9bxSZfZqYiGmdXqaTx5y4voR/A
3ocnxpADGBdzFgv3bE/ZWLnQ0mKZpw9TNGg6Sx+Cs7NZCpA56BOJyO5NitULj0MSYVrELM7oI4IF
+DIYOgRsZlpokUvwviqMdWe9Z3x3kR8sGdDHtYC4EhR8c+uC0SoLV1hTVssDc/xibF3J5v/kpJRg
Ht1JgROnJSh8zOOYjnmVTZbWAZxWKzV3ieyBVGeJ8kIj0MJCOaaVnRtp/ONvz2e1jYbYdZvQz00J
iNg8bPKdMnwOGttAThNSUQtJREpA4gYCPnphUaVhDN9GJD5i8AZ5W1frP2P4jVB9d/LsQGhnYLiz
NPD7ROA6VFbprUu+KDaZNG/s56o4s6fCwND7y9dHBagin0zxS8ykpDmrPIPTYrSBDnGU9nWIhe5n
jpyn5YZHeeMPUmG7px0vVB8tD6vyzAzAMJIQzsEPJk/yJZgd/73Aj+vfkYG4c4OX7P6xDSrL3pi5
dVE9E32tKuet5IFRxHtl8JYEwf6ymCavsKTYxH6hsxaDh0dhJaYqzCFHpBEqNRLspNBEVkAqbu61
IQininyNoDbUVpfYKepGsrBb0ZyZOkQ/5F6As+3J8HigtAGrya93sHgODLNSUTZTdShgHKlAqDhc
mzW7vWec3Zrb+XEmwP0646OwUbh9cxr/001WPvPEnFA3HCCBzRRs8namXFa0IazcXzoGzs92+Eo5
5kfU0JazaX2+UylA/QWkXQNFyTNDRcOgguTbBhqIJWWX8aOm4b2rPiVdv4FvnCCxUJPsu4QtEQML
YtSc7diaAYoxtp3V26MpOSW7pL27uaqR1bjAVk4DKumbrgW6wNDBngb+amv/Cg7GaAwKdyUh4agI
CKdZk1Hc3WgkTnmmfb9UGVvyA3+9y8vQwdsfm+QXwhrIDCXy11IRmxtCHJYuGHXsI0BglCM/EwIK
BntDDQ55/7F8MaHVAe/38YSIEqrYFI4exwb+6jAZJhSQ+NGsvMI0notx90LcbMvLihLHpQYX7vNU
Yaizg7KKxAm/zge3zu82ZlqyiUJQBTHU3VJPrgqOa54cTWF/FwYXlgY5xRC6goVfn+CqSLHKNCEV
eplCYEwhRp/ow801uuG7+pXPz4jo3lkmfZ4cvb9Dy7tuJZfzP8lHu2tX645Z2p24UoOtzFggCMok
0Tf1PG7j4hB0QQOGPKoKrWZRrKXYligETrjNGwR9PZlJGkVTl7rsIS3pDAqcD4PF/WeNVY+AxM/t
P2aNyHKXC/E7N78z1VTg/PvWWFZrKpASVml/2L+svI3COv4DS9weiT82l4zWnf/gzafaWF2N81sS
+rKwsP1JToM6ZNeGu7tXRJGGJT9ZHQlZptUiQDw3rFQ+cTRY5ZQHsTx30hZ/8CkOzJ+RrenflVcT
gZRDMsvo+JkOeWEC09wZFDa17Z9hh84zdjLSjyjPRxNXDc2EdjVCwk0L3jEpksQYv3yzBAPWU4Gy
ZS3mdi/GIwm4K0TyZfogKAPoRt5PuFKgwxt4+RN+TYi/nJHPfMEUfkC+icwh4XJZKd/OddQGjAZL
D/4JNveaU6O4aaKzmuVu+VDVDyxRgDZZxLq0bzxiKoW/N5UUTd+Usaq7E2o6JEE6Z22Z0CwT8SR+
sefxHXbuWIdAumPzsKyHuIPSPCyRNJK+tKHbqbN99cw7HK1QS8bxc2q3jMl1T9LUSlrKbWhqFMdm
Zn10038NzsK0YzqY/Jz6lRTJAiiRPfl7OF5Vb0CfRlMMTuU9Is5LsZjC2yOnIJOrSi8XFbbA2zGU
5uwup/4ndLJBMqM/atmmA0eKXzEeBB9CgIX6gcBipsBY1sqCpvcbWj8TY8wNUTeK3CjnzOr2E6fO
n2yCVEsMEjzawcbeL7qGUH67R7Mwpn26nmRTaxmZnRe09rvSVy0uRYf2x6qgN8J0HTjmGESdVC8Q
WBV025UggQi3HCAer7b+IzcNaVmDZboaHlaMWoLw300m4Kl0wUDVVbeP9wUAJ1WB71GEgFKV44fW
fLOfNNuvxCdwndoIjTO1VGm6KuCCj5bgMWLNlZ4VkpA2rBWjvIIQENhZIA87WPK1fz/xlBdJeS+y
WFg86q5jq9ica0ik/xDyJWBDOV8s9LTQxVZ6Yi+9wmnIBGLKJgqfVtlNnYTGVWYiv/o7ekAy7amw
2m0FakSdeFDNRtgZoLSWcGbEDrv2EqK8hTWC25Uiq4UqTMFl+BBWj7Sx7yA7O1DsfQaiE2LZYiyq
8FlVWqK2HmUxB0rwtf1vXc1fd25vIaB5/FOB8mMcbfQPGchzffl8UuQ96M+Erv87P+0viUSNgA/p
17jB9lsVdpo97LeQ8NacT2+f/lVdkVB/T/sSh+MoEqcIVBomX4kdgK64TaySJjBfF7MxtLsKHfIV
sK0tQAnGBHWFzUtavjhmnac68bYzdCovfvvuxduzOu1jjpqruvGaZVq/RZrPBSj79+iTN7HL2SG0
27NZAwRmVOlcrksfRWgbm1LxpG4i7CQOX/EezRNrsqsZYQe7ZRJaW0Kpek6saixx2HUBNdyAn2mK
9dVYBaPik21QyCg80YVSTZXjyZPvnFYgyEZMwS4Q/X7iZjeTcticBfMyxJVy5Ka//cg8ib1XJM+M
apghtCQnGbDSkeIdqHU+2nq+CKsjVHrnb/JVKc9xfHLyvQolm3zTYRztkfdPXazWF0anzJcGyBH+
jWJlbdCGW6OAKg8q2AnRKmGeA0Fdrj4dEhoJoxyVQe+aq2CGC9QSCrExPUIBxDA4UOOX8x9rvMP2
9QZ1nZQhd0bzNgz5Q0+6w44UoXDHmjBnKqSooBxgEjvsQ1I3L0dl7go3Mb7v25QUuqGxBweZ3+FX
dSgzxBmNqZwMVvMOBahWVBGOGnlMBEJuXSrlFjm8PJ6NKxN9mHkct1Yjyl2I/TdcoOC/EKWwdcEE
maH/F6iwdqW4Uz4OHX4pGCKtjaSUXf6AFhvtRNRd4RUc1nZ1QbDSKHGGCqQbJOx3qWE8QnqYKjni
xX/5+YkQfFSSBQ8QSUiSdHDrirtkLf9TF0tfqUChvRx7rIwpUmgV0Yu1tNdXdyHbWWXhhGd5DD4m
d/IrJZfgHVpU7NsvGvKmVxRHqkOEVdVxajZSA/q4R0qp+SznDb1QO/MziRC9hyFHSJU4aqjX7lma
tOS75cp1hSpZSrsNrp8w99jjnsh54a+nKd5OzB8cU398ZtWrQN8ybj0DRmeix0Q4w5k+5R7Os51g
z/sN5QhEKOnPmtUtDc/G2rMfTKFCHa7J0HLN1zrp7VlnBZZ5c1X0Npimg5zqzGGXODfHhZ1q9QJn
4GuxBAT8Fiy252eQIFwi/p4zJff/VmHZqxp7W1Qt0oogYX2seMHjtj8Jf8eTMBXECK5DpX1MXaPn
gwTW2WHUyLqbhrfGHfM6/hZWcnUjVTbIHR2T3/v9ZwnjMc4fM5vYSfZ/bayBWpRyPpQc/KaSkokf
vz/sXDvvmv/zyOIkpcLiIoNLRGeAbI05lLx6ncEph4qCGClcckSvmggQw+W/YmV64k3EplsKbdBB
qAogFq3aEF3A/UZOX2lvPG9BDO2i5pzcP2BNu2N1ASuC8BDTpBCsXGJD7qRGacbiAIkIDE+wrf6u
u73zSbKh2OWpG0Nsl51u554FRVSSkcLCCEbMGlDpjI/5tcwY133e5e0Xp5pqiDk4fTY/KrXaDs/3
8yWbBRI44aOKKdqFWqFRAn/lBztUDBSl5zxi/pnXFh9zaVpw3BJdu0hXsI+GCKJNd55sOVOU2suU
7WkvMUwiU04Wp1o/6469WcG1qVsFwk5/Me+gs3pW4mp8OaszMGjkup2C55PGi9qqpTf3/jndQq1n
rsioHd7psu933Q28y6eb06RBjlkVhLZf67fryYeLeu4UjiMw+bCLYIuisBaoc5WscIHaaeXzxZFJ
eczWcjqiXQe4gvVjKMIax/uTIOHf966+/V4I/hbNuqovO45Zj0IT1VsB9hFJwvj4QpWmKDTHjC7k
PR/ceuhkRw4v65gUthb0+/SAg5xEv0ejzRkYIqwAPCZJtpyonll15Gx2KX6O4i/wpDH79aGHyVTJ
K7iG4Hhxi4VCrz5lYsZfxnQK4PDyMHHO/PpDcFi/IwbatlIqM12FzXFrkpZWnVMiOtmSvDHy3xPn
4BPNyPqr4uLqZWS51O6suUwOQ4cOWkEBQgg8b0by2Q/1zbF4sIdgQwriT/O/a+kZzzarrf3ex5au
sAH0sjdkNb0Q6EDQEDB7/4kPesWgL7zXeUcPtE8beA0MleCXJWRwOnd8Hgr+PZTRsa66FgtE2DbB
+CW2Ix48xgAkYk41Rn8Q6944Z8SfkNc019X6Xvy3KOxChBK6TPRlX3pedRuaa9Qsp1JAJVYY3UD+
Su9MYs4AH1GuIDVH0SFQaEOgp4h2BN7ATz4binRpL2PrCBHu0gozkvBfCJi3oAp6JzaZgX1gPm/x
iC9WuUa7YbE421g21eskxQq1bx1PKPHVkDWdNknsrgWcAsigKOWQ+vfPJ877h6ALXnSyQJKRq9dd
UR6q/xMveBKfqj3NQ0N2bIo3L3pcrOiat0D5dtsaYuafJqEh4AW9zDHwCyhk3QDJi2qgWRewaeXn
FLAhlmp6I0lGhmaP4mdlgfDo/o7SUhGe0ZrvXwenfvuI+hPuHHjwmC8RpGm4NLcqxzdc7OvjEELv
hPASVGbOZC+0PeOHW6otPTV/sW3LCDYRu00cNLcD1sFGNvRo9ii3+N/p8fuFIWrHxOFkagynRUyB
+h2UXA1CdXSsUqorLHUASiDCitoVz8+yoOlDdOJ0LaaGjev8KPR1BeIMnW9fWyIkAtgwY26AjgR8
ua07G/iS/+Zg/fO73/0DpKaQfuBhE+bhCXx4rMNMiw/1Qt3eeY1PzYaG8iIRWULgGoE8I5rL4tP3
u331N/oO60xlK9n7p1roXis+QxZgWz8x2KIU4LU+uPA/ZtOPFoa8hQrENnu2Yw8D+YQFcU7PgjP6
ZXx/N8uznkv4LS4P1kTGiQrT7mEIsRIy4KGwbUoDYG3lume2jMShStxOOJgQc1pO0o9yBo8Xp409
/YDO8JDf6euYGYdbOOd4xAraY1jHJd8tl4GWU0ULKYJrrPIdWx1cN5/2p+Jy3/5Q1AQhRtNsG5b5
6PyQCSAB+n82D59+NcX7CMz4jY1nj5D5CFbrbZZzMcW89PxZFGMm04kCHroQGe1s60n9LplHc/Fr
JgGL2ZGaZRjYvVpgJ5ki+F1oziyfi7EhchR3dT+h4tePNUcREGLPW5wHguwJHtYCuBK/XiO//CjU
adjKU1SSafrgxKiQhJ8cP4/yXDfJBJj0a2aQAA8XQ5QZkMoiaWhaEoqv4dICDp2C4j6s/AQL1Gzj
EfUHSon4OincFP0WtAtAtWldIMHexLo5n8iB0/hPuq8FuLvIpxR+Q8oNxLlZbXyhzT8H5Hqz02ui
+MH3uOzbysRjRyOxok+v8liNkFx1eRXEE2PgHB9Ac+IjTMKtyr4O1xk3mcp4384zG+qTFdl38NYb
2k2tgtKwfl03I4z4AVvaAoARgeyqhx+SG82T4OWGkLezlZ3QHKoITT+d1fSpD47PkIjUydWxwHBj
OZbqDH2dks6r+j7sv24u782QEmvXFT5zkLGAv7HHfxBWbQZkf3abKdSW5UwcWTw4079FtJLesb6H
DelraxKrxM6zuNHFudYp4inR0tmJJd+fae6GMPEta29JQqZVuYFqYZw1KAIqKpXfCeHTNiecGhGf
6jXgd2Xqt0BoCqxYa+WAYxRZ14Oly5wjlLw60GlyiMkPtMihlczCG1PFS3iD6faOUaZD+sKkACAI
QBM3nBeoONevGFKFEg4Pe/EC1i/wJXhtTSIkR3iawmfjQEXLvJO9kLBEIMRGWCUTeY04sq4I3qlU
+PGW996ID435RPxMFaa0aVawj8wm9WtNgVcRDjKWf18J9ilceVHFfzC+CZ6n17iv2tYR/hcUUUKE
MRodUCOqfiZmn8M28N75qI7nCXx1lvdaFROBuMbGTMEJMQPiLjK/LQtpxGren3CO7YnK6Sn8EJWA
DFRqJavw4SKs+b82mvHZD1zRdfQumqvH5tmo88Z8WO8gPUesxDSN9GBgLKWF2fFqMSAI00BZ1LJ8
MrUxWgU82LzleHyn5EMw8CWd63OFZWMqS2DeHNJYeDA2Zx84jFW5NbdwXERr41IqXmf8hqTaPuWB
jEvVEkBM5gUPKq8M6/JLqlBNNwQp3bCFIYfRt9dC9y7x/hjknHYB5rPWONyhhdTeOhIe7QXSuqdO
CtoHSdmPMd91mII5hjK6qej3DM9ukRFIuDuifALAg2mY5UbzYFAYXv/uK32dAhM4FltiVX2EGrOr
b5JbAIOZSjuY/LJqlJg4lMopdaY9+9/1pslYK5TSAu3MwmZlehPdL0NChJ1ZDiScC0IJ0JxRVtCy
oGsILSYZcQ+RhDEv9066LxwpNL1R6T8Dv8ShOBS65Kikse1GEBC9CwU6rxG4oxqqHPObhpqGaGBt
m7DoGHnfTGF3JFwgE/NsicfcbKzUUQDyO1Y/ZJ95Jk1oyJrLerFAb4qN7bfJpwMnnptV8BrwRdVU
on5g6mkMc15UFh71RnTpG0r3XBdgYfKiDiwSjboRyc0oOG8dGpO5pesqViOAD3DOBUEsu6SPDv87
mD9NvIQBXC0yQ+j75Uqkwc8td3Fq1Fz04Ik7RmUsWIqzPSIoAaTAYwR4hLbZZ/2e2LJPnP7FgfVx
oP90J8/2ssiQO8T2vB6ClM4PEbh9PH881etWhyAELvPqJWqd6XRIu8YVGYOJk2hyx7Eu4BtoPrum
wkBpvPknxu1Nvs1a477FoVn98sXmkPgkkB5U0nbjM++wvDxFPfJ/JW9M74C8cEeJNyEyoBiqK2yu
+wvEa7FPxkTHu+mkacNFnB6/GbyYq7Sju8Hvh6XIFb0avyr3DSmP1IN+nl3hSnr+SJMzOHRdrOaq
f4FPv5VmjzV6/gmhbZYQzfUvn2K7W39gUL22i5tUXGcvbG8UH6urmdM59D2oEdBd/JfLZLg/G9sp
nPBcOkNmL58VtJZoUlVsHe4keSSGldesTtfy7xzmdu8Y8AoD8kcPpfGPXE7Ze48rfXEgHcNOeH6s
2ZJhKUgAKLZRZFDWPs0A/upSkyBHQ423QWAdivBNg3cbfHtdsFDqpqwgVZL86M8N208a7st4Q9o+
1iOzo7JIovYloO7y3x29bY+80H+dJ6pfDZM9RS7ranODHpBl8Yw2eOJup4E6uvAojNWhu8hq0R0A
a0rKxvJzsRTlXpsOjFSzF4gAnX/suxR0wY1jpJuINYjFEKL1Wl/yuz12rAKhnmREApr1BKcYF9RW
hKR99gusuoTerNHPL0qDabIPpH1W9s7T7sk8Z3xUhYq+M/QgYF+JFFIkG7QBmQEJJil2dEKFRveY
omWePREQGhySOJkWpqdN7rcKaZ31ot7l7/1Y8K2Ow+ZJ4oqCEbmyi5TnSPIbHaPPjFltPC6GBM2e
Z3wBiB3YIxyK8iMbW+OYlgMIuko0CGNQj972MK+5FSveQ4Xyu7+8lt+Sp8IsnLZkphAiGrIVFytN
0oIM8C+65kUdeWzRa2rl4H+53HoIxjGxxOIUqrloFqoM/c0D78SYjDq8VrNKudzZ56I0+HFJmnJR
aHe/JiBPFo6kCLTN6wQvR99usJdEgK6dicg0DeyQeINAx0ABwMirgzjRdC8GDwVnVggIgakMCKmU
/VcatLMMFmX2FzZILDCCHSGV/QS7hSTDd2HK6rp5jBXa51IRVPUaBEtMiSuwfor4Ft3PxjCPJ2K4
ZD/umpRKv80kQliiB3ou9WQghcYpiki9FFDBlnu4UoQFJGNkJEBVTBJrnF7dX4TBPH5Eo0UZBJoS
DNwpHfmsnbOuc0fiWll2Q9zyK7xVF4PUhVu3CuBaErY5VKaCi90J8JkZcJRVW/qDufgIDVSvKN80
0ZbEzdyfXmhZhsGKAtsQ9x82qQKeVtRtR+Zn2L233qQWmhg2DtMOG5tS0dqpxOI4XzF4Z87xVQ8Z
TbfID4QrrROTVj+NCBUZ6camAhDnJUhqv1wknGyIX36liCOLLFw+XXoyaGpbZKHIjyKAajiPh+dn
UqW4wm2j+9OTdLK/W9pv7+EQ8UgPO/qg53z/RwfU8xA2OKSTL+LLdOhq4yXoEIJuBd4UE9tQ79c2
A5cIbs7fXNryA0MK32MYwH2FF8KHAojwxB028qYEwkpDuQXy71RZRAdlNQ/9UDk27GRLmgIQvS86
6Fh9sXaQzt6bhZQetXuHQGNeiMbWQzJsmAVb3HoSYCs7RaJsmQKJVhOnf532LefwlVftNVmSXkVF
WMR1xtM1Rf5FfREFD5agr17aH3bjXLutsz/mVCwrDsBTY5LEc15oSKzy0jdHURh1sRN7UrenEush
aRYOu6px50byJ8TDM51OUr+G5kKHx5rQYxRe1f8Yena2UT545mPz0HwdZKBi5q9wFB0OssJOgS6j
MC6bOt5dw6FpeHJKbBT0lpaKWIPKGYLkAJ9+KFSdQoVXHCe3E6eXwAosBh+vVkFLfET73Io6GNk+
D2nUm/KXuvFJLwz+PFh95xjqsUAfNGz4NW+qyPPubSM40YrF3tiATjcXffjIhqtUUFfQ3b2BEgGD
LAqkZBZhyqC+1QL7jXRlt3TgWNv9FFInd0IzbqwG+1dezmW/ASWQIvZz2VpmQ2FAFUFPUQHrGNxY
1lIlTxYmnuQt2rWbxchdFHGVwofEm5794dy7BUvvRCky1F2dMxmyZKM77Stdd8Uzo6D3Q9OQOaUf
LVGMbTPwZ1Jv7zCcw6CU7p6BVs2gIiejDvLS3mbWLAaSI61qYuoXj00hAxxPGg/qercJMXFJCu3C
D8Zut15/BmiB7ISwX57DiuBHF+Qns6y7XgRWVnrvy3EL5FInFpGIRNDt6DeSWQdZdoLkwjwP9UE4
Qu1hNhYKtb+gK39e1KlkQ6lfc8V4wUY58VjQojtP31EJ6Uzkcz9AksHtTboeh1WAwaA8cdAIzizx
J4eEYxknlyaLW2i9xtVFg8Ta2oMWlBttmdGMM64y5qaUdZeZTh4m1SbwNkQ7LVMQeqUhq2yCydpj
S68vx2OUpYs2gExGznLOvIjA0WZie+3z9JsQ67iehNrkmqeoboFg/pqW9BxzZl/ywKahUNuExhHy
TO0ZfcPjiH05EgJaV0PQTlQMHzaGzKoGdLbBPeeeBkUd5OA7iD4YNzMRapydDOHrfuutlmV06CO7
CbQ6h2ZR2hM8umaomWv7pElH39x8jfTYcib4aP0Dr/RzoJS3VjzZXn4rAdX8bdDhCXsQh9VL5D54
KwfRNJ7YpWbxiqCpbrHhqpq3p3rRZfQsY12GeW8KJjEKRLv6zvhxAdUVzmGGFbuoXd3wmqe75Rcr
Bo5jvmXhQQ501Cv4ulyP0fiv2sLjaE7S1HhopaLfIy4juYn2PWSGx5IuJE6rETzlSoRTZroyulqA
aDYW5Wl1AN5gON7QzDk+RTaw03gE4OZMNlsYIvt08BKJeqjA1FVi13XaxHdlLOP9LVBMwlOBB0oQ
tCQYuKgm7mdb87bVPw15FeAtNIksqn+Li6L+zXJB0MSFqiJx3yojhVS1hxnE+RRC5uinRGjoShJu
leJDq1aVYZvKj7mGhx1ocsv1tjbt0YmbBmxvz+J9oWMDlpL0yeCnMNaiK1rjH0XvDM8N1/8d5emH
+LxAXwuigLCKfF1Bw2K/T1EFpm10cwX/gioJzkh86EooOUGX7xB0ePoOG+23RdEIeBRbFy8+NxaH
o/1HyOTwNNidtvtaiBSR2qhGB9hKv89ELJS/gVqoNgCkisM1amnHBAiPRGhF02jUzZwRVMjsg9ZV
E4kHp/91UDy+Ah2b0L7iDm4NOxA5+hUVkM19TgY+E1s9RR6ERiinnrMJs5z+xDym1gsTqh+IQk3v
A5h6iHML2/+X/xFGtbSdUx6hG7YtJpbQTQIMuwfHHqcaBzRi4+wP5eaeGaKrfxNoRSA+6mJAy8ay
RGbA79X73NtFt9LD9RZhP6QoLckfVDzBh+dBIWONNvT1UqoJhfhfZtkROc6ZtnpRHrUgLLKItV6z
YQTT5xMBZrVgmwIWQua+iWdtyr8Hq46NNjZ56POFs32nBc2rAoYoHSQkOK/y1xgajNd4mK/gu5zf
Ym1j8QFgXbZ8kKxENG0tfZSvmJamNblmg8SRPj180U1cEsupwW6CMbZxUGMQIvgghf95SkQNWZSm
2rIYV1W5wPw8NlxnSaLegvO8D+bEJV3xfqnavihlJhF48MixZCe5MYvW9cLBGmYjCBQVwyW1MX3L
u4iTsHUk4xqv+m6H1qZiSpWS9Exv9FjmjLUDmXzUljt7Zk16g2NuhROURHMhrCreUbsj4sPgYs9M
HfqrF9fCatzeRpPQyjmFHdseyIdT1u8UkbMkubd+bdF025oeT70toQS2pqb7NrlxejSwUvvjkfrs
5Iw9P3pTazB9OFf6oFGNf4PjhfoeJdIy0dUT1WKCrqm42hOTdVM7TtAfmJV4PKdrxvZTyrR0BBrX
Dcx1kRFbquk74rKSsWFh+o7HOaztCww6D5sYwfIggx2zP5+9AiyC8l2iDx3N1pw3bQUy978HL4+C
ATeHy87gI90HMiiAFCjr5Yw7GrZtjIl7m2fw/OqiHaCEWX6Mrk25ZNCDJVyNOzACHTwRkVyfEgoR
qDVxUUOx4R/ehGDEUl/bWhAEqiDjQLVQr0z7tIEhXtE1q10j3XjufStbo41xEU2StjQ5HQ/TXMDe
qeSD2Jc3AjF8Fvc2IF2vDlaOAVwhVZgii1HT26XpgiBHENqjfMtGGw41E/KBsPIreO/+hVmAgHBY
2eatqJRlCcIjXNKhl2kppwiUG6WTO6LsROfteJuCwZm2p4nX1YMMJF0SnAdjQBHJExVmbIBCoUue
Y8Fx69dcV0d1uqsavIbf171i4k/85uf5IbYX0nBWMtWEFatJQArchPFmsX3O9ZhODRJGdR1Zm/Xb
t76c/17xokiTu4XxBG3cGbrBOSYlOSBIbaxcgEX9A1roObctS7EL9Szrpsj50pMgQkNHEn5MbB3q
ntM0X3ifzv68gaeW2XrAmIQ69YqGgnsUll/PS1SrwGoPm/EjUnOM5oR3M8yDmVHon0V2uNMvmEfB
40uFYlHd2f7BMtSxoJcdpVjY4j0dAnotbIO7xDoxxllCsDsy36+GEcf/NxjX+/VUEtA3nu8dlj/A
GZhTZtC1BgS6ew1yJLZqqjePrG97lOh4lk3WjjEzyxa40HuJsxqdL7VKz3rH7PeL2J2eUUq29We9
++50QLLzA5telAIJNzIioW0YFFpupwDzk+z95TWNVbTDJK1cJ9IMoFwv8FmXv8qjGXkXKzkAfVGK
JAdz+JNSaulFbkMAejUJPUcwfMlaUYPpicXFFaHCU5TzkARDbkqA08UEbjUGgNwphexuyzNT1W9z
HAtFf0i0n5X4COOurAwTWGXZBPDJbudkWGC+rFmbk8jCTfUYGm6LRTDiiafzmVYPQJHK1A4GXoge
COorfRH0SQj8oaWmw+nRI18OEmx70+VdyHsLOKHy2wD5WChieN0BqJUkIwXLIdO2h6F5jFV6LQCn
aT6frXij+Gn0lAA0VBMIBOeeAoj50rQjNG+qrr8gUXqNai0IuIanm+jUHOPEHlQsSdgl+JCsWK7Y
YUZsRCcSPVIpIaq53ApQk4Uzft4FlIvpJXZDeOnIDi7tr8bb+hCA0ZHuuad/fFW9igzMjRrQjrfh
T6ajY71f/mw4gYDeJkQeOzhofSmOTVbu0CUK2ImmoCdCATG2HzkOZJpMMOXf9uX2OTnl77zWGb/n
6VSd8ZR3yHm9tEyAASTk43Ot8NUAqUuS/f0PU3rip/WvfdKLBExUHETQQtToY9Ycie/jtISpXzvr
M2u09uQhSCcuWZSmWGWtTbtsShwVHByPXdz68jRMfoPZHvRpzDzltgCtrSwkmZb5OZiABsj8T6+h
36W0NWNIOiCTjYYvLEn2VAUuOlGgb/MmW6x0fBgJj6yjJ4eFvNbMxEdIxmIm4ONqaP3qHgBrO8XX
JaUpVcTISE3gBhsC8vpb4kTgZKTy8ITJBRODU7aMa4DgPxTvBS7lyr28tK2AfUCIzvPY5zHRl/QL
7MEB8U6Kr0JSCT6DptYUGEjcbgI3wue70Sk01w3449jf5HdWzlpqSfMgPjMdz8BRD6BrDqtTCq4b
DfDS4V0fVva9JMw4sVx1RuFS8mAEyEM/8pU8YEa2XAkKKNkCOuJFMwB033djymiS0LJPQT9JIgjY
Rgw7y6cIo09jTKGtgNfGYQ8AlGDQsa2av+V/yP4baKXz4UFFjHNjrc9/TFEEv8Ki/dRrCLMsnC+q
qb53phyHTZxpGuqzF46GU2UEGI8OTW5nGRHQrlgC71uCngupSDAznBRxzbMNDc6ue21xLg+hPZlb
KcQEM7BRwrs1PrzpMN+gM36xZC4pK+DblneRDOQpV5XrOaAbrCd5cxxoQvPrKITSz8EH7XFVCvpj
PPjrnfbrxuVV1koWXSAd8ScapjhY8PX/0kYwCXu426o1Iix9vD2vEdDKpgDdsl18G1X4NFEGgcxs
/fTgsbezLEmqr4UwKs6dOeL4D1I0fM1DY5P/SpyPBUFgBohkuHTyIqHJ4agFMoMXMVLovamenl4T
71NJ49C0qdwniMcXTqEU0PdCWXq9hnqMm16GOPS3teZGUeGzBs/gD6lFhueF59y6I09eFPuBH+AC
gLo8UwNWmH1BFZphjJfO28jrmZo7tzrdBxcwvDO0JsFoh9yCAOihA5GrapXruwozPY3Zca30v94I
D79+bGcS5W/DXch33T25V2PJW3RwgRe2jAvSEICynrWu2EuBkUPncG5r1zBWQaNCVmofCq5dqwa1
VCK/PKYzcg9UZhSDEY5VHNvFNqZn3QjUCnT7rj8E8kr4TbXuuko/24+yVSdJGik+d1FcrX9BNAZs
ZppwZAe3+ZAGIKY3+HfjTE/4qV2F0Sh+nZm58O3F4zXrSqCivVjhwAMzbE9FTa3aWzkKw2SR87pP
3N11CsfVrAkgULro8m3BmqFr85ESFbudDG5UBhOSdb3vHviJK8z9tGYnUY2homTdEXvKsAOfMv0G
b3hQg4vP2hcWNlVkGxCQfox+DiOM8SnFmiU9Si0p7EYao4bLH//vk/yVJa5yc30j8s0+rHPVj4Wz
xILBRrgI4mlF/+z5Q8hhEOPIY8bpnVvmVeDkHtj73ZklBUG5LlsPh1O6vsTgeVUiJsqHrdWCdmH1
G9xKrVUIOdke/RUGGlUgiaiCbNMoY11K6MgFHmRt9U5zro1aReA4lT8cAHw/NLNTBoHoP5d4oEr3
wshbUMrY+B7TIMNtyYrxMD2ZuGhUCCuZWuXzLvuEvUtpzN13cT0diNf9UETxMWZa3r3tHFJ+nuKe
FlFFlJqQdiYZg9tFmLzfo3E2KihtIKeQtsN08fUwNUOq00gLHgXdZDrfWj5XzlFRywmqL85UgXUy
q32l7VJwFqQOjm2+xYpMzA6da1On5wvBDZNzxDz+LZgwuGA4Zy3A7AdzQ5UxKBMrkp9M9AkZpAnh
upFnjcS/+ePNyDAykdBx+i0E0CtdRJEPKVjeBtfU3dlIlvHuDLZt4V90aVojWFdYL64IDQNMaWwW
fwn/rvDMnxeP4sI6yND8QLBZUOUDuJspTYOXu1e7KnQOEGUFy16wnS+BqMcGZqFkuhXwRwwrqIWg
29lyZcvbA0CY2wABwmtIksEdTuwJWh544cwS3ByJxLEonufdkSCkTD4O9NXonzLWoiNY3BYoEVCU
n6L0mlXzQG1iHBowFbNMrwD9ywg0MHnY+68w4eS3CRBF5uBsZNRIUvUc3YHXi9O795OndqYhtWti
akU8+fryPwNkgG4wNYu8zytAtEIEBictsNrxa9tXHDmdsNYPa5gipkHQeo+Af57xJ+4GQ877LJTC
MmNUm0OhVXLh4UY7oAelP5hpFmhlWdE4/9Ehpdxh/Ha/AzuSEdYS0SYbucazD8i32bBfSpX427UP
5Ll1yJFzR7PBqit9D0RyrpsYa5KI1moVvMpRz91IQm3XV8aNb59i7i08pbj61jLjJNnYPyXXuApf
S25l21QPgKxA7pHiRbPtIeIGJ9TiRMBYY4rJH3H/Xh0+DUJTF7TiOO0Fd3rPaoGp5hKgU213B9Qk
gF5t9W9eEdEfZSbsypy3IT7zavpTVcY5TfsXRD2jFIHJjXrN3s3LKQBC27IonsVig6Sf0sT8tfa/
+g2MGoi7LXZa4J+19fs0wULQnEOfiNyOETD9kbcpKf6zZ8dD+BtrF3xVU4I885J5QTJ67pJ9PtyB
rUnsy4rsk73k/ydpQn6deywWl4e6lZ8P4qv0HtHUyiUVrgjZ7A40QdSq4TwkRBudBMsxur2iz9AX
HcKLBosk354zj+YjAjN2Xfi/G6bPPbL2AhpU15hVyz6bp/MiniEooqcw0/dv4gw9VAzOOVwh7/NI
plVKYN5VD7iOlSlj+/pUUEQNdXnt1maCG71dBQAqx9oQymklKgZ4QB3Ub+PzOkO4ehwviVQLjHBd
n+nQRlEIr1uWtEIBPjnjqogN9h+9ugeMC2Dh9ZRQCb9qK9lDB2tImTNTycX2uhRjz2bXe2EDNYY9
h/LpxxFdioLtO0kG30IxTZtBjdgrtFXu33PanHoUzKQs8h5sTsi4AmiKHR5mhdMTLtGOqHa/YMDx
IuXMdecRjVcSRSZQuSdLuOY1x/2lvdjZ/tSVp9Wp5csfA3dcKYYhsDPmDDsmf6HmcQf+0H4TFTHL
/buikpwXSdf4GfOrm8+mh562lri8x5XH+7GAD1DlIYnWpiCg0uav+HbwH/BHRjVZICMh0u9Df4l5
F4KE4sRDTwkBY85vt8J7g7PfAzc5giUDi932w7oa7YEo8HJxnrYODdlViMS+1Witq1Uuopg1sjUg
6DSwTstRZzMGB945p2VHW4aQYhuYF1XzsbobO3J8Cdpatd29O0KeTkLzc1X2JZ2vBqwuCjBrBJoA
vHkBnh4yfaPSde++0w9fYr2oJe3iNnXKR+9BwNBLirn61ty2eVNGGKAkuOsOWh9c4rP+PC9NeXnN
HyfyhyeQCui05WZswFcd9gJeQMdJqaxDdQaNgaS05GojJf0iEtONVQiVXfznjDqCxumTDI6JoznH
FF26vKe7pmQNiAVn2xaVzAQ4sQhWgI84rpldbwt9axI2lpJJibV3B5EXuosNVx+mNjh131jF6Okl
K1EvR8Av8/Q4RYZ/nq7gg2eykYwQbsrycrFQ6bi2bb0woAy7xlpRIHMvoGXADg7WnhVSyiRSeaVE
QE6aZ/EQD675sMjmIwMFu6Brl2fT9JTRbKS4RXD7joC+dFmlU3+X8e878IYvbX5k+3e3U5uDAt6I
wSw9rWCQvdFheNoTJEOt8bI6YcSefwWLJg1KyNx/k5RF0p8k50yn6l+JTSH1ROVvNLh5esXSSkNA
0rT3EVieykjwHQOi012h1PiYPyd+cj3wxa4okct+OuSQecGTs4G/orA8iaGSUmUrD/QWK+yFLuRG
t6C/5PKj7UxeQ+ltGPP3Vcc7anz0HQ4VePe9ea3JErJ/Ssit3/ErJ9Bll4zMkDbW+iEhPUsKU5Ed
lHccjoNWzuK9qU+yOCEc08fwkbUkN1S6uHooL71n44Qd6dH1b+Rdn+n3sODgM+ClroJQ6LEuE3kJ
Fj/+VjCcDy0PT5FfaA/XA3fkojXiH91NeVqeQnxFYFXg1jRor6tHDC8mVGlfNw1Y98Pv18QJh/HK
0Ub50r+7eliMt0Ws/L0lj3fwAL6rrrpIfoCQ2be6xW1RAMn/AOYCaZoWbgCq4AoG5XpvL2wYGXoy
nR7whdvPg3ZKK6BD9mRQXZndUwnL05nrsVySL1R8alTW/MldOgvSAnXreVvOajVj99IuXTgQ3JdM
1LTj43+EQ9ENoJ8PflEVLV7tuPRYruetnhMGADwzJziKw0Hn2IlZCnk1llzEd5VW12GqTwCIxO9G
z88FrWTnUPjGfJguwzWplNxZ0eRKaWJxvlwASE+dg1r5eEUnDUqNELpnXIYr9GE/1NCNXHGAGpB+
I5UXEFCjGb/n+JkoLXEFO/CZeKODbhRnaIZ185StKt2xZ97V+l5dlDI/ewFmoj7WHGkboSIux/Q6
uBIYjgDBAm+Xw8E8vuK/6QDlK6yVDA9dzSvc2zyusy/IwaDpZWyJFGPDbqFDDrRqQbYcBxqZPO1w
2opHq04qHYkp7txco8gCW8B2yFbJEjvi9VTEUfMKYH5WEJoHccRXtWJw7orTRNM0GZCvQAyUh1mo
/R11+CcxSHwN6BMzYvPFCWzZkW0FmVibtVHOb6twCGLwymjXTaY7aR3CxebRdpesuTngayAxjwIW
MK0RB+/KdJ1sql21uI8PL3VARCIn/Yyj1ErWpCbvbPOEbASd5IWV6H3Su4i5+Ir4uXWkGYTwamol
iJtE3kHZBBtn9VV5X8vdW2G+OrwmCyUKy35WAL/UelWYjggqjhZDnQi7GSOR+kciKtR3XOZIq9dt
srdZgtnKF4Kx4zN7kiqUY9dLFsSNkfv7fKMd97rJssj+xdZyw4LBkZlZblwYijO+O+s36aVh0YKD
venNACqZuJzjgrFsh6y39sznm2XRduqW/hQ29zjxR/pX5YtfN/bYRvmZqRcIbZDpV9e7qVGnhxY+
LaBeuCu1Vbl+78inBB5MKVkbZDV4f0i2di72UzEjPzN/eE0T8THBjMTzLVvx8tdqJSzvXcn0DT+O
n7hKBeEPh8rNwoq4vJYjGPrKs8vv/k/pYE0Zlg247at/Fwcnhzxc0kvKejPco7IZaTtGngy4rGZE
g3h0XV31Okqz1MMNLk6rKLYh2NhP/zmAhi4K5OW+Lfn+QHU6eRgbvWvjVa4g2uTDDVQVf1WHymmw
L9+QzrxmaZWnesZ1/VLdO0ApeifK3A7eb2RrnezWe//lH61HoH+gW9S+hUaMFQL3yejsv/aMHNxR
BK40O0b60hYVKetG7OgHrrQHuVSnaCQDnTlGzOe1HFFO6T4ihyJPeZGqudtw2nQh4DM0evuv+B40
aW4CoNRY2W8qzn0ceRQvpMXaP6eQZekhA3fcF91LNApn19KM+9UDDKhNZleX+I7RLEMDuCzoG41Y
29RhH/JleuLvpCUfyOfktYO+FwaYOlX6aNTtp0OFwguVnTuyky/frHvMvOUggSYFdgyVvC2fY3lr
TUBaC9YExn+WDf9BvoQlyeKyUHMDetLEi2sxZCxs+ZRl5xt20SIXbMNLFGP67m35Cv0ghM8Y+xMp
rV8FRcqsCUTnL0IcjaHZ5EVcECT3+48IpP7rAUd5YxpAoAGhq6fIwMkGwW1U5HqvOeubsVXn6jXg
KAEYWbn5GH3tnypvKDXLxRudTj371wWWmpi3RbaWmMTKQYhdTmiIv8rUcPW4UdjrEe9A5YGav534
JbnOSanFrCfixT9QS+5BfpRRl/ZRXKtwbxu1yJux+qceypM/isTCYHvDB+Zm9Ke9Y5uMq1rV8pZD
qu4exNIAdOVpmng5PVI6VXgV7FG21tWeNMDACAghe1u/PTFVVutL8q0vLPD1MlHniMkWxE98WsjX
tGwV14YBxIDzHlnDPWJ0ZcJ0ceEcbJRueBRY5VXwsfgmVIgk3IP0yOwJcF2RpDJMzRq2Uv3RxraB
iCoRVx31QoWUQ2ypMHaM+vTiddbe/Dob+LeeZ9FSZw5lRbWWf/L6T/4di+ZTN8Fuq6TOlnRkTeDh
kfERVUjEsozbt05rY69TOHBZDvcJ24OIVMSuSlgeOuQPsVQ31UUL6NbuhWssZZbson1WWaWVFPRj
7py7DqSUgE88SVmReEW424gpdFnNupm60DQH5DW/fNRCylygwl1QWn+oM0+mIFYNJ357gLNy+1OZ
4vWqs5t8YR8xZKdL6RdCPLjal2pJ9NjOyG8RDxcttW87DKpViimQy48sIMGVHpgj5WTH1nvowmXS
sxpWTKhrO7/9P7Y54FsFysKigR5K0DhbrPzDlZc2wFM1OuauzEm4rbNswB1kY+zbmT53P2ZloZRz
EBiVcmZGakn0YD1QxFyUsopywxPl5NzWn9Oc/q6dSrdIe723i/4ApO2x/S6AcPQxvGXy9XXkiaqy
uBDDJZ+sydAJWNwSVlveXYqtfGYvHUrbXhVTvEHmfI9x8636U0tLVDsYJKq2StvuqeRl7OjYeoha
Cp0/TdleQw/w6KZOd7mdB6PpiuQP6Zt903gBhfyh4GtovB61yybNiI9XjhZWd+mYJxGXUpsfWezr
kiAtXMUMkjWoDCFXMOLX1nVpA+YI2EcpJWHt/iqCjMkBLL+HOh7EubFtb5cvBNAtrrucf70Yo/Cb
ZxQu3MvYHjIdrXSDuWKZHSmg3XxXV5MDnt2VZGNN9Tqw4g1sfffVlRmdL6jHR5aj5N6aeOJ9lz14
ab6TuiAfGXJo35oZeWZs/VaUgddgv0NLkDP3M5jh6iM2kvzO7XndWlyaaIoDqIEjmMqy4WQ32W6p
SvjHEapvM4GWE8IG46tBH/lfvFlBY9IlARd/kHlUH+bl6ihWyjJKkIIrgfmv8+uHv31kj/MHy6dG
0tSTtUp7V94uAE2p6Zpz/liUgtPLwSfHDPVKYgP6kp84nwoV4TxnvD992yQkKGIc5c+OvmmIzmVA
pNu+/2SbPJT0GFuP6HcoBatAHDMpq8KgVSS6njbU2ThtRw5bS3KQyy1GKAOH+WodtxpaBKTF4Glx
la1rA6v8jQgdombhPo+0igJApTa+K3Z9zh9Nhec2MbNvoLQMRUOdFQ/Ya6x2TgIJMZbXj5PpKIHy
PM7rEm7wVZ/kAp6n0SM25V0VVv8aMEYtwIndew9NSu1WfBRoEGsRQJMHCDmf0SeQ8UO0jIO9yOh9
+So4Tt78s93aP49hKL8d5h6RbCrN4XPbvJwmSQ9dOtX201FD8YCjaiGcxGkw5gJpleAf4Q0KjEtd
Z1Fa3SLAT9ubkX4bnLM8/yZj0NiBtcBvKBrRdIL8PcZbRUW+sFEIemLnAjmRe6iT1mLoH22wCB6X
VoIF6eX/D0f63XwGiaz03JyfMQQUIcy1JexFsh5rZBD4/dd3NdsO3Bja5EZhIo7jGqW1O+jZIIXm
kVhSpROkXyRgcUwUfCsPgTS6CRacZXQ51ecJCUQJaX7Rft1m2CYu4t1KlGEmmRutMLsWTtb0DMId
jAlOCfSZjs330xKiDtkoHf/wX29SHUAr3trYXQ9HExGRpxJGnExE0oXA1GVBaqsRnxIUYFKLnM3+
+Kprk+1yN0gV5EcA1nKaM08qCdO02RY/e/HZQfIRRc7Oc0D6WlFPKyttiTf4ZSfOjJVq+gt0Rrp8
Tqlk9HynHLB+JHkM8JSFMAnO6G+uu1ur2lXOyj+czWywefOukjc3aaSLTjSPLkBXrPHsmG0x/dln
O8HAljzL6dH685/mkuGlpjhdljo+2g7IjY464Uy2+EgKGssC5FyGMzh2h4PA2ZhviZCikSF5/HE4
gaqROGaovaG149ZZEvGF9Gzlhcw0V14cmwHvSJcd/+eDX1jR5Y9bzy+Bb1UoIz4edVgY8XlEQfcg
zyOIr7XgwZ22jqyQOuO21CfPsJ9XeE6fk0CZwd9wCi+EJ2PtT32iPCou6WcwBDXys19UlozK5cFh
8widfmwYHwNClKj/gCfT4SyV+mGVEIuQlm3dQVCXfObB7WbOLCUJ2HJIwqQo+0V7x4gfh2FZ9ges
Oz0IRGwF9SXbAQ2ersB1UumHkQxZof9HXhS7UiNZciMFMRJ0JDp+kIx0WQfnwa0yAjcGzePLRi6+
eFAI3Ja4a4SuiGFRxEeYSCrLqlcbpQgM139osSoTG2gwU8w76TxGNkztwM5U2/sHi827J463ce10
/TYl2DLmDgn07KHNqTyWfZIqwWLFXW/nbaByg+bS5gu28LTd7mO0N3wTN1uyLhZRu5DVRLv2zq5x
4M84dAlqDIXRjAYdPt357CLnGNGIPWo1X0Uy4su+m8MIxjyzKlB52GOpPurRIBAbjKrBelQttDoc
m5VJ6mButIoANfEQ61w1QAz2sSyC+5C6Wv65V3SWeTox+/OFcWbjjuvp9taEr9Pakp8rS9E98b73
BVaJuviJCtgBxyMMWDLmA6loZloDbJ9PgHbL/BWxsSL3a1t8RDVC8AuAu1amWezvw0x+h8IyL9do
C7DAfpC5sjblhV6KNngQ6wBlGvtq1aCcqSh7cexlxVE0suDCsd3ArCwYMA9w4OyZt38/YPsi+1G7
xSnk669EwBx3LOgEcpTcv96bg8JqPKP0N0LQanoQLmTBM0OfXjnpsf2pyvPUeRhX+fiZqHFkMoFU
rj4WVtHChaqD1s+Zp1zonSqrpHgQyirzHkDKrB+E9uIwMaVmBK81A9AIe4FFosJTAFsqsQGFaPI2
/ZDmIbPriAx64GKuw945mkIrtVKWEJLYbpvEXJb4rtYrpVQoXoapcCnVvGD/lN/2K/cUawW6ZA1A
JiA+j8nhK+XFNSdeKzEiHPZ7B7uflgkwHnKGWjJM9YAu/NeIL5JeZbaZBGBQhrhuMu5OR1NCLtDx
qQvByGIY5JaohQo2AM1thjj2rlRf1A2hDk69wtLhyAywzlg3P9cSblfCko63gMyO4pehwFhLm54E
g4Xp/1oljVDt25g17I3jkpSM+iH4uwvy6slz8l4kRpKjHePGr8REmcUBzqwJTvoKeIT22fn/9FuQ
uBBD5C7qPQbWbkDHh+6y58NUBQBLIVQalYI6lW3ggGSMNd9N7wQbl6VYBSG3dR8cJqOf0NNFmc7Z
QOsXY9eazS7xzxLe4o/9QXG4ouhV1kysO00xqSb0kXXZ59ZZflfD+9zEAt18iLt2Vw/J1WSqWKU9
sew07Yt6eYELHRJeD4AjC7StLjbDGF4u/+AIBIxpBxiSfR2ABc9LvNTJwOzFlkapeLHIrgs9ujT2
C0GrDWmhuvrZ/5XBmYy4LJM9HRyjNuI5T6uAYRrpYRYaWT9uZK8eT9qcTASmukLiQiLAlQsjP3sr
DWh+4tcOkqNaqf65pMo4hQwV1noA/kk0/JMgPsmmrqIVzysv7/rOMA3EIGSYiK8GzEC5ZgkRRtrC
K+afaemlBZJQi90110tya8y9U3okUOY5/nwJ/zTYvkSTR93OwrmEfsG/t8mnRiQUME5rT29IwIbB
PBNttdAXKDNsGkK2lneZZLf/9NkKawTq/0Jygc3QTAxsKjz3Rg0XyGH1DautTimkOl/eyXDuKlRa
Dr/Y1wCo8Dmq2lEMC8ZB9T+s3/yqTPDO8sAF5VcWvoiHhESUE1azhRw1IuWpVyydic21dj2GC0RW
gm7O4doku4/6s9/LbKwbfpuWjwJo729gHlQG1BPZoykyuwawT9/9gSvSVyKZtdy1YAW2zMMRB+di
I810uRfoqwq2YLGb7NaLNrQTcYi5aNBPirDl08sUdnBNfQSVZCue4RSRMzmKKW/QpS6+9NGAfFeE
NT4w1172/8IuZ/3G6KPrpRsXueDeAuIMu08ktwzTIwl98YPkCx0fjyo4uMoybkekY8Tt1eiygWMp
DAG4LU1MV8fenZImCKR3LWsVF7wkgeE9X1wJcf2naXoly/lKOcrVxMx9BENkZepfYvDvRW25ye2O
aw0r/D7/as6zAkbP2Qq1IFlOh43MQnIJH/o7fT1qqax2zrvVdjz/4wx7mtXa4GQdy/8jUVKse0K0
lelBrPGTMOppPOUg5VcNrwEr2JqzwpVUs5UbXZnqxPzKmtz+3xbe70za9p85V9G+Qg4iPkdK9X+P
DLQIgMBPOVHue8WOQtyJtZ3QZBcESMWvkshPoUmfEvU5GrguupRK6MwK4ZKS4wXZrZrULseK29Cs
0EpZMAvILlhQ4JMgH8Tg86audiWxMSN6nl9F3f4965RUbRRW3yjuRNyxE/W5Q3qbOPwhy3xYLFiK
f2/yKZO3MoKUAm9T48zOFdJPw/SY3GVclgotchdRINVQKXE0AyQXgRTandqzFVWQGARd8ifUytdV
JgILTLKnNSFJ0gY5Y9PWCzHr009+yIqxqQh07QKODpJRpx5jkhZ+buLxdjfG0k1WctU+SEA8yhLV
tl/HmTAnJ4nybcf1MeRpRtAYES9Morp5qD2TFSkIrbXkOBmDkokSaa+v1kGZzYalq5rdpne3DAYF
rrisKpTl85iF4/vdYAr84i1ufkDg0BfaCU/ghXefpfa9VOLzE8wDyEJXt/ppfT1iCNPD8kkJ4YYJ
uISP2+YK0VmA49wGpO5qPm5+lJw0pyDWjCHTET/TXdxZK23VqsRPLuril4tWbB4TpD8c/eJi9B8e
TXtu3oBzo9PrUXDnsVk9nonOVTZqkH2LVksLhwiiKqcGYDbeBaiLlZ49K0Sr355A/UQQ0fgzHU/Y
vYDRfjLEm0bJuVmsoQwZ3RZhFFBIhiFUSOcoFeJsvy42BHnXEUXcVZPyeNOy1mCScU5eazz14U2p
08X9FwWOOqBTXQbYnPpO8VVFKLXsM/dM6mNG1svRMQikFnbvi3NFuDVjitf7isudPYXf+dviLC0h
MP37j3jsBDedMTbA5FayM9OPk69VX3M1K6xHTq5EdP100JN9Rwhaxj6p/AUrybyX+zl/Og8dwZ5T
a9UWhUvYp7QUo9kXBkxe6Cc6Mt/0Y3/Sif81oA5l9ekB9UC03aJ+a4yb6kmmZS6+eCar7HNAWV7q
60gxCv+a7h0rBHvP0boiLi1FcAsAjbB3esC7xAkc7WfN8wBGXIKYlf0R5+Wm8TWy//0upnj1KN4f
b0IqRoHeo3jzt17GPLoBcrQHa2XHu6mwmayglQJppyegtJCTTV0BhlgH7PVpiSzSX949lzvHWQ8A
CGjEG0VByC5vc6G7LlWM2YFfgLtJo6zDzpcAmYO0wfOJC3D0DC0APFDBjvD36A8z/uqC76giF4rq
v6eqFd9ys6iTeM4KaLCy6Guf6UDXGTUyGK/VlvC1F6RVgGxC8L2r5fEHqL0V8rO4Dm1O8+pTWkTj
d7d76RLfeOsJ4gVdsJ4Ouy/5vrdlvPKVoGK1d22PjwUNgPkWa93rc64p6tUHkinO1FNov+tbflHd
U+DtbNYNAvcknkClMDA3vb+V1VReWQdQgv64BD0/29caNYnXZ0VY9tq2xmKBcdTROdViOXCFzDG6
wP9VgKi3WxL+F2pt3KAJPkIKIWLbYXDIc6r0w16Vkyvuu23VaCOWe6CrybKahLEFyiFj3Ox1jYEz
z3ZeLygyqmwUuZ7IZOpSjlTWKNnKMcnsEYSBsRE8UeOiBfyLi9hs8qZwhRkdmk9HkAiun2c4GzT2
93fG1sgNO2a8aBqaLHcDz2PKM5+R7KNF+25hP92wtPv4VwqMMPXGZRX/MARq+vv7qp/ftjgwUU7k
atySMOutlZFTC57rv27Hk2KGOnvvLLOUks6Y38JOPXCEKVrKzrpFrtKJHA9aq7csXog2wtp4+WnX
xgslEVHe7WluiPmAnGOZi+uJ7IWfEztzaeWbNlpJErXA0QAWsHsCUWHJVa2KjpO4VnRzJAeYrzG+
mnX6a1X8LaYZSpcm64N0DP7lYkD0/iydKeA2i3P9CT+jVbAHUlEVOG0Ut4xO2HaTNb+ZsaCZPLnA
Ke0MvOyb1buI71qFddolrGVcCaa5V8mW8pRlpPxeDh0L3GoJ8MZbF6kPSddyEotzhHKT9x2a8ka3
jChn1uyQybL3tdl441rnLvwCmewwCUpdUueNU+R7Ia3x1BtdYRKVe/ywZVyu8TtUBwfSk1mLgB6B
Hbr1RKqVN5W7iMcyujkC7CC5L3VwSaWnZI2HLUyYy51rBq92g6ToJlnI0dDy1u4PdFKrGGpetePx
3Jpo3NJgWqnEiWkw87IiSJ9pYmydJFzmGtzKXN+e+mD/Wm71vAEhdyD2fHHJkVV08ulBU+QZFDAc
r+zVipjYc2YytW2DwkVg8gyAsd51fcF4PGl0sCUYUV77UOgDv87TkzBQNh3Ed4KlsVgiQwD8fkCF
VNfAilfk6KsGbT9eBVFtDCv0LiCun8TDkMODqdId16VjmH7145I1rQ9Dg5TCEnjLLWc+yR5XsM+x
879cXAfjApJ5lj6Za5ZoCwln/F2us33uKmYH/OE+FUZ+xBoNHCM4V+cZORaSoGN7r20mKq1owV0M
gSyNjPMHJJDbePXA6pXv3mLUPse4bGPuV8TOxk+GZjDfLQi1Nd00CXEs4bwDA/yG6HsOwvcMya7i
eho6e5JM7HSkbD8VdvHNsvOf2miyRh6hgIX3Buw6YXXOiqTlylk0Z5SsYTMkej3CEoAtLtFWWkHa
n9OhuaiE1l1fQz69U53Q40Wc40+Atet6DJoI5Wbh7cVctw7u313jmKfYBEdTHHJybLLFj9FSwCmr
syM2DYBOMIoesrhQ6wPeOuchKJ3xZCXIHD9caKTRd+NGDClWBHX+9cxw/NvZ6KAaEdFu4Q21FFPN
R2tGJmNyPiCwr6rBn1SLgr+9b95hnOTeL7qrTTyH8kNDJRG7G9RXkmGyYBlQXSDhASQMhaZrxEEF
SnF3qIeUp5gVujVXRcAg2GXZT08W7jSAzsZFKF06MgMlvmETodiHwJO2M4Ne9EXpD5k5oCXK7i50
WHbo+Xjf+kgS+pTT45007iVyFeKtyZqZKBnzEUbHqxjliZT9W747KCe4OdQWY6iMVQvGsmgRUiiq
OeKvn6KEbprcdRVlg2Eid0JAZZwnnOX68gkzwrZG+fPUwoNIgHlTKxfD8wmQk0rYq3kydMeS0Fat
hSNAuQpczwDWZ7iUxIbR4zhg20dgnqkpRY/7ZxbTQxTaoBlDxlwl7bH944IzXyQNIJNUPvBUPLXW
SAuK2PNd3GKvCsJGGL77nGsAXulampxipU8TMlOKkctScMT14LrAIHSDn3UfG6fsQOd6KyhKlA2z
K2FmBuAoLdvO7GodEFWg+H3MTAacaVMnY1eKg2dnrjwbS1wT/hSaVMxpEgei7oUMyXnljeWt7iE8
OGSr7nxrGqWDCnSFimVvO0w7zAv5OQDKOh35KUHNc11ZFLy5cSB+DUOfwXelakzELsFoy0dIwCYa
dHjtI1ozI37j/O/7gGWbtEqVnQwLefaXkJDiIm7vgXruvoE1k4ZTlVGYzvZ6DKQpAG5x3iSDenOm
hwq5TrTEQJbEqL0ujS/bttftZFS16e2qAl8SU2r1LLyrtuCGARTm5e/3ldCf4iyhfNRj5OPU37m8
GhMUtWUBwmFDzD1NfVUwnnLQn1gpXlFlgZ+IO+gR+k2IgWAUF9rq5i3JZzHA4bRZLkV5XquckaWg
GLHt+nd9WvdYfcWaZI+D2M2DGfh+7IYXhpUdO5RwRMrkzunBbY8qKRBuVtmwfVJQTkvtT7h8zql4
wNezB/tl3TbuTtfviGU9+VkILRPgfKWxJ7WcNpLXPSoOuaxWtNpcRxJBqAHjbVZsfGxFUBkU/B16
xOSbMVREBbBDBP3SSiZn3WSAn7UxKkJ1ZCgV0VXF0ZPWdtdslSRti9amjD8Lds+boRAyCDdVi9Hk
MhjbKGvkanJtDoP8b5EImZ5ML+liC/+/4Q0kTUPmkNvjEQR2t3moTvlor+yKMbB1QQ0waJT3dusL
5LjMppYg43S2pD1+kMoguWhVoQmXuRzuy+tUhDqv95TPc0i1yVSvMbgXYgH8oyOwlTscaJpu6Z8L
VK08hxx2RZJbWwsUuCavDqhTvJ27slCdEQn9YltdLro+63lQ8Lneh/zZzjlmOy/66KsqBDRP58Vi
TZsmDTNGKj71NqgpmHOaCM2qe/7oKC3h/hW9InLz7hGhd1ZyW6XbNs/35rYd5Rs2U4BN5swyIgkA
sq7+qmboZ11I+YUsnskbAY/BzOGN47rAOn3BnWfKzmjxDt8MLmO4ZYXNHwSaaZJR4jUdYKnptTJY
hDShAEJ2g/a1wHVMl8IMbdDYfNm2+RXH1RS19ef7e1uU+dI/DFAnAq8S7FGkfEvxqx64OJzBVba6
wXUxEHaA8YluiQrepKdcHTbdtdWeb4hYWf2kVvqz1HrujJrN+5aAa1b8P5nE1OTW9hwCVjU/5r2h
H1I17Iqy7z7ysSFaytt8B3HhRZyjECrOKg2udoJBjFQYcuFwn7lo1qagKyi6l+aGiX3fBlYzzA80
FkuuMZXJpaPbOQamXRxY7oBKIxWcAHN0ZKqlAwoTe1/kECbKSmgvGsdqV+OGukfsWMbv6cwIEB5R
ZgsQjaQxFzuZJ94YprTpo/2M3mxiJvVR6h01RabSFJ5Kul6C9NEiVnb9ht45nqwplSseflPwX6ge
KT+ly1/JbwjIgj+AKIWWjrZlR5nUVah3mG6R2V6ZHB/I57nOU+/Hba5m7adBVg3JGsyH1KCCx78U
ZlthGJz7eFtOYcWU+OKFwPe/4U1t+fVSSMTXsky+iMeMnssuvTBD5RjQX6m61Q91ufQm0esczJrE
nE3XC578sl39hNPj2Q/XwR0q+qAREQFvka0s4CRSs7x2GVnAQhMjpbrp2Yq+4PjAp44+lpNHmoy2
IjxdZ7X3DhlSX9uzamWuCrPVEs+33RtG/izIqisx61i6Wh4Xy7na7wdQPz6Xaq1/mIq0qRBVYQcx
FXzZerPkbUwMZVSLPPQ/bUb6SS7fGLG7H7L03wKCqM7jLSXQy6G6Vg63lCrZWroMDTdal9FyfKDH
qAC+dFmNk4EpJzj17e5dwjSJ7wfZbdLVVsSheSH613HmZUcvGctiKG0ORxST2gHzv0lF0Zd9+wUY
YdxMgsZNFEdzhlkGB7HKinfm1t5kfmp1mKVSQcNJqUnpWA0CAqV9cgSsBHYHfAFS0MWPkJSlw7+v
D5eKL2N9F5Qw403OkxKgqwZd2MFyWAjLGnWIW0MOSURjWC0sFqMGHSFxJ1QnC2VJUln3dKBZ4EZe
y1H/ozgQ/iZjIQORfZSqlrL4Z0Je0q0lJRoMGc8Sq6QRWepbzmpK9OdukVpKUACj5250uIcBlW7o
gVlPi9amvGUjNyIvQrjarxkqGjmH7mOiEwt7fHJ5JbAapu1s6dUDiiZHKTLBpkbhoU1ajA0xu83U
c1Md43Ccmt/uMnXaB2q21POLYnp9BYMO9cETUUjUbgX9Fe4jtPEeWe0OIO5sWwU0Udp/LVoWh4Vq
hwz1VyhPv687BqZ6RDp0PKyKpugqRSeloGmpngFeZgzYMJf06XLyb8N+q5So2hG1dZml+OyFyqV5
2I0p0NJ36bmWzkZaie/IEZu58GLgUr0jwJ1EJB+tpPWPYO68Mj9jPbRDCtVKbdyXb0i1KXd2tYZT
gF9HtUfV/Il0d8Q10FcUKmiSHqgBeiaHjzw3zGy6qOaBsVVisv6VjzQonxLaE5j8VJBZZYodi77l
xRaBJwbBpyJ8lb2wNBRa8L/Y/F/z4HPYfNAH9GMgH+oIlNH772YkQtlLPvJatb8yeKLdy+IaBTh5
8Gg+rPlMf/dG+iovNKzIFzl68LtvOyAS+ttaTCUn0kmZRh8QbsQaxIaMQiuvAosw0WmuTusfX1bX
Tyqt5OM09FgcY3DXSZyM6PhWSxR39c93A4RIPdQpM0fiFineeLMMR0UklXriLmya65NAmIHqNZea
uQ2idxngaSods0SypRMxDFRyFkjr6gWfxRXFlni47VQZGI/Bq1PewA75QVMpcfjmcd/vyjx15A8R
KpsLsjYp5iEgHQ8AX0VvN+x0l2a28eMRoTXDL4rpavz/5ZqyKocHtdLVqPnadRrj/2cIbRIC0rfB
zHnaTjwVcRxBoMncBiv85kbLsy2o9ew/ULlmjRsGUJQcGgpAOYdt0Xhj7J2oxiSuUJX1qP5sTzo0
Q/CtKg+comF9vw4vLLwEubsGCNXBDaIQoBsLhgmH+pGSp2ltcYQLcDJUBdptP+IzZIC5y1nPudlT
Ynpkm6/3iwK8WoyTeTw2cmeIArZfVMLSiIhWLL8Rm18t/PWP3qAClBKMZB+12VqJLL1XT4DSJZ9M
mp3DlnJwKIBg5JiqnYikk66xC2L6UGGOIXM3nomZXz8QKdYQelDZH62HFPQJECRpkQpqYjFTNFaO
6KQB+cUToHBkFkmjrkqH6u245Zq91crORw4+IAuapTJgXJA73vv6B1i1ZYE3vt3vtXJNKWiEGlAH
9UC5lwh09vyU2dzBvZlVcnh+QaXkUG7CT8o2XLMDFDkHm79oiAHQBpKFyaiRAlbOb+6K9ETInSGc
0pscjlG1O6XeQV1qkTgdPIDvEcaSPFtLKTYk7zBN5B9CahWo0Nf8zHpwR8xKDM82ia/NpsqMdz8P
GYP4o2bBUYEFqt/kQ57unAkdss2eVdE9VoZznkJTyOi92dAiIdVG8nJbYjSBy0MgJ3bybHwfWcCj
a8s2iSZcipuVNaJuZJ4btA+d2feBQRsfdVU4b/hVLr49n82GLK0jzg4gDMgLP4rDyd+C2mvrzIyl
ubRlt4kgqFGD9JsTXKbRoeP9aw4WHs750APdSTXDlbfK4/ykeUvwXvHaiz/0CS7FZjniEKWWLrrN
dEOY7iUj9q9ty5TTy8YgHlHwQwh3zzROKtwOi4bbgyqE+YmBqnF0wn+JsPzUMi6iOubuihG/psTg
ibNHdREVKqpRJxGZ5hSg/BmnPkEG8Wwmu1QqvgD3ZVr01DkgmJxcNvgBZ58cvbiSevHpeP78Cx1h
eQKBAcaIcVJceFv/FQygc9+SJquuYYbz2NHYJwNHuKrgPNZuYHs5wqHcd0W1zDgBs+A+2xA5bo1A
iXLDCzrcsd9qpDOpn1Y6x+y3fiPxGXmdGvuz7Yi6YB1C1973OgvH4egMUgZex8dmTF0MSbs1UmfE
JZqtUBQTMdKTDTyQvJvqtiSH13moAoyppJXLdAJDAQetp/c9kh1iDc7NV9BrhMv38Wbw9p5hCEdY
/er4WmOtTtdGYO9A/2iqeqWs2XOJaZlnPo5Gt4wIw3sDBgJMLUAmqZMZEvEnqhFpqJmySGwuJtIP
bKT3EhIW3+4epvr0vbwJdeKRRbEgklPEEtzJ2Y9QFQ8UaEWT5+lo7uKBXLohec+K6azgGZHz05VD
dMyNChQzTI7u0rsp/Qt/cIHKhwUGTuQ70j/+DVFQ2KF+q/tJcJJqQFVX6Ud78yzjRIp7800leUSb
4upduI+Trfqba4s5wA4ZsOUt8U1G4xw4oJ3V0kgEk9r1U+BhDoCl8jJf51qHXicm7fiRFxuDJUMG
C7bDjX08wt7DkqWHDHGVkdqSprlDUNNv3svarT2Rgbu+0a+Pju/gmpgDYjOgGIeG7aWwdMBUNZno
CRFGHqHRrHOl9vXUB5wEXLsHccl74WSlUHDy4XXAgraXqlbI6TO3EcAXjzDpPEqG1thqJjbJ8/7r
pQO+KZ4BHQzQGUrhrPHnjy3xS5Y6m4D+9aD+Zlyz1uPN/oLOqp8j7B34TFNhMm4SjMYdubhDkJA+
mAzbvjUTznleOssKnVLfFQPZr9zJpaj+QvpzpsQJI+900GZP5YWE4SF9VHBBnV8B0hCTiVI37Cij
2/0QM3F/Cx/DwOFlrYyiV1HbJ2HQpn8QqrLo8E7T6pZbYkqGXzFNDNmtoGUtpVmho63+BCPMGWmA
XFDVkVZDsyOhRMIS6/po7G2yctjcZITqR1TvU1TBhiNbfwD7ricLM0Quj/jDpGbLutJqE4DKoVPg
8xUxJDTe5gscdo3fK9E2ZFY3VGY2/QCZEZ1I/PwywvHhHvLV83d7OaeWEG6CEWJyVE2tZJAS9zs/
PVSXwKS28q+5GaQZbC6xOTSvWIb2PMia6Lps6x9/1vIXUkV/BL7J/S7ddAhsamxQQ4TW3BKhKo3H
ERAVdh3bPZNCRgTOKY9UxV0QnuwUMg1WVyF81qhUuvkBFXcTUYhH4AgazamYxtYNMJQ98tLNwrks
O4M/hMn+Uk33s2Gy+w0wfdIH3nDNqUq45qXj4rbcqCBhrEVV30s7SuwWKjeHOpA2ndPRwH8WYcn+
TYphvcQ+U6tKS/CJIPFxnf4O7Iug71lXwPxNdV0ssgSGNy6tbxwGDGTKqbLY1VU3Re2r1kyYiylI
/RzBIW1RDVlRHkGy19AcUaPVlMHdkqxGEfqoRE0XDihdKzUJ6dYJR8WQ8ff9O/1yf3Tn7ZmPWCZM
vQ61BSjU/x4pRJ3A547olUstyDE3cM8rxUijegzsY/KifB9+7xL4ULTdag8m2ieCqwuXATfGMTgu
oh1jLSU9dPYdhhPOrTnapeQ5eD/z6a/AljOhGYMvgJ5UEN9Xta0yiFH4J6cRHBfIviBUZm/+H4pZ
Zu6bRtoUDWhtFYeRnnYdyhYGS2xqnIFVuakqIElm0tJKgCARQBelgREcH7MhiqaeY5PP3KQnkilQ
Hes982vTAJrkksGcoiAvnKDtavUoVSO/iEunVXcfwODM/QKKhEywsWZ0HHscmfh6Dfj/+T6HoTgL
yxEsDIgBTTRM/CBQL/7brVrovFNXgJPzzETq3h4cgkwZUumzGtXaMMN99zmR4Nu132VqT6SYrstP
CyDD17Na2a+YaM+yeHNarn3zlMEkov87Z7uCVFjX/moqWZfZu6py19TlLDTj/H24/ArMY6m92Kxr
ZvInr4Y9/3e9kQMdNbQYbvYmMf8/HPhBL1FTAqg4tYEPYJcgLMwlE8eZJSV+V2ktZes4odzW2q5f
LP29bbPrNwdCKP40gdWCjIuZeoGZEeMGIihwJXbdpwPoX2zu6/0qGfrNRIduqA3sTaI5zUTIXJCR
jbjBdvqdSHyOuOq/lb/VDgN9DdZ+hHzff7mAkgCuNycu8R9vnGNqc24AyX/YpdZY1oNqEQVsImAM
3L//nbyE2rGUlzOCvucghqMOXcIv4hThdXR27qFwHpBCQWxugjAcyLWzw2s7AbfKi7+TfwRZGY8Q
MeDdbuWFq+3cuJnNFgA9gdND5yQ6Ik+guU7yQeOE3dzi+/ECbhebpZgkBpLMrWlcHEko9Zhu04kF
ghPb3jmwSnySaPd+7uAi9k8RVYQT24yzMbh3ntrjaY7h87Dyga9TUh/RrJa91i/3WnZoDEWElhg/
iLIWZltAVdtw3IPWOK9K5wdgh10lJ1tqTgXKUofn1pjxp6XnDt3P76PrxFQB76glCwbcf8vqQl3q
r0lGy3FAQtiUMvgrImj8TdfnFAwbAHdkC6Ip13EDmxmvtfUhZwm3tKoRYGLRbsHjMGuWgmMNL3ZL
clAU0FMypqshNeOejtwWBNAXoQpH4LMWAwEtEQL0y85j7BZXh+u5EL4J2nQS1C3eBAZgD1hu+8Gk
6RRcoE9n+en4Jqy1bjs/DGF19LcbHQV5hY+8/gWXhKiWOpxVn+ANah9Ap8yBa3+su4I0tLjgqvfQ
nZie6N8CgSU0GVGlECIgqaeA+ebRcqxyPUA/UdnKv5Eupg+XYmE7ncvE54b1EQi7hrNiwMdXsavZ
5pOnHn2LnypB/gj/Btgt/R6Wz7fqjy82EwtAIeQ9geTn5l4dYtucR1YE9PxjtNawX9M1fXS0N1n0
mfbtmY/ZJkb+9KQE9lHEyWo51ni1IMcmft3P5qK+OypQBCcnuSa6ijtfw6ERH88qEzTD4ruwWPIT
vEZtJR04aBkEaKYA0+N8SKmYIworIfjmACyToRJKVT2TNocjAdRSdyzmj4oLGNPWnh+1GU6WVu/H
3Arsa41PgNPTbKW41n4Nztz5yORKmvAIO9807V/OKcC8QNMs9R1/QLepHTgfdl8RJts9hsnBo2mb
QOcPCmhTBZT2YUItm7nMQDTPdNZToC5HN55u0lXevLq6J8PlgiPYoEx1WkEJ7As+HJ8zMZhQoV8H
1stT5NsDwJUhCdZzgtpMy7BIGKmh6aqYxp5vQbnlEm/8U9J7HnQ4NMB3gjZHesDl1qO5mgpYvk5q
Md6w44yTcM6z2wviYQ940Q7BphpTVxh6y1fjhckP5CTy1U7Ni7XxZwKmFM0Jorfp0mFdX/6s/kL5
lFLFnq/Egcp3hmESwo+XRjy4wiR9d0RTR6kGyq9OpseF1mRLWVgPzFeVO92olWPRmhqiXoDWcGn5
SITq2WsxNCnMAOqS37ek6Prp/ZiLKklEPO7xrvFH8a27YarB8pDC9Ofmav/IIn8Ev3/9KuB3Iy1C
7/6JDs+JIsT0/KVMYWC1cNAtp8CD/eFM75UXzE9udNCLDCMe67Q34OP5aTgXFWgx9KZWIgoQiTC6
ECzeT1hnqEq1n45HdRP2dZFpAe//yGbqpV9zchHwWGdFJXQg2mHn2NSWXxzZUp29Enchimeaow9Z
IK8V6qTo643+Fa5LGD1Nluy059ifu/CRzDcTNKYAAyQoAB/uGaW8nHkh9jsMwLXPGMdQo4sGc03T
HOCZXEaYN7BWXRW+VKRqAPOa6TynYlWM6Z0UPpLKeBW47Fww1s+CfyNe00XzrAz57NjV32KlTNN8
3tnOEBzI4uwXLgD4epR1yqBdXvM34dH8qQcgSDFkrGjg9JzFpgKBsqncLVvYX7VqZvn5JX7CSDLP
IQza4GAlmNGNmTL0+kSd05WMLgXewm4D1Y2AzBao/qL6vru5QoPKHrlso3Fyh0elGafJMtTRr6lC
azISQZ6UaUkaxc++Zrc9vZFVUHudP4M2jkaCeYqoayJ2lqr0FQcKe9IliDJUHrsRHa9okfRZv+iS
ezFjhRo+S//cNYf+2G4oJTtXwmZgSyjEhNbPdQrE6P1TUgzvYU+cFelPVIJQsdfet4jXC/CJNU6I
NTaeD4ypLCLc9uBA6aAt39dtdzOtiZXnXN20/mg/GzS2izVzzX5EOk+ajgY3qb6nmFLv51RCdJUA
Ph7fMHQjLT8XUyWpJ8dpY3itislAB53lEtYH2R8Ii2Lp+m2h75lPWbGE4xFQ1wBzhkU1I31Sw6bl
LGPxziWkxsKNgqD9z/xclgkPXA5DFVszKbWPoK5RT8R/I39Att26QG2htqzB/IG4OiFkkJV/xhR9
zLew8lJhEgCuZOgvnwUS0+J5bDNMrbkakJZ3ZQC/3aROWeNpdjB32+aOvZSbYni9+oIqyUxqyMqr
UT6vOvKJyZESTYEmcgA5NJvNQRVSi4ZJrjx7JjBM9TpYJCtIuO9/2WG02TOaiyBmkJHpGNhr8hiS
k59blibpONWiLbQ/jbpEbiSHcHK2qSPr7y/qAEbkBWg9vHgvfw3/WLmkoNawYhSsPMhipGS7iT5z
IFLbC5zAVnLXBmasnrGhl9qjX1a6EamaFjvnQ7yogGfyWg1TZDf4RZyAbV6mJ0ZTxhopJt6D12DL
O7i6syiD5XJzyzzJtiuXu099fj3nrfooXRpE69kcDANeVsV7+EvddTJ7RZusiICIwi78eoq4aDxT
JukRLBwmi0AHiPLwZB2zNFIPLClkzcq3aU1FdCTuUyUGS1OSYfvsGYY90ES9j2Z4KTaKQo7T/ftm
Wd+uAMy3L0gzHfdOA+Sn0L3Jnkyzu/RPpdcJXlTT5Km7w6fD7srRvVWz7a2Yiimd7pMqDgRaw3O1
2FugFkmo9pGlMNcFBSFHetSyydQzutPP7og4dfKt85moYPN0tfameVjO/V0ErDGig0LQQz7YBt1f
DJmxyZq4RDDjSeWQfLJCnOKTC+4a/bT0w2A0BkGedUrnm0Cv1cdyRSfQAZdrl2SLzJb8NNvzCY08
XvI1e89KCFC5pj42QiX2URePz4VqRAaOfnp/aQydrH0G4K+Y6tRbuYz0M3+rdmmctrpNqzvb3cYM
um0PVIDGV8WRe0liXwPWRJiRp0Iski6u1mrf4NajOPTmvTt4+gN8FuZU/YwVPUSe6ZzqS6AyhfkQ
3e+7dxYZzSNCEKvnK8DaJuwfSJ3qBAqzT5QpWm+RYjCw8nLSLXbg+Zg4bN1KAuOiJnzUGfce7LEE
Z0AriK3KsqgtdQ68Jn11LCy2nXoYsBNiKQrpKydCSd0qHNZz28eK5whtELyY2xCABaepdVWtmy9q
EUdxOPUgFfjsYn8tYKV+y57mx3mGcKEEK9kXumCBy4sCF0tP9MZMDileBlpD9Ny1nQh1Fp3Xw4RW
J+dKH+iHyZMJCmBJQsta3gOQt5KjVKyvlCwkPxNPguFc1/jgS3ibuTldus+EDtk/+nebTriYysIt
tZC/OsPlvEQnu2WE5r3NuiL1gbudB0oQryeeu8OSHmHx8ogCOsdZPVAOtveBzNiEVE8NdNTyn5BZ
XX+AJcmV4gR0UU36MyRk5hQ1bA7mr2GWtXjvujuXhlwyf3dkKPvo3p4X4a8+l9P9ROBFde/9dAl8
JV9+2XtOFsK3WaOTOkF3RERXdzucsaEAATPXcjhbbnVfwwbWglMDHtMm2To0HIvD2KkoxTDJsfv9
+EYGBvyN+JSEUaL4tMh0n10wAwd/q5uHa1YVpalhCB2TFaBR1FdeSfa9EU6GUck+sqL//SVOwteb
5+ypXFUBdpaJJbYljjUXVxctsT6V9+CyhBga4qSeo56A4ut6M4VFFb29BbdjU3CbdzMElTOCkFHk
Lmty55k0/gddqvv1/kxX+QkYtUChnd+cnVZCZpQ5ZxJ/Cc6Pf1VPZSP9tbnnUZvEhMuFHXDkgOfV
vKU4qrfUEnv/wahITt6LlN/ET0oaS42Q3bifhUy5cdryqa5nyULAARY7qfa6ZbOA+Pu0lZCRiU0y
290W5E1MW7D/daXL1yyprriqZbgVjpOg83q9uOZH64swBYdqZhEAb2R42pFsjWXX6iP8hQpxGIno
tC8JNygwTi2Qha02K0DV887A3q8sJ5pHrvz+nzagqxn4brV++WMtP0Bj0vUMixMFEda8RoiSiAG/
NCUai72xp7SYP/1OLG8ksLe7k8TMNC6NgkwaBjoeqSjMhBpUaEMH67REL7jzVepcFBJwu6YhmPpu
pMF7X6Wl3QqEuJRT9k/DjgLPOP8oVklkT5tYeNrVGr7MAaiiLE7uFv5Kpym5jTFaUVhxa5B77tm3
2NftFAR0dwvGlj21fHd9ZdaWJ1US1a0m8Q6UXwVj10O2KcLI9Pgu61c5we72xs9bkhGdO2AOw/Es
HAoAITzW/ZlMvlf1bJgFItQPHaQjrzMSrGKUQ+4ONDGonafqASSB0cKY1ounxRoVnVTHEsDEKmub
xxWyJiXplCoePcB7yQTicTzJJgtNR44lfs88uPCR/6/Sr3Kinp2OC51DizR8+hp4hfTgrIq+3lCJ
RNAGuFtZLtTBuiT4ImuuA/XOVBhot4lrC6BhGr7CraCbQA//53niljcc57bwRfHuqPA3VedcBJsU
ehjsRn8m3113+z3x3v9+1AJgSzmhnKFliOTSOhUEb26zxZQyPLAbhH2aM5H4KtjZ+Z2+DdlcvrRD
TxACYZk51lqhbdBUCY2lzMDmZ/uGPdxuaxK8xCHEwjwqB4IDAUeJZzRpmX02cSHVfxv0ulaiLjyr
0XXTtAN7mZWml6qynKXpZe7xDjs7TdDdKl4cQPHhZHx6aPJIjzFpAN3QB0czqDW91PieB9yJZw6d
jj/S6G0thNvi4TK1F7HbqNwFrN+90q2dKLEpaXNDg7ZCLq1HomlNxASMBYtezxO9HYKUdoY/LcYs
g1ZQhTafpehgYWTDNH1jrQAtFB+2tFLK2HH/d3xG5P8vkc2xPBro0jMqyhWt6mpIQwNEaDV4b6nl
2wdTNwvScSb0gdLOH6baocUXA88J9gyOyOLKsJeD9OgxMj/SezK5W9efk76UGSVDHuHil20CVxjv
0z/jwQlkLM/81mx37/a/oPyRrJMs1iETe6feWQHiAAoDR1+RXk0bgnrW4Mfq96b7X+y9B2xDrUTd
ONOrOIbezK4dL8KIYmG9jkvFRT2xHo3QregpPTlSs64ZecHZOKxEIUV0mydsaO57BpRqOjzSUvSj
FZzuPcRKbssKLALY7Pi10xljONQm5bmRvKOO7kPXTo8HdT9j/S6FTLZKLbXFLyNK3akgrxvts66n
VszZ+mzTCqUAUgSjGpxkNkxNSkHNPqy5bS4uqsxBqabxXg7buwBzhL2oRhdPT7pN6zlqLcggGg0U
bV33veG9v8ljU9k+PIppK0RU9s6MydNqWw61QlHY2OI6S1st5euNNp7BDHDHMN0F+vMqc2z1k020
rnN4PZqcii1ADQaKURuuYeuZ8gjZnCwLYkE7m1HDcau5pc7Upd3XUZeLmN+4jwoGC/G/3p38vxfu
2tQGvVPTUZAjf1Q7rPRo1ZlZ3iJ1+4xEwa6UHnc99rBXD9rZyDuuMgtExPc4t6Er/oqbB9MjXgJE
nV4GBPQmN0dLLmQOzU5UMfFV8KfGCbat0mk1esYTsTXQSJVIrRqTihR64vDYwxKLFOBpNCuuZ5s5
R/W4i7FDaP/fYSG3fHuE+7pl1ahdxBn/CajeX3UsYQ9f3TzZ9qES80LcatfDj3j2QvlEuHIT2vL7
DmfTmAgVoexWqJulLu+6LiYfUtT6mY9XJYwF5fbqAsOiJhl+gUM62FHm/f3VUV522/MOVbHx4qCV
rBRxqx0VczMkYW1a5aZ9wQUj8De3EvLRSPxWxTmVyX3iEdAQ+pH/aXdU8y0H7on9BEBj3mSGHvpL
AMgcrCHZw+1gpBXRxIf/RocRAR7Z22mmrH+TBCLMHvbNxuAFCQRJvMNOwAM8nt8hN1bRhGYfvAr0
Q6dMruMxjhFC990fEQAb2pKbf++inBno+kXPd2ouZ0sVsx9KLLnQwA0KRNQ77LCwKLxQnWjiyXbU
dptIo7HZaTtC/uRoXEemdc/mZb+dzx3j28fS/pgVSqmFpuzd37NuG+j1h5jj8OqBKKnqZocnVMu6
QuNozmQ3Ad7rq4wChhvzbUJeHdjp3SvD50ONx2dMnhDqj+EEYJoaxb1Txq1J6TFFREGLnBB2f4kc
Ux+e4Z7vlCPhH5KhqXnJi56ZrFL7EOXNeVKEPZ2S/ZVCA5OSJXDStpMRmi/4ftSLK5fx4VifsSnr
+l7nw2I/t7IS5uA+4ukG3gSUhLa61Jw64GeF+nfcTK2oUUdb97w9hcbDJ8b2x/08Zvxtah+GIuFJ
4Vw5mY8mGcNa19HMTIvS8pvHrAtfCrpUrP+xln6kvkSXnDjikjJns5ARj2Qn3XxxCDT2+WSPNlm5
MRileE7pJlSCIH64qaY47Vq9yKpvGDXdWNHLDCSvO2oqLtq9nBD4Biryk8CpfbFwAAzw8igCCAcD
748QuZdhFq8xBhveq/3cBpj9+y44MgmOwI31VuzihYGyNjjgWslnokOy9U1ygY9WyE7oM+RAacgH
eiONJnx2O3tLpuIU+NbdxLOq5RRQKQPjiSDO5nq2IMMr03yUcCV0+mdHtruTozGN/9DLH2CpnYI2
LFMIfqbAkMWiC6M0SicHrs7i5pDJZzo9vllcOUpNTCsSAJI7W1fMa8ocrsqXsFmqcqwj72iBYsFT
bcy/3l5lH2UNJQMP+ZSB3hI0xvk8ah/CRd8RXTdSuBW0gZR1kwAV89PXd9Ck6ykxPANk0kbuxwy5
6BRzGjBI4JtVCHJ0R6q0q1GfC9uorCem+vFyBt93Py2xgsLVDbLmkyN7ojLa7MbxCaLgLZMzOtRl
btDs0BOfMdgecEXyDFWcD6PbvPtvda2njur9mk/qKKddfG9q7af+7pg1OL1GBPvdhdMHAacivGcE
4wAmJ/0opuKnbm1eUURYlf1SFFIoAQcoRogmNPH2Rn2wMUhO2b4eMOIRKZFx2/I2zF6ziHOPcUGk
HfE3r40KQUBaI2xKAZQXoALg5iWcAxuDdlz1XQEbnLSwAIDtTG3L9P4QTNsDojZKdOdLUqhkaWQm
1y+QQZMCO4cisrILfYcMDigVZty31r2he4Thwwi5xxQf1/gIr/oQitz60DSVstYeCMlMNxXSKtiq
ZKbVlHZqc13snSqtpnFZZkWerVZ+lco3ZZTGR2GTY9mqQotiX/yb7mk1nSlBm7cxSNHkMzW9AeBK
S/qbaYPh4bkqiq2pshcbx9VeQGUP5BdzTtGmaouJtf/0Xo8/cnk0y0r7SxL33QZ9y5hm5x1egVQU
C6WNI5cF0WSfeRmbArLXTyobhSTfIRlf3iUFNtjOi1LElU1tLtnFsmPSemfvmvVapTgJhKzAWeCE
VgZWsHTzGXZG7ybW/p8uYbvKPp0ylDlnXnYVUvfcBIoNOHiMQvgy8653XKbxH4jKS+dvArNpWGZK
Hib+t16PJniw3qElPkR4fCzRdTKnq4s3XY6qbIA40FfwNX2PZQYwUdOzIGcJ4lOOnaUI11AqBjDD
koIxfYvYEb57j8IOaTjPXayWoNjxUguBisM3KGnh1Yf23EH0iTGLwMdNbI7lzoKEb10UbH8upUuI
qxmfNV3sjS0NqdYDylZ2sZWcyKbjcvGsAE/f8NOMqBm6jq6ZyX0/10i2hdL7khOjpBJ69JFzfC0x
ci0wEHBJPp0b6C1V5M4VxKRP0AOI9h8t4ynu1Zmo+mrGi2ROD5n+Y+wwA5EiF7slH1gB0a7Ip6eG
ygzHmCmGJeGtKGH2vjBWYlEpe79BHd8o5uqE6hNK8067uT8YO4w6cBhnNlNq/vd0v2EXg+HI36JQ
z1WGbp9NH6vfQrbHJa15gpLoNqmHHZ5YvgZllt6WAryLR4MCMTc+BgjjFFVz9S3SdYTq1UufTUup
3i9K8gSMpymyT0/A4KF9syOpWGWTOY00BPvWl5vnLoytgUbCAVO1LLVt/pbZJGqJ+JjSWCwPI3J4
bcZsxuZXCy5Plow5/hMo+Fr0e8xsYsm/9LVpqx4OcL2EIqXlUB1zxcv/LP2UMe7Xa8LrBflHbpTd
bpLkuOhf+lUvbxCU9+rcaKWdSpvEARCPBh9ho8B9ygwP/GsiZZfkxVWX4FXClU9/FRcMN55FtjNn
bzFRwx+MAZTZXLCoEidNYkWX5imVGKkisP9XGOnqB8pEKCxFdEtEef+L7KMVBjHft55O+OVXKzL7
xLizX6hLcJr9feUz1BML6jXvDBADqNyOKbx66N9FTh0o5d8DMV4UN9wnrBqnwj3L68mQFA2XKSAK
B3JeItF4auD5iTZSt6I++qKXwIK7DjBLNQSb9NxJ1E7jCBOfrl+Ekyn7CRBC8hf1zsODXOPkZ70O
iDJ/fIE0vWzdK+DpExp9mM7zQrivKHd+896XWeMVQ/kiECKNooITA3Sordy52MSOpsL85EMX068U
qXWzSCzAWw0QyqGxvJdwBsYqxpYCpR+7ZSGiYa9fnNbyTgnRFZwaxzqCEL6fOjI5m8bm9N35rWNF
YCU7RjxZcwOtL8tQetweWvLjkaEbBgmRZrtvWnzaVmSgYLyIO1yfnUVHgBu6tM9WyADQWZZe/Fic
zr1hshH74FfPpsKrWcGuuXR/Osn9ezVcHAJ5KFsSkfFIymCj7rYZ+5q0vViC0uN7RMpfiJfGxyU+
79a3ohgCvwpigb+F2iMXtZg6tTi3/AJNNuFxyRJn5F4PfGUugDZueRRCpYwby+Z3jzxfDZ3mrW5u
vdmvPQ0BK2TltGoatDD9jFakeBXJv+3MAHW3HoDJzjOBs243nb2uE695JlvTgNuArynUUO5HQwjQ
KSz+dgBcVQe4ZVWztvuWBAIIWWwA8oB5s26wurl1gGzcMHrP9GMSgEndulG34naxGMGHcXY1U1py
ieQf2cZ4UwY5MSePg65QWXXMCftOzo3hwfXc9QNN8vWCZK/flLobDf/z3PY7yyooRrmXf7C4+QuB
TqRgiYxrYlV+ddng4xmFSHQDVzUynrr5jwUChmvrST6RucKm4TwSzzpAEyTJAQ8HbH16lxW8Twrm
ZQWhB2cVTpWHAYmEXUFrTt/vFizLQvjYMV0UTznaiKOeXgK4UUI5WkD1VdWFSIeFPW4thsWBbcZ0
cD9GOcw0b1knS2i5KKKsWa5i5Lr/1iUATaOeX6tFhFoss0RlgEBcm7OrdLxNwTS3pbyOtWoBeDP0
Do82Imsf4E4RaogwHKgjcy8B1NbmJhOGe82KyPGswBSmpC+E4QW9ezpL2KwI4Aq56MaKe81iPTbD
V+VunwgzhFLKids8TTAZoouGlptWm7iTexoybxV/sJUgo7AkoMi/9l3fdjy8xt9K3oTwErT0Nvp9
7mY+e3iAQdtJ/0s7/H8Q2HUaLZ68jtysnq4HGvc405T2iEsthF68OL+NBnlhU4lV/e+NhsfwgtZa
VU//rmg9mkjPhiPTRrH7jhs7UZnZdpDvnfgS7byBGS+3zqJAc2jegeGEnyPzibm1jQmFfohv2zRg
FElz2UH6p0z3WdkVsRBNJKDtdmfJkJN8JdcVzrE6gkYWi+EgcdSAc8SRdqzGEVRMHXzXKjSIG7Xk
DNtmbiMFD6UwxtNvD0mGRSk8UkZz9JQ3UpJmUg3M4hITVM+37OusD1DB2UqHI4W/hiydV+HovHvF
ro6C8Mah66A9BZVHpuge93u7gINCXdCpa90mei91U2mHx7qF9R93lai7Kq1e9/q4eFwYQWhwB/yS
dzRvFHRNTbaNiTalmVQB2NtVBqEgHsXY+k0HQGIIJAwIBlr+DP4aZhmyNi3h9MwcgL2OYfHFcScX
A95F1r9nNZ5B81V4LSsI4xCM9Of/G9il92oF8zoS8SsZZMAHQpSdG0KXry7bTYuO13sHsMgLsx2W
XV57Gv4CR851CvRAMa6myE0WtfOIfQ5wRJQVyt84fKxh6km1vXJyxRzSiyU89fJ6avuZbmvbUjBH
8dOaG19z1B1Fj7fHIXLBLSNJ/ytonBaplawbHK4DlJ6qASlSWujOIoiY2Ve/aBQCLxQBEmyFGZ+U
cs9cNfC+KfkVWmFGHWj7Nf9cKl9loWsWpuez1mEVDFbXgOT5inQGewHcmDFkVPIOgxUJVS1nYI9u
dour/3QsmbK+nazmi3tAwBIZ3eayhom7uX/IUc7o5fRw3Cf3cy6qsvCnUn2vAHEptBRcgHXjE7AW
kz14/z53ME78yxMUt1BS3fETZtvbe4q1Mexu5oCsz7Qi1ORTiJoVigSnT2HLPufkPIKdJ+9Ipdgk
wgZqy7AqFBo99cnv1hek1Bv3NH1fqVybHfduvhxbGC0ChaWle12yDSSkHpbiKY7d43PnKEYN2d+K
Ifw83ZSi9PRVICOn2Fn6LGokTwZYs2Yq3Y6XWeFLATCkB1Sjq4vwVzJfGky0mK9AOuJeRfjhVhTN
G0L7nXUnkwnkeZ9BUR6vvkxN8lu+3JGySHJAjf5Y3heK8DUU2VVsWbHlI0NOQ/mAaJBJHky6qxpZ
nNq4L36an0CQijTcnckbM9LHGFxcu47/3SbVDjSF+G5HDQj03FDar0JZ9Szfs/6uqi0cqyAAQkHW
SCoYATlS4kWCMIyze6dFTR6Vm/eCLMEV2aqBAkvwa0lfd/009Tn4cYyRwIBtxvHMOcD7lwa7Abg7
eCh8/5eTW9zY4GeGGTRlmk97LI0DLOcz/14Zb4qyA9+e4frZQ+OI5c4kTFHOvVSrdaEJm9ullZOD
cHfG9qdIMtIe8XcaZtDrUoEreePOrN/bft5i3KuAnX6trU06UO+OXeLzQdzBq9ElGFe5Gv+JaCrR
i1uUU0KvsbrgrMXHfPmzz5KGoio0vSvV3a5AjUd4dy9tf/s1UAa5V2kyUTHBFMJEu7n6t0IZANgt
i+p5z8b/utZR6cbJULS0fQaN8FHXFFx5qu7hlPemZszA6qOgoMjSE4TCkKyWSNe67Wz8RTZA3lS4
jIaq0z+qKTxMwVrFsD/LysGeeci01JUSDwzEpa+Pe7maXf0ZTxWMMp++0MAmq5A6FJAvCvMuDr92
ehcKt2GrYy8atl4qXecUi2Z9qwubZkHSCBf3jKt2ScM5rEnj3/VZQk/8rCaujJMq23UGYnFh4a6W
17ulACu+a62fWCUvs1PMexexRDmqc5qRCwC/mSCFBK9yyinUHG2bF51jCaAmOkMdhcgCAfsdVjYE
3YsPLjrESyjXEV1url3dFh+3MNsGGLUDpmYThCxDyXVudBD3ynEe5DzHaroWCvlecsoQOSsXMwZz
7DoG/J29tJs71FJORXXq98Uns7N484Y/GwD1CgMaexUvukUy4oqu6iX9dGosmMIr+o6z4KZ1biOo
+xRuPsgh1v4lfKhXpaocGrWXS4qk6qlwWtzOXNhf+ByhcBmdDU974pOBsmHCr4MworN/Wds3Bwvj
SI0vDKG6b3kVbvdOvPhIK4ae8X9Ry/i/PQNVBThwnA2L134Qi8RWoo/VLEWbvMoIK1NM//tOciiD
TPiLGERF9y3THtKQ7o8d860rzAkDWjc9yFw5YV3r93+yL5rfxyO2cnRzAFM5IU55Pgeg2Eqj/lGE
CiUP7Tsa+VZbnWfIMYZCJlEeUB2WRla5U+sVqWo/ahz2zFNGg6rm+zlbzdMMagKdBiIP0CIKK6Vy
acSUp5NP1PVLbI5daWLfB+FRfXLThEYOVoct9ZwJdAfOfZ4q9tz1hvvXqSmqTEI4HNB8TJg2aOjj
zb3rlNR5rBWfu5ge7jDCUvsB8bP+T7zkgu0ruP9g1DdRC6h+VksbV/tWIFs/fSPNdsXgHJTNRoSm
OaVNX236vevoIOvYdbsOg57Tb0qTYtj7SHKOskkXMJ7MUxQ+JUrFRtkWoYWdH6UrUb0UP/S2DIou
1QBrXs9DD4Dlku9xrU/G8xkTZRp/YMKfpFw0hhwTYAzjGDHI+FKMo1zDFJ7OHgW/v+KfSMTdK6C/
SmnQ2X9l3nrRRFqXyXhK5dBxIwPGJr2dOTcm8aXemN4TfD9AxUzw9tFPFwRS3fMvJZrIJOkh0psf
JiP+RTRGTaOSo0PBkR5uKoPC3+f8IrFPBfvQScVZfEOPFC0w6gWJ3ToSMmqx3cwCVS/JH3evANu6
GXqRJfWqbRXj0Twth/tNu0upolSDU2gh4Uy/cCBgNK+7mjxZf7ZgPPR0X1OCv3rsQ8QGWzVu6+3g
ysevRO7KVodtbBoMPmS1hcpBL6zGrYshLCqyZFkQwrhq0sOBXKSIXAoeGB54CT0yqjkQIWYO20Xo
GcyoDCslwOWFY8defrYLbbnP/JCZVmxQmoxyEPnLl633kwDoEQ3GXpdyoC4Sc2HmrVWd2hZXkgR0
RQZx0NWn5pNAminfeH2Kn/jkHfDCT+j9FAqGRqhkQK1pCfqvyX1IV+j66j1glOJ6YwK2ectL+NxL
vGl3dr7ga3GdHPBoYSTgLoShBQFriRT/PA8u81CW/ganVXNu63RsFnoeoTLSNFVIm8OvHlZcwefi
/1NKByZCLA9d9AR3YQKPJLh7NVhaP/2QISWA9hTt4VTlIhyKZwDxXsXO248WlMWi4Ph0PXwFDPD6
W8bhKsHptnymBYHVFFmRVRed3wpESOKRHHdxYwtZcboxwMLGDrWPJwGUhOBXVPO3B/BAomTJBk+3
ogsc7nt0Y8TZ7JulMvJys8AyofPe6bU9mc19J5lz1GhAd+tCi7T1366h1rAQRrT9+vXOf0qKRpwe
MuG3zSTjQme+o0M3HlLrGZIfOVFdzyTYi/RFSPjagD4TJHwvL8cGntwx5xlhhqZTcFEwLOVZAtGN
sGL1K5RQGkOJK257AnOyv7ipp0Opj3THNPaOY2I0ijGEiQV3kVsUa2OKJCO9uuqxIZx1dvN4IruW
83td4fEhUrj7CFTm3Jt+xJBOwP6ucyyoBeRbF5LPtee9gYQQiZodZp70Hoq/sUm1DB/6bbsM493V
gQm8y47FrIKE//h2kN20eNDhlN214wDerWXjWj/m2Hn9ErfpXLDKOrHPkYAjp8wzkOzSB/eBlEsq
BsB2b8QoMCyItcD5Vl73iTXbY91yMRv0TX3oyrc/FukU2g8mZ/ReCiKMiif3s8x5siBfEuXdYN+8
UA0pIckssV5US0g5XhJAwJFo3qkgZlHK4+QuZdV2oe08mnGnCjpvQ/8COqG3MocEac4yMXOkbkvs
My+lXXtSSdmyO2WO+5hFMBOcNUWCtj7FzAtzIsIf/CihEB9TpyOiYAcIte87nS40pAJlKILsitl4
hdRtNVVwmsvsKIhzbZJsLyAxkG2v0omqfuMdoXXr4uVrQ1DfHGsZTOeTsmXZaF/X94f+VP8V7bFL
5ek3gC5VbQZ3QCocjAiTd06lYEMMbBHj/EMW3QoYtaIjxZoGIsr+O9UuHL446QAqzAh+SY79y1Yg
fI0zhCrUnl3AG9OzcnNDEmG4YPthlAX3A3e/bO8tgHMH6/R19PiLC1MV2fQzPu9Hv8MWiMJMO5+Y
lEd9ohSar+x4lu6VoFEjioYavC67yWAnX5wSAFthoL4874tZfiusxMF2ndBOkWouaeitPMM9j2mf
WID1y9pKadB7vDTkeHGrMBS3cDZlCSw5yU1kNCueUtrTCA/7kb7QiQDvNubY01BPJrXn11ltq6Sj
RPoRmd7i+AOP/MfjUv3BK6f2G0ihlVIotoDK4hHjYzHV0t81R+v2XMp2JUoUTq40xDZ4VfLwc6u5
EpwPvZQKO6GDGSyshHwevYUxo3m7ahNFPkNJiOpskYCUsFxU+349X61VRBsHGUdjmFH9eaOwQGJJ
HfsBXTuGqXeFjYlVi1CRUGKYXTC2bBsedisxcAAlZ2BERVazleeg5oDTj3sskFH56X8Qk3uSWsDT
vMmrzFbrVB76i+saI58UX4KBF+2W7Hi7NVzkWvE0j0T8+mjgSJ8+svVLCM8ejedfeVNUp1mJLs+6
74tFCu2FtGb9PL2XqYZWEQarPDCxUKXot+XPvD6LuDPY/ByQKy7Xcam4Jmsj5/VbHtEoEItAI9hy
Y7Zd1Iz76uUwwKUluFBaBa8clHLN4YYJNAJ+M9EqjmHnhNC85qLexvKGcDSiaBjBn9AgvEx+fxew
Vr1hroIKboreRxBAg26ZdMufIH/JLF+q+yKRGaMV48d01Y4a2KUb4RvfMjQBRBxg4NBKHhJRX8ss
PKia3e5CUsAEHgUVXbSc+hjmyeROmP2kSnA0sRvTpJvearONqP7hqkZCVyBYbwRlqTUc7CojXEDH
FZZsubYW6f/5XvRWCmv5dRU2hjRFxDmFMvfcTFKu96MayzGrprM6va1sZmmELnX7crnkyrDQglom
Ef5J1dso2/mJmESq1Y8MVeLEgq8e2kKeIkbMVrpsGaWcaD8x/UWu5pFr4Mk/dIscy0gc2u89gekL
WIAXnoH1mr1OUhvgjEdAj3M2DCileU5NM43oy7eD16muyaZXGP9ZLiDSz2HEZqlbDlouHS7uB7SY
C1tpPbj9SUY/E4xkZFgPBSNAxJiPHZEorlMcATwuk7es1X4kegMaSLxToaSeCEyNMnxmwehx+NMj
FYkiSuzdoNXB3K24HB4q3ax4enpLVMVyH9x9IBNoqCj+H8d5lItkgv3vFMVlciVR8gDFsXZoqHsA
mkMnYXMmkSEmIVSf8zY3rLpsVEqKe1Ni/4gLawgHeL6ahLNAFkXuwHWo3iTDKmVaXFE1+AeRSTD8
pJUpnAPFVs+vjYNpnifVHCsZW/x6fyHQ3PfotmxEG8XW6srnEDV17SUOAA7Of+vMb8X8MueXh1rw
ScgY4d/5cjXrPVXNJvPu4dOkxoNZI6z4RWtmvUXBcE2ypoBSL6TVn7qysPGDzUUoixD+n19EDQiZ
IxD5tPpdgzuphTjcJF169RVpXqSDKuImlkm+5R31l0+l0YVNH5yOaEia2iFsKiPZOj9ZFqF8hfM1
1lP+kq0n5xQuZE1ZOhcaGt36X9jnoluHL5vS+OXb5zhrmmWnVewZASgDKNw0JjFUaAqzQiATZ+TK
Nnd5YgJ4AyP386f118hPqAixPit9VeAgaIQAuwv9SuJM/PzqHc5wVmVNIJzUC0P5jyPrM0eGJJcP
sSaG22AT+SULbSCVLUpS3WH7Ues6l9P2Crh/06lGNL+CTlrr+6Ia4GgNc6xEjLSnO8ZQjHK+Fnh5
3jXd4+43V3QvRqhOMOEHIMF8ereF22idrV3VuTwfMa4N2hVv3GznQTIWpFTCsCUY59LLob7TrkAX
3iLsB4aAXNn7hgV1T4j9nXyvP3N4jGjFbtDpJ+pWTUIsdr2aINO4znSK0PZqjiyJntUxJVc/rh5A
FOTrv/8ycXUI6OiX+xHUHCiOCzUSedpX+9cPvnK7xVjlytkLbOE4eVc1UKcafJVVBnPThsgLaib7
Rx8VIk8Z7cZ0fgetRxFNhFoeVS19O7WIH1un3SFAw6PgKGHKbMsF06LrENop1aCFIZWJ4Z8+l4AN
ByDa1L0nTAt7KuUL6Z/Al90Sfhf+LFTdirSTY1WiFEphGHVU+ePnO9Qc6yhuSQZhLqEHFDJzohjT
H9WFEsmeE9fWpkfAXRjMCe1/dJ7jSZ4YCHaXiqJoX4MfJhUrmzHUcvJnoqWROyeYg8KVJC7MjBBo
UiQuSlsmAZWbAyRoiJTx0aJOEg7GPcv2pzS/Xyulcxw9kPyZy1AV8D0sMqTFhELEJawPbm3h+w4H
kjCj1DVhKWeV09S51Lnn2lDlrtvBsk8PyWQ26HDJ70I4MIqjVZ2+o34dXjtaAh7erkSKdtU66SQ+
JPnEnGaHRIQE51fFOHMSZ7fWY0FzDDaO+RljkUu1/iBBWuunP+SwSt8027qWYM1W4Nsbh5kE3x5u
lLUgut3KwdSLOMR3nOYcV1sEgZj+SPlc3oqJrKK3HKviaAGKVL1SqI1PQpMOilIL7FVC/DjoloyV
dKviyAPbHZBNUk0rzVa2/lLSk7+EnkVBOC3AsEceXwlTLjidcWKFiA5A4jwVT49iF8L6YPzbD0+h
4Xj6338Q8G1Cb/nq3ljELXvx9ccjzYrRJZCBjPl5nBnmUazB9wdu7p+uOo4zCf3GIZEpSf0bDY/6
ehuwhUFs3iOVyTnOJ1G/CoevEsGciPgwqbL89vYOIQbbeqA0HrfU/pvR50RIfce1380FfrWBTAQ3
m8zAfIXKSFmtWkUL0PmBCAbz9xhvlg13qmlBNDI89u51goQyhEEmFMpNwzintrqZa9V8cp+fJFtK
283yxqmitcxHl59UZciRueVAADJy2xGav6j+imFOJDbq20q4Fxp6H/xU4ZHcYLAKwr2L0Ges7ntC
OpUeH2iv35NElyc30Ug=
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Eb9yXDd8uCgXSZTSBnFQ7R6ymSMAfzAuyQrgooTw04g+toP6bbYOy8Y5xsxyTvg549VEWmifL9ND
eMVhkgtSWRmV4n8w+WroEmQKN9hbgDnUaAJOgy/yJQ20ZVZ+gBZB8X9MG3ER0Z4csubCz7pJbkQX
ITG8UKDXXbwSf2x0Z6pST5L3fBsjtwyPgrAg+6fefgTc4octZPZNSIKQLDdwo4FNNY8QzlpQLXhy
VxzFZAa1x/L3On3iUSYmuX/WzFim2pCk7pju6LEZaF348YASvuSDWE2GWDjTjhh5LiRDgUQiCnGs
ibcZc3voxqpF1AdUhTjO2eIu7CX6swUcO0g1iw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21168)
`protect data_block
ApsHr1X/r5Wnjqd1Iy98/ZFrVRwdo3BA1+/wnM/v48coAV1XZycGOLS2PIlrvEgHa97BHgbCOMvi
CS12w+gExQkIulZB+35L+Dgl0FVfDRoQpJhzF8OGQrCSa7D2Uv08Bedsr8wro5uWpmeNg78D4LDO
RYLM9M47F1dxOgUxTQKlf0yeOpzDH6KLGmqdh82QmBPP7yGd2lwvNhqrkgoj24hYqA9C3Y1OWTER
mTNLDzKTf0c/vq+tPVgSCBn8f7H7K53lQOrdZxu6p7XMmArYFhqWEx5BhUuByolx55gEPXMDOqwh
CrHosWB8ndNddgdy12zC2XIw0XQfGif3WNz6+N2l+xidt7ccXc7Xv6c/aAke7wxOyhz0whmklvHQ
/NqW3SOTMutZW00iOaUNdqFMhKjOqpI/uvUgrCMEbr+N7z3JwKusT0busChwC+9U/LN8cGF3kTj3
PFsZs0mRMFpAUsSK6416pP5wlbYDotwNSZEJqMoP2rVDueIS4RMHvN+Kg+vkBqE3rT5CqGf5e/9u
p0p4Chzy9zJ+hyCK2c6vaa0BKaSdkQvHHZ4H34ZcDYmIZu7XV1IEa3tn7tjgvGeM+bzLWvvbx/nI
2zurheUzq2XmBcWJ4u0ZF0PSppgoYkC6OILmvoq84gJVY9sqF3SMRIXM5R2H35JxbvfW6twMoS8P
GmINAyPAGSp/4W/8St4PEvegSNBX5wtw01dE16ICfwXXC1aEJ18PCOhTV4gg96K0usg4EsIxUCBQ
eV1bQiuz1TdDlXCl98sneefaF5xo1MfZXnbv8LYTwj1No4c3Q+2EsDv0y6LlzBKvHsn+WFKKHd2N
31g/8NZEhls2wFk97L91D9H8apya2AqIgGt6WIhMmHVJNLJfk8P6c1EnKcDaDakkmtkreGnrd30e
ey4p1jsnNp6iTJSRyvvW7KCdr7bOHFe01BUg6VHK45hQd/b4aRve48VU6WAJBiS6nsAi2KSOP8Bx
efJrK70FhQNbpt+L00CIzVOKF4IFfwPgI5MHVHCqnNim26RvjOIYE4ESRNkaaHdPIm8XPijsRMml
W/rCX6MtdygWcLdk5GCXAO314c8hNhAM1Yq5IxniVmDwXwyT2vH55m8HnwMSrhIvigXxvoicuSuk
gnil+ZDK1D3H+VpL7T2fL8VtDDRv6SuxzCZQMlD4HGqld/ZWf6sTtoe3hbX50xOSh9dcEjXkjHVC
Lezs3ePwxbsRNOh2qSohksu1mMRKQyMItRz+k4F4ATDqXNGcm3HZea92yIG+yk87nq9PboIc94ox
+m6UADJVSrCUJyvzuk/Qk+zF7JQDRp/RjudXpkfQvNFuNav6cHkpO3n0ZeFpyCQyo9Lo7Xp3laVD
A5l2ig/yTYbFL88QKnDdXX1FxR0YrlV+yR4Eq/TkrQaol42rTlfcEGKMoU6sDBETsbGIpmgpuAEP
hoYtaqF0yn9MwoOxgWADzkgMfE3cNcHof+g8PgDpsjI5nP0Qe8cu3MTaIPHZuXBhjYvv0sAogdGw
5mTausK6wcefqKXwqmJFZQiYfe10pAbJl7SoIrmC5Y7xASCMwhQ509QXT8942zYsQnLMH+ixPVOl
FmfPKHR3z3R4WHDKn27CnPlWsIul66NedC30xsTU5bLgWpJvahtaCnFN3fcAChmRmcAx56IBxeq/
2WrMSE2aGob9KiAYHvNwGZYe+vVzxU6hjT41YvpzXmbhiKFKEExhzx346OiI5z50T68zhb0Fl9r7
dn48axqOdc0ZDtJActXphchln0KcajJN2Nb/6Xb4knr9IgjNcKfO0IoFY/CyPVKWe0cmSvW/kjt+
BZwnfUq5uGgEyFFqDmvXBdJkPKC2T4kUmL7cShi6XahFvZNG64o3BS1AGjpuVzLm7HutUig9aznq
hxBz+r+1rfbFVAD6E7OMLcZssur+H/Hf+vP33j943MBFNopKd74p1SfwibQaC36QJM8Zkc3GePZ/
aIeo5lgCFkuuWbwT275OR4YX5Y6bT9JizTT1SxlPKonOASyJvLyF92gIVKHpIAxoPbmSxghPH/c1
j/KApkwAr7RaHrVSY/7CDBP7k/ZTkszV2Itz+REeX8LhP9wcEV5jMavp+NLAmygFCdRjmbIpSrtt
16cf3n9a1Ml3JdPMkuWPoT1+XimpWiysG1fRVVPyv2Au3oq1UbIv3QPOWbUIU9pmzgn2M1rhXk/A
TT0KlWaeOrapP5sBhJEU8cnOokGYv15L1Et8YqEWH+d1eG2gaJR5H5f9Zg/Nh7BpBpbwaG8sbCD6
eYTZ4v8cNAAOSNyGVDIgx6XUDrni2WCRHo9NIKz04g4DMtbIRZKuXZdXeeKMTmwUlh8x244+4wZn
xr5ZpEwr71Yx7V0xOd5z1ZUNu5boMzJODcsMBB0ugeLwgYGPsrWQV40k4MkK6X3/CRHLytUF8lNl
b/VuOYiIcwZf+l2P8gMZB6Xo56KF+IdcScOqPbpx/1w17u0vOsgKn7b2ezOZl7zDv71pvkpkrjUv
pJurB3HNuNKkvMR8ahMTZ6sJ1K5f3bm/6Y7ixILKVUZg1rGPbtYcrJCB+Cx5nXpqu19G+M+yv/7c
MlvLMBunmB/0JTAkXbluu12VspWqpnGPcXUWOuLZCR5veyK/ppfXopWBxeffuYW0KXM+LTZagucw
CVyNrahLUX9KBX/6nzoseqZY3uea7yRKcrkUkPaNbU1ZjAMw7EUt5gWjSOkTi1sfm25e1ysyw96J
FZD24V20N8QdrHW1Vjlu422pi7uF2jWO6vaeZNaDYwRAuqkSUSEt6lxJEAy6mKJcahBGJvjYIhN4
bcaTkhQW7SAQMW/+j0yCcUeJK+TslptgeDI1QAP1QVUGd26DDsdCNNODIHmM1vRDDIIDKxpTj31q
m+AhtpkfiHG/4wA73TjJin3tmpzqcO+E5RbIli0NK+z0dbISSAEo7LZrAjD6YcXVL+2a/len91+k
1B87kf44rrHMFag8YDTKlVjQoM4xKL5PRJrreyoMch+ZRmHVIIX6w8wf2lm6ik1ft5GjArZ8g1qA
e6YWauPIePiIz4BTYrjk4GPySIw66L3Y76SkBVfmxwX67igosn9NKorzguUqXuC9guSHMo8RRY7E
lhBdrnYlBTlKg+prndV56brGhShiiCtJIZWmIvx8uR0mc2cX/RBO8eUZhNVEiuIGdmot44+TUSoo
ZE3hBD5EWNAodBW3u/hxWyRUqkTDtqVGscsdcY4UVCyrLH/zWwSnfqF7Yk+pEgBIM4bcX6jFEGEB
ycz3iI41sYmg1aFzzOTUxbjaSZNneTlBHpQDaeUN9yMgQQfpOvqDWc2qADavMKMV+PB7NtzkR1iU
GsnRJ4/0i/Nl7OtWZVEwhBKS0F0EnFIAxzq6MVl/q8Af+F6yH4jcukp3k003mrr8Znnh+RabXufa
WDKuRZiZVZTmXad1F7Nqw5hk8S//tJN2wAsgvM068YECPfvPdzUxcLtJo83CZqmciANY/iB1iPi9
elxNPCUH56aCAeCWpt1ofTH7yDAjDVNe+J4JlrxWlHNuVqqpbso5Kg8eHXWcJVS6sxzR8fA3Y9Yi
N9BFes0ZYnO9X6TTM7PdTiq983YSvx0OAKz+UNkdgQJZGRt+JrsZegOf+qF/p5rs/oETkhKKIOIW
LwV7M9yzdxUh1re5jEVhdGwrU6Mry8hlsinNPU9OmlXkgw5BP/rAZ+1083eG11wmbzn3tUdaZ6i8
ZtqbpSNhUU5CO6dMcSzegJqHsacVTxBHEbaiZcYOt75aTLE7iP1JRtEXiz6BknAac57bzHfEtHhS
rkEM9lY76NmhpOlWnak8OT13W9ijWIo0Gq86EYsGEVnxOvkAteuL7j6hoRoUy33RfJ4PHcp8hlNj
+F4flKHsckMcN1HbvghM1m+nM0i9bnIFXLmDhV5kfT50khZXy29QC08nQc6Fkyct9gAYvTb0DMf0
FVfSe0XuXAGylPdR9rMEOI1qMSt+TT46zxAqFcwliy4GYuWblXpt7ycAG+8AtgnUclzaK4JEY5iq
HV+qn+Z7u0aOJakZnXfESoy8Yy6W7QQOUAcdNr37vb85OB29j478d8PmOyMmweQvIT/QhmJLbFtK
ipIxa55v3oLZ8BW1TZe+fKF++IwhNyo3s18VPIRrWaKHouWI1b5OH3EvgL5ZKnlErj52cC7ucNR8
fxCqtSkYKKOjqUFd0V6Edu8sDz0eWVHOVR5LAS7A0QNIKFdXY+1cItkT4hQxeTrVmbOqT8bLgQD0
VTfSlf7oUK116Grg4aDz54CtCQne6HnaMXaMUubsEON5QuQuH3thKEeZ80DjWaO5rC/RGFg785K0
7gNnh9CJW9f5uFE8wU8BeB2Sx0huDxNpH+jnmuJrpgGZoy0dSKCOo2ff1DQqklHZBXhGtlmQyjVk
SysupC41Xcl7NyBaANiE1s+UQjadekdz+l7W2XUzvxgLUCv+cgZN9n7p7hF9BB4LMMN4r8PSHHlg
CVjWZMchZkYBF+Vm1dRkHiLZr8Zp3gL1FvGqYp6cNcHXuJUOYzcz0wLtbQ0DkbQufHBUf61m6qXS
YGptQUIjFqeVM0wAKIC+mX7I8YZzOLh6xVa0kbPnP5aaandq6iXmoxR/Re6l+cAxtBryC6K0C//R
i9CJt5cY/4XbmQNVARfgiqI2muAmKDa1JCgKfxersVktX0Ib+WbyKWRIzI/rJlzIheiH4rMt8IGK
cvr/txXNUn5VWAABSrkacfMjhXy76skuuan9eeMWNRUy0hcQzngRgrnS7T3NoCsSTKY2oZZU6gP7
FzLqCQwCUbXnG1DVhXBbe7VsZz56kkNsEYmtl4utgYnaiuxy87Fbpuc16pNpfQIzM8wbYC0ec+DH
wj7M33Y30RJtAOpguXR6nCNcjuar8U/VE6BX8l48yJukkfAo/f9wzq/uJk6UzL9qWQT4b9L4ky9W
wIDNOk8+7E2OUzWSt6iFbrOcBVCdu8bXBRgMRsKChJopMs3sx1OrQ5Jn+CM28TauRTcrR6V9K25B
oXjonYYCnJpwONSgYadqTgjCfynldoBo4PLCoRbvatSJaY3TFGkjqJT73p3AHrVq1H3KCwoPUPLl
Wd0c90KiL/uJXNxSC4P6zreDyJfpY1ffk0fl7C25AWhae+LHaK3vrFBGXWnVkvEfIBJzfgrHP885
1mwkv8wAeU5vxwMfObIQr51Dh+2UULjmCffQRz5bWZx3H5aj34FHDic98d1UyE8COSsnKZQw3lOw
IqqoV7Y+HfDbvQCfmPiusutlysvTPqSyElSUcbHI++L7WDDM3WI8dSiGJNHg8lKb1YGDie7SgcB9
Cu5GVmD9O7uRyp1xdF960rbl7w3OqOCcrG8fCBeKFuy1oW9wD3bpwzjoPXItUE4sjL8gsmZBfEDu
NxF4H1ViN/S00jtxBeXqMPXqEzwBZBh/LqxCnnK+XK3e4D8TjKTHS6R2/Zfl+JsuH2BBk/Bq1t/Z
zFhxp78QSZCiR+lKaX+Ui07Hy4/M1SLPSGnxHbQr1x6d/dgkMK3uDW0ssxCuKQDL0wyhttye6GSn
NMFjfMtMsEeKvudgvC4HHus5PjfHSQlaQdQuNrtZzzBiQILA4KEMhFzz9vqpbYNSBN8JtQ4xJ1IX
uScSvJJcGelZHmOLac/M/WkmSHwFzQN9gGFxdt7XR5wf0FbveTVav67pEsWgHam4zqVH1QATxfsx
4pQXeU+SLN5+ord0npJ31WorAOdznGbpYiR/NtI3U0Y6PIA57g6vexXNvINvjN9D2FcZchNxN0OD
rIrYTkkPrb+TX1/0PM6RqTM9Zj1ucc0kN7y4M6cC5CUGiaQDbq5kFIZzzdaG715A/YVtrT/KLb52
fF+5uO5++TVuiBbYe+nn/X5/nOmniUCL0EZ5eMI2m9ykG+YjYGNxbETeOCRyylMN2JjX9dfNZQtX
TZXEwOh6TCWc+kHbbFnbqxQWuVUxHKnJopH8G1wzT1aFkYrCjFkQPdAWuobSgXzTVwXCSLB50Q+r
GyKzkqUdm7TAHsU/NZbYDheup4pmwrTroDqV+MntGMah1q5YPEt+MnNyO9Y5s6ZNhVAN3b4OyV1u
h/xG1sHguEF74FIjghoX/em6+ugQbngi9DR+Nv1WFQ54y4dbkb72n5Z42geqmM6xVaf6Psmn7w8O
XWa2DScLAVMxpUxDLZKkDtJ+ZwY5NhP1wVZjY+3h/asZieU9jGtD2x6NXMMME+3lzuGuejnBfnFi
Qmq4UpBF3xT3U3JXULfAPT8SkXGupRtkVnsYopwE1Q72+vdcknXFWrN7I3jqYLMMtu2mX3z2mQF3
Jua5gfMZxMB1NXYck8Hi+RTb+1HKj8Cv2EmR++TJ3ejWNJ82O9vTU6Q/ywqR7AWz6kycpPzjk57M
LgI+1plxbpVDwTZCVPl/hCjsGuHLJ5jDwpDNoQPL7cu6eDbnq6n09TqkQh153Svgn16X9Gn+tEi4
X7rujmZlHry+kctn1jDdNMD1ZqjKWYk0oJXBTka7nuqtyBrWJ0qt7oaOoE0dPO8c48dVCr65yC4u
pmQ7bky06yb080PchpoALvp3LEkPU1+eTZ40zEo8LZI7Xb/z6JxiufuSMQ2+QR/GvEfMvG2Q6Tm2
oz1vFuz9UDD9h2N9xLxrKzhW+ZeJB+9t281+lE5lLc9Y9M6Gp5dLJYC7Xkdc82XeJN4SBMmjl8Ma
M78YItdDnjOvbWrZLutbWQzsZ9KOoJ3ykSVEu+x8anMqngUL9iThJAJj7tFimzoGZcgzu0OMDjGt
gb9IW2xaRnVayD10/Qg7EdKc2gMxFIIn4Ct3NxFSTYclncpH3DJERTr77D/8c1vO03OnDql8AP1L
5o8geiTz8eR9JbEzGX6L9jE3OyZKPnSqASjYHUe/xYK7ybcwuF5D5nRYIoO0w+kDZJBtSpfXKY92
QO+/9o6PFmYub0CqolxI5Tx1KJ2NqqSfmOtwUpK8YvT6Usf0sOt5pWv7c69JgGtyRzp0FeRR3ECd
Ma/h50th8yhm/2pgGU4ZmeMvMyaffDVEQhN8WdWXhJ9jdRQKqd7hkICpIVuGPIDZ2ho4QiPH/3Ji
iYiN7jpZTiK6K8bp980t56O1aykbaauVvvb+xLYbVkw3wq6Yf8cv17dNrbM1U49yAlsWI6yeXz4q
NXP2OHn1jdCC0ukhU+LKBSUvlP+bcHxaBaFBLCa2pR1VHn4z4ZyWKzZTptQ6gN8jxboDUIe/oAGi
8I4GZ5p/L6q1v2w/CuxhVKPr55k0xQufwScO7nlgkyhsluk35GsTHORQ66JOxiRpPuV+ZB7j1dPc
SyLBF1bBCVodvgS4SL95fCzV+lKTys+F1qSFjCbGuUlVhx1dujvL3lAVVAKsK4YXqwhj1B64Rnbb
Ir2IvHcKKhWauO2vPzVtpSqUiuz1i0uIx35uh/bVBb5Zonq3xRGUG5iOeRMUFhL9gEanMHbauf2s
IjcUsrOS7lTGrke/yTKookIOGBZEpOfJc+p9lJa5osUn3d3dheU+y1Oyb8DzHgO+GV4p7Y9r1Asn
UttVYJErGreTfnnQPMJt1fTiyuoH8cIcRvLsIzTe6+j1yGStkBEPkp1PQkcNc+9gEAqYsrL9UUJD
Qu5JVmlFFSD7nod7r2XzzjmWVAvIpxW9NS8YLrlOl13BRH/RWLCbF/yB2cQGyPLsdvsxWXFviKuD
3E/iDOjJjc4iJLJxqE+DeVzk60wgfJV6uOM3b1/W4fCW5cJ54pTwfCLmj73wezEnTt+XDtwEi9Kg
mM9KLzGlGXDiMb4eT34tvr9N8wR5m7D2cQkRqbGQZkXbIR2+ChwM5OBI7TI8dOiThj8N8gOsOUMI
39J6UCuPZejDDDLHtlFA0fq5FRks/wbG2eRmfaGCxailionDxKbCJ9bpmglIpOWuNGxlIBwPdNKC
P/ZOuziurVispz1BsbLrX6qj7KcsUeyr1JtXGqlWGvoZugAWVxWNtQ0YxrAA8fBR3xdxCt/xlSQ0
1TuQq7f8FRVjqyhLKqg/42s13iGe79eAM4hgUGlL7muuRA+Gxpatak1ASg6Q80auirXn2Lm8klk2
cMJhqEq+vrTwUZq/GOBaeda7A2VBUw3xyRY33MQusr5W/zKWhTJcb1gD2QE9rOxg413wf4U/3tuz
YfjCiIeMAGH/90fbnN2zsdIqwgVCh4DjjVVPvTotEk2i2bPDc3UdGG8QeYGR+PJ1Ic0kclhkBbaR
TyiJlTayhTBbVInugYcD9eKoa1xTJSSFo/FSqJPua8ZwvHD0GTZSKG4VkpqYA2/ztViIR/IoygdF
OQY4yEjn8D6WjiA5kRwUWGu2W4G/2hha/wHLRqMqzfWkvCkS6IgXdsLQkinbNFaqgghbmoQc5XxL
YoRDFwSjW0fk3RJxxE4TKN5sM1stB81VNFgRYBCFkS0TzpcW9YA0lW1CKfpmYHplnifmH8O+TaZE
NCN3chBaUJ87dZBeH9ep5CIe7oHzgNRDX7PHYyO9PT8+8FzSaGXwRoFbItXsjyHF2wEnIRiu4FTN
vaN6gIyTOuXVgE7vWGGcTaA81meRtdbR5e8BrvMTE/OYAsc9SoN//LoSbMAB/g0oItbs0/xVEkRL
317/1uJq8286SS/ncR9BzzwX4nlUmQVM3udtnEiXNUY3nwalEHp1j+zXRWC5jRQq4z7/ZBJcJJUG
ikgMpXAwGE3lvuNHNjGH9Eb3Aah4Pabh1R+40X4ifAia3rCeF4dwOBB03TerSD7FIEznk8C5+kfo
vVHeKps33SbI915eATQRKmn9foqYbkAiT81DJZqCLn49leVmes+a9Ag3p5c56Cgwi8nKNrk0va1+
tuUmLJNXInR5LoHoQ4T4ja6fw8H6JiPwOwTUnUqyvZbSXqYHkz4thHi8M9zr9B8SjAwqjeakjjUY
4s1z/DkR/hiYIswMXijv9lv3btZHjvrEZizg9RYMvDQERsMxX27InmI29WVXe81hqxkGp1NwTqu4
pRYhluf564Kv3oGzzXoJKjzaymuy3BFX0TwaLaLjepot9VN8w/0AuFfi63rdQi98hmVviQ7ApSXh
aaG613pYEp7ciZfG3DsJ4XD8bHD/3BzqM97V35J8NWQuCWZdgS2M9+Qtet8Td17GNbyl7dzp5Xm8
28rHrbC/X50jCkGxSeB8767fkGzNB3R3HQRDElxu6bCPOBBucNah+s0icpsQ0s0YURl8aOa0Qlyt
jzgg8SBGp8uZX/7+1mTRrEcxy4zx/dKOfOtUOkSSBlB1JabY2akmTSa+95RlHYMXn75cERNWwzDD
np5eGqvT97mXZiT5iSiE5Bggozwp/iapjPHHo5jrSzqa+fINZKiNqIZ3lJbtBB7Xic6pXqCnrW6m
uHslLqeB4TQzak2vqPXf8gNBUXr2soetzxX88O+89XqflxiY/H0iRs0pD1iyftNB+PFS06PHEBFl
nu5B309/1hd9NJQYJ4gn7IYiZpFMlATz0wk805KjzKLR0INss6ZVZ3FFs2xiTDbT5Rk/inhtrjbe
xOALL33tSnxUGU4Bp/b/jIDL3FlwK3ogyvvkecXr/sOS1Qbj0J7UbRAJeWRfkRK3nFn/KYlN/tVd
7uwxWi/++eCF9aOUGLuggFSEvaB6A8klFPYGjoPv8M5rO7nwuxw6GMF6g+R8+YDjHgd+qmyMAM3h
rCVAQusz7VKd6mmUBFfT/rHnkeDLo6JL9VIQ8L5H+ISmqHEQ5Et7ecrvS2CORNd4kUQCf2JPQLBs
gadWuzqBrQy3bAzCbp8YYxmLaBdkE6ckDUWE707Kjf5SLezlk/8pF33d607Ycap/3D02pJcgdisz
GDKrseMK73XZ5EzCV4e2WUQqOWZD/niqSBKI4vzzGcviNZahJa6U8NlZ1VIuQFdQdbAddC1jhCUQ
NBmjB1tZS44Zgx9b8fZgM/Yo6Xhw6OXC5sDuQwGoFtvDqD+r30aVhSjwHfipGldrvTeUz3ylisw6
5Te9xzW8SixeQru1esDjKtl7ycyl6taO5Wjivbb6taFWApDUlPCAIctkHmgl9xvy2HVH1pJjIrkY
oXcWnPpLy6putqXokHD+QgnmzLN1pJFty0ixu0YyNAykHC3gK7vef9iaHbtAIhWBefhI/odCwFWE
266af95JeW3G5jiJQa7NzbyXh6SzO7mBLAVx7607E1gWK1ax16+w1nsUF0IWM8+gGa09pZ9Oo7SV
LutTl0L80qI0uLWoAve9AVRVLKUNRlL3hJ1g7ozn54pCtVjMgKPHejFCPGPdtwnGISGZmIuOHHgb
RMjFHQnQtprArwj/HtMqV2XyOLdHRobENRNtArDJwfyGN3sTjDVfni/XlFOxwYU3cJnF/tBEtyHb
fK9pz6B7hKE2RbT/7nFqltVq6w3iP/68Ga6QHJW46vb5Y7RVDYy1M/Tlro81QCBGiUNvjsQOJvSf
/iup1QmwqDOddkkJ+au+xNYy6VPuoRTiHWpt3pZAJGXY/c+BrgJr5kcp+MXBH8UZGPTWGhBl3H/S
nwL8JQFyhtnkEMEP65dJNy5ctm2lm/9wQ446czqdd46hzm1I/bMCNRTRJrR7OyQs/GvdevpOxMQS
NSL+XqWR/xOp7DTBS+mCO02Q17OpatgsqMg9YtuqJ5+6Bq/efcgAqr+CD1SeHeOs86qbVPzNOPtI
MXVkwFuZtf/U44MQ+RrEocWZG2J28bQ+wFgILRZJHY2arAia8ZQE/Tq1HyrmiH06nblFQdacVlYK
X2IkXLPu87+9gIWyRW76sgSl2OPTC34PyjKeRLm/O529+kYeU3Z6Ty1p+KIRvbjNqopmpRzeHUHn
v8GAkNtUGR4+V0dcMAawpRkWuWzFIc8qjuUFnkY9S976YPUH+wOLAJ6wYqKnmN7ZF4XeSFTvr9dz
R004XvYhUPE2hdsrhgsKYCeGw70tkXgdAQ8bh/wQO/tC/NpwCyNqDiz/qUbYwbBs+Ie0qEp2mqSi
qJmdf2iUxnvlR4qKa9wPrTghawh8V8OM+OVAvnYgYPhY8AFJuDNe9YJg6+HfKWPADr6gWL31pHAS
csAIxOyv2+Oe5stFTXT/foWg4wkYoyccckjJasTjoQvpOovXVus8u/g8PAl6jYGUGHgCm4zOqXLz
qVuhQplDHi0glTg71NER9NDHt5e1TJhTxRfU5wJKkgdq77LfSwe4HvTKPlBWjma82I/rxmfVFGyL
PNvYB/VfjZNlwD/jaxEEsh3f1P8ar1PP5M+IGdKz9b0Lv/BvAynICz9DjXAo0xdk1PugJiqFrmFA
qLUOMpe9nt7oNlAHwPHMJebZvIN1Nj750VKnKqdAJonsKyk4WW6RS1sDA8dJJKDSjG9RSk4Er3lq
DObRvvAY7GrBxMFnb1NAjAjT8DuPXX2BP6iT7OkMSTI2pI2JMP/no1f5tnXDo46mzo/n9UmipF7E
TL7vLJfP8Toz1hoHxPcwBFMecp1VUWKDH9N23WIunejHw0FLgHn+zP4epg22tY/gSQeMmSTiftqO
EV+VQTDg9zCZ5kCArrsal7tJ5KeFgLJFT1IH0ulhWT0v4WHPmQ2AQ5qE8j5l/ybh5gnMJK1HnWbW
HhG4KQ2s4Yn6FS771AY23XtYiwOoZ7YR/Zfu5+LltBvTY9InauRRtSITvTPyfAhghMQJEix6aAAR
htBm6wnVMoLzZp+A0HEsQsQmV+hAVAocWfz66eqyqJiRl4CiLszAFecCNT1pTCBvqOFtxRGPxa4/
wghq6ZlZj+ak/Y2gsh8o0fl7e3yCVUm3G0lkMIdhsyh0VaEg6ZsRCekGVOm0guiCt9YE9keliz3S
F/rkWx2i9WXl7b7M0Jv4FULJ4lUxyW/07cS4G+yJK8Q1e1uN3DSMtWcU+c8VoF/G5oUOxPDwt/x8
IoqBBhem7luyw2Sn1OMvMCSuIW8sxxhmMuCu6OfKf4QNNDfnh68IP8fkIL5o3iVUFm2GWBFs53am
U+MHKAEnNsPgLXGLDZBFZvZA2UdSuq2BcLcg6DF3l53JZHMVq9/8S3Y/mHbiODkHVm1SzeqlC5dR
L05zV1zf384NJfX09mpvltE/pS+5cPvUKphAth3e/0iUlqVXfqrQzEg7OTDfXar8EZv61ea1CrVO
CsVmtsQ/wUvrZKbEYlEE44xnaDpsBlo/N4OAzamj+O7RB8StAGtSlHes1bIENkZYiCaPdE6uTyrW
FRbuT6aggtmMnnTRaWXtslAL6VS9JFIiQ2VyEQoqEEH2JQrmFWoprROpbJZKiE1ZPRkXEaXrupeg
T/KJgh3zf2VyxRkPi1Q3FPh/lMimLQm1DL8q+4KRg+PYeaDrh7zTvTVe3yN7STSzIWQr5VWTdPsp
NZRtk5fCJf/wG5+zZuK7Fzs9ImxRSffhO319iZytwfbeaheyH4aNK2rSq2zUw02AkktFjUlwXe9r
cLicnIfER7XBtggtR6ZGNqTf7u6tRoWKBJY3O7A9JI7OjNQx4jFwoUr92ceEhAtWCByDz1hmwdRc
fR4hfMvt7MJkf1pHkXvID/fVOMr2Y2GGfbvfyAJQWRziU565LkAq7Gfrd3dZ/XWkejVUeZtccDCO
72LzxMq9GXndzW3iCamo8X6yg4qVADLBjIQefYq1QuAuJAQ4Gfk+zNNhp4NQZsqREBLBXck5FgXZ
Ewtkwn0Z+qe5i2Ac5Wlyt3Qa/N6ELgxW28Ght7wEVIeTg+uW4kbqEkL1ubDTLnw9dwVeLzG8w5tf
58iSRjOFIdY+wNxW4ZNRXlsoeak5e15OaIc/3cWPqpxADKIjVHXiFA22XOdUFJRFSg1IkoTWHLAz
T7Rt2LF66H2sRErdW75mQIoLjMX5tLnr/4/vDJvsZOJTA6gBreFbgClZHsYRdvZJ3lKrD/7kBm6e
+CRA+3H8haoTwj0pv91MBHBJyQ5L6F4rFQbjx7zhT5BHdeutDOl4buXxvf33mXBezbc/r4IFyR0C
Jct8bdt1CYatoO9tsEWNJ5HKalgLOtnICFsT1psxiOolbKVxGyAYm/HLEGnYX8qSmA0R3sQd6ZB1
/SQiMPzAACDg0IhRf9W0qhspKmoDv/r/tupj5YkHLduckWVrt8uLe2R4muhpcynZefgDqMjs8+Mv
oke5U95qCZEOIZdFz9U84PVU5IfFkovpEVVCq7gZciAx0NCbBYi3PGE/AWEy8kttZ77WVgPdUmtb
ydvY/gkW9FVcVPJkX/t0QT5uJF0wpLRBGoJ5eW+B7h8GuIwHTZvW+WTWyWjJrcPEp4M8a60x8Pfj
Aog7gBjgboLdd+0Q8l+szLwPWJMEotDEyNT8qzskfJAl9NklATqHhCB7mKuKttQmO/E4Aange4vd
cmscPjhGfwynbc31+gN/FMJhRIcHnvt2Ov/MiSFdRvBf4R/cZ3yg8WzY7lq3rPB8f5Ambu6Finmg
9j6yHLfiOKBs/571UjgNRPC+A7VGiiCbztf9DJFj09E1TRgB+FNUV1cQq8LTj+DLRGJnHNakLgPq
CH98oBlPX9DM2uuz+tzux7Kkj1y1idWRm0jz2O+2Ciho7iXuCorS2JwOR4w/KzLigxgI4i4euyQb
Ofnw9P0S0JZa/7Va7ZVXtcVihehDqasPWdH1w/PcXcd0hmGa+bMlAQ0UgXSA6YXjWPhCiEX6nakU
5mhC9fHHCYTbsZpgHI1GdkaSR33IKmetjjRDfFIMKu1vR7LX5FvCUUhxW11ZJARLsckOxqm63nn6
O57otMBgAk3Q6gVtINVcyb7o8hTK4ckQfdA4/VPNTAjq3GG4siZnvoYekqOv1CGcC9O+StcHqyms
n+FnTAdEYQ6lU55PsCUEvs3ah1azmLsioujQKgS1yMH5DNmlZlIPV4PAfPY8kSnpikDjGP9AMO4x
YvUB5sPqseyF4o81H6rbJixVuIXiEyuqludM9wGN1cuS13++8AlJTWiQm5ofXr5RcEkGiUFW/+Zo
uZWTX3T+Iw91FGxm1q+0tyTAKwGdyVeUGCeyoyIL0zicE+vI9F8AuzqBWmNeZf4WDenjRgnXHmDD
5N4MOcfGUK8SmTPp8HRuCEdXGg3x850091SOLDHQ357Humjl3gncBFfICRPAWhilbTvhTJLlzM0Q
mBPdtTr9Fg4PSAbOKf6XSY93NoXRy7xp5Qkuu9Na/xpzRNk/3Kq6luZxApEaSisNuxfGEojs6iAA
QU9XNCaXaYVBjK44ZWVzxYkhMCr80udEL5D0j7aS6xjuWPzBl4RDzlaInXgISDb8by2mGj7fmKVi
3L52hZFxNRQZn8KR5ViDvfX5Si9iIJRg/bOhTaxX3FajVubPe71AsSgCXwIYhAUG/FRRM02SxLG8
eFLmg0xjtQWtzI6Hl4OM8/MlKetKvZs/WQQbhs0iJs+2QPGHWkgXINwnm0Zfuv0JjTNlccNuDKMH
GIkTyWiYVi5Oz79eL+Y3Wp7L5kiAMXvfBFLaiIoYAAEWfu4xnTOBxPnxHsT38Hji25QgbtMFbUxO
GKjL2/+fUWLGkI1ys2Fb13vyoM9XDDIKknKEzpsZRQX54S62g6jClziT8wuV5PbwsdW82L3Bx+Gt
ep8IVKvKX1nVnVcyiKoShWcp3K3Zq01vvcv5sRbFAMOFr5JhKB8UdsIInMvnAVcPkW9kPUgDtYDW
UfwJ6Q8+fPqZNRxr9NyfM7bdqtQIdTnVikOEoZ5DkV2PyN9lIb5X5K4x9NkmsdrKCRTQOZawPtX6
LDq41iRiWbpYPcZ9GbA622/6XBpVMdaLYM2/4lN7BluCySzZ0L9Wa1Dc880L6dXm45n8Vf21cXme
Fm+P1vUm6zqPq/mFPUZMZSpUm/r6L7P1aK+Jf8eGnpUfYD4rRQv0GUauZbiZxHsLagn8DLGhpM/A
9UsWm2bWyoycBHw/R/553v2Ecemf8Z/mKBcOggFSygOhURXET2DMx6jP6a/zE3SwJioqXck4wSyJ
8fP+LV16AmPCioSJ8HogtexlAa+szamNemJMzPBy62JnZZam7w4KiV21h4NiJIuiS1+j4CqPmFmW
4irXJCgp1rx0tF0GsOg7YkuglZlzAPxi7DrrivGJbzZVyobnmQO0AHfn70s4Jgh1OpqtYt7kNDzu
lr1T+qFmjI8NZcu5/axSoe7MINoXGhMbgvW5JWXQn9kRcorz1TFjhEgju2UWBHULQZOV/J3oLjGl
cvzhCC58uHlAX5Rli+UhuSPcHbUzjQOw+wmN6cy0HXDsb2rEcsYtOb+26y1bcTzXA0aiqs80WS+p
ga79KkhX/qBnJuEFEjzBIFSvMfZc5Agh3WbdS8zuRokmUYNrLDKe/NnmPq/BvpmKz+CoyGuZlGqx
PT5TMcSKsunn7qZVLV/zrO5/acecJCmGr/w7bO9cy9Wdywti2ebzBJ7QoAs0nQfnzPsDuYFacQG+
OcAQdxTt+oSZBgkpjuHIYt6MNbTElsgYPye5dOe8kiurb2R4ly6bjtVqWcz0DRZ7olZ3RrmTmaII
c/lO773ckfhoxzN90z0fIJGdjBCK0BOoPyduuGwGdXRzVrqt+/RpfHGyg7C2RxW6XvEFOQWrn6b3
De4GEQKEX0pBVG9XHnbS297ddHbIDwsuNkuRgXeRt9J+8UVt1tNnswFbpmzYVr3K0rSu8FkhGYtO
fM19HeBJECLwnD55nxNXclOct0PajdY/h7DX4X2AhNpMRmgklhknp33FI0zeS2hP3XCXkbKVqy5F
ce0SCtpIeJnFpmFcnYW3dYDKtp5eQxl63r4oC0uXriYKXxd04rwoYS7W53aX9En+hyedLTFTfNdx
BL8ImY9Kf1OUHt//6xU+aVNe1CFgt0APC9nqPhKI691sYb1vYxITT1pIyFamvO9TtK/lqx+Ns/R0
h9H+PO0QgUSbbKMZd7/LpE0fPUn0RXl6YtUsthsDARuUA5Ev5Wifv8p/61QPscswoWXV0qrtoWnn
6z9cv8M55k7UogTKfpRPIm40W2emeR41R8gGE25rRaaMk3GYGbu7AHEZQxs7sgmXKY82Fw2T0F4O
Hsu/2wHLbEdkIonXkaDFvVLhWA97ukzXt/WuWZ3OeiYfVrB/cxyCBm/6tNHL6MJVXXgigK2gZlcx
XjuH70crLFQNirAGlWAAKCy+5xcqhr7BsUfZZwmZCJQktjbJ3CDd1BHRvgb0XFrNM4zZGU8VcbgK
z7h18Yu9mhOip/omPeOAJcFYM2b8efCu4EHIWk5woV33BL+I+qsmzmkDfk6dfOOUM4fU8Qfdu4Y3
ySge5/cmesYcaOyBVQJ9x44/H7RD3VT2tghF8XE3qzPcxJnZFuNeq2v6ynho2jLYizDVsWNp7+nL
FWKbce6owwcbk+0F5v8ZBWITK3DCNXyHHg23khDxai4WSCpK0ozn72SMVRmnc6/LArddCcRtJRZE
8k8CbqvPXWb+lvt2cXeWD4iZaKwk0oxWPz9UnvnSjHzoa218V7gvN1kUf0J9j7pmpRGffjL2kTzD
QY2Qrx4MpnWG7/2DlF9iMLi1yaImAE7esEXw5+ol6uBZjweGRgPM+bOkxj/FpeHsEzEHiKaiBQFp
WdCRm27l1t1t6uDlH72bZkeI6Gy05DQpp/wnbSd7yU0Yeot8X2Lev0fYM22h4l6F6C4DaKrhKeJQ
VPELbAKWBNZ+zewRd+RA2ssB/FhOFYBiTQM7H4bC/QcA21CxTOruCdW/E2HSdaNPP7nSoZOZJhE4
ZCknE/ynQbAAfOa13iSD8lRanZAAbV97ANdaLCb7q+eewYCDYm2qqnjDXUHhf5GAmgK2gZUZXdcE
uO2djMhxtssAibMrzsdUSUAkB3TU4/9lbsKnEJxrHxalfGxO1ZOMfA2GyddDpygTTLbIwgddM+oJ
e+sp89wZw2KnZ+mjucsnZGaRleESzlrmC982lPduJW5x87y6XzCw31nNd7q8fiJNF6dI2lemeejo
h5uUHjc83jLxnxPlONH0kst70qX4zv1pcKaz9VfKtuUKKo3GOVSZMiC9iF/CFSJmIy77cSOA0+lr
jrY5Pw+3mD22Iu5faXOs8T+EllfbWSwqVLDSUox4Id+AqIwZfu5pUXVzcAquXh65jbCc7OfLAM5C
UgoasT2MWS6ARgfU8XtFYyiL+mibHMcvnLfyPoZckpzmvMcfzjT4DA1vuW7mKIhDXsfshSsy+8cV
mtVLH234WB/rjcuv57TYK9EAtuhB74iXZ3a4udRwCJZly73K49HxnwW+uAZWA4TGTo4jrj9R5oxE
ZpG8g+zOqBx0v+yJOGi7qxq0MQYKNnFIK2WLC85f+CICiVnKVm7cx/pUnyw0oM72v9NwGDm2GTnt
7VPZztH0/A2/AVKhTDvzIYJdOw3BypmLFoOtnCoa6fiPet/ve3fy3AjKZUw1AdG26RAGH1hpnSbB
PRTM7C1bnasdJpURL5/uKXSn64LbMwdN0nsw7pzbDRh1OcqanlTY2tVhEsKD8bA98L5qPx4w6G4e
F80usav8/wdou/Ch20gfX8mV/JR1L+tO+GBumfhLjtAONX4eXZMHSlW1Rml/6Pc3GYpXXEngfWDr
ni00b8WZetmnGqPmSDYkd1sp0+rLTxgEKTpYSmA8p4M5DFOuFAjRPDD9Qzk4ImDTO+DWMaj1tTUs
BPasS+G+qwXxfknPuqRgAyi2i0071T5aekZxBsrAdGCAjJHDNkawuhvAogYb2Dx93aszprzys5pz
7uUbrli0DT7xfgI+jvII+04ovDjhPE1qiuI4BNWhpD+28koWWqcSH0b1uPHNRr6o6uadVCywAw3g
Bxubafk+fsUDW5OOhR6gt0ma6h2gyosKKgmi1wf4CTiT9S3GMuB0m/mGNGbopIu1EpsodS675BIg
Y8rRLUEgzhGPqh3SiiH/H9Q+sfW7AjmPGheS52X3Jgjzh/pfPcDA4HRUtvOCjsURPyUjOJ3cLTAD
uzgtdg0lxueXzAjfP1fC9hB3x/KCCqP/CUKidFtGWzEKaqa+RYQYwa8cepJgVHBhjcZRa90h65Jk
0V/gW5XhHuTESqVKYsTepymjEKDP9ac8fJp/VfOIk9+pE7OiNHFqvvbW7NwYVnTETZ9NFsBZ364W
QpfsUxtQst8a9OIqJ7bu1d0D5NyZ85czeryCxUEBJfX2wTD7JxgAMYiu4AIIJWD4zx0i5Serpb/P
AgmqikLo5l6PjPIVKdLN99Iz3xETFx/K3m/eF3DTLVzg+lMgChCMlxFMC8S3lPoW2RfB8+YtZzxy
qBrOETGaoDXryD+DIsqnsxitoedBhVrlotqSONE1b9RuIducsqpb9Xw/MTLckOxBlTDInlGUdTGK
45mestrHiEz4jwudlDUN9XD0v9x/9avuyyipwdjf3yb6BGvveBfHvxnNF2eFl/v/1QwtgNW+2FFs
b0nhJPp3QLWJ/TJ1EMPdbi9oL1wRNbr5O2Dzgte5isS0yTi+6s4vNfdjUpyYLy75OmPBuY8zhlnJ
LIyO7mdYEUfQuLT2jeNEvd3V50sulHpItBrcK0wCjlfStlR+SZEZqOz2eL83qqEPn0uhy7hwc9yo
sN9xgPw9wVmNB+me4zUQX7i4aDtPvkWThb00OxKWe8yYG9zAYPd7rHykzU6FKeDLPoNi+RmMwp0G
2kdKBblz55jkpMggDwr6Me7KFct3kT8OX+b969y1h18TUml848pVAam4u9HZBnqw8RnOapSK5ozE
5i0lzll46DZ/ZN6Va5b35DLUZaJ/THCVWJe2UGjBHgYj16c4ViveiAVE6D6X+ZTZ48PbmCd7IbVt
rFgs9WuuylldJg6rs6HlpPZ5k2pyEGUbG9WB5DbdsUdb4OhUwUXpuKWmy7nMRawrNfj9MrUPDJxm
RIPWRmEfo4gBmmWe5sKov5TQCzeUAibD6wslhH1agsZzUu4a4Kf7NDDQsvQ25pNv0rLj3lNxYzRo
zLTJqUaWauishbwwdSwAWdLSOkk+CQP82qD6xhTBy1ul58Wr/oCoE5dU/tkpOkIzXHsDzPpzUCii
d7MqkVJbTzbZmA5K4p4dzWUGZfQa5ddprpwB8gsZn78e9qvefgVvGsqGOS8fkvktZSHFssHKsWYw
7WQwsr+FXCZgBePtneGCRJevo/ei9naTcYTYIwqsrdYcNN3XhMS9hAFrCNlTSS+2NYaIPW0C0ek9
kCgR9f5U8MKYKWg/iHqMlWpEXFnLwfeDNqq3vhRkyngvFUwY39FG4NvqlaLdFKKQsdrwv+Yw03xa
ho6sXte15Ql8yR/tKY81aut/PfaJlj/3jR7Lp3k5oYgZknWGsSNta4XU3Z5eXbv2ub4VKU8ZOCNy
/j7a6UuteoMdpYSn+GabjPgSdEFNzrCZdgeM3SqeO8AJE7mbdO/t7+IZx/NDqGt6mc53VgLvcSuN
jd90WrRUPMazw/+2c+jG5w9nBCgaDnNxKNUs3aixe5L3cA2mtehLcCIPm8IuXegepjsMkZ7SKc6Y
+6gHgzKFvBkK3cDQljhCGbMPKY04Rp4NMVgG6GPYYNHJnFdAJhdQsMXtxWd4beC99X9zIlDZopPg
nRx5mNT49X3zJqogzGCM6FOrkEaj0Hka5nE5qnQ5HZa1iMVZ+WnPsYsRc6uIUCrzXmSOE6AY4wbn
XMuhkKmbcI5CKptKCK0YlqSuWDYFHosjSo9Fv4hsJulmp79PbulPtIpm/vv567Pp8CfTgNcjo+VQ
ODTB0INaQyGHmDpDuIgjjGx+MWhZ40FtBSKYZVXrMpfaclvZL93URCDdlp3n4/SVBciqFRDckUQQ
LVQ1tuIX4/0RhWajcgHO4TzSXyqiggHwxlwGqwQoM/pxKC+C2tkRPyIKbY8ALu3x5KzZp0sDxOCY
MwpumTPhYr0m/2ywLVMEBs/zqksX3WFUcjbnj+oSVUkSbFjNfEjJxYJabUiZeoc5O3h9XmCWfyfW
ps2DBlxXgmYValq0VRgJTXmjvOvRko4MszUKNKCfiV8ZRprMvqG6Fulg2Iy4qtu/s+Z75C31mtWd
6bBJtZaVrkh5oEQfG7OKavhDdM5t3XGUspCw1tWIav5Y4Lb1du94FocBbcjn83tBaXg1wktBVhOE
z2JDRBSZmqjpN4SNg+NXlHwkdrPFz4obnJlWs/xa3RN1zjJD9r/+/SaAAk/WWMkS6PHIAXOinWYn
ISSr8FVH5q28Ol73VEf3Bp+n/DEB2W1gQjZzUjqcEmJRGBSYNJmpgln/CN4X+PjGHQEqshF1cUlY
izYlIwIo1RmU6xjD1N0TnbgmTa227AdERbn47LCVShExI6uQSEVAX+nGoJSPeR3jmsJOVhGZ0Xp0
V/kEXJimZTZrBZIIdyhPEhlS5Qf1bGdPuz6a2lp4WttyfTQVfTj8YgUkId0BguT11mSfpM0OOfhH
+iWaPkQ6xa7wZd15Haj4t9kVDdslerAPkqinfcb94dzrqnkd7dIADSjGOpHR4RrmrlAGDGO61oxR
7534BPOt1eDzmuVHn1ph0lAPq7/MEIv3fV14fV6mXjw5AlLqc6uCAudS2F3IBpKIObBLbKSaikbJ
kNLZf717Bhvse2Lo8WV2KuuEKCN5w/SuQv5EH9Uiy2cZa2oJCWAZxDzjlRczThfDVcjiR/hqTOlg
X66abqjsLAxk/A3QssrIpDWzbCmXQhbCtyzrzVcCbp3i7++7nVSDdN+BwNE5tToIXTatD3eCGoHe
4HJGjkyFdfQFrPXmFk5eo6jKB2wZ9u9xikgh0burPqCfgOc71McMOn7nj28xu2hZ9mzYox7CuS87
f70GrRjZIzykOv40R6ACJUHrwPqHldhB/9Ow60WnM7RJ4ZHT2zwPAZsespGM1XfugLEQ/0JozFy6
axX88DvHgUQc/DBdsAnYmK+Cbu7O/2EAMLuzSaqWfDrDp0csSABz+fKE0IEUZWKfKGcCTvtuD8nd
/k5iv6h2C7DcTeK1I8raMwIn9+z61WA3bFvBBfPsDm7xddcYuKEs/YeK9tmqiKDPotd5KtNE0HjR
hFv/jpqu7CQZgwbIi0p9ENK/9mBKVfrpscYz0L2JINzBn0A1h82/410O+MAnKh7CS7TJQ57naqlg
IrxWLlFULaxYnayXUWtk9lm3gaq3lmrB9Prk6LDUKzsGfa6tjoqJlaPeQRjtJ4yaCsdJMSk5M8Hd
aBVMdY6H3MpLwr0uBK27IN2nFeOX3Jw2tawbgEuwnNska40YgSfIf+/Iw1qnMuD1HAD3ISnU0nNV
m6bKpjN3G1xwOyExaCFJrtaXWnJURT2w3z519VIEXLB94PjjJ6tdkc7nteDsIXND2lFeAAVmg260
q5JqClUNrWmaz2rZBmtIneTfgPzBBAcWV0zWy9qZqx4SlTL21kpIxGgpiTx9v3BuU8c67Q1pXHYw
1EO72V6Mq26TfcBFc2r9xkZY6AWSAlnlI+EmRELl4JrScto0Mo0f2dYpd/o1wAbDcUUGfdGW/R5o
Hzdt+WHKjo6xK+VAsMwTuhjC/euhwcVhdu3xLo/np6m+WQFcLk9kD3kFPrLVA2BStMlYCFIGWxxW
lr5R61qJT5yBlKfixMhfdGbVQTrTmnTHFv7AdT412uE5EaCUFw0wuhX7aFRr6zeinn4Z2Nj4Ty1c
rVuL4U6hTMM5dWgrvq3p8aipPpDIVvOZ7NETFcaPOwsNUuBBVVWn7mtF5/t/ual3/8MFNcMSynfy
arT6E+4rjHBAeMSmuu84ppHNlSehPyH/dMligFXuAH7tiU8svZ8szIHFjsuSyLTc1ZztXp2DOZHU
il4NVoDQWD6qloasTzHdQ91sMbltj8BN0kNHcoLYZLCueVVkAoxLnv9ha0Yk3po1Y6JagJxKr4wG
7hHXnygly8G06+utNls3erpegVxaK30jH6Tt72OA50zFPWfJikBBYifI4tTgq7bjG+a/fl/aoVMc
jQYw9LgAzK0XrLCfs/Mau3FIAQ/sqhMtXfqg5pFNmphpBBMBRlprQPqbt/3IK3MLu9Pcm12MFuIM
ck9wc7ASUwKxeefYusYx5CEG7WdQjQtQQnOfINa7b9BdzeRbSSLFJGjSYA4udY9661YY6FgpeMcz
ZVn5sc86bszT6NNTMrKebFScmawR6XF8Z5zR3xgAzZf7wUixTBd8E+JM1BXdjjzkjsO+VJydKNZ2
0j42hXhMct47y9GEV+S8bA18hAFvPk/Rksre7Zu4uzS4d29D8/JqipaYBk/L+YJjmd0xYAAT5d56
oPXFpz6CyIgz2ZcpF1TKg50xxbLGFF3US5AYYbigo8QYlpJ2SfsCBEPTg3XaMFc42ORjRXK6GiS9
0XoFMmv8gsPZuugl7fWuS5XQdWQbTTZImGyk1QTUGW4JipBarUikpS18Luvkx01Epq3pQMhbznfu
sNr+FokrbtTop/f5JDhN+Mdzr7PW8h0zI3R5wGEMGk7a1celoC8PKjEWjK72fbBuoV8BRs2kg9T1
RGwVpQhRo/pOlXN/iYhTeqyrxFoPqq0lBlDfPd2Ngc85ifjNwVMq+sx+CgalgoK79vWVcIg1qnP9
+7jy63AZSCiKVu6F7riKc4v7u+ijjsvsYMRtdM8M3N1MD00zCOW2QA8OHLSfmn8+9eBJVkHriYTA
SnyKpjCLqOWNFvP8wZcWmHj6ruEcCw/MiPv6WfgS7GFt3RTEQ9fuVD5FqEVHfuQS41K2XzzZRfa4
/mqeXBrPbQ74z8asKnordbq8g7tC4xh9E3ID1Puno1n789u3nwj4Y0T/0lg4NFygtu7/OJA2nFcT
qWHSbLVaXvq7NFXiee4f2JgPeUgVj6tjsiFKtCwRRxrivzhoJGFeNziIpaEKqG+XaE8K4E25ecXo
zbALo0WO2LS5Fk9sj9v9eTB+RZ9Jt70kQOt3P/QtTb4U7K9OXCQG40GAkUqzO5k6ZPgDmPZRaFYA
6qECQhYq0ZunIfQno3vAXKnj+/tP6xH15P/3gkXYJe17fbQHMy+2eWEXeu5epFt7hUhRRFqKlvGW
ht2mvIcmN1OQUHbRppwqeojIxNjoxw5S3rtxOhvQ7rkJY+Swd3DvbmjQl9T26+SJ89nqdVj66dRq
UeNCLv7CK6VjFX6TSE1sPS4NzL2/TPjuMQwJOmRQNQkP6DTgXxqxPJQiDuz7D6SEY0KS6diPz+ps
zb7+WTeKhUp2kB4SQOYA5Ubr9WJrtdjNuTUyp9Wd533JIPrW2hljiUgh8rmP90Qna98sI//fzdHX
Pp2z0AqUN6WtsaZy/2BghM3sJ7a9HlJiFZw+qEbo15dNv+u2jKhVs2y8acMkTQFtdB5jMeydH/OA
dXk5coiuwQfdjzMVWRf7ew5/Bsrs5wP1lndEm2ZqPX1YLEzXaKK4yfpoI+PhF7ICEl+ycsv+6kSX
64t5pIuZkz23zGqpzhjWw+bo6E1Y40H1V2o+AoK20oEpHWAVRXaW3SCY58ebwRe+e+i979cmHL2X
w3AkTUheU4ftTXpfPzB0OKty9Eh2VT+6IyywG8oQWsUMVRZ7n5T1HtHdW8XSBvI8QrXcPsEzSwpc
NcklAcxd7jl5ZtlYqXzVnUOchqpjeClueyJUQrmP+JcXZJcrzW7u8rzFJzdZIZDGibp3hnFnTmMO
7gdjmoXaSdFslzLZYTghviKNFGD40+PjqkyqwvOJv2u1yPI2zkFnAo/dCussO7pNEizz2b5CSs8G
gzD6G5k84WuOUAl8oLiy4f7uc8DNP2uQ7lymX5/nHpFWZ1HVpKgfOhgK/nmtQP2+CB9W2l2+pCvw
PCZNOh2LMZDCamPsy+XqN5E7PdQCmtxonH3M8V842ox0kEwmR91U7BgkVQ+6THZJIRQjKDQmTES5
Oy3r1hXGNLn0BBfEmKStHOlcIW+heH1LU9sxKsaw/0ckEKnfx4VTW3BCMTICjgXYoFcz8IWDTFV+
B+VJhT+sAgw6aADTs3Tsg3kK6OToxMhlP2eape+SNOb/oGsxVzfGiqc7GwJSDQ5SdBDHBzeyC8/Q
oLPBSOzBLg+9Vi8JtpuUMyKKy6KwF35324ObdJzRwevjzDInmUAOeU0R90CnbjPgkqftdj8+lIRL
NZyOgD4HShWiHY2eDDF2VGvveciSaBFp6RBaluWMAqHPhtVF8HJWysLAHobnKi3xWGq2zJAMTlkH
MdlevIUGu/negNZyM6zNrc+t0zeGbBIFOzYb/gGsOY2+GmY/uhjgMJttiFfBv0DCgKeYbdZZ3DGv
2WuZnF0/D85Os6BTd8SA661zLwsedQIg7N2yPpLejrybpQFdNW0KcNOiyPfiE+yNmdlHqEAc5oJ9
esdmAJ8q6d7cfbdgzwSxw0AWemlzmk1Qjs0Lt6Q6DucPpaYVaxBc58WJof4+QUj+aGV42Uq6sQJs
+7Hl76tL4DxEeo/KogHa1A72fi/kQvrRQcdJxo7cGYXV6TnuJxRbKKwIPvm/nN4BMuspiHUr9JSm
AJuMXx7uGtMBkuHQwCyMUlSnNp6+9iCBBgc07s46kdHpUaaItExKLjnWG4Fej5j5U8Xyre6g9xc6
bZOyqbVy4DEqGh7/VqSiyrh3aAem6Jwa2FYJck9HNrgJ55/cg01baEVdlhZ2tg06z/LNMfFquFeM
gpoPLEKk5mNIA8/2p/0+thnIfdLix5swv1//N0XYAyQGtAI4mIzw7ojLvzJCxau4m2J4oQER49WM
0kbnQUUeqoqqTG1q50+VGjXlA3TAaraWKdroOggEmFhBtGNFBgXButcJGit0RUA2kP4InM/SdfPS
Ev60ALK2T/aPHPA6cXuHdHuAtqY6JJauGd8YZAtCGMuo/ZOYBdjO1L9w/+VQPuyBQL8WimA+J8hm
hgpuqibf7czCkr47hm6DMnvhZsrDTcPM/JYWhTW+tKmNd9JFmlFs2hXtbSMdLb3HKy3V0yWpNagH
rEwIAiOS2LXviakI6M8Ul8YwdFwbGrDnYlJucJqh23ljP6RwaJTdYb0mrLj8H5BUgx8FunT9Q60S
jz1yBrHjBS7mnTxsPWlTJ764/U5LBZCbqnCvYFHhrXti96HSPgYLSLVwrznWnl2XULsk33a7R+tH
kR4Vwh+JHfg5rhejh1It7B9FMRr3l/Ge4P+xlNyKEeJftYp7JiewtBgMtH+MoY35WAeciUHHmEz2
8Wvh7BlsJ6vdA6XfiIheX9tE4JFZMtQ0/8yWFB3IgVGvw+Ax8clUO5r3jApKLk7Um0DzJs/gkHtx
waGmRs0/qypr7Gd6Mo0XlUwUFipLhJdZfsqwFl9t+Gk9vRdQjt+TKfqUKxPjb7o3OSPBToR73vHD
Dr+PtpYTOZdOad9Nwj0ho9I5DaGfX183W8K1ZwBuRLb0Ub4HuBu/9pTyIIzwNbHCOQ+Wg2ll8Jo/
h8QwJWcTJSSuxqoaTJON7gBlnHhvO0uZldTnPIf3ntvYREWq9YqZz2IDbfmkkKQ1YjMcBKaKaHdu
oxMWYGMVxTwDvn1oOukKVisIuqtk8p96nGWIsqgGLY9nCEFoWe1fl5Iu1cgVBn0A6Irz3zV1GqXg
fWWS5CeXpjxBxbz4nGPaNEEGT7Mzrn2IpyfbeAZYnryX6DQoEHIo0TsdWAUZYAomHNcGIk79Jnbs
bKgT/plpw0oE9BTO/c5QWkLzQgBNSlXB47OCGIoe71ceRNvbp/zFCa3JRW4SUb9A2/nPtqND1dtk
1enxrJZXDjL2JKIEFPOgy+lUgdJSMx/N6m5JhwXtOTsNDDUB1n8ZjsrQN9wmzH1t5tm5zapo2FXq
KAuS0treyeraUznkH+MLYf9DnQiInp6PavAapmXIpjEXy/lHMdhUZ/kbzJnlwE7vG4Zslj453oxG
OptN75M43ciLr54FQycix1oYTleNaUPD0GnO/xqhzERdcrrvLpH/Yt+Rb4io6TmZIb4H3E7gfcaG
UWC/rAg3hZkbyzYjage+EUHL1o5xVBlhXO2yh6gupB64Gwuf+JKjNNGpALbZHE/mGDtJGDlbq53O
NM+23vjDgWG7hogi5PPSVG2iGOI8EWkYkfXotLlqWI9a0PsdAWJ9/kNGGbQOPt+tISUVhBmJn8W8
eDzPYRRbwPw9ykLfa/gFKf3/ZKUP1TMRZ7ERgFOjXZXTLqSkfKui2Hp1SinbYoYclcJQmwIj6i0q
QyNx27Vc6kvu5VBerK9h6o4t6XJEYs7YHuNUYmVSDXMZ2rzahrxFREhyWQqRGhgUanGUoKSuo8+f
FoUXOs5AR+jhzUQkKOefoMov06l+Qw9LSse8s6qpPNbOYQHcIkfORMUyOhqui4vSERzXbvAPAkBk
NDy8YKKbaNV+kz3/hJx62u5kMQ5FdNJo6DE1rwegWOZH37bxn1FaI/0EHZ3NzZCPLdT+fjLL9Z0Z
alQ6WOyxY+0TETMBsck8YrG3WWPLc8ZCiqkxza91ynCO88gXsziPRzaIJNeQnwwsSBa6uO1EGDFB
/NPgngjz3b4xlcCgVJ2MCcK7DxLr0ttkHYMoDZ+FkqKfyiKuGMt95aHd/a2wVMZcvWF6utI1k4kJ
ghYhRsTtS7tzRYn51U9SQU0HrHvU3ufrpjnLSt/2RQFiAHIdIGVGNUJMbBHMqLbD1qCegnk9bhSH
kidOlWyXdQwkI4DYxhEq5QU8CciuVD160QRVpEWCJ63LPi7dbFMAhi1sRf3/OIt4upp66FDL4RQk
AAD04fi0bRY76kpVKy/4Uhp4OOHKydB1WwyrPJqwIeXIfqLE/DrSyATTKPixTaNMS4ZgWCEk1Sfr
+G/UfKP7tLhunXmImyDJeWKHqc2XYisSKk8M/a+X6/OLaSlzGyybDtHtGiphPriO5EHhAOg9Xas6
m1KmjBcUij/BfMXzE7CvglnixyjP/hgOxW0QCnNVSQyGGESDErzl0Gj4m/4K4miGMKPkLwkTfr+a
S92DF76Urnxl/CXbCN5CWMnkLwtcivrYmAgOELd7EUxWfhni6TabsrT8TA3GtBsVLLezkknMzgAF
Mu6+fxPqSw8EwDxAppgaVsJkkfmYPOLaYhhqqg/BVMu6Kzh7NWPf+e1BnKWwvt+KxUpzkL60dVJZ
nw6Cy8qtvYhdTgEqAzbIkW7JCToYg71IuUeI3I9hL1ecGsaW69troDdT+xGWdJr4k9hw9Zw7uIrT
i9GVLbSzoQO6OWxgDRidOazpDy+hT7+afvgO1yRZRKg8STaUOUOKDrk/5mx/neFMQy4tcw3Crl2j
FvA3f/dMghAiznjFYzIBJYrpDwby77YHZxX6+bCE1Lr15iH4yt16Qbnee4ZYu0/HZ6o+Ym6mejJO
9PGRt8gUhjAfWtbzphnOWL+ThiV8QjTxp1XSsDYX1Nj4NuNDBKm/OIWzTQXCHerGE/ksqrXKlCBr
VBzjYHQsOClgrCHwHuBPGGqaOvZLgiMyBAh5sEzfTErnIuReyGIPFZGaaWcGAt+dggxPhyqNzhGY
NyDSgL5BXv1QN1ThH0CGhZv6FxOJmGeiKT4KrcObpA1PCR95HpAlIY08LTFvKB1qRMM2RCXqccD/
CV2dKOLZ2USpl8qOov3k97ngBE6lQ3qlHm3T2rZ0izp738wvcTnL7guivAcqoqr2tnj+KakRtqkR
HXm8idd56M5Y2pDr9XULzi490UQEW8hDnRPCcDIjUtGBDgvUelJ76BSYlUCmgNhe/9WFN0XAcG1F
ApgVTZpcCI4fLJLED5NqpICact9ZmYGsbsUxDoSr53bIyn34Kab6FOsJtn9fMDiL6N4xYns6t9d9
SuuSGZutIN0vx7Sj3jTxpmJM8DoBfw7DVpj3zfdVrlk1RRWCAu1IaWM6kzSrXy8QDXPiZeJdmS54
cbGQ0URHHiPDUD4qiANqcFDkEowluGgaZ1Gy056VCLUgILQ+TsIAPHQLBtq/S8uLY6ryxZ4T/ro+
sJsnDv/k77VJazEt/7GTtP7CwCPtEVio7oFi7fQKt+zkXL4ucUROPW7goDGrvwUnluwnr/JQj5Q9
SKiQ32++5BUddbtVVxcMqVuP+oWf+wkycuIMbFH1EdugfqTXkDr2phgvSBAnVXChca0bMZ0OftOa
cZMXKKjcHReoZ22Rf1y66eXwttxRVpSJXVGOgBFL+n3wq04QiNvrvxvdgO+pTFyd6t6KKY/uuMA/
tQhSW/daQTjMR2KmHQDxzXXEkwntpl4kB3SjvH9yoEXMrBCVLttOuW9d43v5NhuOXFALwH6g0Uob
m8uj62UFQjXsF/qKibkFM21BhOftVaraS/cj6i9YF4h2AUNqPqTWcutgT2I7CPBSYhd72aZMd1uF
pGFtlQ+GXSH5J3AA4gLR0pZsbwvRfsjci0tEmHoktkS8AL3ODrly2bGza2QGnLrRvcLPm7iAGMoe
4ERWrmkFmXHu552FVuvAtIdlUgzy
`protect end_protected

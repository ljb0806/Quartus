-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fnEUx32KJakGC6GAHo7B51pW2TW1bjllsEpJikj5cshaBCgWgrhadDc1FySEuEcepB3PzFaA6wMH
sU4qfBQzRhDvMqxRSyK0bMHvKzgW/xTYmJmlm0rbGMY92RpfJQcRS/JTf+tj1KPsuqrBSsqVR45f
i174dLF436WHhKOmXscsWJ2gCAfFFmhNo69j6HDTSWUai+PHQcQKR6YsgSn7i9gfpLzjq43PSe0Z
Re4VR6krdvXpJIOirCUK0zFytlgpaBoXP8wxiSaFHEwY2TgNZmNDqrmt5YPchmEduSlTdnS6KS7E
wEg/vzLnEdZKL2cBWRGd1OW7YXvIhzlybpgkmQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 72832)
`protect data_block
WZGZdO4Yf96f83JOyHU/2NGAaUgiLYNnausZnde/56k6eNDVi2t63HC41HceqmIhxktnlKSHGwTv
/uPAoCSODh+0TtXL4aAtguo8mnFr8Mpk1jaH63uIBdj5Tlgt5xMpObPFYBO3gkRkdYG5DrzfnVWF
2Y2Ozyluvr8OiLDhS6CYiKVv4qboDm3n03Rt/xDEqPJ6bAj/6IKWupOIAmgq3j/SwQErKsOIRaKr
CGYZZpi8UN06vq2CFuLCGHB7ucHfBtdJmiqyjjST7YdYoTazX2Go8ZnHlLKTYT73SSEW81siaEJE
Dyasl75MSuX5rFWjrXa7QXYtvFlqFqv+f9vYRTmqsW3aurrJOR+tgwTIL37pUwh8pyZBcRUdrsgB
7V2jarghwBNAKTMIZENVqFZ7ufglZ3kKXdoGAxwwx7J5AGiArm8PTiv9Jl3RgjQW3Plb+5DWntwq
ndmD5qVoULUC2PGCqdyu87HCO9cckJIGyK9HbF4NNxXIq0ze4BeQ/qjZ0zWYTTK42yj3xoqOc9mD
ZcSA7QZqJ24gcmG+IxdvOkTf2BzmFH0ozvko5YMBE8s2BDrKGjazKip6g70GOlLFFwPfFE55OW7T
0hMgervvVU/ShBA5F1JDGALpoqMNHQI/nkNEf58J4pPk+nwz2yF4iNwwTMGjqhEpBdpQcWpge/1O
Qak2/16XF5KURnip8tLzyQcyPPojwlcmdpJME1iO2iwRGL4LMK5h/PseteYhdD0ldtwbVGC35zLH
lODTLOPSE3s5TJIxaln/clfo6nSNvsmhcVFMaEDdWYwGv03/dRUyMqK3LtZo91vCJPdg/5KHJeep
7J56xR/1iAjsz9zl3PnyI/qjw+hdhbxFgqI92N5H+HTBag9riC/V9Yb7xLpRMIk8kTA6l4RVwLdZ
kkTt6ib8wUIridcgWshfIvnMD9BKHxoyKgD3QKNAAfF4Egqtf2UvK2Zyte9mnRGIVjl/aTb8tftJ
76U94BrETHpB/mY4YL1bR6FvSbN8qlaoiMhRasQnrmP+Ni7q2zAViTHRIzOiE8eRMcIyvU/Vndq+
tyjQOMXLxKPWoGWYgiSrigGLalRDnSAc5zcth13QcBAVFKN6lswDcl7RAF4p51Igv/VVCfv9volG
YQ4YdQPsdjVSnAKlfXJBBL/PFC4l2AYLS1UYG/TGpw1UuSAgUAPlTCxUpoHm29OoatOQ8smpHYPv
tIfGOFfZl79g6fFIhBJwNb+AzRBNyIhq3ZP2Qr8W9bQ7t1xr54WnqRJXM+Q+9ZOdkr5Ine4snzgu
N/4KwtLnc7HozSmc0BYQkHT70zl2vp4QRDU4DjJHTvSLlKn/tAyzCmoUB/CfGUO2gwB8EJYlDACn
IbEmtd1mVyFZTLepHsH84Ho/rVXZnr6ZBm24V5UIQ5OHA5KXdnw9awpszfit2g7S+f0Au4vPRe16
ZLX6rXnUWGQVymMEa67cng2mdvpC3BIMciyxUwFkmtawO+aGB+psukHxnR0x/SLQWFCj/h2EmLEV
19NILS9KQ5BmmVKuU+wMhuwKX2KmhyCOFo05qnE6dqRWWWeJ4tOyeDY/W0P4kBF2FLrsT4FGY0IF
b9TzkKcZVAbLAxAn623aQ28z2vM5C/d+9qE2U47DCgl7SUW6DjnONwlgkWnS1KlY1zvL/PL12+eZ
tXQIBLYJHFh88xPVDmr9yjxdiDK+5pRnLRIm32DFvJLCM9dnbyD48w16WysDEEn2uojoRi7NXwv/
/4fzAn6o1SY6qhTTKXZBrtDaILZ63OsMmV31nWF/4pIP8H7eN39rpS+MNbS3WSDX0c5KVxEb9AST
tX5Eyl/1iPZzQ48GsWFk3BzcS9/MyR3Vkn23EkS7Gdvm54n0spigWuz9DxGPTO2USF9Sjqm3E+Km
nssaW5uthdS5MFjTaVzz+ObLiNB10EC2B4zTSWEXfyeITL62WKITdC+x14Q0RTNNypXEtFKhN+PO
LSvT4kWiTififuD0UmuSXDOnSlQlpZUfKBIyFWCb4sjNLvJK3rWwyzSWm/qNUdJkTpbZoXI/56F0
5V30jK65y9v5H+n4LiAEm7ETwlNY54r6aY2p9EsHoIgZELVxP7+Ubrv9eqFPpqOLV71pndHU+JGV
rdfHkx1+/4KPNogJG1R26t6+uLUIlJDLEZk/ltCyt2m39E39mODgFheQQTUtuontQpYWTMr2EKTd
NsvEjlVOl/9zMEzLIO5cWiP7ajDCy6IY6kARIEqhvbO1nFgAHlGXoyR8UkEApdkP3p0PAGPZYib+
fCFblaIBHjdK/EXQU+8kyYRmfl61tPfS51r4F3P/G3Z4l6FP16gBLBQB+uuxebntUiwQvXHqIsFc
SCf4SD9F8RuA9qJg6RrPt8emUnngVr92vIOTEj2LY+SY6AiCwuCtLbTdpzOZREaAW3Vu3860+6Yn
nZHLXr/FwhU6ktszfOkQMrzz/k4NbEDrJ2kBD6N1MtO4MBQJd+DXizM7bkyYpKaSnpRxoEX720ho
zXIN8Byc6TcTlKAiilQOLxvstfwwZ1AQjdTNVfUbfwtzdQ7b4QzvHgtsYEfudy9h3faT5nDRe5sg
2+iN4F0ACVd3CysDGPXAez76DCBtGcNSFsA0vTgDxTVI3ZDhntLXjxkmC9mlwoVHvterKzeA9xFS
Xd7hXcBkLbZghpLrSMJzjbwenl9gCQMcPJOh9YxdBmzHIwvBqqIOWenq3s3ZCsKlIdDs4DKdu27A
TUCX1CT7uTLwKRWp9W+fwN3q3Y347ltmKXdUXMx13mdMQkiDPCot3n2tqYUZmq2kkPIqUiQSKqGx
aBZFQSNWZoxkkwEv16dr5RI8OIybEgsEbi5+uf+KuTW7di9k01b3IDDobuF7rcYcSCp5Y5CxOKiL
HCFGhlsip2GzF0PzhVwxsw9vcOTBVcW+u1DO34mL7FVFvXWAZusqQ0rqMJImwdlWnbKuWtPTcbhk
9SlKxs3IttlgyvDsuxpK/nfSLYwVhSEdmpEgg2Lcv8559RWeEE9g2GF5ZzyawXnRqclYe4tyjrVE
i5ybm3UVQBt0DP4HvSlCUmAwXKTqok+KhJgFHA+5Z4uCuIu7sDspQYRyaAzXcYrJxFstaEXeN46A
zipGbDMT3MJTZc+JUqREWSxnjUtWPrZhlorfkPFZnHYYm04yyxjWRbZEX8BojTXFmOeFf6R6G3L5
0IF/hB0K7V0i6Pyx3PK27VouqmYluY+E8xmg1XRAgTIulLiBrWqMS9tx3Z9GuOCiAII1Evenf7hw
r+Le9Xf5uaKPgvvxbk3v3dYnbjuBcdyEy/mtc2N040Wd8WaXGTinxCsCcbrVz7jkPeim0Vk5et53
QipK00U/4CKpwVNw1YeB6epWE6ULg0mEh3cPNm4W9ZSGPwtOGPTjcw1YeaMCI9Erm4YcKc96HPHQ
yyo6G9/whtUOe5h3Oxe5ql9JC+jMYVFREr2IZKxDwOe36rEtz2HLlEss2GKbFiYKedypDSb0xWWR
ovl9wkj53Ky8NIyL4oPyXYFb2yVb4UOdncWbN4ZNgvFG+bhIpHsCIl/lITded1X/aYEXsPMZW7Xf
3jROD6GoGIPnMPk3ECkM8ohv9+jjjTbOEv5koLEtuxeY383pO8w8DFGJbRlyx347EOFDY+iuRHQb
8txe7ER4YhVYWfR+SKZY4f1BYzkRVnAGiWyJiA5J127gQ6XuxvdaOgDJBnLGyA7ragpadlfysPQl
7J7t02XqUR3rr2h5XlbFsN4D4HatQvRCGZzj9OaM3jF77lWV/Orf7M+MMR4VGOcFErWH6uj5SYCe
8KXrFD15hEYkhNSRMtiKse4XBSiYTxEnS5CClaQbpsyU03CGNXs9/3XkiDcmDurSg1BWElHvPsVo
mT2FYH/SotF8a89r9opF4PQHBbH9kfnC8s17ezVvn3hpwd/qt93mbDaTIAYfSQ3u53nXqLZsfnAP
OE4NwdYRbV+y74E+FFuLuvBJm4EmOiqT+5giYrrd8tSHDFF2QS3obJMTCJIVQmm1HS0N3Y4MjEj2
XtHj2ikpKxJc1MifYk5ElZauHOfjJev+iTZ6l1XeX3RQ0DrXrDGLVJLAzpYbWwJesxvjv20smpAT
6qVUbIUi0osWVyZLHMTY6DV6uCH06HAPHKAhLlsbeAwtss4KZbKHCzPZdl4UFEJQn3vvjeD3OE3j
1iYj1KEf/ZulzvlVNMwjhNlRMsXktSjGn5sFRfKeyWz+GCZKpy/IjyyYUnG08/R69w/MnmYYFxRi
UdISIaKiLihjJYOwQPU3pfsk8+4KVQ1sNN6jj4QleBbe7Gy0BTwYI1D841LCI9W0b5AKQhQ6257F
EIOt++ihEesjQ0TVVsA+z3dLkt5bDz92RHVeZ8359r4SeysB9gUw2gLJro/YF517xHQHo5ayKvK3
FwSaH9BIT16pcC8hW2xYyHhXS7WFu9pPCtR86nfOuZ8wIJIMgfuXyJedoR6wqL6zmyIgiqTCSpDY
bYcE9HBkxYaC4QjvOzVvr7RIODvn4bXcmjnhH0HE8asUNd86BuEgROXNSJAKWXF1TanhBmo3jXB9
4jOh8QEGl1lKziF9K2u0YobEjt0wONpdGwtFhtUY9LU8YFcR6YWNf8PG/0+vPYMaCRRWUdZjxKBB
9yBAa7l5m1S59sJpcxouuCuy1QJxWaJYktmUbXnMfhbf8DSWfBlh04ZnJZsW7/po4gLSr9JKP9so
zmk/4+PjkIzpWyUd8DJQFBmlTSfcKk6jZc/zXoGEiIlDKVOPDXrSoM6Q/hvdgFmOoN0u4PMdgTmT
bdQf3lsw6lYrHXRxFaxVpHALLYQkXoksx4wEOePU1Z1oCzz9tX0OTNtOdkQ+4ra4XMMBKejETkuh
XFnV2VY6DcQiCd1OJAjhhzu/q/Ys7Rk4Fq+Z5MsDDzrAxptvqFDE2h9/HEtlCHO2biScGVFsC4lm
Z5q7/zV3LUbIYl1YMl3FQTFv7kumo7sV3/dVxamuy9V4C+fbmR7rZpHF12ciOrfTlriVUnL2zc1I
+ounDLEf5HR6yKH+U7KmX/SIWrbc65WVIWpRCOgwHQg8JP/lBPvIhpvR0UpFTCNQuI+G4+HL7MAr
eGbIgzn9ckOeOQthj3RVP/0G6Xm7BbAhYnFPBmQZF6IRzdjhBC/CX4D8PG9og04jTdvJ57ZrsUGp
FIzV34OVZN3ZyeJ3H0yAylBhO5h2fWv0iFpQcZW5EP7YfxecUtzHUfIPEvvISr1zbTrHoYpjqwgo
Cu8pNUIwK5sRnU4dIxBIR5wOkfw5h1+my858l2EwdedYRtbEk7mvPsA/rfH9ApPaI7I0lI8p5omj
NE7q1MIi2I2u2pSFFBQ+E2tsBoU/mbIo8/xwJC9GU4L19jJIs0kjdARst1uIDIsnnJBsab+/xOVS
UdeuPNug4s614y4P55yqQ/r+81vJ6FQyD6Sz//H3+8+c78gz2OTM8/oBq3vWiBjwT54/LFmIePKK
EFvRPTV+ynw6Bjt3aNdfu+PepfE6r3XpLyccauHKydtRqFFMGYvmveV46l+IYVCJSxAcbyB92w/d
wT4+KCeYjHgquJky1IKs8NHBPisnsLLRI/nAjdoDBK/QutR23l030C1mwFTJ+yJyE1ESTEjdWxiU
WNMPlgBsgHQvs29d25OI9748HMY1zvksR3gDnIcCY9/iGWqK4p5iH+vAenL6bo3Zy9rc4BJ1gpeG
RmkfLygFVOmYfCZXYpxAHfHPY1U3jeHkSrQBtFTSXhp09cAiTTB2oj5LjGLB4jqH64NyxBvAQJ4k
wqWn0eDJD7JG3n6KbqbmltcXp46uaH53ClKrTBeDCHGctvCKabr+w+pirkYo+uRwf16zLyM2+zMt
UHxYFox/K85FBC1PiXyu9FnZ081sJX97B96uG7buvgCif7KafkIwO6LWz/s3ukoOOX0JRVfCg9Fv
zkaRj8fdBnrNLc7NoiumauZl5tfDqGzDrLnahBtB4X7odaFbThcSTUqHJOMHVu57uvoRtWe2RoOQ
rB/e4YEat9Tt6q9lEJi+EfQrjRIFwB5AH5hPFZHKZTQkMFWJrel9E8axyrrrDnohbtD4uFDUDOZ0
q7Rjegbxu3dYUH1BbGpSYHAYqSnfS1U8NBTfyMemrI65m7LEC2NyYD03U7bSUk8bFjcfyk487Nam
CGelCe8Wtwo4jwOxtX5MPIySHtus4KGqtwVWYfDHOr2hePyO80mjIaVHFiTdx7RmknendrlVjgw3
ysyxnKc19ZUzVoz5mUobJh405WtJvwz8UdBHc3eY/616radILgtWdCMsDYm0Z0wBdRB2+3AkqKQ3
xl3N+ijHPeNS01GjkUsdNl+53m+A2HBF+1bqrwSi6AlQVWpItC0IuPmsDqTJC/cO2IwzrfjdT+Bi
PbdhnjymlugQGnaopX3a2LwJp3v2es4IZd2zHYmtDI6ZCNeJmdDaAmpMyjT6tNZUs4tAoan6cVL/
mT4Qy8tcX3ENKQgYAlmksZhgYWQFUuZrY4KamHAGllDryrhkEBrR1lS7FPabvYNjFGZxOKj8Y/sp
WguJB93CKnaknZPl8gmbBYMoGwvTmby+iRU7DeJ/Poq3gPXyE6hjqs0LOSKgMrSv5l5hid2D7ipG
GEU6FnlG5e+Py6DjR0deuSkDB1FhBuY9k+1FWd8njy8BGJLaYnaZ5gaFpUE9yq3rHryQb/nU/n0L
Vg8LOUp9LVIygy5rSXWE8WqciidZN9VOYJhY5pj86/25F+LZWJDxtStrg5tJJW3ex8GmD7v1BATJ
ihLltg1Yg0qIeJPN+ZSHiwuCY2XRxWk1HhuldTj85t9zobfZnvVhAwQOMYZh2kPmpbnZlEMnsQvT
Yv7VDpz5g5jPy2W41L8PdjjGYA/MbfkhHMTK5rq+mPc2tAp9FqLrvFrUewj38conkeH/AwO/zHer
TH2uGViVpExow9FMIZpZLdICim92zssho1bITmcO7vQWVb4biqFmv81431RSv+Faiiftgy0N9B9s
IO0X/mnsS+FMOs8Ffa6bIFaIPs7H6HKe/97mbbxrCPLF9/k/P4/L5Yctic3N+tRcQ74uNHCba0l8
0/UusVb2iCWyQwBJfHlofWOef+pDcNRcSX/aYXqWICHuwvh5L9EezRQGjTDwp6MaVI8MKsqvSrvw
7tRAqrf9fmOygcGrd+XroQ4jA16wrlmwP6bwAo7paWqHJKWUsBhjLcHaMW5KtoelKBwgahC3dd2E
SZN8SyTIDeuHDh+CtxnzSnIeGQYq44gQU0CGouu1NawHD1SaWVBvYZsgN2mFe9n3Zo3utQDCoulk
ZQOQ3uqhmMFd5zJMPVI0TIyICxQzwai7lChiqcD0QgYXu8+NttC1L/SPKDXVngi4kUrZ6oIyLtJ2
np4LInXMY4+BZ9ndateBCAYCT5tvCH6L+oJyU43y6c28qn1B8bzFmEpRAb76vsNopbZ4C4HYqDuc
p3oPfBwJcK3QLxXTQl+z0TqnwLYCTf3NCxaaS2SV+D7qCjzCnDEZZM+zy0fRwlUVlwqgK8cVMKYA
g6fzFv4XBZH7QnldeUIIs03iEZW/u9+a1oDhdxY4GymBe4QHa9EZYIhT3lLVp90LCol6CO4rTzea
IueyWrl9uaYYauydH/0EIOnsjj6pCcrM5ADhsVXE9dI1dkgtVh5jPb02edu29kZ6lBl/ZCTwTeBz
H/1Xplf/CCTGngnFOHDqnxYrd6cStJvesR17j9LNFbEZI7rTkp16WPdK8tRYR74O8TtTBnFBvZWj
ea2El/TKACpH+QD4iG6ePKUQOxYNn8irhaTqJ2M+KpK2JoZPKTqJqq90smfFtpzlYGVMoEAGbUtz
3KCm5se6W8ZlULgCx5m2XZEaDWGvubsE5kOKhJNX7VjzpnKsJMuIyBGEeDB7pCkP/hpT/xMFSL7i
PH94RqiEdDb4iMSmucgdLdDf4yJHFqXowiwhWkdwzu2dJ/L6/hfpVkfhWNQgzJ6D+OeV/58Uc2IE
YZnVpUyO3XLqbAAJgD9hA10xQ31++uqwGrFmyUVccKqWJelH1y73hlSQWBtVcCF0UtNvMvHEofLs
S0ljr+dHqsTrxnzqjyezuHt2NitUR52o6wejojbBcQOikAzNM0RQsgZI9AYjDPRaXcwDB43YSA/t
Uh6wSmQPPlh2xgq2Sa4gqFESy5rohm4gyHQzHosZ6vg0kG+OC8vcJXduj20Rs5IpI82EonMZ2yjb
YgT0IBakxW0ybW60mOxqy6EslzSM4AbcFG3IoPEi4FakUQ2NGg1u3BXQk7Zcmvu88ROWlD50xdWY
nSKKq1MONjF5fzJX52fIy+xvHcBKCFTD5y99+QUvpl59cG9EZ2vXkwnvgJ8bET3KTJ+PRStwG0lU
2LMLaKzX2s/bizmGIxwN/ZEKzhrOwKoUkP/NXe0oX78byeyAraVl0MokPXjopcgosh9QJlr8kZ93
jgRXXIbCmIEf+Pmtaay77ZXr7gazHoYxvHPEX/ZGRWWbSlY8N/hvusfGOVFEOkFvqfXJ94PVIzs7
wGJ2aEbGtgADzmJshBsvtkkahcP52ZX0wTjMfuIQ8Sgyxc3mtDN4r9eW/kI/UZmCdGLCek+IKkeL
73Nq74FfjbZXhBd46be4RzeK3OYzRtijCRy1cq7y0lkMSG7j8pkoYoq9cBZM90QdoACw0MVFh5Sb
+WehOEC4u49xtSJh5Hwi3GSfDZKrADkBUmSzT8zZ8+bYcIVJtoh6cH74RI/7dZyIyLALkn7ZD5Xl
n6kMs2diPtmufauB5imvAMongvwcouohNexiPZt4AhyRN5OJRhSEP0x8BXn22BgLOG0n6MI9AVl3
ZtnyxoVl4ag9PRQwsRzZQu7aOW2UzX/+es+PuuTARvdkMrTDX2TLD+vMIJb4FWh607+7a8E1WP5q
toIWjgl/vepl+R9SADhwq71U9IhH8rZZH1X4pgMseNnc+3PWCJIhx57KU4aalG+D0m8/DnsIIdXk
Dt82buz8pkFGxY/oIKeiSohdjFNtxQRrd/OjLTAe2pwdZLu8DmGb2EV60zYSMbiEpD0+e44SeDgh
KzinM6P3QAJ4fHeWWkI5mhfT0eDtI5hhPSJDA8c8KB/nb2hBl+76onfCWKwsmZ/YaeZ1hP+ELF2n
KjTexI0/rRIR5YDzPjkvBfvWWCmYTj7meaZuX840WbiC2UIGCwMIwAkwuxeR2SbVoNIpY9NVCAdJ
HOkVdigk/UOWtf1gmA292+o5W7eowdFXL9rXpHnd05yiPzbmTZKrIs0/BmMv9WWhCJGD2nPxUTmd
MADYrm7cN5qyOWSoehegAjuQ/5qyXlJC8FI2Z4rI76lrOsIJHWZNpYtaTfnj/RqStTXy/8d3HY3q
3j5SpEPAzTlT5rUcJFpVEzVhlVskj38u00i+yvT7D543Sa535Ah+jan6GKQ2Bi0mOAOtBGiGIycH
eFPUgOUUhjgCJW08u6hZA6cbZWDTQWOHk923F1EFK/5/p6rVS11xU1nA+runcdzdwSxxadS1quOz
FHNFkMv/HpiVau4PitWXZvUDXc2Bkee+bAH08DI5DdcuS307xg0Iqfw4i6qTV6yeRZvL4xIBajYH
uJU7w13/1WtI7Cr93nmQPi+zw0y/niBr78XbGg2mPrGwOkjtG09HmwWXteX3GLVU7Vd3Kud0OEpe
ICQv+hRfFBaahvJHjNAjqkxG7TnaAdo6wiLI22exdGeIugZIQw07UftaYtYrL6egfvV57mF4hQWt
sBH/QoZxurkoW/niQsacG9jaZ51Y/Kpqwd+5eRAvrhqZDJgr40nneF1fcxvq881jm1VYiUqwd5yL
WxktTDvQRk4NJkAdLMMywoTCXmoKs4Lq/9zJb2IvZQHSXQC0oD+klJ++/ROCzXSaAkCEgnhGwFQW
z9OdLmIg6cyjzhD5inoG0AACH20Shy7LSh0dx4h1XL2/1mQyRYfbkNOgJQ5CrDuofUNGMb0KOvRf
JrRuIh1dlOkW3gr6ZWut7YQT+0SgO0JHEJHo8q7zjus5zW3DeEwoJneRi7h76FZtEMXLV/sEU9c9
YWFjhKXfVqXpGyScnGurMoKOw/5PIpUTYlpLd/UxnBJXiz/8JwpYrQapl1JSy48x7othZc7mRuNy
06ujYY9k02UA8dqIdfUrt3Aqn3hG5ObksLiloJeIjK4/lCXCmqJlz4K3lDeEYXAK6UIJlPYm3yCE
hgypvrdOwAIV+07mOPFlxMUuaBbWaC/Bt0zsT7azM5/z8AELE3+sugP9o0NzEsTEH0oaDh4Lfz2R
UDsibmgUPT345Fak+tr+j9QzCBNLEFossJ9jOjVoftudWPfN2HlhvHVzCXHPptO38fcEff3QkXEV
34NJ7IbK4TnXCzjZYeuvDSObr5Z9pC2bmrBMH983dbo69lDoxY2vCJACbBcwU9+JAdgXPZAqb/qn
UrG0lv2fNN0uK3omZeJOvA1/EyBm7UdyPhwum0CyMlsHF3lHjzXIZfCGn+nUSYnkAsFhp44FBfQa
dVo1KkPZAH/tH4FC4BRWD7+RNbEMtHmLJe0BOLSu3RGDtcWm0u7JMmeUdHnTScKmpHUdL5jnZswn
4wiAoZufU2ZTOMhwBuO/Yc/UrcFocJ3wehI8PWa3rbZqmERkB3qd5FrYVwecvdSB6+hvnpQP42pZ
DsYZqYnelFikXXekSeAiKJ3V6l9ZR4rDKLR5uQvigP+Ni6pKu9hEX44oiECsTgU8YwGPlx9ESc9F
qH1VHbxoMeu/e2alGerubDXoerHv1ZjTYQb5alw8SdrkBs2NKU3YokG3bQWXhwVi1ZVb01ycKcLG
4Y6LInFLD15xB0cC1Cl7wToBaFnS2PXS5bLsNHX4ELI3HpkQwBtjTYUiwHOCuPrdbfQvD8iVHZMN
hcJu620EosTLmbwxadPPJAuO/JWIy4RnMP8Gwlf3vu4iTrV+Y9ZMgz8t2Lley6JRcCc6NGwy1CrE
K7xufRE6iGB7fbP6sFtYg89/I9bZmlFcGxwQ7SrbFL3TRnJHqng5xgLChI6nM7MCLVZ+cyvwpgGF
j4RMfw/o3rl0mRaV2sI+aUmKPFPzWXT9yUpuvCb5V+CyhhbPgyD49UBtXQK7rra3qDWA5KjPp2ju
vGCcngnm3gW5E6fXed+mybfZRAVp1jnnHQDOs1HpG9Yf5tHUJmLm+F6BWQDsBNBCVcJ9ge6PElYh
IkXkmbX0QSlniE6E+Q7oPXbMUxpkn4blQHDVsBXDa/2/PnA/CHKuuor93cvIe4/Q1+WIo1cMV4fg
nOwaXmw5NpgX6NDuW84R9LqNDzkfjUu/Rh91Kw+SLVzqQHs+683oNrEbFJ6AmraA0fIMdTUAJ4eO
UC8je1j3z4f0Wq0EyLdz0rOnqj9OwbUeR/vwQGWyV5ecrIGGZg+MSNKlYKrhb14MyZdJG10j0quc
fYr59JoS7llhu8FxZzb4llg65/3sZ0VzSIGiVi7Rlf+DtcAHiJp8y2VqEqnvXHsvUP2360qD/lGt
O9mgIgiazmL2fxydZr4jDD1hnONLKnOx09/x1Lp2N/zO3Bc4uG2w65ywq5T8HG38DgdUxj03tIQA
Qi7VPUX19Da3sT/l0TLAlpaErwg6d2aJtUWm3pCjD4ai3iT21fxKfDuB/ZKf+2JplqPQPgEaS2tW
q+t1wQgVi8QJWYrC+JeWyKmBrsrby8NTQziTknp3gsdhNBoCYvXSI+GHe4Rn03BI4RnnBaIIe69b
0pNuD7BlFAu/2f6XBibaq0XvSSi3qF/3BMJIMK5R5fT4SBbwbjAP6L7CkdPehMVOyjadD9YrYFix
NeRrUlB0KihlHwB8unKH4qOdIQm/3FRzzS62PIPGN4BLNRRI5Fkecp2WW/d2latQ81myjvs4Dn6N
uDZv2fIAP7M3dEaYMNa6uUl9vWim+yshTeHnayqpN7SSB3typ+Ua9XHstPJtsNkvgalzLR//pBtX
nHWGT1VDg4F7gup+iLliHfvNMwfdwriS6Yg0sRGDc5VvZxbr7NtrYknhVt7exoE3jE4aiA7G5WkJ
SqCU8W18UnqocPnhiKXva9dngBc+hrfx6+uRPMnHFPwWNNxIw1wO1dqAjdN108ZMN5RBiZdGlcdv
fZ6pyw40m74AKHGPuLHEUtrSOcVGlFExu3yc1lOPMsO+4Od2EuO2z9bmReza3Ux/wQBNcRt8JzYK
c3jdHrzrCC/HvF3z5rIlfMAmm/eo36EBBCeBXFmUQKPhTgONxdYbkYt8+LcVhWhCNjMkf+oMyKi3
cSTEfIRBD2apoQMKHF278KZB/ivsX+FCrvb3P4+NaTZvX+ofSLjLhn1LQ/nu0tC8yhRNTjFw/dHY
acUFufCwqG3iowu9TBAQgskJd0FZ9rC9p4hRFmKN8xDLO6mJfoROR6TnwfMJfgQ86JrZ4CXxKKRI
+I19R08MFrzjiAd4PFT+CDQdImjV4f3zAc6Pk7kKlmxm/RebAwnY+JLWZ4P6517ENEy+AWX1rKyO
V4yjuZjx/tM4NVum8kU67EwxBz0qcfK7mxxs0duU8xT8v+fSJbJB9KsB9fDPkVqKoC/6qZIIgDTu
cN/g3w59tLNJyZaz2go6JuGlJvQDffViGJ7ji2HbS8Jj0Fr1gE1B0mcruSIEJPBpnymnkLZmTwom
SsBcXxr5+yn36PmWmoH/2LLIIFnyzzCRGXsXkrkOoK4gHzEZmjW006jcv52cL6W8ECbBPzSMA6/r
dd1O9pg3ZEptdGCogfF3lvwRorUmykGPFKDCEJxqEZ5A9P/9Hw7+brPE26CmeUJbEt5bWKg8G2Lx
errTZpZa2H4Z8LcgbNA6aPMa5pV8JuULUJCWd9AQYzursreG3BKEMI0PfT8pyXmOlJ94V6HBl4gl
fCIpARP1MlJEbJNeCwXvhAFQeZwfYjDk3vxEzsyvB0NjWLyyM/q2OIHfOMNVz08dscjghRGiDRHA
y7mN4pGgZugOMRBgrVHpxOIOXnYYiiY071PMEf7TvNt2S3jr7AvgnFSVm+C6rTpYZVHBzxfs8HAJ
GjKmBPqQW6bxMDDHoWBQ9dgs4eGQgPx0bjtr/c8liJ4PZU0gkpu++OcQkJ5yLFgcZqLGUNzcdTJY
Vy5ZQ8LhdIy1vofHYzZtXSWa51zfkQf0eFU8gaekEYCOAfJOEQaJSoqRhlH01aEbt+GLtLzYj8zl
vugIGWBhXfqoo/wynW0TqAW8e5AS07QEih8l09p+SuUNtTBToEi0FtJh0uw4s7CBvom3I7r20TAr
aWh3FkkeqwGSJ0oK5+9eVNeNvwYJ9rHowqtDy+iggE1Oq34lCapTdq91J7pVW4F39xP84cUagANr
N+Mi4PAby4oEJTSpGfTdUJEGuNm1TvtYewZQ/C1WX/Q/9oWy7zciSDOiQYI13t0G/M6PrnHN/4A2
OYrI9roVumOHtb45WMBx86FFuXK6HgBJUgjFAcQ+o60GPHDK0tXTrJ+oqCQDxuT/NOxm3ZHM0YA5
HUrhH/VFDbOTRERG84o0nTPTx46P/+6QxGHBieEqMBivSCd2oX5SHFFZANGE9XOPON97VpIAD5dS
dswx6DE3MZgehxCpcVLgOc6YkuFU0nHqqQdCKW8+BwQaw3XNBGQpHXv9OQrBsw3pMVh1DSKpB1Zh
bLtNWIB/3gDtGIeZ8UyvmOgXOigGnAIVn7dtMPRXYPT7sVg34xuu2lAnXGI5l0sJnHhB43EHZ3n5
cp9i0Wth+IevirrZ30iI43R8olp4WYEPoXnHBqnG5vdSu30nmbafv14zLWjIPnI9j4N/PsF6B2k7
T/5iqSumcyHPF7TqMw1rbLp/AU5ZFDLaYACJXI13OMSG8QS/HCQ842pns7ampb/0lXayrS8tCs4z
FeGk76SZm1AJudkJquUxfxf5yih/OcXd5qnR6rwpUC8qpLbWyCpTpF4So+OCCGekg3haMvnBa2bu
TBobwNlKDfiBTAgQv6YZCi5cskD9g6otyK9+jmvPsMzvkWhgNk1QecJHFoSVrBTb6nXRAvm8wh5R
VCyha3CA4bwQwQ3TGhkn4Piah5/BXd40gaI+4Xq1cLGQvcCQfiVvfNMOP4LE3YYEk64ZNZjaK0yn
eLyoX0f41Id6Wtlpn3c32hAZ1RZ/T2A5KX2wLF7BCnWZScMMEDxwvUju9k2W2KXfoXDJcArx/a7m
XJbo7WimpK34oPq0pcsmUXHoLODlrou712NwNMzUinx8FOCxgHGCpK8vsytp5a1BehnsJuv9sAke
OUf+eYeOIWGSEIH21YGau+eti0L0MCiDjWiMZdWT6Cf1m5YvxMJpbT+m6PpYtCt4e47Gn9F+n/0k
04DHoEru6VV71zSvRhLjs0HvkX+EP5zGRaHhEllk8bCE+J1jKoj7sVIOoBWlUHWJT2jBVcKOrDYD
HyvoCg869eP9vL3U4qN7EB771z2nhjmqrS4ezXy6nIGtC/sUX/lN6SRblIulCIQM5jnNoZoLvFiv
fmDN5dQ2IftFJlh2+aFG2ZxaCnVMgKlWsymYszWqx51lBbEAaDou7PZFBDX+MDayzNYW5c3zTKnj
dWvdfFa4Hd7MCtJ6ne4Ll3LzMToQBL687dxFlHbOFk7t8Zrfd7gQQ0RgHbfguNbyPm9rV/ycM9Pt
9RZWNvN9hTAoGXuNWhrIsJcvdUrGJxpVc3xIK/aIg74Duntivn/T2N3i2la9WhdZDjYPEqDTrlPJ
/kU2cvQ0ReYffUrscu8FRJZF0IK5QCets+WvXGfp9sObmzMDBxFcynDV9QHISeODXx/jNSzMif1b
ooNghs05c6MnT2UMmRJ+fnyXlFukAnRyWsNfjhAc3j8XAviPFZjHq4bC2V9haBujKL8E2hk5ST3Q
+RiAYq+pyAgPf5zs527Z4BxSeAD2AAE4Y4rZ1JB6qRC0U9pIYNysMI7lLoKnJbpjbNhnSQ/7uDU4
KE1ulRcYg1IX/3DZd/8I5vx5Ry1lBiENItdr4QAdt1FLLHH8FSofVR0VaDrTRW1yEfTvrQTXZ5VN
WlliYOxqmolTU0fS3tMx+I6n23kn1xiQeeZVCRQ7wiRDxwDcN1l6S+WZe1r5bZ5HXfxx7XjXiCut
IGB4Tx3MYScx+qSQMf8j1GDtc2oBp+dJabiwAssJADMpwCmhfV33G3tiSaY7obBY9sX8eTt+jQBL
QGtYa/R4N8wzQEZT8mh2sEhBG0xKaS4kmiz5hLB7n+1Wy5p60hLvbycchSImPmt9ch6b6R2NhsFH
o1ykwT2HYqpgGJCn6dwXTpErfmzrq5P85YIXqZ8nlDpsolUmRuQ2bJkqqIgs/T2qmQvZy1iBzQn3
AK3uvZJL3HBvzlJIyAg7frGQaryIohPSON/lXle/FiHhOpx9kqfcchjyI8IKJ3En6c4kE5aBz8KM
UcW43HAOPUejGsFS+k8JPeFWWeCgXAJYlfJ3e0KKwGDX2jQTYqCN5nfulUfRp3viYsN02WYT6ZJr
cuMH5o9Iiky5LhLeQjGZdFAQnZ3/ueWDCcSoCfmIAyNWVqZwh7StpLjsjyfxGKBJ4bB8Z0JMqEvT
NwnQGp6GDFiZGzU+kZLSPT6fISr8ac8wntHk0Bza9GNnjyWHh4XfraIAtdprYVZRhYRofKmBNsO4
FV4Q+85tzmmqVzkN+Xs6URh5oSWFd4bl5pTp9gG2O6MxuaXnlKuo/JDZbB5fu/TAjfaYuJt1JCPB
PBQf5c7q5gXBejxQEjFvX3va7FAW+ojk1NL1RzbI1PPThBx47fWPtUwvdILgH9DeYZ5KAxETzkyO
dPIlFb5VDwf9V6LaSBUap1DeHaUU4u50AunZwubK6hdV/sGfVB7jrVMLw1lp3CI0DDQgsAx9zCRA
3Co2Vz8u1XOWmytr1xWWzPdr3EtSHI/M1RRhbw4ckb5ZHZS6etxrd1Mpup9UL25Ww5dH4hArq/dP
nH9h2fETt4KrdMSJGao/kirecUVBL/rb2QTdjd8wpMtpDAEsww3NFPYy1FnX2WR+63UnO6vgCzJf
PNG3UWlzzy3jSWHYHf80iTHqL20baUVLVRfK8AWzIjPmx4xkORyh5aITM7+Vagm8gbmJJJpN20zg
lt5zdnP+MyUd6BABCnlzGj5zqwDVWTSmuiVI9FuDVloUwJXIV8EDPHFyr4E21lCa2VlHKPRAC21V
KpB9NaqZd6tYydQowVJxGkQYlPEsnJB2JWV9ZQCvXrRVND0YaOjdqZct9j12bvLgG6uPU8ZmHp+z
7v8/ZOUz9TnZSgrafSbNGutG2ifFfBol4xwCr5mkPJHd/m2fdaz+WPTmfS4L9yUTBHaeluih7u8i
0g6y5i2SI/3cek0jkJqmazG5NEpU8e0SxX7rZk7ksTHBH+HPwlRo2O/naAwLN/Fu5Sssg9veIwJj
UfJwoixv07udbdlwToj/xAvbqp0NDXezG9YBsUQKH9VWDVfVO24lhyYMK/8aCVo4LwZ1XE/4f961
b+gjCl2oNnoMvrs4CBDdPPmW6RV+m0ftoKBtndz1kOJU+PoK29UBcqbFfmlkRCNNVk4XiLxpFLyd
BSt6A38BZ9lDMkpmTWu+UMe+DIEQjKIb259ArhmgVhxZWhlkNCQeDngCzGl18EJsjsyGSkkxxm2k
h9Dh+CYKJOmYCnjWmDW6juRSkei90xBjMhLAMN9HZe3GbXwP0bmS6/88TB35qu6T+CZ75WDOTUYF
JCHfQTn6532QP3/UhpZHj3vtBV1q7Tun1qOTYJ3A62yDZk88MWw1DhjzAOaMmnNHuJz/8VQQcDlN
WeIN3EtHhNFZlMQ/3lz34aVRpmN1NNCvCXhBMsHbQz+qZZYaIR5GrFmBjs/o1fZdyOw8hIkYthG8
VjmoUMe+5GgNETkbCsWkeCAqQNmlcCtNE/Qm/XlhT8FT8z/Y7xaZPR+/AU45siRa4+UvF/jNtwOp
FDMUq2YJOSIKfJhJqtJ0DZIehdrMR96qjklEE9VzPELPqg2+HEYDskEqkfXbfdNPRZY7M4rnrg5b
P651Vb2Va4X+mBXJZvPyeewKjE7SnZq+ucTDvQHKzHRUInrh2Q6Eq0sLSxD7vuMdXYlxsupDM/f+
AbN9Cro8CSuZON9IDK7eNf3Pd9BbqYIfFPR9jTsayT2oD3zNZY81yavOCvxkO7lkVji/iruqM7Hn
oCIitoTBMm4lMdRmzRxvA4AIuctSOO+UoAnYXEBHi5TaZiyRL/LtEzhl7ePVyndKBCmOHuSCRJjO
39sWiaKlxAn5ygFFDdUsnD3Ulr7Icvr5AVtLjH7hELePPtscqxgDbDy2wLx94yXxHMIMk/1wemdN
YW+FU/jQlX3JxUjlgp5w+GmamzvBy1p2VzOge9IPI289Gg9f1TmW69B8Sd4OI72ki4IrKCSLfIwN
BQWO6/YNXhmdA6EuA6nTCh43Cy1KHdLI7hMudyNpRjTfwP+GOuAaPG1dn4WUokfnYX6no1AFpKhW
/ueIqm85Ke6i7i2VhmM0sOf/MYByi+72h3aPeC7ITJp9vNzDzWS7siO9bKBX8r18d+vSHxJsC/ml
QG+Ct+FUM6OHc/y5LoUndtuKPyXVSduYqBs+9G6kbCMQN+sNzSQV/1G2bbHSJ0uBM1BcZ1Pf+ZP4
FsP015uL1TLS+WeDkHounzPtYu0xjOsVHfHGaE92BbYIYGr8vXYGAeczlj6j3t5Qbfm00k97jidJ
5FkIS+jCVC0e6IpEk6dnV7/i/5u/h1yfMLLz/2pmrdZ4Na7FSnYXVjXLZcufNmt9EJCuh/cjIR82
GCNZnRu+ok454hVbUblw1HSPqsZg3deSRP8N29XcmXNWhR1jYYWmKcpBJzsaiM012XU8x4ltsJQy
81narNiwca2L/AgT7vXSAQDMbeFhK5WbfXaJqHobNYg8FspwMbYOM+21H6txu6Ytg0n8jsbi81ka
5WtFWq2kWM8EPojmCmZo94vVRTQO1Z3c9pJ4TJ7D7NMR11bokJbgSCZ+fQ6nnmtDknJWz4q21bZq
Ll/oEf5xI89VchsfnMhu2UMjnudBoCsUXq7BKtORyN2zJO1A9yPxDR8Iz5cqYB3fqrOE6a4QyiAO
eBWiMD/8xbqG6q2AWM2CaQqk7GW1PJ9csKePLdYhFdOEzKjA6ot8LNDBsbQDzmI4n8ys28XgCtJO
54tl57bjlfwI3/TRpZqkBjLkJsrheWzlS270qiciGtQy1a3NXNSid/SKSQdMa+6zm5Zf/1laTHXR
diRruQL/awEfR+yQdv1eSBlX8Hc8GHNitpPxWTvjx8pM2NuhnkJ6wbzJys+c5Xs2a4Kaou/5j4jI
NuuU+HdlacCBSk/pXQmd+syEi5C4l/20OxevtpencCJUDeNpB7OUl7MQpZXsvBwBXf1hopS6FusS
fzG0LxImZaEdcb9CJr9zkiCQSaj2zICohZqu9YB/dnQ2KXE/ZvVlyfHKQ3JaoC56tEGM10pMsJel
7WaVekRUCXSvdHXwNvoKQZbrsiYNEaN33NIN03Gac37yxKJZuix368OaIhO0TbzWWSdy8wcahcwD
FlWNxoOhySAbXgMUkm19xj8iQ+kGF8je39IWDF8GV14go4KiXocF7AHhJV6gDJ8xB48gX5LH75XU
WaAeWYvTMkRUyqRePsphrVhjVvcjlM1Uo8kx2ASTpYq/Yrb37F/ANe04E/ln09I16M6x0Z3M+TyD
kjUASP0BaVJgdPbww+A9SxX3EGkv2xZKhaguOq3eao1rK/5vhPoQnk/s6Ace98o+XGECazTQaYti
JKnpo5tK+hDFuTAMuY19k1E2vcTtSQI9vhntQeBpWYXP7hmopOUHJdL1CcDkMRCfTRXMfQg3Fj2U
x83P7czn2S9xxXcttuMgXJZmrd8eMdSJkJgKQIxUgjvo9NDyyw1c690XlwIfigPTznILwRRwkGjs
P9W0DDy7XqS9xTcK3zUHnGuieyLZD33y8Q15eb5/sjFaTFbJArK065F7jWsaaIXAkAwl1c1dgkqa
7XPtYxqXIKWs6Of2GOEXgFgwlCmxtKVplcUk10rNnEMAbTOtegQN4NqWK21mTJnORvYq2BqV3PUk
b1i9hiX+fMmqCTPbmxikgx7aDp52a0NvRMJaP3rYbMQgZ2CujzxQFIqNiSEC4GksGsdRbxRtpH7y
89ZBzPhIwljxYZEyhr/iOGj1mLMni+v8RKrNCQswW97QvQvRpc7x0AadtttXiQq4GqI75fB5Menx
FSZqRvSadPmxEdbYtUyGXK57V/kJhWWDYsL0EOLMTzT6divmP/mrWgED6gVXRFOh9JTU0/3Xi0Og
A1qOg7zZ8vfqHgh5YX3QNKwRWjEdhobpDm+3HqLRNMiHugdoljnRRCmm0GnBMLcohWnfaj8WWj++
897WsaUisXoj0D1YKOt3nVy5qRsdoJ7teCB5UlnC7F/C10O52zOKf9K8Hk5k9S7AerJ1h3CznpC4
wnqQcjaQmbQcOFAgMd/dmQsSHef6+ygbcO2T3YBITrUm8PH/ASZwGlRBTM1ARnAYT3+0A64+jqVL
AW6uiC5PvV3mI9xyYXMWwIgBXyKaKL6tKbULqKwyK1YuZqyfEDUxOA71dreXd7dFUteDQL7xJ/CF
sQ+JhCiHrqrPWXy863mRgPpvkJnRQgOZHmN2LJGFTRfM7hLjeblIV7RHxVtNvNbLOjZ5NQPTpaWZ
NH2OYsIrwdNjsIll+kfgjFEiu9hxDtbyaxUrm1BtEjXHek4oQul7fIL17+pdZqgETk2eShMo+C9O
ODhIiDsjKqzX8DsoEa5VQXltcAxiPQaUIbrNkykNnk+9IGrzTqZV7ZrORAtc7RqrQAc4POkr/giv
yBgKvJgMsYP/C1kKpImGuPGYcpPb6cS89wFw59B+Qnb0hAK1watMish4Ty/zR6CgCBhbCLEorwQP
q210h1RDpl5h384s9PrKM1QUbhz++jGEP99D5w/uXhfTjJKhdMX/siAxHQjwR88u2THtZQURuDqw
7+c5mf/5lovWcoo+bS0aKlslELIeaZxU/IoIg29gXc9fE8YiLWcvl8ee1FK+ZjPivCBf5UE0bSmH
fFsDjLHpKncTSsZHvfcQnwuF2CUv+DH634cH3CHqOUwsFrN9xVzT7GPvXN9QEMrGywXcZwXj0cIs
LqVDb8VUiS0aXcyaA8fkVRDfuFpivbYoYM6uEPYyNqyYnpYWDXRS0nf46816h+EFENRQ4NOyBWc0
51yju7qcKIzmSK7+OV+6uK4Tpqq/X5U9seAGSBtvYQh9yL9JkFXzE1PYakBG6qyTroRfM5FkksaD
vVgfoxYqzYAofGTaIcrZeHTsnkPQG7YODSI5+Ctld9mcR4NA0WzH741WI9RB/ZNonSLbXUBzu0ph
dj5e1GaCQP4Hd/uEh31nBMXipHO5YYu/zrZyZo8BKsNcNmPa1FLXpkxdLWTH1ubSlW2/k4s3JVmu
VM7rVwCyk1BDO266IYIS4noQLqo6jIQLzSRWmblGju7OVZUgYU8NyR5bzYjq5ILHGeukfOB3sT5P
zpiQ+mTuCGQuQXXMWHOUq1L7KhgUZYpYTST4cJVx8fME7QtTdSoNsZqtG7RDnFaovxyKymRkSETx
SBN28vE4r8PRJoBRXtQXwpFCyO/01eDcexTnQDotHJ2eW06Rn2xjm0SiWzS+3h+SJi3aeX1jOCWB
UbVhBx5+q3iSN/ExEUjz8ZIgNYMqX/3Aqb2DlJVQNyYW3nNp4dwZfyGRG+9jxkQXphpxscHrY4Ng
LhnCcJo6of0O56HSK1Cwc1kr/nlXlhQwB8+Ls+nMOsP3ynSf5lkwPZK0UimeglbGuJ7d1camzpPO
TV2p8Eb+ZxKn454G1km6gr8XztrasnXf2Gi9PpGpuTblAFPXGReFl7ShDybNZpCVXiUvp0MWwVoo
zGMtDfFXxPi2olYZd8gMsP3mKPyL6T72eJE+wIa8vYwlHyb5gXFcpyXugnKqQ4txQj092krtEch4
Uic7vlSA/BEPGmC48PN4SVglP9O4/zoq6bbU3Fx3Z/arLG0qQlF+c+glfxYDbJkV/XnqcE/Z2eTZ
S9zLi+85CYvpiX+Hvy0zubp01D5D85zESQmYliOj1McG9ChFGUSfhcAtz6ILzbwHrDOzYMHInGGR
fYLkn1ucpRWjlrgnatdDSKU7ZcTzrKiSJv75W4itJIEvOSvCIDnU2dNoQbhzsoaxBfjiQP3pfb1C
c876J3pevpcFqqhUEkglWawNndsC/WYikbblXgO/7GLHo8zCpmUQarDb6QSfCDyU067bsb6DrzEo
Zj+5RC4dABwgpLZd6Ws1dK0TYYvRYH4dkpp0Wc5KzvMayK1fVKwdNGovnPwpk7hc6gGWgvL40Awb
+P9JmarizP2sX8arQaRlBpOMBu/bApMM7yTJJIBRu583X4QSVNj6/EbNnIGGury+EQ6dwaPTQmpS
LZ26Tj3I1SUdNkeDkcsrB92ct0IqpNETez8/9qBTSDzorwvF0SxM39AvME3Te6ji0dYfUKbfsyhp
hRr5KlnTJ4me1zKGcbjIOsimk4PEoDaQF1BGW4oufufdWEeJot1mweVCokyEPpTKszx3g9g1ruqj
Xv2yHec83Uq7EAnlTQptKtcTb7mzduAs7ogcTQ0D5u5/TTFGTY3m2slXkgXyA0IRumZltAPQ1piv
Pmp2aMvX02heCppj80nHPiarc5J7FWUq7v7A0cOdPZkLH01fi+bF6C4/hmMK1Cn/SaluK3Lrum3u
IGR1jdEyJBqkzbzA+KqbkNSwq3ZbsQYfE0dJP2MAB8JOPN6KiSpvg4CjpMT7L38fn4O0vJ6aksD4
e4Z731JtuHH7fuX+9R/Sa2kiOy3HOCTdEWZPikhUDbaT/0fKktzdAkk8BpxW/vqK6QC5lexi7GiH
o5BBNB1klj0ssmqE2hqamP/Pii7tJWkFrvYe0daFX+6mg7TEGKWDovU4dN8LnpXJGB3gVUwXwp1U
hzXEElT5IRoq4UD1ss1HfbA+shIEgc0tAGvp5uhph+xk9BTBzhVn9Asv/5BOtLQnLCtkZXzNLyrt
3/dUxTHJ+1GN+Tfa9mRh9ZihOt72MxE0Kzgh8/KfXpbXpJbkVueeMzXO370/WxneHme2h/cRJQPP
mtXgMSZooOu/g7b0MwBRD6jfum31O6psLq8Gqg2mdfl0IvzlKn9J737R5qfYAYZbK6LYTsBPk7MJ
tXLjfoB4y0mFy4AEvfzoRM8UKZziDTkH2hgsBdEKSZwjv8I3l9JXA5oBfmTKBRZHiUFQc1Wkt3rp
l8/OYtInnj1GCH6urD+q4zOe8Z87XVYY+dgdIDAueIUtLyZNbynS60ZNk+w8cnwZLxsZmua1LkAS
L0ooGOC/Sgu6cESCsGcnz19+pOWasbSfPSiSN7TqogSmu6TIiHqW+rOHWj0K+bxLKZBT1Dqa7rzS
ISHx/Dw+rk11Qbj/vlhVwIkc5vi70mZp8Z1LhhAHHOlgV0YSEZ9Wy6IZxNXglzU6OxZZYtZIFTEI
h+Oy6IHLppECeZm5u9OqCMKySnXk1a0KaLXw1IgfRo5kokUr9lsqyIGgr0Nwrdw2RnXt8yBGVNPB
5IZD0j75BklO7BzsSKx/ASSEagmv17Z1uOnBLQ8C+RvDgnuYwug4ccKDKrlvbVY09UxDxVzZfj7E
2rU1GMlIJ7wii+zE0BlTla/Dk5SC3IZxs+WJO2j7MLFrGnu6D05fReKRl+ko4Bh1Dh9ThhfZv/iB
Mq+5v9NSfFUaliV4gT/ji4n/EDS7M6MMIxro/f3by1uU794VcqJLBky2551S1K2Kvn/B7JFWuyzz
UDP1JVITBJ5pH40i+cBNY7ZHdTEf5zChf8Crh3nD4gOtcfabZ1VJ/dFDXSeORV3utogMzOWmBG1G
Fcf9VKQbEKyQzD8eI5ytVrD1wONCIL8xrtyk6bb2N5UnEY3N4KcD8twgxm+N0aiDA8PuvWh80x+O
pho/ZWw+9NHH9wI7Fw3WfKcJcAfE0Nft1XEpgRiYDxz9uGn+j795Er6fJXZMGuc2Cxj5GoE0gadh
SGh4JAmJ1sWZFjA4fMcMQ2gVzHDwBqp0g52LkXSISodxI2s0DIN0GC5E0XMQLkCgcGTyUvGZ3F1u
Kd2CRX6R+UuewPdKClhePL4S5F9pcnhZqZ1LsaOlcs41nT0ymhdJ8l/VWRMB7l6vtN74KeM9Hapu
Ep4r9E0VQj9KfdnQ48ZZ7VAQePduP0TYKAKE9zaffPIu6MqDxI80Yda0MgIc4J7qNwinQfDzakXv
H6iHJmOsh8h+AHxTRjja9FvYHDNX3bP40X5FJpOzracDZ4tcFbCOzI17UFkK8L1UyztYvfzobm4h
Td79NuTQxhRGPvzL8jOlYpEUDKQEp1VWs5p90MGfxEI51lkXXkdly+GuNg/BjSTh42kN88VjG6w8
AWhdEahdXtUBb8py+CGHfeoumX6vCzZRJNDjPqVgmD13VeH+/wbHDwkeaC9ACijjzFMANWDiXeaY
50u3yWFw+TY+cg2Pi16TQ1BBi/2o/m/WWIdB8i8H3oIwXsAjEOwXDqicBQ+xjfNbJPdJ4bI64Abe
9ECjldi5khExwCvVJwRpQfCRYWSThL3ys3+fL+dbZ1Z53z85hhVzIRQdjK8SLITX+rB38LG5uvs2
h5UBBMJo6BwBZpdBAisoh39vu9kh0Uek+YE6MlVTcufY4MNoAUQ0J888+TMbOCtyonIk1fcVALFz
lLFae2BUmnAQTQwyMTZwAExLdFj+2YRFScJ0ZAnaKTdA6jso2VzD0Kf+aJy2WX1qFO3XihB2UfXc
82Mytlf8SiGrBKO9cpQ0ByC98x9vFOT+CKmP1mYgXIn3Up8wbi4Lkn2kLpHTB+a4L1kOLB7sCu3g
l8w5L4MCW2UxfgRYt6sMOYWNAvFgkGxxRhrJTqoAXUCZDYV7K0glwrVE0gKHtdH7JVx+sxHdVeJA
9oEJZLSccyBFQ43RcTUkcen1qkgwBrHIcm3b72+hUlIuOT8BDMu43iczklbU6/pvWnd+kDU5fMx2
D8qVfB2MNIr2bgFT64Z21kwUOmo+bcTlDU0p7sFbJufETjRdVohPZar+LUTOXdqfJXFAzRZVm2p1
Rt36llbvRy5pgI1T17SybLWZSt0S8iCOBUGbVK2ZbGWG01kEEiIp4WZc3KMVeUG/5ngNg/vuJOQq
+TdvvdU7s89FuTLvr6H8tsNjgwvgSQD1aqCBvGXIK27k19e2A6RyjLv3y2FC2JaZvsyS0ywB2n5w
qYkJLMzTgbpSsVBwtxIJkS7lkQTAdRFRM1xrTXfZ4utsi8S0lYRGf7/+qd1dTUnptdZAUKrO8hYy
RavyTqotdiISe12XyHegtOmjseaeckTje8JJC+NWOxwliiYVD2ii+uw3at30ZWEnwVcYSSvVSr7Q
KG5ZwlW1Vnc1JImpDXeibEIX8iHqyjDhbUQitpR3Qim301SzDV8JnSOzh4s0Uxu80660cuXp3I04
DCbMc3QQ/hUUHl0wmKh70b/BXIFf/A4FYHlu1hS5ynmfciaoiPAYITVJ6dBGXVxijWuOiou2c+Vf
NAxzzihkWvn+GcbJM+CYFmtOpMQ0m/NCliOH68wASzcFHPLHWp8sQr50XVjJerMR9F6Omo1PF237
ImVhqZ7kaKOZeUgOiryzMywp8fyCt+VTtyFWSURAcOvCF9ixEOnqJbSOQk4nyf9AmW5sQNQOxzbs
Ir8iB3JU4PVzEjlAXg2uRsAtBMzZthNYhk63Lt/7WRfFcrK+4lHQoyYSsSLr3Z31z8b51XTUbiyZ
aUUxXUvc7XKnzKZjLve6A6rbBmRvgPRkyNQdwejX21CeFbScdAhCUKBE1HHa8aUEx/ndcajRF/gD
eNULBfZ2lw8qPqwFpyperzyKZN8++WT0sZCQabKzug+mV873jpZUjh8NHrx7tDC+Pizpjpu57nBP
Q6c0LHgTJK0RC99eJ0J65/ZZKyzoaFmGchJlXDha6RWOdpdtOElGTBQFEwphXdD8JummKAtV9m10
kwiWaKtphO/bYapYtYTNA+NttR0cCKkAkwgRm3ZgronXpC90oS3I/EE23/K/Hp15U1roZ/LimQbr
c1hggmPNsME61rXjKD9lFfapA8WcKzMqruObk3QuyIYI+jsAzwHOVKxQlxv0nwkt1tLDMg2/iejd
mPB76rUAQBjFP/EF0FbaYYfJ7oBPNxwTfP64sXoYGaIuLsbxMwduTXnpL+64/1YJwJT0Hya38a+h
hH6mpDlHB4VBoJS1shXfuiv1bZYNGNJCUz46SiALaQ6L4+5nijySZ+Dyowlj3QiWkNROzCWA3sMM
yqoQw84zXOyFyJ3AqUqCdqOKoPYCeirsZv6j+kgy2G2exBubyHGiDg9xa73SLzCFBXTpsIi7cNKa
tyw+fHRn/y3LQgp3EitpwFn7AWyMC07h4R/oTg7iIukE6zW1zLEqfJ7Ajq95/l68XAC81VvbPrNt
4LuK1RgoTuFeVSRxm+9VxYLwwc8XqtRYdEuYkq7eb92BaOhAsBv3zHjEdHGhbhlX4YM06Eld7igA
y89zrZ1zcpi/8r3I9NGmkFi9q4c8PID0IkX+zFFAtegx9qEmo2wvIpEq/cgIG8vp6vNcowHvOyNU
Mit7vj77Ti6jzED1vzdGFpjCzJX8iFwTHSVNUS8CZlr/SNpTHHuuC3USZUlVf6bf6bMbhZvvmRiR
fE3l85Th5352DMtmQMqKNzifmFVhmgOcsQE9Sz3Rz5SmwlvUqwj0WONyWHGaa0886UdeQp7Xsepu
JRGwMm2AtEZ0euWzHrNlMwfrMDblyWyYuOdKNT7ukjtQ6SI3h33oVCytPhKzQyvb/ykp/j683t41
dfmsVBOwVf3dRzrHmWQVcZooH2IxQtti43kp+nmo0CMRfALuXkpAh2J9kFYEK6U6cvXlUQySMiFX
87ED7Dz0naBb9rUpfAuZlKMSz0ahHRzcj9HihB04Yda57mclg55E+aU7cpp0xV8RnJmuUIxg6OCV
dsJGW/WbIaXvjSw8dEd4a/f3XzM8CWBpckl5kBLrT/Yitsh4cyYHinAXQ+TCvw5KKoreRfRBCFbI
0eHKEte+lFncpFIao2sJ4PEY/K3lw0uLUovF+ZexjCGkfTy4sqTZTxtagd/uHyuqTRrJsmIMZXkh
vnhZde/274p22m8zn/144KhDMELIEeqTy9u2CtAAQpbTWkd8PJkgSzVmFKJdQFf429KylpZGYjdv
cbbPLzg+4GfGlAhvlCUSTZpnBgF0+ZJBpFe4Bvol16IZ1GMPQ1GLbmHTuROxF+UeY0MN8rbzxA84
yuF75EchEJ0uFPz9471+tgDfFQ7hhzKir1x8nfUGtXecL5PoukLkuVfRW5Jj82YbyVrZu/s1d4pM
5Pbzd9QiWi/3vYmRVrTnpmgXSPOhrHpVangmxJ7E8ZvjjWvrZPhPltEO6cYRNcNv+pbYyOMBrXwh
bZDOW0unX6L2b15ZE+Xz0VPyaEQmNYaA0Ai/+XwHOfOC1814wHqK5CKHsAyRqijKc6t7fbxEnfg1
RxjTsJNwYDgqDsIHmfyTEJqdw+ctixVSsZMzW1iRRCoAi3jxf3A0Rxrr2YUR6a31oh/Q/iaHPVmg
qMZmR+FBQrRguzAPAjgJSbDlr2frBzKaLsGZfOvljvOC3GX+ejOQ+X1qHRJcVrEiljTC3h1fD16Z
2VBYt2vvUStJtxKdCUNnqCDUfu4GVgCplBySC8P/eA+Zm7D3sLYIUrR2gRMXszG+gozjbYd29tDz
XdK7xf0k6OkgzY+nxLB3Hq2iiO6mP85JpfEzDkpWidN8vvI/KBsa1PNpJIvAUaS58GHSAgbGTZk0
zvK1SUiyuik1H965I0Bscm2CALDQCZ8hEkYLjd14Cfjcdd4mzH27Vu686Ozh2cEL790XvMOW3h3r
ARV2E8SFbbtjJSlw2C5UCpcHVXNB1eUkF3durnBYhlpw9CAHWuaSKlRkKJGRRkPYDKW6HhDfjej2
nrkXmWQEgKUbyNyB5+mMSBqQlvzhrDlKjGxicyVvC7rVre6lcJts4VSDUACcUQad6cDMa7i1mg0p
tJgkZUYFYeaB5/75jb598mRfb315YgTEK/JMezM7OinIDFPB1VAqulfEuQElxvtaRC5m/Vhxxf+S
hSikTGln/aC1NjMqVeS46HI1GdbnxuC4Z5r7hCFSU+GUkFjQBcOwNuOh+bsMK86NKlhuXkyxJwBO
IfQu4H7Q0aEFhQbTAFO+qtxyWnihHiZRG1IhOenymzEne+WApwiIvqOprHLBP1Wve/G+RsxyQJFj
aJMYEpuZ0E7POO9Xe36/c8pK1Yl3zHZ9Q9pkUCJcyHFstT7oP+zHKMClm/XmdWxnSlb8Gr/Cj9Ym
jsR9HYlFFBBfNnR+gW8dTMnx1kOLV3PRZKI6LLclj7KIEu6erj6esjdc1HsBoMFbPu7ogO0crTjy
KQTvA95d0FyGKXJkjpQoOtlK90wEsKvEa4jGA7Twxgulz0AB7w9Fr0khwLe7WYxI/D/YKXm9sBdd
NG5romaJlaOgJhd08v63icO4nnXj4pLk6B2JjJpCQmSaHN6mAuAn4TiaUTanVtJhKrjgmBRPfttO
UcYCZJgSioIQzQj7ON2vxirbq+7BqKjHyxcqHvOjhcI3n0R+Ylo4SfMOiUea/coLXqbZl17iAXGD
+YzYhOcr1ZQtKl5AEEVNeox/FoOt4fmiC7XgavmyQL8pt6MvgbBqN0DtqqwF+pGvNgsCE7eiuiUR
65Eid6Z3worHDZnQ5h0TPY31ih/YOCNW1OITP7nPSOYUlBXGYjeDIXQ/0JrqVnOJwqGNC3f8enyn
Y7V5r40lO9z6y2d1qUMq5zzaK4/BEPiMDrikBPp+SdDgd/bXrKQqztcB/HwazCa8zs+Zb0YlXe3V
NOHXBWQC6MTb/zI4XUb4X27H0HBSnmSfo8DzDH0ZNwqNaezJLFgnTJirrU3ks8m9O3RIvMk0z7dX
rEPNwQjWe4DtsXIiin+zY5qg9rnXIUCzl75k7VgJXGTUk9c2Ig4rWoRfcvd5g/+KkUgJ9ilXpz1D
IkcGPBwyG6uJd32RR7V0q9Da1/kdxvs6BNchxniOvxXbVxE83BS9unDP40S69ZTS7bEaiFe1urdh
tmEcGwdZCA0Go1JyF9iN/pp/CocEG8VhWFCJIXX1WTaptJ2lSWNINtNpF7XQ/BSj1+8CpEceYIFJ
Rbq4X3n05Gp3IgQd6iz7LTvIH+P5wuChgz1oPnngMopV569u1ZvmF8YoSMdzE1a8BTS+693yCJiB
3ZtvVbFCfrOnpNLuuffsCCdfajQJgkp9nKEZko4WDMJ4wdtA1jBZgb+2jQq5GLqxNIDklOufSQc/
Dp+sVylWI7Snu7bfxoe8irrm2PZo9+d2K8Url4um/BnaY+GDnC6RyubSWx1A4iq/A5XK5MOEBbCt
7Y1HF4brFmR4Ko2JaD4FkYJl7lpn7fpu5VlbS1v+TTvNxorgANMw7uVWwTHyskwITDvPwQZ6xhhp
D40E3wiBovxF3ym/P3wxZIbPrHM6z/EfhP5rzuc6+w66mKULmTQzSDnOEfrRsKnrAKFTXIZqWzu8
YHQSzYq7ggf1QfktNYkBuk1r+jylm4F+GuuLapkkx4nBSUjGz4bGZjrI0iBOU/piCMtUPbrWAD9i
lvoxeTYnXYtwUR5NzTqULAl5PYrSfL4SgSRNgNLZBCYuWbc3dnAlWWzZLCS2MdL4pkGWLa0g53V6
WI21+ZViFVuPf1pg0OwsR3yj/b8IdkOIRt1T420RP5ygwLnelhOgc/j8/whzDuxtAVaknC4+N2X3
PcyIYw5cSnBTmQgJVqzvkgUXKY80bsKyYT4I2upFvpqLSIQM93xhfRw5yqKj/fFcaFBUMOOL+WK2
suVMXxm8hXI3uJfa/te1SqnMC2EKIe6Rq2T/ivuIkMZ0dXmjMwhz2Q6UhWzpyX3oRC2dSWNdEvSC
qLpWktMXBWUYYaURKUtHdo0FlAhJcmN99kJZokA98YNSj/2JSrzyUsFmKysXs7EyDCtCwhPL3l+L
8Si5zl5P8XY4aDOy2mEVGYI431HhH2vEbPiy9nheCey2vKyxRSRPL4l9yfzQwkx5w/yYbuM2oRCh
6xnIBfxhF058OcFaZiiw2jLAcaTDj+VwVCEHIlWvXp8CaqMQeSXk0fIoW/Y0n7X2lAaMUAgQ8lWl
jCXVjgkvr0wFJvngZLgxya3KyAqU0ufg4nAdKxlxv6ZJou3z+L6g/BQDxD0DfqTOjvHFlOUU8pMo
oF40kUp+jWFNMj/J0gRyYgXjWkeTLn7ZzyDpJ7xda5ur9nVk9A5PqgBuN4UoXaoPu3hwNeCmTDIa
Gj2Fz7ZK90WE4rf1sFTDgf1NLyV/PZbnoK5hfMZWjvqBo2Mk6/jEXgrIa7dTl16bACTIMQ+Vk5fI
OGUesRbQo9Bp8dyvxLsxxS13GNYk3gbnAXURve3OChEEte9NoQl2Ax5P10jtijohz4zO3yslXaHz
ils9CPgCcuwlOh8yH5g8+4HmE1Pda/uGgnLOOV3EPjmMP857eXrK6AQfHurd3nXjgw13QiBFeLGW
tXLWmamwkiHghDS4NU6lu/p65J4nWPVma5vwlgU85rQkoAncGLH1WKUwwC6kX33dPQQeDuXb1d34
TtQrWPOliOuOmz5/HcEClZydDtd96CF8B2cZXu5eBTdrZZpTiuVcxCp5Eir4qUkCyiXP5ZZcxXJ+
31huI6ajqowATlH599sbld/X5D3cRAe/qo+4H+RCRnmJwxEV/aOSINIefrQEj01pAQAQUuH/PFBH
LAASEGcrE5S5HSE4V7fvjKyl6IZkRsH/D03sVaxIR/UJpV9tQQNhPfu58Ln7o+UUFP47zgAxErHx
NuuY4fmiVjYd6xTRf3W19Ic9Hz+6dNlVrrsgZlnZKWLfmMNfzdAZo3fLH0wdw46DcuZMP1H+A9HM
ZIxuxWgjHCCAUQYHiqnOs2v/pKW+ExXZA4TvbQ/Acbs4/FCua0QJMuY20IZlZ08sqH1VMloIhXQE
fW4793yJkGiI73CU/H6dXSertXqwQYSFkd/kgtj+udA9JQ56h5bwE+SH/Uyb6pk3O1bKT3hz2xqF
rmzQSn5uir0KQHZRWAgI4GlDQ242sGmmc4kvAEhOw5SIaOdUgGrKze62IxfVDdokIjCj8kwfEO6g
En6axqazqYmooRENlcxb2CarTgkJrbOiI3YrTxYZQsaQ7YPZjM3XYQafwVOgcS7IPHZ9B481SXRa
mYgp5hFgrAZGr2asHELA73i0vqu6GVND4jll1Q2LDNTYBTJlmLEGQPbjZcw0495TCGFIqpiA46Di
RHMDeQbqt2rrCO9LDxJrxO7uoiR4NJJdmd2q92utkUwFrkP5iMBYdUmyjGKacul1GoRt6Hj/hodP
MIs5xxS5PjQE4U0SbGEVmKGQd+mvs523W+djWURIaH1voPe/Qb1bB/Rw2ToG4lERKvSGtkSeMA4Z
j0SHA7z5GllsOCuNjMQ+qC7ViwakMrCwvwg0AvTRhtqdSVmqc43qt96VuxeYpsvGJtdxGgBcRqh0
VrDdCfBiOe/sE4qwl86D4KRQyT6WX661VyOVqLPbp4nBnPxtiPWMW87hCe99vQEoKZMOqEk3VTca
oa3bQeGPgbvSnLPZjTqe7dtEJst+40nlwQdJRe3NX1ltXAGhDnjzC978XGyeUm6QuNbu9WMA5VVx
YOZ3qWYkSRmv7CgSLC6vMTZvTWiDpTNWwqb8bNpOIzxNs1O7CcCWSNO6GMUD3P+YoJDPWIO4947K
h6iZzuhJ7sfBK1rRXurAVxN4vd9VDuTGuTd7hI334Vx+DJ+Wh1Y3prtYrJcvw6YY0bQdD5CVe4nA
xd/VAHekSL5xQzH3RzVvpquB3SmZw+zmMQkzLN8fsAP1KrzVRTgzzKdSGSzk1qgrPanIu5tz4U8h
k2oVZ9rh6AUbiROsZaVCiOBSDb/hfCm7aTrbQTsEqS0lUI0nRtPVUsYt0VbA14lDhdxJ7UmV5r6y
y1/OpIW8w6bQcCf3aH+d5AlA8uxCdRcZSp9AtOZ5hf+rPv9qMTssoG86cbftZmmvY6fTa1Q9BrTh
tiz7AXTzvgdt+ROvxh5jM156Ri0YgEdybVYXPLDbGT7dFCHi8ANW0SBWFEbf65Eoeh8uj0o2O/7a
zPesXJbrrmUQhqqTLk9B+qEM1Z/fRCW3KN1a25AH6PKmTelmjj7zJNmjYPF3c8ovjlmsQBFwT7fV
AGkUOIAyHYIHaQ6D5Eq+wkvfdeCIIcytIT1h8Qk4cGBtcxHBxy6CtkF5vUBF+1HfComh9NZBaeOS
8nObt54OtbakwV3/EsUsS+EUmkey0JA+3SsDg4RVU72T2KSI47TRjD435hXW3KHgyydws1BuxK9F
ke/S9stfx0eSMQbb19k0OvfVO+KVfndIxyv0G58XusAwcXKNo60bKEKFX7t5Z6oYBEupHIks6gkr
2PUiiXb7zv7u2gKbUHnT6hgxuqVYu/FZYvmsn+TgfrAfDLpJOO0p9B5acM1jedtBsxX1Bzc4kckg
5kpZqrmAndqyrXWC1dCT+kV+FjwA5BAGuR+9fRAwD3nbPn+fUj5z3KA4/O08D6p+zkIYm78B1tbn
4mDSTsfcCXUEm14aWd6DJW5twttYElvo6iu1aS76wms06vEvbdWsu3sW6rXbp0iIYgXzRjyFOzR+
9f0P42foa2MLd/GSF6s1rco5h+eB8FeS2oPw5OY+2Z+T9flTwiVd3JKsZNZrfPGhXqM+HLltp6rc
tZoLTxmFcME8t/zWWfBTJJmkKP/W5nVzhoLzhMYGl3n0rWxAxXAlwkob8Iphq3griwFARYB5KPKz
W/zJ6aZ1z8u1nlUmpw4u2nOYgqqkBajrhpK6xFr7n8oO/XDVnPsR5cSm+dwO2f0raxLY9RyuaGCV
To3MjcIdwAyO759pmvvGpC0Xu3EoYyc6xeoTV//f6s6hrkspLfeKuO4/5bbFzxXzwgQx050TkRen
TxaZDCCPfPj8LBxQ5OY7sdcJTA/hnIrNklVJjCnoi56TlOV6pKi3fCcAC790y8+/nUsW2RKZAZY4
7tpRKLTkvXiAS/SIBPAoo2J6mMAcEwmpSOPDc+34D+wQ73ru3gUhxs60m9WX3FACFZCFJcDQl47x
JxK4f+TgD+btH3xQQoPxtoQ2lE96ercw2znqGjQLi4mmV91qDF3MBQL8nrtl1OwoSKPKfFqGswXu
c3PE+sRscsWyn3VNIQ8YYG+VCdYPA49nFO5iAIOKtu5rl34waS2Ivd+tpV/1YkzOMLcfwGXYxHur
Lsp3pZhm2kOKovzMXah/Ri5ekJ+06Zm1zv2qS7nrMf+ncuttRJhcTZJ8An3sls7RBSl0QIEW8l7I
1wUu76MO7vTooHda09Yi4xJPwtlru7yrTsirNvaZB6lxdKtvMPFdvKXvLuCOugZwl1BBk3IC3hqx
UJ9GNJbchRE5qoldn6ZgCd4rx8Ceh5YU5/P56lAAW/gyqJv+xq3OqGUm69o9obyjpdIc84TkqsFB
pXEuGkXNZhmPdiIV321nz0QzKXQeI9jrE2PP82Rzpw+cTEuOeDRQI/qlLM0wZpnN941lvn2yA7oj
1ilJoMvxeZEk1eTWO6QHtgb+CGTcDA1meJOK5S3vvSOrmP7CIanGkJmaHbuMMbv207oba5Bhg/CT
K5D9KSDtAaVMDWULG6lbM1TQ0D1qiXtbfMyg/6ZlR6kQathwqGpQbbrfoIZswQ86ioU6ptdvaBGi
fk7of/3Nxzo/m9RvZnVkELu3k/DIDlWH8SbkG9x45uwsL2jeWeofQ/MvNXxFVfYewNE2fLVPpN1o
eiEIjHrmscbB/GYF+9xKweml4jSNyjDN9MOl+mw/ZYjB0O6C+dDwxt6YrwIKbWWZCAluPD+ws43y
JoU7VeWntpiG3OpnKsPNe6pAmCkR8pDb44YyIjA8AxVOMUcGdoGuMJcBL6zafXC7vYA/qYYLri72
MaBABbzXGC7vccJONhcpv2Le5A7HQFmuPvQjPT1Dh9EX5CAjch7sgOXVDa3a6MIrOoAS1ojbV+e+
ZXxcWMiPfIO0fMMo4CooNA7ucKvDuGLPvq4gz4a2wSQo2leYibBKE587HVaQWSDhO3cLggK/Um44
xvXUwAQIF5WtA9di2sZKZ29xMM96pCYVjAYFPESQIP1CMqxJ4S6dfrHQT7f2NmCA7gTOwPV8J915
Dym1mg1HSwZk/5dBtrOarP8UV4t137xqifbtbVk79XL+lOmGGmXqkIIv2u8Ho1btXASysz1VfV6L
8Qhmw/WQopAQUfOAsnhm3l0J8/VeObs/YAH7Lql0917Kv6X8Z7VxI8FO/k7FBs4BdXncAZRSj1Y2
J8USjBudwEQTsYUF0w5CIJ0PkwAclUmH3VShMzOjYgVIxacD2cVx5jsYJEEL8bwy2JnGxFDQAw0a
R5tZ3e1BnWO1kdV4ELFfeCAf0vrnz82Bj2Ew1hGdN8Ssepn7o0X3x3JWduWfSIGQ4P9M50gLPXUD
CDI/xMuiWNx2P4ovNgdvhAh1e+Q6im0K+xUOlrGQWGqRlDli2ukrPl7DBBa278QDfbTuUL3NEfTb
/J9lthl6sQgbqFQW43KCSI0oN649duqZeLAjXHGvzgMS7gJrbrYe+YaKMmeHn+1oSRnAoeSDd3OA
y9HlWk7xRZgAIcbyIXnBvZDhH0ALCzwpKcxgwTQw7Kz+p+Z7ogGHh5vRj9qrE+13++Dt+spV6+ST
vmZY213fQUXWnVT1tOGw+mqaVvYTjOSvgqRbmG9C5sA7RrhPYkuGRxc4nu2x09DFlhUF8a0aFU1E
6Wo/PEnkWms5lbTwELbDRVRfQKHUJHbxZ9uYtWNB8Vfi3Z/oU1OxANlE1frk8l0navMF0Z2gjc2H
i11gznx87EZlGfmsDxBYW9ANyCOyKqnUPWMku96lQyXdle08eS15zPu2XM/1EEOEQ9GIRE7gxiyr
etNQc6AK4eJsAnDBTTBrvts4E9EklF3XB5zEYBHd8r2Cj5P9zmzGLRggu2XY4Ru75uQeaiKK+Ky3
xQRtV8jTHe3MYCdZDAKYxXszR5RieO3HBw7XLX7EGJliCdzIMjwAokLCfA6UeuG8uM7SsLoI4RQ8
N+Ydq1xq8orGpHHTMHjOKGu1P5rHgRRiCFJoelCxJqu5FXlFtW75/RGUYtc5ILW/I+E19/p5bUPp
cRk/4O/j7HrrVn3P41mLTsrPlYLTwEyND9je8tqvn30cyS0xWapLs9TMoCtf8KRtMCD9wlZDX+Ip
bOhspLJVDL29yOKEstaURcELbY2xJjHBabt/VYXRi/PnFgZzJX6RzGdDgGZIwMw39+r+Oik9HLVA
eLl+0uZ57AnQNdKdRZubifukKAfLOAWRTQeVk7mVUxrJUIpiRTyjrpZ9GPHVp2FFtV/UQXAgOycd
d+ZvjALl+dys8swaGLqS6VajdbMfXVpyv0ihPUyMOaPgxnHb2fuw6vaoDFh77Zne21R//TnmOv8B
7tWC572iuJWR1Ti6OPB1qJR29/zzvKpQrCPt+N+OILEnRejcZ2/Nz3/v7HepbwU2JkIeTxjGH0Dk
vXQPzkaLlNASRWHIG8UuXIbAug/QkkX+bMnz+Q+3ooi5FcdIjyM5TCFSXPKuhPxdNRTPHrRpviIE
6qxcq+z9QzQYMUWPedk0/7UcMAybaogrY/zWtscn3OkJ8bI0KCRRS2jnidzJt5jJLSkqkzO0gDw2
sxViUgH3YVmHRPT/GRxfffLxv3BhxryFsalmPkEpD9TwGwP2mZ2s4S5d7bvKvz1E4dbPmZMt8RUE
Uq0BtGMZOWNsN1b1IqU5b47GH0RK2UqrVCcFbrs0gh9mm+lLOzykQEqYx7SM0cxtmCerpy6PokRB
C9cnLHxFoL5HyAqO0W+zQg8687YmT9lZLxWKkmTUGQOCX7Crn+FdkkVMvg2ePA5bb9oTpY8cc6Z5
O3tiuP274+rfINd+VuJAXLP2DD9RJGZ/Exwd6cY2+kuknd9dVmduOitKaYiIOiJ9oAVQLj4Hy24Z
sBKUTP7l1xBakOVNfioeklqNFOe6JVb8IUyDcHKJG9tkfAwUVxym+H+acdeHM6iEzmNQLxlj2pTK
8LDg60vinSdxnNcvlbJ1OksRQZTlhBMMlnTdD5/50FfZEttH/pXGWGPRIRYGXdPqUBH5pffvocvf
MmL7Vy5Hw9o2xS32UTiyMtjsPogdUiICehzfXOL2Dqtu6Wgu+KaxFdB/6Yt8SO1sYr6ZplYwgnnc
B/hDX1iPOfepLVMGhglM1DcfvIR30i01EFX03Adq0p61c3IxQC2CEP+CuLm4aWZKMKDTfdT/3bxA
LXOyhoMl2KT4WqNM8TrxCKmFiWsaxtk4r/ojj4feI97VKbG6BHNBbn8Q4D2oC9D0OoYRXQkLwnLE
1b4Z4m2yfS6QHYUGJjc6nXO2Z4CQn8AO5r2ttNAF9GemAmt+8Y5ZEPhIY8DVs26onYFxl6kVSXDV
W9iSEkVYpc/w/+2z3npcLjLD30lm4tETCvZ35Nrr2XBYlQdmc8+c2JvHyVlaKahqtm8u9m6YxxJj
9JZNLY//QJEy47E1ZGwFAmVeri5XGHH4V9kfrVyOV7rMMK+ijoZPmaHrppA0DRg1/PQMLC6ecVFT
fGwEo6u4iUBZAx3XMhs3Ahlm2/aF1Zr6Ugk1YFqYcx6m2xgGfTw24wBR4liabYzQBtbgvWf4bLZq
e2K8UPGgn1eOkZ3y87AQ7COt1iqFvS8gHIzVhH7OvVCqewslErMIFmVy6NDb5TVqYk/5Pri8EteA
x87F5nKVPYFq9IsM/tDPYdwLOWZ8lW85UmWtrbciYEMlpFaE989smRacvxJ15o27FxuEF7h7VNr8
yqFSdlSYmRXtyuNjtxy5SfZHyVHOOw+VWAj5GwP15PWfeQ09MqdB1v1JmdKoQ3l6GxFLPc9ZB2NQ
W3bQG3SnL8eK3r/mjirNRrROqf8sSaca6rnAyy08zNkXc7ZJb6sY40WuJbLByup5JKCbkruwfW5O
XD76B5i4dERtRXpm/512nrz8Bt8Xv64Op52chmIPYti/DNfDReSa7o4QGG9xVMQW7GxWnQWQOYyq
SvdLq8i6Y7vkdLEkKi8yaghOuSB9ccFAPtLCQF8TJ5On+PcYMdWOwKT5993H3crbvEcwC5eYPGVR
wTgcak1Y7aVwUVUy0ZWn9PTbJ/FzWzSUmLGu5QAdUa/jxKnPQHnkOTosKb3+MGEK1jt0GdGZXCxK
8YjVNUWxj/j1ko1wKhICsEqCMojbB7MdvES9W7fQB80R6K2YXl8YMsf+LY3mQzu8Jy2xVWGEZbcc
RWwcST/3kA91esf0ZVxnR2+R0J5iqF6DW4aM4DuOPe4IzRr4m7uH4gfGRHjqZBZULW0IeR9RPH1T
6GKHqF28R+fjWskksg2mobDbcO1B3crwBG4+zlKqzHldXUqOMi9ZIwnHtVKRkr0c5D38rOASvAwe
5ZkcBGNwrsEQLhgU1ZoSVJjKajJUPxW5QbleNerUD/jPcXhonZxY0zrSyEb4g7lfEFu8LwCu2zkn
+xecX/Upv5bRB71IpjaOCttGU08A79YtAuXTeQFlyPadY0gs32Hx5KKXdIG55QAxTCno46LMLo8F
NRb3jIKxaOFpjJ2qeh5IjVL4VShzWtGCgAjB8XeEg1oL5PilU66viXvfNwiF4Y/wpsn8jUIIf+Z1
ZgmWds24j8Y0UvhXu3ku+Ww/Js4lxdihoHvtL9SHLQOgRcWCPCgzGk3Lrd/yKKz6DtteRtxdczeD
NYOWzHE4doXPkTZfv6d3/QoiKsy5FB1SR+tVNwXI2IYVVEU5NBdh3HcUG0uT1zpO0lC3YFkNcyCH
9htHkMbYbS1jviv4tc63oM26wGRXJHUhl1NzqWAZpQyRRONRvMuoDimyMcfX3muQ7mziGAFqwVWr
Q2U3DLEcI4jHqRMxJZRmM+NZKjed7H8yCJhsm31v8C+ZWwBzUWWffkWtmtuMZSWrTY1AHAUBltkP
YqlMfVcKufeDNkhCd7Zkz4HZLIMswz2m9+t0dBHaKdrO0joiS1F4oYyYgta0KA51hd5mCTUHwj07
8UPYA0HsDpb5frAIi1yPnzx9yA4RNMacS00U2EDSVzjuEh5x3elcMJoll3tBWcrm+YQH0leeGxMl
7FzE/t+zQnNyTCZ95WIs8a3lzWyq7Tt9jmieRHlb2cA8ntmHPhYFARJnj8GhHZbw/s65nKHz4v7O
E57u/2CL3c/ucjNwlkGRaqKPvUDM95Gk1xb+m3XZ0T151S0DQaL8B/cOi90Qvuckjx9L5XmNl3Zv
bEGOKTlpH49K6uBFNZXpjkvTfYy6NaHAS0OQkHhHFCzIPqKLsbu6gNZ2zYW+/jLHd3W70yjrTs95
dAbB/RD91gdohNgGexKXeI6/s077nlYQ4I02w4vAyWjfXcwsP+u2k/UPuJ0MmqB/TcuqDNaXnB02
ikhYs4PfeAK0sEY8mldYTgpBVMqSAqhNQxauqd4yqX9EvfzyG6e1PYycVF2lbDecZHGD9V99psRx
T3o1GlYxXFcP7j+TeR9mCxkh+5YgzZ51N2QyaFt3vZnvVT/x85g8dhPzfwPdavAtkwy6sGyOI7yk
/zGV2Vepe6CWQJXK8PugV+6uXJMF8SIDxhRIS2KVnM/sJtqR9zucLxFFAmCibVONmmwjH1XQHDuu
dozw6PFfgg0HkNhizeq3lICMcBH6hiDuySHJOR06ePCR6yQnf8QlxOy3JDcfgi7cGlFCGU04OiHz
P2wLGejM/wltKeGJ+yNmJI4vQy3B7to9L8FNLCz83UPjstwuig4W3sbN4aw6A3vbSDmeVvoRHVJ9
OPsU4MR4thndt7yWe9xm2el5IW9lU8rD1dDT5f2QZqGvzZ/inio3X3oMuvACxfXy0Qj3IAmSmd/v
QNVKSgBjJOXGPMMyC6j6s/MeUcqnXwRWV2Xd+IL8PVfPlu1BQGiDd7MgdrHGFBSjCWmACUERIeN5
NGwNjg+jxIlaRHq2SU6KqnQlI9j/qKwouXB+eRQ2/JqM6qic/jR4s/8W9+5bJjVF3V68fRaLM9K1
i2VKZY1Gb8QPtm16A3M1QmF2NjDwviqvOK9doZ/PpgottaliHd5NyO/Y8/bgSepeApPQy8q3TAfE
H6Ipzkzfiwhtjl9X+t14EGLG4qDW7tQN3E85625uucx254W0Ql1NmFNhCVjKyORCa3tWM01RcGJV
AKEkCFbC8mlFip0fFC799s6H6kcAEGipY5c17uKs7VwbMjnMDmmscz1684MajPD6xrzqygD189tn
EfVT3rvRY793XUoBtuqZWTGaJtHPzbVGbOGI0dSPFuPtJxjO74bYGtgUW96WwDURdYa19xfhi+tz
NAbMJ9eHFfAAALSJ4L6prOLOlVtVqGpRmXYvNVzhhfNBXPvPHmIa8jr0OR75Wqs10gveLdtPyihQ
c6kZh/3R9CYJmX6bzK12ZBnDIoleJWUeckObxyzaKG50r4KmiUAjS4zFTR0WYgdjTHS0P+Mzw82y
RS0Clm3F+nZcy8wltUCcLxuJOynNKbV8httle9Ny9V6rx55DwHUcssUL74vFmZ0pklRq5Zg6R/KZ
JbWJi0AphXWXW4KXED1s0G+3eeyoqT3iyVE45sItRcvBOd5fB6HXGTvEms7G24KOTrcv8xNIR4iy
pDBOVWPChgeqO+iMVThS0TETSiyLpfeXnCyq/W4V//Y0lONROv3+qhNhTKdMkO13jftjeOlyvOS1
FD7hvLGfYRCjhw15VpHG54WFto6EV+CpaxVhAgV+VFxOc209SQcDuA4KjsdSGhVwTSoeP29ppkIl
MWNDJ93rN3UefQEQ/b3bXwRFRuLyWkSDJ8E8QNFbEn7nRIrK3n9Xx6HhpHXskYtIRWGoCiDEYUqp
jYLS3LzHtqxQZ0Lby3oBELTw/eDylqeaZS8Z01lCxrn9V78NrdRoxHJF7/j/qKgH3/L30YWwjoiD
cFdLb9jbVWfoMne48mVzRXknDAFwETi18bHAasM8azVd/P+YrWWwy2GSIa1NLsKFUzt88NBe7OPL
OdJRgHWgnNwf3GXVjfUXSMv2NOOfKsIdj3GnCNHxSR0LUiebBQnlNe/qw6PdeKzotWZervqCYwTC
Yz19/oVEgVbzV2+y2xWR08x78XjdXAnSCR9aPzaB4RgyjBsP1cY/Gwibj5LUPBl45XNwCHtX2BgN
wWa4rgTpnJd7TdsnZh6XwTeoBVfo93UK+BEKIMT/tIjUYudyG7Upc9M8IczZS6N/ml3DNBcjGzMY
aXD+LwYeAMmaeHEsXOaiH/IZHgsgzjp1NCuwqF0LJPY5X8C6JOnMW9yw41zzFbPogS7r5aKNu/p7
sgFjxBXE2LWbNKRRVAJrVG8EgEYbkszGCaH05jAlaEUSbayCJI9aTdZTV9H+Vnz9oKHbIevDK4qj
tfiyqOm2nV2HYthazfG+j9uqdJz+5o0vNpdZ901oBcgOmVJa4yaEEVPo9Fguf3z7dRpVcHiEkQqo
OW2knN6+sGdUqJjZiQ4AKuhwg0OKS8mjH8U8c2fFd40oxdEkt8AKVqAhwZ1tzrEXrke5SBzHnIuH
QA6ZPfbPxReFaTcBhw4656X1Kau5RxO4t2t2vU4nscqcIitOjrp+p+GDKRknw7mNVpJ5M35y6uq5
iq2QhP+/3g3d9h0HWUVeKG+IkGrjEJrc8zCIGlIpgTv7gyYELlclVsnJTHUxO9vMA7SdHEO/vo29
T1UqYFvrlSYE0uLo+FuZInPaskHg2yktu+QC0BOgSgF7cFeKeYIt15ETZKQcLhVnG28hOH3kZNa1
t84BwvqWm7q8wfEtS43aOk8p2n8sBgMmUZiX9ml4UfDKJzGxGnHFtK6EQKK8cGgC7O6r8hEF7CDO
D992Fb/1JNNLrqHM4TryV8KuFTvw7DD2kMMj8rPEJUVNQ9FNVbC9wB37+GWJrcifi5vEaobbvt2w
5PoE5KciXvNaxl8fZ90HKiUY5QrHaCDvt82LCsHdBQgp7pWJMphrUGFPU7m3HPOFIrNFiRw0fRfa
UZYTDVA96nUgs6XPCAL50dWxPPZtHFjfFHy+ujQxv9bf0rgIwH+l1gNiONcGp4RhsHElAS03GS1j
yobmYjdpJbf0ve3i6NgINc6K5WjC6K+dRy57bGpW7fMRFvZnzb1VI5Bk+0EF/dh4unIHY91K/5Zt
egdgzFZnzFZMkNbco9souh7hB3nbSTPgOaAyNuSmm+UTF5iB96ayYYi3n3ouwB0FqAngpiOQ9PBd
1gl7SIFkOiMuLb8llwm4hLexi8Gzax6TPzOaXU0NLJUz9hkm1YUIrbEnRL+Z5yq1UDN/+XXZHd/w
PlPDgzeWXj/Bm6kciZWpKvCVt/Viw5SV4eE5oXRiexOLbhw3CKw0Bw5SuTJoTPQx36uKCQavWgl5
CpesUxYuHNfeVJWTKRXw/zqXWcthare9XFVD6xhGyqjctL39UEYfjW+Y7IdkJqI1ObNGEqNncNd/
os5fRtkIXlX1dTfLCesoFGVjxksJWZ7wKsX1E+UxcireinLIhYJ5eKdDBo+P1X53nRqvK4OC5j5Y
W9m4ane5smXZRdneG6YM/MKav3O+0lL+3IxkatDu1YUZgzko3bn1+Uy5ovF4+N/pZwlLVDziES3M
P1i1xOojdpLra63l22NLdV6EK0YrVSxyFmkRKTXqLAn47BI//pdQLFaS/0jUVYjRdy4ZBFr+P9xY
D4XJdeDjhYgbRp2/AKVth32CV/1BbMc/Zy3jzideuY+kPGP7ugcowCbhNFV3B/J/ktAFWfZ1+por
Yve7zZXBSk5/dq7CUgCg7pkcqc2hcekTiUl0P3CWk4dZixsuwlnsSjPwP+2I0PDSqSHH+RdOVNlb
/oEHYz7g3yrAt1jJ5A/Ew/6CUKsdGEVrHsd6ckcKjba9QNgMSUbtfsJ0ZR3Vi6dbScrt1zbJ2EO/
8osmaPH9cKuT9RrPn75JKYHRC9uNmOekrpin+DwUsAivaw6vZx9ZXDfYTxihaepNdEFJCAhmMnqE
WeLxIhLcYlTEtVVaB9biZCMa0Ulf0P39YZffMXhUcP3kOYxgji0awYNUmfDRhh4vllwGChBml4i6
5dQdsGuMi8Ygr7ZeXsyZGF3KD6AyB6AnzkGIKgyErC0ZynrZP4CtMOTVj2BvKCtSsIXeSO4tGMr9
eFlgNN9ksDox2taD0ptlKEJXfh3uwZXhTHCjTQnATWfLs6PxbroT3cb7UnlVcS+t44zJoq12sFyg
yShgLdtNICrioOLzZCrGtvw/PHs5VnPOLT+FDlR5cHB6KQ0h2Z0HQOCPg/L5j935SMwi/SFkWl5E
UBffIVnTStnqkEYzMs/WI5e6JOGGFdTfdP/hg6mgTerAXgJY7X8Hl1yPuaDC5WQr89zF9FLLiCTr
drVdRgDZSa5/n2xhW0E6HjMx6x0E0jjbXDjkQqGvZXc68sHJ8MPzwIHfd95hRFcdAAXln5Gyp9is
co9tCLlkSVVsV79EdNOhF4YKgBSQMHO3AyU3aDatAIydTB6p5Ekl574gBsHA3LqdbPBi2k4K7fn7
iZHd+PD3ii6+3wJJ0/pj08gUOv1j6M9EpjNPAlfIQSAhjxvLQcHSmKnvCbU+NyFRbi6IdyJ0Eniy
/nLo8j+Q/AZnTauteYqFO4/FGjcEws2/h33UOIB/E8AKMnVTRdTA3el0DPvXX4vyfsNg2c79fYRo
OmHQCdkWrazK3hdVJfGRiPD3N8lNolBXm0Al7WnzrFaHz+QrloPXSbBfEeDq+90mxkn07C3VY+PK
nN2I9liHrztP53fk6cgh58Cj/nxh5D2+FRtAaNgY9jGELW779XWs1O1ALHetBdOtIcQ/FkSauGaQ
pUzWR51Cwo6aTVH4I0UUfoQ+NvMEsadx3wJ3QaV5L0a7QFj6LMRXUoLS4Jbh3q/hJc7r1HhPMwQu
RpcGmj0rO//UMapuVK7UpUGtTZuxWAEbPGYeHUmm7Xp/EzNSYy075Pb33J7MBuhRKd3/lNJupe07
YO4Ka89vgYirOW72/CvYyAB9zycQqSGWkP2PADjn+fWJpOsXIvpFvxkBdu6S4yy7NyyS26x9/JBA
r3suyEM2tpPMmGtqAjeyvlMm0MJmhFhsfZzWrS15qhSDi8iTUPUIlcEnGhF4nW81jbk+ALLjTRVB
+MNU6wOglaTJnjhSQYbLpIPz/NY6RjDYSWtiyGv5+LTy4GhBxvX2mTbZPrX3/ybnBsguzmbM60P7
KXa3jihoMbOu9PUBzmOlaZcceV3oZF8nSrAi2o+U4SUxifc0Eu1BnND0Bh4Vz0fAyoKiGNVQzODB
MgCxbA0SxL00N+xm8PNbRqNJ98H/aWwwksmL71KzkNvQwk1GLx/pV92Tj9he4Jj5QAzWM02hzDe4
8qXm+yiYYv2Ub/597NZmeZyo7CR08Gu6Upm8hiymtmIgGV8N2RzqdSzWEKkobUie32uoIT0v7uQQ
QyKOvQDwEai7+nCHJPdO08RBoPK6r0P8ZVNlCexuNxuhT4ZqGH+67BBuIwTkI46F863vCoOhe2Hp
BgTDTJ9k140wHJdFouKhnVrZZ0ouTfu4kcod880U8MCKszx6orj4yjmgFAnekmrhTj7LTYz8e0x5
zolSc5Z3DrYx7/pk4uQj0N4QapVhHKQvMSe0PzIZrLNaJT0gTUZ83kswAOkuHLVpr3/WU5ts3wRv
QgOuuKK4r8MgkL2ZLXXJBFoIYb1K1uQobRo4GfKvX8qagHfqXwgJ6b1dgWunTeCQ8lVaA+Vp+9lM
COUo1jjCPZb9Ah8DndJ3aktUFHuPGwmDAXYfEbvKX4r2l5MgwE+xPcRZrw1499U6B70wnp2pbH7K
yQpC8TL2Y86nxaGSHDGr1FfjSGxQRVutz4R0xLuswnGCvOc5m5ljwXiC85n8wmfgtbmBwQuc16tT
kheN8Zem2B9Sm4yXj9HEqAWVkwTLqbcolEpt2STf9MsobNCZyJ1jG98YL+2xiJPZkr3Kvu93GdIg
npy2cv8gTN6cCagpa1P8PN71fei6ALSvdU9uUvx2SF1nxEKwaMzZrISau94gbPsDh+PIUqVfLt1+
eBsQuAHbE52QkiS1Bg/F12yD30HHuK8gtW7vVSYrJ50t5JEpJS97dr85fsHtyr49wTeFJJQmyAIP
DJ5R7qX906OZLUGTltCcUkdOQ6TiAYKaobSeGQaqL2QtoHBYVGapdrXykcCyZd3EmwLR0fU7i7ol
cvHgrt8ckl2HPK7VIKZEQmS+ArRNN9E+30dwD0LaZNFvUxYOqPzgKSHjhJqUE3mWT/uHiBS8s289
BzLfihCC964GS3ecceHhe22e+L8iqg3D8PXloz9gl1HnhmbEDZtZ9c52lSRRiXlgk86+TzYpDR7W
BDzpS6Sq9VnUzQY4jtL90Cl/fmEcSieiWxpggTAXYEhSQ4GdYHkavyZvnXjmH/MoxHMksIob1Jbq
eVdsjmY7o8H3GHkUaIMer42hBPyLSp+BjQxl/32IugTjswiu0suH0Qkqvq3MM5wytsJwllIBFfd5
uztKzDZMQ2MdWwDAeNHK+u38fjsg2QOb45drWCPVYpWyRROkC3eUhBH7Sr37JxvvX9UR5XbsWRt9
KcxyaijKXEX5Ae1q0SEIgnMW/+ZggJ4KXlqwojR/B+zoWOYNyD2cy2rNHNeI5vstPSYsI4zPd3CX
GExX7gIX0j+e7FAAIXQ2S22UYNRaFJA5eWkVKa89qfAPY9asV+GXiGlaAWZG3HwYwQZ2eEmv8jJy
Pg8NjQ8SRC7/O9711ZqPO1Tbwvnc85slwxDuX+dt7jjeMazQxroLFNPRHx2ci9tBp7cUqLyN2Lsn
kzXHvjOGeZrcAnqr3uQropKlAneaqkJAr7aKoFxpN7yLIJsN8OeZx9d2vfa0YpnUkbfymGODzZqg
8opgd55PnGCw9q2itfw8jQ9vJNycMLifUhxSkTylSKZQdQpKVD4C4DKOyr5z6HnfPbDK7fxYV/7u
1peaiG4ruUrua761FXRhaX3OH3y8XPWAjhDJ2GInFfdh4+1M5JfrSKrLcFjkHglUkuw4awZyqiVz
JyBM78JI0qwAdpdoKmG9yWmxX0KNlU65lAyd14gtmEDpTM4gI1yITKcHArDJ+5VP81VnhYKCThbT
u6jBPDBxwwM61lI1gluEH+nMdNM0bpckWiyFbZh4Y4APn0EqOAzu0RYQbAq7zCLWBTn0cjt3ANEf
QyN7D63zU6Xmz8SUl0qpEcFUYRDt0caMjTR+0jQ0PYmm7W1QJkmKTKPeCFiJ6IqpNJOhz+XLx52i
BbHr8SGozA1wjQAQZnavb+vhQi1ZMqFivP899u+kWYi1zE7MTdm4n8E+jdVs6jkECi4aK5EeUXGX
PpAbuzkctJiISDHZFc1h/4kWkmHuJI9ba/HfOYuC2uk97cRM8c17rXWlgCX4imm19SowWsoecgYx
vwS33GFvNkt2C4mQLiCVOmaA3f6Oz4uE9qGLRiA4b7cS+KCahIidCfV4Zjfm0Lu54z751FGpnvVQ
qZkLlrRd9GrTwBwxk/YWn/VF98itukl6H7f7cb+sQugfKYQxyMKdE3dUq+3tYfbsuor9xgQTTvns
vs0d37XKz0hLyGbPNoqd3r+QNPjfHswTWhLADPNFG4aqd3fOve7ZeTzNUEWed8vxQivxfjrmIRcL
T/SOsWsgzzJQRy5wyH2fhgrspuGPmfjCV+lRpvd7XTjMK8Ll8JAp1zJeSO42L7W4uLNKBWOuneZj
R0xCyEk7KXbg9xpWWH+SIsYWmIfdnHW8nuF5R+gugUDfH+tMsm4TUz+0GdLcK1Btiyz0ZDMWcSMQ
8betPIVuzPINslu2bPJqSKo/HJnKM5G5pYP6GR9FvOFE/15GG2bby6LYccZl7YXcHiY/1q9uRRwN
cNBZB6nC26641YDDVdJa+B/SAYaAROHOkmYzHgprWNgAGLTovFp0jcTDv4ED8xQZZAxGCSHZ598s
K3a0RJARBHjwCzoc3hoqnVA6577RVb91EyBMHUk1nrww0/j+lNNr0J7qfM8FOx0qjDBmWBzlZg9x
eqS9FdyOZcA84BT+JN20D9UHNe8j2L2MFjyxW3wBiS0ZWqNgle3o2MOz0WICkLiXMNUtjsVhUZEt
Sp1XythesgJ81+lcdq55U7CdXYu7+2vhHN384xHWUfcMtyggVLDcnratFfie5zs7WuF2sPkZmOaJ
X9DxrH+o9fi602qe0vQjvnlZEXfXydCwUDmnZKx2JwsU58wsn8RVCoEkurt2hXIaECn+QeESnGbI
sKeuQvcWrMoHmJ3UxF7PcLJBEyn0lcQ26fKYC/AFVhidMBgkx/nh17SSPNpWf0THCocMUJJDKqfO
D/jZH+U0JNrnxqduo5a49IbYDAvimLHWe7/Gh4FJX6vMxztBrC30PkXKP3m0PTRe/JXmpEsJchxB
RhO8h4Z4zhR510TwctykJZ2qbGsKgLsh/qbItMPAonKyeUPfGR7DLH94tsii9t/Zf2OebovQgQzI
zbA9QDgAZ/yMa5yGFt7CWwLCMbJhVDuAWr6GheW/xst+bUK1MfCt2EvYR/bwrE9ZyLzSrnl+hFZG
hMDN3oPjjwWlpX05jlHNRCbnQ6fuyPxPsqP59MESGJKib4olujnJKejkrgYh2tUQye6Cp/6/rP7K
cbNbwKjpB1voaBRQ1U6fi8uW0XePknYj6rSSyQMC5Gz8HvHz2CSuEZmCfxPd1HSwuDcAfd0blLgB
1paUxqIcC6R+ztbi8vtp4IwC3A/r9/IQUtABa8t5wEgpJ9B1eWMiKbGGKT7nLUcBOYnHZXOn6DPy
VYGodyWsW1ea5pafCGw5jNt7aTd397XZcfQO6cCn0oiH0BLo3gYJjH3DDZmdl7jiag4NAirJN8Nz
YUCpslBfHMB1AB04PaISJJB8MAfl4ltj43Tt9ZazvTY1+ahC0Vcfa8HxjN+2F3cbSbwrpedun91c
bEyXgoDn9yPPCq658yYKjgeIiwCMFS6VwgRP/ZRUVEEaknvQrZDKNHwB0eWONYvEsAQ72hoM7N3E
lSdQbLtMUfBmKesMRbkO4eRP8TOL7n1R2B1Q6yAELTGM/4yvleOToKY9j0MbjFwXlCOdrwIwDHeG
4zxM40mObalQ3pbZmSrpn5mCWXAEbo5qrR3N4Z/H0ZelnXufi4zg7FuAFwcJMzGyy2wi9uqHEgcF
UBl5GNgxGtzoHqNwpQv9FYs+UCJ1KK8V/NN8Arv8XYvHT3gY8Amt8PcUyiKqAVXo1O5aQMX5+zbP
zYMdtyKRvuI57gFbKUtiHy2ONcEK7VXw3we4jmcdVVPMGDMMSP99TQoPQ1BmJzj05V7n2scOAnrh
wXq5ZSrHo2KWjFDU4w6tu2PFr8kYC+hY+Y+E3PZ88yvM2Mq5BtejsfhXYl0a2cxFO98voYR/Op79
NgvOcUDkBCkRz4z5iejUP0kIwt8wSujb+LILKj9cw3rwknvUjq+11baOrNDziwxwywCsJ6W9mcdr
mQ2BvGPhVWZjQk5KixzMZiWe967meBaApIDgH5RtZ4/ltLkDpwNz4tV2M6H3C6hVn0Yv/1Ftqn/c
1w/jHxZM6LEA58xZhTfF7VdPz/unrbA1Akm/8rG3e6KqZfOLxsbJeSB7Q7FBUtVK++o8ELEAAn6b
DKPxWRdljb6e1+poafUnb5jeQD/BhVTo+Bf7aowBeIrJUj0A7qOCrnCH6PussYZYlZ3OQU0zLV/z
ju83WxrOGtIvO+if4yNDDRWm7wODPRng4+fO71oA1cY61YWTyz4NYhzn6Uops0qUkfoLRWA6SBuq
JSGFr44szrNxsMyNQTHiZVh0gHaQXWgPabVypZXP8JHePvWmq/dAXEMS46bzXUILTs8UHsbAfcYN
lQu8YaWwXR/XScYkiOfD59gH/xsUa6uObkWhVLVAYAz5ZF3tAnmmg4fl/b713neZE/EtOIdgiwAm
ZlORh+RGdvhpxx9+ZobaRsvqY5cIF9ZA1rnKg+mHM57M1yx6piqWy32rsXOiiN8t1DFhl0Hr73OJ
dMqs+27Nrr8Iv3b1LGeAYhU5aOLYaZGNKUWYZRRqbimSEPsPa4Tn3lol+1gVDijh4UpKyIWf+UDK
IF+M7oeRyD4FuJQFdhZBQWTndjJfWLkUxsQ1+HnEj7yYqkFsx5WLtR/Nqta4Na7tuE96+zcxjhp2
r5CHPbtimrosKuDlQHK1qm7Jj5h3JEPEIQgNeD/1XC4DD9tLBB5K0bt4uMcnecNnQttKOxhiAcQj
d/om2movwAHSKPH62c04MyQeYcXmoS4xxnjPPPi4EfhGxqzdbih4rG9BAOKN8clGopf+8mgUNNxn
+HjH5NVyNfXdVdujK+97HaFEiIDtMVU0lfNlQB1HYtZclV79o/EKTnzxqbTD9/s16TrsiWEoB7Ir
3WEPZBBPjG+X0+M39hUeUs0n3bC6DaUEJcGmWIA+nAXoczWnaPMIaBWptKiMDadwsOx/yZeMJsgA
QgCA0NAdDI3V8XL8l5+jELIGf8nDXRXL0TZlbB2qdNu0DIolWU0GZhZTGfAm7ojkcyDIPlMsPwfA
7t42isVeNMwEzWL4kD+TQ1yWZvpK633F7qphhIS70ntrJITggUu79TzPP1NGUzejL8y2F8TxXikf
vl6ujfybuLrSvj+b+tuR8aHow5ak7d0+NdUnfoSemizAMxQjpr1/kggWedk2aeLrxq5j0MxYjIei
1D465OCQTAhYpklqIgoAFwsY4KRlqTg6NixIiHG6k8wBJvaUCcX0x4Mvb3C9DvliRMXhq5CL7oD+
2akZ8yjg6Na9pPubR8KncgZ/J6RpoSCfcmjVsxqP1XOyy2GeWeOpczpwh01jWVbLVsNhsgCivsem
gofSNULEfFh00dZDNai0oA6B9jHoEIYu/LblHTv+tzvoSYZr3n259QLZCy+4Eb0Dg+r4XqwaI5hk
igCdVC/MlNzCwlv8tZ2kBI/d5STrMMtUv0AcJnex4wOdC3qBhuE0xixL0eB7HfCiDXAytwN8Nztz
K3Ep7LW/7uZezmRTxXKH1sdcZ3YBN+p6pDVPaHIrNK0/iRkdoS8msfA66N8mzKE90EMQ6jgMzeQH
GEIBSB6qO9v8l8hBx4xHS48P97aG1JSJnCSAv8Y5z7ybcvZ3/X87jQnCm5mwSIBeFdV+IU+GhHga
GG54c/dte05/aoimavvuSi/PRqqVvlhl69IxZ+mFC0n8Cprn0EQh7auXeox1a99wSJLcpszc786i
QVfKh+vowxtbtQsWcuocfM9KDB3+fPEShkPkERBb7xlo/IMIcIU6VoXstR/l6y14e4O9eSgDwP21
q0QM7xdSQ7/U3CLCdt0VxXpn6UceCiZEdMRpGPQIw4ghSRWbgimHvTXr0YiNws9W/pSYPebRh4Mm
mFVn2YHnv5YCRxOzLATVETBvBZDwLoRVPRdtFm71yb8ASBPS4Z1xTKQlEj4cYYK6Kmu5+EN4pg7E
wtg5doOjfJCvcJ2ioIgbX50IAMmWfenZj/4KCKoN8FFMYF4jlSTMOK1WYWFxmYoK3A9EexEAqcvd
xqSu0VTYA8nCfDNKajiUSM1CXMmEkr4APZ3zjNBAwXFpE9MwdBdulGSJHKhNYPq0TY/2+gn/Qzpf
3i3fDu8EghhC+3ZNhU1vyWS/tipwBKWyJnKBkE7xsQpd9c1ThzFbzOjbAehSGGVjiq6m7pPNuDDd
0rOXLfma6zVWB0+2xuBv+3YTbqmDWPWKGZfYjmwlAyk/1lgI2CSRqcswixbBVeHQdITKuwYTiZmG
DS+Xao1JoK/xisUm/+wwIC3TuscM7KWGoZ1uRhEWd7Y3xOM8z3/qwpJ+ZgUpDqdwNZmehYQJ/JK5
Hycn+TC7Wb2PtFatB+P7/tWvUeS4oP3fUGNU7kUkpXf/pcHp9yUxWHfcpf8iV4quECs3Y++wmXyL
psPO6HJrYC50Jeqzffx75XSZx800zUt8Fv7rrTS0sjawVRVo/9oycBzddW0mCMGV/jT7HmSdb8nI
2jjoVIiX/lY2uw103z0sBV1Qg6I+wdBKxIj+ZzSN2upFI6DYlNX8e4PMPa/vxTM7erUXocWrY24q
4xEBtmmYNiMmld7IAUbfUy8U7NYPayYpoNfqChpHSaLFkOzb6P1tC3juakNmuF3m/J7u5Rt/Md5g
SQLqF8MvMWAExzWtOgawCMhwsQWigNyINpe8P1Ce5Ii4VIJvmodXpfq+hcYNVoTOcJJD6P4E0v52
Gv0j3x/0/AFdiEkO9OWz9rapDsd3+CcX1VJwUsf8W5wjxbM9J+Wb3LYNfgS5H028TrU3QoeM5X6n
JkAH5VVLGI3NRSzZn076ZxusmqqfuuomipV0mnfIJJguA05kd1Caagr10/8hwUkpR1OGb2q/M27t
NGtfRuifw3b8xVe09gVqYHcbp7gT5nQhEL1rsfLH4UVrqHTmQxFQe+fQVoBQid/9DO6sdp5Ur6AG
66i3NT32xY3VwFbTP6G0gwdvb4v4rS2P6BjaqNFZpJ0rhbBtmXv/GvilTAIcY1nQHhm3l7iqkh//
GWj3ZsBOotTDg4PCWUDF7N7g2JmAr5rLvMuPIRTIDK0NEz2UfARnIQjnqSL380ZiY3z4aY/AaKII
Ghlvrp+kOjQZW+muBeQYsJZmq7F+wKubCzw6UFpGjgnJ302RBUK+U9ySzX49rwuxnRtncrtx3dCV
C/ofi9dRzUekZSqEGBzXi6xitS/gmg5CeMSfl05Iu8sExgIDnbvsta2dWBFNai/tHW/bHxN3+hgt
OliJrsduA9oMqzzCN9wmgAEbYH7pBDhIieo0hg+vVxinWgPwEfrN3xuOBa8r+pPqxNOvdSwhS0Ii
aB4fNwMN6jxh1MMyuHYpdSmyqhZgPa+JZh5wxi0vovrM6EbAOq2JJDkzuMJfgQpJwEnOtA45pqiP
HKjDpfLcdexppowwgQIgumXaa9H3GdhW2Y6JDxPBDBAlF+WkArrgNog4nooSCv5ak80660nLRFXB
rtLr4B+sh71/4L00wmP4oeXp0zTiC3vpBSMCYJFjnYxyF9ooWt2Di8Lq5uTjshKuX6dxTm/V3b6p
OZ4e2RfnVcEnXU8Enky8urSyb0PteEl+oGtqadz7k5k3553Qgy6EG43VfG/T2QPdSUn+vx5iY7QM
O5+vO9NBKBuKSjpO4zTTtvBQ3QleR9DRA8fA9crSai0JXW1sDCsAHF+bqGJ22a+LTCg3hWKmvNbd
UfDLEKJ0FKgZ8JQiMVLZA5ioiE1nMSfpD6tm70lghe84xPmdCKtOruVvirUB69E/z8HyxpM97V+z
lDYvQBLv8mVrQJtv8CwaMu5jMlodPAm+k9KhCsdYZ2vmKKKfXAXlC2BKEP6EHOFpPasG5GfP56TH
J70XLelgapoOOk53z0rS2eLmP2zv5e0Wb5UXW5VHWByZ264IjWUQ2LZ/SW/RBvkWx7NxB7P0mnMJ
NEzkh++1GlUgE1rwfcrT8RNNGavdz/JCBPfI6AoRKjirjadmNh3nO8IZHhpIWwIM2Dlr6uMtb4hG
BzWs4yA1bWSWZjg12djhVR0JhgYeexfrLWdV3uJtJts/bXrPdXQqjZt9f0FAB0FIMY8hrwfwFKs1
sV7EFaBkFFrlPrwaO21/4DYaia8Y8u+5uWHduN0BuVMhO668fVTiPqtor17JFFOCWKBqBRKEUyAk
10JJP+zbmjQ11PTg6ZNpxtOO9m+WmqitB5gaQisbn/td9ZSy82c/m3ZFrEghLbFIm6FYe1eWnj+t
psbxD0Gtitj+5vLZoZmX9Dq4VmGz5PyPwXmLhfdNthmL9tLtGS9ePUb3Kgv1yl8GcUmyHtS51vrr
u9PJHbqZ26HpAe5aELtCQhae4FthA4gn/mWvekcXUY5WKI2wEvMh2VwOCSTyR7IgvDNB7qJD+0xF
Cp++RtdbgfqDI3T+ZN2+jEEJ+jsiIbfGHFPdSSegOctfSBSmmjtiFUUicqEyTWhMS5hvURQWfdsj
lTyldWZ0RuGQAY9r1vzB2lG+JzdExFtPvcH25KR/ngl8ji+epatbWe8UofWEmhgSTzdhpcEh1mlZ
Szh2MZsrY0UrhuMCSFWgRETdKF9UdGWU5WHcGjhx23nz4RPMJRMwfTn8vOXisxK4VlLjbmBCzL5X
GbMjnmuMgx29cMsvm43+YtH8VoxwGuZM5n+5g0gRekC4/jX3MUK6u4uald8rTdJoWmISvpXkLUIz
wpZgDOqy0Y8zSmY0joUtCA625KXQnRzPq8cG11b5nUIFkAVgI7E5BkpGHxtxbzOISrh/1Fv1SDNL
Y2SfAXic9DNR8Nop+hs0tBOosbrQOy6Bc6pmgXjFeevd7GfNuQrnKcVx4FSolJyY2tJqLpg8rPLM
mNQ8fNzH2HNzstyeVG6w60R1KrnPpBp2ZstiEN7SUeMnytptJ5TCCoTVU9l9b3pmX64kCvRnQkVc
svyS0yjyTjX1/gGBLXL1IZsASdIAq4yi/znsiYCC4cvN+RtAarSicthaK3MkX/+KMpLoacgLimUQ
Jl6PFUiJm0wIp5TomLN2hY7gjjx5Gbpc9czhJFKMwcuBPIa1F8j/6ErkS4ap4HLafXvY/83mWZ3X
/tBwswGElwOa423a0nnCIJML6/Dj6KLE9x9LOiYeaG9nVmgrDmht8X+N78HxPc8XGUrXQ9pM5MiS
/x0KZNoUTAOUGMkfkOmKOQpveO37GIZ1FyRYd1DrfhYMxJI1qQmJ7j8Kwpv4k/EpOtgqSBE+iIxi
K5PBfg6osDBV44sWi2UzIKng3OS8HmUKA9d7u00sYf2UN3iXJ/xxRVHbUQ7TKsspTnEXedPjGNBr
ON5NpnnL0UOj7ErJj/LnRlBizQyApDoZQqR4k3lg3qHCJPKoiq5tfvAhDroopjIjEuKp6+5BOlgV
zrSzGWk6/v8fhtrl6SCzjOHVvYa2pyvN3HeJZKB6CjyZuq7rdbnVIJ2GFEv42Mq2RhvTwMtuQPqE
jV9Ac6rVyUpHVvA32F9u4fppLDqnYalAQBCqP2uvTi9s0eAgGB+jCT9xOxR9VXMyJBVWVrplSQv9
WPjOOxvNjUEQBuIX/UZ3NDCCYZO2cXDfqdFHqJgBLJHea4h/1EgjuvRd0kjgyScFn26P29g1ztSL
2uM7Ohzrv/M2s6i0BY8NlzEp+CV3+O/XqM9UlToksDThGamILjdIjwA1UzhGIiKlVnssTbhQ0sdo
C3iJA2W9RMxFM6FKBLG3TcZbfaS6OfeE0o8rwaXcNruo2WxNoeC+Tj/1XRwPhgsfsrkjOeC8/ncX
oeUgLYFzOOuqIuzikXgOQcVtpnQwQq+qyVahOpY/3SURsBfV7RFRe72HHs1HCgQYC/fPQ7LZwWSp
shy3LQ0FMnIfD8COEUshI7F+gjsJTDlMD/NiLC7I1xMoIU9Y4yyPrKBHrenOMI4djN2ymZTfpJJr
DPpKMAUMTCORD4w4IpmSFKzKZigY+siTA7ejEuhADmLyqfOJZdYCTRljIYqlGX/oBzZusfQekcq0
pP2UQU0LU49Yn70ylHtWtyfweNVScuIduYb617y7BoBklL/zKjmb+pDWfWHcvUXhmCVDba6xuoz6
00866wlsvmdEDYAj091FlPmjA7DWn0WRsbRC/hbd5S6pxPWGUAPNhOaBH6z+xFeKPnGWu7OB2LOe
trD783oZ8bFLas93nJ59sfkjl3m+VziTCZNxmF0kTBVflJxfQVfKl8+xBqK8ilMH4wwyexGbKdEv
kb+Yn9Vsg+C6Bwc8bx1aCdMjvJMsCsiCNYYAA8fjNHmBLnMnvbTESQlMJkLPCmWIfa4DiB0Ifv9w
1i1uQ2zTHG9Jm/EVE4Y8dCP2Vs8gQiyEzD+WI4m63veuTu3V2bh0Vl4gBC5WW8Gi2wDTYRVP2slt
xYNVkrMaZi480GpCoVdPtPQurJFTxa7Wgriv2t5RUSeK23uutvF1VY3yRNl3UYK+6VXFLVzz0uwk
wWzx+wUV8QGcHE5/PA3CbYlYi1R1tzYv9aaFr6l2LlEqJbc8diFgWNiMhivKtVyfZZ0c2b4Ay2P4
HFAPiwnyzRX9JqSGXCI+193SZXFQl9XGoL1vpyZSlM+OOK0FOYbr4WEgW3h4Wx351hldGrEL86Xu
GpXRs97Qn0EkdRVguqx1LXncjXSeYKSFTW4vbnmEGzXKq5JmZdpPCRPGlBthQlPPzPIfG2bmO6JE
qSkKEBO4lpg0d5eb7Y+spg5AbXcGwtacd4ak0qcFJXWpKpBKs7JzITuBa0NGa2heuD66J808goQ5
mAE159gOigGYxyHViVznwXhgPCZyElOZ9XpQ+1+2J8OzlKcysk3VhmosiVMVtjK8L82P17naHrT4
KMNwz5/sA2C4iXAqyKQ1dR6ULesJzhSdvECEMxCJZCRmlsgLT6kSSOIq+vDAOpdgJGaUO8xhqZzZ
fQLja2wkvgRef04CrqHACGNhTmebYcqDPTckgNxmgyLxXhJx/BBxVtYPH71WYcKzlTuZKUedaJg7
JnDv0yxLZ82Lns/ZNbeD+n1IFeSwL2SYi7YSwPcV2ymKwFlAVEaV7L3+x9dXVKY8HLCQY+8yPm1U
4r2kRY8rxmuk3xzOZV9gBbnSct82J00JwTCQIOFKSnKbR563lOQwE17m3ZK7SkaiIkeENeEFCiCQ
rEPxb/Gb2aA4aMMW+KqE+KWZ+oDB/mbD9k0VniNrq/cijzivYuAaDbssYBvvfN06dTlSVVlHBbFk
4Zo7W7xFCAe448FBqcM8VAxl1shlC1IuFoHHixOWPByfyH6ptpk59b6eIKqip2ZZtNv+P3gFWgKl
Zi4r5ckdkJ7eRK0v/u4Yah+rBQwPmUYv5K3mVHz28UaxMgob4YB3F7CStDqNPUd3UO07kO9NUDKc
MsKW/IzCuScg5WRrAeY10rivIgZFS3TBdfqlWkfHDlYo3QY3tz1lyrcounQtvrw9qUhCl8Y6TMwo
ahI/KBe9bBbwRh5CqSsO9qm7NpsYO8b1mhHE6/NBpGAN7iZfWTiWjQgXt7C4fI9Bi6T5DyOYBkHN
0s623NOKOy/JyocrPaN+iiEgYOdYfmClX/FwbGLkK576VEpvtuID3j1fLEDbshL8L28lyrJHKkel
3GFqOvdk78uXrBhZlMzKY5rLzOznRpM6MPG9D3UQphsHwAEYpCMSW4B36EBq7sYDRAp7H6yhoq/m
UYJOo676kpJaQ0TcYb6W3nPXZyHGhUQZgzDGMHcVg2nWEVfP60+j8A1HHTMMqNskTM6ZLRiq936M
HfKx7CxsRY3nYjILoyeEmJfVqNdK+KKq3OinDbTEglLY8IGVgLleF/Ed4EefLK+CrkMtVmxDo1jM
SrMTKlJLCoyLzbV5Q/kLGUiTtzpydMwXe4f63pYWsxrt9fbtOFdU0oyQ5hznSGgTyRCsLomK4bgE
U2l36i164AfWTZzlHwV1FFNlzO5ATrDf4CvNuNxVrdXVE8ZNNTJ1xpJ1QF/6uJ7O6vaos739RabP
6rr9bzqb+IuJWAApXYXnwiLAxjsDSL8XB+j2qqrHMgr2tSqeYl0YJpTREk/0K1VZbg33xcDWv5qC
BZFRzLfHmk4LvjAw2Lz2+C43qGllvDbwrzGlZisaoITSK4iDFSr9aI9CM2aCzp77kniv6QPjoYKn
bT5KostnEmHyPvhCBRU1hap2kIim+aRGLEy2QFDVKhi0YYO1TaH+t1P/Don0uDGHFzsx02YuDj2J
Hm8WeTs9Py5MKf9G+m4WGqq24B1w/X8RdhQcqgPKk518rlIpip4IXwLIwgjA36HmmNJc1iHAr/sA
r21Hh4hVfhXC5EY05t/TzkGVI/LSBRKJK0OR0eBtC/KXkahs4z6VrqjFFCiXVCYibbnZ8NlQq0HK
UegP/zQArOqnbx4ZMYtcBK3Tw7QqZqdHcOTUxUd0Rc1NEor2B/lX1J4/721EY2P40sTgpnzgeqGw
9zU62xvG4TBOQtR1sMZ7TOb5db5jZI7jwyONnkI6gKL/pLN61A8VLqps2FrJBl/8We+2LQseHxPu
3oGD+Fm65CAW3mgwv4SqQ3UHaVJt6/tqMuCtTzEztcpIke9ng9FlI+qGES8bIFe8psQbdRKjNeBj
wOVS3iVaANA86NXY6/h0JEJcBJbXXTmYKbvNRhTpLwsqg/Abm0olkErWU+8nwHE6eOA9rH+jBfWq
U6+qSI96TkO69bWFQf84x3DRAiJJmwNC5m7ujxeZfz58BHygBP02Td8d6ImtE6CWuds5dUi7CvjV
iALIqCBypkh16C71FeFaMPB3QKOs0ONWVrqCvgW8c6RYzhKFapHoX9dYIW82zmAoLBzT56m4tnUx
1bk56zWnkW4JO2Pp27257FprOf0wRaVl1sze0/z2fCEtRzIe9Z2VZIboyPSBIXjY2J/OgoG7mZr9
EJxZYPxfAdfKbFQ72M9scn+dkHJ+85HMaKJgc34dJIgipplD9BqmOdTdHjc0Z1tZWjnwTaX6dk9B
kmvEXJNgzVTKCWHDR6rlZ3mtJbsFyaO5kIKvx/p/S++wwRiK4Bpg8wGeVwnqNs6fPar21q/RTUXJ
jtr4rkO+lDv6QNWbT9c6/0AmRqXMV8HVrNlCD9DKPMwnGNsmQ/8HpXTpKjqcf+qM8hviamkavSth
tauxA2Q8o8KrHcqljRegWwVB7LV6f8KToQTujIaZMLxd7SkefsBObA40+x1NY1Ozt1/18qZjkNuh
xvfoV9/P1cS31BLrjY6xgUQYU9yCfO/DDV+6jjceLLfg/J4V0MRFQMtUFxZOGZUizpzMzW/R1PBp
CwpeeJSkem8/CXCgQCdP9LZw6TNODquTEBZrLaVrksV4J82J6+jl75U2PHK5lJw4tOd9KQR+b/t+
kMFWW9d5GNf/wX6JbVZeRevUQKWdkDUXnVckvamM0G1hPs+2Nbuv+zVVtHUiEMSlj61n83+b7KYj
Qjuyuhum87mA626qZug5F+Q4OftISwVMy65hne73VVtfF5yyW3vBRH5lN9O58Yj/6x/pQCz1t9lK
ZTCl8Dy/qEWT9yNad9zwBFLr+wVFjEbsQYUWjo7k/GfqiVG9Yg4VsKiNH99fYtBISy1KGsLN+dVQ
0enHM6lifo4RL/atTYmb0RcH0F+nMgse2geCbyGxzzigYNNxKy2qgJchOpopO0zgr5L2mtHaKhFZ
ClKzB6jFFUF7WlD1n3kEjLUbLXDEPclQgivll3dS30nIdJBWL+sYtELNjZwoQ+Xdb4ovr61iXd5N
9u3EnnHLYHT6u8d5OL/bPZF7gknP6TMu5oojIVi64kFYhCmsBJlC+kgOJdP/hmpU4SXIU19qJYfO
4L1TO6y8qju/5Kjz0vWgYjDHsj5RReSD+YxwV1vGCnviWhiuXleffAZ5WeemwYp18CF3zkvg+5Yo
XiLqolHMWkoa/tvhJUZqEJMfWLheEcE3jhRiQQBZyqt6+9cFkQM/+EOWVuLfu3XXhjnouYTD1OEY
cOc7u446FRTyynwkcN/SFRh2jhaO1tiSbNIcVdrKaoY2SgO5e/XF0xdnJojUQHYM81cYtU+mhTB0
E+xlQcoiE2wjzEhG7dajrzCGFT/3IXU8ZdVFMr3rISdLwhItbPJgNMh0wZqjTcgCYNO/Af5FOReS
8pLpUMoc/7O4Ov6dZ2CdcXfg13/37m4Si6j5Wgk3ZOrVgvXI66MKCe9x0g0trRGkK2ELZ8Ci0+Nf
CtI0+wfamRtduQVRW3fN8IbiumXnhhXo0YkXLx0tKmaSS2YDujcCnyNbMFibpRDvO1nrxo/DnSZI
6n93A3zOH5ntgCIuD1UZ8P7r5XG2EzcTg/SahAcS0IZ79ToqDeVcUhpUuMfDU32CQkpbTlNM0gG7
XLAl69zQHYWzx+m95On9lfJZ/fRHXFGZjXIzqwsEUFOfb1AJVAFcEZIOIQ5N8Vn6exteCkEuohvb
hxHM51XIGBAYOM/ScZ8j6Jce2NuafwYmUICoba2OLGJtU4Aa8xuIZZV38L357ezrBvavwUf4DTWg
fKSyFsq0/gC3Kvn8OS3xuXxbmgjyKGuV0LZd8GY7xeaZGwnRLm83/Rya5PkWfdg9s5PJJ1+GYcxO
UQXTAN1CoSn+PUDeCIkcmURCk1Lw0o/0MBVNvtZcwvRJ66DD5lvEQQL1EzhEimdX/kN1z/K3zcvm
TwCjwE2Y7hGxEXbKktl5XqUsBJigCVgYrkBDcFGEjjBxkpaLcQKX2ANImupwg1Hq0fqTfi6XkTaE
YntmXaVejyk5TYL8HfRD7zmjUmfpbX1dJP5xOOJcjZhX+tWWC+sE0LGg//kY5YSgvBJ+bOGrVhrq
mmHdBX+tR0ohNLtenjiZuRS9lqga2UjJBDE5bp2mZAE0PRo2scAOH2f0Qkm6iUjuFuf5A9e3jF9k
1ZFVj1HBoql3F1MSw9jKbHL4OmN6K8nNTd8Xxgsoat7E0VXIuhWy6O2KpkVULUQujfa89e5XfwXh
ItxBxLKTVn0+TL+VwZXwFfOYjYbwur2zNwcQMsyzaJSFyJzBN2+GrEpgonbCB+jawJUxVcUkTXWV
AO4Qik3DSqu8IfebVaH33vBGLJiKCrg9GKc0pfy1tgu7Gn1YGu9e3EXeXLI2cQHcyTI6skp0Euy1
zp71JbshrFwM7bOKKoqcH2CgjhsEjaY6YOpTN1hclfo5Y75josrtJMHPbIr0A36nNH7Vv74Kx/55
4TqzPf38+eVzn9QQ+lyHtTxzrBvhFboeok3lgjfjkcTqUCXxxOoZhHbPkkP/CvY3iyJ2RANsbIqz
mwZgL0vHpc4ypucInRpXRYyEMvcBc6qu85nj51ky6DF1HqTFZMiRpWypG3r0bo6b6qX5I+6G26RP
drRGu7tX8n80DT0ejF0p5e3+jTYrTkBJ693bOnUSGHrqt+gGTo4pmt9GqvcAWsPyqRiIDxsnGVv/
EzN60MuPC1esnyCp7aFUQqnM2nBKbC5F7TIxfjFvbBa9x+YREqEM038EipbGYSKh4655JjTKFIE0
2AXNEtpHw+xlE7mKte5jwNnQ65W/CnnoFpQlLez5hYsY2DxdOFa1eHaP86npPkBktQK1Nl0hEjO/
z6EHrRWoT6iHPyuOaNSnbB2H7FecquGhseCCfQ71B3yGz2Uwy52IZa1t1N3vsXoYTWBiFhnosi0n
TMmK2UhG0oIC2jKp2YAr/MRCVsXFJLyDIvO3DMT9fht8uGUsnSy8Ff1KdTPl9YsGAOqjHEkst+kQ
7A3r22FXWlePARGGNTp+5eqcmGFXBOMzO8GMzEKHyxsrxEh7T/hRLQqU7NiVssudM2Ne8RNXJx/4
nul6TNB2FGXXR8eyV/LfoV6/Zh/AG+ssoNGxxVMMTZ9jRbIMrlZ34WmOCJyvyF9chj0oRmORNez+
o8VHc05xz8WlWGlYm1FuAOfXaORR+YiKxOA3JkPhEn7BXaSOif3aOb0ZLmoFvS5Zc2w4zZxjSmi/
s1gkAhZYxKh/gHCWe2QiaXFEg/o7xvuB1Y8oAv/P99hD7GLTaY39gwKSXeyQbnx/vsic1ErLsHkg
Ik07ZMWrd3yyhZiNCw2Dpzscg+vkpmJB4gG9a/k8xr0wpXWho7Z+EO+ljtHzh7sltRbLeSYTscsi
Zgg5jm9wGmKVGURzyZPuM2FHCaDPw8vK+qWV1GIjANXySqEAeybXRxPvPxsy31huO6Qa6wWt+qMH
SvMeChB8g+LMN9y7iOFXNY39PqKO8w2iljB6e6MAIFq/8OKPakgDv7htLy0NZ7BHHkn8VEOK2G37
t2MOe8VfDPced0u2CIko3C9wlzDBBFyAKb7QXH9rx3cir3aZczJCkwbs4F6O5W041av3TGLv5Luz
I6rB5AoXP2A+XF75VHKn+Be+MyTR5P5F0rRrI9jlr9z/C/wMA9vubAvjYpJsh6O4V7l/Hd5+ihLm
IRxEpEPRLrP967AxXCbgVdgtOm4vR60Cz84LMY2X9apEX796ZXUJgQVfQ/0V9Q5WP/8Ntn5ckcnF
7xOvKQfMGBJOhhPZBbioRlPPRCn/5ueAUmWCHrwrYlBuZIQwpaQhjGXJ+IK51RteiUIoTrQy2u57
4IjxHKPvG91AqZtBOpvuvuMJwMsnlpaU1+pdMsy+0HbdpNwUoicO7/9Ic5SHeQD9enRlTsvxmvZT
wy2M+uBHgV6r42qGeSfm00NgoZwd1rbbTTwPxYX7xW1+a7uPyVHzzOEO+MRNNj349eC5liVGrQsp
hK7CORVXEeUCqZHPG/h17Rz6VkpkQVaf26PWLiLk1SEzSALiKM0ysoxNX9s0akYrcZZroVcQlQVk
zzf9SK/Zy14eeq8mj6HjNywD+GE4eLNu1qD1YSogGK+9pykEEQVmWpIa99HVNdTojjvejUnBJGJ0
6C1IXJ35PM+q2COlcZxNia+TuAlkY+gixymx1FMFfL4bp1p8Y/r/IiJfMuGlwacmleWCYzdB85PS
rXHqHvXvEbW4iRQ6QEmYXPNJmA8+64AGK0uzy+eNCs7YhkqE2Q10ta11kU49ayJFBKiHmNRVrnOI
allDjKgdRvOKjGc68i7YMueA5rtaRm3GzdCdFmgwfDDII9ERIVMw9D6BaMgIpTk1SdewFlRvVbde
RRqBLvXmoJjophy6M5xaxzG1KaQSisQOrbtjqQiK6cMojYgoAbMYm4hFZ/kx9WxM77XWI4FEUhfr
Q9WWfSAEckX6i8yQry5MAto48I+rORUv+nHUJr8KuyI87ABjJD7tY4HcXOE2oWn4oidfDfklMCZU
N0f/w5KsTjmPxEzjASzM//UkYKIMd8JY+VUDDB4vKRgQpghwqRwd3QA859+OZ4f6Ix25Pec43lze
eg6J1fjaUCtDZ7JaI/qbbALbRUsQ3Uti8QUFWKanj5PaAIdoMlA95v4QJjF22xPTIQkFCeOb1awV
hoychnR2xWSN8GB9Rk4RDMrLlzvxoQU7speMMO0IDMwjSYNcJi8WLjjqzlzt0N3I85KqAc4aPyb7
CG2OfUkAKTG3BjeKt7lKFa1tIofYsRAzPTV0jWg7ErNoaisk47/rnxB6z3VH8hphnjGyjPpsxTjy
fRmMjy3DKS1c3pgbiln9hOnFsLJh/r4Qqdew1MqiS1MvoODFc/HtkD9zd5yhe1xR0OU3vSFwuYs/
nfHOZ5fCKO/CI51F7TtcfuIw5Y6y52LY1ujShWQ3SwJ32N8Wtcj3QI+MkoUDbDzsdw3kyJQMu67h
PunfaWQgfkULr100bvdL4tcxyDAB3T72bi7TkQ7xjGRBpV8kymurK/OtNtt73GaL97PMXqEAzNWa
r30IKFuj85bWk6yaLsMu92VKuoAUeQnn5/ytJePvQQ9jxeRng5Rh7/C7TsCYUKCu+1uIwRhRtE6/
kdJ2tag5xoaUgdIFULr//LMKE2hUPQCZA4O+g1JYLFlFpdROxnRrOTYShhZdVKyS0wNt6JDcNztT
/JRYYmad8wYG5k96EHLzAkRmLbBQlbudNjDLlgdV5iYLuGebnAWtG3Yi6vTqizWjYYOZRuNmQRLS
jm3qkbN1VYCX/RRbxaaPJBMWiavRtk+v4eZHpZoTXr0tGuAlwpWbxM1zQosExXC1mMynvZJl8gCs
VDpte9BNNNHAbsxFWcoLCvY8doesRi46QlrSN6/7v/cLcJPIarCnVjlV/D/hEWgkANYW2n83ao/T
ivSuQ9gve4DtKL8m0gwY9FDDUt4iXWpIgZo45HjjjXOpelNzocZUVzBm+Zb322wg7bRnjGDp49lr
R2HPDQBLjQjF5V64Fc/Wz7fckNZUZ2qauBeC6KJdHlSeibQtaB9PF1a1ElrIRTpqQQC282NwfpLc
lXtZHQ9ZWkFC7KM5GQv7AHT2g+Lur4+7OXnANMHIE8HHw5DoPaBrux0OcrJoglebQUdTdrU6uAcw
mffMVPSe5Nh0aClieiBilbPcAo0yIIDaEatQabhHxzYsWt0lxiq8kcQmVvw9NcH6vW5Zm68HeiPk
S4uwB0eK5VHMOsGQsg85UYZYjcFCJB4CC3wKILyf0tNBW7MPAxprFMHi8/JdxDi3Ri5WqnqpRss0
LSpvfe+YmYnsZmLevmhF9OmNc/KWM0S9sE2wIVehrqqFUPTo4uetxgWB/R4LpxgjRW1TPXynxg6f
gAHpLq3GNfmgMJucztVDZxYmMm01IhsdAMvu+YVlUew7Xc8d7H5SDOHzDhIPqiPOAIAAIWnnNdoN
5bUQTt/6emwi/91ZTZc6vvfdJ1i60Re2xSRicDUgeeCCW7Ir8R+YcfjYkQ0+tSZc9BPyl+yUyokS
Ql4XmsWMTsZZ1FPD9PEGvTxd1tkPlLacXfJeaqt23dZpTHzjYP0LzcaD7SXEF1BmOgJhNL7l7MOV
ycywZiUSu7CRSE0l/NMVWezMfQaL0xAOprA3O1cy6w7WmWHPle3RxdMTh3YeakB1HwW3nVJyGmHt
wTka8deohLq3lQLtPya/YKXkuDolNMgRsCIkfIUuX2kx4OC0jXmb8nD7bcaZu3Zfsc9MzkGJHsXr
G2r02hiBYdZvKT7rpPa/hY8Bl9aV0AiUV+IAJIGXo6DT+pdGxC2xqZ4kcVrRfv2K1FgQ+C2ksBRS
K0yjU8gJwKWONIvippMAkKkrWBntxO2PG6QnfvjDIN9E8KK+oV6nftYeGev/O3ZLxwtfkmpqJgEJ
5Ex8kINQY3t965zb7PmUoH6BfjVF+Ov3fEQeNJf/j8xi6xLCy7qh7NwXNgiTmbnbDxIILbUjJymE
L2uqCv3Y5GcvNBIzD+IvAXCKGL0ZrfNiHPDCwrQ/jZGwcuMISJ6NQKGwrALjNx/tmvh92FQ1l8C+
DNaRbRipe2HgF1ggW84sgO17cNt8qw687Z/WNw7c6QnBGncjVeUB57dL/mEBIgTEmSdmydnbqOTG
PXhjskOcyryQGF9vMkxjXRX4x2SSdmy06eweo7zlJDDE8/0wY7cOXtrUVun7RDG3+bZj2zanag6F
sYf4o4KUYq8jGXv+5G6ASR5u5izaACdqXe1l5FRqs+oHsgkoP33Ex2+AMOk8rJoHBzMN9dHhCZg/
Z+zqOAqsZTvu9qwRizBGtSaIb3lQQpmJn1C4bJu9eV2102x4wqRqFhlo3E/5+WmPH091LD9aelJ8
FgT3ZpGFH//3yNDPL/eLWOtVvfIfk47vWEuJcbvNvgeladJemd8atc8Ut1utkGr8fimkw0WeDf+V
0yBxaiCMbJx0odGKhwDOLHlcGxP49ayBnvtQ/QPYbzyNqelkQZLCj4S1hSj9qJVvz4yfQnL7+GWs
8Hz4+AuuBQfsV97/8j2otGooxMZD15fJ3loBNadGmbF+06f1C8m9DCLM3uf8MeWwYJsg3+qd4GxH
mrGlZ+jGdgwBEJ/vh6ZShVm6wLuBD/eGDy/XMxdLE1n385wP1tA1KOg4VnJ6IpcyAZlqA7UEn7pn
rf4VZaSVIgh4oNHBaY1kph2iv956enpreCy3gJGeUFbhxp3DqqDqSBRmfCiPPg9ILhVQwAfGEjwS
6JuwO1aiLz3dROxAEY2jdwYJu1qt0Fh/2FM6+jEbLnHPptuJ7AJoFi+WbYk4emK7hJoCBwPMhiq2
Ybrp/65lR3cv8hXlA9kiLuc/Dn6Dv9pQWicBuWeJqGPZQTA9636m+ZSq3whdTO659jDb97+LMYLf
RVSeeCdfs6PG0pN5SBfqp3NK2mLbUaA+pOTwt3plwNgPCyHOcUq/H8RtP5SDRqmfsdFfEYMnZ50W
LknZ3WetARRMjoCZHbgBY6Pg2t6o8p+DmQjpieiyD5Q/wTlmTC7/EvdL77MWrxYKKTQykM38noCj
1IPQy1U6/fwrVAPn5dwnbsc2CQW7mSvGk4qQ1gO1kmqhKFkaxFqMaGBZ7CvFKH3qdMRWU9HvAYNU
tQUwq6MNV5AqdPAtYvcPiuxSU/E+EYyUPO74regLFKFJ2UBZ8I8sNENk6EXkrr7jxt7vHUiVJ9Rc
n/9GH+dcofkq4xdShHwD51uWMwSe5oba5hdA4CGiDghhjb/DukvSNAy/7FKCY7ulHd7SGskTc/4l
l9jHSjofEhy/QcIDpI0dzK3VyfgBUkJthobwUQu/+su9FuwcWi3PDxPkAuz6lQ0j1/IxeiM/rAdT
JxZlvcHDh8pJKgbpWGQaKnPcgn6dGcRCEJodZsSisjHhyHhcK7Hrt67bKcqLsER6ULdnyeNKKK9+
65L/t4HBk4tb0x5YdKQWvgDn5qzQkTpKCxaCY00ZWFEn4bH3CHed12u0ZCk991TBYTX51DRXgNLl
z28fFJdZaX4fMGbgYI0U4x7GjmaVs2YRdPkBRAfzlVUVPSUPDn/vCclAEZymROYp9frhxVxR42FN
fIgWdVWJ2HY9YwbWMGW4hTqFzthG/OxdCjJmOr3nHENp3ZY6ohuhEAjuaozAhn4ClieBxKdBtsVX
Ic8NAUAy19Il4Gl/rwm5+4+7Zg51Wzy70Pr0vYTkHdRHeVfV1MGbKaBur3sE4RLo7L8NivRymnDI
JHGWjYeD3yjG8/X1vKIWSPYb3RIY/YJ7G4hdZj9OYBPNZ/LGtbkWyvLDSs6ZM+1uSuE6Zla1Ewwp
AyAN5DkeQ/3x0gBm1Im6pvWuABdiG2k/llEBcFkjWHbRPm0+usJ+xQQyNHGeBE9V1xUy04KL61S0
dE2b7/SKbuV9p72ayxBwoh3uN4ymqWiRzp4cJrKdOTGUjJBUJSbeTjyteGOJB5AD6UXMY0rn87sJ
+JzxwEgvCcIqwidhpV2dxwDLLItwneaupaOnaI47zCpejOST4vMte7LfdaLELN8+qtuO+ipJohOI
1nU97ossIWuk2kmF0conFdCFpZOVd6r+/i5mxM0te5Mi8CmOyhYQdNjEjkozzYSEvFGg4sb9Ik2b
NvVL21trZ9lkmLQIdXrcHMQXm9sCzPO5PDdMh8XzPbnWcVN0g3QSodRd6VIFqRuadsW8r6RtBI99
5Qj2U1S/qAxHwHv3SQ0rVFKzGWAhqtPY6Bf1CWfRC9kqrSyfUgmtAVWpUfKpy9BSRQ4Bs2aHbQPb
NsI/zLIqc8IhbrETSKj3s+koUDQ87NdrFlR378Ct5RqudaSzHxx0hLrtyXWIbIqxxS/6ScMW1jxa
7aaTZSEQZjInxcYaJ1YRpbDcg44F+hd0pz7oY3zrcup07ofqEfxtfZUPvOiB8rtsW6+sFUzu/8jW
9B47sMuX0RrWg1p4mbXNCGIYsAXXIyPZfpY3l2pOMuxE6eQhg2xoeKZbs2RcJ/vDS6+chdLWw2TF
eZhQM+gNt8yMSLz0WxXWMIAME/QE2HlPS1/hShyOOfoxT184kkWn69BNVRxK9JMt53UEL/BERv5t
by9TJpPnqpCoevkdzGqQZgmXsIwMvNsrgPLGwM54A8qNRTVLaVv4TIQpvwmZ7a9YhDe6Sy13kQVD
qA7MQmFQkB18s+lqtE4a+dAt4L0JsEAKu/T5KLKWfSk8rA9heGrGl9VT6+pVz0rF0k0u+0BuLDSw
tEtfOnCfUabLD7emVbupwkNVo5hyG9GTaLoN3ns7dQRITIimd/8aRZYAkHSRpFqsf//c44MYF/I2
9cD2QBQkIk9U+VktbDZ0KwnHQOmfbx4wtzb4Bu4Y9wm7iFq4Vx1McDNJx+sTpShqcFx4wcwGl+Ki
KpWqErwclDlnwu96FbQJ2k4WX/OoWwxtAmoncUX185nqabU8DHUf1ePhmFhBeAS18Borpj3hAEzj
GqlbFJQc8jNc7rPFa1VGoGkuoO+HDDvDqq7bEFSeQGOjzW0cCwcRcrTZfAvRJayqtvfkVRuTGSK4
/DnIllnxh91CuiqpEkOlv0dKLkiJBT02zPDIDR9pRmeMIZrgx5aaHoO7sbc3EsN51c2n8pgcYlFM
U4ADfz4DbuL04dT60B4WKZCJbdarndpqmAuR7md+k2pHnsxq17km5mrnDflNFtF/nddk/IrUojBr
xZO5+v17zgC0Xw+AqxAYapieogWngcvBYfEk2z3PyqxbrTRZC28Hj6AaTalKAnijnuSidZQt5/kz
qRuc+7HUicmVAAfbQAIM4bJm1b2tpJFQjQ/kDR6EHS9t7PtwaCgKclFGvn20mLyNB2ZurZwHD4F/
nsU69VvoXLuQiWdlsRq5ZtgRXkYs71kXHXCOZ40FqRosZUwFDT0fVLv2cynlhFNnyutq2XeiaGsI
neJ0Nm/sJGCYNblRGPPaHMdfTXbbfzPOGP6pfmDHyMvvMBBSOLYmS5Tl3ghXlzrpQ6NiZHtW+M5r
xf0gf2F6FOGJh+t8eOHvRTKKcIARBf+X3qjhgcm/4iO8q8fTYOZa3WBPc1naNh6+nX7vNSsO9F7y
mWDCtFuU8NB/GK6KLKxMwZHezSus58PmCD3r14FeI1jl+U5oq3v5Bktbeh4GVGO5liGclnENA+bj
MzHBFcir5TJJPDtiJTO2zxDvks7Qu5+vS2z42d1UqvmROFdQ27YqrP+YTBCwPqR+QakCgRiI7shn
9A2YL2v9727NeT6wocIN9EbHO3/qsSvlnhEFdrjDDPyH8a47TFSArmfsGddwB/GOoupwTEIrH7Be
fo/paCfuYJz4USOtYZ06ZyiIxzF6bFD7FE5wddc2m6yU9ulRKTQKn6tCoTRjqH6WO1M5WTc9CJ7X
foJWIbePbx0zfaZke5QsOEpBHK5oo2TKRleB+iTht1KhxMUaSAVUTA4aHLa/7KmQcVDKCVPVpYtP
SzVqJr8nzF8erUkUxli7Cd5GC34+nDKMebpNtgMrFAexIcftNsLrH5ZPU9HCYvmbFAqlpkVWxcAx
Fj/56gbQbt1FuQ8ZK6VhcouqutYTUiwa116RXz27H8G+guplLPPMTfXh1EV3eywzjWZ7IAqZRBf+
585W7WzPkbFFHweD43IxX6MtND5FKrMut1/rRvARrIELKfu/YERuSAr7xyK9anQZ4tFvRiPllMpR
lkW1jhro/RLef0SbN6p05jHBKazFzvUIO2YCUkgB+nlrxO8NtckQI+7744xwx/uWnlV2Ru+4bBmU
fanI+7AdiP9FgRYV5MvQqx/aytghrwinuzYFyeLxa768Fvawj1fNmgzT53pa1eCI/2qCuOUzZwkJ
OuX+2AWz9KlsQGQwvFqyUgs9RiIfcRTH8KncYiCAZ3XUHG2hI45+PWs1ReQg04ZvmVeoFuP02dZ+
5W4OWSqtYrlkp4NvPZdPgzguuDn3Mo877DIPvonKtB+5WJzuPgVAYGWHrbWqRcTiJNQKSUrGvlEp
V56Zzy0VNrmwnbOLSVS5l3tXIqu6c5bJs9254yrNZ/g//rcdSEx9GoUfkncJB/Mip8MVu/f+A8nS
OivSroQiXOaowfTV5NzKeoCLPtYoXtdCzQedWJ0j9hau4ZxevP2JFskNDMkQIuFdrqrmcgSkbOGA
skoUYXIl9JP3ZktBsh6ELWjurtx5DUt12OMZIFdLj2nmadCFoKA0dZ9ABqxjXvuBxm0x3JMA35eI
q606C9wkfu8djtwCe98L5PWtYfCrgxLehTZbADruE+WEt86jIJStVyoavTR+cdbFD4TvXu4Bzd7o
PXe/Rqo1N39CG/Ix/tGYXDmuBqlTughFVMZdDP+pQAbEpfjIQG/9N3FgPShJZQ7fNaQFqSKhcxMT
2aVcvKlEi75t0gof/Q6U1K8ZoZHuJZ0wmdcshNmD5vFg+ay1sKjTLpj9lRhA3+scM7jT1PYVgsHb
9wyCPUy9l8p1uvrt4rQXM9+otrRZ/dFrbsqjEyENskAkG3vW7NqXmN2Hyfn5fw5p3emxduYqcjVM
POFE2VWbNUrOb4x3ho50jys2sQBm+5/g+hdQxbILsAdFYmTanO9TbkAVL58OzDqHH8x/G1kNyLs9
lNZy/Hw+koXzPVk6GtKlZytEl2JKGp/hLAFnB/Uzoap1omVFFB0vO6ljANEGtYvZw4CjS5CtXhkg
L+DyEgdpx3k7w8UlM/2aj2Bp2ebGgyDNKRfXnMxtuC0bw1KcSBb35H3lLNBZCHMwrghj2qOOLPN1
F7pedenvUUdh9qtIChSj3NTPMMQP+0uGzRAit9nk+CBA5Wwbf0CxQxkHhSsVKoJkeBzzBHoxR0wW
kc5D2O9LPQg4ZkBM/pvtBXhnnSwtQ0J+utb42q7Pmxk7+uEOib8RlWoiR/RyTuY5vX0OjoBx44OO
WekD3lGLkkkT82Hrd6aVyAt63FrVnR78Sgo8VNZD0G9YIaqR7VxSECyozonSTABrkz5ghAhIHPbg
RF7O+YhWGVInXTe1XVfmp+qYlr2XjCwIC6EIr4rE6RdpDtkhTLBz8cfiYsZ0BrSUiKlDu+wjaQZV
duBjLBuDcUTg17nF47sdpgT6PxgwyKAxYRR2Aq0FU7j/tnztEsFTtFvbfNWHrlIFgZmSFUvV9ZZM
/Ly5wcchLb0jfdEQIlbR0K32+J/iaIJe1n8flk7/COVOyKhGkzApx9Q5JtqHJe5FO2jWS/IJqZFO
Khenu1hwwd/7oHX/E4OJ9SkBPLNegaWMUSJSI41SFwvyPOEPfyAuxw/DEqK5iYjfGN8NXJtQTM1B
MHvMEqLTPtROyzup/aVC6NEiOSmCRZ1sABL7jC2jmAeAg5vXiPxiM3dX/vVPerQG26Rx17mopQvC
kBrkMS+XsoGzoaunZudtkF0cXA3o0jg4sdexdAGVqYnagUWy6G9iEAXihFm3sYzqrHyiQerJFyGX
t2W+U1tyk3SQaB1GrnEzxggshuX0BMG4Y63ZL12PTdCnwsN8pLHzVpXgh0YqYsZ3d/9b/gMzYS+I
2sCnae+em5a76p3O2Tpqiy7Q/hD2EpW7JvCipRBD80HbnWjUxETZHBhhaL/BQOAEmpcK9oyby4pU
A04X+aF915T9qX1jeH/1/r2i6HKJ4D8T6t+7ewdVeyNi+64JiIRIyWVk+yMv9u2EUeuT63+mds8v
0Ot1XdzjKJk2dau+Me95P/x+IpT7eVhmZlImseN13VgFtJCdfbyY42iRMd2VTtSthGdO7gF3C51F
HRbs8JBUOtdQeO8IZNC/i04h3rFUfarAkO4HCV+v7sPk0c/McCGUP1T7eS7Rb2B1EehB4x9m4wUr
UC0Fs2N0wYCPhUM7dRSdODDDaQrxdS2GaQVDamf7f9G+sWIrfxufOislZYGgY1KkWUykmfyPOU5F
hqParujkzYSyqHKK039hDeQGt2cGzAhNQ44O0HKKlsiEjnISBAlwdnfZDoRnc1UWZXD/cDMDn0sh
/8TbE1sjB2Gw9FEuUHjl/nyKFLKp/hcu5V3HNLd41bJPLmJVE5NgervrazAaSURnwI5cwIIJ7K+0
kS5qHhLHtR61rqnu96FjEU1cWX7p+xeLdX3vTYoAUx8mAQQxtDoMly3m+zcTKqESxqC2zUPvk8/g
KPBV9UFATSWppzcRykSHdzxG0x+NbQ8bA/5a+OPKEAs8mRpHQHh1J4/0LDh5xz66mlIomfJTiTVO
g/+kplXh3it+4YAtwW1ldzezZX42a05PBF0L3T1YsoIGXeYPO4HVlsbcjktu/yaz/LmrKBtq3tHW
A7jmd4egc3zx9KHwb34nzXBPJ5PvYEC9MRlabiuOzNGGMNjOhswOW8WdbKpQTQa1hVEN3bizVUOD
xVHHu+cManj8byEbSjvh1MlBdL/epxPp5HNe2RhuXbDN3qFJHi5tHibtzBkf6MKKd58lX0p+4ZAm
4snR/0h9ivoXeavJG4CtOk00OHwYFffw7xCaUv5CkUF0EmEKzEa+y4HyKhAmQqF46nOTmsniAqPG
cA2PatsQswopyW54Jh7knlMJHLm+WfVWukudw+Fr/nUCt/uJi+ZagrnzeihH0X4M/Q1FEAyqx4kO
PxwszCaoohEoqpJW6tyRP5lRU2he+F7awxai7uGeIHCb6OU0xbMxQ5AifItublJ/dQ/QkjKq/fLK
lj5WMOGcrk1YD1SGIhB7WVigpzLhnQ9D/dk2gdl42pZg200Ch2k4X8SYvlY9y8+K3SIO8RXKukJw
LrNBsOePiYR69gybKUafo1AsH0jbZ4x0PSQ1b38E45Z9qVanX9wq5fjestAfWnmptKGK41jQ9juE
+rSc+CVct3IpJyGflhgPID7R54a42Jeweee4pqFMYPMwc8a26BvqLEV6LIA5ujSk91cuNVZBKjnc
65hYi7681hmgf3VCZ++OkYYYPwZbCM8KmeutyEzJUxHAl+5Y3uiTJvh5rWiI7YehRIvFElAriziY
f5uw8ATio1uMLssRxRrKi69/1PAYRMlhUjjo8kzzTR7vE4L7DdGG9ZiTHD0KLlZjsA1wK/XKz2uu
8aCRVy1No4vkj5TiLtRcf1tVUi0NsSgay0nm/oqCSD8hQbMooEae7aDJRZrfuIdGT7eJcv7BYF2r
HjFz1pYA4KVGU+Adbh6cYRpI/A2cLK469atojLKYMN3N+T78q/Lpw2Y2X8psPjTqzDWeNCpafyja
Wzagd4CIECfpd//m+pMEp9SUf/wCgcEKUg5Li4W5QQxePbDCVtQD/pLCR5jKuiRWrQoNntekp40y
Ep6BCfg7qrje4UN2fJ0yfM5uazqTucpi93BsJBFC4uTJacjDbRaxERPNShOqPu5qE0R2+GiK4kYv
d8x2Nd2G+dd1LaaU1+GsaGXZeZWWt6Z33D0N0AVhfTURojSGRm8iKs/9u3DgaPdSyedE1PxrN+7O
42mcBdk03StPblFr6gi3gVVvwnUGJ0ZR2wIJPYMkK3D/12UVsruBCFHRTd0ObRJQzpzql5LE1KVx
bIPD3c698dmjd4rP9LuCcI0g8tnFNx6B7kwBewQ4+XakxoufqzfYr0Yz0pVVOK0cOntmxrY0tDMH
nk9J47le9e9sOHXkI3mTbiQl9aIwmMWrHTj6VUecLaAe5xzAZD0bjXomkXj8Cjr5ApMOjwE4b4tw
G4v7vrG1VUKLRl9xzrNwp9X+EYMsm3fDBYfxe5vbP4mh3gLpkPTdjlNXaAez3L9z2HQKV1T8WLzV
LfSj1fXz1DqYjoWPizqP+eEtbpC9uDRU9E1VXBO+5bXUQG+DaLDdfArQxnYCRXAc416jzSKhMy7x
AtCruo8Eyw8hCwgKkSwyqfqNlamiOaCJPONZLPneBPXesJmXbWmGY4Bx5JFIdE5oK0ppn6UU6tTp
uCGqtYrjoXgNg2AL53glsk8Iyg1eAJPrWfmYFHi9mxx/xiuYyOcVQwsNQkSa1rRYG44Z8LfxxQvU
r/zkYvhfWGBmskgYzXhnua84ZjSKQF5mOm6qQMz8vItRPb0k88uhn9EiI/SDaSEGBlDmRx5eh462
6gTU/w9XHJ52PpyB77HBKwJyf62cAGAdyLTKy3kpk/GzsJA01cqLx0E/gn6C4NDYEAmEoXzw6CGL
ot84+xPU5lvj4QeXxYNtNhUY2Q9g15StGD0x6fWEXK5WU2jRgVBAsWUpQObz5qGwnn7Puw5oQjcV
54GgBi+jzpe/zSEq6ZZR+ehOSvGHsXIHEBZ/STAgvxMaBlj+BC+O9ipJg/Rda268qN4eExUlJy3f
jHKf3a38O5VcQx5NBNi1L6MWfm6kt1FbYFXmDKP1TZ+dob0RtkhlQ1XCqXMmso1bTKOLoQwvth0K
YinAdKYH0e2wVIcCaC8nAWF5aBIk7f4pWHGlqKohKg5eDhd5uLc1aJ+r/CEipNCzYNqUXM3xVduS
AuH0gB51SLZPOcv1yn3NfYqYP7bCU4Kk+Tr4i7NewPKR7YFkW1wNygrFpPRMv0bZptSFnKLYtgp7
0Xa3cOItlFlGBUYssRBrhXxCGay3Iq9SyA/Y9a7a7zensadYcHN3VqlT3Sx6A+q92Q5/JQNyqBkY
geR2Tzjg37J15+rLaZfCz/lyaknJsYRnusLJ6lRcSwXdmossGPSmdk6a3cO6X+elBDRIHhsjIKRs
VPqjbzmvkPH5LrFBOuSYdX31BqH2aZjniFcvl/B1DjXfCwnVSC/p4JK+D+YntemXVA8fRtDGtTqV
VYyg+xOw8LHnFtN4sYjeI3jcNw7VoNUHe/j7Ke2SBE8ZgWLO65w4v/hqkcbinJOGtkCIibpGzwFV
M87KrQBkYzoEwlxS0tefV8u9E+rOwqsr7MXSxZ+nNzUJkHDLfVAS0GWYXsoxVB4THAu716vcnZPz
lWu5nbF2UKQEbHUjzaGWoqZrzDQ5jIKaLr7AwLoDCuNDnqsD1jT32BPmlcCIGwNnHLHGMGaAGkWm
SLMpv2yyVTO88TeHm0Vjnm++t4ybNFgn/C9+qsSzrDtFn4LW7CkAzve8O9Fluc+dZ6BOoZIiQXaZ
YF48v6I251LUPVRadJqUyo3Do6eSotF9ULXFyrb9RoKYEV780oR4iWCQi8a2cUf4k/oqfgiJxcxA
thoujKFXRqGh17TTq0CmjPsMdUthLWkSKkszqfVx2RnbIY8D+aBpJ/EQ0h1UOMlQI3ety9Qz+7HL
u3RLw/rLHWnv8BnxT4BrQL+8ik9zNc1W2rKf5kefiSgR7cAUMnGd768G5Pq5uW9ffLGoRh6oL4L+
s3VusOxmJg7D9nX/YuWBn6DoYOWRW1It9y56fGa7LsEFcLr5NTgNdT8TdSdhE80n91mEFMbBTryx
MXAaFx3UG54O7+aYA0a42QBAu2OEsc/x7Z+1m1i6kgHMt68DbpuHE4FBoAkcG2+MHMGNzN/98fjS
iWRllfS5dtKpcPP4a4lNInNDba08Xm6zBXabEEaZDCwn9ji1FRAv+VlSDfcpl7CaFC+qdrAdzTu5
4AW82lNdQ65UmKyb8zDs73GAn8bsLi2getJMoAyAt70EEdGbHYlDezUICbeI6ja7KhOzRt4ChQQ0
s6yC1MJ6/M0umtb2DQi4b4Cd5SZA3M6ml/awShr8Z/FGGU+xfQ2jkyNZcBl+Su2CssU9wouNsmeT
a/7mKJEq/XXTXyjdLzICtOMZejmGHVNQBukBdsHRiCHfSjx7BafoObitNmiC0uqiIga4GlRv5Dex
vt46DIyM9/hV99O614U5I+IrAAM4N4tTUUoSz9FyL2+hi9CQNS1ecMPLd0ep0cGgpy65FqL90vsN
lzi1QhN2/S+QAtlJcWrVNbpt+CK32NA16mymgbwFmJ90WFwMw5J5SgA+9iBCKpT1LsnRlsstrvuY
vxi6I7pgWyUdcvtPpyfQXv50C+1mg5gbycv4QVKjk8uArNLbp0jNW+HFTG1XRMbgmtM8cy+DJQyK
VLtwoaRF+7QKhAZvfoQWXWTxWj8KB3zIZ9KZDb9szdFSTl8969WIZ3y6myhUf6g7uiNqJSZpTUlS
N5rQohXApVhgc9dNkB9+f8CITZq97LgRCA1bnw9fFhgEsxRpEHKsWPdH5GfRepacGXApHuF9Vo6D
I3xy4L5YfnGOn97qaJVYrZd35Pwi9jP4F/P05tI4TWQ1A6R+iEEDOI3ISOF/EnAmZbi/pMGonKTs
dM/DGKgi+oqhYydpt+MNbAMd1MiJztA5KsJSyYgGdv5XQabOntzYXjs3iEuZtRf+08F0ve/4gLRm
VCnk4VR4+judxlL/oHZpyMJN72t7cmdtgh+uEeFFyaqaZrOlm5ez7Dx2ar70vcPV+wvoriq7Q8cv
Mkw1BTA8OTbdjZjVl3Rg66BGsDlfRczjUR2iLR5jRuG3+GKZ/wvJSizNcVDRpHO3N6zw5KNcnwm6
gK4/lFhnOfcSWBeVKSnKWdClTHeFYkBorGQmTl/VufXLad2wXoXOSZ87vFQrr7eXVEry84Vn86n+
NXgGM/qaGFk3rBvCaW7FmMRguS6uI6C21XOQP2s1VCaux4tGjxUu9rA6YUjlLWRS9+o+tfvN52xi
mD8zLcoXNxbNu715yfcRwHT/VfSHsm2s/CXA7OkSOBb0+NBF1WyP9l1pjv2KvGhYQo69TIoaxO6G
BQwhpIewA2AhgBmu0IQSOV1607c2ddOnOo3kD2C9AuAeXYp3tQop9QxUr6t5Mw4S3qgD4W78EopW
702t5kId/jXUniAZGzskYm166m6TV1d+dzuqT6JQZ8OmM8gY+WkXrHUZJ+7lpWVjqdBvDiov9aD3
/2hwa3SBL2uEVjehNOuGwv4gJ5wsi7R9+tfvOLhezDzZptMqNWVZpY73WeyI5gqEU/cQnPufuWd5
PjhBDQaLK7jS0gssPsXxrdFmgGMDEXu8NRgELJqqR65uqbPRJLfJAflHBLQiA5eHKNH+6KS0+drc
dj0WmvVwESXMRA1OpN8D5Wnn8lNWYzO960Z6DDwzMVjqDrRlWAcRfF+dj8yuS6wSgecYiOFgjJLM
8x4cz7hfiV+BCPnNa/uqUgJaxbPMh56ULggbhvODd0efYXPSjuvY+IcjCjEh1K6X6PYRpcJjh+Y/
Kl3mg3u5psaNbmhsbr8vSpYjV9IDCOPHRlu9fEm2a94VOlVAH8V74KAuRRVjFS7nbfiyrvZzcjvE
xCP+M3PiZ2TTJeQ350axdQ6QEOHn8x66kZqzBjhI8SaBwFVdIsLetpRTUihsBVgKNS30NVdfLTdN
wxyP8aTGcNC1HVXWXIJGMMFMNVN8IA2EsucwbUZT8RSKYVxWWkrula1ZKEbkP8S/SiGFuj7qJYNw
QAdoxZ5+CEFmuTPPGEZUwY20jNBX/dn4xbPdRDRVWDQXltOtO1si4vqNhIwRtbFFRr57HVIAAfS2
xDN/b5kSnsDczzxBckc6P1/5GXGZLFDwl7M8h+iL1jI2mjANmV43EgYSn4eABrUtA6/axKu1lVcz
yzUsT7MNmXKn1qSbZvOihwFQb2g/ekkt1Gte2U9pDYyuYJOwt6Nav7c14x0YuR/PJeyW9AGTDqoV
gou3ydY0oPu0tVz7zR3sHRVuC9+tkLw3ENcnn8SOcBX41AbyWIEVDVYRBMSoYnee/1iNk6yoRZZb
mJ6KFshoQeAKrwb2E2lB9MMNqLNx179+lNK2lAeBzUGoDEKO2XeavKVY49CTMjdEBBf1T9iipGKa
RYav7mPVL0SSkQgL0NvmiTb+TFegf6UdG7BPgkhlDnD/5l8LTxpXQXzEeBsnWJt4DIjJa4Eqk2sk
Un7eb9DEDHHmipUVW8bwCrkZuTD/7gb/USelaewJ+tNkywpAOhoyPdY10nYww4ue/mTT/CFUlp5/
Ab9LdSaTiXuJYGDfomZtIvEW2KylYKlJh5kfWybk7nCrTRHXjc+IrRKsfPtkJvQxaBOa1oAMUXT7
7VRi3mCLdqb/o0w+HZO9CUsZDy91Q5/ewtmzk2gDcnfR1JH2y8Tp3FFRMPEu6uI7bSrDmC5bS2IU
BOlZWrmq/IJ7wUCug1dWxprIqz1eyTIVgp6U4J++L3pmfjvfqaNDZI6uknMN5ClHmXkP0ThhDEq7
2IV8S6688zIg9HOz14v2hOum5BQ9prY3fx4O/sKAB6ZN4zisvWpPPTxiwo3rZT9b0fRXPFwDPcvY
Hen5Lk514ZjVYF41i50qWc0VjfRF1SOJXwaiVyWrXrDyeCJDRgs86Bp822lAu6IfiT8yv7zMM4O5
AzQ4SXrnc5IPNU24K8QpnX2eQWjVvtQqQb62bKsGfWKTaEwPoVUdvj6h13FQZoXJB4jhZCT6FoBv
u+XdPpcCfY0NLbBvKaBGw3spj7d42u6ASQOSaOe2kQxM8kSh5MyW73YPeouEjx31yfIqj4VtjCr/
4N4JmbXvlmdq+G0BIxW+0gxWLLDDvbTzRZDzfdJHiPqdtSf92GTOPDjqGIECqSoGfOdlZpxFTN2r
GtHptZqSp3rCD8gf9OUGXNudqPsN1wHga6mtAWpQosUcmzBrf0K2cX+rCasCXfZqJrEeFF/XAPmQ
Ftw0UAnicvwZuxQmZHlMFhsxIAIhD5bJNHD8eCOFKIABSFiQbESXwqTca0LhDadJs2Z22p5fWBBD
cBMY0JqJHDuRMVVZrAM8rmLEYv8zSPUH7ERsy3TgoM3D+7KkLHpxIACSh06EFl+5R69EJlig/l6q
SMaElCRaiKrzRYF/b8o5LH7QzovYIrtjYlUxLFV9Z7J/IqxIbJ+V+S9bpA412wzzJ/z+PyV947Zr
6ZE3HPA84Jd/WpI4sZxvCv1mHOHm7Cg/aFqYewyOelBGbhmWOgJCDfXKP0PoKsO/xJEfHAnj7lnG
Xgxc52eHMgcZkIWgOK3WNoNIEzpWupNOP8Crg8pYv1W27jbngHkNY9hJMWBu2p9uOzxVzQgGq1iW
5+nuUbv0t3fJfXktXQfnxxZso7KqO6IHtV4q4lj3yp+tjW2bbzLEEQdbiaYXpZOVL/YDP1HyCdfu
KDkP8ogKwLxJAhxZDAVDZeHr/NEMM+6nM3P9lMRwadnRDqBcIhFD7odYi+O5cEuvaJ0PR+xUQqvg
1BUpK/+rM5Ct6dVbuOk7URI4sn2gxB2J5v4QvRVBtDxx59bfTlnaFfiqBySvWjza5SMHLmMjMvcJ
9i4YYFcFRLgX8lZ287swWeAvthWCQ0gL++Qs88wYa+fT7/NhLrvaX6+1guek7/jF243OJoRpukkw
pjZrfbNvpkMnDHg8n3/Qmf3VfFYGeDnWMYrFIQhkS4CCnxFQXofdww4joGn/NbEhs/mV2BTs9vTw
tcQqy4c+T/RGY+ByDVFY1yreJV71PUVTCmXSu/OQ4NLX1a3lpWwKkrWPCrWI/j5kEmHX7Bqjvk0x
ha0Svthi0vcPU+0/irzD7pZvYKF1ISjsXvgl0xU8x/VYfYxra7BHLjsMViTG38aIWYyebRD9pJq4
QV3oqd8QsbGg8+tjRZZhG4+RdvuY2SrRxSgVosdBUkUSkdQ50lmo7UEpbggb1KBl5kdhBbJDgw3a
I5aInysGuZIR004QpeShdHfw4wB+RPxOgRG2E+iDXn0q0PVwPMF9tJrFVdxqAWT8MuQZ63+96b8b
W/6OQLiAUiEFpOiVWGrOj8UetpLtk4cF21i8QHwRB14jLwu3lNbFDQfqGY676F9/JqSDwGve8H5O
3/4RTG9VmWLm7lwMkSsqRi1eyHmAMC7BeqUxiXtUx+N4MUR5qBeSCmK6D04McH0lwYS5oV/uFG1+
Zy0n6ciEgAyrHgWWhsI1DgvrnhZR2A/jhlkwkDFjGMpitd/UwUbvzelab2Cb2SmVqmgwHO3k7QoV
mFQzONVCf2d7hCa1adK7F+0KKFst/0UmTGzZL+wQfE9Bbj4jrIy49U6ibZCrY2bT+edkU434lqI8
HioCDiRyFeXzv7SIB7wkgxs1Gh+tFfuhRPqbjE82LYPldE33hxUbVSJCIoGjfYxVYZrtDugQKSFy
CiMHXCPFqD36+RwD0Oc7L9KjaHYTYeUrb28GrOmbt4L4sUl6A5U742kowOxTUwmP7+s0u8PE2qxT
TpRU9DpsNyH/7lLKWCXyv15Qe10uSYAbIQUIKcS8VY8T8xv+gONewnmx0vv6K3LsUncacoLTsslr
8Qw7JIFISMz6zpEW6q7QSEyffMH/uR4lX4eRfIcQtaOcyYaHuvSdVDMjQT/Xx1ahY+C+cYVPbcm4
OlqEKqXkRVMWlptTNVakKqYPo5WiGLyRPRAzir/Ez/k44NYHFaiMWcEVi4djU4Q7S9KeVWLNdFmk
Lz5I9GbNDPnbO4GmBxCR1YxmkuMwZ49HBXfliXe08gcmX1Kp8yXml41Pfncrr1Wjv+5cUARwW72f
dcZ4SE4h9lQgzdeeWTSUzoCvXix7FWiJUUQeKoVgc9bJliPrvsmPeGxio1PgvVkjmdA+elNfo4N8
/NxMFwAVBpQnJEBcJ62ZDC05Q1ct2akOcFASZstzbBd9ZQqR6rgNGCKGEP0gQmuG+ByFA713lCp3
t9IDgSs94ebM1V06l5yzBxcN8XZzWSc9eqDSpOycidM5lf4RF35YnrDeGwDP+H/vqxBpbmXAiykl
//+i96ulwt+jVwSk+zaSVVBWT6jxoN4ngDNe5sar/crUdOZntr8skT9+I06WOBHhFg4KeX7oaRnA
+k9TQ1CeKKKQ8M8EGCUzsBaS25UqsMBUBGYI6z4MI7KJGIRmgH3gVpXaLv5Ph/QM1c9ir0x2lE/L
sqIwPyB8WS9J56LdzdxnYn0PwQSBP/MUsWW782k54ntdJv4qyGqiwAMx0RhmsE2huYrflVCkIcvB
4uMr74hFM0aZrEij5k6Oq273WLoCLyyzXDhgb7IXWKnA/iGEVY6GJAawX6Y9E+Q192fKVaKIsadn
kfPxKww5961tY+UdJJU08+Q1MyabpV6hZsTccK5efPBqYPbF/pZWkYo6OdNvUH3Nt6J+lSuis+7j
I5TibikagQjaLUTvHWaGRHL/o9DD2A6E9eLsBj4SVjmKceA7GcB7NOWWutTLGOxPgotQcu/H95Hw
38IskD+5mW4GMZ4eXmSzaCGuXSL6F4wNgzFhRR/pgNBaDHdTWipqQz/SKXQi1msvMQ1bfjkXNvRJ
UczbeHWmfo8/gR1f8BycGICei9IbkBpLeUkaeRBc9j7yi/+QXmfrEBsxM5g+Sz1cnMfLwc6ou9jY
g726glh7SSkZWK8UEPIpxLLIZYHiGObS+qzFXw7t+xaM3vvz993rkUASc75gZvaQLzoWy/1MZsTp
xQtgXPHJnJJdxOwbpgvCpcrL+pdBlVvlqD+JbVkb8TwVJQrjI2a+2ahhaV+8KaJi9t+ErM/tMuNz
xpOhjZfxBOP2cpwJN//M+g20aNN38fxTJJcID0t7uZqhijWDa3xmcnP7IFCa0MOpsTkuLu9vNqnP
CnphIEDpENXM6XC6DTcToKybC8l1NO02ydHkCe4ng/clE/Pfo9FF9bXEDDgamlz6DKLvNVPmnqiO
XtWML4bn8lx+CRMhnyP6zVTV9eflSEzJXocbyd+PLD5/vXCGrr5KeYXQOZCE/s1zFDcXErR+rDG+
iVn0cncq5hZa5g4/BxQ/rtSH3CoU8/2r76CJ2PTOmZYHP+3PQ/OCf4VbRTUOzwJD0dUEp0hxXHc3
gZcBmkxHR7JiefGiPnt2NENLhqSP9B13WKJPQPfLmtnKtBW0hhAbL0TsR2DRqnqMoEvDYT70L60F
AdoO55s0XbJkq4WWuJoBJmHr2X+XiZ9ma00ci/htjmJJig7x+H/PKJYhz1rrpSlpbnH+DmVA+NDQ
PLLCpv0AX2FgfiMPDW6EHb2z7Urvt19GRC6BCXDaLiT/Uet+XyFU/RFYENLHJOmt/dTLqqHqwIP6
6ZEMxpZZA7loJQUioHufftPKHwNfIBAJHdNDJgXJ8T6msCNE8f18ykR66r2/JQQjorfMdlp8F6c+
twuZpOpE4TkY52I/2C7IRCid2fQE2GwhkKip08TcUmn7FdUDm3Tik2RJngu+hlMBuETw0bALpeuO
A2NNM86gQRAzDZbBCAnhdsN1pbwF8WZIh4EUCyd+FNAAhCK54IioW092HDDP7ZhgxvlMLToYU+rU
YwDzGz9UBrfnd4S/B24Vl6PlF5ICnSejRNX2wmGAlLBbAhrspvzReBax02KqkXLjwrzjB/ykqdyh
dAprC1DO+LO6+q/R8qVZPPmq4ZZ/Woy1Jd7TQQtv5eTumCInH1j8jzX/rlvifP0LfBPSSe5trJc8
gkDwG0lAIOqXaokQg7OOxYB4QmRpiymjkB4g4TpbqFu28IEak3uUQPawLc2uF1ZyZSK0dMkyMCUJ
gIquj19fk+ynUSwDvBGuvoGxLOmGuC1y/3x55IbvW4Oh599feXhrissQytWn+8HZgIpDgqMRu4Qp
PQ4lxMuCGE2fRBo9od+z7snTVC9aE7PfJ1ertSU2IxJdd6G3Ux8r5Zzj8osjxQKKr6MJTgCNhwG+
65PYacAVGwcB/yrAyl9KqzmPbu94hZzJJz16y52zA2OjNO8+cswRyZ3rBCfYbLzI8WlANTKJpWuv
ZeU8ZiQgPCQPQ1jf//M0D5YOcu3meJ29gELROp55GMUQ9GNv5ADC/mCAJ8qBhLJWSKOad02E444i
Z49UVXdSGkgg+Slnvh0f572P2Lo8L0CTADuKRTdnu2yXiAN7gExXuulmLMZcNiGiaGTnSpKiyiie
OMhnIFr5AtZpnqrYSpRKo40ZbsrXsyT/EF4f6xkgxyGyzO2wmtm/0Qp90m3y93/8lNMoB3tOZpwJ
a1E4l6BEceZj7AcQrTD/s+8UO0Pwu54dvSWtUULJ52h/TCulAKwBgYAh3Pt5LqgOkpVirkjOzPyy
aRNqvXJonUdn08rIdlWcBS29MN+Udhq9Q2GontX4j6dzG+gP0Cg4psKL4PaMEnwHT9EKGmqBuZ34
L2YC2jBtXoTxJsRMsgvWHdPxXokM0tuMul+mql9PYVys4GU9m2BobQ4ygaobOKtuNnhbfBxfsQcl
VjYNbbIci2fpBUq0lhWrAsYOOmUM+YO6yWPfF/3xXotcLmkNWcDUsnHhr0ZfRnQEfXfQUMIhdSu0
IfWOK6h7cIUYU5OskcqiOYqDCyUVATvF/LcRSEfZnPAWXrE2l6eAhk3oAT9OiCT1uR53dzZ8sZNC
qBuRVCo2xc1glLIsse6kG8QshlA2AUgPzf0lcmvJAc2TsxaChN1uUYpe/Mxf8rm4fvI/yDXJHhjc
jVPAt8QqzGh/oBpDMONrPinAXQJa2xR6I/9Y6JBXZbaR3PtItAj0SCbAf5P6fow0SA+vap2ynzDJ
ZVNr2mAL5mf/dumvDmDn7Fm2CqmXY+6ZN68qRvt8dYiV6T3aGo2XeS+A6aYHGONKJI4c9pQOgwh/
mJcz7sI476cwQ9yxNgwEfmlkB1HwTQQ0MdkEpRV3orKwH2KU0//xuvCG6+xRQVA58A5X0zdiMLHI
Zbpp9OOK1PSekTbWjuhyexrcZeek+7p6RhfhIIlQwg8nTuBt2fDVbn7uCsu+wvmkcKNDbfOMiUig
Kv0c5/tOcyEgMPQZSd8Mqd4uuRNaCWG+iiUHHNzouEMCFyr5Hl5ex5D0xHEpV9bAz0ZA9+s50riJ
R03vonXgR0q0yqVg7e99zM8xp5cYkJGfjnSCeSB1CN3UieVGI+karPjkzL7tyz07JSsj1fKBcMXd
dwvY8rpPr+8Lq7LhhA6l7hvBTfQofjiizZuSsX6831HVcF0jhqqPfL6xOxXKvVX9tYuV+v9YxE6I
C+OYP26+dXLVdeyDrslJFdlme6sIH0BrgxB2BPdf5HsYX9v/vSVzD/FltejObUS5MBAfrPoPr0TH
vLdtFSpwjfYA529cXHNGYJBH1hzkuLNvTtxcm41rnsiTMoa5ckIaBcSvlyP3y0y38Y+KUmsiacPt
at4Y1ko87Gx7BKYH7fGSHyic18xnGIS5TvoCZUaZp0psCJhgyWLuJqXUQEZzxNrF7k4eKaO36GLp
RQN6KDl/9Qlt4CYkFut6EoUo0aabVXtA0ZqBEQhhLo4ABR1v3HxRpr2WYG5u2xhYiwGnhzDCdMGB
8qKaLFQHBNmMASye9lyHoLs3kYm6Q22zyGbNZ8U408TGz/o0M2M4ZQO5JhaombWx5hvs5U2WR4SV
En4W6voujA/2WnTRalfIo1fLQZ17T4SSAaIMR4W19/KMLV2/msC8cOrBZHA6D1wqdzY9EFa8ndkc
jpl0clA/GBilIa1YM3BdR8e0uiajLRIoBqQpQz7eOjv3TI6t5wiFBx/puCmtKQTDfyJcWSmprIju
L81//FvaXw/6LVmCUg9eZ25R7gyHgri4E4VxaK0/GwVF1rl12XUia4MQjGQkyE0j8DuqA1EOiWj3
xTGyG26RlLavCDDePkWpjMqxzl1+dyv1VvILt1JPUAo1km7FYJxeB0/hsD7uY80Udk2hdFE7zfog
qww+UpK1LXy+elQ3QKJa01zK5tSIPqNoZYjEVHjR3/Wbhc91GuWmxfiDcYUCVR2r6uEL9Rd/gq/X
mo77N/KP9dymDOwy7N8LUEBigzXCSMYedmqJ3MmFksdyUJ0nY0zLrKp3eno8Znvic/Ej86CuzGYf
wo5mgkxELQ6SNBI8Sz3ErEY8969e8sG3F/+rOXlLfCNf7P5t2QXvIFVEufioyrqeEWC63y//0dBe
09y0HXorArQpweakzhHnyxPzEn5kWaSTYzQDGL7HFvuDgRzBEakTg4+TV8UFh/24nY3CTGX9KpEw
qPZ1BjeDa3xtYznlLyCiK6dkWcjjwH02jibokjkb+136CpAsTSEhHTWNlIEfnfDlBiAkb1xo8Zbi
Mw119X+px4qk9yM+m0l8RRnCwmlmPxnxltY3boq3p8wZUYmrS+M/r7+6pFNf1Ya60IueAEb7MPqH
+M8zHhAIqx3os1L5wIe1L+BVOm48vlGvVtWKxz5UW54eYDSqz5Usi4aiqXNOFUJm5b5ACk9gaG8w
LQ5dsO0rX6qktG7RLFAz4/qP98k9kxh6OWXFX6errSiUDJfcIHcSoTLhGZ/nC7+jRF3EBHBBvr6E
hUDWzfg+TQFbXNi8TS9Q+ojWpK2UmTl8lTIl1TtguKp8Pnh+R0Zjo3YzxL5HddYUY7ddfN4wqjnA
hniqDNshHshdqfu9hrVNg49Whl+k7I7w6K9y7Y+VxU2mny7ANbmxhs6VKLuXB7j4BpTdwySbbI7W
jyn77epIWzhemMj7hQLzkPdMBD2BuPW7a9pC5NEO7QYfGXRO4khcENfLipteKYP0KXCFXyCTlAw8
P+LS26DoHrUJc7Jfd4cYWyhrIBM7bbPoaYuZE8x5fJCbapkrY+kuB1orEkYSR9nmdoXX43ppA4fu
V0XMiF4cdMGwPAS5jFr5HTmK01kg/Mu0BDMCbCQKcUbYjrrcNdA/5DS9qHcR8cCbXkLx5nz2oxLs
rkJOcSDB3Xb6q5snoIAtTRkC8yOw4O9v3QxVRilXE3qs6smvhhV4kRoStLC7r14rwkxyJeFHplBN
nCp0F58hVuQgGPihrl8M0w6oKE8cdz9YqF4ZXUgfYh5K7l8/lXj43LEMPz+3HF8ZOCFgo45ssl1P
kmFzDdd/1wor2h+re/KK6rA1YTuoMQQ8L5O7LmWjGovyfwpQUbg4yUvxi/SYJmrYaIiXZ4B8oX/6
G22liXFN02l1DULMPf4tYZyqdiFgy54AIU9y9XTPA0XDdKVrZiUNIeszmO+7TOEI7XInRE9wDvT3
cJhDkFa5wf/rrE7EqTuCu20rFVWVj+oE1svxf0SWpYoga1Sm5VsTS2OWkMa8IGH21ZPPiWd1hyHE
+MwOUdKTOaUEpIEKyMJbXbujP5Hbas5byY/a4k+2DuOof7mBpkCDqTm9B2IzaXXyOhByeEu0j1fQ
rRd6tqJptR7r2+8ZzzZkwAnHp3CXyQzjcRYcObZI/A43WI7VBiMobgIAj7oO4gjJZobspJQDl9Ww
bsEV8+rxqrnHFOVK+QDVLjw3Py7vjfJGCqidcTLM/jw41j/ciSiSnypB/zNJbrovoR4/VTX4Y4TB
e6DWp27e9tHGWfDfN5i52qv71+SRTfyCGdqmPl9RXz8CcsEinm9Ex3jmnV62O760UiWfAoPl3+7g
86hkY7xORitAXwQjqRwHg70r1YaNKKnsI+XXJpFFFvYlbASLrqXNevhQG2Q5c0g0TDv7D+JURQ0i
jqj8r5ZZ7BlfpOSurrX4l6g+l22IdWqU4YBB+bMa9bcSmCIVNyR0jg8X5CusNw6/YZMNtuWxDZ0F
+l1hCxE9lhQzfjpix49TMl2+WojYolf/L0wSYNlI4TqOZfWnxPHQrgLuxLDUFMh5+fPxgM804Ynw
HnNUXMFmvo9Lu95dLZmrDgJC06I5hQAA9f1AYY2nyjTwqS32XvdLIfoZd4978NnGNNjs3IE86uRj
DuwFoMP6OiJsOV34Td/5iqcqzYBHzeZhEiU0ISNJi5igEP9MAw0pI4TJNxw5EE6iECLC5/80wjWY
CR7eSnLgeH/Nc0YAoTO4BxdfsoE7Ei+5Eo3v6C9ngVk0CevAW0dI0WtPTTnTRLNrcIBFMzNhAVT1
DkbRLhneXsuJ2S6x/ROCfklqiTISpSV95bINYkhSo4iwN/NWOSJ2ReruDdlJwQvakbQsChnhqzQ/
8KDGF8rfTLn9kpZZNCfD6paT9fMclSYV9yfeg/uOdnDZE1gM3DsSRy4aRG01lhOGXhb6lMIua0Dy
s+v9gGS1mGYrA6UzHD3R8duLOZWvX8AwZg2FmVrxT3M3ry6YX7XFO0Q9C9Q13iusq41vveXBQa/6
GESRQu+jDUh+SJHYwReIQ72Td8IsEB12uFTaBqEgfBLZIkX9PK3WqDZAJwNmEmM0V/FmfZHxCr4J
cGchpx1UPeg9k/1P6aoqnXyCoJdiIAUCvjxfqaDoCCg22ojOvYIl9FLA7LwzOJ+bHOyJ/RGK7Fk6
rIwFXI69QzzuvlTShjNRjCTDfuXiHh3SXukU6PNiMD6gj3yTAZKjo9R4PKQG2fmiIN/ROdJZPbbd
ndCsTEhgNsxGqeUA+51RDHh2WsEkT62pRml4x/TWpIkGYk7d/ruF2yEcj8pr3RL7NByrni/UXQ7C
ChhyBgM9i1WfaLMAJIlkFVgP+zsqfZrrePeEanEM89aSU9X/KpnCnNw6hDarwgaOoVLfErW6hQeL
oQW34ZA96eGxXtDRKtBO1uGeBfszdeOaABvzyE8XI8CoHHctj/qgV7XOhaC1cpTshsNyvBo/STA/
+WzRxP1Anoib2ldvyBfvZShiAs9K6iyyQMqqLyr7qMJKuPqus+cvzIWPb4cDbXA5RM+ea83NPS/M
RpXCgvpf0vkvbfwbZSQE7pKtifM4zekg+Uo8T7oMGyfzXR6fB55zVGUSzf9V0wPHI1JSTOp5fQNX
Jb8NZZqQpiTlNgB8yNlk5KDzoxQxzHSnFuEChh8J4iGk8ziRrnC0wAcc8KmLU17M7mK4atuFOJIE
Cy/x/MWAqabSRTOAM3cNnt1K4PNb7i5T9LN43c7aEQKhAL0z8z5vnbxrD2Wmf3ndfNM8IU2JjdZW
MMsvg3MNDkNQGltoHg/3GsQWhDGzLYOo9f3o1JxR++tvYA/L4j3Hu4vJptKOo1yYkSVUpw3tAN/X
Y7gZODU2QS0a0Elz0DjkLGa9PygL0FkGvw13LiX+LOkDq6j5vtZw8EM9H76VPy4XrMaL09WC/acs
0XH94PeyRG6Uh4+D8crxjqhimDiPtpfHGqWimgFerap979EfLGXKvVyMy3HJ0YYkMBjJegmavKnl
gHUkXHgLeWs3HmU8BDqqxT2n0YtN51Q5tCfPG+B/+Tq5nmPYfSq5wHJJ5vnzAKzdT1e2pCnt5DNI
ct7q9ik5oHcqe4esZwHyRtQmuLRy7FRzojCXxCUdWK63ndMH62CTj7iTXt47iEL7wpF9gyQP0Opz
gFzL6d6yzqdua9XVYyQA7QhTbEKB+ZRPQ6GfeBw+kobeiWfr0Ob1sHB7MqG7Dn1Q8/KiuNuFbjCL
FHbcKlxvAAONWtOPjtN0b0pftTcmqu4dCsPOJhFIhpo9Hy8E6Iy0KRsShdd9j3V22dVOG6TFiSx7
nAOEafjbX2UxUdGetsH1bG7K9lfmMTFOOR5ELmyjzSuWuv/zwC4G4Z1ucbhvLrc6Sh91sH7nMRXF
1vCbkZhkJKkVkwEw9nMqzYmGDzNKW0Ptsfjkbly2uRvu21IZPEPZmK2NJnHlwacdAy6YwjSJ7SNw
lphrewYpUGAJsRKvZzoKWOlner+mLPvEhRhKiyNCE6wnQi/zhuY7rH5qnGMopEcSd6IGPFE07Rtd
8b7P/XWKYST54jyTQazIT3AR0l8lEecKlv/cyDdpLBLFqEzTMqikHWkSiVaIiIjv0+TEq+g8YSC8
ywzPFZNb9QCM8WaXAZ9jNKPiBeTYzxuvY1lp7dCpyPikF8brsBwxfxdLNcTynbrcY3eDsg0tFy4t
hG6/rzJ5f9HPSDaWIGOAuY/55zz63nDLXRSNujo2YNM/H4ERMO/CoxvZ+Dv9GA3mO/qokaFsq2R0
UaqDGdu87zKNA3NEkZDTxvZdRbMAzX8bhE1oSOlO7bxupwYdW3xDmoj0TciKDq6AK3ipVDTxTeEh
SoQAlBqxW6zWlL+r+nPqvED8cotleok9ASQkFTQI/o6MxH8576qjRk/Aa4ECPVSUPRefZeIiTSkW
ouFfglDAL3kQGRcXA8mT7AvQujIKfdPiIIW+K00MQLtAPJFDsFZbWRQh+WUO6X9p7itPRBJ0rzUF
nThziC9kLgAIq7TyqwJZz7k2QcMI4JlwZGEFblyivTh+vJxe7EY+ZWKtL2pzxnLX+VHVirNsx1pf
eH0eqh1WeBHYVFZn1g+LDTK97zNy5QdPacOTbpFKpWPzjgiwH3qAw1aEAGzzfFl7iCnrGq9Qjv+a
PI+XTg5j/VCeRUvgbHy1cfLRAyzodk4NGh1pnI+LixoQisW+NfF9qUBMafzd9TrcG4+ZyFZKI8vR
2M9i2sLm8tpfRdNkbjXKo5T4D+6/aE6dfUqRyw5g54qWv0ePjrO3aTuBkns8J3KxYxpyzBxrB97a
+/AtZ35Q6+7opVJWsmsGkVozKIEehd6jP3eFa2DJzyQFklTjK2jpF7YrG2H4MAWSt+0JKfK6LcLJ
GwhfdEBWJWa5ksZrhlGXRqRLcfqEx+X4RRay3ZGo1DSppzFHKkOrW/OiuDfr6EU9yaf9lcibBwf3
PSSnmoB0IV1rJzoLGJ5NT6BrfqBZwG7TjcAcmv5NZsskE2/Rreye3ZU5CAemK0vae9VxnBqZXtZ7
hlf63ADVvA8eXPxVEfoMEOD5Hnq510ruaB2gMtDif0YtbTWcsV/bk72cNdd+wj4C5HGagMPrQs7W
UFYnEB4iUIDXmV0lMsThvCJ80V9mwUP1mhSgZGuL19xf3QN7WoB9MOxa8lqsFp+ewDVxFJ2MIqxN
y6MNY/InXH1a2BGw5EDAgKpQDGxSoESEEHIiCLgY9RBHnISreK4mgdq3inXVjdAPkrIMrZM6TAIZ
xigwO5Uog6KmKmfsDaOlRNfj2fYsODv/2LP39b2afhShf2PA+S35DQ2FTiIMj19a8vViUhdgv3X0
PZJXWHzMh9i1VjVJVxb7Y/WFCT/EW2jtLZhFdWZPdP7WWDkRtR60nrQMwYF2EUJI1tFTRWNotnjS
dDkBBX62oWlWiMpn8rAI7BuFm2Za3mkWiqTdNbiL+AV6wErbrooAlH2wMOhco5rBGmtvnsNmL+cQ
O1zJO1IG6h3QGmTlzXZqLXnkCXDnkuGQw5a0NGGmNl6bdpSTJIIcu+Hi4HSVIGnqtXIanXec9mmD
CV6nF6b3jrpwA0+sHOKDrb7oqrKk2W6xF1/AkfuC7N+n7nE1OXN15dY+1hX2kBHSBN6pNJXUAwJb
p6ZC8zbt051UIDcmm5n8cW0w2596s6iY2mg+So/e9GS7O2LYvSdzO2fFQYl08bhzJGA3y7VdsMMy
F1W7obhyLosi2CzCCsJIoaVW02Dze8j5vkEiilP6s9TCsUQ3YRY7LGlbRSTx9XhTlFpKCnoIpHEd
6uIWxOYTz9bKOepwvA++oKUrU0FHH1KNL/Dyh56vqFZpCjSqz4QqwcZ3jZ66abA3cAc1xVEmASnS
lCAvFCR8n/U7Nq2j9QIgkAOv8wP3W+pd+cIqeVi0BgNxOLF79jN6Xdcq/RS3iP1p7hInrZ2M7iPK
oetw5COcwMLbElSCu0w9HDejAKlm/UzXgvvi348dXEoIAR5j6NNtALIjF8l6+cyjRYLLfVKgeD/s
/BOTtaRtgBCKFustxBXHxrW40UjQgWXzY/lByvLcoTIhXSh8NXq2ehQKLGDur8vMYJhNgGpNbwMv
G1oeUh8t2I5KnvnvLnUmzLkD3gM4AmEinZFhoNl0aweW+6th9GDqvN0N7QtATuSkgFj9UQZ0JPcJ
aOH5dhrup49nr7Dwg1wrwwjQkXTgpMZfrxg7D1yih9g7eKQy40xIZsHA/OI0V0MIiD+NMi0QQcZE
amGjrbQXoEn2Dh56zA+gu/xkJsdG0ZIhSP6Y7uxB5MEY197VosgcNWbI2yzmerpB66NbikHcaFIX
GyJQWwkVlcc3HwPhxEPPCFEL7WNTTuwJOpwXjucrlKncBiJ/GKWVM7q0aCoU9md5gCeUAEVQaS19
PQ5Bg8HGEljdT+UAPgW0vnry8lbbIM7CoGPZvYlkuA47UFUUHdU3HN9Ned988r6ROYp+RlSy2z1R
jalcHqYd7ca2j9QpellAzkSxEh3+ZQHtz/irHCm7vNcUPPPPk7/DwP9lH7Umjxfru4t0mMAlf5UV
thd+byTxlCEzGvSrfwyegCEwh/MRSNpm7Zk1Cf/19LxBCxYA8A2leN/MRDMFuSwQ7898rWkKCeLB
+lxVmfdKxRrhb+XwGoS/zoEKh9YQGvWKOQn3SKVL7kXJ4Rd7xABbo67TOfifLYk4TXXHWMXZ/20I
E3LobrM4+LAfMOznYnoqUCirf/ZtQmqoZ2iL/G6GwxrcwJdEDydJI8N/Oh4tJ2ys+z5LnvG73o2T
x9RP+D6HG58w5C8wUKavqhcJdktj26p9+BhSPXQp1emq/mx3LUV1cHT61gHrlnWv/k5KtRU2zjZ7
v/9h+YtZgFulfda2AZ6tM+TGjmgwlOsr0GLnx64jHChg2U6gh+VzcSUAG2lGcMN/mEeFf3XTJxmx
JzrKw4ES8eBVm+bN7qzYA5b4Cg0iNIlBARqmtTJEBTcflWPgHEhVwFXM+ZdAmrBg5vdLtcJdWkgm
DkwLvTg0iefI17oP336HphnmzMwRr6EbJDAIbIp7h1f7evtUfNulbnNGxRKzPNgMz5H0oEk/h2iB
2Prce90bdfCUA2409Ldhbpk5/c8EWrkQ77AMSKovXREhxzejzC3jUv/tlogu7RPT4bNu73QPU4Qt
v2Yuv5gtcycQnoFHOmoHuq7tyjVsg7I94K1++RGykbb4YoagzQwp6fhHtoCtc7k8oSc2RMcYp/Pe
sqaXrH0aYQeTlmSWaSfssNMZarm7SqVTDyScqyXIcIjV/7VSZK/qHQFEWVpxSZ1/QIYAwpORp4dx
K751/ilASz9od2flEqPeq05KV6JpbpKbERAO2N6gUeHyuKsHNqlH4EWk1+77isX5VzaspEahMZtM
8iFG/EhPCjRFnw0X9Uuf9UxJuGhfQHQPy8k4o61VDumNbMw46Fgh6QwtGwFKZm7rkd/JNBo3KDZw
jF9yRm+FIxbA4GthIH9NxnBhWMVYIQZdAsogpKx/uhEXJXTH+O3uTTCFcQw+ipC3at+y152FxjQ2
F+oblw0Txi3hwANEMjEzCVH+jKOKCHcn39/PT100GR3h0eUUHYVnTyG+rFM2Mtoo5kbop9x90C3G
EMeNlV6Y6oUkZ0uxox+17EaIK2SzMY/GqNjTu2Bv0qPr6t1Ubjg8GrDErwDGMUImYUE6i5LHapDa
crkNlk4VX/OxAhVJABGYrStNhM7EOSAtwVvQTouZWvGAS/y7mvP2bRpJYkCr7WTNAVVZVwXqKrR/
6pkqScCA1W0anubNFqIszqhrvwWESq4bkFUp+t2FjISI73Ydbnayp5Uo83noXRONQW+Ipfe38p28
+UIgBfWzeEe587YkARxNnff05B/y9yvIUnQCBQfXsWgIyvkkg8VkE43zq8kEkWGAY7gRFvRQcbIx
WsyVgLQ+RBaJ5zMzj9xA4/LkqDVsqkfutBLyBc3xXexF70nuvc+scXuybRsms2t2v9wRUsA06OOb
Cw9VxXishvHa41y0im3h4PTfLetcwfuwZkqUhntDv1p/ergl5usiZyoFr0wo/znz17Cyd+Foiolv
zDJBD5YptnSsKP8kLtdrevCaw9oQBp14yaS54oaNObafvkYU6ehhuKLUMQ5rV2C85KqbOmJpVsBe
V5ijxSPdBJrEKaxYLT5btvUcrVYPC2zF9XyYFA67gR+4TapxDBVlYDLgTpddjhRusuKN2FZJz7jJ
oquJzl5+hv6CH+Xrgco4B4kTDz9euW6MwdQkLQme9/1l+Ddbu2CY/5SzaDKERsKPzkG/x/1IxYDi
PqbCLSHmbWGrg0fApL8sl3zjyGQGOX8SfJBCUf5KAJ6Ql3S3gPP5oObrBiTWiM6m7xVKxaHD23LR
RN7qwrZiKcjKldNm1S21hAkH8ZDBshLXquFx2O4MUdYwNgV/v9wZ4bPgPke2lLf3WxdUsbnjZdW3
QadYFHgLkZ541xjbGjVHY6jIcBaBSiAECXUKpArlE9w2+eIJVHu911MsenkH/wiC2mDisL0dHOSF
9BGG9iCGehqn91SrNMA38N74Ah5scLBS7bZP5W/stKu2GmIZZPKk+O31T6K7tR7AessXqAO5JYFu
JN8Zq55IjAPT/Ljw22eGEfZdZpW7HMBBfwkg4+Ewl8KNfUhJ/R3KcnhLpveiiVGZwd1BiPal8e2U
hOINTdUrIM8yqvVUULxu+ZnRUAA22wZispnMj5NuIuLQdY3gyEieaq8WMUn5JRBxryz78odVRIMj
OQC+AwH4+nICP/oNWAcBMuNh2uJzXQAdraI5rSfkG8b6CgZycPoRAUg870Nl8F8LHMb1mXa9T3Bt
hrE9BYhV+y0QsRsjclQa9na8juy6ICLQkJWe53GoGhqsr0F0Sj8KXL/x7CWPT154C1vwR9Xmqrnv
QZPMNQOcBUa2HofvaG45CdDjtFsV3Sdw6D9NHyjzN4wEgsRCFkhPLe5UzpAHNdEic/Q+uRUaI6Dj
bn5UhVPtvNHy/4bkzsd5xy9hMuvrL6HpzBTM1fg8dYaPkXUkExQoMicDXF3PyYeaKf/n6koN4MOM
H/w+XmKsywECifjg1uiJY/9YaE1fz0hgIeycDVfHANQEE4kUArKSalSTc5DPlpJslbu5QbgUEytJ
5ZNE3NNEdBsZ37HpwOSchLCNYRXcLgAbEk63rWVlGb/RN0w+1yuZTGTJivaIdf9n570yybwO4Z27
8o4233KIvuFbyPzXilhOJDs7m9OPgXdmxkeurB/0tSQ4ZmqgZihPXgQVWD727svIkR1OyaodIh0u
q3yRWO9blolcoc/a29oCqkMePBYUmIsW8GDPh03s37Yb0tOJVbRkjZ2A+gvwC/eACYSEsRXTieeB
HDjgxP1KiiqSLceJsypBqosbmjrJQXe0gQRVddKNRna2OOX9zstMpraSGAERLfHbMXxR8v43p4BN
ZtybN/P15fPa9xgqIA4C15EwuiqORC5xCGgGwPijDClEvA4+lfu0JXifoLVkZj2WEje/1LVwVQqF
BKzN8/mP7Xmaym8/vjPGvhTZUEoSg9dB6vo5Ef8eP0zcfxj+Fy5pqv/cIM+lJZOB1wtKUlW24C8w
uwHmiBcXZpM8KN2XLOo+xo2/3/54YXLCwdCQRzav1lzkRUfzhr0sAp1LODMFhgZRltsszI5pg3ZT
d9pR+jM64u3/TIv5e6x68rpvJcYQoH8rPCFTkjt6FrXDvimu17PGWftC1YkfVgSYMo+rjLZr9Iin
Q8rjZDI08L1y6N7Kg1xq5JWNsEgiNAOr4p2BsY5vh6mONm+XkI84A8TQZujOZItLeZVYdW1UlfQi
dAoRlikEnsSw8tjxY9tkjsHJMctlMOJbgt9nWQ9Bv0MFt6T4hh9KJBvXnBEP2Frr3MEmg8e19tMt
5vNK4j3hBVwMyKSoH/YsgrmuFdTJ3DxD5i6gsLJKZBtjWah7/YsSZxo3uD8SmiiBofjCQvLxCwRh
QCj4xAIgFs/0KJQLp2C1TLg1gQjbxY3uLsbQyPY86QHBP5LhKNDkXclwFewk1uVnZxoCvCzlWfw7
DB38QGFQoXYT94kdgrUELVhXOydp55fiMCx5x7SXj/HGa/t5rnrTjhK7Im1iWW+fdfYuvHwEbl07
yAzI2dL9rdmzEayl2ri4rafzcYaToiM5QR3I78ql2lueuc8dFCJXfkGJ4StQQ/H9uWFElF6bTS4x
4cmBo2dz1yU2vj8l9s45FKR0XEA6NyiULYoaZw2poAmWQFlzGZmQoMitZvXHNqRZ2yuUipnclpUI
mFoDroq1Xm1lid/4TDongkjGbdEcww6OYBWNRRxws4zK6h3rnbXk7TAlH45AErhh7yf9fdtpY0iL
0DaQIOYKThauU76lCZPUxkNIlgSnHjLlj17YoQ+8LONGFG254CLpUKJaZ9cd0IHMEFTFBzGp/fdI
ZEJfXXk6mFKBW/v7991ewk8q72gbNXxL8g47/9H0eGPwSwOxuFa5X9gGKqqSyo+Ml6CaAitjYomC
yP4KdC34B9081gjFqtu+75AloTj49EM+xwKb8H+L95rmVvr+gask0KTdJrPE/NgnqJsGOzbaJsyB
FtWqNwyl+8qo23EBszmhpOAzy6kFbDuz18sEebMPpV37EVMPo2jb+qawnG3PbuJfZvj44LNo8laR
SsXnqjKyzKoXG/OaafECFRzPc2UiuweAH5KZyhWEzhimheSCqfSywjC3UfknTA0IbAIxDiPYrRvu
9PlVwftFJLYtQT9JNfM1awTnquqeELxIxXYgAc4wgXKqLTXodCLnuGLAgfF3MpN8JOLdWa+f8EUr
psWYRY4BBOwAY5Ibr63Rz34eAnUMpkx0eWU44YLAv69rRPWfXsArbCmCOK9tCvF/KUVncOOURzwJ
WvrTsd/w1E2SnxC5VqZp/V4m4x7L14aP5Vp7V0UiVp5Rwpv9HGSqYYtDjcg1B10NL462x8Lxjohc
zKAdcfLxwW37BfW+09BlNuFzHLbJJYz9ZqqIVIqFh/Oc0QeDsRXQddhrOBfF3xvORe4dKcpOmcpq
8MalAvoj4VXiqCBf9u7vVXl1odCRn0FV1/AkURapBfW6XsuldHEP0cPf+Gi6mz4XIDF2mWlVVlKn
Vqhpvl7pe/Atr2mX48kCW4uF5/alHKKZRSf1kmM1BrcZyHA5w+KquY7xe3Npg4SfaLq3DARMKNBo
uU920b1p94++oXbsgIHjrT1X17oxsUqUb2SrUmwRsm97ejtY8UZ/o1o+HkW39SS6HjR4NXIjaohG
A88JyIOwlNaYcx5GmOt/OfuyA2Fn3PMPJddU8fMLBUEKFrzRoOdAwwq2bcPJCYcztT4Rbqri0gnm
idWH0x4tEhQhiwwaPrOuBKt7ai3WCW53PC6hMSdwOd8r5Xge7U1xDLG5l3npjeEWoeWrYwvIq901
AhwvjzCtviKP8FGxWTVlkcD1821lMBlY42na5gyw/bkHLohwxWb0cFojh08N+WwJFZ7XX0UUO4bU
NJ/kl9qgIA2ypfLMvIGN2soXQyxPad3IO95mZh4VLMrcSpRDhqrpCL8aW11iKfRsA1HuyTxQGhsZ
/vMEs8YATQ+t3orbWy3a/HAN3QqZPB/lf0TjzRowawyvWJkd0T6jRIyZdXqjKCadLC+fk88ikmjs
C+oWBwyNXDN9ZaLKW8w4Gsh5Q9fit4FY2hiltooaTuqLwMo+2uRUtUaP4PzMclRjQyhIGKG24WyX
p+QqT8V2Wpvg5/glsus5KLGVtpXPqqhP2ll6ugwr1qnUnKooTM/JY3FyIPhi3YQAaIWMcu3JA+6F
n87qOfSb4sAiiM3LAVLz4lt9cmNztkQjzhhoJAHYbp66I25RYDM6Q65HomHLaoNtJZY72i3NBx9Z
MZoiuWDNflKG5+meAd4BClZnh9fwOsCwG8uOTvB3ljZPMFvSoANE23nQvyGYBPgWpMc15ggzkLZA
BIX/4/cLGsGzXRwoX/Z3122RfS246ivC6n5iDIRwykk0ajHVUCgXQ/2+IKAtXGvYwMyKG3l0RY2e
0yANK7L+EmBLhjxWb0xO+0mkCVZ0gmqKvbS8c4ES8mUA6Nsa9reDm/04nLCdPI/DllWX6Xm5gpi4
Xl7Od4zJgCp9DP9/3nw8Kj9QkH/36z0iKbpIhg3FVit+nuh0dtSYb2GdeHVR+XuoDeMgPatMK1HQ
r0WmkU33R27ueAguvAFArGHaCqx/j7lDdFNFr8ykHIDHlATC3aIh+Pu1Su0b6PG0ZEfyyFYogcnx
D2lzxjv9jgADEyBkvp6K4CBhYG3pL1EHsD6UEhAI4i1MuV/S/Jmof3209G4rXiuzdYWdLV90/u6g
n5/ba77pBRm3PkmcXwdawl5FkyAT7DChBZXY1kTfvT4r0/s/VSk0gn2hYYT/1hWcAv0XiOLIU89+
pgW56sBScyjWgFgwaP+T7yG+nVi4JIgL1iiXuD36+GS9m8VjUwmzNt9y0LknXpOuA4jHjFQZPqb5
RsaL/dBkF9hwkNRO2rD8K2kCjVBRyw5wlWNJgtSo/b15kB/5n9F7YxlYw4CYu4RCFXkdbvIcpz4t
or993ZKba213IFH8EXC6BUT7BXIYt5GHfbp6+y8IaMrNNWtFvJQp8QJLeUqSFIWaVeb1PppOAFAw
eZVJE27RljMvupL+NLhJUrj4FCjp2T16QM2rtvHyirtHJej/CeiZqNdFP570zlAGTP1lnWVactPc
+etyL9dCgrNRX97C8VvN14zminTES2XeyQEAnla8VhW3fVce8Ak0UKY+dyF5XLqsD9n1S0kjL3dG
Ki6lSuwqo1YgsjK61x+Hk6W2apblYxNFTvYV8Te4KU46GYlfnkF2yPviK56ChV091u+LyVhlIYt6
NOF8kScvVOpXFbQcnMCIB72lYV7NhdF84OSWg+qIGDDaesjF/q3v4LcP/VZV6TZPDbrTP568wtY4
2QdyNoAnpCi+in4PwEmzUGxi3jx7YfIWgWlwTzhoJGNOzyLwwaFsqZlILw18h4Tj0XEpouGR0z2c
xq15V4A0Dy2JgWYHRQ+2MWQSyy/W8wh8UWqxL66599HP7DS2uE8gtPHWmAvFmXUPNzeIiJdqSDRy
r75S5QzgQYvJNs/qFrxpsTSmTI1wmanU3cGLcTXLmjNAkXg1OWtFqbHCKyvb6oYRSAfvdHeV4o1y
aX+96hM9NMaKG5UMfExYV24fTI4WAkRvOIex90sjPTdCpYUNBTSaX83rOA6N9UYgYrwkU/Qn4Huy
HiJ0Lt3ZkjQuN4gUDsjlPyINKuxtGcuZ+ser9ZHVQahipF1Poovt9pu2tZR7IqE+PDwcyMLP+GJt
goh4siYVPLZir0prLLongDA5CatJQ9McAvC8t5nD7tTJCf/MJIERvwfwhIlbUHMUE3YCYyGjqOcR
S7Hc5VPfku1xVwFVuybrmz4uNY4E4Lf1r2ZfyaRB4v1a4poVMihoaJEIBO+8sTSRaixfpRa25gLr
R3/ZdKcExczBILpdPYblsHNknFthq9IfUvtoqWMZ1Dstj36FYArzVcDbr4Qu2r15Dmw7XF8qNvmm
KT72GSzWwypVY/aCnnRE7c0pEcvw6JBqTlMYWeOpqn4J8QmohF5Djw33xC0Mi/DmySnowKyhs9QQ
xAysJtiIfsxAtx+0JsReA1G6b5lemLSL6h/sTp4vouUoNF1yvWxRJ3KtXct9Iighav2Uyl9SdpFM
zAeQZnpBohV8CPRGe8chH6nVBL/lWTaZ+IMNeArlVP0rMNCTzFpfB/KLbx+FXWiCA+xV8x7xfuPv
IoUcnzqRRtTp/5hcpbGppZ7sMt7XWdIKDzxwzROADD7jwATNqV3iifjUEIJ2rja9xcdqGkQZTQxb
zMWqK2oL59vIjRLuxcBXOH7xfaOl1SBs5elWr+lSrlPDmVl74k/ph48ZW0kY/ZeaAzhXhsAgCbV4
IaVj0QO75V72u2CZ13XEBf25A/QMqtIKX0SZdbMoznUsw00X7elNhaErUNp1SeFo41ww0IHTl6Tb
SR2/xAIx9yT4GILxjdnsa5LmDo7oTAjmxyUMl+Ckro7VLl5CT6gd3BdHCM3eaFdldkyaR23RB8pq
b8mz4t4yu0+YHb/EQMcCjp8U5iKawltOQsYPsgsReLxUg/F8CSATqhBA2FXXq+VVsXofywlgPhkq
1qEOPAo1ZrAAvrpaRpLZCjBbC1qBoJ4dgMaE4IG3UpOfUCgDUQUl/MuRz1KwT23IGcwe3Tcsw7bX
9rzbc3YczAgaqHwHiZnQMjYUbPm0noFhdFElZedi/s1bNSe79FH7FyApx9IxOAKVAh51cbNfVUXv
LyVmNoOZn7tdHCeqq1HZcdooX4NqSXZ1fa1b6l0/dKuvcb/zekagrqsgc92Rxu3CiNIduTvw0NOL
YIjrc9BZF4pAXtZeHZPTmTM/TuPpZc5/4ixOoM9J+nvZGhpXTwnqqqmR1PW8Npb8JHuRoYj2ZYNR
+VzD3wqJSrOslkJnZ08znSSUACrRD8jmXLxoge1JL1rNZYEVdyCIiqkkxdPL4E23EVy5aXt67NHk
LZGJBYYAihp06EUll3VtbNC9jF8zQPDBkLmhmHJ32tJbisjRy+57oYw0OXa9t/0T9+kX1fl45qYG
+aqlvyJbJ/iJ3huSZKi+/EhMf1cMSIRpaSb+yT6KgYVb2eCj834nTLmIByFt4659wc93IfWaOtNB
dC+6hH2Ohc95xFnU5WzPXTULRRje9+aw/DZI5N+jy1avDXXPwpC2av6xFAyQ/wPj3wLRMSqJD6+K
k61W6SAx1nalxlufWcCKW8tb63lnvA7Du0RJhNSXO+ZM95dHzqwg6WHGlrLtl6CwA1JohjqAqFvb
O/ggAMLhav3jB2skofdd2bHRxNwqxseCWfVRwDB2CVIL1V+H2iq/zNHvHSXduhf2UUo2k8Ro+bEw
wHrALTdgAyvuD+PN+uINb4BJtbeb5JdXMBWmcoAiC2zSqlN8msw33/rpAGSAB0mxWbvRiZxN/0vz
/7j31RvMsVIqukGUWbo/LLXY/mhCLomMzbNDueGAmk1p6dHCybnShn4uc6sPuGSxpE8eaPquDus4
zZ4yRqFt17xVlvdyuJf32I6dyPpzCuSFd/ZsyjtddcY2rxXGdatXFYsi+2u7BmgP3S/35LysVFjY
r5vEtPeht6GB8QWctxw+ca3FnI+BlpfPi6Si5SAD9wDwn/DN6x5bdmEqYsktS0bMRYxj+xdy2vn3
J0lkx4hBW9PgajDk4YyW4jcqZleVTKjvGLA4aNWsANADYZF9piHKIASURrB/gKuzw5GnzsQ7F0la
aDnKHECh4mpgbcLbNrPgNMSvOByWKWRvvQk3AxOod5KeC1N/dsxBRyOtiL8LVv0M0ddyIz4U/JXQ
kiWBJZYJR7beD4TODAvc5EIF1Y69DW6TqcHOYxY0Ly5dKevfnhdfVma81cXnvkySBD7i5N/MS8SU
0KK4ovmbYaPzxhgrIFZRJwH5VCzyZdWnN6zFhwkx46qN8LKnTTkUuqRIuEPmgh2bDwtz7fUOYSsU
pbKEdk5yQBeNposgSHuEId245VFscHpt9PepotC1eUAcIyQDZa3rjrFv3iRJnV+qnwzynAW3gssK
0Oc6W49kYnUpi7LJVvJtnMn/rfa3KBfm+S4LNOs06rl8lzBVGBFrq9q88vt0iOyH62yZrYTBbf7t
wN3zHZdGEXklijOYt5WtVOF4yGFRnjIS2v6V5Sk1+NViUnaeDYXekSxyda9YPA6kPsuMc8C3qr34
jIT37cWgU1iEM+vGOPth+4h+RuIJsqG04imLqUjBU6EBmGtUC2uztyhVlf01LClNVrG64AvVFBFR
dsSwMOI+UgnZhOQo2QJb9JRrYfsFcmPb367Y4ItZ++JmGKnIoThr90ikPW5UWIkAkVFLjJftSU8n
aELL2lvjGg9Kb5IPgRcybSxc+P72ThbONLGjguCei59zKJNvz1ZdA9rK9Sooez+Afv8jd5xlxkUD
iiWYSYvY9u3kct4LzTg2BucdjX9C5Kr2sXA2zws/qWVl8+VPDYlEA3MKRtgqB8JHkBreq1JzTFhi
nfDniB82HFLgO1Q5GdjpDvg6b4W+ptJrZq218A8zeq6O2AcCJ2pUgloayg5ar8aJDuHB36G3gMIh
THdzunO8ESHbMeTiXX+WP9vmmfMwebixTAgBtvfnGDYiYFWzGt7zFaqvCMV/atFOCw9yzB7p+jQJ
uRGruZ5ScSX2xcCx5/8Qo555CFsi7zTeoYjJzFuG2hnIFVm5HTwPZhrRtGs24VY+WS/QbpIBzuCD
1XXzqDuRu+3dZJgXuVfpD6VC9yJzkEmu/12mxdunMzy4XxnXec4QsxFTuF/Z/wY/oBieLhF2Awnb
dzjMQo6XfNnXsfAHLHiUAkhcO8G/DGGCiQ+0JBzC4A7WPtt3HeJ+C9n8r+EEDHyxUp2+LTlm2pEU
mxJXeAgC/iQ0wQlFsa/bAYMFvsKLuZDoIlJUWciWqZdw6jWFx0OJB5kJNhTDSkUwxzpKNVMkZIHa
HJnUeEuZCMqJmnEJl4Y6152waCpPFTDZZDyrYmztmV4iDM+nIQSPpJrFhXmZQUkoQMz1o5UClZfJ
1piPUKo69lyKRWwaXEteARDdJh/IrSjkzl1yDWDRVwmnJXc3O/E/+rZGiqE/SnsjCauBbnsPS74f
W9lxK1G7pjmrbaFU66F/0f7PYHyvzcUzJ2MtWH0/Nm/b8drvmWeruPIlDQ==
`protect end_protected

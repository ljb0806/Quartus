��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�C2��~��?f1ĭB\1�r`T�Sb�p���0XQ)���s�f?(k�J&V�����u;T"�i;�T���z{����,�+0�;uO+�,�;L��[�-R���`�-�<�S�ګ�D����"��
ԟY�S{�!]��|�?3�_���ά�zVY�)I! �4���4�bq�-����O[H|J�ñ��ya����r��s���v�+�]�	^	��,WM�/�f�g�UpL G�N����Q�x&F��D{�si�>�%�`�.�\�a-i���2��5h�/��4*�*m�C?�$/C�˜�BH�q�x0�S�t`��AQݩ+2�[���������pH��~9����NouWe����O�(�/�ս&$�f�Tea��+�~ E�<�-�,�l	]������v���L�K�\�n�I��f����ëow;خ2�Q$��|�~��g/�b�+������sJf�>9����^
S�v��W��㻏P8�D񹊖k��e��e��;�)ŀ�a����(���hC����BY;� �zDçS���-yQ��N�J�gYT<��XŚ�l>�%��쐠!6T,�/����қ�j��5�wPIL�),�ΑS��DǸA���J�S��7T�1��h�G}1�f���
�:uc͖o�U�@:�ٍj�ĢD�O7ܺ!�}�L�8:zy�� ~�Z>^{ ��ܵ�՘�N�������Z�ڞD[o_[ፇ<���M�j�:ML���-�شp��Y����d�����'�	DG������������7�~�햰�zC_��-��a���`�_����4� ���p]�2�E'��N�<����V*|�*-� D��ׅIт�m��H�󉕡�}
A]���g��`�����q=n�k�c�6�~�$�Gv�$�_kߣ�?g:��4��=F��Lg�	Ԟ��id1���|5gO//!G�Чb��^�:-7�:�l���E;�q0���r#t,�[��$����nYn�Miq�����ӵ��I3�=�����$�}���|K�^�vW(��yQ��G^	(�����J��㗇����cM~��I\���ܺ�Jق�E��SH�a�Q�9�Fj�Y�
��w>/Ӥ�ݹt���p���jt	�V���9�?�)�(�5w�c�ħ܍����z���T;�d/��4O��=L��]����;v;Ra����Gk�	�g���fo嶾�
������Ei?�|�U~�Dm��-"2s��i6��M}�h��� �g�����O|���K�_R�5���Y1.$`݌0�(r�.�G֨�����g���� x-��t���N~�!"�Jd4��O8.2t������PQʽ�>}:������L:�q�3��Ka���]����|�$��H(� hD��A�%�v/**�X`�5��Z�T��L2�$���[/�/���7�R��^l�G��בͻ7�F�+xRw;�wQ�FH
7�H��
�C�T���I�N���{��_�,|��$#'���Sm_��x�~R���]!��P��	L���Q7(md�5A8�}!8�ų�� ���&皛�G���c����q0��7UÜ�z?/�b�{��x�#�Y������uM L�84�&�K'=�y�?��+!�?��ePН�O%�$;DY����V����v�h�
a�E_��2T��C�Z�=���X�5�]�A�Y���^,�+���n~Sz�����  o�Sld}~��}�H>����[�m���bI�
�·�Q���GR����	�"&XG>^�qX�H:��9�;�8eW�je�&1p�7���%{�:@�^�Dd7��؅����J��Kڕ�Rp��B���O�]�0�ں�V�;4���3���)�];�υ��S��uxVI]�HL�x�ح@~�)9��A���2+6A"+K����!L `,i��P�Y��Օ{����1JX�L�>e�Z�����Uo,�E�>y�(s����Y���y��c�ʡY�>P���G��9�0ﷆ�?j|���uo��n�ʣф��kA�\�墱�5�գ�j/b��J���/�n�N*�Ƣ�dĨׯϛ�&�Hl�:�����f9�r)}	�2��wc?$bG�ʃ(ӮI��g���q=�zkp_���K����?TRr�9?rd �hU ��v��
pHݺ�������в�(m���;��_o{��$1L;u�1�?��!K���ګ���Y��&\����$7�K#��ΦFh�s��.,-Ƥi� ND��땬+���*���y��BO7�]8*n%�*��@w��l��[��&D�*��>7U�mI�e�V国����6��7�ᑅ7����$x�O��Ж##�k�y�@�N��@h��7�x_(F�aX���C�Sl��J=9��S��#e�/-�v�2�|�� ��W�[F?��@#���d*�9����%s�^ha�q��������}�����!G�0��)�yς����;U���x��1�/�e�>�X#��W�zh�'�R_���1Y��)��t������l�m�fޘ�e�;�e%�P�(�>�Z^���9��]eC�eeѴ �";�H	�o��w�����5���Yc��e5C�����Zۅ��A<o���$C5)uw��%��n������i�i�9n_���<B;�ˢ�hMl_���<N2�R���x~{c@W�6
�����ʁ3�
�/��qq��[�1	⑩Bk�u$1����{�P��p��g��E�xs��z�Tގk{��<�/nj�N�h9@��B�4	Q�A!e~8Q��&`����h��07���f7��P̓Pܮ�@���zw�΀n)�����}0]ǚ��!��W����k�d� 7#���
+�ڃ,t`T����ʬ��(����O��w�6�T�U'�bN��ޫqAl�'M��%D���r��x��z.�����XV������,{��Rv6�@��+��q4�TQ������\�?	�C6�?-��ޢ����=-`D���F�Ad�IƤjg��X2�x΃'<oIST��6Ok�ۅ]aZ0I�&��)����B�Z�	.r�I$�����kX��PY�8uMo(�w!��$�Ь��7Ρ�"Qcui����ۢ�qC�d�u
�t� �֥�V��e�䗔^���"v�w;���i��3���}"1�t���d�D��MZ8��L��cW���=Gw,�:�n��j��l������dcK��n�l�<�w^�Aħ���|h��fd۰�vj�|�Ɩ 	{��\�g�$�%�z�����x<�~�tS��M��Bh��Ƈ��9x0���j����M��5�&r�_9�kc,}]��^�p=h;R�_��RB�E�-�%��ؽ����Xu�{��'�h����V[�ºpCE���i|��a�簧8�w��7�D�2[���?`ۡ9�.\4�9ZRHJK�HXCO�L(��T5rTJ.�^ t�9:E���_IkC�o]D�Jx��o�s6���*4��Z�O�����%k9J"��w�F��I��Wj
o/���
|��W���4x����ؾxm�@܃ ���0�:>R}��"«�6]�����wk�w?�M����QMӖ��~d/퀾w�&�s��BjV~Х�)r! :v�\��1g�*�8�1L5R,�Z��^+�	�2�A�ήo�6��2�{���ݒ�'^�,�d��3�9���������ÿ��gH<Y/�-\�'2Q5��D�h{LJ�|�(J�0~l���^$�B/Q��������9`׵>@gu���}���2fr���D́sR��~�	���w|˿�H�*z��K'�B�}�x�~��f�{3���b%l"
����Q�L����\6����jf��!j��_����sҋ�1W�}5
GtdMn>�`��8!³�A�a &6=��le͊JS,��\�q�#4��b8O~Ⱥ;�U�a��)���(t�sh���v-wA�Y�_�R�
�?-x �Q�B$��t`���_�j��a���@�S��(,+�'�	VgP#QI#�s=Y �Q���r��v�Ѿ���LP��_��4!j���w"�jk���uc��_�
-�n�oY�ƣ�V!\ʐN��ȋ����l �Gi���Ak�{x!}i�6f�C*2�t�`~5D�'�v��pΐ[�ˁ{�X�o~
���
��R�ڄ��g�	ж�WVk;k�w-.%	Z�6�%W�.}��9ǟU�z��-X�>l�,���DOy���.�&��Sc�-r��vB��vL�԰�s�w�!)��[E�dP��9k�6�}�4 K�`���:�s2�����p��(}	˼{��d_��h&(�%�MoV 'sb���u'�,c0<U7�kQ�G�h,�~�?���	bq�/��[\�)wt������j���<`��K����E���F<�}�����p�زL��7��.�=��_QJ}>�Į�B��b�9x��.�$h��Us$+*V��[�W?$!E?����=h��uV	���?*��#4�=eh��Bxժ�"�L�Fы�T � ��C�2�ꪠq�*2d�ճ�54�m�3�f�2���j	�UHT����t��y�G��I!�uP����}�c�ь�T�"k2z�������6�Z���)c  ���I�3���E��1�}���te^<T2�Ɂ��
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
m9poasoODkgqGfefPzz9iGh+6CB99wIY2tiA+fEKEAoQ3REfJWogjHk4zDZQUTFNkpY79oNyawU+
GMlZl73DxY7PJes5/20H7AwHW+OULgsAJTSC9j4M7IXkYVkt/cr/NUMt5PmYhPA8pnNKBm4ijzQA
OT+VwiJFvZ4C2XsImrUJGnAIsmHVhZE2xd1LZsOATEahZIypd6EVJohY/CXcfo09/WacKenFRhu9
hi+VcjB+y4QmiQDlcMQcJuMgiQ6Br9JDVVmuD3m4PTxa2I1S5luXM2L0e6soywESnK1RzjDk/MKi
rY7IzxAv99psfbwAP6rfdzWpLoQp02nx/YlnYw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13440)
`protect data_block
0c+2oXFDDu0GlihaqQUW3s0IVSPe07a3ptlYCoy07Nyb2JsT3QIa+2MEUtBuHdkUWcYqwemkvzlY
7AwyOoKeY/MVue+0dL2Wh5QMIAR/4vu+gxEnPjQNciHG+moQTpplhorFDOZjkxWhWAz0URL/3c0D
8R6nxccHIsrimZuCewZ6BIIfACzcO/QzM+wkT8Vb5tRZXkb24lbKD8mi6JYIcFQDOVBN0fwYzu4J
YWH/nk+ym3aQ3HhNk0y4fnRjJCuPBv6pems57SB1NZfI/hmVNDoqJrs+4oZNtdCO11sXJKOnIyAk
C9ziFoCTSCasOm0enZIUaXZSeBoRF8kkRPAhJ1WiiDz/BaqOSUgfzVadrl5LnynJB2O5TCut0abs
mHXXQMNjBL5+uqMBaVVCVN12L8NopuAuHxgouelMsWAQsdX/O/GZzKJOEMbB+7dcC2tsKuqMLopn
7uYAWccKDju/5wdRCLiEfJgwyL7pTvlVrvJJSmFRO3C8nSZIj6IeQKyLpv7SgPRZqXAUrXWjLFTa
OcOdUdLnSNTm3/LSC/zZRmSazHiCd/TTxL4oi6KxaLS6nUoPEN49FwYLvOv6jsiRtVivc8ORbwfX
6AUJ3f+qYhZji8TQmBimsyoOQIHLAhdVVm+Q8VHOLF0AHQqCVSC+ZLjoCEHjUeeE0B8emVx4Ks3r
AZ/oOh6MwxsVgI77wZVDBplMmfqz+iWyJgy+gOex5wgswsOC7axjxPYfaxMeknXW6zHG0Yp+vDvE
xdDnmzo1LAYCB7wglvUaiJoCiH6ctuNdxUqAFlJys4yRs3Da26R6ZBq/wIiu8OISeLQFA45fbzut
3oR3lwe23kFz4THlmocIerKarb+dHnBYFZqMOCA75Z/fnFjEz0MAeMKQsAGKCXZVBreMuswgUYx2
6PzbHbdt5M7PAYSb7oSfFeZ7g9NcubuhqDsnFLS+qBnRboGnR6Zh1cmTgrHKOt9/R74XfhxBxHLE
6WwTmNXlgnCFcmsv23cktkgoIKIcVu/my9wXpV0/+7g+JqHuorciFMdxl6ZQUpUUKKvi05wxdZ0v
mKVrsv6FiX5Tey+UJRr5fOhIUfUHudZAtfTtKWhUV9kKtxucNJXNCiMkXimVqJNr/frDUb+mG337
qeEdcL/eVLs3AhFpBvCdIJsoqtBGcZ32/+905HBekedKXKy2FtLIXq+FDf1NxYuTwbNhdOeOBOx4
FPC1rboT/7uWNaUMP0EW6gLAj4R8FdM04zwMqBCS7O5uzog78fZ/gO9vRQd730cTJSsnUxYxJQpL
owcoXmdCzQ8wAFRdjnGBWAgw2Kfp/zDBNxxSDohJ+kRtNmjOm/g1ZsYoGa2JudD8B+w6AQI20HnQ
6H2pbOGFUVO9ClCE6tbXzYqYuaQV9IP/Tm10iFqA0tJPlFHmZ9ONERRagp3S2qaPxw77xlQL3uTL
SIL7vm4cJOI8GnNuWdkmGQL6IQ6jDVEmaTnsRtYt9JFkwKPRk36ED6WJL0VtMiHNNUfFHF/Fi8oJ
Rd3jhesAUTFNzb82HU/8PMTNLa6YhGOHIFZIqz8z4g/+6yv+hH83FpFHjbtLDdKpJJq4zVENBNlT
CY1BD0HWU9kWjVztYMTI/fXxDKiuvd6z/RJpxssvXRUaCJ+Ejkfui1kQfJhrZnPtHsZatn27r80T
kDRO4wrkplPpdSeag18ldN2JflLaKQckJ7gwV6QltAD9F3Rv4f2MfxteHwLw2EoCc24oj1uziYFU
l+DDUaGA3yWWRdLHyGzHMKq2wsilnPqtoRq5erCtW6eFA8UMkEym6vhenUDhh/z17lUvy2nlT82t
WZ8mziINVGbRdhvSn3ZtmNFjv70/ud5Zul1K0x/5mkXb/LeBMaXzKjNVNzDyrPpaEdRI7EllAhY0
gtzbL7wNb2d/RY/MygPY5G7wXGHMkKjf0uuC2nn3qeDxJGXg84EBihqlU+QioxsQI+ZlVfRh1rPu
ndKrjzryQUUFqtq9ryZg0RGyHGKa8B5VMM9kcwV0JdPzxXuXLMbX/Rx3DUyshQHglH3vX/lLRYb/
ydpBBtSixXEBeu7anxMIZezYiEgunjkQ/Iw1u6/vUloJhJtOzc7bsgxeNSLw4PJZXGcZG5IHCZ0U
nDZhG8d0UnZv7yR8CTj8L354C7ardV8b/CMOQxAqEGMwb9LT/8L9+v/ExkWPldC0h/u2+b0+jMiG
L90Os/GlNKP/JTWyNjAXH3Z8W/f/0Crj4RuB4us1F3+WfTWc1lXfP+SZGILLiCKPOoNX6z+1pB0X
QOSLfHzbdYZJSTr83dTP9q2pJm8WTcC35xSo5p86xol0HHgNf/D+jZ6JUc4APfExzJBfyG7SHSfR
G9lndRYA6tJagf+QZcw7E2I5lzA6YqMGIW3FB4sU6NEtTHuqtYeeaEzsNQhzrjuWHXk9Q6sf9N21
m6LyhVNkBekzf2qyUSO4TNOj40vaE/QLNLaeb8yZN9j1oBsTtH2B4B20NOBqhkhqxJEfe7bjW5wU
nDTDABEdyRHdRBN0kI3+F4sS+V9/PrEJqt2Ayh7Gta+pZvp9YDtCRIXxy28N3o9npIi1ORUPwWnc
3e6AQsxq1MluBF1D6atUlcuEkh+qFeTZk6Kp8wgPiKnuPQ2oHprykiaH7HatJ/uR2pDgqkQCll37
C9BMa52mGy2VubW4njI6j5h3yIE/xivY4a18hybhbbJT5og+tAxA3iGajTPz6b9bGo+SELkDnqHf
nIA+X1IlRoofIrKBzXsnDjdzitAU+HH9rKDdYNgAfE4xwwH+bU/JJb0CZYPJcn5NyfxBf1nZeHYu
J8JJ/qcPViQZ7963b+poZ9+6Fnq9n3zuX+ckzExyA475KHQK6tX3ooNlvNdUv7vaxn9/A35bz+hI
qdKH5pE6UfrgCd4K8mEJvSdAbKGCk3McYOLtXtuNwhS05GtGW5fAHkzd6LSmk0B4FXlBWKbI/TLw
sv8OPvFKdpMLzbelytehAhbPCgR3PXduwxafFQ31m/y71rkBOMeQTylZRVQ3+S3e6d4z8I1ZSAcb
Zb6AvXcZD3bpeX9VQPgB/7SiilkPy6LWIMzq0EDgz04WqhLkLovfRo0OCY/tI4QCIjMIvxT4KuJ8
3TtDcpDr7adi4yEnhBw+C85OaD39k+TyGwIGIr+zN/etHI9YfDzKrwaQp3wapMWUrvUKJuuODYXM
S5kx4uJKVelR6/RzQjE4pRWtEj0pma74fUcdqZJV3sMSfUmLicjBUyQx9cic8+JrMibxATaxczws
hC3ILNhmveirUXJJ8uf4BmVDg31jZk00b3dOAw9Hsn65UJNrIYYofrqiXEHDAzkgpUYp3T1uauUS
LDWd/NCbV4SDqKunABN6t7YeCPw7j+2yvLXMSJ+2Fw/Ryoi6fLBWEy7MVQEGOdwWnS5i9fcQGvrd
1SFaR1QXOdsCnu1MHxQNZHAt0hrNc3GLfErNF5/sAbznmNKlwaqwMgWDL4yNBdQCstMluBj3jqh9
1DkK+zvdOPIYQAQOI9EyuwgpQFyhMsMT8FAq9/fil1YkViwGJZXYXDntXuRgZzhvxKYfe7BAn6wR
PEh2LeQpl/xfrWV3b/0+lpj+LD3qMMvdGyyCK+xu8XVzs4yc47mTBENmqspoJS4A3GDOWOJMvrUu
WlwDxglSJU9Tq0whkt/VTJF5Ka6dxGx4bjiAP/8luYLdsvNwWl8KEEgLswldMZ+27fmcLw+AUOKr
XR9Su7mY3vgYgHWSC4MztSjpQqiB4HTCH3d2ZJZ9fnfLgLuGsU0DuzEpSGpqUcat4DeHUL/tTuqu
VbcPgUDLDw32GY1mlyv9ec0S3wQOE4EctHcg72Uc4hB7GpDOg3ErGWYrBjy0eho1dF3lrV7DJa6T
UbSXiL92QdcBr0kz5PJUkNUNpFD5aj/fADwwBwB7WmNYcl2DpK0563LCkG3LILVB0Xf2cS4YenSV
dGfOlmQIZQBQie5cMKEoN279+j9agN0DFg9S5DIIizkI6DVxyi3rhi5JneX9jQGQ2N0za82cWxRH
95tsh9E5yUzfC5dWUYn+J0rNBMXbjDuHE1t30bA8suSqAfKo8WnIbRylUSFzpxP4ma6lMRE10LRB
bMRU0qis4C+Z1LGbEwPo5ZZuANAlemKAmvbJQkoy+hgy0GfnCG3KvlhGxemBOPNC2JNamhLlO71K
VUD2vwB2q2SP/0EMKU53W5SWF1HshmebGGINEkCbApFHAupVHLxSx/EFPYvGCEnP/juWh79QMxCi
ITJEBRFpZqYRCM74PRnGHnch+O7ZrO0SI6yzZt1HHI5+Ku2RVeu+BTJvPuw8VCsN3UeoYLUCSI9d
FczqciHpOFx8l/oZx9+1J0GkGJJmKQq8sjM8gVn5IcjrjuI0lzbT7t2JpWXfFXTdP3KswEXM7IVM
z4oER9SzapQK6b30OYjI3nYZPDSJIKJWYi1XYvGU4WvvOkxc2711+8zbW2rZmpqE4YCwam37FimW
KVibHZZc1GEfRNZA/cvAhmhKSfz5LnWb33lh3iOAhr6lqmcieoD3XnQwPHm6vivnL2Q6T/JdNPYP
vBtVmwUabupfc2cVzcXGKQkOEp/Boo53qo80wvH55DtdGKvn6dWC7gauI9AkVLTUumvTiwAOUndG
Bn25hS/CnaSOvXIs/38DmqyMNA7Kwev2UutAD5Tb1U6LUf+H2qOnAaO56qifIZxOTWUj8WaR+pGg
4abJAsqzFa6LJnO0RyKufYuQ0UFPLuY/axZHvfdEOUOceDbo5KU1nNWFS7fSl280dtPlt1Enufam
8K/IzBlDQwIlqczw0gpKkessqCKVaDDVyV0Yex8Y7n49MXoNyBHZSApkMzV37Ilk96W8+MR8Na9i
pD9uyOHKb1SgRUrOCLH+rFLrNN3zFgtXdA3bb/9rQpPmLsFBGfcaCyikRb6JhqeGW3UeHNbf/tGb
/3qGrjlcVc076M6Agm81Shl37T52wat42TeUh2cDuvndiRCo6nm7gzUfS+BnN1XTVvs4SDyKE2id
GtrG4uYQWJmn/W2b/Xv4WbnGY1niOtJiqeeHM9C4ObODyGMDTcgpJ5jSIiufNo92BFYhRdXG56A8
m/FzbBgh3+beklLW/s7S27OcnbC2bHBDiGHxZKbFcBXxvEPBqeUceFpHxmt/obZRNDyki9Vxl8Mh
UTar1br47SmZpOPg9/T0quR7GcO6nMNUP3jhQMOfd6SosLpLRE5udJ6KQORU6babm3zHz3DCwaTX
bPPUdtkuYuHgmQSFVxW/c4pNPQOmtgyY7/KuPu6tm+3dDXdw/0A6vc9w+X9MAgCcH2LNdo665q7Z
ObLa9PJKHbFCQ3/Jf5BGSF9uRm5B8lX36rN6BXtPzRFDQz7XGfCEh0Rnzf2dy03Jr/WTH3jw4uKc
rYYhuA3HMZjHWeXG8seGh43HP1yJAG/OwoAN8K6Rwt/OvVTV7wvPlgfXSIbKMgtsNQmZnoLDBppR
EL6A72eyWvpZZw3ZNkOpK7hLRtV/W4CCEW8quoH25vmqgyR/oLiNOKSEZvcbwRS+G2SgW2WKAD4S
Nvn7/UKmy6SqBu4M7XOJykoFIYrPcINWCgC8oX5TJv9HHsAphzOd+pOXyv5qLDGDR9r9wOZhnIWT
Wscmf1N5ELo3J9UccJ2GH0pU2vJgtx+NvYrh8shSgbgEK8rgt+g92LYnT04dzQ4kQmZETcXEINgw
flIUoF19iV35DIQVzGfO2UIR2Zbi4qR1qNO3aFbktzySZMrCCwXZe0poF37n3+BEn4/73yrMTTHQ
AHw0g55wvXCkIDVE6Qy05czPGTtG4im3NleTbOrBGuMrjA00S2Et7iP8e1aO4ZNf6+POr7eVdNYv
vF8hFEYTZ48UYKIYCpRdV7B/Sgsj7X36Gm571ZS4LSctLcu28w+FA5wmJnYCYyuWtqQXU5uOx+Db
rg0DqzPP944gcdye+QDklw4e0bjnWPa3PG+bEkxQPRVFeHMPx3IYvM9N0gOi7+4/yGw+XJc09dC8
QO3HwsZqjMSsqL5t6cSrVv0soOSYaFALveBFZY4t8bLZVDHKsJjcEdd5vaSyaESOUY2rCGDmUBRn
IlMxpgPlcsEbcro/bdJqCUCx44VYjLTaXoRpROrkcLlW3LaH7h/DaUJ5j8JKYnkeHZS729vqOfF6
K6S63NLYnZn3w+AuwcKChFw/5KmvvSCPKukhcmJk1MSCsnyP6/rX2gkLG/fF8f5vL42ugXIO+02E
XDjdNwSgqFYAeuiuif2/9x1iJKrJCl+MEzbTXSBt3HLVvhX7pgG9VkpDRS5LjTD5d9FarGWO8tKN
ZJcGuqCOcU5eiyEd44EHQBBCOtrTolq8ccWh8z+i6cdifGYNY/Ogx4x5aGuhfx1T90KtsggzG2uL
oD433kjM9eU9S/kreBzx6M9DaSaJsJ98XyA2mKMggVyQtACK04uGFgwF8stEd7lfFSSg/O3uuhpS
vLRRLtkmA0+VdKrrdBEVeZHZYB1TXfppWlZgq7vL07J2vT1L52E+Yzl0fSpGJENfZS8BG2RDcYWL
Eveq7ueRHpfPd0emyoiI0OwLWqX8RWbmdR8j3xkHUu4lHpA6+CtCDMxoEISTPSY5vhaQv02RK3Dc
ncEQrcLT9CmNcbhKiPqIP9s0O7o9+Cu9b0pjdDpmsWPCFlWqGDGZOCwAGZC2bXh1VuQc+eeb5qqT
wg1UF72QwHmOIQXtuazYoRdrSufdhN355MieRJC1TvBmUyivL76r+gSo9YWW8aJ5HJLgD67zP7Ul
4qoly86MUGEVYf62bXd5ME1Mk6i9efZW0OdQzs9cdqyiOONbGyUtCUDAxvG84fIjdhC8vdaHb6+Z
rMfC9yWmuHA3IWVi7uqm/PXcBOTWCpOWP/liotF/J4K6IloaI77vRd22E2Kzdqi9HGAQb/a+wwai
k2yrK4+wUe1dtOFc7LH6tmZcf45TiqjNEeTLK11sUOUohqEAElK6ypTXhn8QdRA+41h8hGrkoUmY
LwmuiAl0d5xryCBADaXxNG2w0tXg/yWrUgBW7lZRlsn4OL3Jixr3ZPfqL2kevE4imisfpG7vToYg
sM/O2WwoTwCXozUYcnCkwUSrAWdQOQiyQaphfQAn29O+6O89j5CoZrHDCwQXqG101BvJSEdDbRjh
bE4Vl735vncRK8/W5+QG+XdkRwDG4QAnaw3AVVRSeuiYlyKGoAsniHfdqLnGiGXksDlhRIx2UV5X
fWyM5zwciCkkx+XKI0TfTelq6y4Kt/W0+XULF9yTC3pNCCY8V3jXExDqIXkI6FwjUVofrtidjZHo
QfXAPIlcra7FEWR7HQl/eZ2Q9ti//IoF9Wr0yauNFl0HYnd494cin4wVSdeTT2Cw5gGTKyFk2tbu
1xb40VY3mSuhRAaod9Bkwi5oIt7u5Yghu9MF4rahjIQOb5zAcRZzblYvWWhPxYJIUO+sCSp42/KK
9990DDiq4vMlwhjjmIgk4gqlbWeNJ+xB+6Bih8GpccnHDxcnZGoRGkoMZcA37KDxd4bPJ6jsGXkb
B+Aa2KcdjKAa1sYtYJxF2sY9Y/VSVG3XXGSjSaeKtTpJTy+a7/EuEyRj9uwZeahJMHYPrN2pvqYx
5ywpo0LKnKh6wWPzHEo+u7Az6ANyQbU9xRnu4Z8NhXmkTdurIoMjFfKBleP8BgGXNbD99aeoHM4o
2rvPJU6Tc0/xcNZz3Jm1W58ZQNDUM/fbknijcHg8taBKj8rehB+bxWXoSPf0sYTaWunDF0+wLCA2
7sZWb5D0yhSGd73Ow7WQqWChnN5YiRsahpJGgEOJeYUOxxQESwLQ80iFa0h+BzW/MgbM/vZRw5Td
K4hK3BxeF+eR2RiRdKbDrbrQxjMbMoTvVXmkZq0DQ94iJlCs7ikpTgYA7ri2gZb+WaM0hcd7Q5fP
GAkZi8mU7iTRnks8X9yqJs2DZuLOrtEiMfkHK5I7xKbVHzNRpz8j1lINGLQyGKRWbmFriU/O6MDH
fJSSD+TrNJ271lKXiZIcJZf59ig/wRky2io0APABDapsMwRH54G+y8Icfp42Ifmv+L7/9nJP4pAF
E84zIiDP87BdpXG5sqqzWOzKTIObfCIwCC/Gj85pL90exAQ4vDrlUX6E5SB1hTXu2vQFAV8ENCnO
vxj3/nw8VnM1YiELISa4YpVP9aRCYoSUzgwk+e/sEzfytqoNiRuSpeSIdOpjvONk5c5kydwvlz0R
YcullkZtZ5PeXx1QsSxS6mru1rR1qQ+EXSlyO/3R0QJMVChmEJ6bv3KUkKGZfnZSVMhxNe+co5Gv
6ZpyuMu83ZLhrEGDYHlSPB+fdFf6vlpWlFDADUbFOIk5PJKm+IZrp+ARpWuEGy48z9Zn0te+Un20
8SXWLRc5fZsjDJkth84LkAm9bIN0AtPmYuTfI7NwHJvIBZ/BVO5Pa8ZW+kYji5F1COe084gFyRmM
Jw/PBEmxF4IzILCtpkh36AM3aqRJlHhwp1PIHVNccPd+YxO8PCYxwi8kKjYOv1OA5WUDDDsq40C4
VSQfqMBq2VBhWZMPzl+ThaGKPxqnAutcbSlFwSc0H4Jw09JQvCZE3kayI0uG73JIDwWIcChm94Vt
yMMv/bX2oNjg+yVzkI/apG0vb+lNaF2LfgygNQdb5RL8EaRxnyA0IYSsb/yMbjI5d9WYdIjSa4e6
v8b8T+xacWiWkfHrK7pwwHy6OhGgf6aw4lq1GciY0jCrEzdaE6mxIT7/BuJrCDOS7x6hFKCLjahR
viytbcYVUkKCldRwDqAA9JFQTIh7vvXdSgGpmpl9L6gcy8cv3jLtuAa0krAMH19NHC9QyknYr3qE
AtkLPR4sGr700wDg+ArF+6mqH2llzJQlRtA7NRi8eGBUDaqkzRcG/6xVA6B8Ty7xPaswHqm8qEGp
uYdP0j0theiYSYuIpIMcxXWm9O+P9Qk+q+M98lnKtz6G8Ekk4nKIFo6+/qfviJI3Qm8U6APVFbWp
e+dfB6j0X3vZM5I/JIHREBoXxIoOlpkqLbdPMO0DyQ9dmUh7/7IWz3qnJlCjaBddgj4vdUp79Y6U
9xv9NCaCkZb1pDHAzQ214FFFkH4b+ZWf6u8fUx0r+vpU9VmGGqgTCMxT7gzeHROqR4fnjYBqW4EJ
w9dr2h5i/FtP3dBRVepqjv3neUY21WKNJFu+luz3qbytcoO3wsYBRHtCHjH/CV8iEXuYr6qrehKq
MsCcHWMDpzSQOql4GQiuWmClrzd5fn1nudAaiaLUZky/b9+8K2W4wzUBtye2ksFWZB3lN8nV6FZd
S1f5Cjaj7QDIsXM4xkGVOTPJvSyWgE9SfxIaMZkX+CTjggtlDCtSlx+jG1s2LrgYcLF+TyDjCOgZ
zIJP2JdYYzLfXwy2jg20tb7b4Tlvave+peVYcro3F04DdVsSociUarlx/c5E29fwhSRgvjdYaYoM
LIn6ZjophxtxT3pSUXH88weNtUZCaMvDgGm80y7ND0o8b+O93flGyQE33NOhKV7/lQSk9BRo6Ynr
pQzrENeJnw4lQquOlmJuk56rR8p8y4mbe8kTRj2AWtGA5CnimoDQlWeVIO/Qlrf4a3Z9911A39B5
Nv9RzjimnYN7uENgwURqeaiFP3S0lV96KKDpJK5SUux++7SxxLlzqGdWYDp9gbetkzyglrSM/zv2
Az7KpoKpzIdaUleCZaEbkd70Dc2L1x4RDk3igQ37U9K5deUYKby0bFDbL9F6XelwE46x0X7nJUZz
sAfTEo62lZlbuVUctrVzI+XqvaquH+kNrJ3WpnJK71wpYTDxTcHTCRjtNC01sS6x+nvSm1KrnvtA
UTqPkZStXUMeyc0Zdqu2BoJwYGU5rWcM0iGyFisllMAJnIYS325/0xOUx3JWgLK2p2vThaD1oS2n
b3uE/umPNxuewTVbOMD3ei9B4KKQhbZK5y+xS9v5aG4fAejgBPK1xpuq1uUcy7zrpJ5AdUSGiUQC
f0yn/5NK06yqBRwqt80PLgHsrBcWJ67ceuT1ZW9h8ZF60r+bFCG0mfVVBguKKzeFEhqYI51AKZLY
4+xqTpxcyJlRw8nGx9CpuddXvGjeRguVl5sDsTwg9g1ubnZzYHThYO/MbaWC9wQPn8dy/qi8D0YL
89H1wXcRtToIkguV+cvbdrWBWkVl62yBRzPBo4PgpxJMuPyJal4EsmULByztAuTEmr0PPsx28hCx
u1+fh8yexMaZOK+gyx0UgP8BPGCN426bEk/p1DsFxcsQlq5m3UpGPuhdaWeoAxnfCMb8YUc6yg0J
TfKDta53qyASGBdo86UWMRtSXXSbGUgES34hOSnQwqLcMKYXKDkAKSKJKoUbT5vZv7z/rnqP7U/+
g1gSuJhdkKWSJUhfwz1DCul3IAPSes3fUddVesQ1DT/rl+PGXiyw9oaKT+B9HTjxKt6u9d/QosZC
hkCWT5VigQnds3sspnC9FkuOF5behoSxE2z0DVSOe/YsSbF/Zo48V8vmFPw+dlUZOX26CEM6pEWZ
GlSdluFqEqZmp6ljOYfH9NnddioaQ9FzZwoaOXyb31dUSSrYUfqUkTdP024yl/j7pkhRjGO+DYCj
yaogBBX49HWkF5jGURx6LLwoQwyEdiXs/O+NU3nYJMXAz4ViF8uOnxgmcjIQnLyJwN8j+z6Goizn
GEGDq8TWYBzgRGB22oLiYxI2xLNbggCfXPk7w1HyMBmk5JAPAMsf76lW9PJ8OqjflsKPkg7juo4/
aWHPgWXYxSpp05c0qTojKizARGzjxYQhdtU4SKapgldb/AcSddn+OgI2bAo4hi+207MgD/2hCDzl
D0hAwDFLaITnzlnFGHaiiJ3BbU5eGwrm+p0MH/RyeR8k34cuNgbFW/iSravqqOhxQ9AiDBaLAHrp
SDUJiYBqkcVVuaQMuLXQJQyqJHZC9a6Dv3kLphZvVj5W6NCri8bBLlEcUkfFi+Ea1JvLs++Bh9kZ
y3nML1w3bOV/Vr1wzPsRUiNtvERzYc1VI2343MHg7AcBTgxgJSID1ooSMaeW9ZppSbbq0Koivg7e
Tet024hamA0nE5opv1BPcUCFo3XwLfeK++wcDqOjMYM0aIkaFMThJDwVALZD1atD+ZtQfdDzCqdp
EWB1tZ18RU6wLSYP604OgZ0bMpq/cMqZIZXQCAiG95eNWyFNhhpwH9lctkQ3tX7kMhx79ntq8Iv0
4M4idJ83QVeJewCcwzV7cjkei2VLMUXSi8KU6euKiq4VZeOcrX6sWB0JWWUk3hcN5s/9cIj8NwXg
5dN+K8q76xu7GeHYQKFaOTOu92rZHsrtfOnF4CteHeXqdySAPXdgzYBjGF/qhNN/FBlhpIQTJrL6
tfFBZ/aarJ1AroipAKerku3J3DWkJD36EOzq5BLl481WNssAxK1T8hxfU9ptSmT6bKIB+JyazzF6
v32bhToFXmHbMm/tMtNLjmXmLrIYw7z9E/5LitVkynyHvkwE3uMXLIgnp8GRgH0M5V66icF5VExk
K36pWELJvyYUx9WJOxusFV+k/otoaDOUY5gwIbbXVv0a5bDgXKypkj+wWNmgeQ3jKSBFSIwjacN5
baDzvm8uZd6IzI21ZkzYJ2IA3UvmPGIBtfWjhu2kf7cEkjJnm/H8HSib7JhKzeQEbEVmQuI2jVhS
FoDt/tIWxhO2Ls3KPHkYIFNBYX0+mvI9tee/Ff8Po3hh+NLp5fctq50GWEVUnTaenpxCqsf0BgMV
TSEC4kfgkw+9KO8hEoZ2EAnXzO4cap0z3pQBYYWMbJJaSbHWXgBFEqI3BMCLeCMzLSmClRyxOoD+
Fiz7FdaHP+KNxVwbtRdJsvGDEURgKWeHH63LXUbGllurdsEaGIO3Bw8vICRk8tr36cZ0KAEtpcH3
pupKq8vT3LP3qhotsc4ah4cuB2P3sejzJe9KsFs/YOWgpz5zgRs1jZ4naw6+j2j35MpJ41QYmjKH
5pdWdyzQwgDB9LHKngkcKh/Ar+kfCnTf+WvkCxK+0uv4hgVOb8C9LN7mYSPIgu6ej96eaCbCRSzg
SvGjGKt20lt5UNaLCDsnrKcmWKX4gYnyNTc63XiXbUP8YFFVazwCHR+c9NS3LjUknnYIavqb3EEQ
kO5Hq+B2pTMzSjxRjMG1frHp4/h2BTBRFMTFbkOSBJJe35UpxCWqfQFtvHhRl7LgKDMetCtvhal/
ZwewAIRtcUJh8/5JTZoWE4d+oBl3osEga2Dyt4yrpfDuCvvo71aWrYYxYNQKJPwNP5AlFv/Oo4T+
avqZbEY4gw5nmShlGp5Us+pJMEVTRJ7ne2DWK2rHm+ZUA2i3prbBrJAQmEEqPAw21K408D/4KD4H
Ox/EoX/J0tKyVwn3DFflTQ5N7WYV2ewTD1wxqDBEWPSy155HTqBHkDOMLx1qSTZBpljhMgLM8oLr
BTu/wqoRbCWyltnB4i8zybncnQDk3jZmvoQPSzvkzkG+REFaJZNYJu0e8fjl3R72Pd60AVnxbwet
Vojx7knvk3eoVtQxXee+e1Iq+JoaNxtMKmXYxARacj7iV+XcS1lq5M1NMH9XEXkG7s2ADAHFz3kv
lVXD3I+Bliu+XT8LUppkulob5ZcH6+W09P+6kN+uPQ6kdF+Awy9rfrZzOt7SjoukYY+oXu6r1fV7
aPIrhcb8qUEEM9bbPqb9ZNTW9W6uotljl+cYsLzK0wpxdTdnmcRJkyBrP0w1E4i3b/H0JULTZRaX
VrcWeEcvLLoCbiE4zKtLT/Lsz7zjnioHaaeOqAVr6oSYUPmClpTkSbApXoJAyiZHJlWC1h4rRPtv
zUVVlTO3Jcq8GjHbH5AtO+wMqSWWvtDT5HApoQ9GvJj5vRsiMpN7UX0Bx9IbGbyKAa4ZmPtGzq9Z
4t1b5h4bHpvGQO2mS7IMpKD8rI/puuJILcKiHiSfKj/vR96fpwQkggRlKlY8uQwcxjxp0nibgpQu
UyZht1PAxpIMh3fPh8p1v0aGzCa+6j6KuKOXwAnyiqgXu/fYH4YUsI0UJrQKvNG91Kxu7DLAC4jp
8KiPI6l2de9kROCHOkPmFxiq1oRuJDOWHjHRqU0QTVrU1clYUEz/Dk0QyWPVQRQJsgYU3NcCOukH
RYh7+eAmS7y2Dn1uBnfSeEJougmnoLok01GnNRvckYgA0F97eGmlfWYanBNoZsl9bzBClKdempSG
29oxTZvLWEV++CFsyFxdTkl97o48SVdXNKllOpTnv95Kp9t0LIswjSEEytAsB9n26lTodA7CW7ZV
wH2he5OeNQmpDy5ZhkpHHjcxWkmdT/SQhWLvfWP/wU0482gs1bPPxU3sKiu5mLnmsJSdyWIvoxp5
Y4kdPcxfy1Y/h4aWfhekngwF7n2PSmcgw68nXIaPKMKn6as7hyLOLKKkIfRyWjdEAYt0tVSpkkOz
9gVcceKhvku7abdzaUZW/fPUMxu1r8M/CVVQuoAHs6vTsKXlAUlbV9Z7i584QdqZJJYSqkR8enmE
X9axjycjLEF35rXFCBbxL+iqR+nZnwzCZdOtxVfpPAF6iB1b1sDO/fPnweTNfCShpGBsR9iwrtIH
Agt+amr2oL8ntdFtbSP9sB3lmNzl8wFbmrSqz4weqX87OMQb2+utDJpvFrge3ZwoFNIKqA3aZy/W
GhQV0qfy5axZl1D46JffsZXukQPPPxtwTO0gTgC+N3P4pKC96Y3uD3QkLHh7/kXYiYg3La3fw6Xt
AOqa5dbVEBXpLBR6y/BY5+d0NPftiHFP0GoIlbcRhrEjYmwIUvJ0TgkIz0iTNQva6DXEZ+uCoBec
IJ0gZhvcf3Jv9W9qK0klKlOhVRNsSU3lpUM8OwOC9qObxyidafqIl1b1A+LahiSI8ljdm44YN7BM
Hs6e+IbuMwLOnNTQQTadyzMAIU082cTAtEfcHwyX04rRoiGdPMonMSymmhfwOVwbwdJmVL/5XUOw
YokJmJd0X03Ah6er/EyUymy6mg8ceg+IbwnnTlvg74gEhxr3yjYa4RKcTPaP0b+NqqXgUc5JNUBW
uldMlIvJDNoIGW6qR6g4Z5qlx9RkzZPqK1Py8kRsANSxyYpQGUkyfLR1MvouAXqNbPMnBYh9Jsqm
S2YNfKxpv0u/ee+eq39DRh1vXMYGzuwsKEt0MJ1cz7o3EFGgnliqEimL4+WBqXm9pAXdj/QpIHH+
v4o7vl3zQg52I7OAV+cSI3ox0Vb/La3DmoV8RBHGBg5Q+d7BVFV/M7+Y55cBswzDo0C9HQG2uR3J
3cc1nklk71mU72EwQq5PM6hd3i34thiP0BnmMAuJsigk5QVsz0LaOYs87KczVUbjeOP9W2pX6AjA
G+9aIc0RZEfNWi0K9LIqmD/ndhfzmQqr+hgLSF5qBCaKA+bT9FH2HzRraBUEU3u4f6Hb19V5n9UU
WleJ5Y6FY9Tf1EBTuIdZpyKlq/p9tAOukzVGHlwwQjzs2PF3c+xoe1J090VW5/RYfGh3wVHCnjuu
T9h+xXDKqGWsTmZIHMF6ReMXPxRXzlqYSOr22xRnpoPxqnTZ6U71rjiS0c78O5IbccgHZYlGpxqB
QtC1PjgGAHa7H1lprJ+fEnLwKgt1HZENsNceYafacSzCNPToWhHSLi7WP2IKHHb3jU2GT0WrtQdb
4dQNXAptaGqmhglyfNrp/Ho95PoSc/YW97Qsrqdh6RQHTIBF6Vv9uIv2+Q230efVzOOt3iL/01wo
4t1NSlbGvr03aIV695nBxEDSvq4BxSgCEx3HFwh5sf6rXBKKK1LCljbhLCU1rS2njOQdNHRfHOOa
oZhgDuUTlzxOJwrsf8Rar1ig6Fqq5wU7ncCpxAQs1e8UoydjqOjhjc5l0hXHJA02GTIlo0MNnN+S
hZkN6JMx2wIlI6d1I51P3I0twMIJSxTb0yvjg/Ih0/NcuZ99YDmYAzOleyFTmtHbD1O7oeTLzhX/
OAlSx6fEYhsQC7csolRxXZwRnCLE4f6pih9s13Fx6eC72EapWYXoNWldge6tpbZqNTkhssnX6NXG
coMlNatwwSP81sHg9DQT6rkOFhBLCPAQZZb8LaTnxxDXWSx9A2czoNVFSiaIV9ZlKC7SOdOnv5bP
QOLzm7TeWmpS/86V94H/ckX+YSHuJKgdcyuklK9BaEUEl04UWh4RUKM9Iponp0ctGn+p1byHzYPH
o76wW7JkvN88PMvkAz88sguv8dBIpZ707OEFSYx6ShVQ7R+8/hQ6a0UtZN4gnmIxAk50KfbmiAW7
VLWiF8B9naIXYRaMXgL/Wrra6k0fm9Fdo0YYINmK8JasvFvmgMZzV5podf0hFaQlLhXccOqRI3Ep
ps1kk1H16gni6t9Sk4f0ZxSCH4URjMsuMKVrWxIkHTJeVw4vUkTZjCcZnlxxdL1nc6r2ZX2kTr9X
/AbCiZMCEaaFeel8SpugyjOyXmhWZ7O+J+r3fPj3mHR27uueHke4Cr+0NOWF71uy4OL3PEmyO+Qe
0kRE1oxA1u8bB51ftN8W1H5qd+XCkkqm1J8eD0PPWcBQfzKfdYwG2mpAvaaUdq2x/pff3+mxh42Y
MnnyZ7JELp2PEvijEWr5XBVO0RlnK5jUUlnbedYlniAjI3LexWuU17MVaDiX4SRYUWgsypMHh7uA
fN8eR1zJWhQwMhCC2RuO6D4fRtZT5eikQVi5sLx1QNTAgvxjUU+XPAdjCVxFBUxjwME/sgU9epyb
qe4E5gyq7rJSQd9LE0iZbbCKBgwrFgkwtoM9g2R24qlrKHga3njAhB0s642wXe2ge+GNMGjcolY3
7HxvydYISgnQSZsZMjmBUFVNI3Vhhc7tTTxlYYP+nAS4qB44o9JZ2Mu4pDBkQiMK6rp55Wy4b1Ko
ZrcbXwcxo7a4qaTdlsRsfzfTjqVC/BYpgJchGZ1cQZsSGoS9RCb0hDKUoNHpOPpcCqUnEYKXELzq
d+0niGg3kisArtyR5DOdyZ4CqBY7pokq2sZqtHVkzu1GU460OUpSrf2fm0xsnNyk4nIB7cOwHHSz
3OaZVmV2WBtClWHEfVzJUvKbxZ6VXrxRAv+/EluSAzZFNdcbM4Ff6uGtrmnFFpYlRO4RVxkT+2kP
ycO0QVsGhxgpLgtgOUvqM2i+s2JDH1wLgkABANHSlAvkkG+KpgFUR68FbLwYUoKdOpKSx2VvNRvG
Ufr4gx13F+WwgNyyFdSe7Yas9DX1jfNuJvz4OtSxdWFnrCKl7MxPwyxNf5D1BoDuHupOe7ocxJmr
lHYURSlhCvtyj9wcczzIpt45RqLcj18aTRTxRThP6ImVrWqmymawXFKvjKnhHjSO7eBniHj/R7IX
Uf8reewmMbfJ6XwgvfKp1DI7A97B44dlT6PzmT/Ufi19sHLe9XS5WhRqMCagZ4JQRl7VG+XSDh1Y
bNFvHqf7wUevG/+oAK//aXPLaddrzZiqN6muPnOoFdk7u8snSECpnvSIWXWOCse/CyGUcxcgP5Mu
EsrEM+noJtoBp/9jbRGjaK0d29oNzBna7h22fMP7fo7bjlGlllOX5Mrprp1kUhen7nIbJlXwYyFf
qy4plO/zSYLTXx2Bd7sI4tD03+BIl+Xg+2736YvmQECRtUCsUd9vLpCOaMMGsPoQTb/G52+6xmcf
3n54pp562LKHxqBNa0pbCY0LlMNDCtaIYZ4aTovRH74MrTKOUM6ribWelRsEsUn5T3OBnRAy/E8+
xF7E5WwSmpe/acDgX5FiRuKE/YVbMt0vxgJpVgsrE6EPzeCvICUMqwJAFCOiXvwsZ9PhoRIbFvao
i2Z/N6o2iMkfh1fcTa8CgnjL8bPxQREbTHkZaBP3no2sIhn8bah/YHHL0XoCxKmQPK52BhrqdMOL
2SaRx4QOMJqqi+EY50BNLDqOEbirUdTPYN5roAKGtBiE/pqqWPCEn+T4ddK2WrB5jye4M6eKPCjS
p+ROya9ErofpsWeHtsYqURZ8XW/hmSyZr6E7/wWvZF9TwCItWUADj2LJ7bwtGT8VDoJF5k4ZEhYa
F0+VG6MmPB2q4g6yt+dzYwr5fccSrLHqSSf6Kad73hzgVaonhNCAZNQkpWQFywrSa5UXm0Q9OcpY
fPH/2exjnqZzh6gbOB9KloRpQh3sTxX/+ONsZLxw5ErGn328q3Z/RwXHqW6mWObTPvTU9V2lY3uS
44c63ASoQ5r5mFnTORGjDnh4ajF16abNv4ZF/a+nbZpHM/wSffhY04JKqVnJA0/LSTMudBA0hoia
/onDlKGKquNQhkaZKWa2BhSXLpn2mfuQuP2Auqu+aKapMMw++gSjhy3Os/evaXSdfoZWyVH7DerU
w4LPZbaxmrchQ+dmlvGXc8qvZ57pvAaQ8Bf5du7Y3yORRyFMYiAUlszUOtjmBBstpRxZrdC5/L0Z
6EKzGR1PsR+vCIRM2G5QQXSplk1gOv+Iwz3ttiP9RRiwqrI/NJleHQRsjuw+ycGTXktqomN2P9lO
LvhupgRZ9MILeprFxdBTtF4YkyuYAuUwtbnBja+DTX6ul8TfbB1nvLTWR2V8LzmWHYla3mENEVny
wx647ibyGFljFaNl2FYf9FHdlpJ70cg+/wTd6o+NQlg6ZqJmWEGrFKNgsg4Oe+3/R/LBJ8xZ0cVc
CcZEOQfSHYSqn7GhDunnd2w5dmoiOfmlW00zhAwriRH/dPEkiAIcSXq9gbig/0vDSjRFxH25MHqR
GYRXhS1HgDNbud5vSuFCORtdsSaA83AK80ZkmKSoCkLl5z9Udu0WdlZfs6y3KEMCjnq4BjpvVSuZ
Vx5u16MQfqZiiMr617ao3CnQ8YFSs0YA4Qo+9iEDyrSJJ3vEg6SReCzS/RI8Fvv1G+9iSb/0nL8Y
maITqo0f1PnhMkMehiUzdly4AOcTn7tHYua/9C/7/pe0s36Dt0woEgv0PcXljk9VaHJpw8d3ixbs
xcGeuLL1inC0a5wMjJ/cKN+TKKmJAc8DkC0V8XhJs1rOBvBF/7Uebz/GYBJk
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IWy3YWsFdnYW3quA8tFmWWyxEpCeCXnbQkML4GIWmfvbHZFk+1+569Zzen+0g5o8pnGxrYSJzdeI
4JT2sC7eIDw7Xdn0mFQ7/MQSdVxabUPw+JFb5+yaTF0J97YnoGwc1Elekbi+w2GsQWO9RDOvlcX9
VzlT2BAxvdc7kJall/+SgCHjxUugB4g/oH2O8IqIrNYztLkFW6XWVhKm3ud+TrGKnZ+Hg+kc/Xrb
H2r/l57u0vJ5gje5KS3ZpmZ+6rqEIVuS0cSan7oSFO7zhTHXLoZwfjD4U7BHd1Imi8DH+LuFMA5k
+c7srkRdlz34/Mjx4a/6s/xoU9nqaQyKF+5ITg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5296)
`protect data_block
On/m3SqXyHrmM1b0Y4IZizL1aHUXGdUY7j++MeG41qhwpjHmMaNGCKkEXIS9nWJLJF9GzOaFrGOk
0HiQGlp2AuKIUWEVJAj95514Yf4CpG14zBQ6InPj2cuv4vM0L2bNkQIvN1tQ6bvDgMCx6+TjjV0M
QWdCvYuJUfwfKSVMzsKfsAcBk2iwo5qlnhwshGeAK0hFfqmHSENjAc3wG4q/Raq5caQrCkFeKR+5
uBuxg7ddfE5J4ABDKdN+xCo4PFHQIZkcIVw8+9X777kc25X1O9qr1+sT/gCGdhTeRuA6qIRAiwPt
hboEHzoVi9EoOSwBdHGxhlx1+IyTJqaoloN5VdvFF/JK60tbCU4xC9Fx7dm+B3uBHGh0vZSbL9/E
bx4CLsbReMwaaH9xpmK/98yf8wvdOP7Kmb8XfDHBP8KCFWtdQklgC5yDZHpPyb/uhslJ4aXTmgw6
mk2D9cq25smqn9baBSreeFPtKhoD7BT1kAmCGLW9bR4b8LkDKXA/C6nEnuYXJen1x48hb6djQKcJ
QqnSnVoAHb9h6bXfa0oulJoyKlXhTlzI3uRebdFjObnRH2M17O9b9N8Wo1rn+CaOd/ptqEft5P12
ei+Ns8g/5By20vuHxEgwd+5exTyWwEUFkHeiOSXXJ5VhlOcE/eE4g87UPHbN45nghgA/ipXtRbKR
318DvVnj2MxZxaeRMddCzl/Nu/SLzibApjgthDMFhtKXMwRJCzUjBTCphQGCQgjQxL/JRH4dyPPd
xOWbzVxpGAo0Q1j5TjKbYMSYwLPZE17MSk8z1JnYdPELM11kzglCBevQqsvqRRBqN/f4XG1Pt6VP
xHJmoEKBLqAHez4KsYKwnv4nniX+S8kBezOHTBnA7FXC3V6YI6IFTLiHL7a8e94Z9lMCnJDoxBhk
QCvUcy4hXj+TDUT/PTmKzIRUQi2Wb06EBZmLOwrvPq9KG7WC/9gzj5Wls3rO3Vdc/Xda7aCqhiLm
0ZzGp01UoEXa7fYdCH0vbxr1easryPr/iydNPnNG2fFzzND3P6hia2evbk6/hEuFuOhFDAPcwNWJ
cYZmYPuNLsooxbeCTs2V2+8xw/Ihn9YlUPh8NN57UI1yrkww+RbNe0jNDY+XFACSjoKydl/+3RhZ
7r52c5qlPp1PdDhFD8rpxGZpW6YyswevFp9jU1s5b2NC0SYeigVHmZrjkMviWIavNWTAUH8fxgHL
w1b8TOb37Y7AH36CT1uMSLgYH3iSysrwfrDFje9KatB4Vx1i3lBctZcytHuD/1lMWWinFVUeH4XN
JgF17ZrgvylrXDK3kivxwwAKNmUsuOydYWXoqWlQCQw6VK8jd8npfxvTxH0rG5kvOHHtiqzn0lJQ
AsqqLJRFnvtWw/5CEpFlTj1zY26BllOWOQECEqbt5GlYs2kNDUmWNI5frmpXZckGk+pOjHBKcBIT
dUOkBQ94dBLvcqPYoZmdym9yJUsdT/PIsOvcoJ+oP62STG66qGCCSOP+atWMY0TMzIO5Ttg0Y2Nk
TN8IjddkrTaJImTNn2m2kgkhwyFnapvmTI3U8YKtK4cAwtoJgkWnAOpkSgQGfh699pfcYnEmgFRO
yhZ8JiVbgK6xj5Pqyyn68NOVVlzgTqfC4pyNvlwu1e5I2EnNUYdTntfX/gjJRPHWS7P3WgPfk4+d
gxNUb4vM6edIXg7iw+1h8CeJM2mJONLs9H5yWwrfHYN0eoP85Jc+mmM51W7lbjzkBI1/g8xrhUby
uXctI4dIRQb9jNatEB4wFzRPZpxYsjGJudU2brgU7A9QayfuB1LJkYkvOcEWw7xmJpCUjWflCuMR
I+UI5APsXGgwqCsYf166m2ZpWZS/wkrYmZbdNz5hNmRi+7iZHhJ4T0Ii4c/VTdbZ3qCzyJZhuBOe
Js/3tmywVmZMx/dCfhX4IJi3WlOCcScbeY0qL42uNIKJ6l1yZw7NFC2Wc1XNBSBaSQV4S6+nnakl
Ix177+2NpQ+6y/zS6S7/V/mz3HNETez1+s191D4cbPH74hIHmsymY1ZMYWWrc4l6PvOZ2g4/aHgO
X5dvOugi2asVuX4D4QJA4W8L/scr7hMhPMyEB+PJZ7oriymD05Dt6yZ9SNOyRT/R4M+2OZ6kjrnG
J8WUbuQLsY5daow2HzvA9gwoZscvItR672gIDIAwZ9r5J/0gwLydiGvBvN7e1XZWuqRDenCPu3DI
7ziD3eJHKiqsjqO+B6tKxtBr7vFiF6etyFUQTWgrnX0+CNjk0zqxfQXTNPErIbmbjHhKSyHNANRL
Hh5M4Wpv3mOINn4fztfH9AXV2YZpW6RTCCxGnGU7ia9jvRQh9KPqGeSA1ixhV38opJyDY97INfP4
pCg10YweWapL3+dNt6fEnExp0GFH81A06DSuNYLH3YeEc7teKxVwsH2eXWc1DEuXbay0k0kaetKC
VKAHSF4RwKg2yB32ya3SQlB9slgl5O/5cgfjrwikFI4EgHHnogt5YBHo3/ZwJI3g+b4dlzs+CKre
lKHFH2230N18JOfIEIPjzV1qrNxYGntDwF99XOLn0XEYedQB8Fj4hjxso7DtzkEqU9Fq+p66g1D2
ecsU9D/prqpnru2uMuAlE/vEijsgH36BiGX1I9zBBBI9mZdXSODrtNUK3PQZ05+/i+2HwFLmGEtA
ljAd1IOiLuAeNEnqTO2m+nVn8y3c3+Pl1Sa6kPpTo85aiNooSCvpK6xFg+bz7/IUiH/5Fb2tw6qv
Xe+bN2qy+PxJ/qJqhgNxvjAUHZ1JJ4en27AlbqTLtwkfRIs7piexnykRmUe66TaTgZP01/xiJqJ6
YVZKaDZIeBLJHlgKzArMezDmiBciLpyNv/e6urABaZkb3bzMm4gpoBVMnWmgcRRn94jcawOEP1OZ
M6rJ7xADMtaoSViNVsaVNEsjaGKYU6nj6xlP94k7zZRM8wkOCenHPuGLYCxrNOxl3+je+ra+Rg/y
vTZGpdA1AbS+Rs2INc1Bk7sjVxQDYpaQEyHlVVMRpqfCATwW+GOO7EPQ03hAzbjF8r6wW2OjrWcO
IZjdI64U04HcHND6q70Ez4tceMBTgXwqw1FS0jIEr4+iMer+5zn/tfwSQjHk8e8JOjW/RJW2oNxx
FOb8xHfYE1wV7++Nt4Sr6EfJp79mdtntVTqEAgKw7iMMJmD7l+qAApxCdGwjPY5t2UTcaMtegdvV
DNKVTtfrDQuBKs+sZuJ+ZIJQVAoJtYyn+LEKwJL80++nIf8hPJ5bAmO1s1TagCC5LH0DT+tC8Qml
ib7fIcNc5tJwUQZrnY1BxZhEWz7qrsUSHpCgMS027X2T2BUSy9ZoNxXmAhoZxHS2FRFDsMAyHrAp
QXBZlo/qugHLpRr9QpoJXyMBSsKG4Xf+njwUo1xqkTQ6JO3hCe3P7i7YZyXzZ652K/X4v2+GcptR
uIdpdImceqSc3SRZCdO0lcJKeFRax9Zs8ODWNl8qPBm/7XRVYUt1pvVA5+LSIA3DaBpSVFmpzrKs
+M3h8k2WZIHYL6tT4mHz4jy3eSNFvMknpxZAjC2FxOpzxA684aJBgwwGXZ4u/EXbFTd92AWbgoga
OnnqMsStyhHRAwq53IPXJoMgmSF2bbLKdqqbIvD1OQWFc8Xf6O2hzlgQ9PSz4Ybf5s4Ru5n2B1cA
1fzrcVjXeiw8gL2pN+HA0dWo8IlInQWzyLOJ8Gmlbo6vL3u+r+eTPLJPT8A0BBTyEWkxcAgoVz9Q
ulM99d+4rdqhfrtQTFyJ7pfk5QeVu1x/0epTh9WKhNJYJ9hI5EmVWrmOkzn/7lFPkSDhxE6xa8yV
9EdY/r3v125Rj2p9emlTLFneC1Rb1rTKnBlY2bU4Gu1fBv1XbdQ12PHafMuDkMJjRlAHLCTXvz0p
duFyrjLQ+6uQ5e0POEJCU4rUh1ingnhAlYkR/uzG2DYOUXEavOVmlm9WwBA3wfnG1RlySwUCffbT
mtZUwkeiPDi1ZBfuXYeb7Ekd2cIkGj5PMmWFUb7CztSYu15P2lNZ71U6A4kK483VQKH7687Lw4/5
TMQmndfUjiAwXuJHnOGJC1rxMYKyl/fdf58XdrlJYUXDCToyipMfmQj2rIGa9qiqbL0K/Js92Ty+
+DPEBuv1XthjfeAn06F42+LzoycMhOnuUzMgy1SzCZZfzZ5/J+fNPdJuYHQQ/cVgkuIatp1+nujD
z5OkVMgrKuOZrQvXjbq1ex3IhidXwpf6tmiOSL/ZlAeLXyNr44hW5PJ8T2T6WEWS01eYo4fslL6K
FcrRkqrCJu9sOVkaJX2RyxE+54ab6oxd6iXM79zWoa0/R7QzQvn4mr4GV3KLBeLQgCU2L1DqXWjb
VVVxmBKyJtUFaB7t7DjQtPn+wlYlvizK1E1bPl0MtvjiW4nsoVnCKxsgz1wEg7kcAUXMFB72IVMp
vgVDXnYQaID9ip3UWQrYoJZgtMPkwVpo27qanUmN2xRSFZHDiiiZjWNTOJv2tkc7ykIu4BU8t4vX
NfNm1djd7pa2dT4BwfGiuNSTq1G743O8uaxFTl+iJzRnq7bHcbmqmKXi888k7w3H3V0rbEOEIg08
+ZiQeRemnOWHYt9SkvGEk/xxvpYnciDuI8vqFDlfCQ9f798aKmNThsXLkktFM3/yhZMkHKan1x2y
6xVbv8eCuaCi31iMebbpJCjG0R1G9oZ1U0hnBSRjXfSAF5dd4v/aewZOEqkthPKNupv1QDH4Vw3c
UxrJtSK1QsLbDKGnf2P1ra8F9rg2hZ0YE3Sro9UFdVNv/qhg++OIJyewiRqVsJCpB4QMKIU33Bow
/3j9sHcsKlwl38/9rYkhlRxiiRkp2kfAInB5WwvpPCuVYRTDSN29BdyrAHtx6o0oOvkeBJvZ6JKA
RhnL307/HaPVcDcbmO45Mi3QZo/D529ktS7c2uYOITShM6TKux+B07Zsf8PAOrG/3OszO7oqZh4r
xm/fTt7YCi3bD7gnZrSqeeaM9oXX3SZxZuRzWGBi8qmmf0y2T2tpiU5Ew0WipP+cG4KlTXSejmpY
s00AjmOCf8z81W7WFsoRRGy6UDzAiKixpHNgdcd8uACPgCclh1SRAoh9o9UBR+PrLCfjdXhjcZUo
Oro7GRgWShVWaIQOU2i/XdU2kNTUD5iUKL54yj5ZaQruv+NZs7HCcfA8D9Jih6dvH8Rp7hy7pshJ
k+5c10Aol02VvPt6Mmdo0+zPlwdsqbOPFJQryfU8XgneFyRRLAg+18ty8OCQPZEoW1i/F3QvtAvu
Ihw1fBaANZAWo5inACsURJgpS8w5Xpas0/JGp9fJ7hXR763c5XSQOQRXM8+QqK3JrPTD1juS18Lb
tqC+WZv65V1q8AibRXCCn1CqWimb9ogMzdBzHv5zmJmGvl9m0okX9S7YheiCXhl7h+qp8Mwedfkl
aQSMcauwq7x/UxMIXY5MUuGbgC6HSd65fLXTAy75PIzo2EmfzKFUTe4uV7uyxeuKHVNrmwenVdnu
vLctQBcMTxmIUj265g/PBZ57YnfVFi7A91j9ehq9Wf++tL+cHpaOtbldtF0mfQLnyw6+6my362JH
wpz4Ut8JZVTj3KUFGKx+jbF6iYBiw2nNKeTqlM8yhT4k6EYpW0WgO0L9LYUsHYzmD8we1xGF/Gg6
QLEVyafpPGK3RyWRSTeV0cBAMWhdvZv5/G6NzbyDTogOEMG2umtQAUNwGN+8tsuhWIqJNzG3cPD2
/BbH0Pe0+4Itl51y+HJFNpd+LLdCSUvTqX/VuJwAsJCFxjArO+SBFAQfU6gSTkKOCIlmIFiFnqab
WtUYVAXiE6QZwriCQgh/CojA5kukHqVER6DRFrHvB4mY4fzqcq2KchZfaO24vhoj5I9GyIsh/lHM
gj2YYBznanCXiwmGn+dJqJo6yyNmhjPOnKjoS91TEbtAWZX5+aLDxS1G9BxsBK8Bsx5HGa3ttqy8
vmefipTyUdjg670vuNR6FyNbiJBGrA6H2htKRhAlxV6zvZ0GqJ/IxQlAnn0Nor/l6ui1/A4xtYBC
eR/d+L49pVX5JaZqbnELdWfs8TFGn0wjGdUpRcNGj+9vqib8kAQ51WGPJQFCDSL8jm5j0ojqBppS
j8gUx6fj2vyi9V3t66a/+u/VlE6Bx0RB0KIEsdWE1L7qwTsdlemc6bMWG38QDpwlgwPjRTNuB33w
ddzLa3uBSOVRJZ2vI4ZoXKtmLrpNweMiotOSsz6o/3Hwg2srBHstpuIRCQ15QKAt0CXCpUqwOE/f
w4BYTZ/+hlw2n+pFWA0Pt7YnCOQeBSrXo3mGJHSLp4FRML6Ki3zA/TQJJICMvazUgSpwebhJMzAx
F7WZF3drhFK2IEyD3EhDBMLvQ3d8tQddxRbk17ajPiZU8raBHFj3NzAauIQZ/GywP4wRoiVX9HX8
LSe66r0s9IPgxj1JZbX3JH4HAe4Nm1MkbUn+NLf89wccvKGIngbIF3lRWrKZq2wL0qM86xZuZh5b
0hQlKESEhUrx3iFyS2vpJNh/eQiEyMO8zNrmakMiWapRiBuOTRbvxsFSpUJopjjSre5S9POAbIZM
txnyEqK9tNWfCNSeQiocV7jJji5E3sfNW1L857ECOX7Z6rfjuB2i/gL/63NgCPGanC5IvguVmQeM
wc4rRwocPSiMzPHdaradfde5+u6zRwOjq8jGljZbmJN9sAPoXccAxG3/TzV8qmoj2sIUiqWIWubQ
SKuCdPTmvWDMR8bj2FN9yxMmdw7+Z+KSdsUH+gQNb0GTX8VNmR8AKtfn84yZa+frSeusN68nhols
hA+ZW/oCWxJFDjrEYFHFxRxcRx4gxh/QWfcAUSbfgZNTlf5/Ay8AM3Btrqb9Ln5JMgeRUr6EnnE5
4S27uhdAIahH5r70ONimuHY3yx2HMN/dWTm8KDUKI9VIdgj2Vg4pbFDvZZdIbBVuMO9sKtiHb2Wo
hE/xzQJqCjix0pV4dPt1l6s08vbNy/DrkIvwpi+boh7jCmoaxRs5E5BUx3vJtGRyWD7M+5shCJKe
TCVY7CLQ0hDqWqz8WfLvHqeo2WD2wQ9d/bEsxzus1L7tFS+8bc3HlYOfJr9y8YHACIT3RA==
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Yj{�?�Np����wf��@pl��}B�(1jVe��S�I��f�yZT�����J7U3�?���y��Z�xPӎs��y�uB�]�ۍ�MO��N�IZ`Ú��k���8))����>{2O{��ǃ�g;��q0�U[5�7|
<�ДL<����=�dC(���qd"�덦s������ ����7
��|J(�
���XL��ep���!�+޽��BBBpɒu����1
�*C2]"�(\���ğFIj9�@×iO�l�����ȸ\�(U]�/<G~��>гq���LSz4^�4@ﬂ� ;�ל2��a.FoV�%K�g\�0�&�#�i���6�q�.����4�� 6-^ �o`L�R���p��Z�_�ZI�a*uH�j,ET����7����AZ�~-B{0Z9�w�J�83�JS<]�F&|�`�y��w�aO��x�Д�����Cv�x��RO4��6qp��l�9G�2W�{0~�ߢ��_�j����3r;+��ʴϏ�?�V5���q���F�)��A�s��Q�=�_𾊓r�̔L? 1
�\`œ��v%9(k���^_Y�7� UTЊ��7�8{�F� �B�DC�	 "�R�CtŅ� �k����pXB2�ޔ���\tv�S�T�H����Iϝ!1�p�)E���W<5+��$!Co�ʡf�K#��u�I�<3���:��ڴg���ޑ'F����I~�(3 �%�=�����;sl�Y9��,U�EyC//�t*b���'��ڽ�n��GFuQmR�-���?�^W�R+囿B�'Ĭ6��ڞ�������Z���"x.(B�'R�)�bu�ˇ�cX�S���z���9��䰒�ˮ7{I�þ�FDx<f=�39t$G���r�`��1�/�\�լƍ����O�?�JԨ�q�"�!�O3��)Ub��9�V��� ��ͼ�	��.D�l���-)��Ĺ�GKZK��a��׆j\�MM�R��8�AjN��1b��@
8��N���޾pwit��
����$M�k,����p-�+L7rqF�2���<])��k{�F�<Ȁ��Y�0U�C��.���_q�_���٘�)�?��B������2UuG��O�J1c�kB���mf�u�����M���"�j��'�W�����M��,��g���0̃�ڳ���S����]ǩ�3a�}���+��=�;a`r*�`�Lr����a�K/q#	�8K�?y�S�<`���5�)`x%��X����Rdt�6�p>�I����	0�:�m�H��\�Ҝ�gL�e�M�"ʚ�l�v4v���!//B��������Ŷ�O��q��RW�ɂPtC2���9���b�����=K�Ϝ��1�C�w��8���`�,c��p4.�HA���W~�	&������<���c��`���GeD�uC߂�fIlJ쬭 �"�S6��8ƈ�9&7E=	Ƌ��O�Wn
��D/�ݒ�猄>��p���v�V[1����F��g��C�QgPPc�Y�ۅ��F~"��`+��JG�����`:Dm�e?Y"��Mf��C�&~"�K�,���@�hH�6WI����Lp@e
ҬO�p�	��e9a�ؘj�������K��9۝dS��ƾz� ��EU�"��C�0�〻eN�nڧ^�(�V�lV-�y<��_ɭ{Ls>u�n��:!�D �!TOL[5��kY�q����i��
��ל�<s��vy]�F�5v,ҫ���x�h#K<QDg����X3iWH�Q���EXI÷���tk�s�\�<Ǻ�UR`$O��#r��zMLO+M�e���\��+�:R3��3��\�Q'i��"���x���Qu�&�.U�}��m���f�ׅ�쿙zϳk���E��~�� �_oH���̤�	dG��H��(>��s��
hʁ�y�,��wXp}��Ҭ��Z�]FiJU�{�ve|b';���#E8v�S����H�[�tj?�F�`;p�8�Ri}� 1�Ԝq�'r~r�\|�v�i�CX~|�� ��+��K��do��]�r��o�@���DwS4��U�u8Z�A	ߐ��4�4�3A������}8m�n�/ӯe�
ގ].{�OȊI-n�4G���SÐ�G�䕖*C��H��f\��/�R��L�p����o��r�����DT�q3�|��zkqr����]~��=�wT�i��e��AD����<�g=O@��i#���3G�Pv�+f:�R���$��0{�8���I�
}	��v��F/�A��nb����Px�rf�b�y����%$hS�S�sd��՘^o��=z���9�v*���k�� �j��!�y&��8>!͘��D����T��p�?3��p�h�N�H���6�9�tq �>� O�]��L���	޾��+O�m
�����1!u}�}s$w��H��	w��������E���0��8��T�<6h�CMf��DM�$����EB��IKзHH�p+�����^����ܙ��2@ "O�4'�z+s5O���8�t��?fm�`�]U�><�%���̂L=k(
�y�I�_Ö|�^R;�y2}7����k�	���Ȇm��6�Rw��Ҥ�:���:��� /vq�h��h� ��x�~���E+OC[b��pL9�R�����XT{Pp/d�0rT�W)�AZS��E��>+2�ﵠ�-�e�KR��4!ᑄr��d��Tu
�Cm�;̼��ST�h�T����oBVĢu"���,A:�_ih�8M�E;�1i}\��	�~cQ��gi�I�g��N��J3�B��Z�8OR�'৔�R�QC�;3��A���Φ�̨N�wӇ�������mT���]���ň]�3񓪇�'$�.��.i���=n�<;�G6��{W:E'�����&z�:��A1�K/�d��=��ț?�`�!r�4��`��p�<���y:0� -�N\�X��6BHnk�]F9��`Χ����ѿ=n �J���� �<�{mr` �����m'�"pT�g���}�gy�9~�f�Q���������bj����ńԂ�gy{3'�<;�uO��j%��ӵ��?-��z���?�X�,��%���m�t1`	a�ʗ�����o>��-)�㩣���K�\6�G��m��I�H���	���h��п�I��m��QV�$��8zAǔ'<�}��NH���If��Mrp���"��V<0��-�k����9�븮mؔL6S���[��d��uӑC��⬧�E9�?l�e�J��_n�{���ef�7}s-�,WB�6|ߜ�`a���w�cM�@k��t��}�{>)!��R���;��+�נ�Cm���*�hcB�0Z� �f�_�:���`�����H���`"�9$�uU5���n"���ڳS�C��1͓�F_�u��[�U�ASO�Mq�[W%�ňҧ�:'Sp��/4P�����	hǟK�����8l"���__IE8�Wj/��fG�`�c��	>�:��K
��F�Erʃ�`9!��I;W��pW�{��R�5{I����B�?	�3z�+0����d���"�P;���K�`��Hcq��,����V$�M�;)����l"��� ����v���e �]��U0fZW��Q���\~��!up��b"U�k��#n��p��Qv(Ķc�֧��j�e}ྸċq
W�.��r���
��?/���뉑���z���̭vbs�
�����X�B��ձ�.8�|��R?�/���Zoq�6.,��+)��~
�Sg��泘��a�C�V!Dp��!�
]��;����=Ee'�X�3o+���ʈ`��&.���A>���({J��;�,��./�/ ]��ş5�?����EqBD
-�,aB� �B���y �+m�B&L�0<��ck(H	���e
���*1��P��*ȊU�8�$i����� v��11<�P���U�q���"M��<���{�P�Ϥ/ڰǋ���w/�S��(�
5�)'���m-�YU<Ҥ�+�j��L�9T�v�c<9g���nvi�w1��@�Gk4��E�O����������RJ�1ʗ���em��g�)�Rf����J+غ�7��N��S�n�Za�yiS� �r�;��,��96\!�P����X���]��Ƈ)Vo�̱_�i��.B3 �/�W�"����{�|��X�и�nۤ;!m�42)���݆'P�A��{ ��m�a;I0�۴
�|sK�rZ��Y�L-f&H��w�d"��c6�%o/ǅ,�,d\,y���R���%`"���2�?���������I�/�L���g�5�[�����.�w�<�<���ƶ�,`�A�њ$B�1/�A9��X�����"��j�J1؝�8������-�$,�����eNT�%QQsN��Vy���l��z�r�F��@v�7ǠG3��Ί���[���z����> 5�����&�s�iW�*�	�U��P�%k�	b�|y	>p�V&U�i�Yۥ<@l }~8��/7����FCV����;�<�%b$$�7*�Wv�|�����ټ�#�/+�[�s���-'Y̥��F\Y��Q�ļ�1F+��~���{�4�뜼���}������w�	/��`���=h��ɭ�3���A5{���ٟ䡂J�"O�ru0i`"���	���_����&�\��z�Ӿ��	P�a�� �ԊB�X}�gpOG	��7�<ޗ~͙��w�X��#߭x(�#�y5ǳڳQfNq3��[K3��^"���y�2?�5>�KJ�������!@눃�@��|W`�2b8��8�P�Iy���8��xg���z �Z ~�E�m�t�[�"��X�/�i��F�ʶY�����'��l��󰎸��ϲme[�&����BfH)Sۊ(��	/ߊf���"ԏ���{L����x�0���߅�ޯζF)���#��=Mdu��t_��.�s����MoP��$h���x�U ���э��q8xY�=#�̂ [Zkrѿh`�YZ���F(��a[?2�����@v�
�x�5� r� �|�]	��!#��P�ThQ�$�:J��x�n�VA	����Dzi7_��� ��ܛ U� O�r�v���.H�."��;�� ,~��۱�7�H�s'	����O�2LO�1�JFn<�RmtB �Q��[Q3o�DtpDq�d-�gv���o�T~Հ��<��A�z�%����Q�w�L��>�k4�N�on?�{H�]� �����uC�%�h#fµ���� bc��-G���N�?Z���
?��@�Þ�p�S<��c*�1vP�8����D�7I��I4�����RnB-B�{;�C���0k��
v�[gGVEU���"O[��L�oKG�膻1|ru�+1�����NS����%.�x�p��E���zm��D�9�[a'����������#w88�A���ZK%�1p�.jR�,fΠ�s����V��'��U��?��$�W�d��B�|�D�|:�*�C�CF2�*w��ʻv�(��TސX�<Q��}�sS�<�U@4�%����1S+����U��6��	fD�����-��栠��;�+	�#su�'�Cxʏ��bk#�<��h/������qn8������S���Vl)г��4+
آjK}ϼ`��Q�Gތ>�W�X��K�^B�Ζ�u�0
�{w1,r��^d,/�`r�k���p�_�h0�36������,C>1��\��D�����/�դ�K���%��H���c�EЮ�:������[J���ަQ��)-q�lE�_2���,��ظ~i�|����/��6�����"Bj�D�W ��#$�`���E6'/�S�U�W'�� �/�~�=DH�V�x�����ݼ ��A=&��ZN�/I9�FĞ=�`h�'�<9�=~���{�|榯h�=��L
��$4�}&�_`\>�/�I	��!x��1��WH��5L�s��H�g����o�J��V^JM�*��lv�ߞ�a0dA��*Fw���lǔj�P2y(����aѼ�+-�eEŁ�0��#��;����wo0�Hh�Z�K�8����3v���8N���34�%�^�-��0~�8f'd�%�������'4 "P�Q�!�+��+�p^���Ė�ؓ=�.�S(��&<����^�(^c羱r��1I�6:��Pf
�9-�eO���0�|��oa!! �%�<�d ��!�@�J��2hD h�a�Y��D֗�}�}�#Y�h=R�U��T0<�Ӎ�1��O�K奘]���hn=)�50���dW�D��X���:������B�T�g�;oq���'#��a�J��)��X�����bS�2��IX"�����G�t�o�8]���/1�A��9�����z��Tg����[RS��&�	�"2���J�J]��K]�3�U�3����-ȥ�t����U".҈�_��e�˥�s(�t�嗊�%�H���PV�l�U)W�7�a6u-,Hp���RM��8$��æ�Q7�T�V}e@4�ǚ��:^�R�yÐU�	�;����zP}��vt�X������+��{+;@W���g?�|�wkrк�!ِ4��;��3������4��L@�:s0n"*뽞r���W�x6��	%���Bvv���>� �Ԡ̃-�>^Qv�U8գ����1�Ə������r�y�i�U��rƾ�� ܩ��u�=t��>.�D�����}��ևl�
7�n��݁"@�.����hh>��*!J)�х_~���hg9^MP2�KIe�TmW�B��B�yBJZ�ȋ�tK4�	\��&\�]��V;���j�b�9�ښ�9�0����hk�ju���F��U�+���vj�Q26�Γ��Xܝ1�h�y��r���ٷ1е̉�g����b'���u_�\�����r��^�8H�	0������
ng,�~/;��TfLq���D��_�?�e\I���$�ߪJ;~W�?�s�6��WJh���sM�+'�a豾�A�z^���6��r
��zkw��pE&����{��������0c)��t
����l`�A��Q5�(n!s�>�鏎p͘됔d��F��E^jc �jl�#@g�H��j8q�Tv��WuZb�q��~���N�|Ai�/{�t�K��a��]l-�B�����J����d�/�iɶ��;X�ƭ��qz|H%�7����S|`O�9��'Z�u���)a���M�Τ��N���L�;����C��yM_s+�5Y�Wpq�����1Z��Q'H�i�r1�C3�5|�v�ϦD�{lH)�9��S]��q�OS/p$|R�af��Ӵk|�9O�\���
}B9��>��{c��Y�@�PZ^�s�[:'����s�G�.�(�&�<�����|d�v�L�.K��-2��V��@��z�Fw�aipĳ<x���&�&�e�a2KtQ`���Ґ��m/�)W/���Ͻ,�"⩮�:���X�/Tz}|��6會3X�V��,�U%���v�$=Ig�֟�
�-H̨3������օ��AeF���KQ�R�{�������/����3,r�b����W�k~�[=�3��G���q7Xt�=P�	�ʖ�4wA߰��jJL�n�5!�cH���G���w3@������2����>�����p�F��.������H��Ė���	��_�)KhTZI<>Ll��	k�z��)�#-I	&�ˣ�{�G���>gB�QK���Y���s����\��~d_#ʌ���S�+k�xr�T�,�槨��BppL��ad�aq��-mZ������A(�R��e�Z�K�!�G�}�\�"Q4����,"��e�JI�^��V� l��\�(��4�F�7������27q��\�2����"���G���?�z�!!���Q�Tk]�u& ^9�gz/>_�'o��%T�0����E�k�vg�A>�:���0+�|*TS�Gme��L$m<�)� ��TT~�wz�6C�� �T�$��iR�bE~.������Aϲ ��am/���zD�۠(
D�����hN]N�|$��M5y.��db�C��Ӕ �`Q�~3��>�d� �3����&��Q.����ɴ�7����MML�z@���	(���,�X�5Nq~nXM��ud@X
$��`��&�ƿa���R�z�;˕�A�n�o ��2�>tX3O��2-g�
�6*G��_�\`��V���������%E��0���L-�m���\��-\��SK.���a${�%V�ch⪓9c�+�T�nZ�����Qųc����Z�m��\�T~��|\��ukU,���XȖ,zQx��NH�ڌJ�C��<Xx)�2�͝�0�q���X���H��as��y�������b��8VE�Y.��E��SL%�`:��6��p´�)�e��)ɹ��K���5�¼��.�l,q"��tޞD�� ���9(�1� �� ����� p����q���	8P7���[T�W.x�e���>�����k[�$�#�Y)�C�����v��?��� ��h}�xwUɶuwa3��,n�&�x���_�?^@��f!Ȝfչ${�gru^��(�G�E�K��&qĽ);~�z�$Q��0Èm�B��,�h�
\J�sJ�T�պ��I����C�wZ*�?��c���ށ�煕�����M����߂���L���̑b�ū��C�f*�	��R*��H��*f�_���P�s�z*�z$H���� #S�NZE}84.C~����U�Zp�aqr��k�D�~��A>R.��p�G]=�TL֫a�	�6�/X	U��I���eD��Ez�(1@0X��q/������.��QC�d��z1΅,�J���9�R�UPV^|��\�*��3�[�u��W��C�0,�OP۽���7��bT\BP ����^�)x5���/"#�ŀ���H?��p�*���u J5V!Ϗ?p��nB�Q�im'N�D�Z�^�̓M��;/u�[�Z��D�X�qR��K�m��1�1�z#�[X.�<S�	�sY�1�6'j�'�:=&x���T	x� ipW�������J��Uy�
""2�߮�ګȘ�3Q��<#<%�nI;��3�u�[�}��b���F�=K��ظ�f�Ͼc����kl���K�͎�a)�;$2=��~1�Z�i]��M`PD�VLs��U�He�<[ հ��^�|�7�K|��gЙ> �y	�����<�f�S�m:Y�1v'�*a0B���B��w穉�yڷ|Kw��%D6�ݔ�Cy�5\7���?wE.5Sm������"��R��5;�ﺻ`��/�P�s�M%`�]@O��'�$��@lo��"�t�6� O��uT4�	���{�x�Μ9`6�4
DĆ!��֠�96�^[EV�1sz�}�{W�(�F>��R���*�K���~�mQh���jL�'�� ��7�����:�Uοw{��`4a���fW�����	�Dn`x!�ۻ��t�`�Nސ��b�2\/.<�|�a�k��5<g
ȟ�mM�J#�(m����+���H��Tg���0�Exi�Y�ҏ�@�k�6{*"fp��p`zꮡI��A5��d'Q*��U��Ů�sD(�y�*����dN�L��0��q:;��et{��m���Y����S�N~o�_��+x	}:��l�����P,�� �5���դ�76������͡ ��k�AE�wC�eȈ�i@���yx�� ��)P�1��x�0l���H�5�Ԝ@�1���X#\K�k��AA��59���A!�Z���K��1NڭkA��9S�&��d+�(B��,�e�ثI�2�p Y�\`�ƜN��u2���3ڠ)j&:�=��6�-�voƪ��ar�&�Hqf��LW\.5x�z �������\���5�j�&���t������r��ݘ���'�t�{P��*�hg����H��aV�$nG+�B�X�O��{'�a����������������������?A�� ��L�df��:�xSA������r��֎)z��S#�v��.�1�Zi(�}�L�A�K�a��*ƿ��,Y�s����w�{K����?@�kp�wYh���e���:|�h*�e��&���p	�X0�@p��p�/��R�+�]�� Z�T��i����ݨ���Y�yh��s�I�&CB8w,82~������+j$ዴ��Χ����K;ͦ3�e`�E�]V��RF�e�(�'����|GV�R����'/�u����Hrn�U�!l(����"����)��,2Ս��z�*�����(�5��4A���Ӑ"�.;�Z�WҒ�.�M�#�$!�,@��Ca@�� L��/�$je���軅�{�[/�f�MF���V�T�F8�����,�\x�ϼ�y�_�Y��Ki�+azh�+4����˛W����?�\��{��P@(�+y�%�����C*zk?��K}���{F�-�jb��{��7��q��,;���Vj.1 Gx��C�WQ2�㷉�̻6�;��	Ĳي��/#��^��������b eq�Ǻ� 5L6l��FL��������bՎ��;��j���)B߱�`b��%Z;�8]�[`���X�~��6]��HE�����[�J�~G��3LX,���ґ�E�ex 1���s�0�[4~�z����D����{��tO��ҍ����w ��@y�{��^s���� �\�h� ����g�EB�����1e��Oa��s�����bVX|�ȯ�r��A<�f�5ag�f�7I��m�}Q�~rڱ�%���e�~��ӕ��G뙯����a1�	o��_
�P��;C����!Bk9C���T	�~O���y�����9�߼�>J��2O-�p�E��]\�^7wp�Ų���{�#����ޗ�:ň�Oc=�Oo���\��20�_)��_=�Ξl����l�D[t�@~�����2��!��-Ҫ��=���r�=IXQ�W���P6��׆�����J�9�.�d);�4ZT�3�L��������(Dq������+��'r��j�:т�	ٜ�v0M*~A�������J��GP�c/���N��\.q�k����R�������ɰ�_��oI%%��=l9]�cv�x?�O�� )�^���^H��E���}*�z��g�F�*��f�2ȥD&-���ͤ"�Wp����Ne�@j7�('��^nzc*��`�n�i6� ��X��J}���):��� ����VY�_��_M�}��W�_K�m���h_.���E����-��XK��}�* =�Rm�\�o��Vn'	�Y�;�r��R�ό� �L����ir/�ޤ�F�!�(8΢��Д�a�R��^-U$:a����x������9l�D��_�і�W�YR�/4�~�,�#�g���;y��d�(9�����A�y��u��7Y��D�4B����Ͻ�1~�_:+[�g��9��cNZے��ׯn2?�4�g�Z]�����B��K�2����^n;ݖ�8���'�yZJ^KS��ƀh<y'��4�#��)��U��H�
�;�~u���"��|ι�veǫ
u*��ZZ~�Xw���4�8%H�:������\Nc�u��3��D7����4�`�g�6H����s}=���U��ؕB�LC�7k�͏��d�8�v�� �'��/9P~�J�(dg5lu�����=�<ے�� �1V��
и�Q��x	d�rNn߈	���E�)Kv�2Y�ƚ��f��H��(�g��=hg�`�c���S#�џ��k�ߩ����f7]�R�@%{P-�9�\3���9� �B���0��	K�-k��;�/:bU~M�Dʩ�xW���>~1�>�bY~z��@McM�sK�WF��#?�G^�K��(��D���mX�@j1������CmtZ��P�ƳMe������Q�S� �K�i�c���p�z��+0O^���]IU���s3�T3�pEUft|�E�8(��"{i����1�_7<IB�\Q����W�_�S��i���(�0=���f�Z+G$�' +Z��|�rt�#3F<A>�BH�x���)�t���XMBMG#<X�X	9gê����M�BRt��|��4�H~X\g.��d��������׉u�(�B⮃_���,�z�4��tf��0@��(g�kk��u;�~��9��|,n�∐=�Ԃ���*�s* A�d�K��Y��&��_�-mLo�lc��OҴ���3� �#�0OLr�lf��8������gB[_���WXy��`j<&�a����<o(���q><�&��z�Kĭs_ݛ~0p`H\�]��m��i���+�������s1�Ea����sp���K
p�A�F��_X1�@������n���4���Xlg�����N��|�����8/ ��Jzs�4.�wA�$����%D�*O�;�L�_�~�{0~�wx��V�Ɨ���x �d��ˊr��r�陻)�)���-���mw�~�?��Tn������B_���
(�]5��W3�F���+��47+qU����'�jR��媅ɽ�_�V�:�պ��4Z^IZW6��+,�NC��!�r�5�B/�S�t�O@�bUW2��`��%���6c����W���3M�{vv&nJUލ[�sݘ.(�)��i��K�]��vcu�J�L\<���<�����։�4@qE��/�������E�O���4}=�&s��% 9rm�-�i�e���$ϐ"a��8d���@�?;�a���ϓ�o��F�$�ꝹF@�:�����$HӋ^<H�Qr�z$�ptdY�Ҟ�g��9NLG@�)���e 6$m�@}�	@W7Lej�6!�}n"������������"��#��\��s�q�
�8-��m�k=}�� �����a>.;�_���. �B���Z�^����}��|�n�RN�O���c��:T�ө(���>�C�Lݙ�DS#��B�d����o���7���i�g~O��G�x�Z�fn�69�oo�To�զ-\��Č�ގ�ˈn�6le{�L���f7�KpXD��AW�rgO\~�珳9�_5�I#W*�Ȇk*=g$4ʾ1��a��E�� ���)U���ف�m��������e���x���#@�ﭼ�`��ԫ�Iz����� <�m���ʄ�� ��ز�0��ō3��`��ŗL
,Z��a�N,H�0�e�d��ś�U�NēI������UU>M��m��A~~6۾�ޥ�\.�3���di���'�A����ϩ�mަ�b�)N�ȣ����\?09�Z�D���d65�)����v�\�������qhN��\Rgj#���!�,6�"^�QG-�J������"VCX�_�l�N�J����R�TX�I��9�{�A�;m�i��:�F�P���ń*�:߲�E�w��S���L�����yf�� �,[1x�"��1N�(􏁫c��+�)§ᇗ�p�U㗣�fX��*�,w釭�i|fdϧ,�T@��(��#.>�r%���2U59���"^� <`��%k�݊l�P��_��%͛�:<7[�	o	�N�ڪ4���2��V��^���M�4����_�R�C1l9Ӷ��$ ^Ҡzy��DtI_Nz�{��\B��m�X2�S��l�B�/iixU������9�K�<3Y+��L3�rF��T�?��Y��b�JS��&��P�M��nء� j�SXӼ��
i�x��,e��������l���H��0d����@o�����c�w���]k�w� U'1��C��`�D��T�+5�qf��T�~�f�p�Q)������c�&N1!
�c��  &�r�����U��Fl�R�r��( �r~�*���f�<���=r�����a�܆*0)Ԉ��e�����ω��}�b��(�$\y.-���d���_��Q�O\6�K��K��f��GD��sM9.���o���ɖ#�P@��l)�r "81��j� �v������Q�n�w�$���Q1ݤ�B�����H	o���!|�W<��p�z�����q�^�!�tc����'�d3�ܾO����T<r[�P��-�OmLV6� e\�l��@w���vPE'���N��R^�8[��$u�J�/�E}�b:F�A�}]RyX�	40�g���dt��$���0pf���������(���C�A�_bH幷L�w3/D��R��@���4�~���
A��2\i��ʝ��*~� 

�C�: ��>f#��.m�؋����~�?n���XY��[`�
65;�ϡ��]�R�`�>3�vQ�D��xIT"*��@n�������7�)aK�m7�XJ">���^6EJ�[��V_H|�_v��c�V�=H���\xG���v�7=f�^h+�=G�t�}e�A��@�M>��ƈ#���ÿD����5���>L���e#���< �:V|"���\2��\���!���ޯ�j���z��Y����ކvW��΂�n�ne	e�DU�S{1
��Fk�}]��	�݁𕀻���m啙U*pB�yĀA�yE"�b�N���yƂw�d���?�	w���~�Ls���gӎ��.�d%{�q?V�.��ߖ��t�i;Wkla���k�6Ъ�]}�HΌl��I�d�f�"��*��^�u���c�����]���#��B5�Q�۳,^�춐�~�r�x�'�-<���0,�P �Pًi��"9�Ưh�
tW��k������L2x�@��(���g�	�k��x{"ّ��l�)l0��v��Q�DcTE�C�N��eڳ&e��Kׁ�jVm��F\Y��c��{9?��@(�����6#����*)�vh1P�nZ��k��	t��ܵh��9G6>9�Q=q9�4�P�g��A)����-�Z��`���e����x���Ol��x�Á�_��n�K�Viq�$�٬ِ2_�^\i��g��<�=sw�`�2�*m+��w����D�k2��}=�i���hj�T�RlJ	�>Pn-����y�	����j0��P������S�t%�ܪ�������l�Tr����ˣ�8���5v����7}�ޖ�}�����]"�<_����?�E��JmEP�Bx>�G.�Dd�FM[��=�݃|���PB/0����T?�C�I@̗%*ǘnc$��t��se
�Y��}�M��t$I`5A�T�'H�N��P���2���'��S�v�ԋ�mҧ��8����$��D����$ip'�������R#�9��Z����8���bl�2�pPN|N	꫞W��]//!��=i`+B�nH+���v~(���G7=����-{W�X�7�G;;�$�|��o���%ul,�i���3�� �~"�������ӼgY��5Z[�O���U���SW��G<�ʦ���Iq i��X�I=�Z���X/�&9��"0*HÎ���"��[1�|��ļaf�H�T��Q�M�ȍ$�!��V�"�W��"�(G�^U�<lM����%{�c;�}Tʟ����9�q�C�{q` |�3$~jx�%j��*�X���M��1ʔ`��?�[�Im$���i?ːn���~/��������u��e�^x�$x�=#��a���
W*���3�0\��D��|�tözqzD\yW�5]ra5��|o��wP �@~�0�|��)��AyP�O�Z$��!��[%o\�����R����R��y��Do?�#��c���tѨm����u���<Ψ���=����NsC�&ŕi&����sJ��D������%	�`>1����.b���YG�b������P�,ӗ?�F;i ��r7A}^����Ͼr�9��*PFlgl������W{��ӖHae�!����]��OH�φ�E�������7o)�d��,
z�,�XZ°�$?�Z!�(��}�C�t��0��l��������k��l���Ω�4@$@e��\���̝�Z�^劽}	u�����]�|UH����#�	���11�l����<�����Vc�����;� ��~��F���.�ޅ
��#��J���͸�Ɂ�y�����B�&3��f�A�Ԓ�j�kRt�X�"�£S_f|5Hh{�ư���ͩ/��Ä'�X�zD��ݭ�Qh�*�91X2�Vx�m���7c|��,q�Wg��,�"�����^������hB����}�kv��:�f��xD"�z�UB*Z������{!5����^t��!�"����<��*ݬͶ���K��3��ǚ�;z�-S���P�Qܲ�J!s{�վ���]^�I^��¯2?�Q�
��d��.�o��������(Ѵ!�`���*�f�#�KV�k5�t�C;s��e���
���KU��L���+��\FI����9(���N�_��p�RU�_��)�<XyY::�:%�:�a��1~^�����,�KR�s���Cϩ�$Ϋ����\��ܜ�"�3�iY�M���+ �������k�ᕭ�����@�O�<y��
kw�9J}m,�1e�`c@��>�z{�Wż@�K8�͇_[�k�T*L�Lk�e+N�׋��k��NGk�=��ꍋZ:����m�F�*�l~�N�+r"�.^υ�)e�����°���x/Y�*
�Y�,�a��� ����3�Fn^�[gL���;�;��ɖ��ʵ�-��}�A�'�T�?�9��uF�y��Y������Fjlѡ%<��q��/��7����ٮF:o��i���������l�N�<�8��v,=ȝ�����B����|Po!i���<��|��[?�F1�]3iM�l���0�A��Ї�Os+���67\�5x�y-+��!}c���F@��t��n�Q��ګI�?庛��V�wSgӢ��z�ǐ-S@M4^5�/�@]��FǛ�6|��5��}����˔N#co�{u+�j�v�4(��.I4�����">f��~BG�eER~�Tz	��r��KFsҸs�N���^N��v���i��A��H>�N<��Ӯ�vg��p%eu%��
��7k�ִ3<�������`	� �s�{�u�|>�30�%(����mQ,�NBe|ͳ��� ��3���u�B�_��{mJ�i�/�9�U�3��ǝ�O�sg���{�T� �<	�nڧ^�h[�zV���F4����i��s>��g�d�A.��s��{����U�ԩ����>\^��V�� 87��F�++�HZ��/JU�?p'��`���6=Iĸ+oQt',)yG����
��W/.-{p9Qh��� �����WZ>]�Ru�}J��*n)�<1��Y�|��`sB(�0S
3>�<�9Z��N ��A��ns��6d���Z�b����0E�8�(���zxV��iKX�������yQ$F%�=�f\��Fo�Dt��1�6���HS��7�!,��qw$���qp�q[��u��V�o:W~ͦ�(��iOX��>����V�Q��&^Vz�ż;��VwY{�6��Q��/J#v�лJEç�d��qa8��mI������l>�	����i3�tp��
 �)�V��_�9�����oH��i*��N5$�> C��и�� X4��-�g���?ȱ
)2�|mB�`B��:���$ذ�zPa��v��f�����i�)ֈ�e�D۳�S)S���Y�� 3��e�j��T1�1����QWy��O\Y�z�8�O��0��gy�@QY�;%���:��ފ�vԶ���t-_P�r�_D�j�t�4l�J�t�h�$G@/�R#t�^�x���9\a�c�ih�n�w���T��ϟ�m�{����%5�"M��輡l��q A��l�+@b���ic-�+E��_�#HA������i'9�k�ry-��hK-�m�=�� ��0��r�QFSQ߬�/.��B7�����7���<�����` ���� �i�I��]}��(�5�Q�9ǂ����%�T��, 3a��C�Mx�h���&��JkB-:Mw{���,���Y(\L���	����2q�qf� v�������4KP��3S�?A��͜���Z���>�C���%���>D. �_z����K�|��)��B����ҡ�M�b�%�h��:�[/�^��d͢V+�0�2����u?^�8F�!B�K6�ޅw�<H�uf��ї^)/^[�(u��Ū-#�5nk��K�t�>�3�?��[U�������x�%{r�U���Uy�xAB}�� Qٜ���9�=��2Ȣ;�t	z�U����C�k���&�f�k�����o��O%	��Z:�bH��-��Z24߲�mN"��za7�`6�ڄ�5d�E�u���ni3��t)���s,l�FI%%������^mI��ϭ(�4ܤ@�`�{U��6�K�>����8(�d�F��d7�N�]o=aAC����l|����l����qջI�8�4��Rz+lP��A�Fo�g�J����Zs�����-�c��/��%�k�4C��D�*عٵ���H#SNu�P*J��A��y���������F�cK�'afB�ޮW��(ŉQ��� �]��P%�C��Z�b�{ :G��R&��~YpC����N�p%^���qGM��oAi���ב�V&���trӳ4�l���m� ���V>Z=3�u�a�����V6��b��s��;:ƅ֪�ʂZ	��\�����Q����ʐ1\��J#��8� ���n�Z�ѱ䤊Z�`�}xO��m�pn����Q�����e��d��T�E�Q)WX�^�A�\��+��U3oy�V�R�9<v�I�&��,�_���ݹ�|+Y��FVRQ��v��4E��g�D����+v�0�S�	owDE#&yL��8ט}=���{?�(w���@�� �֋���y�,&a`9$����h0z=2�r��)=�"��JZ'��%�ɻ���$c&Kϙ<�y;����
��jDK�	���"͐6s0�Ϡ����EC�۲Z��3�=�C��-������X�!Ze,�0���}V��Ac�*�嵽|�1Z�ʻ|���~I�Qy�+�ܔ��Zf�>Z�$�Ϣ-��i�/�ta8�хU�ZB��H,�fl#�K���$O�M��e�;�|ޅ�|46�S��̝Q�
g�T=f�1��C��S��r��c�����)vXa��&q�Wn�#G98:�m�I��u#	xRC:vWD�*7j���q.��OƗc� ����BQ1VP����!E))�	� ��`�jW{]�K��S��Au���Z�X%�BBG�48�O���@t����i���]*s�V�
��׹6���{�R$���6!Yù��¾���O�Wm��l��e���d`�6�x����v�Q�)q���Rk�.Д��
�ډRS>ɡA&���*�>�\�|�r@)�U���i(C�ɨ�q=�@0rjg3cf�L`-@�n���yO���:�b�г]s��YJ���w�<�y۷ry�B��Fl�7s��*���ʳx���a��gO;]�[>���XU{�e����4H:W�����q�hq@^�;�d}���[��ӗ^b����z�!v��ai3�j�kG�R�c��%Va�B�x�D��#�y<�qʙ�!�6d�^���/ޝ#f@~��:��:K�}[���������	�����|qǍCR�#����4��g^���˯��tU����g5�<�-���l���U���~q��P�霸���t�wj�B�B��w�T�B��0��#���8�A��IeSY���X��p2�W{i�f
�gE�4�Z��n�$�n�H2=����AgJ࿶��[�"�ߌ�2�2�J ���z��*�6%��-�Tss�:^u��r�"�2C�*����@�����J������~]X�\�;�ݳ'i##$SE�E�fz�c�rv���p��� �^4q��Ig�(i�����:+>V��6#_s��n&))j��^�t:t�N�$p+Ov�;a�`�@t>Pj�%~S)�h��ӸN-ttn Ԯ:)w��1�ɴ��ӂ~�o��N$�^Q�+~�)(U��$G�u�
K!��ck�NylX��q�]�R�8k���i-���؆��K�Ɵ#n����.G��k�:�{�.Ǒ&BR���q-p�ewߎ/�WP� ��NQ_s��Y䦥K~����,�s&�I:��Kl��e_��pmM��r��e��5�Lx�`�-�ă'��([�H8j��Dp�#�UPx�W����V5�M�t�Y
��h.Z�J5
�ڝq��$Yh�J��=�B� �Q?�H;���,M�N/]�!���{�_�.�'A�'+��_3t�f���Gx���J���$���!���B�ڊd��t�U4�� ��:�K��������cy�A�g46�����F8J�����b$X�f��	\�Xf��5�Qh�������NX�ӥ
@VX�B3�l�ԉ.�`�\�������O�r�^����%�'!)�V�����(��Iv=ʺ�(�7��mcr�zK�?�2\��YW�^'��T^k�3!r>�.�u�bb�'�����Gc�Ũ%��a��i��I ���(*�+��aO���<9�c(G��z>�p�H6�­�e�K���.������}ԟ0�����.}ӷޫ�
h���5��4��	��E&��MZ�}�y�D>��@Y��G������C��ӹ����+N9R��J<��!��W��s�i�y�eC3>�l����[�#\E	ʄ[��=m2z���-�$�0����2��6�>B�g7����>��S��pWM�>g�iJ^�(�Iճ7�@e���G�{WH]�iw3_aۡs$z,j��Up�,bܮ�P�Tz���v���u��vjT��!
_
^U!�5p7V��?��[���
�~Kk=�̟)��y�`�b�\0h��������;�� �I��	TVA�(+�nZ�?�y�1�F����z��?��������N��t�kFȫ2���a衐�7h��^F�yE+V�)�E)|�p��"�v��4ڐHZ��e���ȇ��t��{�,p2��D}�KA����?pdJ7m������"sB��ZUZ��r�xn�u^%8IQ5[@��I�%�ՙ�[���m�F"O�Z�
�$4���S�\8�pW�M�Y���{�YOdKũ!�!bk�#�yZ-�>�J����� D�a1����"��ƈ���h1���&W��3�\&�6}X�Ȣ>a>9��PQR�d�ÄA�П	z,L	4-hJr�a7����e�v��1)�_����K��ϖ$�|�P-�	ȵm��8^�L�Q�����ݓ���|԰��zc�	b��G�K���?�/��C��8�~P�^��1�_��G�*p:�����,6U'ڬ��t߰���*7ww�#��'C��F�S>�_B�J�_i�kq�VZ��S���J�����Td��
!��\v��Ɗ�U�C?�ݔB�o4�ӵa`D�.q`b��&7[�1c�5^�^�,񉀰f�%~w=C1T�j�_+�$�����$o >������}���*�fd	��#k=lE6d�`���u��K�<0O�P�-d�
jT�Ƭe
�8�@��4%�B{T]�-��o �鵤�n0EYw˱K��EzgH�!�"�^�v���k>�n?�0���B�#�Y6���	J��^#/���`��Q�8�Ǖl|Ůn�h���SuW�B2G8�H�T_��6B�X���v�H��ژCr*�~3K	3|������7 �������% ��0�t���zΊ��/�ߪd�0��ڢ�3v����58Tŀ�<��N�� X��ez��+2�D���s��֠���	��e�2��@��u��L�h��XuA���}%�J��g���5���
+���'p(N+_�]؟��ٲb�g�CY��X&�E�o������M�OQ��]�ȕ8Q��_Xw�ڹ�]w�5+!�|����@�[�`x�-� �]+�j�mT �pX�E��P2j�Ѩ�����.�>B~QJ�L�����<�#;�8ҁ@3������
�pښ"�;T ����S�=�M�-�������znt��L��aQ���d�Y!R؃�(kZ�%q������;y���h��� �K/�q�kC>y��TXѩ���\&$2B�H�⩆�i⋤��S\jr��z_j�t��cZ������umLgRT@�r�q���.���W�BH���U���T��Nw�p�z*bϩd?�$I���r��pET��˃gd�p v���S�N�9S���|kh�fݥ�KcT�9���X֪����b&'��tw���3 U�-�!Lk�m�}6)�\�1��QM��CS�}��#x�`��B�td� �iѯG,����tŊ�5��Z0���Y!��.��금�����^A������7�P�x���F_0�"r�>RD��Oj���P��UcV��$�������9�,3� �l�����Vc�����I�g��K�[�W�q�I0�Ȑ{T���	̋�nPf�� c�x/���|y�d��_�����4}UJf-�6t�HY��O�HD�/�� �|�Oo��ͼ�� x� Rd0;��R�V�V2;�ɠQ������	Zȿ$̖���*uY������M���ю�؞���
&f�ν-����j��@!}:�hY���׵��V��5V�!˃n�v��}����J��e3���R&a��S�v!���J�6ഏW��%���̛�9��������d"I:֓�,3Ԩ;;`�cg�m��b�Cq�Q���D�J}����s9��x��h��6���-��9�ʘX�C���|~�ل�%N��"�,;��#��.I�
Tס���|j+�ٖs"�W^i�Q�"K��M�Of����{�$.��P}e�Ǌ� L;b�@��%������[8rQ>Mԯ!�V6���*�{-�?�z�4��i����"j7���Q%����~��+#�F�Oՙ�ݸ�%�I��ڰ�R�ů��]�SW��d�x���T5g��Eˏ��`I�Y�
~#�+e�sҜ�5�O��G,�>�1>e��T+��#�i������4�m��[�	n�Q�����}5���ܘ�@�/yA�sIW�jh�u�'=_1e�l�4�������
�&�sT�2�A�_�Ů�y��y��D��B�Ȯ��(C+�S� �=�xQz�[�^�����������JvK.�
f�R�Ez�[�ɐl��% O����E~P���8Ȅ�����9H���~fovI���q?gH�@�@�8E#�Dj%�F�IP;S�%a��{Zj��zI�Kr�X��w-��s�ꟿ��k*�'���5�m G�g�ݷ"%/b�4��J�����;���&j�U��M�zO>(�S$��~��7��
\���*x�>#��~C<b�[�h��z�w=L���Yg���-yHLx�( �zLzH��0-�/�~ �bƕjK��y'-|G#�hU~�����m��I��U:+�k��|Z��	|gL� !��r�
!&qy�79G���r�t@�gAG�#�܂��)�'j6K�����n]���>��-4Ϛ�q&ej�� ����7��9����X#[�0훽�	�Q�Dm�����D�	�֋���{������h���"�;^���vK�щ����ʻG���ָ�ߖ��fn�f���=�J968�K��>PPQi����:B�/0n^wI��i��	$İ*-���*��iĚ>�H� K�� $�o��K��r*f�4Y�� vv�x9�:�e��~X��=�OG��P�R_�V|$w�h2�9��>�W@9�aw�7��m�o"���p�ۢ[d���R�f���Im�q��e[�7�_��O�Rc�2wb:� �R��=5�Ag�Ns`_5��c�=z��D�L$ˁL��x�]��_���e��ya�v��u�t�����c�F�C1�\�p,�Ö�GH������{���Jk����bZ+K�\l�-H�R55�n� ���w���/�7OQ��W��`���g{Z�
�/1��e���q!��v\��Bg3=�ʨ��*�S�%�i�����aG2���ʗ�� �[��Gڶ����|֙�NP2��O�ӽ*��X�󫊦Fn�(��ǿT��a����~m��$~aX?��U:"��/�'m;7~��/��C@�}_N���@����D����؈����8���jSX޲��7X6�~1�Z\��_\4��:̫�s�'R�W� ��栾$g ��p�T�i��,�Ȣ����b��R6 5Lyjw�̠[�����V�0'�O����5�@G�C�rlkԙ���Y�S�*vY��i"	�l�i0!`�l@g�F��I�a'�U����\��&c�]}����Ygz%�$#��}9�P$*y<Ӎ�]�݈���Cc�]����v|�՝	;]V0�p�m�sxy�]�FL �jC��m�y�%�k�F�j3�<,�4���_�V�Bzv7�U�TrǨq����	Ӱ���G�-y�F}�.n�@�	A�����t �Q ��&��p��:�;`���ԅ���m;�w�+H_�_�Am��0 �����u���B��J���ñ"[E��>���*�'>��	�:}f1Y�B&,|@_5pf+<S��"��5%1;t^�M����z��8�a�#-9��vrK�v `v! �s�	�1��.:�F#�P2㣡��ޱ�������{e�e :xC���	ueP�'�0l/����+*��}r���8Z���>r"A(P�����Jb��eJ�k�!;۳cz '����|:1�r�'vS�G�wr�/B�Ov��)��f���PEz
��q;W�R��h}���D�@����t/��G�¡N���?�y�i��j��e������Jݧ�d1ω��?���ߜ��R-|et�/�V�!��m1��2�V��v�����߆�AAybЇvS2L�>5wཱུ
f�[?�"3+�Mw����L��ȜM��� �׷�2�ˁ��K�dS��}奔�cl&a�mj9pe�@��$���ƣ9/|�P���o/^'yͺЉ���1�|��S��n`�r��߲�·'yx�^ʳ�1a4�=��"nhGꭶ͍�k!��pfbj�a��$R��
�x�o���?�]jY�u46��,S�Ps;-
3�,>��G'b�gz�}s�T��t1�}ًD�e�<��0"�Cɔ�"�ro���>&��22����DZ�d�Q�ڜu��Ne.�C���(�����0�KB��� |�g���F���g�J�t	�'uw^��FcZ�h��eۿZ�Ks
b��st�-hP"�ұ\*��«�����I9mϢa�'-YY��r�,���tK�����@�	���ςC������jM��:]|v"I���}��0ۅ�A=�fr]�\E�g��rz�=��x����Be�$�"z@��y�ͽ�#yWN ��ua���趮�O�ȁ����r���� �rm�=�{���G��*^�?�2����/��nE{�q2D5�q5�|���\����k��`ڛd
8[���}�ΈM���XI\[y�忰	ǩ�跷�������{�� k��a���()���A��U�����&��Y�]b�v_��pQF4�F����PT��~^�#6/O����{�Z^#�8@�5�A��=y��H�JT���W�c�N�pK SI\N�f ڷ$��{sg�Z�e�eI�bx/��p+�䁰o#:�6&&�nn�I�3$��Z{̐�t�I����U�{F<*���g���"ִ�D�c����:�����ƣʛ� y_ma<��`�[״CM����f�A�!C��QQ���m0���l�l�S}��wp�Y��m%NF�Ld����g1(��C�L���-����|ů͟���<C��:��0�U�qLv�.@�����m��z:b��#��U�����;�7}Z5��pěd�y�X~��w1�1�c-]ρ������N{�~� ��4��
�A!��2!
���D0�Y.3�x:���Ճ\9�I���Rp2��K��J"�_%O�-����^V������	Y_����Y���D�-�䑄.k���H�;�ȹ"�8�m�X+6�ۼ*�rY�@�Ї��&X�`��G�U�&�N_��AU�H�.P_��&mwÃyj�Չ�&C�|}ېn�+���@�f�40�B�'MP��^�Ч]�9�bd��m�9��Ȑ$�t�|�]�;��Ҋ��ҷe��LL�5�G�?��:�CRܤB�?03���o;hW����I�"�̎�$ȖDq�Uy��û���%0����eQ���,���m���
�-�L
}D���j{���כ��$���P�2׊2E����
��op��K�բQ
��G�Cg#�g�;'��C�;N��#��r�	�w��'�n����EOrPު�O�#�������\�Mu^�Eu�إ�Ez��H�/P�n ��)�X�I�a��^֭lT�Y�OS�U�3��Q+�1��[J~�ٸ:�e	����P�q3�0p�c��@����C��>@����8���K�M���_2��
�(�h)���Y���yDqBl�P��"?�a�$�xV��#��u<�(���8G��p����5��G�3���G)
꣧�� +h2�y`r:M��`��nk�G�Qt!nۮ�ڌ�(�30�#�B���R�\���z�� t��lP��'�5�|��'e��3Qo��d9�	$�`b�7�O.-ٮ���2�~F�ܗf��T|�|��LO�68��D�5<Ʌ������"���J������,����]AɎ2.�&=���]0�D�:'{;[�o��Ǐ���pw�ul�yܨ��t�1� ��4�PPzG4µ�V짉�a���S�(;�כ�`g����	D���K�L�[_e*~d�}���k�,�-�V�9�^��\���wñN��G4+-����FM��Ɛ��~kXm�8H�����?�$�����E:)D��ky�{�p�+G@�uR�n�XM�X�!l:�:��c,�}�W:�na`�!�8F0�8.��r�U?�)�����U���n�$���-�45A��*�5nm���8Y�ig{R�Cʊ�*�万�(�Y��}�%λ����o����R�׳Hy�u�I��.�ntv��gi�*�����]{PKU?3��*���S�-���R`׾e�!�s��QJ�Ţ`����V잼p�l�W��=��H8�T�=��=�4��`FzOs_�f�gg�q�"��hn�E�*����1y ����f7���K�K%��`�sK:Up�������y�)=a>>��}�ͺ\a.@.CFF)�L��p7jw��d)�ƴm%�,�L2�"?(a��z��+��FT�:	t%�@�F��5-�����M��:y~��*ɳm#��Q�Lhmz��7�̸�
�װ��ڐ�S�!��
,������r��D�A3}�TBC��
�a�ɔ��!]z^$)������%Ǣ�	�R��mp7�X�VK$��L���a��K�{0�mQP�r�s����j:~�&|e�jqug`�}�����q���B�{i8m�b�V�P�C'g�"�׉-�e���&t�Дk��ߐ��X�K�.^y��?k&�d!��'q��i+�6��0�����歺�惍03��Kk�Eҕ�C���b�j'�@� �S�x�7	���=����F�5������u0�kr�����������%K���~���3cR���-p�&��?��e��ţYR��;CW�"�ö���iŬ_���K�8�6�5u��6KG9��8:j�v�;�(jR/�)�o�����O	ViE�4uzPNA��>{o���XEc,��3.�Oɱt��Y]��ǀ��e�)ћQ���3�s���ţ�һ�R7��Bʖ���s���8 ��,�ky�V�3��%t:�ڮ�Пp���{�Ӽ�ԧ�[�v���D�c8q���`>P�����OvX䢄��0�'B�=2��]bR��g�2���;�cq��55�ì����Ǆ���K���s���X��v\��{k�ZO�:g|�S��ѝ����j�l�꫽�0��Z�����au'n��pN0j� ��5���W|�Q�F��E�����G<㘋�s��a"M����H F���B�,ҞZ(G��
��_[��$���:���w)x�������i��}N&t��ܭ���m�:8�?M$Q���g\�E1�pG#Y����nӵʻD�z�� H*ġ���F�F�1p�&��T�Y�pDRײ���{�� �9_��I�����((i��'�QI{T�\�c� t5�	wE�`�&���9�hsX���O���Á\<aJBuZU��ͺUL�:��scGl�-������Kl�*J��-ӝQ.�;��"������>�:��iQ��4�8T8(_rΔ8�s����.W�;� �h}N]Hޮ_줦��%R񓆖;�1 �'��
������Vd�t�¯�e(�����8��b��ZP�RH虁�a�~�u���s��D��-@��*�o&b��u"q-�΁�k�ЩlR2=
�9�X�x�J�x�0Ɯ!�����O�h�ٗm�ޟ����b��n�����9����p� 6Cr��fWU ��X�Ma����D�|��܈����O�-���p�?i�GW�M7��ͫ�.)�E��w| �Oך�];ݧ+#
��mF���ְ�� ��
��8�F�p���˭�\��~�@h��^DQ��\� R�A� ��e�b��r��!��.[SA��g=�g!b��<�/��-����)�i`ᠴ�86��A�����B�a�z޳\�*Xs˥��P��Rϯ���#�����������9�L�A��A�/���_��w��GQ�������Xe���[��R�|g��(!]��h�BαA8Dm�e��4.$�e�I���f)�3/�	M
p�ų˨~����l�����0򸯵��j*� ��Ġ׋a����hUu��Ul���P��
�E��2�*�e����=��9a��k�c�2�tଶ�B�O�����,��
;2�T��Q)
;����K����[��� �3Z"�v�]�˙/�G�������j�q������F�5Q_��R0CzE����� ;z#�l#U�b�*�tj�QǉH��J�H���n��(�b��
���*{����t����.;.�F�߷�d��o���J�p�`}�Fx�Ӵ��T����ue�ju�������Ϡ�����o�m�_s�7����-���$j�9�4W����a��ʉ	K��m�H/�;^N?�f���9��\�@S�5���;�m<Ɋ��(�I�]�u� ���".|��D'0=���qx��œ)�b
e�9m�˷���3��$���}�K�h@0��o�	Q�gZh)���]t�{�()Q��n�7kK_��~�S�v�ϕ��	��s���u�n��~��R�=���t���
�R?�7 dP2�j�f��Z�8��I�IOQ��s1+\��N�
]8	A��F0��cf��hn��:a1���r��� ���h��F;�������d�3j���4�[ӡ�KI�����!u#��'����3�*����ݲ8�z�Б-�0����*��L�'gy�����x*[^`���l:#7�����_�2���5���Ð�oׄ't���G�y��Ֆ�^hVi�@�\xz$~�2�ڥ�[����ƛ�g: ��&�	��\�����֊6p�Y���U������)����˔���U_�|;�7��.9�2�0F������k9QY7����(��N�]�D�qi�A@pȴ;��끰�5��rwKy8�rk��\�y�|8W�M��Q��R>/�]���٢�̩0Q{��O��=�*&�}7�\o�i���=��1�(�Le�Х�y�#��r��s��+��N�����2{ؔ��yW���ݍLi��_~仺� �ǵS�t�.��.HǙ��BN+Hd�I)V�svBְ��!�d�$�����/�3�Fq-�����G���c �<��Ν��R�+��SxY��t�Fز��aBſ$ �դǂ��@<�z��{�G�H΍���"�o��L��;8�����\�V� �l�Ѡk�����R�82&�ll�W��9x�
 -+|�l�_J�H��(YjR/)F����>�7�����$�G�-t	��j��p*�_ML�����L�4�����M���>9N������P���;a8`kO�f�-u��O7:��	L���[ n�:iS�HamR�����ϿWM�k\"�U㝣�;%���:���Y{}z���[�H5�M�3��t<��ӋP�-�9�0f�Xڹ��m�OI���zz�@�Y�?M�9Ycf�����ʎ��oM�m�a�+��ǒ�ݶW�9v@g��C����t/j�ڪ�-�l�����T�&*��ΰ���F�C�	*fG��=m����c�Ҝ���V����ݭ�`��U��T�NWO�x�8U�u`��~a�!X��T��C�'��ƪ8�[	e�1�׌�	Q7/�[�sٗ&��
�0? b3|a&�9����-7|3i'�p����B!�񃑈r�����ciKp���0n�����Y��l�\m��j������L)g��~��|��*�ɞ�,����	l�|�da���F�&���:w<347�@��+j����x��^��U��##��mG��)�|�z�2�J נ�]�ɞ')��͒��
l�9�N������V���0G��6�¯s�>(7�ǂ&��z�(H��aT��(��No6����-=�M�"�0}Yik����F��TlG`��(�+�!Nso�j�$��β��l�ɮ�)����Rq�F�B����{�Hև�����~���6�{h��}B♵��1��M
�gY�o?帠7�`�RcX���>�����)\Ea�;a�4>���|�U8�A*�b%���'+t]QI(��O��<����dj(�L$���o��w�n���F�Q�v1I��J� *����"�vF����f���2N����Ac�n,���R�<���Xߘa��&	*�-��ia��J�q����rH,u�B/��Uv)�1˗�v�ke��Kp�+�Pe��*�����6��&>�ď 31�a���窷3WE�jm�o�����,R�K#�ܛ�W�$'���+�]"�.���c�e�/��w8l��^<����2؋/�yNx)�=�H�aE0z4���^.�&b�V�BV���Ѭ߫Ȃ�\�V����T�.��*�%h�,�����x�_�2�i9�;Q����r�s����?�m���6� ]f�[� 8����ĵ�e/_���˼b6t���"�w�)�y읻>��h۝)�GѨ�3�Ll�
��SRx��K1Rh��Pa� ��},��l%i/��ޡ�\�쉆�ġ�Zu���' z�gG���uѶ��h=ކ�+U���;��.�����t\��vKv�P�w�!g��H����)egH�j���],Z���^�G�Zjʆ�Аᶻ`��ԩ�#��'�A�*��ճ���?Pm�@�f�+4{\W�0�Nhϫ�/��R�/g�b 6�X��5�f1M�����T�P{�jxW"*aT��<ňN>X��6�w�I�U��A�E��g6�w��%-pjfI�㤫�<��{��b����>1�v7��d��-�z��0�	�S�/�5�����C��S��ˈ�8Y�]�n���Wr@[��@��{4G����2�.��!�z҇!4����8V(�%��{(T��U�^
�����n`�.���X�բ��C_��Im?Ռ+9�$1n����>��^`��nH#$d��x��X�bw���a^Q�|)�����P�E��d���OI�{��X�� �C��	3GIr�"���2�d5x���R��;�L�:�wO������Y����ߠ �=U��;�H1@�~j�n7%�qH�qz���v�uFTy#}��k��ݬ`gϴ���$730~�s�[��)����L���z&p�c��`=�N�@�*��3B��Uk*�r6�;�1l�rL����@ˏj�4o�F�")�D�2<���@ݏV�P���G&tk1�τ�p�Žlr3ℴ�9u{�j���곲�!�����f�S�0k&�1��{�B���*�Ю88W�"��t�Ͷ:���I�8��[V�g����Y�J#K# ���R X@ڬ�4��N��Q��r������S�G	�x�&��*��pܦ1R�r�������6�(kK۴V�s�}�S�w��\�;==�p(V�g��3i��`j!D��YW����	X��4t��.쟒�Wi�TQ��̠�N��}������H{�|�?���/ ͷ�F�f LF��?�DI��1&X�Q�����6q�����N�v��Q�����\�MA;�Y�~�2~����RH��H���@C�7��+m�=
|�և/���~��o�0�,3�� N��C���P����Xy~�[���P5q|\*^M�\���ΓB���,��"ڌJ�+?SH�v�_)�L�Y�d���AE�*����^��A
WG��#�:��sٵ��ObK�z���7<e��0�~sI.�I`�31��d������N���0�g�1�J�,l�匟Ql���r�DT�+���g��Ji{��W���J9}�tQ���I�8�`��Ж8��@�� B/5��"�^�?>v�Ϋ�VR�P��n��[n��-��r�[2QYU�����|Pl��	�OH�߻p��9N�i+�N��{���ɜԪ����,u�)���{�����AV��8
E!`eY��,���f1kğ$#���S�>��=wF��#��[N����t���q�bЭD�!%@z�3R���\D���2@� ��O-�r�6X�[��
�&1�F�M��=l-�����<K��uE%]>��H��}SX�Т�^�T{�w���}�G���׍~��Or�ۺ"�	�'j=�����'���Zf����"�#)�YJ�����^VBX��9��}�'+�H@�'d�Xg鹙;�$�[[����V�t�8�w����tX���q�������]
�n�j�[�Gok�|AF_0q���kQg�h��p��,��Z��+�= {2�L���X�q�\���n���3[��^ͨ���xw.�2Ɉ<�1�@'B-��n��Q�x�Js�ֻn$~�H]�����>�9����/�|"�//���?6�cϏ���0��X��f��{��P�f���~̜�o��5����b�II�m��-���֨u,'�;ᨃCً15�J-[���H�
������~*����vK�h�M������S�~B��<[�\�2:L���G���P��=�W���f�>9~��	�^�}�����
����Bd�F�A��I>c0TS�ĉ=Kn�;y���4�;�H�[O�B�Y���a�4X�0�v�\.^�~����~������X��7e��t-�(?��ͅd	}�+�Z����@.uW��|g8� �"yM^�#k�K�(hH�|A2ؽx0��I��W9U!�,�5`��^Y�E.�U���,�ZV���ccӠ��q~1�_��'�{W�w�'nK�`R�|O�"͠l'<�`�q��Aw�0 �x�G"*���8 �*��0O*�&�͠������kw3 =��ml�8mJ��b���Տ��mYf��������MPC0�q&�J�X���D�a��J�幚�Hs������n�@�,wc��k��Gկ���=�8��S�Ɛy��lAVX�L�B[�r\�������&���jb/U���9����$]�m_��]�J�4�rL��è�6�󀦌g�� �� �&�k?�tQ�}�#m��T��/G#p}�K�/�f�UOB�����{{X����.8�n�@��8�ô�����B��=�7�TǏ��J�d�����2����.T#(��^�nܞ�BA���jb��g�7Ƒ^��I��{���KI��o/M�.��R��1��_7'ͮ�"����fc3�����S��ɀU����`���<�X�ҍ�Fj��;��hU�c�4�/�)$w��c���d��K�l5ѷ����X��y�?�T�/�^���2�5⃀��?�F��et�1�:7��r�DSja*p�>�g��Č���n���N@O�o[xgI�� �ڤY>$���j^�:2Ƶ��#S���l ?��|	��_�@�`�������è	�s�NM��5S��1��泰���^,�J�ˤ�KY�7��ci�����q"�YR�@�<h�lI���8|�r��N89.�2�*Z�<����
�O����b�A3���D�����k�>@�c!
U���N�c�`�hW��������	�%'�c����,�A���2��gP���L���~�IW�
��j���*�� �=�;�(����N�z��W�P?j,�`4�.%Jc�Pb<�>��4Lt|f��I��Z�̀���Dyb�� �>n�������D8����E��3�¡��A�=�P���6����+m���}����~�#A�g��{�kJN�Y��$!�����p��Í�B��\sٯ�p���-�v�=U].���d�������bt�����4^�䔫�0�B�a������c���s�ٍ��%���:P9i�D������ V����� ��>�
qjb�Y����_�jh���Z������2N l���o��M�����m5�7�JW�咀g���?�+��rNÝ��t��H��h��쾻���/��h��$��u�@���}����E�-�-'�T��.�C��I���^��4N��&�3I�;�w��J^�Ã
��U�Ϣ޺/�1��6���O��N�1���4�.�$[~��jy�}�iS )��^��J��;
���%�!��7�P�"�v�U@^������z�PA+w�fTk�p��{����Xvu�y�Y�Q���ĥj36��`f��� �#QWm�KL�V~��Ջ�QL������JYP����2��8͋[4Ve�'�s�6��ܟ�]>2�����X�%9$��L���r���4�`/��B[]V��q)�ݪ!@R:���%�.t�Ո?�� �c�q��K	�#*�3t�G�tǮ���ǰC`�G Ck�sD
��+M���������?�%�ܳ~.ں,���2��>ĝ�KG3�X|�wЯۙX��^S�i����"��u4p8%+�}-��<�6�l�d�nb�N0�I�d`��l���`D�E��ȇ����GdsT7�� k��E�A���������9zX�\$�C��/[�K=�gP�:b�R�7k������҈`#��[�rI��k2N��I/���,��D�R �&	ƾ�MS��v<��i49~���qw�����򲑾���ڃt]����d�G��x�����W�},5ך�>E��N@Rx�SYnN�����a��	Dv%	�!ط��|�ai����7���T�}&���fSL�h��0@��vx�0�H�f�	[ј��р-���1������G}2U4��f2���5<o_F����NY$����RW~0����NZ�{r��]��=�;���ע{v�=^tv�z` c��]h_��"6&`��)�1ƄDZ�M�._Jۜ����5EW����&y������Ϋ����ι�Jg���t1S�'R[IN��{�te�EB;��S���l���� �k��Y݀���Y��;�1�(`���M����i/���n1p��,=ըYm"M�C��a��Зج�K9c�����g�ٚ+���-YIR+��&��Sb8�'�b��[���rQ���.�!=�钌���/�RP��y�� ��L0L»�W��u7C��
/�\[�7�}�n�T;�����.-�hc!U��p�?6�"AC3�������M��v��v\�/	A�p}{��d��O��/k��v���=���K���Y^���8�8�༺g-q�-�1�,mx�?�)��:�Js���/	|�y0�8��#�ӭ��6ڞA�W�Hx�]���N����8���B�������(�G�{�inrb��Ҡ�>�xx<���\EN�5����܋Q��p��2�1���ZV��!�[������b��VG�dA����(���D�޷��-ݸFɡ�;��z��� �഍�J�ra��f��}\ٵ,�٫��7�	�+��/W�g�%'����(h' 75ȳ��^<i:���Gx>R�

�
=p5�SD�"ԑ�Q�xш=�ic��(���x��˾t�P�u>�����-r�_W�� ����v��uDȄML�t�z���ܻ���Za��_�^�Laڝ�3��sA̺�uK�h)v�_��#\o�zk��#��f'���^��)�9= x���,t��2�!�$�=G�)z�9�J励������v� �R�2Ze�Ao"�+J�.�����(yPM(�Kwr�� ̜H�ByiV��5��q<��G2P��UU%�@�q�3:j�s!���XO�(��_?�Z��M;* ���۟�"��z�щ�6{s�1��W�}ja�����=�$�"����w��L]in�jB,��N��~�F�Iƃv�I���ě�8T#6�4�V���P©L���64>���Щq��%��c��&���؂VYu
�p�����a��	�t=n��#��S��S���\,ۮ��i"��j���HJQ(W�&�`_q�c��;�9ȗ-�F�MA�H�,��H~�d�d�Ĩm-v���[�G�������X1>�j�S���mf^�WQn_�1ՠu�� |����C�)��1^����d|��,�$U�:�40�>(��&�)��>�j��@\�>�C�����Ӂ_�*��o�cLo�~�`��*��̈�	�>�7���M|,6��e ��CI�MgI������%��\}�<R(	�!�������K�eTg�R���h��^Y}޴��^�i�7u�H�lW��0���Rl�wߣ\N����s�y-[N}J6��=�<�Q��>��&���M��Bv��D�Шi\�ϋT��.���D;F��+eq�}�L'���D�������]�aotf@i��-�N���s�˯�H�|"������������(���0������0%�����[E��gbᘫ�y����ٻ�1�|l�R� (�������x0�d�y:��;.v �@�R.j����⚥�,#� _ƙ2���U޸�ʑ��I����e���Ieڝm���8}U�^�Y�_������ZP�N��Kzщ�h"���"�<V���Hu�J��j7���N��$F���3�������I%s�V�B||ǅ>v,���:c����<�&����WU�l��P���mݒ*�2��5��aU]Cg�
�"�2t�׀DY�X;�^��I�B���l%�͢���3��oT��m�\~�1�K�6n�<�?��=��׊ۮ2�Z��!�y-0�R���VT�U,	��O ,~yWkǸ�R�畞�Ɲ�&�#B��E�o�j�rj����1C��8�0vj���Ae�rv���.�J�2E!E�$�}�L��	%��CX��@���m�ǎ$����+���k����c�=���BܙJ�SQ7���T���R�����Э�o�XG�-��Bײ:pƘ@���+�҃(/[f{��G�Z?�R���$!�\t���h��.�<���+�.��B�ڴ7%*n\����! $5�c�q�y��Y�`����E��a?Ւ�$wm.IT�X $?>5�SӐ_���^,�K	)�F�su}�d0L��+Q|���Z�:���Ű�gF���D����4�:g#�����u�Pǥ�-2{?�R��_"6Τ�	�=�U{����������4�u�y�1i�#\��T�IW�m��f%�#��\�#�S��6:뙊>����$����jZAX�X�/[8
�"�����E���{����M���m�O�R�A�ƾ`F�8p�B O[2ڹR�q���t�׬����������偆��p=��3�o�_F[���h��K�^/K��Y�#cJ�f���>�7	pك���AO���w�fD㉬���	�<�)b�?�/�9O�����Y��^���V���I򅨹[�ǘ�hc�0�����hQ��ϛ��A� +'�Z��g��V(�j�IPo���_��;mo�I�p�	�r��oo�q<J�I��/i�����S?嘃"� ����^4��
�V��s�Q�]E�����U��������n���U`��}:N��8����K�^]��
�����\�}ᒤ�-�ѴC	��:�-�fr��l���HM��Uh�m���M��N�Ç1/T<A��^�j7F��[6�J�~Ñ����G&Qu'�oÄ��9���u���$�\/^��r@�)���pfI�}Iu%h��m�{��߮P���cZ��,��t����u;��赢��Q�4�B?*3̙����P�VZ�a���ex�0�G鑇���4QH:�'5�d��B;_w���5����$q���?*\�����<�?�RX��@L�����C��pp:�c7X`f�mI�@�eUۨ��P�:d���#Yf{`�$ B��D�Ҥ�*����ӌ���⢡h%Se������a��7x�z�jN1�Le�9&� 0y�4�E�E4hY~���DL�ˑ�^��B�_Є�e����5eX�+F J4��N`^;]2�(��&x���!�z��Y�"ʡiY��YҴ���\�P]�B͉����w�L�����2`���r�J[R�4pw�m�=�?�L7d��'�G�`��'VxΒ�!8�m
��T0�Q��x���
o��>��$��ee>a��L��F[�GJ}
��l�x-I���N�(3�3�Dct)��[P&�֌�����%���th���d{�ea���r��-@���-\�jߒ��ƫ�b�;��v��:�s�	Y��k��_�-v�u�6��,q6<�͜V%�]��g2h�ԙ��2���E���76I��$~�'��NT�B_gRX.Śߛ1�]�+��z�-��T3p�h,�㟪��*�"��p�+�a�l�����|��[Mi�>;�\hI��~M^<��gNf.&�B@9�~�Ad`��m�cj���$}�*�:h��k9	Ac7�����Jn�۬������R�}i*�i�A�:��b���z��>m�F�6P����ʪ`K��/.8LI�����nD��sBr#.��0&=�)�1q�(�x���1P�k�݉/D\��#Na'oʛ|ظR�����f�������dyM��<���q����e�@������m���RZ��2V�y����CA} _~�Z7>�R>Iw<���ޞ����W�,=g�s��N�6<P`�*�GM���0#��.#i+	~�C�����G.���Xz���{��T��:3&Bd8̇��E� ��~�>:��q�7��(�'_�*�r�p���w���X�8�	�I����(�/m`���C��(r��a6OIC�"�`ǤL��7�埤��1yx=ӱ�{�ڡ��?d)N��J�h֑=���G��o��fm��λ�2��-���6�s
��PX:*��t�*'V,f�<Jl�&��O�f���ETu���z�y�U�`�
�,!���C��&Ӥ3i;]�/ն� h�oq�ް]�/�Ng'��������%; �Y�R���5��YU~^�i�}'lg�{ F�O�Qٖ*����-i1�٭ay�s���:�#� ]�y����<4��b�%�l��fޢ�üa{����_�py�5�e{nT��s�k�ۦ�'ڵ������9�/u� y�+Du�0n:R��ji���@�o0�v�)������o����ǲ߿�A�^��ԃ{i{=�=d�.��E���A�M�7������>�y�F/���F�X`���Y [:�~T��=5�t�V��&�)<Q`WI1��Ƭz��j�V���ȴ'm:�8䢍y��+Fs3�~�q -�@w���>��l�0	K�>2�q��
��|��\��{hJ�}1!�U�Wj%��r	�Q,K�t��=�0 |%C��O�ޛPһ�2&�Χ��0M$H�
�Z�A�)�ho6~�g��.�wym��f�T�=ۀ&�D8mk�ˤX*��$P<|r�A˰Pc}{-�N��aTOi;�sF�'�*$3�
�2�"�3��C��S��e;�QH	ohk�N���k��7�+؋bC� m�����\�3���n �z�"#p.�_��	����SM��^[��V]��=�5���:�,�]]�9U �u8Yq�
!��b���BL)� _��K�����_	溏�$�:F4: @c �+�nAs��c�6"����[e&��p�-|[�z����d��&Z�v��Mc�eU�P>�DgV�:~"%�&]6�NVpk��	����B�}�ު��TCq2�׷dN����K� �?�Ak��K�x���C����J�
�\B�Z�<mԄ�!��':����7ir��w�>1To2�^��$���DD,j8$��S�<\Nj�?9Xi�"V�g1��Prh���'B�&cU��@�Os�L�'�Xǟ�����p���']��'���Y�-�o[$�+Y�G�zi�V*d�]񷻡&}�.lt�Cl���x�1���N"黎�i�G�V�������]]��{���r���Ƨ�(�i��#M� ��������/T�+ns#�)T&�(��G�l�t��̽�1���v�}��n9�k��5$��2��c`ʱv�*1�}*�A��(ʷ���"��Ad
<LX_���|��u��նd&5(%���5�5��GB�ȧluĨ3ѷ���'�m�L���x=>���_|4��q�aN�{=$��oWV=�8;.�Ɉ�n�Jg{�ֳ��\L8M�
�<���y�#lJ��1��BHr^3����z�s=�u��_<�f��ZN�^21�C��;������_߂��GJp�|U�� �����C�IT6�I�w�L>
k��#�LbN(��_��^�x@�p`�V����L�l"�J�D?�N4�䍇k���C�@��ӽ��%DS�����#)���-�ˉF�R����Ǡ��%�܎Ǖ�[Y���΂'�nrڬ�W+��o��^D�q�z�? ��U4f
۫�jGC1���`(�8z��j����I����C�5�?��t�PP�A�E��#�����h,�)N�]�P<L�
C���X�s5[����P,y2���-�&�[`q�;s���������k��m8[T��?���=�s4B�礿�|,Y�"0��P�Xmz����t�EW�F�*3�T c��;��rF���@����)8�(&z�sG7þ����P�e=%e�j���?Ԁܡ٥e�.]?o�9��rs�$��_��stcJxJm�D��ε3C�Q������LO��O<3���	��0[�:��3W����Q��Z'���@&���Q��y�b��I��(��?�_��^�[E֭K�&t�#}\R��1R�5������V(V%�?�j>Gm��^�=�H�m�>��#>�DLl��[��d�[L��.�N�]�'+��|��flfˉN��fS����{%��,:�3�+�\�{��a�x��My�W��#�w��g��4�p���g|�Z��֥ "gY0,���Q�)6%���i�)ϯ,�7�[�fG���V�⌔�_���S��\�����=!Ӊ�X5�W��@���t�`�G�!�8�x#��4�\T'&��}�Ĵ����	���b�9�s0��z媴�����_�-����S�a�#���������j�=Z7#r3/(�<[YH%��O��]�4�[����
��d��&�u�=��$�v4��g��7�_������0�u�r�Vj,�G����J�=��c�cP�ޕة���(�����Ћ׊)h�e���<¢�7ׄd�l�s�e�$A5܍[5�X�Ȥ�?�zi0��H�)�xG�:I���@(`���k1��N��_֊R[��� �]�vk@�F��Y?�_��[LĢ����Cl�	�њ~�%��A�'�I��&M6�?�	�.���Ϣ��?�����q�s}�:�W˨ V�@��2*,�̕ML#�"S��M�C�Y1V}�A�4˫�~h�R\�"�"\j�<)��rB�!?�d����W;����p�s�������Z/�&Ë��5S�~ܗ����I�x�������[��/����W�숞r�}-� ���0�ۆ��nDf���ϣ_��=�߯}���䛆�8X�2u��B1��5>�z���_�stI!�sN&E��4c����1�1��.꽚y��@�X9EO|��9Ř���{"T�uC��nrM��"��R�oD�DF�A��^R��*��Yi�9%�PTB;p��	�n	����n5d3���gT2$�-3C̈́>���O*�(T5t�F{���D�_[�p�L~��*�x5��~��ג���aUd2��0��i~��y}����"0}4i��X��_�@�T�����S�a�t�����|��?�F�c��k0>mpDb
�_	���U9�4j6�̭3P0����������%��ht@�r�N�Ϗg�-K��I=�g��/����'�j�R��N��(a_�Z����+kn��1I���ϕ��� jX�G��q�2�:���6/��xN��9�C�S�ut>�'Eb�H�~�gfM�φ��f���8Z6m�or%�2m�yr5����g����8Cyz�������t��3x�\�!k��m�&�Y�Չ�'p~�G�>?f�v�o#�54�_�J�s�n>J<��`�r�7�7$y�ZE_υ�O� .��qu7���G�G��
�z��Ѱ��
���6��i�$�m���1�=]_�g���yf5v:+��%���Oq�z��M��H��s����R��^7�q[��L�F���+����2��q��H��+��UM�ghp� 6�� 5y�2M��Z����/�m��k�U�#��K�(�"nޓ��b>j͡�6�x+;�R�Խ��<̏&�P����%�ʇb壯p���[�S����IF�bk6�,�����u3x��S��x��p�r혀91K�N>���;~W2;T�w�V[=�܌}of>H�Zܮ����i���p��%��_��<�����4�T����?sP��
�*̘�B��f���rU�2mC���h�X�RiT���Ľ �(s��?�����cEg(�i� sn���Ba����u55Z�(AEf�r�Ưq}1��z꒧p�x��1v�
dn���T�e[���i��1�L�k0uɺ��!:�	|�{j@�J�E�s'���d�����M��|�$�����t^I(�M#%"�Q��v�39��%K�QH`���ʷÑ;\@ 	�$j1��a�I'��uS�4��qE��f��ޗ炐�$W�����P����-"҂�Ys�]�T��8"0w���� _'I�*2/`��ׁz��*���3ڴ ���m��غH�Ł��E4��%O���TN��B��)�y<C����H\D�1k/���R?z���'��т�/,�{�`௖fdMT�oA�������P����a��Ї|�#'1!��d�ag:���� �U�N�n]�n��OE܄��5P7�P=�G�J�������*�2xf���J>w�{B��\<ڑ���������V�:�J1���pz�ri��p�8@�P	���*�];]?`�&�x��ROk�RM�R��\C�3���_<Q�y M���Ro����̯�H�_NTR�X��zE-h�&�8��Um��X��5F�����Ly��\%��Mn:M�G�	 �Q��?�d� �_."�JWA�e������jg����6�%��I8�)r���� ȶE`ĸu���ýz�	�^�B�?2u��z��oؑ�n�#.c��<��"*���|�}�zJ[�׌��^s`"�9�:�#�L�u��Z���#�y�i�� UU��V[=(;�&��P��?́���\�G���a�tC��v�@�a�7r�Sǆ8|ϑ����X�D�8Uf��uCWnZ�S�ҧ*&�fO��8Y�0 [�3Y��Ӗߊ@2�/^��3�:.���7�}���a�	�33q��}@P�ue�k��S��悂�),e���hl�~�������c�ѹ������]�"��]�n���l��A �|�͸���¡[gÕd�İ�$�7T����(#�2kR!3�H�����Yc�( I��_!	h�tH*�b��@�<��b���U� �8�ff:"�d�M�:p\�[q��XvJ84Ye��Մ�␬��8��2��!Si(
��=F�\'��O^�%����6^�����!c�M�ۚ K�s�`Q[T��@b��b���gT@�4�� ����#"La^�O㢀u:��wxn?�e�/x/6sP���sĉTG�s"�a �,��!�̿��7|8Pw�a3�K>�-��o�/e���4�@�wՖM��#�Ԩ��`�Vc��)���%|��=��AC�[��)E��8Y�������v���x�A��JczmU;}��ob"�?�-,��OJI�SRC��5����Dyp~�-늃�)#^ԠV4�Q`D$2���gvV���l�]��0<��G�y�#�v�G���ޛ���ވ�	8����ק?|�.�E��~���{�/Ţ��ֲR��]���
��g�DF��Dˮ��V�^��ӹ YY^���������:�>�h��Vec��'�`��UP/(=��'���iU��P�u7Mj5����ߧ���N��l�1��dV�P(�K�{�Ѐ�=��
��V�[Ģ�Ԋc�#��L~~���r���IKZ7t�c�\�T�Y`�~1���V<j��`�+�7&��r��l���?(��v�qX
1{�>���1!����7��u����x���Y�b�_���X�*:�`~�����"I��P�AX���r��ƭ-���>~S�/M���	�~�z��j��,�D$OQ6�"?� �����gFY�Ÿ�W�^:�`3
��ŔM� x)��wn���USLV��vߒ������/�Ni7���!�VvO5�J�� ����)�5㛝�^�Z�#�v�������~��Y=�Ww�%Gzr&�_�2�����v"�]Weǧ��i녩N���*�ƾf/�yf	8np���f*�e�˴ۘ�U�}ѷ5�&&��u�Qw�7(1pj�|,�%8'��t�a`��+�MF]	e�1�)L|�6�ԄY���~��_9N�������7[�A��a��k��gW��g8�(E�^�k,-��e�3�(F\�
���%��ꏹ��Ҁrag.�
l�]�	ַw3_�L���N�񸂢�����Y�;ԫ�V�U?NE�A������s/9�� �K�sG�)؃���[$�֥�vg��?�����]R_h�Ͱ��$�6Ӂ:צTb��������r�.;B��1�I���BR)y)u{���+!���	��pH�0q�����pcc*X���J���S�7�M$�Pf���Y'ł�QvE少X��w�<s��ی�����Vܼoߺ����3��i|��>��B;�,U�� �w��߯V�>GZ*ȵ�"���;Ijw8�W]�X��V@|\h�_hv�^;�L�f��)�U{�%i�śRD�~���-�j*��|���W�Rgx��w胦�w0����'{زtv}�Ql���/����?�	�̹�t��7fj��褔z�B ���%�
�k�O*&�fA�6C��Q�MN�����F4�[+��J��e�g��Z�g������yg������� �G��$,�W_1v��a��AU�i����/έ�Ks�9�4$9W��)}��4����B�ԡ=ClL��ٯ���n�w{5���]F�~[*�>(g���cl��=��7͖O���^GL
�*�F�y����a/ǰ/�R̭��,iډl%�Y9����`�DwCh����e/�בߦ6����6׊�I�*����x�+��}���r!q��<����t�{
����T�w	w�瀼��q|h�z�Qsm	��%�Lh�"�?�m���1W��͠8Ѧ��dc[9�n�4���VsDB�.=���~��g��%E����,�	P����4��b0��1��3=1j�]":���f�@��\H��'�Z�b�a�NU���8DB�Np>C��o]�>��uJq��"�c� Hn�Q!��'�6wD���n(�Ըj�J>�y&`����$���J2P�	����C�B~q�R���{,��Ϧxx�d]3��{��E~d���]��$��c!��V�i����o�F+.����m��B/E�ۢ��b保KE�����M����I7*�;H���K�|D���/Nזn�!k?�L�����y�9фLTS���
`1�Ŵ�3�����9�v�� ��m(����}����?��C�1�������3�_��jոY׉Cbr�����n)���C�3:3k�y#̻�8�S�5.[��^e��͔��:VJ�X4R���__껹�0�!��g�'x��ӽ��؜Ik����*��i�C�d39�!�@�)��-���9�2��"�r�JƘ4H鈟�U�uʻ�I�u���ƈ$4�*%�jn��O�ߛ��^l�*]�l���:�i���6
��D��chI�v��)�  ��hb���Z/l \�*�A�E�ߔjS&��?��@+�R��n��b�"�
��m��,=;��t�{����N��;�[������
)z�%F���4���� #��rC�#b�<"�Y��t�X�Z��Sn��aK�J��)�#x�q�
��ho�ҩ
����Q�}�:���a��n��w`� ��i�ܙ�dM�*��_q ��\��`��Le�9%�hd���f*.7QRs�!O
1SX���]�T}.��[u�x���T��2|ھ�v�HŶUƨ��,�*�|#z��_͊�� ��Ͻ=w-i���hH�<Y�к��������j_ق3��Ȧ�/������I'(�c��I��F���0>�ȁ��͖@�良�ۣ�alT�Pd!.?*3�dss"����Ь� �,ub�̟���;�� >��DH�3A��Y����)����F�B��a�-*���BI���-ME���������QZⱥf������7}k@��y?�˷5P�j2�� �j�(��~{�cToA���E�p��ԫUQa��៽��u
�V�Oj�iT��Jb�B�!���m���~	���DH���8�K�����
}2ލ�Qߢqk�o:��R���x�����5ݴ�93����n:��@K�圄 ���;�]�ޘK(�J�dE�Ԯ��ضU�K�b�}
@%����V�g/VjQ�������|�tJ�˻�JWE�Қӑ�H���0��6�洎]��Lrd�Hzb�͇�9���̺��}y�Oǩ"|�d�*ZP�=Q���n�:�L8.�j�����U�r��Zs�@�򛚘���: �%�&�tU-��4�##����)x�$Z���ʇ2 �S�!�`��c��� s�{$W�F��8��B͚ZE���gvS��CW��.}&4j��q%���&8��T\
O��F�B܆K�7C�ESQ��,��ő�ZA\���7�M��ʟLu��<��Z�2�UѕJ��J��sP�t�9�-e$I@���@���l$��1.��,��S���g���%1����x�r�I�#���'O�h�c,�`�c�
���%E0��\���~�W�旧���m�F�\k�L���6���!��50����g>$bh��S���nΛg�S���Cx��U;|��(!�%���{����J��b�<z�᝿;!�E
�4��R�=l��t.r �-p�Wuv�7�$��,�p�};�Ny�#��	.���J&��wk=��%��:WQ�q!@�:���/�l�0Nnк^@��^u�4����D�L��.�&�Ȟ�|݀�&�F(`01@���O�#���Sa�*���m�h�<$�|.��Bfa��|�(��FQ�8m$[̀��p�e��q��g�f~^���6I��h���� �դ�~4���Ɯ�(���Y�AQ�X{n�&6D�
�p�
s� )f���#å9��`b���%������D?i`��L��q�=5I��<FuaB��ձ)1 oڎ C?IǱ�`�A�}w�+Eڰ`ŪA��.�W/���;���.W�����kOv4T@�yZ��v�C�ID^�4l;�k��1s`~�����}!�u|Q�aO�x���|�)�\9��{I ��J״ݩS�ŷXǙv���#<:=��ԢG	��@�*K��,�ye�j-�u���d)p�F��E9����q�v�6Ջ/�6{��?)�9@OE0��Yx&�>@ΰ *�QT�"̑��Of�2@�",�~���[͔��Jb��Zy&����N�4��?j;�� 0�U�tοX�)+/��%�uGX<��^,�g�< �c}�J���_Hȉ�*C�ޣ�"��ʞ�0O��4d�����dHj|�����SPn`�=��F.������B@t���d�D���s�[�荖"���^��v�π��gv}EPe)��3������d�D�z�}W�5�{���_0�����,�H���6"6����2f����3� �ܲ>�j�Ӽjd5y\U�
=��Q�����+�����B	Y��$&q1`%�*ߐ)SY��Y��	h�Y u>�r}�\���")��6����l��_��q�eM�����j�g��.Mtk��0?B)c+�y0xw�{ 3�B@�wW���*)����-�.�Ӳ��ޭ}��Y�f�E�����Þ�l�bD�?q-�	��_t�㢏�Sl��ճ(��с�gƻ@��
eDhj�_˝g����z�sU�Y#Y,P:Pv�oNq�,l$@��0���1hD~�0��u���՗���o��������)�2o9�i3&�0x�Zs�D	��l�7-!W�jMe�IM#��,d���\X�'�eOO���F�}+f���\��1�T���d���|���
��JS�E2�e�U�QB5	��`�we�2ڥ�����%)�!�gɕ�"��mtP�ٛ*�V�OkC�Z��(���5�Ɗ�D;��3��A�k�=��]k1F����ji���5MK=or-�_�Z�n�����MX�5�|vk���!�ߟ��m���!'qzy��P!{�i?�=�ݦ̢�k�ې�����<=��?Z3�%�&:'z�M�Y.b��!"J��ѯ�S�X�e� ��d��mH��K�!� 5؊��`��
n>9���D[�#�wf�#E�j	r��W"<^c�\�fz���<f!9���Όb#���p�[�j�����v��ON�a�����Vf�x���L�Dc˃(v+��N��?O��L�؉������:��}�"b4�ޝ��@1]����������$|��m8��.OA�5x�B,�mO�� j�ӴoM
��Zq�믔��z�,9c/p�^��	�Z��Ҝ+g�:����.�����C�ki��׍��5�	�8~d�ۇdt�V�E��=F��HJ�+��i�j����0�Kޤ��&���"K���8V�����G�˘�� Թ�h��uW�.�D+�}�z��șK�(��-Um�Ү��X^�.�>j�t�-�͛U�<�1� ����p2l�U����z���1T��R~�b�Q*B-_��än�s�ޝC����dTgV���y����IJ�U��tЄE|I���L��\&����F��@ޢH��!(v����A[�wab��$
�~��O>W��*`��þ�dǼn=��Wy��p,y�ZV�N�=�ߒRQy��zIe�2Q�ZHC#I�}TE���$�i՜v�$�4u'�C:�,��; 	=�S�㫙J�� ��w&���Rчc���5��4FW�/(w��gY<=��R ��t��0��4������NF��P�L9E$־��l�gZ�����n�u�ʡ�u�|�Ap=D���Vy\*v�#P���W��Q�L ֟�����G͍gPD^�CM�� �����a~.�z#��'��E�	5���1(|;�'ƕ<|2�ڗR�j��T��S� '��
x~~ޱ�w�6�|
t�<ґ_�KZ����6�Q�(m�%h3�S0���U�`�%�T���T\���:�3�Ri6�����J�@;pVEC8Kl@.;��֐9��#��K�rEM��;��,��$�\��U��W?��RѴH#�3��n?�B�?��Z;�����>�'j�>O��QPS۪����w;���e��'��vT�@BdY���c0��ju��g��!<$�xҋ�ky޽�|,7k�\��צ��G�����+]N�m^�<�'�o�,�*j��Ǆ�<�)@�2���p�����GKnԼ�Gi5jγ��ܧ|���p��LS�=�=t�1b�v��TBx���-)I�Z�il3�j���c��t[p@�H�ȏ���"*a�[|��3��y¨;�Ji_�fP�L��Eh#Cxd�n�ll�
f�%t<Z~
4�]כ1PЊy1h�s�!���	s��|ČZ~>�<���2��E�t	�q�p�,�&���ȟD8���,�3�j.���?��n���*�ԲL����'jF%f}�LŨm^+�CȥW���Z����[�'͍�,��jI�qސ�N����/UY&S������SB<�K(c���l����N�.�z��m�S�!�vF��'�4B���EX,�Ѵ��6���S;?��&�S�+���Ke��q���ͳ��}�CѸ~�q� �?�L4��"}���U��sַ��WP�\�\gҹ~3�}�M��@���Զ����C�J���}C�v�[>�=u(�3<��c����r�� r�A�X��]��S#�:Jt��H{�"�M�ѓ�tS#�0(k)���eUR"	?�\N���of|��+��D1Y��<��.�!�'m-׏�@ٌ��/�T�����_Ej��Z�����/��>�P1��`�Q��N�`x�듊Q����(-�=\2�\�0;ۄ�兏O�;�+���֘
"��HN��0q��䀘+�[���b��y�3IP�����u��#�"��Y�7���9�@W/�|��Q�_���O�[�Ee4��L� ���@��x]4�y^�o��be�a_��0���ۊײcD2Xg���9�6G�V�1�P�FeŻ������(yo'1-Cʗ��&n�yc���BP�A�{��G���C�h���"֩,�,�?�4?gS��"�r���w��ڒ�����P'��F����uI��bG��J�M���+��GV�dP�p����p,ՏF��.m|u�/=|���iR�L�?�]����㲆��U�hZw�5?=��F�Q���u�~f9�B����:OV��r9)bEk���/۱3cM�����B7[��f�H^o>`������7.�E��}+� Epт:%,P��@W~R,��V���d/8�.�)�!��9�8Lt�Xnp���3�R�'�\j�U��X�B�2Mgg�����҃��t�񔤛('�QC�]l�z!�l�M̧8	������`:tI�F/�lm�+���8��qc٩�d���ݩ|�3O7��ok%e���#��ce-��;��ɀ�W�arg�Μ���Guհ���?i��r&�dPpm@�Ԕ�a�������ne���Czn׃�a��@F(�<D��	�t���G���o�s����Eլy'�?����
��}e.����r<��6 `�9.{��n��*buf��0�XB� I���CqXwH�s�T���3˩��ǫ�(ӥY��Y�؇%@�Kz�^.���w1�w�x.;'������͜�[ �cq{|�"��M��/S���B�V�  T�걦��!�52T)��7	p$�o����_W��u�
�-�����:����*��t`�M��T.�b�A!$h�����A�AN�4�{� �1m�<g=� ���%0֋^bz�Xc�p�EҼ2�����=g3�I|��	I	��89]A�_��:L[A��F.���#fR-�k�\�G�M��>t:K&�����Jr�tW:�ʩ��&�+u�i��ޑ���DE�+�f6<��`͗�*^��B���}�(�����ʋҀNv�����'�V^�B��*-C��A����|+��u�a��Ln���i%p�7�f�x9��JP����q���'��e�����������+v��+{6!I� �tt����Z�4u��V�S�VԾt���3�F��BR%
����$$ ��^/�:�F4\\��c�4 ���|/�>�]�z���Sp�����aS�m�95;�~�ǘBڲ��<$���ـ�c��m /��O��6����1<,�;C���*�ś��`acvO� ��F�P�o�_��*��9S��#H��f�C�?%�<�1Ш;N�껕|E�γ�^s��D�u+�7p|a�z�'=oثL��ž/����������w�<�*����;�,��WCa�Ҙ�~R5q
9]����<���e�E�(���φ��t}����+�aw�5�!uMi&���vyeRq��GE��g���72�%8�A=@���<�/�0���@��*Pfq�b�]mHq"�D��F�o�R�{ZG��P8s��Q���*��I)
N1v�W��ui���۷7l������ҁ�@�	�yZT^���x`Pv>��i�Z��O���,Hn2�[8��\��#��u���+�P���Z�����n�����@P��)Kޘ<`�s�{�V��~O%N��?�-�x.���b0�R�a0E�=5���^ T�T�?;��U~���I����s?h�	z���mϜ>�@�����G�Pc�:��W�����\��l&��O����Dgaݐ�\U�a�F�ĸ�>�E�K&e�q�K�R�B�?mY���:a.���,����e���1�$֑��~���ܧp_C�}��,��ޠ^����P�P��I��Ke�O�W̺9�]�q�|�vZ� ��I��FI��_���-��X�t���\���S����H��w�5H&���R�6k��+�����(P��0����k�)DzuhTV�\�<���X���_K��^����s�TۤC�C���;�:�д��2��q� �C�;�����J_�\&��檩���wҶ����#&��)[)	T����u68��D�Z��-�_tH�p����
nh��v{��P`^��<V��}�7��|-�vԋ`?�~�����S��B"���$<fU���~�y�G�௄-t�]%��˼n��km,!0e,��w�I"���Z��<s�-�E������b�舃�Ţu��j�>���p�q��Y�!�C$	B�0���q*���D]/�n�+ڊ��+��E֘�u�8U�!�ɿBCWo� ۑ^�㙲���5[&�B�Q�W\M�+�lek[��v�mnIm!�A��cЖ�����[�ե�-47j�^���Pt��E��Fr|���FBo!䵖����gp���g$���v�.�٘�˕A[5k�����Я	�H��_)6�y�B�iH������}�M��������A�Q��#[�ۢ�r�/a��A?=$�l~�����?�E�T�8�@�ݼ[x|{S����;����a�o�:JF�;C||�O �]|f�wۨ�	,4>���M>�Ә }Cm���z��R͡7�:��S֋|���hh
)bfZ�=|eVJ��|�~[�)K!ڍ�G���E&��� v~�S?�Pa\�F��e��\d�[Alș<σ��=#�[qQ��[op[�����w����4TMI��688��tf�p�Xjͺ��w��KR�!+s�_4�	t�ê N�X�^ԩ��x��L�s?��6��Ȏ\�{W�&��$E�b�ك����)?z�]�f�4<'�uɌzIK���: S�-P��(�y��h/n[w��a�C�2��j�m��WqQ���s"�+�o�+�цx>�_U���1x����ۥ���M��F����Fe�ĉ����>��f.�!PE��H��*(-���[8Y@cl:��]=?B�܀'��gF	*���}�L�݅��;�O�m�ºՁ��6�z�N��# +��?�� �-��낤��Fe�I�ut��8O���r);zq��@�Ӹ1"��w]�9���5�v������ߥ�@��#�8�EZiɝ�kl-��m����~F�-	a����AH���ȋ@��`�}��p�j�\J3�4�r����-	g�G���s=R��]�{��"p�¬Q"&�l��F5�艽-p?����CT��T�����>�6�
Z��6�w
.�^���w�ȱV*�@���,���7d��N(��`i��Iz��N�Z �se�hAĮ���Jc3Yֶ����VB��sʡ��qZe���{���q�J
;��Y-w���s�� �Q�ޚ�� ��dX6��8�ۘ���靯v���w����`�I�����%���t�V)�ؗBG���!j�s�|������%q��wa�$�u���<
-�(R۱KV�A��=�$Y@s6�,, �١��@��E�����[A���eΊh0ǰ����| ��^�n7�#�O W�A�ƺ�*��d-����a����&�E��a>[⛓�Zg��1���[��}�	��/3��&>G�����!���%L1�G��2�l��/
/+`�N)�D��c���z���8cQY7���D5�����¥2T���0@��3Xv=_v�M4v�xq���% ��	<UϹ5o*mR�cϨ$��%0jg��2o`�RK�����̉s] �Y6J�qȿ�Zk��@�1}�:��$SY���u�*i7Q��9\�g�3�5�yUv*�"Z�����a�^��4���'�;��"�v���r����]f��j�;������ۙ�w�R�B�V�dI��+p�[���6�~�-�ME�`K,�s�/�R�`s�\귇�>��� ���FZ:��(�h
FM�\Q�-�Lڛ b�� �)Q�OAF�i`)�-2�\�1��5)T,�N}x�Ă��b�{���.���?�x��q;`e�(8a�
S����	:3�����j2$�H������ǗS���y�̶~��O�h�e�+ ���]Bܭ`������d��)�]6t�1�R��=�?���_kk�ö/�Ú�J�^�����/ ��p�7O�盕���o:���ȁD��B
��\W�Y,ۗ�?���M���#��W�'XD;g�Z���@����f�I�(��;�J��qqI�R��GL���ұLjs�n�C����-���@0Jpq2�?�x�%���u�Q��u�g��Z�D�ēIب(��4l�N4�FR�[�Q2vu��{�ۜ׭ɥ���ϥ��>`���7�'�k=��f"�hCbE�&)c�*`n���@D�1:f{v}\���]X��%�P*�s��[ ����++�Q�X(�[��V�^p�4`��R\ik�B{���U~��J�MI���O��_�Hꂓ)k͟1+��N����إю�Z���b9����9�I�����O�����H��Fj��V���7;w�]���N"�ux��a�Kv;8r��T��<w��7�b%9p>Sj�$rF�Љj�-����Z��Ԫ�����$щ+y���8��J��sXbEY�F�}��ww�N�2�S�a��W�x��R� ����)�i��AE�=?�i���1�����C��wr!��8/T��O�����S�p�F�LP䱋���q���g۫�8�HF�3qPS��*����_}z���E�%oV��?yVJ��e`��h���U ��tIm�q�Hq)m��ދj��w�J�	�8�q\UH������:;�	ҭ13±���K xgZe�;�:i6OSW�1�x�(�����9x�5�_���yΗߡ	tn_��c)碉l�4�� ���o�Z@@�:�ЕsC	��$�[V��<΅��y�	O����yY�^]�����V�+�[����ϱ�����"��.��3�{.��ܥp� J������]�٘�<hN�Y�ã�d�a��B�suV��K�o��\���I]f=%�1�C����r9��̡����Qu*]P�AVw�+�x�j��|M�/��nz$��3�r4L`]��4/�� �|�������ѣ @�Q)�i�s%{@E����h{5c��b�L<�c$=d��,��a
��U7�%	`�^�ym�c|�闾M�[�Wrcw��H�r>�)�S�l��n��2����ص�c�3"a�$iq��'
M��瞛*7�b���V���x��zx~�}��9�˓8/n_�֮ZE/Uᤜ��A��P���b3Ь�;��k�&o}�QAaX�|��%o��Kk_�(1�+c`](��
�۶����v-�x4�Ĭ�R�|������X����4y4_�p}��O�H6�°���uRt�=�=��v���^š��#B��{��y�<�z�L�eU�^�k<����'��k�0H�kն0�
o��&�����܄�v���ȟ8P+���Qi/�Ŀ��E@q�MPe憊Gk��u�62�L�dy*�ѹ,aa47���*aצ��d0������3B{�N@��G�S=��oq�C��4mR��z5-����i�Ȥo��2��ar���ne�Z�Ș�
�H���Qk�aǑ��Uov��2��~p�_��"Q��=5�B8�����Y��Η� V��N�E����8��q߬��}���P�\��\b�X��Tu�ܗO��� )�A�.$���:������.>1L)�R�XeD��	�B|5�i	���6�%a���a)0��^ɚK��nR�92?�7O�I�W��@���6�vzF8qDrŵ�����w�1�#�g:y���z��d�O�M:0h�e~��/���4�0���[=/ޅy���ѓ�t#�^���l���;�w�x�+��8�ٮz H:vb��3ύ�r��s�}0��Ɣ��\Ok�U,ۢ'̟%l�[M[ScQ�*�i�{i�}M��<D*H�4i��6�Qˬ幜�����@�S�*E��b��n��-mwmc���KJs��T�� ȥ�*JA�^T܃����C8�|Yc�bf���ք�uǜ�߿��sV�F��	�,�~����-��F���,%=O�"_!���O���� ���w7!�)Bئ���`��i�>�mK�1�X^���Gz/��2�n��L�-5H�%��hJ�$��|����/L�u���Nġ3�M�$R��U&�l~-�Eo?��咳�-
i7}#���?g�`��D�/��o���" ��������'��*�xm*_�Vj&}���s��z����f^��x�\d�,A��Q	au9ќ�4 -��l5 akr�83�d!�֭��oU����=�&�ƕ&B��neP7��C�H���3� ��D
�ҩ%ކ��2ֶ]^Y�i<G�I����Sc�bk��m����h��
ܖ�W��{��ҐrL�ƞ$>�W�f��#�F)�|�˩
zN�(����g3-G�Tt��%������<"�����ϋ�50���^��+�(���W������sӣ�;�Mw,na�� s�v�њ����fB~ܥ p�f.x��w����X�
��z!�*
6��ǈ����7��V�2�߸��[M
;���0�K�r�$6Xc�F�F��E5��:}`�s�s"�aa�TݯBR�7뭠�]0����>��oIfKCQׅ����8ܲ����;�6N��W�S�c��9N=�l
�9Q�j�:��8��9��h�7�b$���H5l`B~L�4_Y|)���y���['~���7ʓ�[o�:r������|<�3^��9m����[?0YM�Ƭ�"6��� B�$OqBy�KZr�ݽMB'^��:%L�'�:���{}�U��JP�v{ܢã���:�m�!^��,y޿$s���2�K����sq�� ���%7��i^�4X��jI��yD�+�U2���m/i��XI�T��iЁ(����z�y��x��#ֲ�� ����'�INNd=(dG��jC�c>�v�q��-������H��o���Ɵ&�%H�w�2ah��3ع/�"�<l��<s������%\,�K�{f�0��،v� ����zi�����A}W��)� "Qc� ��QZ\��Ή��ܒ{6!���!qD�W/ؘ�)a�����uP�W��U~�e��mY� ���$����q՚h�%[3�����H�u|�7aH�P_�y''�\�4>^y��F�!I��?�}Pt�TϏڗ'�[8V_5Y���N8 j����|�9�Ad�,~�F��+qp�i#M+���1�=��=�VH\��G�����Ƅ���}K��J����\ZP�6�T9�qN-�1���Y@W�?�&W{��?8Y�m��<�w�FY���b��� �,��rh��toWE~��%��6��MLa5�|�߄�t����B��`���3p�=��ղN+5mEZ��.ݹ	>S �9^�ͧREil�Ӊ�S���7�h9�����58î<y"^�Ozݏ�����/�pTW{��)����ؐ+94�d���9�&@��8��Z��0��Kx �7LA��b��+`!�s�rP7�D�^��:�D�U�6�ߦ�;�tF$�`��ç��1�)�p�����>���H,s�`x�q�ny<�����yޟ��T�i �`��\4Q�Țpy�n�>���zP� ��i:^Lmt���J�XY���(/vd���@n���ْ�g:�sj�0��"J�5 �;X>s����w�#��o�1�zx�
��615"*Y��i��w�S����
�6�=��)#�������l�΍ӳot��U��:���#�%ڊ��{@x_-U���Zxt����;M�k��*�;�����Wa��������D�#.�)W�Z���E� V܆��+�\xB\\0�X�����CG!NNV���p1h��XZ��,fBd4�a&w(�@��ӳx�bҽ�%���n�k6�0��6�l0���Pai�^������]�hbxE(��xi$ƌp�n��JWy~���-����ȶ�
��Y�je���D�s�jt1m�~�Nш����J�<�;�As/x�rgi�Ũ_"�E�;�&4��5y�>��=�ĥ�$��a�s\�_�`ѶE�б>y�0*��5�ߏ�s[/g�謭�O��LVG��ZQ|/ԡ�߱�����M��������V�r�+��g��R�_at}��'�n�]k��dh���] ���D�����!0�_�8ར��
���&}_h	Y����&{^�b��~��;��]����g��5�+��]t��Z��D�`�����u�*�_��yk��f�{�UY4.�@@3r�\�/h�ʡ�QYh� �m��O���$l��5��댴f�ۉ�w�a���W����e	�n��H��  q-�eBe�2'J�
5[��m�����U�PR
�F�'Ll׳���]p?.Stx>j<�j�>l�O�s�j�q/5�E�r�
��B�G��M|�ۉ��t�x��)�UN���QZ�p�1��I�I�/�o���L�L&�X�5?,��B��i�d���zm�ӿ��rv��=��0�	��,���4���HrqۆӃ��3�H�~Za����8�q�+"��׍�� Y�S�?�4���u��.ã�>�_���=�d��ΰ�����)����<1���w�P��W*�tZ���ΉM�w��'f�bO�r��ϑ��1�L/�� d��&5G(|���IA٬���~j��$S,r�,D�/�{�����R^�����k�6��wb��
��& �]YF�%�w\��K���ԛ2��>x���W�Y�T�uϥSie/`����݃�5�0j�J�vJe��O����3c��T+P��M���@��<{��xP�X���Zm�!E醼j}B�Z������\���7e�XIU׶`�/Kl�;֒��`���*���Z���pL�&j�"��J0���U��pjG��>%B蔀R�3���ڵ�3AX�)$��t;E3/��i�!Zw������@mX'��zk�s"��>ܯ��ބ��������eB����.7�Tfb��Ǭ\~/.
1��@@G��R��y��j�Ik��C��J���c�Y��Ų'\d���ن�A��\>k�w�u�9���x�C��7�IV7�`���<�� ����먍c�a[	֎�,�̮k �EX!�+m��Zq����:Av`�x8ə���	y36���~�;G�b��Tbuaɮ:g��f���<I��U6��J��q1�ָ@G��ax*�E� iџP��������_�u<Hy�q/f����m�J��M�H�W"��,HR���A ��?!��|c�j@����b*�槨uMm��7_����"�_��])�ՙ3U';���h��-/��Ļo�eh�m�6�J��<%ѿ�'�X�=+C�<)�h�Z�1��O6�n��S���T���f��R�#��Yyؿ���0M 8H%�����$��"�B#�f4*\����J� �r���d��T�Dt��1���RȹM�E�tNB�HjQ�V!G�ȼ6�K ���M�83���̹�"���km�(�HN]�Impl�JL�3�����>�$�b� �
�z� d�2���?AB	_I�����S��Q��⪆�N���J.��,�q5���}�#����*F';�_�����xI,c�81{w�d�Q��;Y�p�����MH��/�M���Z���H�W�+�W@c�i�����7V"�?�P������r�c��R,����]�����a�AO�z��]����t���F5b#��,$K����@X��"3���H��m���P��P&�bns��5x��¾��Ixx�r4�9�̏<������?C��Y�%���=}����/Վe>X�����Q��Pp���s���7�'/�a�+T>�ϊ�-�%�0�4�4�ҧ�Ef�_��ki�ap����;��g�F���YF��/$�m(��Dyj��'�!Id���ܰ�51�/a)~��b)�CƓ�R׳�6��ÎKs�C1��^���=��f��ͨ�J��G9���D(]��%�g5�t�²�#e��NF���ϩ�y��k�������f8�U�[D�'��/)ק�Y�V��k��lV��;������X����RTBK���A�3��z�9�:�+�@��R��y]��?�f��Cu7J��y��u�M�r����%ڮ�Z�����u�Q����=	/��G�V.I�j�la�:Mܨq���
�Q��t�\�(�lJd�
@ɻ*�h9��̩��K�P�g^A�=.�&��yՃ�vl�:	�\۔����z�A�������	:A�,��k�����@':����<�L�LƠ�WwT
�$�+6ל���e���h��l�EK��Q�"�����4�b��\@ф����6�L������i�Pux�Ɋ1��/$D���o-'3G57].�L.�v���i�t�$�姱�/�F�����9ג"�p(�L��j�q�� �5��@��K�*�sc��p����8�eFvZ��-^��߁r##ΐY��o0���c�-0�j�{�3�e����z�e��6o��G��	i��3N٣FL�(7Y���yU5n"K�ƭͰt@����ǴI��H~񳼪z�7��y%жɋ<h
/��$��d��s���Cd��A@w�@����]�B�!@L�脪�$��N����U�/0c��d�W0i 2�"4�������x3��\A��SB�)�+��~b�T�����m�3Y�$��}�+r��r�v:̃Y�F ï=�8C���$6^���r�8��A%4E�$�P�0���N!sg�ln�{F9���0H���(O xc�RD��|�ػ�ŢG��i��9�q�K^w�B��"���A����J���/V�k�d,"�(�x��ꯝ6��W�`|jb�N�	Hq��積�F���{����F��n�d���5#���e�ңZ�L�M���t$�I�h��ǒ:�LZ����:�T���`�0��E�|�����,P�s��)��b���3m�)�Ozf�������z�zuԨ��=@鎾�͋�D�2:v�i9�x1벋f��1�<����y�j,����9=	18�$����
C��J��w��~o��d�:=mu�{��R�{#*:D�m���R}nb��73�~g0t��m.���|L��~�r�4LV����Km����8���|�j0��D��+�sÀ��ǉ �$�Ʀkb�"�%T�r{��8ئ�����{��b,&G����y����i=o7@�8���T�{"�Q�	M�r��HI������ga=�QE���43�-�]����Y�
����r'�3Ȳ��2��\����nA��D�`��D��#��66�j����M�Ǆ��|�q����乶���ϕ�
,�� �$����M
�H������~��)ޣ�����i)����*�-v4�W�2�P�Dx���L�H�8���	LЗ���]�A,{��a=����~����%���u�7���0\����{%��I�=N&�G�Cz�����=8b��YN�\�/�~�*��VW�A<������ o��.'��F�>3)�h�}k��Z1��9�n�DA�����k�L���s���E�%�nH	6[���Rh�c��j�d��<�l��0V̼���"g[?��~���>j �W�H�2J�p� ��&�I	���q�{7����M���P�R�3�XL!'ɰ���w���/.J���&�����Q`m-T�`Px��+�~՚�YU�V��n�N��������?Jo{�i�Fܠf_\S��
p񝌵�{gJ��1g�)�QXi�B�:�M�n��k�+�8�x���P1Q��Y�on�s?�⊡(�;�I�Y�l!��s�>�#V_@�Q ��NN�\�Ҁ�Q6��1 򄀈�M�o(S���a�ʟh��l5ܞ��Ɏ{֩�����@�)�H+�c�$
��q��/�ViɆ�'6�H}7�r_ٺ~��a��#��L�N�U�ӔiCe���������/�8� [2	e��VL�r�I l|$$3�M����4?�ho�1B�P�˒T;6n?�_Ӷ�z��\��<|;�������Ѽ�O�c�������W���#����QM�
�t(�vfr3N�M��§Eߩ���؛� q�@�������M������`IE=�vA:0z%S�q^��NZ������;�[�p��^朴�S�����^#o�}i��pb�ö,�l����dc�'S}��ȇ��ޢ�����z�����z�����q�� ������7�,�@�2�@A�Ͱd���l�� Lu��Ŕ����"�̭`�v�s�J;�|��Շ����x?�j���ؑ��/��P�eo�����d�i��O���+�H~��w\1�x��X�-4R5��6h���(ygE{�׀1�w_:� ��d-����%�
�8�uwо r��SSƀ=~U`�t�x�<��@��(יٸdJ����p�~�cc�n��;���{(�J�',�/J{� \�M/"���	X�$w�����!th�"kV���� ����¤/仸��A�z΀�i��q����:����xa�l����3^�#Gp6"�ؒ�Fϸ��>��״l�Հ�x�M�L�L#f�:r���������'�
��+_�5�PdI`/U��sor�����H;R2-/2z��� �N��-��?�����k�����Z $�:tUe���W ���}�B*�⡎^^�@'�d�����&.
X���LT�j��WKLkp_�0�rc��M�s��ۑ�w�jC�όDRR�+�\�7@��-��&�d�P?W���?/�������\(��1��Kt���-\�%����i�7��@E�<F�*��y���+��42���b%�6�}���.�/��`�r�h������q�̘������5!D���r����(���fʨ)���m���aC���^Y\�7@*�����%�@���;J�fd��pr��5�1}d7B�XR�Vj;��$l��<�s����怔�0�$����4h$a����=K�jH�� �^��:!Z�Q��1��Ƈ��pF���I3I{6Yztw��V�]��;��&u9��
/F!��$������@+�њ0�\��J�l�fa�-bm3}J0�m���+�滌J�o��	X��0�?j�/G��8���p���ze��Be7m*cp�g]h�>����\�7����m�C���$��ɚ�W�v%��O_ � <N�
� N�&h(�madߓ�u��R��I�ON!�������Cv!��e�1|��
R����we���y]��U$d]�	t<�P�W1�;r��Q}p�Kɘ����n?��,°�v����,j��O5�x['�G��q'���d'��9%��Y�>7���k�#8�� �l%E:E?sA��'A0�G�J���'�i|PW�2:���x��ߘH�}�X��cĜS(�4⵵�44�k��4�_kk��!���X<J���=dn�����5�QLz �.��T�]�W۟bQa��}/�7NbGF�Aa��a�anɃr��Ǭ��O/�����eg�`4!��ǶI�`�D���8fs�f��t��]���@A�@õ�T�!����9� �v�דIX��ƻgw�����P�@kR��<��qC�8#0�b3ބ���Sۜo�=�p)Pr��U�v�Lf�Π�2���B�U��r��.�`\���,��~��~��ڝ���ǵt΀O01* Y�d���m��p Y��V}�������A#>��ߛC��Mm���z��1=�2�U�`CHЙl���L~�I���-lǜOUeyj���zx�L�~G�|�ԭ����dY�KMt�+f�6��.�$�k� \R�4��,_�T#.��z��m�G\W~�5���K7"Y��uT���o�aס�N+NuK�?SlV�<��yb�N9ԯ`���ռ(�KU��,gx���Z����T�Y<��d]]�~���1�I9+��֌���8[3�����Ŋ�R�D�b}(9�ΜA��E5�5
��ڼ2^��%�lG�t����ae.f�NFD�V������R���Afj�I���{����Dz��R`� �z����]���P6t@KY$b�|�X�w�Z�zB�D�2w�i�JZ�C9,��&ºi�B�_�
�4wrj�k �wΩi��
OA�*�1N"W�^}l��4��A��p�1\�A[��T}��\7�4-��c��P�W�2��q���.�vd�o�VnOD�bS��0���"q/5Ϥ?�}�)z5V�3�ڃ��·ʴ}%z�9A�ǔ�������k���� q"O)R�mߣ�VK��id�ș���
Hj�	���QD����hJ�6�ď�Jn�p�?���C����\�n���lO�Z%�1���{����+� \.�>T���������f��v���{F^�V��ժ��/ I����g<��+�������&HO���]. 2�S�ki~#`���U�qm�hm@�]��}5�.	�n��7Z4�SnJn�A�l��4�V�z"`���>����N�D{��z0D���<�e���$%3.���l�I���6���G���;syVkEh��吁�%A�s���9kS7�t�`H@ĵ	.��~�(/0���3(��Wa�{�,��w"��p�]'����7^f��o�B-��|�8�!IM1W%^�1'����Pk?t��\}�������CNK��e��ɷo\��/,��å�G�Ȟ�z���~}3�g���!4��<q����*��������ȡ�$̚��DF�����%���6n�l=N�V�"d�����ZV�2(L�<a�!�HR��E��c���������bW �X�b��ް>�)?�l��3*ֻ���sm ke�$�	sK���6b�**|�űD �b�����C�ϮݞʿE�%B��"�_��wkhd-IE�	��)�q8߱/G�!(.��Yl�+܄��n�+!d��2�rlcÛ�a*#8�N!`<��{J;�q�<���c��\Y����Vym���Q��|�w��.f=@��YvO��������Y�/WV�:P[s�GvD�j�n�[ø�|tpn��~ȳ���'�X�������;ݬb���`ti��&E���b{8.��R|����C�b�qJ� �a5��Z��˧yb?�&Ę�'`�<��|����Y��Z�a
�r$J�e��g5Yc���u�>��`�\n�S�{02`�x�F�n���>7�:a�Z�}�^��o�X� :����iœ,5�A�9i��n[�qDY�?�N�N:GS�1��i��y�µ�H�B��5���@�^�$��-P�m��2�!L������N0��W��.���V��Bc���7嗓.�N�n+XQǈ�E�)o�W%Qd�Z2�d���1�` �FK'\��ے}�0��S��'�um���U@%������&;��ٌ�ġ���,~�6���&���@�e;9,%o� l����H���ؠ{ #�.�I�0c>$���㡇Ɠ�^e�R~�e�D�P��'ݰ(���E�a��pG�f��
0*��ux��\�h9�A���&<[I�����+j6 ��Б�'�k"�D�&Ѧ�o6JŻ�+�X��W��-s���{EBߘ��U#}�,��*E��F���s����+�/� Y�:�0�
T�/�*��t������q�;$�}��z������z���:�_w�}��M�O��a{m��3{��0������%Eh�:9��G~|ѵ�`j�ˇ�#�l*F�v����E_���&?[���jn)�Z��w��)+�}�coN@��h���[�R%"x�:��L1V8{�Yt�6�n�;���h�Vݘ��+ݞ��g#����J9�z��m��<������ZH�oՓ@8�Z�`�,��H�X)̛Q���)��Be���Q�B���r��<�󩣪J�S�<
�5r������f՘@����Ҹ�%�8{�
��G
7>EUb�=Y/�-5zB#4���	a&�u�s��� �yt���}2G����h�5���MLW	%,&�[�k���:(��>�@�<��l:��n
	� ��sP`5
d6��������Z$�Z�t8��P�REp�?��p'j$�'D���y�ag�x�PZ2hX{�8���s��z��`������VX�)�d֍}IU&���Y�7���ȩ}��u3Ic0� �����+�w}����hx���s�$��Rh��Qb��u�M�'��3��(q	\⅊匵[�*sr�N�H`��PV��B�a�Z�D]Z8�劯 (��sT7}E���ʟ�PA	"���4W=%�`���ut���hx��\�[��2�s�pn �0��Yq��N��7?\���˶SqPk���m��s�ΙC�	�$O*гIe)x�v���hŕ ?�j_�	��ka�j%�H��%�|.��H�)RB���or2D�!w�!n�hq���N����*[zăQYN�G��������Ih���:=�k��'Z7�݊�����=���2��C�Ï��� Ӵ�S8�wCS�,pG�� ��F��q���f~���(��I�I���e��.�V�M߮������O2`���q���W���,�`a�m@,��TFNJ��{�޶�I�W�;�k�H$EH�Q����Z�i��N�y9��x��z��p7psN�ƹn_x�R��M�s��S�}�UOY���P'	80��\ ��*���e̤o��׬`W�JH��W�(�@�J�"E=�X�0Wb���y�B;�PX'�4T�((7�C���Ĝ���!*{@r���1ժ	Qc�`2�3*���-�4o����
,�����k]�Y��8ne��<�����\�ǻ)g+�dAK�&�h�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�C2��~��?f1ĭB�h������^��}��;����rPnE�CF��~��9���ؼ$aHh����k���������q�b9��'Op`�`�����שC�����/�5\�Z:>M���V�L��8�H2�7�f:��nl�F�2ǃ�K&����9�+���0��Чe^7!�E��#��t�HGf��58paw�<������H�@�N�I�t���X���ũ����7\�Z3̿��q�����3�kXs��a��t^2�=����@_cN����R�&(�!����KAV�ڙ!�=��Q�jm�1Mk�2UJ߯_�>�'rR��#��׈8́��z/z@z۪��p�Ȕ�R�1,= �w̹/z�{3Wأ�r챰kk�=�3��m��~�#����B��ŝ�V����"����E^ј����Ҙ��&�en�Y��*��U%-���A]2~Դl����܎٩u�¾�x���4��%��Đ4�Ѷ��f^*��I�
��Sב_�k=hn�a��1ʥ��I�o�'� �v��)\���[F��}��8��4F#Cn�6Ǚ�Q�Y��0�sJ,����g��Ҫiݨ�}�Zz\~�[��
�O�$�'~}�7x"�vwߴC��ލ��t�	9�$��q���,G7_��{�О�����`�b�p�OFr�������u�yW��=vVC�]]3GU
�����K��ZP��#�{P�z�5���_�ǏI(]�f�PmOKI��a���:��1�F�_R"�C��}��7��tSO��=��N��^��+�ָ��#4]u��:��S����)J"�.o�A��q��� \�t��l�jX��f���c,%�DE���kIvP:��Y�|��~�8Ƀ�,"im���"NR���KG?�-�[�H� ?��x��J�%-�D �$ﮐ�$�J��qO�s�H6z���_�{F���dQ8�j.[[F���4�o^w�Л7Z���X,��6b���������Ez陠����0���PI�wg���N
�0Q� s�E�f��;�)�Բ�.��=�qi%l}Ӯ�> z���1IfU�kԭT��Y�Vm��dޘ��L���N����Gv�D��wU�;.��:�
B���	)�RPuP�DP�cs�[sa`������Tn�����L-ݬPG�{�a��c;Z��f�`@�l2���*I~���_6���q�J�~xcuF3�2M�.�@���9'��'��"L'tëw,i@耈�/_���� ��ܙ�l���S�	���T�����SM��U�C�4���3<οh�Xo��J�7�|�#ؗ J�{�4\� [����|_�6�LS���S�d�����$o&��6�@{�y��n�����L�I<�SA�vΦ�P��F���]ZS����T��Hw����^��7�F�����YxR-ٞѴ��v]���@�ې&JQ'֕m>��'岧�u��dn�qr-Ǯ?L^���-#�T�Mǃ0��W��*�c��&\,�1_�6�����į�)ӍR�OuC��q_��ee���+��l+p�頇%'��a�����K�ؤ��B��G�4�s�j3y�w�9V�<�D+��Vb4�|�NZ�i�PTz��oA��u[�Ź) 
H.*Bt'#E{����X�2�Ytvq����%�ɉ�P����r���/�v�W�D��"�B�ŕ������x����8����,`=�������a1�Y�#�P��4��&8sD
��W��B@�&��+z[ �p$E��A|{�٭G?�v� �_��� �&�<�k��H�ϐ?��x�冏.��/#��^)��(U]̘8�#�����k6�Ľ	��(�팃=�{��-5�L�<c��g}>��h9Ӥ.���)��*�w�?��o����0gɝR�>y�E#3�����\��Q�,%�b�=�L~�z8���vw`|H#U����uU�bFE�ӑr:z|�;H;�cS)i&�B��U^�T_�N�,2�(����
�����HU���Y'��<�Hz� ��Tc�^�iW���&�o#O5b�κ��n��ޓ�r�5&����d�{�:R0hZa�X͚X�|����x��G�@h�[�a�8r!9c��B�+��1^1��r�A�o[zn�H�vh�	h}���ڽ��{1�Z����ҋq-O=�(2�p�õڮ?�{��V�Y�������{[�F�������4�1�|݋=�O�q�*�[ҫ���W��3�p5
8�Tr�b^�v�HT!1t*���y�@`8qq_[���Y"�*Ųʭ�>~�X��FҘ+��w��&���#pٛ��3�3@��cu��$��=2���r	5�xe�*�}Zx��S���e������-�{�a���j�ښ�!k��������Nw�$���m�|����0�/.���`�����	+V|��ɠ�1����)=i�8�NJ�癖mЂW��	��~�g���2K���Đ��8nW�T�ȗ1+		*ŋ�0�����R<G+��4
�x?YfA8Q��#:RP���TqB�	�t��$��y������ʲuȦ���ys�n�oY�Ֆ�ܥ�M����רV�y��@wCØb8Xl�`�*vj�ѯ?p�!�U3�U��RFzv�<�� ��#���iuA3)�j�
h@:Ly���&�$&1�,X���_~��\��FӺ<g:Nt*��G��/�u�V$fx�[�9]�]RY1<�dy���3�x�H"��)���N�����4�Iv��7���XP:�DU6�Va�������A�zG*�4�����\���Ӣ�5 I�`�y�i�.�ʮ#׋1,��E�>FL��eE�%�!y͉��Ր�*D{��h.��sD�Gd�9w�0n�5VÐS^.��I���8�A�"39�����U/�`�L.{k�q�A�P��(�e2��a$�uozf,#T& g� L1�������:�N��<�j��)�"qXX<!4���%���2CVS'?�K���o�\6�����y	�+i��,M�R/I��!����s�g{~��h7�\n��Q5�d��P����$��y%��7}搇#r��͚X���	���Q_J��.s���(�ZUn�%ehZY6���܅��,W�z�Rȣ5������5���K���6LY��@?u&V{v�M��@9�xRRy�V�[k�hb�>7��>����![�h7����%���;n�?}���ӌ��T�|�_��(f��% ��zz�o�����͊�J���.v��֋IM/��C`��8�d5'�
��D/�q�W�k|C�f���["��o�c2��?J�]���r��1@-�,��̒k{����e-;y�A�.]U�5J�;lŗU��Kh�7'D���k�'�����d1tKq���z�������GB��-��sp?�~����݅x�ah�M�W��li�,�q9֮��@�`q�졳������w��p�y��s��*H^���1s��{��^������ <2 ��#�dɑՐ]7ڎ2S[ƿk�P��ߒ#V��
��{�Rq���'	�⃋53��Z�A��8�����`����n�tJN������''�v1�ַ")�&o�N+���I}9��t3(��u/qk���2��V&�=�6����e����a̡���Q����c��?+�eH��h
2B�d:��C����V'/h
BbXGn�KO����v�Nl�[ 7����C�_�i�[eq���60�*����S8���
k��t��ys�!L��7%�¼����f��������*a�oDbg�;�m��*�rNuw��L���2_���u��Uڅ���x�3\��������b�6m㗝�2z	>&�^�o�/��J�$�7���&=oF��%ʌV���+P���ŋ�bgQ��A��a}�]�d�q{��"=B��(�@c��H�Э�)�gb�\��H�H�gט��C0�T��������W/�&b]=���sw��:���Շ4�������������d`�������*��s��� ��No80�͝��:tV�%�j�䉦8r9�5H'.�_$���@JY�㭀-�wQ����N��}|�7����y���v0FC7�ZDP��F�����m<�AIr�� ��ch�P��t�;��������jQ�?�{L����ڛvuc�M5��P�S��.qiZ���Z�Q�:J��)D��]��<��N�d�E�6�3�ȓ���n�1���q'R�]/-;@�F� �%�n�6 ����۲K'��J�nW�=A?��-��ɀ$&��ЍM��0!$��\U��ۉO��Q�k�
Y���ӿ�Zķ���!�4( j�lS�o6�~<��pOKt��e!��~�.Tվe Hg$H���K��e�L��3cv�:A�=\��Y�쟙����ߛ�2�^���ml�^}���@3���lc�>�W.8��r�t�b���.Ul �?cx/?�i͎_ݠ�Z��	�������G�?.��զ�e%��&ɵr�����:�كS�,���;Jk�T#9�*�Iɋ�'�@~����T�����=�a8���1��%�d4i��0�U#h�	�@�J����%����e���J樽�6���Z��$<գErFu_",��42p������M��e�Nȁ �.����{< �' �$�1���N��$.#M0�נœ��p�5f��1�|s�'����l9���f7[r��4����{�w�$�a�J�<(VB�à����5[�⮕E �
B��n9Ou�|��nI9�qe�Ou�]j<h�ɏ�s)�@=h�E�}��;��
I��x�҄�H".[�r�Za�7`��꘭����W���ҽ���.w��:k_�5�F{�N�[&P�W�g�/�ng��  Cܙ��T���=r�dd��󎾒�����l��f�����yD�γ!��4'��B�:�횑�[T1%g�bWz��*ˮT��<� �ІE�-Q0��1�V�oѥ�{������=�5�V�i??G��&f�����y�=��$V�Ɏ-Rwl�=�Wᆅ-���M6���#���p��m���S_ ��X��ߺIO���I�馓Y�6T�	�6oc%���C4:h���A��@�1�*3/��%a�[9w(��nF�Rt�����;��D%G٧���'�fUHQ_�Y��?:��wD�����@B2�~)���3�@�˳�;�K>'rn�Eܱg���=�4/#X�����y��A
]����OY�)�cjU�4�AfG@����g�������[7���4�R|1�_q���6�i �|u��8���F������Oa�m+m�i�pP3qw�(�xk��O�<�Fh.5G�s�|"?^���A����^�X�X�^�;�\�'�<2�ap�MU�u`͸�ɀ��=��w��<5�����	��W����Q�I�F�.~sK��V�h�8���>�,��tv���`s�O=�k�����F 褲��b^̓�g�}i54J��P�JǮp>��9J��	��y�Ē�gi��L�4��ɢ'��悍Ո��P������-�+s��0ۍN���}�x����:i��U[P�#(X5'e�y�
����)uv�A~2��U�<ҩ,w+���_�tD�	����9f��K^N"-�WxpdD|�F2��Vuw��K?@�V�$� ���7���L}v�v y�6sS\�3���D�n�仔�b��H��/��>�y62V�-�ND	ʧ�Ԕ,���0I4	�m��XF��$#'TK��F@L/m]��:�ӻ�����[��������h4I�U/�'	��;ca]���6|J�p]x	���/f��r>I솈�"���W�TPG�h /Ϧ N�vpnzw�9W�#��g^5nb}�x����4� ��e(�X����ғ���A�l�w��RV0Ml!IuT/%���ŷ��-��N3�g6�3�n+JO������(Ztul���4*K*GA��$��D������Jy�Io��Z�4,��~T�ȑ9� ������w��V�C���+¸g�%��Aj�d��Ń���s��j�\f��Ù��ͣ���N'� ��-�Z�������G�.*68Qw��G��'�A>��*`4y��������/�4`~|��~AU��[�@v;5뗾F��A|�<P��E���[��d�u�X)K�c̆��>��x���֞_,��>(��6}20�<��1؍���K&�{�Xh�^�]��q�A�M)�
QX�}j�j��<�Y+�?���F��N�[���2C�M^�+��re���yË���@8ȿZO��:��h|���w��6q�D@��sAc+�Z6�|o*D ����ڑ��a��|-��#:4���`�m���ޖA�������`a�Y���Agd`�~*�4��ɱT����K�B��^|-ψ��������t�飗d��MY��X,��Ԇ�wrd�4�(lCj8e�߬O-�`�ye~�!)�8'�NZ�lB��U����]t%;���wpFc[l����y�Q��M��ӵ�+K��F*T+k!�-X����2 9VL0}_r5���c�>d_*��S����ɨ�sF^=8¹��)�n��)A9.z�I#�y�*�D��r�._
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��F��g���}Yz�䦍�ŌO�H�k9����"Y�(E����
_>!$Y�#o"k�����*|FL}�z���!�W��8Y2Q���z�������i���5.���sH�<��p�}PH�5uI��9�+p�5'���Դ@ݨT�ԏ��Y"����Y،�
�V$���XP'��xƯ���{����M�39>�P7���p6!��L+I�זh8GL�lbB)�/ �yɯ��é�J*,2
��2�	�wQ�T˜��oPD�7��b���}���ٳ�=�f9�h�$��W��%uw'`�.j��롐�)BoPQEm���W�t�ʠ��N�8�J��
B����f�J�+��lǎ �/�"���4��ww��mN�9�+c��r�~�Hi=�u8���Cl�M^ǞHj�7O0
d<�k�=� �"�\f��߆	��9��;�_��r��������q��3EiaaTlm� ����0�?�]�ZDxr��^�u�<�Wa��֔�x�3�.yI�V�PK���UYu�"k@�+W�F�'�4�I���!!4¤ыFL�����	'�\�T���xa��Pu�"z��Zƪ��35�z�B��Ac�*�&�b�w
�32">;z�K�����q����Ji%h�.��k���qi�W���D�JRs��	��k�;�y\�_�<"!q{oI��GO��SW�4㬼����W��:�KXF������S:�]�T�wl��0���_�F�`?^�:�R��Q# �6�Zgr��]�8�/�0���/�=yo��m�bA����I�,1f�@UL`	�I��?�z��?�]���(K�����Z���i?f���0��(�J�nU#�*��C��"[�τ��.f�z]�IQ��s�_b����0fnG!��P2���(� V[W�ZGl����"mQ��a:�2쏸00�I�a�x���P�w~�I��D�hW�$�t4ޟ�,��YcJ9#�K�7��y����Ҭإ�0o��DC��M��9�|�ŕi���1���9��2S�>��*U+a&W$��_�X�G����h�`�)�F|@�'��5)W��ۡ��Ǎ��k�2��j��0�d�����rU]I�N\�g��p��Ц�C�o;�D���S�U\a���4��'B_t����x(���}�HBY�)�M�vXDDP�,��8����~b��gߦ�=�Z�t�R�iD*>�;�I�>�i�[���"�_�6�|��}���	�o7§{SŚ���#��ޠ�'���?z\'OO��􋷛�\�Q▆-\:qU^о����6��.!���pW/CB,�@�Mo���Ȕg}���"��v�lŬ���̪�F�Ͷ2���"��8�-�����4r*n���L��J2¤cy��0�j�i��	Ƞ�U/3��
D�Gu#&����k|��KH�?H�.و<���%��R���"Hu���x���^/{��c�M���{M�d.!�ޜ
]�yA'��Ş�����<ڐ=j�)��{ ���������y��ɪ5����=?������o��SaT���v��0�@�`���s���b���t``�����kGwnd�����p�T-�cu����+P{� �u*P��>r*�~�W�LtT�����f�=`̩ ר%�F�P�;8��A� /N��'A"��,�=��w�1lU��9�F{t��Lק������X�3ӄ�b�vs�l� 	��H�oa�>λ$l���!�.;ܦ+�1��8�q+�"	�j�xS����&`����>�D@b+�X:*!�a�c%g7<�r<ql;��|�h��9�y�"f�G��^4D���uC7?�"��d��m���s?Wm�G4��Q���R6 �+[�����E��Ւ��1���mэv�ט+L5o�пi�s����P�p@@�Ma̔�ԢA��u�8ߠ�Z��fR"�6��#��Y��w�	�Nع#l�p)&*8'�E[�*�4HjC�|8�褛G���ظ2e�l��BԘ&VR ���:��J%��;>Q��OM�w��|��W=w�(}��e�X�]��J�?������ή'N�,��E��0M�o�d������ڧ�����Y��v��2��n�	}K��Q���ܯH]3��Ї�@)J"-Ix�t� i%���Ȑ�*��"�X�:Ϭ|Q�a�-J�a���|aF��e��=��=��J�C�P��X*��4J�����A��vд�����$=���U,�2��o�u���bJ}C�a�2JW�#��`���mBZ	N�	>R/o���),���tLi��]�u-�q2�+���&�	�6�a
a���W��mT/����c�q��<^�Ai>G��7!垇����s�nd&s����C��z�8YR%�:�v%�tD��ͭ�Y�����c���A�s9�8]U토$]�j���)�Ӂ�2Zd�k�^�a�6R�
���K�=%;�.��gf�/�T
F�g5�IS��Z�z��u�_/{��kL C� 5-�������j��2��pb���oOy��DJ��Ei�%��r� =���Ĳ'�ن��_V+��h��Q�#�����i�G�*����#�Eg��9dU��	��dM�Y�9-���y,���sl���Z-'K*�3��C�aO���4w�J!�C�Vc[0*$x��>����[z-5�O��tS�.�WT)�]������d�1.�A*�bg�u�*��Fk$��0�A	~_WJU1��t<y~�)/�\Hjꄈhj�#�E��5�l$��!k�0���(Z9<[/�R�#AQD�ѾҠ(�����xi�]�`M�9�0���ѮX]�om�1��5����Ҽ���Ԅ�|jQ��P;�e����� (�bj��J��iR��FՂ9�HΧg�+o��oj(��㏍dxi��K���|_��%������>c)����Xi������a}n������$znڞМ��[ڳm[�N����%��v�=��|ɨr��U�� ���e�W��b[m�<�ogC�t��$�k��������|ޡjv@�������
�L6ŉ�ʅ��K_{Z�j�)F�0��Yٟ7��i�1"D�qހrf3��+�o�-����ƒ}�g2�xAt���` ��dz��ѣ�Jv?��;�5)Q*�o��x~��{,�N���̩Rm=�:�ޓ���ՙ�|`�gM��5��ӧ�z��ʾ{�X{o�~vop�q�?�GՐd�� z���s�j^6q�-���[0��S����X��I��p�'��yiC�]���&^k�|w�^�A��6|^�%�d�S8&�kA�����	�Ԋ`6c}�[qpC}����ށ�p�}���ȹ\,\�0أ������bZ-֌xidD���fg�$�up{�jx�
 ��|'��m˰�O�,!�1�i2 �=C0�6��m���4���QԠ�#`M�c��?�ަ碌l�+��Lb�&��gr�IV�(g?EW��E�L mYc�D��{
�4�QII�
�,�+�."\���͓��G��N�p�2
�S9�T6n�[�Ӆ� X�a�NG�u	�HX��PI-�O|�������k����!76��\��I9��k��KOU�u�7��d�֐.�X���0���?�g*�>zl7�X̸ďVੁJ�w�ov��]>������(!e����EcL5?��zg�ܬd��Y��4��*��q���y��o��9e{Z��5i�NI�٪��t��M���O
h%�@�al~]�� ���Q�m2�S�nM�K��1:{H�P�?��zV�x��-�8�!�nD@r�㹥�/�/x8�3�uˆ~�i�U�}�`!�q����piי v$�`���S���#Bhd�J����/A�ƹ�����>�ZN���GSS�r\��3 ���H1@N�`��S
����n*�����χ�P�N龢$n������{5���.>���#�
��Kq(�R�������4�.-���`��qP7��<hͱ�Ӈ0=������h5ʥ`q�dӸ�����,�a�>S��G��ԩ�\��k�p�}u�Z��]%���A�����t���͜�A�ߪ��!�o��eK:�����F��?��<H��ΎҞ�l��'u�t_af%,>n�ËVqA��:`u���Jcok
��0Z`���[���r�Fp$r���{��i��S�O��Q19�O��Pv?�j8��}�Zm��K��<9*�'���|�˙Γ!����S�荿e?Q�
�L��w���G�)/���ֺ�~��aLdM��KB$�f V=�	|("\'>����h�p[3���Lv��F���R͋O�"$B�a�fH��=� ��ȼ1@"�{ԪI^l�] �a+`?P�j����#�|t7�k���HU��F�UM����}m[�&��켍�넮���{����C�Y��)a��*���N�ϡġ����!B�9﹢���Z��|����*H��G��g-��� �_IЃ�"��㮌Տ�@���{gǹO�w��m�=j)ij��$R��)�D�/�	��`���|:�GȌ�`3���e�o������3���G�Kw��R����{�'���ͧ�D������D�̉k��?���@����X-�Hr�`+1uz!�lʕ���_d}�Q��:���~�Tj	)y�8�S��fz,��u�$7�"s�����c�n;w_������K�l���ri�xLtyB�
��N��o����h/"Fd�1���]����;���G��`=w?ZK럞,�o�	����j�7�B	Ì��Uf-���g�z��B���TA㘺-b�\��K���}[ୣe� H	�b+0�~��nn:L�	*ʉ7랎�Brt�y�E��7�z$ 711��)��/�RD�1r��LIFqQi� zn"�ҽrȈ���aYy<�+�yӾ��xL�L�"%�8�h44ӕ#͎���ڧRUY-J@�Z8��Ԑu��}��W�W�%Hp{ڣ�jS���ފ_���T_�_�#��>����g��'�l�֨���(��|����^����h����Vssq� ը���t�{\U��J�@�S��>O雧�#���tPR2,�G��lR;����48��L��
qn�(%������\#â��rHm��A5�:�r,;��iQnB�ɾ����F��t������������{(�v�s��%��MБ�������� �S��4V�P�7�����(��cMC��5)V��u�f�dGQk���D�5���/ q6�_�]����H�� �?���-�Bfl�e�o�$��L/��=F ���ed�ݾ�'3,F	K�%�������L%���ڱ�o�E�
�F�����8��ڽ�E�t�p�=�{�7I|����� M�����Uk����JrĆ��R>m����ͭqઓ3�%��Iz>�6���i�R�H8�]�
�?���-I��q�z��,P��!�����A��?ӋeV	�6K���N���5h���O��՟��	��,�!+>���%×u�����_��>�0�ҖVd��qV&��EL����Q�p3Ob�v�F��yx��z৹��	�&<(�7�F�ϫDo�x���)�r�n�xy{�/�9gV()_����"�t�y���Ek��3�p�G'J���e��5�Ӧ>NO��n3�4�G
LQ	���㕔�3��\E�֣��M��`��!����
s���*������T,���Yu�k.�M��S��H�m`�!���\�q4���G�+��Ǌ'��n�!S�4	���͚�=j�	yZ/.K+h����M׀�o��K�yr�,�e�z�*>q���t�`�� kԖ��C~�a�<>OyP#yRexn|B�*"�-�]�Z�c��1�e~��W�7ڽ�hƣ��jQͭ)�G��b�"b�*̵Ȣ 	�x>���#ݺ��GA0a-��r�X�&J��ȍn�7c%�`�Q�0�����Ư@T�##�:�u~q�i)I`.3�A�T M��I �ipbz:3J�x<矃�&*�,��(+�J�Ds^����7����'�w�0����'������H�f�:~���)�10пH�&�p�h.���N�0��� ����&��8$�Ӧ;!I�ۗ�+��ޡ[��wu��[F
��Sr	X����X��'S��[����"�� o?r�M�Ȁ.n�_��:3σ�r3Z��G<�'�$˱"��/�n�e",qk]=)�s۶�f�1�*�\^~���}jN�hq��W�7|ą�����0�[�8<�2J�eH: ����R�h����5�ѕ���vz���Q�i��=Yz�n�b����D@7�u+��S�N��eАI�i��ֽ"y�r���X��o�`�O�p����/́ �Y3�qƨӽ������L��B��B%|����48bo� k<@S�!o4X�靆�E��@�S��1Ӓh:����QHX�p�!jG�eJI�Ȅ�{�C�a�`�S��)���g�7����T �#��@_�u?sx��nN;T<9���u���yZNڧ�is*ݹ���)�\��c��^��r�zO>�!�����m�(��C�|� oQ�q���'hfD�}�7:��X[V�`"9ݪ�Y���g�1�w�H�f��}�d��㬶y��3�,P��� ������Q�^-�XRVt0䂌)cQ��K�� z]`�a��3y�p��U�ny+��i@N��=��x��y<� ;�?�obN<��q ���h��j�PqNU)�-��|��A0�c:�ֱ�Oe�P�Ҿ �uM��"��S�DDm<���a6��8c(@�PN�@Z�e���Y5�f���.���˂ *`��6�o�p��۾���I�nM�\0�����qW�P��9�s��l�,��qL��T�^_>.��B!��t�O���ʃ�m��M"/��Χ�H �sS�X@i�5���u"��3�݀�:�����C9
\����'/>g=��kSo!��x Y�������<����u!�n�O���b�/��ز��Fy�xG5�2�0�2�&s�uaW�K�wָ���mA��#�q,1Lǉ��$Ey&���q��f�Y��:w�����g��֎m��I�I1kD�8���c��#��s�m��H,fkZ!�^�����b��Z�7�,���)ĳԑ�>iB�wK7x���G��_��+�)0�u�b�|X��h��:Xڔ��}����@3L�2C�~o�I���WOg�|ͭ,ߝ���ۿ�g��\.�}u�O� ��c�ХBh☸�mM�-v��g�3�tP�|�m�#:�5�0f� �o�9o��^�Q����>=����*��'wlP��WZ�d9y�����'�u��CkǊuf��߀��Xq[%������˾�`}�M����O�����Q�"��2�s1e���ۑ�l�je��nG���
��3-�R�M���3�=j-���\�My��ѫ�l��`����nɬX��c��\&�d'�m�A��9��B����4�/#6u�Ѽ[EM���.�./q�����ӵ�7���S�)��N�o��ĄVG�{D��ksd�0P�I'e����p��܏�]�_M�r�kDk��cS�C+B-�d��V}�",�=���F��"��In��'!�Nj���� �o�����	
h�����x�o"d��-��9��f�a{Y����5D�x[e?�s3�PmTÍG��G��$%Ǣ)8b��7�UW�
�(Z��,(uT3ж�����^��o 4�sf���)<��14|�1C<ԗ41�: uz[5�#l{'Ý@�q��9q��K1!?�X�,��\]֖��"�}�V��[︾�}��C��Ŷ4��d�dw3��X���V��F=��m' Z�Ul�l�Lؔm!�-%�+#�I���=�q_�?3�PV�6�J�Z�V% �?W'���k�V?\�a�� ���Tλ Ղ\[�D��HIv��x3��W���	����T��L{�f:�����)qj��$�Z��8��z��6�č�{0t�>%��ݤ�2ǘ9�,xf�|n�$1��3� Ȋ���Q����oF����f(؇��S�[�����1�\w���n�ϻ�cp����޿�~�{�c#�\�P���U�TW�/g�7��ICɝ~Pߑ�E	����G�+��
�L�.T�[��E�[��a�6	�`Q�� ؈��m�5\yؙ�s�ڍ�H띕^Ob������q16@�q���#����?5�d���:���I�	}szh4D�4g��%��bf�|%�	d�ط�>ЧeV����+"h!ܐv��dx�U���~�؆3z�EQ�����^�D��*�GN������Ԟ�4�@�ȩsĽs�-$�_J!��_ȾW��g;��14��"�-YE�E݆����s�ٗ�ӱ��o�F���o���J�8�]� 0FmWZ�[�O���D)P�$B/��8�͵��H����ܹd����V��8~ܰ��8�qA$fx��Q-�i[�m�g�]�9��Q��ŌV_�����mZ��I��$+3�1q�m��`i� uՓ�,^N�%a�ne��y�X������T��*����Tڛ5B/�$���@�7Ro�>�(+���L m�P�6\��/I�q6*`���z�#�s���q��vb�v��"[���, ���}�� g��N,?7�l97۰2vh�$�ZC�������-�j�v��X��p._{�>3�'�t�������n@�r�z�jm�x@�F��o���Ew�+b2|,��o�8��l`��fq��0��[�砂g��2�M�X�����dH�%�@N,���K5�����"|�w!S͐�Xf��g���	��9��o���������sǭS/Hn����*$d��_�A�<�B_�me8�_�ʤ�4�Q2����T���M��t�T}��saC�f��ߧP� "ps2���6�JJ4�>��&��hZP�a��(Li_�=r�x�a�8Y��!�ɯ�|�M��۳�ܶ������J��r�N�!:v�u)�� ,uՆB��<Z�����4l� �#�'��;##����e�s(��Z��k
1%[F�g���I���_"���@��[�]� ��(.*�Ţypu�k��5�!a��x+v��m��T���9�ظ�9�~�T
Z���������T�WyR��g��⭳�y����
�S�	A�s��ge�����d����]�䥦�v��(+MI`�'q��Oc�πj�O��>j��c�>F`��Ufin�>��:�!��� L G;��;R��t|�M/��aS�!IH��[�O�;�C*�|��8��?���Hd#)J��T���.y4�;z���ȩ*`+��#4A${�t�#�"�B���;�_�=}�C�gb���("�y�W�O�Xj��UlPx�3$�3�XN��1tE;���;� �݄�ˈ"z����'��K� 
;&},h����i��!6)�6L���d��°���~�U3�N�}�wKu▕���H��f���pC=��CC�U�?J�{gZC8O穃��t苸��o Ρ�<�6��mг˟GH���w�/�gو�<d�6�s�=I��"|C,t~��?�S�����^� (��eq�^��V�!��}%t]���Ϯ
v���������}�)M�m^��\/<�K92��)�rt��^��� ��o�xCg,��	� ���^3�`�Z�j_ݤ�ǽ��8�p��!Ypv�{�x'[���s[�&�5u��[H���zQҶ��o��4��ȼ�Ӱ���Xd���f#F^^2ٽ6�8?<E:������?��Z⧭t��.������M;gb�,�c����	� u��K��fPȐ{���)ө�V,�9�}Dט��E��s�z:v�¥�p�����~p�G��6���p��j�yk��;o|;��@�}x�G����@Y�&W6���������dO���8��?&$?kV�g9lYj3��?���GÈ@Z}6�`
a�ėj�r��t�b�gHy�mv�J��I(_�D���-��
ɼ�#�ך-=�3~ �{&ny�P����ېA	�OB�Y���,�Xl�l��-{���7�fgŠy��'�r� ���q�RWy;-���7|*y���.ҎǓOFv�W��_7`r^6����ܱ��X,i���Z_�Dg��Ps(�C�*1ë�4{�Y��ƴ�4��4��Ph�M�M����Q�V.�� ���+�.��`���ҿ��h*��v���AM�����Өy*�v@v����LJ2c��T=؊Ն��#�xR�C���zuA�r��m�P��oX��\�	 +��rXO��G�Ҵ0�ĕ�ƚ/���as�J���}�6�щ�Ծ;�����C�<�K��+
��M�:���	��L��mUm&�z�Li\e�9���
�QOO?�לI��+E�'����}���]�S�Ru*�T$h�o������8w���h�!�)Y�}±LZ�,���y;̒��e:���Ц���M��],2��,�;K��_<I������3��I7P:5����`a�&VdfHR3d��U}�{�������۳c2���f�b� +�2@���go����ړ�a���c����ԙ��<çZs��]5�pHF�CY��~�e��B����\��p=y����E�%��DfV�:�Y+�3���K�N��6�Ͻ����~|\\�^�_%Hr�J&Q*u��{��i�8��[����{೷��[���`�R�ĭ6A]/����HcNJz��݃:	�p�[���Wk�P�w6;�c�_�Q@aPY jdp<
�]hr5m���n�Ƨ����2�}�4��m{�Y����m#^4�ك�p�k��D`�i�L0�=��u���ch�v�Zs�Y���f�q��U��6���k]�Xo���K4?���m��+3�Ԟ�����8�W����A)f%��[�ldN��t'���҉�r8̌kzw��q;)�GR/d�������x��B#@�fZ�5�f�\�U��z`8�"9��p�w� �k�D;z"Gsk�1	�� ����K�)1$9�"M��e��r ��Δ��M���Y����n�����tn��92��n CT�8�1����/�� ��:��9X� &,r��>`	�w�ll�hnq�]kܐ�
+\�ՂWo���E@���7�r�X�{�V�>���\QpV�(b����ӓ\��h��X�Ĝ�v�	�p������R��5��W�p�=��>a���эdr�If��G�Ȋ 7ܧI� Q;�����4�-���P�?�I�O����1�k�FPb���d�ɱɭ�U��x1�Z,��Ⴝܟ���û�P�*3@��_���!=A��X�M9����hl}�����Ov����������8b��d$������e$8&9�l��a2�Eh*�ð��b��p��:��bQ��1�r��(���]�K�;Շ-�8��e�c�xT	�@P��S]>�)�ǜ��a�2H�2�~��6�3�a���H%�?z� =�BYƊp�a�r�ݍ����:�̨@���۞uRn���[(f�m�	�Vu��H�
��"�o�W��5����SW���86vwX婹�)A��k��H;h?os{a�o��TL��N
������<������?� �W�,N��T>����3�?���P�w�;���Q�Νe���'�P�A�Q(���Y�$YmiJ�q`�?SW��P��W�z�@��ʶ�ףl��X�u������ݻ�L���FͰ�2��w�8����N�c b!����۾2�k�_;���|=m�=`7��DA)���E\7��}Q�.����%�&?��sm�p�MBʣ��9S��9�.�|ыE�Ϩ�,��7l��̽��ֻh����y�V!�FTFfR$mQy��x�RP .6<��;�x�'ӡ��L�I�K�0^w����1n�7�g��H��s�s闱��E�6�S�Ȏ~�˃���2���\������{�f+
B����>�?G5w�>�r�,�r%Mqw��./�8�nfk�Q+�P�Lь�'q��t�Cff�k8R
P�������7�1>��U	8�B$��$*b�K.��x"���:�Lp4�l�U��4ϐO�NN�d  ����S)#y^'+h�3ʲNpFOz����(0"}�J�*���O#F_��ә�@02w�:������s"�����<Ճ#p�<'�R����M�����IX��{��A��y���D�tZ�n��
�d���E:���T�3��nk����l�&𖞩H�Lf�*�C'}��Z�>�*0�wA���72�Ǿ�LޢG���U�r��aPo� %�5��$�n��^�<�c��>2��� cXϋkڏ����L2�#�բ�Ĭ�����L:�x(���1,F��57�r�f���>0��;���o/}W �Ցp����sSiOׇc�<�u��LS4���T�!�@� FD93 �:���H� 5*�~���䢭�{�Z�&c�e�nB�"�lV#n\(<r��8i�%��Vp_J]������Cv��I9�������H�ka;j��ܺ&�`�&0�p[NI2r�|[^%8�),��v�ǎ��$��~j	u�����o�t��˙�������+���~��*�I�q��S<ҍ,*͆�*��wV RpC�3%�@¥��PG�Z��m��\�!W�y5&��6,�jbK8/�zE	�i�������V���N�C,��z,�H��:��x%���fyQOY���7i��:�ZW�0<=���;=U@�C!-\/ň�iR�i,�$:��9��\�Y���'�@��ޅ���#v�W���?��I��!F{��46l��@��Eȟ�G$�歏�c�/�h��B�
RG戧�<�n�:�P��u+r'���╪[P�n1Gz�����X��nm3?\�vY�}����H񚟳�c���;���ǟ�]R��[+Lf�Fz��ZF�<�a���<�J|����'�+��"jY�+Urx��E�f�jS�Z	x>?�z��p��3��:@>��m���B�
s�^�\�0�s�����t���O�߫&~FD�	��������aǚA�`�}l�I�<�-�1K9	�+˭$����k�/�<�-oO�!�?�y�m���D,2�?G!XB�~�/�≵���Mi-gW#�ۙm��r���$����K�*\tJ�\֟���jpG��Ƌ��"Mk���	�@�4�:ץ���3���H
Ҕw�Ϻ[����T�H��z��+ou���?�B:5[���i��@�Oo�;R��"K�و_س���F�8�����D	5�N���vf2J���=]�[�����,Hu�^ŴT���dbA|�jzY3�% ���d<ذ�<nH�?��WH��H������{���G��G$8��$q$e�w��$�'#�b��2q�X��g����\��j%X����1S�
w�l��1�Z@�򩽢����iX����S�L)ݖzH���i]R�8G�NԚ��9i�U�o�lp?�k���(����Ҽ���PV�Sc�;D%^�gD�F�tr���]PE����@@���>�Cp�CsmTi�Vsp����'W��W�>��7
�3�˖����A���1��dp.%�9�ַ�]_�0�"1>��e��$���$At
\9�7o�
F^��*�������6�~@�!�������؋��@ԃ���4\Wb���"i[��H��p8�9�+`X�$;��0�d�y���b���i��`���p��n�[���4	tִ�a�]�(��(�s@�h��c/�x���7\tΛ+@��K�RHU��)�ֈcZ,g�"�QL����f<{*(9&?�4��q���83+�̬�_XP�u�}�� �##��/�{A�!�j�#ƃ���ԙ�}nm��O)�k4�6�E�D��O���;w���]�����CY���ܸ�5$HgV�Y���gH�h��bF��G$�/+��Ɯ��߷S���h˴F���rv��t!`S�A���4e��p_.Ԥ?N����Q��cF��|�M.F�k������A]�s�kIzI��_[�4��ెΟ_4��ۄ2�)���%��M֘�T��d,G����Rv��dq����I�'���_����"�S�!y��P�OB~`E��U�[��?p(?b�b�y�K ��|ڹ?m��S���v�C�<w�)YRq�Jj��]%�W�]W�{�:�Π�e��"ނ�PB+�����;#�D��aD�闹�d����^�p���F�А��P�L�+���Ua(�M��c�ڽ���I���p���/1��?���#/~�/ ���������i LV�g�#�6?qYc-��#_LW髩�d�lV�����8�����郋�riB�>��v�O�5t2#}W½H��I�3�9��N�'���f9,�#�"��T���U��ن�V+���@���5�8�p�.����٠��,q�%?�Fɞ U�o*zCnI_�To��Ⳅ�k�RT�k��!���D�+�	�S��vm���R��h<�����7ms�a����Fl��@*�k���w�W�;��/'+����-@�0n���י��5���p�Ce>7�Ѽ�#0Έ-����1]l��K���.
>��ݱ���ِ�e�n����NPa�:�)��J�K(���{H�����;���1� ���>c����L���5x���z���m���y�+�5R�6�./�xD���~�yW�vmC�����p����_�Z�ׁ�
�xK=j2UѪ���8��l��}�ҹ�R�@��P�Qyf����A�vo2l#��RiZ`��bd�=y8H|i�nso�J��z�.���b�3X���LP�)Gۢxw3�h$�n���plj�DL�?�Qq\�':����%������{,��9�6��Oc��J�g�LX$7�J$�R�򦣰Um���}+� ��|���(��
�ʟ����<8�L\���� ���Խ�����od�I�� 'n�a��v\��,��rGsV���s�Hb�u���w�Ur�t���4��_N��"�:ތ�h-pkj��\�@�^���uH�Q5�XUs��'�-�&�Vd\�2��+.
+�zL��`d�[n�ŏ?e��"�5�&󫖦�壻Rk�[�Ku�oΝ�V@e�� �����Ǽ,Y�*Q/16����F�L@'��y��fd��x��A2&heV��ﴆ��9�J-h鎎GU(Ku�#(���.�"ehV�ى�=���j��Qzz����)HGv$2�Hl.[�%�u_�yX���)��j8�7W���Wz��K�ip����wĉ�kGQufxM8B4�P��_��!��Gmg�*�_�a����=�oRq��s9�X��<1ú����x��y�0��o�R��C��5��-1�K�������C�߆���Q⨿^P�<Ml�����9�reJ�����a��	���X�a����eɥٌ](��E�X0$��l�
B�ZUÚ����V3� e�|.���1��1�v�?0�Jڑ�ޑ��J�À�����޺�p�Z��`���.Fm����ǏD�u}�w���ҽt�$'~�ww����JXY6�m��Mwq�Prg|=C�!��qR���F�B'y�:�����gQ��I�?^�꾍ƘP;~�]���(�W��k�lk�?�$N�x2p
��fz���Z������ <�S5jod��6��y e�A'�T���70�]�po��1>'���������.�%a�[d|ZXę���U�����H�<�.u��j�`m&�K壂��H7|[H�� qȷ�9I��=}t�۞n�~�9�iOk{j0�55y�k��MO��w���HKtE9�K�VC���1����YB[Ε3α�-��,��(�#�ACAR����T��V%��{���蟈�X#(t���&yP�֪��_�1D����[��!n���M�WT�`9��|������ �ʿ�֭Qxg])��*�;xF�Ѿ�������w���!A�U�L���iHb�d�UC?�xV�2�/�͆m�x�mk?BA���K��ߏ����+�e������u�i�ԁ�Sb���'aZ&��~|���:�̙ʌ������4i}�n��'��Q<WK;఻_e���qC��İ~��#�(���|LJ���2ҽ�����9ָ�����4�A�#UM��l��úvdS�R�6v�w�pi~h繻�o�կLV͖�/t�[Wtk.��#Ӡ=�ѥ,JR�6�I�0�c�/����	|��������nJ�	�L�[���Ì&��p7���¿r����gQ�r���$���~WO=aF����u!���LK:�Bwk0�`D�{���풫؏���q�#t�<�0�*��hf���a6�{��_��(���
�`�xf�Ԗ�ƌ��,o�<m/r_��C�60c�*��O?�N�h���$������d�U!dp��ŐCᝃ���ϚE8N����d\�����`%��fe��]r�sN����"��k�c�tvLhB�,��i�ȉ( <v�bh)���[Y�F/Τ	�A;@^�o �c�➴Vc2����9��qѝ�
rz-�[&M����x:qA|L�=tZ��U�a?��@@/����OR.��vy%�4ס���e�z ��l�&.��� 8���6������S��}�7��g�K�N����-�zuFY���_Pغ�O3�7�F=D�]o`�p����ڤU�I7�!ǡ:-#f&h��T�e׆j|���ċ.t�
O�GV�L��׹�����{ua���JD_H_Ȝ�G���r~�8��<ÃD*�\s��$d�e�[���}�3��ߓV�:��9��)�&P�}���%:J �Q�E1��(1Uv�8��l�r۝����mim�-	R���9�jq��>���Z�ù�����k�w)������ �/_��x�4:�	����8[v�~V�W>�� �W#k�S9ĳ��X�4���^����%�N���'3�ɮ���8�JZ=��y����9\A�߿и�>�|�g�&Uu'��h<RF��9����x�9*!��^ֱ���!�_Q�Q΋!c���`x��E�!�96�.v A�i����]��w��0*^�dx�(�Q(���Y�[Ŏ΋!�)g��E��N��K3�{q��p}��- 9K�`{g]����x���Zuv1�X_9	�Z�\gp��O�&�^�U&��ҿca�"Կrb�X3�������Oe<��Ӏ�5�,͌͟�U\Z��_'e6��4��]�i�����Hj�8}�	��X�"Yx��f/���}��
�!��S7m�x�]�-�'l��	g:a�\�)7�̝Z@/G	�spV�����A˃��k�~��&o*a�hv0��y���[C 
m�/��ቫ�O�'��c[1��:���b"*(&b��N��z��~�٬�>cD��ω��9�>�
n�]pt�}f�!�����I��$�p�H��E㴭�~��,q��^Z<���%I��̒�fi=�������|(�N�¼�g���BJ�
����>ڃ�AQ�᧥�CqDrs~����^y ����u���X˥u�c�NV���,_�`���Im-U�Ċ�G�w�miE�x]H7�&�H
�s���� ���T�� 4z���!����O�����"�}��w�ٲ�S�H�Y��ɇ@�T=@*�$�։�dٓ����v��C�g��颪����啑Dz���D8���7��P^"{���	���x��]�u�ި�W��^8q�!�й���ZCr�!Z��[��c<%e���7�PD�a+�V�G�8<�[E���Nm���`s�2��ae����0��CÓ��z����%b�:��Λkp��O��?ͼ�o+� ����:S�~�/ 8�~�����o��MN�-@�@���O��|�t���q���s� �dۺu��v;�S���"I��}Jǲ��8�qi4�eJ������/4T ���z�3�.ن?�j2:�Ъ��o��4�ܼ{ӳ�&@������W��"��u6���H<�=��'��b@տ�h���han�V�I���K%��.��Rf$�m�r}OD���� Pb�y��x�'�����?s:�;K���m\y��`�,U�M��!(DU����vs��G|F�<�-h� C�[��\��Mc�ʺNq�b\o����/^�#+m����T�0� ��5]��) �
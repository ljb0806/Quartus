-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KpyAPjIkZbW1nr/8h+N8AiXBPxF2OhmIzQ4dVxnve2/71uluQ+xYfpSXilUKj/No/D9qjpY8h+f5
LlhJsUTtp5C3DtLtoxFKzPU6ILfRo1kEx81qQtC8r4kI5ISJ9pmEyHDUmdjRDb5KXzvM94VNImf9
ve92TAODk98gbXFbYghqPQ7UkWPfxE0u1eJX7+5WpL6ABrWfxpp+jG6cQooRE7ROZKvqEfBjg1JE
l2OeobfWFCRIv+MwcXhFkHaTOUjffEDGTw3sGgPQgMB4WYwQ3QHkmrkEPP8CeIIUDnATEMClOtBc
uUV+boSAvUR4vtzVQ2jCSiWRyRsNgz8/YdcSTQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6656)
`protect data_block
0xu8TyUo/jTZS8yARHxn3WZ9NIogvwbreZcAKO+h1QHOf2Sqf8Xcsf0YY7+UWLqJSQrUvArY+WIi
ACATwja1VagA+YwF7SDpeou6MQJQRAHHRpHZZp6kiSVd1qHDO/z68KknSbb+R8ZaM9A+fT0L6c4H
S/Rzmbh4xrJHrqTlKDEiCUfeBWpgmEwpVME7vpnz8fSKdzK2LGMzjtsAmy64cO+SBuVN1kBndlyz
7K31+58IEdKM7NC6ApjEJ5GFFsAJIH8k5ptnjZ7Fg8n+dAjUxttnCbt27BD5IukrB6MlGB6UgLEC
5+8qcbDNvRp4ekWp1zRfeO+p5nHdza4UHMqjx8rTqIUxlINo2JiQVwscXX6d7YnY+5RVskvw+u7S
k7hmJy9fEqkWcp1Zk/mpqeF3oOj61IWWZnmCjtahZCVyloInh9TN/XBM3KS4zdBiDj+yh4aNCr0B
B3C1GZccmTHWtE133u8Ps+Oi4+h8Zq5HC4IRKuBPBFtiadB5Zvxf0vH3iWGtgONk0lAQEe1XQLce
+Uec1cJX+MY7No0l/9z/n+KT4Ud9sui+Nex8VIr6ZXq4rUnB3FM4s5HpWUtuHnVoSJrgcFdhfXyy
0pyBDn8zfI6ncgaZkVaw9WUduFRk50cJAKrSjTzHOr++eWh1Je34u19CHvIcEjxj9gssNozmg7qt
34ceyx3mO+8tGB2sJYJaTctNTbOXp42UpNLzo6Ax3E+osQWps+ndDhYcdpaH25/KuYgppUbQW66+
xszxNTULAU4uuv+QEd4YQL1CFBNFceNMa+gT/S9PGs+QmMlLDs5hPsdXNFG13H0moKANtPrNaIfK
EGkvSx1uBDoDXztoPRYSj1gPViTw8suxqHI6uYZ7bGANZu7nB6MdTRjL2Rx0WKtLsJC/jpSekJBB
1piZQMT9OzcMdJ4yzp0eEpMz+B1ndR6IHq/g3Q/fMbwcv2ezV73AcopEI9skpvPHEbTIDkh41WV5
lrC94W03EtVnyxfxHXpXxkSbihFfMuyp/Og+X0xwfLNkgd+4MwuOAvLUk79cgOsE5H54bzmNAnNA
gURAwJC0NQBlv8hbO8CXTV6eIEUb3l8ifCTl3jo5RYfyljWkNwQh8pnQ0yCQKfcOmkHljfdF8Dgu
BtOlxptZORtytz/hP2HlWbhK7WeUBoVIcrQ02F1BaB2dlUoFjV/nftvFf/9hTXpXfd7mPGsGmosf
rns+5A2svi7D1zdK0eDaOvnnyfBZanAMiLJnBonoK8Zjja3fEug51H7FHAC69+JxTFJz7x/1SlG7
aQLa9ufHGbQe/2d9fTUW9WMK4nN6Inhdn7ozTpaZi44/23XOhJ7JGUrdxjrr3TswX17rjjkxjd1X
eakYoBjrottPkMQ0neQDtfu29bosDD+1s0ojecsKjHgabqtlRtRnTpQ15bAJ1xzYvv8tmCuJSCPc
vdhYvl+OcaoWZ/J5gR7ewovLS1QzrJ8QXCc61lkxjJfTYOeaMV9yZql8HmutJVsp6ZcQv9kIFmhz
I05ohx4478uedvRDRKdZNMEjK+VlUmMMSzHQbWWYwN9KrPsczhagPquG6G8ycTrZIVhTjpYHXjcq
R40XK819BSMmwCEkui8RqNlLfcjF/haS8L7hKnUI0YuFwIl/RVT1EEqjplNoH0pOSZ9kEr9IcHxM
PHcxOoqojNxbQD2LuBZNvdkeCswTp9ZLkIh7orFZhu3RUoLQQDbz/BiR+4AlIeIUtblLw85YF+nA
LzFRrCBSHdP6tiHYoS2HeGuZs7mcBKEzwirfuJqsv+QDDunFvro9whxdgbXVzjV+bK8gHMU4US11
PuJgXGE3pqRiCEUnd5gyzmx32aHZOXnhqDkNdOe0O/zZffwJNsMrOSsVKzx4OrdoDI/Kw3Rv/fDq
O0oMkXbiK2HVgHJVoHkVsZSz9FTdVYDBPp+QN6Nhgi272zxZHrFC2nw1q3t5fNAqZltgk9WvIGVS
QeEpjF4ETilvjv4OBNMrFz1/gQAUpAhyf6JWkddvqAboQZtaw8sNZ6nY9Ic/cRut3xER3fiqt6pM
6YSbmWm4WJXtUwZm75yd/1d5GHlgZyt7MklemQgy+/h8mz/3r5GdNYgWR2g1wJH2Xh7SEeBqEZA3
xPiSl8dC2fl4yIIggIJyeGkF5Fc01J6NXLHiyvOG2Wqa8EOM/SdtZ53NixkoQOLK5iY3nKp4aDPf
ND10npsyh4w2maa1SbtSwpTA3+1aPGRHVhyYHOPOJl5hn8VDWOPM8eQXdgL2Y4tnHL9zD6essSDU
0y8MwpyhLt8oET99anTMsamAkxveV4dhYQ8yi7O6nZzKxVE70ZDyAW2EmfDsX/Lkv+XG6/vcN78V
KEGg3wbd/hlZyooOw4S7nAwsrAeeOgQWgGICfyK6PzFpHfbOUknrd4YDhZDP5x7tQEZzhgzcyk/I
8xE8HNTg/y5qTfkrOtfc7JCJlZj1q2p/iYLox2ddg24wZoz/XbE0GdPdzKFjAUy8bF7oBwQW6G/5
nOT8V3sZ1UKU2O3Bbs77S/FzOpsIzh0ox3XxrkdbsgZ0pg8yZEbqZcJuRNEHh5j+udh1Ib+yyhF6
0bJxmX5jXJAvmM9Zqt/5PUhAI8PggvfUttIJ5mW4na/9hcvFevlp8DgnbAIB13m9WrY9r9E/rd3Y
qj+puP0IBZF+WOm12YM3u4Bw7h9WLOi2eRt0CZTRRT5gU6ITFlGi+gH0INouIsw5Leab/lC8e7Bc
8r5p460j3jK6ptJJSagSPFRZ9zK1EonQTbLGB2B6FvegJP9hbNgfKZR0f0Vd/njh1F6kF3pFfwxG
ETeifV7KxX64A9hDMN06twSh3xNxKMDOPRsE6C3vk9OB95LVgpU8O3jA4/iyRzT+hIycvJKaAmg0
+1f3Z5wnoKl3IrnrNllJyb/LrQvOQQjOCYgBCxbbUmD6b0TVFX4cbeygKHnBJvD6RJX+0C3Uw5pE
UnWrZ+wIMDXUvsStJSeoAN1up+Wph+TjnxVuZJhCOqGVd67z6ZMs98fBdo41vpCHgDhtmGtp1Zmp
IxhHHj2neQQPxh/xnOJlOFYOPFZPW5EAnVw7JgurPp89j2uPCO0Mk/cP/EEqBUhKS/XT0KPgEnWC
1tj5sE+/W2fRdT9nYIIy8IX5wArL0xYMxT9rPBYgZYlcZdBdpgs/f0ghHsd39FUmIWHDoS8auzjP
228N3w+LXB8px1DjPH2nuLoCYokSv9IoxAbzCsZFyvNGLzfulTRhfAheEjUxavJojqmiBBAA799y
xyyfMd13BPdMfpBTqdCGWtl62PwWtUgmvUtYfpB+LHp1dtxBNynSZuqnD0kESZ7mwB7YzBSTRJVg
6M9NTCTmBvkN9QgorUKHU1GZHgwRt6Vq8oyxrgDNPyBQolXVN0x3C8tlm+H8fnaFFrvIt1i7advZ
YRfEHGsoc2GSpD1pYKFb/jqmIUU+Tarnb+wcaGWf/ThX7ZMQQT329SybYSX2cXMtRiXrx/lOvEN9
0kSP36TmFukeVh/vHcgn1D9MlEEwJbgqrPitJjCZmONJ6jj66LO7OnGSgyl7k2czabl7n+eqRlya
Z8cdl1e46WrIGNxHuQoPAIDj2snRl8bjU6AgzZRhrzhclQmfBdooXPLmElvz06jgOM6nkWuyeSAq
mP7R8/kcZ/uRD7M9LXtKp+oMQbNNZSf5dnEBeOoyiuIqmhdWueYCNmRjl5+gozA5gPXYrkpslqT7
GFhluKweA5GlctqGxO+yeXFx/JmvmC8fs7AOc5ESahOiebKlyxII3OylsjxFoOiqTuwjmtP5OJpt
rCbhyHN8yNOIoTzw2ufrE0kwD+orQHvWKztL7NCZmMkK3xuzYEgkyg8dwh3JS/lVeeNwMOZENjAr
4q0mL4RHVyq0QDbEw5dTKLPznnmSN1mGB8+0Rf0ANQmGKO+FOe0S/imgVix8H5yKYI/XkVxO4dTc
c5cEcgNxCRqOI+gl7hVWt2GBGKlXAjpcnNH5lAwy0Y4mll0e6SlMztHXajX1m3fv9dIodgSQu80r
WsQpDDuW2NxTj596Q3Kcn0djaMkGW8T8HR0kk775vn3Lfw8m+SBJKEw//8+gTZJbqdx/ZritKVCg
TgqZ/NLK9dih5b/JfEP+y+dc+SIUsvpF6kTeo57lErIeY/T9See2gRQnzNF82RwaaPoKFJ9TCM4V
yCsno6PnPmhmKbRvVTaimgttIghPPZg07BtTXHlRBzUdeKeje6MCgPgPpjELupifm5QEpnQkJrn7
k4Kkl4TuuNHIW4W3+Grf7XOSGYvHV93tiWnQpILsNTIIPbIAF8tTpvE9k6XVo2xo5Unl4bbGFrs0
/vDo4kLg4YtZ6L2AdOvVXz+qWncVWLnfILpXjyavpRUBw42T9l4cUQKEmmtcEhkhWwQuvu7hp7Lg
FiLabZMYWpNJOwGmNfw0qCpWvHg4xzDuLoGmEhtuFNAC+MxA0gJbcoy8uAcWDUijonX6X5IT/BTe
PWwV//KV92nswpIknmh2HkI7iySFiUzo0Wi0tRTy/q0pOYUySJrBqsjAAv3xeB4SFF9OsuECMGLM
ufMtSwEqhzycRT/68zQCz21sUbnZ4PpT3Y0xUjX7t4WcJbB91jh9hvtBQWogp4NggEXqsP/gIfiq
BvvyqodRg+/a8mGxi4w4pQTCKQDJMa3boFbr5nFMH2ocrDj6FLCujdjC9mC2NIBmYkCCywZrhrZr
Nkxz8JhsquOigxcCeYASz4hamEdz/wVFoyRrRd3DYYfx0+6CZfFG7Qqs9sIs1mDO+VTxq5Kkku9R
+COzxte6NJHthiJekfPQ4ASyb/6WqlFsuWVl7xYh/meQ1gOVkJ0lT41spCySYJg7psZtCZWCwhfD
A08X+BRkfzxCLKwoDPXjrZUUKE+nV73eKcYLGymRknxTUCs7WDrgGwCUHSUUDEaCWZU12hvSNqe9
T6CxMLULpvRcZExdqAY6QpnNVL8IF7sx9/8PeFMF5evMQU7moDIk8t7/+fsZMt8wx0JYmkp5Sb/h
xalIrvwLV21a5T5K8dvWTJG3tLARCK8oJjvWBh7lltOs/JP3ahS21Y44e11oJMuhDELihEWB+Juf
9JuJT+llcmXZgPEs9zTOPp+UtMWtYMrECcfxoFVNQ6/CCUcn3txYtHs5PZj3SnFr9kWuxZjL2AKS
vX1Dhor8TBHpKErBQuF0HvfRmmBMSATmyFiJuqmXcf3Yhr9UF/T/gVLSvs2q33tj7qN4B2nvlm9N
3McUY7rIWVXmlheeW4ioSR1SUyp59yTlwDvahCrfsK+6vhN/Hxgi0w9xmSzWI76kJCosVgC4JhVd
kIMk/fI3AxzaoXxeEG9gZuPS/hAp21MHlxDJ4aKHiDRseInI3Uf35FBXYu3Z37+sIzPqkSXGJLMq
fwt2Bd/pjghE6z/66fC4hzYdwB7fuwLS9X88lrVWyO8J3XFfUHPZfQU10qMwMrj4ZQLm1rhcZfq/
SVDjF2UtUEetEox0DyqHN3neiD3udYT0ZMvhqmTp0x6x88WeEIXSt7omalcmy1xPFaWZLyWnG59a
St6sDQXnSMm1lvEdneDRiYxJIw87ov9fFeGiSDBnMcK1KZp86N+dS2PCefC2zX7xNyKZtTGD8fmC
i9Q/yyCw9zTn9wDquU+Y4WSrt16xIeiH7yyruIke7nwlh7UOuWwG2qVqdEMWlWcWUL7XiTkfiski
FlvpFBeIGDSe8105EG19YrJl7TI6S1hD6TPbpBDaN89lErT6N7Pm1YmeFNkt7bU3DqFD5K8FnOqU
LJPuTtIguVyd+92qtXn7CX0P9/wFsrgk7bteBXV0peOb2l6bW4zdB6V/zmiXgx1HWvGnXPbbNgmN
dDgz8t9A6t1UWTPkl0KhdBNieF5QkPBgK6itY7rukf0lqWmMWZPZR8ZCOnBL9ZBb7mPOb5IVWJNi
7MmwoMOXRluUr3RwWGFqKP+xzYnA6CUADtBArIrPEYSyUU2kZI+SnLPzoUhn6HSkCvvfz3oC/ptR
7CqVDk8XO/aeAIoBka9OuahZeoPZOt+tfGSXu19kZBuu/xnzlGLgZgzAK6go6At3IzmEP3Rt27Fd
l7vC/SyX6qYC98iQXvSsv7envSMkan3qWARKqxzPbvb2uw7Hjjefq6N2zK3T4Rl4YG9FnMlJZiYT
OphFs+b1r5oaBvfG9ieioeLKnlMOCep3VJIHS5odXBtZVcV98SAGu2XAf8mT1zA4b0bAJbRoedR2
Yt80IgMc7ptnVfbpXY5XVQ6PIVZyyGNkYdYgbTGq730WZ519b/xL+yZxgjsXCWob5NDD5RI8Z232
elhySunCqAcTMTM+H04xx4BwmgqSkXGouDs8wUPhWi0RJBEPzIrn5Hfe8uMzd8C6qEiFtZ12wD/T
SIknG7YFnloS1IxoBOZ7qrwChJ0R3015w3p9ZXz9G8hsZ1s3H7U/qGsP8fzG6I+CA3l2ZLm02SWH
sjBS4m3PUXlfqgb67pB66jCS2j5z4O+JG3FC/3L84D1lYrq+CkxCXV3wBD2fOhDp9VoRJgAkWabh
Adn3JXQb6EWw+8wrSwFDnINhk47IMo0OzCBQQee3XIoHQPtLiaj5qijf+sk0+yRAu95OI1pMQZWF
Q88NXrK9JZrH4vbeZytBI14d9DPWE7RcJCr3Ei6fiRzERKlLHDPGMKBe4VhMC71Y+pAxtAwuLRYz
Q/aScae4X9x0hZE9Wgt4vVu84WDpzcZN2w9Saz7Xp8HT7L4IqEcV6LraexI6vj0pNRcO5nIKrsEs
Oe04doQzzH0YWykLMJ123m2Vu4fUhlxFTMOh0cJd+xdYxNbAc5I53bHgSf8eSNzLOh/lSyfY1xep
y+iFpBkCzxDayjTrQeBTx3Atbum0FPOVOtXqyzNiAIox48Ctx8zcOSHB7z7h+1cjRKJ3hwcN7QoP
0B/GSdfCWpIq8u9I6655sBhRQeyudsyAcglQ+TEMmc8qcof5Dck3LBDk66oRSL1tUNFxT1SrfNP3
yo6UUsWo2dEwgHBAKbLuTY3HOqkt6HQXFK7r+L8RsIU+4rqrlnyrxN0B6nKeT6yK3x1Rnfg07kZU
jqs0ZZNn2cNMC5RgKC1EI1y+xmfVHQ5OUq9HIlszSDLyGRtv2IWVM0Fe3nLvZKKFTp2Zn2p46Keh
HrpYPPaVWO8UC5+wEEfAqpE7DJkJP3A7yxd1Vy+4aqkUCLW+4qSiWitjKnvQ2Z1kpMs4EVrEFhOn
1R2/cua7qErmLjPom8g1P4jPEGsUD76o215vBjgbhmB2LeY+ITieYpWnxC2vgF3UGOwnrJuFpmI0
z81Snx5WNufY0FksF0AwR4BO3P4fK4VwfkgMcvT/IWVYFYls4iGgpDIC6ziTNAhg1oh2wcHkSc/A
2qENqWyONsspx+k2Mqwu/6WWlygEdf3zhHr8UaMHhRGYYFFKOq5ROuUuPG1mctTloE7u9AvIrfFB
2qHbpZLhYyY7Vsl44Y0WArsh3DsxSz5R1Anogcf7XJEy4UbQgiMtuRqSSE1aL2dUB23Z3G3WEr4S
bchDwbr2u5MeRSNpzuXezaAv3eQAk8chQQsYqY5A3Mf1JI56VmVIYVEgrN4jK2+PKNXoMdQ1vVzE
AD1eD6LV/adUnwovoM+bOtyfoBvf+t2fqATchy9VyrHIRXfxdPEVKAHsVKql+/+x8eHdj67lH8kq
MIurLWa/cupV8Q8LoMPGV1FMVeIvLxV1XjYmdgcZNv6xCfoBv1kaYne9OZ1TIC/+YD9y518Fubfm
y6DJP33QmgF2Qj1H7lu/rRIBNMXVVayqSWBbgcWrMM8v6JrfJz6TowS9f0mMPTRfcepHHnTN0N42
qhZB18Iy3us1/8T2S+HJqeTM66yaUstuvR08mRnDafdehyzGa3RlXBU83rYTWweOtIVpit7hgkbT
zeN/2IPVeSRid4fmZ3XNtPym7PaVfc6UZ5yDc7FQdEnB06RIurYkaqtv2V9yy1X0WyjwJP1qlwr6
ORGuCRnv3q78Icw29INdCPZU9MxI2p0f3GQld51F28L3cidTc+dwUPCiIT6ahc9r20m0YfKlgGRE
Eq0QlC0/F/brdPw98Wc79IPPR+dd4s5DiYiFG1P7M2HZBgyiOuwDPEEBMeNXk7TqFtFX1HYxpLzD
ajHfp/TOA1/o7Jp6+gpWz+REh07Qeh9wC9NlW33sNrHrznIo1rVcKRoHowVWRt7dmuzJvPT0Xx3F
y/dHvh8Y7RHRCK32z9lHtvM+1OZGXo/JnTXzt+NOdCipikG0CfPoshF1yFnd7lTn0/9aRB5oBeSs
ZMrcJ9oqonfsD3vTBE38g76bUuU6X+zYuCtKBQ7H4mRA1elKlb3LBPIxaaOSssMzJGvurgwgYb//
jDA2cGse/bgWNRF2WYN33gI+GezHiGGQYZr/uG+LzdBUggl0JJNOYfcS8oo7GwkNJpMy38QlPCdk
907XZF+/LAab34+DmOIM4J8X/24yUPqQDnQkvWZ9XbIW0hrL58xIKnYXUG+tsdvYhYDBE4vbwjyB
Bv1DSj1NrmFSvTGT/Ur3YflDG78kO4xY1kMW+EwiFyg0vs7sEQElVlZqPqYwIiYnhojBQG41S1vk
VkrrjecWmZx+j3N321khn8Fl4vduv3pNQjDk1dGKhWsjznszNCiVICfCkKWw2qs7jVUnkYhsQ2sO
z2OtB/CLGHFE8douUiv5opRPknJX1yD5P0ooYt9q9hwSmaxFkIFQ1Ttofr66diZuF5guHfuZnp1v
gGUFTdfXbJFStwz5HczS29VOnT2DZQlH5PPffZKj8bhWvFJFJzq1MiwPnKiVA9PlUtgRs7ALmbX/
pJVXif3FLIUIuuc3m+IwgQkmzA+aY53ZSn5beWn2gEZp9h3hY1y0HFyDtOY=
`protect end_protected

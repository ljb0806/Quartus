��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��F��g��9ht�)|	q$�)�3TS�r*N�K� Ў�����5�n�`�Z�	5/�]�&n4{Ч��116��8?�#8�S��S�,�󉺺�����L���k'����9bFi�Q�A>Unc���XS":�~�X��r�L3�V?0�E��
LEڐ�l��𷳵��<�}O	�k��M?����ϥ?8�bڠb�2��j�y3�~����� �-�e����k�^s�̹H�k"��{��O���6��V$�/�H#���Ho�p�튿}s�Vv���_jZ�N!��P�)'��n������������I�@�9)n3���Heu>�oY���3��
(mm��?�drχi��G{��� ��o�k�� ��lEs*r1O�D��I!��ǫ�đ���^�_wڇH�&��BE4����#��n��àw��{k�ۜ-�Sl�A+����W⥈�"�M 3��8�[~5��~��%C���_O�c��a'?#��*G8�3 ���=ߌ����c��E��5߄�� ����h���"���z>��Ƣ��Qe��Ʀ��ʀZ��i��d� ��4N=u��t��(>�X6Q����E��`R񅙮[uo$�����Q<^�.��y��w�b�e�R�0mB���Me��y�\ �N�����]0ф�<l�;bVW0%�\ݶt���x��|0�Lk�����8V�˛G��7H4��k+^�5
�X��hJs���|9�#�-�7/�im7��b��&(@^䞉TI���TI���L�Z��f�x�ׇ-?[�)��iTa�	
�Av8�?�ϵ`�ۈSr9�r�� �l��*�iS��a�IDw���m�	����5 ����x2~��[�U�x���ph� �(R�(�ky�� ���ub�i�1��L���F>U+�9�
V��Z�����-D����*2����V���a��7�s�Fϐ"�����):\�v�T��q�OS����Y�V�K^�o����r[����ņTZ(bŸ3��R�ʿc��l=�_TY;��iA�iA#f � ���Z�7eqĆB�He�PI��n�ߵ�Si��\kUҳ-��$V�yW��v�/���0#�t�i ��)�����t����_{�4�40G�tj���N�NQ�*�~q���B�q��B�.'����=������0r��BDO��H��,6F��nRX
�_=?m���#��e,V;�ݵ�L�3��
Ų7�I��|3�c���"����`Ρ��)�Z[�:�hT]����w��X"֚/�7f��lQ��K�Z����3��Z��S��'�[ڽ�tY\�+(�P�N�����Ď�83�wM�+ $By��t�Z�y�!q� ��9V11�kr.��⯾����pīrR���[� �=�~;~���L��<���m�q�����8$F&�S�!QY�?r�mi�!}��3��(�+)t��XN�k�W��^�߭��zc 7o�[��3݃�b#�*�	�ϻ
h��ӊR�Ӿ�Ol���Wo6TD�L0r�zqҟS�%�&�$�}ӷc��!��蠈x��Ә����x���mѤ�'L��/R���Az�7U[�7(��3c�c9&t��5����]M�*��#����n�xj��k�T�
�o���>\���u�����2+����:J�ow���X��r9��'b&�s�W�ڭk��ح�"�ɓl��3����dm��q́J��L��PB�>0��.��W��%�s�1�^<>��#�"Jm�j��o�f��=���^�[t!��{nk6Z��2�~�ԩ{���	x�4�f-+�;��I�W) n�͉����~C�R��"[�JS!%�N��n�O-��U?/��g1�FR���3J٣�V�AM����;D�:�E=4�G�׶�O��>�'J���eL�k;���_&��R_��/�r]�I�����;�)�����2s�@�'�l0]�8~6�����+�}��MՍ#c�~���!��"��N��,gKs���|�A�^��d���RiP���K�6����˟��_��n|�jt�����-���j(���f*Om�s^��~M{%di���#u�@Cs�鰨<BML̊�5X:#�ϕ�u$`�3-��.���wio�;S}���9🍂�IO�#�2���9��}�h=� 0�[�s���7ӊm���՚9�iY�#1�*f��[��<�"p��R��{�d�ޱp_�{A�}�t�}�?:��1	1�XʼEw�6�&?Z�;lv7�XK�#��X���/7���c\I��K�w-O�2Pp�Fpk��ܻU�WV|4�hmC�R���Q�V��b�+s����h_�!�!<d�R�#	��J�|!��7cR�"���$
��j�=�8��"�^���NXA�ј��9c���
��>��Ŝ�B�Q�k!�k�cy��.�j���P�rT9-e��䒭��R�y��L0�$�jZ��y�}E>&��x��jl�#g��R��Z$�m�5/Z����Ц�����}���N���J�8�B)�.�
.��ثN��� �Î?���GL//���Qŝ��<m������Ez�|��I3>L�3�ε@)��GM�4�mW�˭��D��c锑 �����=�@����7��c'����Dp���&�;^���7C���S��S(����봴Y�G��e�i�h�r�#�|�E��Q�㨚_y�����|��M&V	�H�pZPȒB�c���¥8���KC3�q�{�/�bEk=8m$D��ɬ"Q+�@��n ��N}"BzU�t><{�Ғ�z�Y� �r�|�������(Ϊ�gYvW�g��Ul��,�:~����=mpM9[ގM���ߒ�`1P��~�	��9q�%|��K�������r�ӵ�1�]����4FA��$l�&���^��q�g��w�[�#�Ƴ�ە����(���%/	�;�GY�Jq�*�9
�~G���.]k|};o'�\��dNծm��cfн�xDErQ����1�����<O�eF�����;�ep3h4�U�̅�Q��\��h�l4=H���)U4Вc�P�$"�[ZX�{ŝ��"r�-���#g�l�\]��Bf�^IUW�G���Ue����:=���E��.v��>H�g��K��W�@�Ëp�L6J��J�>����\¿���7����l2*��nTi:Q��mb�9��q�*����.>��E���*N��. :#�����9z l<Y�sDBɅ��	��-��W9��"����� ���2��wmdY�Ba[g� �1�����]
(7Øq˽�ۜ�5�X�'=)E
�d6qcC@��i���f9�}uO0�����]N8�jX���mf!�l����ܘ�a�Z��)�������� NX��j�v�fv�*��?��y5@A�ls]j-�ސc�d�^�3x뷬2���a�q���m}rU>ʓ�ڹ�Mo��|��^�R�~��	��l L]Fv
�`���Y� ��I\�SӚ�I�3js��?i����sA��\�@�I_Лj�����:���/6뫫lW��
�Bz��.�sX��Y'��:����!v|<��l�o����j���>���{"w��>�o��ֲ��R�=k���7�X����w	�>c��Uh�z#x�<���H.����\�Ld���@�R���VR���Y���D���<wy��E�~9C��� �p�W����W�iOV��jF�D�`����\q}"\b�]�\�Q�7���B��O�J?n���P":xG�B��]�goY��}6�L�\@}��-~ڂ����o��j��p�Ϡ1&-�{�Q�[�۔-Oef)D:5x&ŗ>)��d��9��?*�ZO	͘�_���C��s�{6�;2�y^�������"�7��[�[W'��4r���㳔���:=�&�~�Da���ļ�ͪ�\�^U�#++��^H��\�K�Ӭ1)p��I'9��s�MKV���_u%�r����i����-qY����/N��b5Ͷ��o]<��Oܢl֚?��IV�3���ay��f��~����LݦrU7ҕ�Ya�rW�����eT�[����a�.���適��{�mldp��$�7`ic�,��[8�2�K��6#1DG�I�1]{e�#�E^�)E[S>,���O㥹5�%��`�t�5��橥q�ͣ��c�jyE�¬/�e+m]*����f����{��rJD]��5��4����hG{R���÷�O3�2�l�6����@�������aP�t7(FM�0��٨Ϩ��3�]㺒�7�cҌ��[2䶒��=��W`�;�Z��sE���[Kc�!�֒G�|Ղ_�k�N��9r�p/:���mg��X��g���!ʦ��ܿ�;�[R9�
*�X6�܃���֚u�\� ���Q���if�:S� p���8�!E ]vo�(���n�i1�J���0��oL��~�Rw!}����7_@�m>;K�pb�((go����ş��x�^�ǲk�\�t���ޕP���%��-���[��^i_�v��J!��i�Z�.�g1vݤ�����Ҁ�YV�m^u�V�;��_!}g#U���}��?�5�b]�ر��A���h�	k0̅��8;s�4�+��e���@���'d����'W,g�G�Q�]v��w31�X��&n����e��gz��Y��R�* x��3�}���-2w?�~aJ>��/�
�;��1/��{�?2��Q�^���(��	L�b�������g�o[͵�h���R�P!�R�%�:��E���o�s<;���4�.�.z�0� #ԧ�6�4:l �r�[zro+�S�W��ٿ#q�����ץ~*ucSJ���&w���EJ�58�*]h��Rk�6=� ��-M���ַ�_��Q��M{:�/J:}r��ₒPW�|B\����^�c�@�Ie�v7��N��F�vw�$�AY�[��8�a��K#Y��F\f�����{�PLi�g�K����Z�[������Ϡ*%_�Ĥ���Ӎj7 ��8¿�a4�,�l�8�m��w;Ҋ�ظ�b,��X	�n��d;��L
n�����M~Zrv���<���2/�1 {�� i�ik9�d�1�c�b_��p�#��+��{�G!3��r��0�~��*�C��&E������� C$���d��SO1��9�"s�-�b����&��L��M��wF1tU�T��j�����j&��5��t��Jĳ"��߀��.��_EuM������̏�Q���'uws@��ڕ.�y9�?����B7��.׆���憡u���C�%6;鬱�iZ��7������~.��lܘ0A�S���Xq�{H-�gv���^�{�6����P?>��G�]-���?<�}�dsiK	zYۙ1HU&��x�����ܰ�JbE+�OU6�hj��o}��Rf0�$�
[q��Εܸ�XQ|6�G�6LyFl���̆�V�݈�]�s��O<M���*�ck�E���3�w-�u� �ѡn���M
�v��ifImLܲݙ���F�#l�0��M �7��ػ����@L�v�4;Jc�\݃�ދܮ�+�S�.}�v))J�|�=�Dzը�֕�;�n^܊��ju�@Hq�u��������GW�K�,x�;0�9�+AӘ]˭�8�q)=�M�B:�K�O�? D�f%�NU5������8�f]��ا��ό\��P�f��M2@��/��7��>��ڀ0����H�@=���.
���c��+?��rx��S �9��'	�5 H������"�:�|z�w�A��Ͷ��Tuf&U��@N�,3�A�--�Κ�f�h�DCt���[�"��%v̂ǃn���zw�Y8i���J��ƩzRdѶw��y�W3���y@V�v@��re�Ĕ���:]�6�Kե��]���|6=��VK�)o� ���c&�M���vZH&��a+?h�ak�A��u���5�0����hAD��Ь4x��%�i������Q�{��X���M�|��xw�E#�[��䕧��TE�dA�$W�y�LｍCߪ���!9��_ή��>�Kd�&���s���	Z/�L�@.�qK�19��Y��Z���_�A�0���fQ�H#�< |>��|4�Աw%М6�Ը� ��jI��{��Y�:�������,�yv�<ݭ�k���WY
���2�v-�8����)���`*b�'��A'�I�����{z�dmY=l蛟.@&r�aj��-i�h�wB��'����fx��!���J�]�b�L�8����oK�M��O�[lSǌۚ9A�3�@/�w�L�s�R�Rtʚ�[����C)gʬ�5�����W�4����͐�wSFLr�2hz�x�V�CW�p�=��C�h�b=�<�%ò���z�}to�l���i7p�#�݂]�1MK��|]�Uii�ܬT�Ko_�<d�V���������m;t%��f���z��F{Bh|ۻ|i���Xksab��*Q�q�}8��@��	}s����V�r�;���P%�$����jv܏YX�߹�����-�:\��STNBa�@L��0aD<p(�!��Q׆�S,-�z�p�u1#Zc�7pX "d劾o�����\`��$�����K'��l
s�{�y�˂{��X�|J��ƛ���k�n�t�ƪ-I�̂�\-��V�јw&e�T����d"!��΋��#)��o6��ƷF!u���_h  �����^=TN��U�� �A�
��wr��ԝ�=�׽ev�\zԈ�o��<i���;��_`XX�BҰ���g�g�й��e�5�_�x}ʒ���;�q廥bW���?�D�j�=m�	Z�t�w�p; �ј�
$�Ţ�o��w^�F��,R�wAnPF>%�U5�MI����~~Cf�eM��o��x����z�82�&�c�`n��DKi�SX���r��l*�obZ�9��z��^����+�^�e',�DZ��%��Y�����a�~�g1{�
XQ���dM�Xu�]�a��'^�� r�E�H� :� �� �[���� �+l����!�t�)uP�m_)���rm��@$)�؈���㚇Z����[�aJ+���g����@�A���
��0\�ە. @�̾�n��<0��ĹJx|+�>�6��;ٴ���2f@����hB��L�%�J���x`��4���`LUp��ӫ �*k�P���>�Uے�D�܂Gɪ��lQ��wy�N�5e\��SQ? 	9�h��I��y��O���+�h5~��R�g�Qb[�0f����bC_J�5f|��ô��r:���w�Red���E@
�=�%u`@I�,G�j�D5�*;���6|�/0�J�<2�`����Fv�����@��#y���J�jwt��w�-y���"�煌����b�6�wf�*�L8�
�N8�=�%��ƞ��R̮��WB.�Gg� $�}�}�9������?��d�)�?y�2���^ U�j�K���[�vIdpdd>�JR]m,V�HWs��ȿO�T���=�j�m��1�H^J�H@ع{�P23�Ah��D;w���K&'.s�| �n��5�O�x�/���?�Afv��C|5�0���-�^�Eu �$�D>�k����d{��K��
>W�BH��a��p<��<�� qy�Ս�^�ts��q<��O��B��>�WR�_�<2:�����j�7�����˘ϱ;Yi]��D����4/c����(߽������سew�פ_.�����B��D&nA��(g�͕S�$��5g�z0\�&�N�`CA�z���Mxh���2��X�ﺷб���x8#�E��yw����.
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AOpJOnc4maU+qGGfqlNiy4uvIHxtAq4Cbkng62u8HiYoS+jAuBZkjrxdPruF9uLVi+50jhEiw78E
idvQAeEs0PbX/kQNTxOpjJPFAvh0ZyOuvgKfZGHXA+jQsTS/5mIp9+t8SShFIb4PGU9fdg02j6KH
UiLt5/PZh5x68W373DjEYGUFBciwVH0HhlAG3F/KFaIuid/XFMPIRf9JlFdekRhwVOGIi790UEAm
76WSzN+MwfXNtmW/Dlb7ZMeob8VkLS84DdobhAmHWM9GGDp8ifoc/zekBKfVV7l5zH/WQBicfkOh
+ObodHsmEjwxc79fsIpJCsnDxgXy7xrLq66eZw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13296)
`protect data_block
ZlEinQ4vOlVbDnQBeC+bKFGVKtoaiCrCioSt/VOEbGz6RqoOmHj21Hn2UE1Z6tmXuYXhQdq2XJxw
6f9RwSYwDUDq2pXFHlIWHqb2HOeb1fe7fKjmkl9WJr7FQzKmJU5SSAe2c6MFYAC0ZGEkHvaJgjBc
F2A8ifHFOO4hVMGmbzyabBv/1+HnEqHg4fWwmxbjSkCbUOl1psYVjsQNJcG1mEtHKpiSTqLw85T6
/a8CLPP/aHDgwx3qH6gY1e6n1EhpjrCw69h1PeNPZ5VqXG0miJXn9qTvWYL8O6KTUlhEPUVdu8Rs
pOYSOd100aaevDXD/gkVv2n5jPPUEgSu8Z5V+aHjr0M2djURcc4R8uOCZ9MC+YWSFwiPver/0GNx
RiwyoLLwCbMOLXlscnOUs/SakEnfPkKcL65V2SLydbn+9KA2XTyli2v7bFF+a/Vj8l33bnDOqMzj
Re39uHCdHDgwoCWiPiWzOdVpKfoBCHpRCUh3sH0pNI5IwlakqwnXezEXKUxPj6QbXwdt5w6SGRAN
RltM8csj48eXtjZxRAuL62wn8+Y477HmumHAxF+6w4O5I+OQMhVffLkqpU7yMpmSOOvUheg7oYXM
/l6PsQiqP+gMi6Xo0tuJ10js+cU/npLfClRozouAZxjf0ZXipGI52timRAsa2VJEYl8S4LIZ3l95
p2PmBLBINWOqQqeGENSjgXtKzlgNHwlkWBUBWlag1mi7lpdzSEPD6+Md/hbA0Mqbjkio58ZxVk7+
girKiCZ2aBBy0oJbVfXmF4Z8BtvEYH+XJIUECmBvEAmjIZjuv+WXBFo+QmBwVZpf42O6AaHFkVvV
OJ2Gm+NjUsp0aD2x4aNWEkZgioOLYaJPxdgQEWGcn4SjyR19ReBnHtxTzsIIupbOl1wuDDcFTC+T
Og+mmTNZ/q96p7cmRl70roCSYoNNrItHWkl6iRFJqI7v7rle81fKmCuTUlBURN3TVi7hh2toSjfX
gwbx60SBAYyeqJivg/N2fhnRcRiaJflAVzTnfsx962M015pNyYWVu/zJ+A9PxuOskiZ0nB2Zcswa
t2bxO8HAKyoOLXXNDGmySyjJNYu0eetDB7/oY4yBnkUwtrMiBuMszP0NYoSrLjfSj89KPSgTSTuj
FO/2jPQAEpqsdLecoJ5F6dAadHSBwFvicILQw7bqhG77YcXo3sibFXn3mCbI7i3mh+wGsYAGwa77
yK1OiELoxsPbzydaq2L8tC0VMAeN0y304raHuEAv+YknuB6rvc6xxC7Ks1Kq/BlqstqjYloEXgCR
YXhWTOBxK8ZyNFhYDsPGAtfomllpVGBw5024gymb2SVwEjV3VG/KoeAZqfGqWSIBoTmR8QJyOByB
iYEXJcuYtVqVX8u+nqLqTvQuujGiBmIJExJ3D3MFbua7aP+MLELzbucchnZFnpyqjonGfTIQqqY+
Zstzks0ZPYm/k91UaaT+dQS4ikSE1P9npMStuHBAues/rtCQl8yuphgv5jw1+2MEPnlv/uYxeTtc
6XN1urpsZ1Lcr+DQ0/aiBRjJh2MyLR8i2ulD7j2OtttajVNphI0iNX+kKOw4agmdKjeVk3cUIC1K
yzPjO/kTvGT2PDwB5ETqirvU6SeEhrHo62osLNlyUrGpOQnetmddqgRzU+rQjFNkExPp1QRplX7E
HSBpftYWwVp4+sL0lxsgjIQUPpk1uaMymE/WyDQe5PGjgxxp3S7P9A8g277oWjzYW+P3wewVeHoM
FvnNUkxyqNndgk0noNa1DLpmAWbxcsmE8e5i3PJLzMfOm1XxPSbCs+SkkCAsTAdhPPoBSZx7tQCQ
x5wU8pj9OQfMuC7eC2K62G5GdiVRPCrSqVifHQOMGoyCvDS4sOqlyM6cDuX/xgNxX1oGGg+H/F9w
uigY2BTaO5g71V0lTKAyyYeWwCmS9Yb4+0AQsGF5ODcEuIaGLCwEtILuxHpdbmcuPlNn/j0Xh31x
lzngugde3gP9zBYoolU+v+1RJ8Ktxqd9fPCjJF84NRx45F52nAWrrtYxUFpQ9UYX9UXmH5DU1Xi9
s3XjkuButieInOEhedRoYDyD1xNCt4CA9PODOFGK5D2sW1a8mWchtBpq0rjZaHG/ASPVqFHHHDiq
KUzrKNPR6tLvqXBjRUb4jaQGF7yu/zf8MEL7RgD38YiCi1KQAJtRmOp1RMKz+Mr3ocO/naYAHlMY
flK5pv7Z7SaVQVZ3EuWu0lwgul+RhjRYNcoz9jNALKDL0e9k/aHuWYTRKr4alSlAYX9eIXMqVq9v
ipOYXFrMdDRGoboyHiM9y0147tsku3Blv5oKLWIH57sCPMisc1bOysTo7NnZvZ9OysVl94n+TE12
WyAZTYpZmdHxQQp2zbsFJmvafctYw8I5X4gvtPZaYEplflYn3QTfFi/zr/K7cUkGRkVU6fedyqm8
TY4IxjYMPwa34W1n3NshShqOY+62oLCzHN4BGqgYV7RXjYEAI+wpcG47IhJ9iP3cVCfooE60g/aG
6zQLl8lwAN8nxgBckTQJJR/iWQ11LZgCuT+bLDtYqUzCt/2Uw9XRqvLdjQYL9+QAP6O1RkclYh+2
CI7kkexHAgTC0oQmiWiG9JrD6HlRg8+Jg1gCMH7J2Yhqf71Y1V0RINLUFejPgZ9hz6UzwtdFEr7N
c3010SgPvHQ/UUZJgLeykXzaDkfirSYK50bMP7OYGi2k6DXa/539lv2i3b7NCuIC+Z9CQ9VRQFDL
jIxaSMl60YDvBxLIDq98ObvLwQYutlwbiTCTJvc3OuT/+quJ9AK01FXhVw+/6IxbNxTpzgnQjPpz
ysLeB8CBfzZlZMmgidR4ndZ4qQgbmGrp/T+7ToRfexx2qrfPCZvMWBpv6t44GQHJkTDDOLLOBs9U
8Lxn9bor/uHU/O+bHca9VnLa2pGK2FNiKK52xk05sSgSVk6t/zN3R1Qq5/vIYf4zCYAsk0H/NukG
wWhl0JcqHTZot6xDlmttJTI+koFdrqRkaSqR8b3HF3FNB4OGNMONB/sn3kKTC/5fEadogOWBPvzG
dXZPVy5KmG4Don4NECso0q6/yjzgn4KMhVtm5RrrL8lKeGM7DtG32nt85By9ZKxv5Lv6cUZGHyzd
jGcMpy6MsvN8DG0zKh+UrjZ5RhhRjKgxWiqTQts76wtPameJrWC7aYzYDyESL4zzx1iV1Q3mzHxV
K8bi4Y3lTLwLKpPpCdH0/cVFXCaKdy/8i2XNbLmR7OoMz30hUSeWBEhPApieU31FuXO6Mw1UgBUu
D8N+5Y7Q52alQSF9edV3Y4kAXAxElRe+zUTP4YIG900hGmD96f2KfzwkkOU0AOBa60cKmcSWpEWS
kj+Hl2lkMOA/wcoPWi+eWO+cn/nBAH3pI3LYaN55NQXTrE/Vy+0aM9lE1gWxzLqrFVYfuPlaLkae
ERoC6ApxKZz5gij9u2F+vggSYTgFQnE1hKKhBDhgxTvssCY3L270aFGu/PyevLpCA/4JjWtWZ5qR
UIiJ78VCGE9osjDtvT8LHUZLAmNGdEQNtDjK+DKd7e6gLi/4IJusVjK5EW6m7vpFcDWKvy8ANAkD
LTiVqJEUawlC8tW48QVOWc1/8Sfr4Ylr/0T7cVHAPVKOQZvzeRnbkvfn6HUU/PdQCbq78dDnGgDB
nHRKSZcz1ugP9PH8xDMU0dCTBrL4NNOr8Ir8GMfZWK7dGCu6XxK73IfaRlqS48jQ44HihsQI3t+w
jrm8SVWZy90cKDIC0uZ+54q6n0OcQnBGLQcxsDxEyJv/ARj/NMyMnPZU2jZqm5HuWQcngI5aj47Q
b21wQGpbKw6TCMO5hFpm60rYHohiSWr7lv5CaB+py5WE0cNeloU0NcHD+7/WLrttDSqgqu8XHdQl
jAEmWWm6fGzRdS1pXNt7UThEMy0s3JfFMBrDS2MG6an8ZQEgIfzzZejoUQw9Td2zQa+HR410L11r
oe79HzjqCuGXRcC3yO6CYF5pzrFSd2ikEY4/fB7Fr4EVKwsl6Xt9EvFdSl7fRwzkxH37NFwGdoNM
O7PEjG+/6GTjS2F4pUkFUeR7/yLRReLbJSU3k0mtFw+HF7o1A2rFxOccJTOdqr8T5KH7V+7VU9VO
H6cOt9147hzSDlshqoa2bRzrTZCN5sv6behNwCsvXrBfI+SAN1uzRChHAF8qUQK29TZ+KSMZM7PS
77Qp29AxxI/nT3ZEla7v80ixa+SC0PwA/d45DkiUj6CRhvWxXhuKYLjVofKmG7+PLTe5FrH6sZTc
YGMKjQo3Efa2V9UPk9w8L+qe4vYTZo0P1pez4XzC10DaKkRpnbnEOhftOD446UYve897HHVSFjUq
7qNU3EMx0hLC52Be2qZk5CdBJ1QZPZFSkpPtZ8dQPmukh8yCTxWrjCp01mUbfea1xdTxENF8Pe77
KNULH+vu13uFkCh59pLJsRs41E/n2ehEw/fGWNepj1hwllkgjmTEwv2AsC46xJaf6ylbSpymyq63
4n+eSfyFFbGQ71INfqyBBBfOTjbpEov0SWfm4kgJp+LMtExd96mrEo/kj1DinhpGR9Nf3y2t0fjo
Co48XYFNDxDTd3vHMHbTmDkRYE/lXMrmbXa/pyBo/Q7riJ9gYfSQURbq9XgW6XvQQeQjVFQahSwf
uBTdAuq9dupTBRMc0jTUda1OpO5SllyUkmmzXEhJk+yFWvo7DnKDbsRr8PQII8Sg+y/Eq1FmOoay
hnMAFCXw0HzOJ6x/6pQ8q1Yc3mlVdQjmAhAi9k3vrwleDdpuEy9+KDbOqyj6E9t5lR58gaoYKi/4
ZgiG6aMTKiM6MP9A49Sl29PvK9C0dFNujVi66A3vk1n6DUVci+74zZ5GpE/WyAY53R2+4nK0cFg/
YO77Q1JnyWw5diXX6+yOJ3Y3ywBjanTPdj0SxR2UrAeHmR8rA8XQLhmsuUGcAJ8Tvf+BXUtUJWe8
UZ2goJBJSkmu3KNypFB7Cha5gh/9HcW0PmjnBNFZMIiA/3qb3EoQqdutS7h/WJ8tRgQxaNW7Q/Wa
5R0UY36z2GVatbVGrg9T3uG7s1BnsLrH+LQYS9iBkbr75ZSvdKbGtUq5BEDwoYzofAszOTc1pBM2
sIeZdgbHG9ZKo/aXch5SwBfmjPkWBSzY/jZavdZjJs7GkkRPY4gGBpY8hyNijpoACaj8TX7EllV/
CbjVkFOv8JCZNjBObztgtPYrNOFT2ptqHfSrM8Jkb2+Mo7nX/9k11ghvFSMmx5+FQ61b7ifSLrm6
JDgTZXs3UFGEkliuLw4MqjxCiS9LES+d5Pz8vWIlcHjZjK5K9ybT3ZTjemRYhLEPSymYzIgAHLoq
x9Pdp6nqE7V7BDnvlnZ3Nsa0AXIwAGdi0S9ezIoWPuztqBpeNu8gEnoF7tVF4bByZYmubFLuiV5L
U55zeYZj9GIKTDGIAP7caMDbIwGGJ38gZRjqEGaGBPjh27/zgKlzTZA+cbpmFTARGCHpK2hStj4+
1Q9IKwUY14u2qCoohw0wlVjhP23n4EakxhIwe2qYwAaGUBIAzkJLqCcWxOow7HMHfisGN79N2Xnp
ADPqI5oHrFMlAuVaOfxL2ZiM/1wzhn59mEbsqLZFXjaBUJPZLdyjK9jwjH0HfgSx+ZCQMdZN2rvW
P7SuG4UjzdYQhOKB2meNEBLM+MXX8pCWXRcF1vhYBQNkF3FlS1k+yZ71XLU8753CQv7pxRSMaxj3
+ZIG3JwG0jdyODuTwFxLOJIrmE7PB+H6ftUsViJSn7KCGe9aCllJiXFyVwGqzjL5GQTgIWhZO5MW
EYnZ4nlIofBTxR8+vOqZ+7PuPupmvN0NpM2XcNTUiM1m9ZMctAIMfJnl1vECxbFmkQnEJv8HstQU
z6Re+owPBjF5ioen9lMII+Z1eBDf2y8i4oSpC8DDVyfdSC+TzwOkaRhW1KtAyfQrJx8pqBuNSP1o
nzTO2c6EgEz6yHrGL1XvMNjjs1rT1ooU78K0TPfOY40lisHCnwRkj2SjXCELunKm7iQ5CosK8KLR
fyfFkB/Cq3+gyjdh0lZzqUAFgvAwV3qPAWNZ7J4qnAL/WPxCRQBGieYdcEUbEHLjLKOjCbsnbqqz
jCCmOM1/Zja+ddeOR+dPWZp1vA/d8z2m4do6s1AeldgVwXybBRpFtbiwyEWPyQH3sekW2TvnYK8a
idKYZrumZ8O2uyQ/vkgm8kZQBrEfd1NpAHZqZBa1YiwC9t2YnPjc9aN0P7Tkx/EpAgTyDDCDxeaI
k8zSO8BCfFi8yJ9V85bSYCiDB2+T6f3Bx4WFN6jwoxHpjw4I1AveydZronOlMb7R5iYOTRSDCVEi
iF1J/R4hqbP1186VEuHqX4BfKaqyXsCYUCkN0yfbo3XheDqCIfw4UP68znVwM2t/mssqmScPn8rf
1nhKGTQnYREIG4j9WAJpm5aSok5MF4bQKIoYbu+Ik3gmfe38twLSyuELR8zL2mERZ8WGKoaj64VR
bBK5JNRjH9Y81X94cni8xNI2s+hzm29sXbv2/L6TUd6J2D4Mb4QjpcXLP2cxCubhAaCApuEQ0YKW
OzBnutSoDxkBzShCYxoEAww3LIPITJwDG0iJUW280o+pSrfOqzkvaW8TnlY87xwwouidqC0mmLSp
tXcACbeGbZqAA3no8kTfL7vSY3BknXs8QWiRn6TQYYf15FApuoFJER7ZpjkBMSfuy4l0C9VBlgIG
EvN7gY74lqnAP3/iXsLtE9ae1Wh/ssquGkBpqTdU6Aeqz0ptdhF2opUIF88ZhyR7+wg2GJ6HFAab
JQTX0sGFagNJy1REK39ozDlgLS04XzSEnFRL11X2GaxCd9xEiRmh8Tacgj25ukV9TC2S327dXSBy
PQXyVr3H8ffqJhejKtZf/BjtXlaWqyNqNQ3syhMfZRpTv5X7n070BizjQ/7ko7ES1Mc+Eq9dy2ln
JT7gUAoluZGHk9X+cig8AZxLiFxCYGwPBc4mnQmFzEbW4txBcivWUlbNOjU/Bpch3NyG3bnHR89d
jbv8BwkNLydo1uJSUMqsZbE3OfOl0MR5nLxlyswYX2jyk7S/dps3s5UEq98j2WvIlfbMFqIpC1rB
PwViKMsP6SRMnydn4DZig1ynH8fW3JMh29xUXUvhZN5dh44g07hYGoLy18wrdOfp8+DTBEUPZzuN
KYh3RoQejBfTVT9ytqp0t9CPX2BHEAestRemdoWfDVGZhhT+Y3Rj5YMvYz5t0whOGWpCB6L7DAxZ
zz4YLvWPha272ll1zMIv90JdxOFkEhCH3propYWpdwe7UGK2fTIzNrifZci8gWOQG3yoHEqmIs2E
jeEMJtV6GmLc7utEwds2QlwNgmo5wqtWWtLItJ+1X/no5NLURV23HyYjdqBQUhQpgcauQxhcBv6k
+CMV16sK+aaPqn/xZ1pSbzviY9C4Jo3D939pTt7sEvE9RMkEC+I/4ZjFGOXIKTQ21btsZTQQBjHf
0geSTrKU5vR69WzpVyDaPQbeRR9X5xuqHrjJZ41UfZWX5+0hfqmk5nBlK0jj6lb2wMdRs+PmCGD4
N2kAtHroKYUdiaobrJJY5nRUEbBn1LZqISmVwiRx69v9FbfInVARD8QnS/dXuUin/QrjIcliBnbV
n+uzCBcqU206QESLxcBqqAvDxvzYepwOHTCHpVanUNM0rnOUWW00U0mcpR1xhZ+SSYNT1Mk7yBZi
hCDsgF5obH6noqk82U0luM12FdNmYbS/Gh1aCrdJ60G4By/lcv7LSzwxieYMICGWINWI5OZ67O9F
8pFuSZw72PqL+LGpW+duIm4oIo21mKeEA9eGQtv2xMeWKCvHwSd+d79cqNUY/9Xm9DpKUfSOp3FG
bCuwzH1CWMRPTCVuiNL6BeURuKYHWO9CRwbRJ0nfRz0k7g7EJ/Sy4BzgYIghWiDgTO+eOnijc+6G
CiwZT/Y98XvtRY8oV6G8tTpHRYLaiyFe4jNcNyAlxy7gd1KJBMRZPfGPRNV4vDC+iMnl+9TwXPDj
r7I4lXVGfvwM0qDC1iWJleOYUXPkVKkO0/xn/Uv8s7WpVDrTfbyeaO44092jekNS6IgMxciZdUkP
Di1tsV0HfXJ+n4iXTNF8c9sR8xNhGj5sclqLEuNN75rWxTJo08N0ARIIENoqqoR2gUshlqP2WsIq
Q8Y4l9x9rmu2hvb46Jw3izAE6NP+ruZ7DlN0Sl5aSAum+Roj/oaD9XuQefd2qv5WF9dle2UDvWDL
j79SCi+5q9ZJIrrP/66Aurabep4ckO+aAw2b/Z2OCzSjmnON2W41q75ZNrSyrS4vhUs17LcC748A
shKiyaSrgmaaDnwB3DAMIYAN6b7eJa2LgjTZunj/luE8fZQmpJf0h4K/fbwlFgS0mgubYUthhzlJ
f60TT2+9E/1JWjQ07BeBXAucJx2g55kh476Hf5uQVgQJuc68TQcwNHkrbecXmgmU9jpLf+ZKm37s
8ck5Agsxcu9Bo0kajJwJUK6mrda5NlmyH5jKODz7d5WXWIlla7GfTIAPYyx23/uvYATVNOBjkgQ7
kEILPr2NQ7AT/crTtT/qoGlUqYLYvRKGfOsvV4urA47IgICULGwu9gOSqX3B2S91ez7WiBkhUij7
diZaSg1ESAEtPXYIb9Q4qKTHfvEaFMClrYOAhCb3UQM+MBhWoNib+D/qzGkG5BHBt2sgKZI/hYBI
p47rfAliVV09kZiCQvaaZT3p/tdAOl+02d5JpJ6MfZmpmKtA7y63HjcGe7pfl2eANGMo/lfSqJoS
8UNMuS1H+3J66QD7BzCZzzK5YuWU5c0mhsejxQjLuool1SvL2UVE0uxPFy/pgR2xXRoCk+bA74kz
kOggisF2L+MBi7jfLyfnu/aiQLYFmCeQfWi+5y+PUA9N/f8Fe/bTuCaiW3mP4zPn57mp/ZXc7+qd
zUn8K8gR4czJ9J5HabGIg3vQeQA+reIvT6HkFgORqf6AHzqOe0sgCpkwug4s79nFsLLNLabfsQQX
NJN1N34fWQZuAgbB1gO1/1TnjtjgS63LHP2FnwRCzNjdfkqka0YrOO9X/Ji8DWOLBFdCiEFTRgkl
/ddE4B0+JDz+xMVVg6B2owY6Thlado6t2eCBz6ux8H8RxgaMNBJSP0sfYaCgt6+ANRgcbcX35VRg
IqaIe5BazysXxpJKh06sE8KfLq8BT05ohy3BaE4NIf9HwajpB8VRtjW3Z8kU0/xyRupe60cHYO7l
VnM5difpg6Nr/BP5h5EDVqW6GCmg/+l+YYTWAIgmFozs7B5A4j7xmo9JHduyW1eO9dMkeHDBWPp0
HvIQjlFQ9q1/GVuHahysyqLFdSPGVjbXwct5HCFgkhTxqWSqlef5tB1/CkIYDvM9HnFnj1NvXLkg
RcH8fgp4/W9HiIczlQs4Uuv+3ELlPBgT0lI1RZG96NH93gfSEifJ+cMllMWWjYSHCkSXNL/BMQ6G
qKSTZ6hPkcLz8n30AOmAi7Zu/ktjtBCe2raoe6vApKM4DsmSB5gVCyQjd9aYxbcpHV60nAmRlBBX
ZOay+GwK2R5oahI0Q/OnOiH2nMZ8t1f68Rhf0Hs4oQs0zRx09D+oiyiJ9prTX1/VcpvxjC4F7Tph
oYj0i1mDQfsi0I27vvEis8MfeJ7b3uwIM4ZyAo0lhebqiRrGd1Xy7+n/x/4uj+OMZvT/NIa3slA1
CZmAGJJeOA019ffn+p6l78cGyfhiYNFvkcZaeR7kSgEqc7Sxwmcc6/B1bckwLltTLb7PjLSfPFwR
lsKGw90bPtSW9irdemzmdtY9P1/aSTuAbv1NOtyguxJBtIUPbz5/lLIX6sk96DwwBRA+6jQXo9JE
G6flZnGePFIDLhUZA0C7A+Ss8GSWp+F7hk3eiRrb/s45O+iUpO3ZybJVu+dXMwkfcItDvKMgQ78W
8iqHKaHEGyaAfrkytLXnueK3E5zJWqux3IGCBdBv6X7Hvq0qJwfhfNdz7j34T6tOUtLZ0Fi+f0kt
K9lXIlriik//Q3pNRQCUT5jNa89xULtL37mDV0CXNW1d/fyKcWG7VRac8WD+6LDPDcEQtadWGfjh
EdcFnHrXPutu11GJiGEe5XX3q1P56Zr5tIw3s61WMKu/od2Kunm7z2DoQ5WqASKcbdDooHEyW5LV
pTfVD0J/mrttQ1cy/wUUSZH/cLNn4p9azyKlwAf8AIpuoU84plhjBxMo+jdM78g3aDEzBD2iT1t0
MRB7Xns+d8TNU8EgTIl5G7a8GusOAELlMufxxCgzAl+t4RK+d64Uy5PvtzbMHJlc9QmZmnnix2cX
z4+AXO82L+Tbyb118Risxy4rE6S37JsrTWI93Uv8pBUiaHMjroWqv6x/f3/a4+HBLiph/qk9c+n9
dXvr7P7I9Wa0Q00wDE17iRzxXjOs2lkLW/FzE/O0ebCIwIDD2ifK+TfXZZRaTuNr6QgDdfF4Owvd
0kVa6LAy5+Y09KXiAN0FODfHobB5yvEq2KvZqE6gu/lqOipfQyrMEhPHfvTvZ6dVmS1g1q94O04r
QPg+YUMIpUD2AAfJ0o23ZQZldNyenagqNycRNo3wC5Ff8sHz0ulRmybwdjewe5Sywrvn8lhxAqs5
OGx/NwG3OFq5c1pzGsvJoGoBFlWfUyT6c2fIVti2SatfhInGfsP2sw8dynfb+LkVKJmxoyx88KKv
kRL4p2OS02rRA+OAMo7WORwWihW7SyEyGIWH6jv7VBaxep07hXT0oxfmDdsa0jLDgvVRtuZKKx9s
9vz4s8l9YUgb6HPlsR/izZbiBNH2u3mKwrwyPzBcO9G77KT2caus4vrfiECGShl6V2G3M8MC5BE7
tQ2bBOnuQF3L/4qQ5ZnumIc8FKusmAxvBng0rM79+bAZn7xi3tnTsHpOa3dnB96G8wubZPDPL2Gs
Nv7ge1nsPNmaYvDWNlSKUNgbPb1stYAlT964t4I+Ns9sWFWDDB6rMWoYwiZPlN35Fs72TkuNh+1j
HxFXxeJEoV8G+n2rPAxVGl86GUgRZHSlrLVWugjgjK0VWG4D+I4PBPUjnF/g8SzVJ/e86Bvgv3a4
Bv6y4FzZY0qmQdVHq2wFGbn/i4vV7j3TBbgoBR7dq89mbE32XlXU+f03kIYGbg2ySfpy64KLYGnU
Q8R8gENsmvrwRMADjgTnsai05uMouezeT9uN6wYCGitrc7bkpgXSv8oijZkEuYU7pdjJYA7O83hg
DFv8X/QFKU1L3kkCSWL1tSjLh3ctBWda+zwKQxR/xVgcVwixJRsIyYirQAM7hTNX2nED6klcMAJn
qpLNs1s9geZDlXKfqpFl7kKmR5ERcF+qH91fkhmXjai5Z8BW99H7VFqD5Lobp8dXMfawdQBLxibs
KbuWvQxaMRpieu/GG3svYUX6NPQ12CHEMOATrYdAjhHAQypKCNby7Nwb/wz5J6/qVGuYPlYKcJzp
hs+l/k5iEiqMNvg9B79IiLgjvIaLCOrZ/hqo9vf/RLHz6TyxT4aBeSKDSySJx1+v0GV//XH5E/Sa
nVSaboFQwAGA0Fd/P0bG6UYv6u41c8stx5yDmiIThjq+sx/PIUWl3AReYm0zmSYdMKFR8bp1xnZr
EgPBnrDBsi7pO00LGAhApAyQAyU/UyujGgqE6S9oVzCcPktfSoreWzosKD4C7SOgxTf9qzoKu/e+
aJa5DGw9bjXQNvcAxA+9b8TvPAIW+T4kWNrf8dg5WSVAxf1i52Zuh9BVz0SiUEE8jleGMzLUxres
0zFXYJizG1v0Tksp6oqDsk8GqM6nV3Z1luy9csr6mewK0YQ8dQP+FJdS6LaP3gFHDXJG7dzel9fB
2I4LWUpXrH8rwEQbSBabwcSE8jXDp5zhpZQ6JQwaAiMkvRbfZcSSInXKwoMvey0+HKWA8j9C8JSk
oc0SKcLZM9gSbUb6ZDeYJEPw8x2T2HVkVbKl4DWgQTg0xlEomdgfWy2w1KxuyT+wnK8pGgKQb+Va
fw2KNF+Ai2EOF16KsmY9fQWbub1Jk1yGb9sAeKJ1o8PM79G30+zsi+ThFsOKB/peCQhxN0yKhzgU
lcQFOgyjXcx92TUw01O1x3PxdWuK3HdWVqWl0gh31EuyNJVMkTkrI5gJnW234PDy0jGaUjWUa2Os
9Spj0yhDvRC7FiPpunE4m0Nn6snFE5M2Z5Cbc/qEZfj6QDr18PEq+RbRIAXWfTF6gL0SQ/T7l/EY
AL7vHkgWpQEu+4ar/JAnpPy1WYVxGpEq5dPeTvIDOO6Iy6Oo2TUbAMC9QoPMVy1/WpQvK3XWuSFg
EwZ+SAOMDBpxUAiQD7XscCwBzAY7GZBYDeDSwapK6/KSnSUdW3FRdiuXJ1neqClDfOV1d3ox4Qyl
sL6ijlSiJLHKys9KlxUmH8nBZtQYDSKAhnX1mKL2Eoc3/u2SwhwBOPgSqTc5edu9gDYCawm4tAYg
d6RQGth9uFli+FdsmKQh+xmVoOnb/WdXfjMMaowFWlJX/Cyr0SxOQL8wCk2SaYX1rUTGTmYrLjUs
ZU2E4FuoqGpcYAdCKKW5V9tonJRd7knwuMfu23jd8B3mCLQROJ8BJGimygXv7r7nztMAeJlyZMse
RVVFPEvtrTeL/lOKaO+gIXGtek2Cx8VtGqwyRAp+bmeU0XA3U8euq9HEgvVhAbC916HXy+6pAgKo
9ANgj8fZjOKg4297jf4fS9/BnvkVHFY9xB3/wm5+hTwFtfKdiRXN1F0OAjQNioN1VNitJjsTgr3J
/U68FQCX+5l/fX6W2RE3p+OzinJwrTi0zNvmqgoCVD07yotAlz3S0FiMaM9aVOAO4tKipFmclmXp
V1NuSAJOnDv/Wy1R+nCleT4Ne31zJSC6iwPjIawNsBcodrRvH/9K7WpFQX68JsFesOh35sjDWJPl
Q2QXDWwdjOB6CJKQKZF5sgVgGDy7wyh1FxMzClmE4yuTylGM0GmD2Gom0xwyThWd9ib3cuqKFmbI
E5KnM1FgaEeyizinj0ET8aJBlSkXEzFOOiH3IIBg0+nk01lp7m7z2hMZTUMNrROfpuBJfCK/AGSY
gCoTBcDlU107eh2Yi9XsWtSjP01/4gpt5pejT5l6f9AsUimiwwcMBXqaWiHmcZa38X/8TKtn16we
yZrfHgsK7HR1UvaDsD9yF6KxXgEEAxvrOIOKoh7QdP8fxCDMncdmZvA9zTLPYxJNLaxCBnx7orso
zOIoGNhIiW8B0OK1P/dvF0+3xVyrUoqfftc9n/PE98n8Sj53HqDHAzk/vo1i3mOiUfbRthXsBBo9
ZJTVEw92NsColC+T4P34XFsryONGBWj7cfSqlTKtBhK9lTEnTE2BlrCnxFFRGw9ujgX4D/9HLhpp
G5Mknn1KKWFECdGgyYD/7rIPu6dj5nfGIlfJuuIY6YwwMVNgNvwdA3o3AEluZ7IjhkctVYV3VMrv
MrYVQPF4glFfm1atdY6rNxUSsqG1orrsUjb8U8j5Hw1rWMx3EVI508IDJkZzd6sUQ6cLNmbSycK0
BYrnZ0W6XFPR5z3zA8u9+T3Jm+wwNH4BqMGcNPMe3Oxqkal8rzMfbFLEhqlKwX8aDXC8ZSmTyiz8
vlcfVZKC/F7M+AzOUiuldSFyT88tr6q2NQlukHp4O+SmAGQK7cu8NQMNnEa+UAjjce2FUhmUAP3j
7zeehUcqoQbym49OY+Y55rDdjRICzMH2nPJMpIbGHXTvH0Njggt/G8TK1+G5IyY0qDXFHouTixUS
OBdzVnkSFwfc/096yBPh7EXD8iHDcnLEM2aIFPDYwkHey3jfFVmFdxrWCgV84E8na175hez9ITBj
D9LsVHH77dRODWpEjvLmGPH2aIaDirIz7n00URtpJ/Mo0UoApqWHEuAw3pYiGzmRp4pKi/VlIN23
fWEn4cbLBoDi+UANlr4AFxaVZtFiQWxDax4m7cuMUYL60t4zSFcLr2QiJb0S6N7/NU8GPNLuAmHA
e90khYGr0pjIPwnxV9hUaj0rajj4QAVA2vvRb86MNqQ7mvv3QNGRlDyiiWsZUeZM+SOfu7dB5Zgc
lJvbWHOpCEhYCrRQz3A6dEBslBT4skFcPMRddRJaffXfnLyI/1+0hKQm/ppSPcUTwqhT1OPZgZ9S
PppT0IQ96AEtAoJ81KKj/ZqgRtK85Hn0U9TKneCrhsi0VedSseFPhMptPCqcATdhdf/ZieJWqyjO
dddRD1hG+AamXjkFnbhbAKCb7baWEIWMrgRCulIiyqvLFp5OpnsWTXbz24NWYpllxymzfxBrQg0T
6BQJy1R3KnI/enFI6xg1Rxy8/gBAUHkYiFkI8Vq0wFNpKGX3egnJbNF7exxtW+gw3JtRI2wOqcrF
WuBd6CzSMYSuNyjZMtcxdbDS+yQT3ftF7ZGBitoxixABpfvqTPT302mDFla10NxrfBkkUQdAbOw9
+kI1BhXO80ljbFeCxpuYfBqixtn9+mrRtvtBoCHo4iZHBAnEH+poMmhG83jyT273hGwdPNE62oqB
lOUfLY6GQ4XMauuY5oPejAnHT6ZCPOld3xbwiNW+LzGN3YC/WaqNaNg6HltmagvdxVGZodkPaZuI
xfJRC9NsWYaLn/q6ziMO9mfe3JSLi4C90/n0pSYOqSMsWnNGBVtXcZXqWsDodpyTxzk4ANfVsVuW
9uhaVvG5RkYY3FNArNI3zd+ZgrAzCNAPzDBTPkMLlwcuXGx3qYQmbIRCdKPCkBiRk8l3SnV0CCm/
yxmWl8Fgh+AdGZ29hDbSKteJ5IKdC3W/lfQik5Ehpe6eC9TdOB1w9cFY2RZDE5kKrNgWBQkVt/n5
ZJ57mP2RMpS6LjU6IZV7DJOMyzj8EHSIY3XgLHSpfQC3PwWTQKp/TIGRQ90LMqvQBaRTpM6YdQvF
VQgiMGAneeLNEGeBqYb5poaNPXxpIp5Ns4an3AwUIpNfW8x4Z/QPGRn85ILBW+E6kPcfu2BYSTzO
j5UXxCBVmP48hGs1vyVj82EkN8gnH/MqKtZvdmtdNfqPjD6epeccbJbnfFRZexYYGYVF6x3gR4e7
A2gbcXqN82YizJC9z7lgHw/r2PFegIyFR20Hfx30aYnI8c3gBKmfidwTg9A8Y3eE9rjrIso1ePR/
Iia9CsqHUUzaflAy9aRTVdTg7IfKlNdzhT4D57y6u6InfpZsRU+xeLCGpkMZrPb+K23foVNhhX4N
M07n9lnzNz4cLuW0U+qk0u7Od9jt3SWirahuoUub32bWzVn7qwiUXFKY9sNx1UNHSs2DWEjvYhZw
DO6Qrfaz9mtiJ6Wf4O1Uhrt1mZDyzb35CS2QVjq3YngosrzGPvnhCFPrSfTKVRYe/55yV/RAD/px
keT06qHu2NYBuGweiQomgrZCAmZbt1AnG2MP9Anzd6zgdxE0eH75kK6hLe+herBZlsRYbtdf3q0k
ZRlHoUSHNnL+itKi/+96rdbnjsKGuJBZLdHWqt0RKOGY+R0eWQoELPL9KDKQ0d9cdk8yuKz1GD//
uegryxzcS668jfaksXSuIqdRnE2o+36ai4CFQZQmBmaAcJ+ocULkbZc41bLy/yA/QMdl9NfMfC4l
SOrRN7fJiZVAyLBOwDJtLiUOCWtV1641YEKqS84xkuXpm/0zCw/iGog8V31zpRvIKk2Yuk/FpSAI
rsdZsvtLHOP0SWccEITFxNc235+WlWEtpUc/RQ59wLS5hf2I+5AGlTsnkxDBLyzcescOdTlXiqMI
v6lk2FoIWqwGKluiRLCCW1rmVU4hyU0IbJYeU7R0O6KDGpJmt78vSTmROTBHoGH1NNB51pOVo20p
UooFeetgKHn+c1C/TPNjR4iV/9II93VNc236EJcr36DM+b+Cw7RYGqUDt2Uql/mONv/OQuAA+Yby
KXcPcivpRe6D7JyDX2xwfiYRXPv0p1O9SQ/MyQYqrJR5IZyB9zjNI+69PpBih2u9K7MyPIrTud1j
VAZIJdRlhT4An6Evmo6Sad0jEnDHYCiZdgYQ7jvih31kdCvMEaWXPX1HMCQ8g0uiNXrLwI4xpx2k
XxBkN1JyaNL1CT/Gm5/zYb8lqY/DcYRKMmuAOZ4Co8nne7dJPNqVci3pE1N5cfn0+qHIWxyPA+N7
M0v4O4VYp5X+xps9Aap0yvWhgCnOrLlySaerE2t7tluFWEdN/weeTtpJYIYs0eMR/B6o8L3f8oxm
i9DP4OAGMlj6k6TvSBp+lzr1OzchoAg65HaZ46iErbj1du5e9DXiZoXlz8I/LQdiL2zQptNFyPpL
1w2/FSSD9bhUXVrgKqtLCI+PzugRqt+PfnHwaboEvU6Jy+N62blRYYosD0nlvLMxJzvFh9P+86ao
EkXQLZ7BAfywJ6pKv5CS6y8CTOLnftyFsdi4NSBt6+mT3voD3SE5VBXRG0z+r4pqNPJjwkyYxeXx
01A7CMkwqVtITm0urtRXsxnUkNjzIxdJcvw88i6GMLifKnONmxYgRZ6HoUJi/OWCpT/a5gpU5EH8
BhEI+ZmALIulE3IECVQZqnh6CiHrEGCA8msKqeL6KB+CkYizl8IjZ3a4HeYmku8qk1YrhwbzfVKW
OyDaqXHnCMbWKv74P0MhnCSMlnCC+YXcTjImthZshJYgIGL80YPYpHRsJ45mCefnPfyz58u8W0Tj
vQAksF0tzVuIUsrVj5HKDKSgX/a3rss0d2EtZ/VDDyk8ViI1sq/IMNcVNz0CZqPDgO06yL4pEb9g
SMf9Phi174TpinnTyQtii9qhgzncuH2MiYJSaZib1LdYKzeA8UedvPNRDXgbEanKZRbp2FtnOooA
bEENu2P8op0DmAlZ0rlwRsFj5Z8AQDhByynrKyCyUxhlhs37DZBfCLAlFpN/Iixp/CCIuGLpCyHj
R5a2Opzeh2bLxtr1faMx0hqu6pQxcmwePTYSCUinju2JMaTIo9BqMauAmzWkMxtCszbFRKYQ1/mK
arbbCsQtxYLUFzIHUBW4NhnqUF+fv6HbTn7oBrjEjTBVp4eC+3384WtRQFcRFPPgrm8ovqolHNne
i1u9LwGn3uN7YymxaqUQjjr/W7eFmHtVANtoK7VBRB8mCb8wF0lGiOAilEKx52/O2P+I5UntqPJ0
IFuqKr9EPnGbcmjdm9ZB2yuC6VLmHG/fbpTazzHUyaMB5ZnYJqLVDucHTNwBK/B9udQdCydVKQO8
b0ZTF0rCAWpKBp2d53HuKXmo4a0cALUrGkseObLY/7lyVI8CJ1l3HEu+BrfRv+4Ks4ec+3rkkSRY
iK8nBD47oXzP9q27nZ+1OkzkRbayWMr3pJvuX5rOq1Bliqg+uDwPCMYFdHRJTwY8P5GVMd7zIl4I
coVOOO/aNEQdRcgvl6SD35UXDUWPTA/GsXxC74fAilZ4puWcEqBY+OWMcqbn+AnRq1oaqvF6RTWC
9Lf/cMdaCgAYWwHhPYpSq0cpGwno5GI1NVJgS61Dmz9dMpsBDIWYSp3jdBIsnsOINs3twU/BajCM
7MA06wTTEp61kYaiFztXOSSovSgxKluB+VmVD1UBlSyfcycE5PlVWU9Iy5dlMT6s7wAua9egEArt
9vlzeEx4w2mKq/ciA6gbmqcxuEFUJFoJqMALmba/9+ICigWjQNrgWyzdne8+6sRFFZHI/CHlIDAa
HDiCcra2JX45NgIUo/yHNcZt53mETxBzDBvXGXaEvmS95lXSYd4zXrgFFIW6I8cAf5u7riVaFNNv
LdyZ5kd6ppYRXptcQuL4nlGsQYiLa/VwIlNg98G0H0wGhqfcI6cobfKXFjCyp2TLdRLErcnmnlMb
mWa6ypmK5NjL4P0eMyPd
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Ym�7���7.6��u�� 7�(n��^���hg��/��lSJ܋u,B}<$1L�=uj�H#j�'b�!!6a�i�.�{iq�^�[0nv��������䡱�v{���s��I��j�X�+���J@�ԝ�5A�un)�H-|���_��D�y�.����B��k���CP�CE9R�ѳ������A�H/��`/�*K]^:F��6�H���*�����j�?&p��`(^8�z������ӧՖ<i�j�Y����Y�Ӻ��f�:U�C�Z�
�K$4lF��uvD��ZU?hnR���G��!�en�9e�3�k����E���`w��]�i�����Md�f�k�{O�ٵ?��԰N+��*Օhgʨ74��}-�GF*K��o]Q���>���P�, ���˨u��q�&]ޣ����Ao&����c�Q��k�m/.�Pt�/�-	�X2Rz�a�c���OU�NU�פ���a�Q2&��Ϭh"��_`�����>�b�
D.��16�P@D����yF�t=�];�T�̿4��(C���9�� j���U���S�BsJ�y&����L�d������������(����v�n*�1�1��͑b�C��WҲg�)A�^͇�ј����Vk{=N̙��o����֙�3-c��_�T6PQj��u��� ;90�T�H���F밃w�����ϦF�/ʘ�*�ɣ~��B��n@
�tGc���ve��)�k���´fS�z��\��0޹OH :�#��� @�F}�SD|#��/M�*5��yۧ��˖�z�'�D%�D��._�N�i���=�Xhڅ��B|V��bE�t�b�#Y?���U]�<5,�W����P�S�E[ݭ��m���2��jS����M��	�!0֜��kz|)�熡$���Fi� ��G�)X��"�C�@���,d���⊞~:�D-�s�߫��Xx��F�{��-S�麨Knx���BN�����KGC���l�yFh���//�>�{�a��,� S�{3��v�ϛ���N+�c}�?�YJ��~��:9�~�h��bٚ�:�WȲy9r%�43?������)s�ȍ��`�!r�N:�=���3N=[H��	.��@5 	B��&�-�<�^�&O�$<����^�L.�D�iK;�N=9�����:$-:�A�	.%�H��&[����D���w�78k��c��Հ@e�q���+���S��:�(8�NrǶ����F`�V�C����섮|2�¹����l(��~�MSf�v�)*�}�@� 6/��C��
,�%Q�����n���tx�A�a���[���{�PYa�?8:bX�7O;soۦ�T��t	���E2��Q1?|y��:"��nϲ/x$F�p+����V��N���I~��R~���nX��(H��$,�h��%q�A֢�M|�����1���ݩ4)n�B��f%����r�j�q
��eN�4�����R����NV��/�@U2:����i������E��9%@ߎ4�~��P�WeN�k���*u0]�O�2p1mw�gMV?�XF݀���~�Ѩ"��f3��H���������$K����u~/
C=��*X�j28,������?��, �c�zt0���P�\�(��^��&�n�$.$F4���/����ߑ�{�X�0]�)�m4T�-�o<�yt_zZ���
�՝�}���umʂ�=P��b�*x�[#/���{-�\�oXEe�+�R��$��6����	��.��,�\LMY��%bl�&1\��-�iX-��a�L�?��E��@�
�:��ɑU��>ui�Ţc��T٘��ǌC�ؑ�'}B��A�T�})Y��mlb���D~�'�N�u���ѪPp�Y"7�j��[5��� -��۱�)r`�d�J��F�K����}��l��#���ε�t�O�ᑾ��Fu�a����k���!�[��i��ʦ	�@DG�fxm�� A�O3��74��B�ID|5�@��J_Kl�5�.���M�:�	�	7��m�|u��< �5+�
&�V�����@��0���~�������-��r�Y߽�jV��΂8&�r{���(w�C��	��s k���_2��g+����
J �Pa_���t�lMhCDQ�6K_�8�Ë�:�S���`A�7[�θ����Ҵ�}QH��DpF�ޒ�ٹ��fZ�.�̲�n��H;p���h��9\�a�����6R(��!�L�������b�ꈀO{�"��?"(zn�n��}M�n�
ɝ2��H#���e�G�X��U�K�<rn"�&���?�NS����È���zR�%_�9�3֨q��<1`Y{�5.}MC�����W���8�E�v5+�WM���9o���J�B������ |C$�Lg���y*H(�/[���5�R��$V&���U��'L3<��fF�&���dJn�����Z�I�3�~R�H�H.l�`>!B,xLa���e�d�5&w��(�s��\��xd�lxL�y�BL����
"Ğ�^�}���f1�����8x|���*f�tt���4։�3�p5�t���n�ԋ��XU
ǭ[�������f~q� ,&���Q�����8�/�9
m���ö|M�N��{��9�R?4"�`x�U��$��N2�3U�*���&��w��Oa2�~6�慅���O���.�L �#M:������@�>˖;T��F[�,��a��.�䛚;�M�\�j�&�4�M���U�|p Dl�����d���R_�ac�pڟBa�v,i=6�>J�Z�Q-�`�%`��^�5G��Os)�b�c*�~�C<ŀ��wj������h�~�����"�ET&il^�$SLH�kK��Nb�K�E�Y�S�7 ��83Z�L�x��3�_�8gn'c�0�yT��r�f�շ1�{�.N�c���"�������:��W"�c�� .�')�
��aB�V#ח�d��(e��d"��&���O�L]���@&�/��p �f�mX��Bmf����$���Ii���b��̏\8R �@�����j����vB��,��z�Ƞ�|�a8V��"�|�=w�xE�wh� �V�r{�w���w8�Ǣq�;t_���h�<&yX�z5�������_l��,���v��Wky{v�Q:��yN�Mo:�{�{f�Ux��%N&�˗86%�
�c�t ���4�<��M�y��'���
Ϙ��u�dB=����uj�W�t��8R~W�VS�sQ��D��l=�N{���	�0���=r <i��.Ǵ)t���s/#S���;)�틻��d] W`��2�n�Z�	�q콚���P��m[�6୿� ����T��
����w��wI������M��FV�[#Ņ��7���I,��� U�=�����TBM�Z���d��	k9�m D��j���V���@��}�U���X���ۍ=[I
@$�(��]O�F�ma�v1_�g,�����v�4M�����h��m�X�9姧��9����C�:g3,�+��gDcuQ3�2�ޠe6o�%�A�|sS�h4���$:e�g���m{��O����G��"�S΍�&���-��Z��`ϔ+�u��wt� ꦳֓�fv��E%���.dl����v�G�n�1�?,bJ��4�dV�Fd�N�O��{�+��'p�S�'���
=jú���.����^�m7w&4��������v�?�J
)�Q�<�E_�C��vύ(x�J}��%�A��(hd@�X��j�258ذ�Yf7��ف��j�v�ń�8(��^HZ��nE�.�@P��$�/���!���6��hX�����A%y���������L+���Z���c�$A�R�ύԨ��ef��o��I)�����j���,�ۡ3	�_��GB8Ҥ)R�b�2t��P^�Ҹ����mӫux,E�:����3�F��A��a��:2~��jgzp�	p$P�LZ}sV��~�"��u�(���n<����ܾ*�E��𶥈��n?V'&bUi@Y�T?K����~��'�?�6̾[4�!�|y�#1�)��6���Q`��ػ$�Rg~T��|�j'��Yں���u Mt�Vg���c0�&��M��6��G�y�)�e�;cM���&���cwq�������h~��Y�>S@�,N��D�������~�k񬟧�%ܸ|��Q��-ήq�i���ZNI��d �$������f5ۨ��]pZ�:�x�Fp��OJ�zױ�y�B���rO�CV���,[�V*���\�@��R�����ɲ#(�Ų}�R�o[�N�,˼,�����7G$f BNT�b��g(Z�l�aN��g�A�6+h��u#F�����D9���	K/b�l��B�F�=4��h'\�$�Y��y܀kS�>��m<M���HHE�blJ�ve+�,hC��<���wC�H
O��G(�Nr�]�pJ`�,�!���y�%���B$��@��"\"G��٨E,r[�'�$��0�X�>�Ajy��k9G�!���C�
��-���0�2���.t���S����~sO�藁P^�'k�:�?%���ϾE��V_^��#��t$Vu��XP�Z7�c�����Ԣ,��'�++C�y,*&�E��T�	�ؿ��k��J˾:%=�O�]�B��PR���`3O{�Ԑ���4����|�̜Kח()��;s�6�m ��X�h���W&��jVV8��@�����O�c���y���5���ٚ�˩�^�q+wD�ǆV0&l�Z��2�l�3P/\���e����q~�ǌ�r*�Ċ��ڿ�=q�Y��O/ؕ#Ȁ���!͋�#I�N, �	�����p�l�4�,Q���׍��c]���3�&�lApa`q8�])7ۤ��=��Ky��cG^!�XB %-��E�.�N�c����{��iy������1r���&��}����%�jO���Ҭ�P�˽����ST��dV.�Dg������ފ.�*�Bβځ;uI�_���XkWK�z��c�	;���CsȎ�A:�̫��4���+!�R��1�<�@�=�G6��~�*�Q.�l<Z/��Q|�l�C�[Y+���-�{��#oeC.[T���Mf��B���8p�_'����]s����o{��M={�M��CV�pؙ<d8���f�\�y����|�̭��Kz  �&�c��Z�ee�"T*�&����]H����x{���(0���H�ke�96���hk�%���r"�%I��X�i��e��?ߣ�9��}Ӷľ-NГ���T{��PN�E��Rhz%�O)����s4���E䉌�����S��K�}���!��|t��&f9X���A�F1�j�!2
Wy�:v��9��Q
}4��*�xäJ �nQ80��r��}��g�V��U��Y�C���la���bd���AǤ��ZDfp�&fVoB�\�R�9Ny!g*h� /"(��Ĝ��\j	,��5��3�K��\8����ay�m�U�n�G�f�$�U
�Dc}9Ϯ|���	�~�m]p{�F���i���&?85q�-��V�����A���ze3=:�D��j0����G��*Br�ማX�*f|����f��ȸ��tg)B8�����E��@9���2��IUl�tYR9��ڮ�~��J�쁎���х���1���VM�ա1��]w]��SY�7&�KR�I#q\��􂐵�57��-Ɣ��N� IS����X��d���koI��f��q�&�ѫD�ө�P^n!FH0'��Z�R@�f��'��Vp��H Eعv���ݶ٭V����-[2��
|��`0��C$�ڢeU�
�>]��(
@jM����K��n����"OƉnϼjw�aB�1�xxV[B'�;�p$�&�L��z��6�]��<hEI��ڕ�r�s�|Z�����8*�M���"tlE��%��ȄH�!����c=Č��i����Y�k�1>g���K����Z����j1&�w��m��OF--����~Sⴾ�T��Ž����b|�z .oŕ��!`a�/�aĒ���L�ѳ��*�y�-�s�g=Lf�~{A���
�������-�:��a>�)A��\���h[mi��s-e��䭴�g?��w��]�yz�"iǟW����0,Ֆ?���(i�M�'$#��~I�w���ro��;�����ǖ�]��� ��?xn������w����/��MS�fA�R�1/��>+�kF��E�����k�|��Emk��aU)�</��4P]�<��b����o�y��|쯻���p�w2�N�o]J�qM��
�g�X�~����7N�p�1�a���$��W�,}�Md�.�*�'&s��O:��%i�sz|�m�*��m@��c��D�'}<9�yp+���G@����>)aL/|yK��$��P�v���j��i-��	Ӹ��G�\��u�FAC�d�\�N ���=e�r�=�P�hP�~ �Ù>��BL��^d� �	�w�S�h�g���V�gue�g���%�(�$h<L�g��pjo�u��|�O�N|�������E�Ħ�����Q���Vm�U�5S(��]��h�v�Q� 	�V�v �o�N��Dv�h7o`|�)��S���ڹ%�G�[u�mi�C�H�H�p���f;׆����:q���r���{>�����s��
��6>�OsQ{تB֗�m��3?sm9�ڷ���s�� ��1�Ⱥ�u���7����L;]�q��z���o��Z�M펃���x�ykf����k��#���M�g\j�$UZ(�i�3�⪫K��[@S-�I<�Lho��J}���HF�B\�(�J:	Kș�nc�D�ɞ�4|n�(�x�lM˙�o�	�Y�-w���+���� ���.T�0`-sƫ��9���Zw��Y��O�a���(�Q��s[s���
�z��~����c�@oȹ�pp"���Wĥ��>!�u���z=���0}Rr�.k��g�(�,<�@j�:��>���Y5jǐfv�����_p�+�Q�8n��B��y�cW�%:�t��0��#Gr���<Pi}A=՝��Vq�Ќa�yI��T!���g	�\"�pxV�A��Se+7 ��@a��Rh��߾�1�h��q%~"�h����ֹ����)�j2�P��Ҡ ���v�o�k������j�!cY�����3Yа�ۚ �nĳsab6��
hT9����\�ԫK=m�9K>��c����b([s�,���K�,���Ha������
�$�E�v��2��4�8B�DV���Y�����dҮe*�5`�ښ�������y`��p>��>�}f���d�$�%8��A)˹>Sow�]���'�<�P����/?4k�b�`�;2h��*�-~�u��*�6��-��f�˴��f��"w��y�\��V��)�����acݰ{;D��˃`~���Eg���`�T�k>#�Hw�������f�rH������/���}y���:�����V�~y-�k�"�H%�i�2}1Z�!�Z�Wsj�����O!�f"�	W�g��ZxĲX4#������H�8��L�*��XvD����EB�O'F+��e*�������X�.���]�t�G��f����mBFw���,c��%��!��0���Bw��s�<f�P��2Du�q����?J�FG99z9���-3}�K�V.�gd�T��
Mo�bȁ�{;٠5�s�^��I��>S3��,yk�@���$w�6=x��n�k�Q�.I�?���qT��1/�4z)�����ߧBQS���)�2c��r^v:��v��=tJ��� �n h�ryJ��6]"]�?~V6XEL����gA	��K�&_w�Ep��Gyy,�B�Cu~xV0������p�赫Blm�:bv���b-0�v���&�����L�D����d�-|5m�����?����H����5O0L���&�Z����n|�3�YTXoY�5}d�-}�@�%S]R�7"9r��� 4œ=nQ'�ي���cwU�^���Sg�v�+te~)A-��$�O�j�C��b��9dM/�®��`�9��vN>��R�5(RޫL��ʍ�ݼ����C$�ם��=	֠`����CiTQJx��y[��qNg@�A��`7l���L@��A*uO�l7��h�Ԅ�3��g��'�ޅ���� @��=�\b�*��z_g|Լ�M��A��i�#�ҋ��@���HxkT�6u�߅�f�W��X2�<�s��8�O��G��3�K��M�Ibk'��yX���݁�HK�Wf:6�nqx�Li�8��0�AaMt�4�C^�-�3K�0�vH,A��>�t���~�Ĭ��Fp�T���8�:��A&���W�~	�G&����ǘ���4y����9��.Q�{ϛ/��o����A�mM{:7g��xn;�e�䅬�4
���K�	|R(0��]
O}��*
PV.�7�d�Uv£\#DͮK�\.i���0�{�ߢB�ϜCkD�w�ǐM����0�Q�d����"	@�2�����3���p�B`�#״g�L�L'pza�#���-�f.&u������rN�I%��\��K��$ "�6��W) 2��E����� 7�t�xC���:Ї��N ��(茵H����0$x�*�c��]o%�:d�F�2e�_�S��$�_���w������q���:pR��A�"i���{�7��g���G�ĸ��`�Ul��?�Y����B$���,�ߺn�6���BQ�)�� HQ���#OeW�Jz��&�nl�W�1Ᾱ��	qm:Pi�$��vl���}@�W��h�� ~��=:�4&��{^̘;ld#�Įi�_�/�xp)�_����\��ź�_*�V����KΝp��h�+W�`hciu/�^6`��7�����K�C�D�A���T��Ts%P)z���79+?b��J	o��1�c{k7c��+58C���c\�w�<	�������=��ʘ8�q6�����F�<0� �姛�"�"h���v3�j��&���*�.��]EXڹ����Oh�L�����q��1r=���D���Ly�ɯT�n�b�"���Jy����
�h���f75�����\"7�g4Lߠ�]�"�7�N���x���<����H�(��H�$p.?�4���9�leRTd���PB=(m�$F��	�%L�,N|L�����K���]�	�)$rбb��?m���I�E�^�aZ/'�nC]���E���z���	����{v�>�}��}��zV�5o#���NQ(���~�*��Jh[@U��F3d]�:D�B�в��f�ql�^�������;!�<#���d������>�M��6I�H5�3��m"�ݼp�N����Jo���#R�e�)w�DJ{~r�G���FV[���H�\�'��M��*��+�@�^@;�U�ZUr�G-U.W\����葑e��u�M�AmmN���&Z���T.��j��������g�ɆEn�{��Z�R6nt-�ّ�.�x�'D"t�,�����6��6`_Ǣ�}�}\�S���,�8�}���T��w� }�:�)W7R�� �\T�8\X�f���\k�Fi,�2	a���b�G�Y�KZ��AD��U�;j 5l:L�~7��ν8�����j��$~�Ad�v^^�L=��m����ƍ����K.&V�����z�:D=��|x<��n�������i�q�!s�I �J	ې�ґ�p����;��59�G�|Q6�ݾ-�q��|���:��nT�\�[`FrތVP{���5�X=�C� *~T�$�U9A�wH�dt4�\����ܮ}��3ri�������M����]��]I��&�����M�aж(c=.<N�@�!Z�Q�X��O���_����L)�_�H�q���.�3�i��ބ4�!�n*{M�tߓnC��U'���x
�F/Q���"zj�b��.� �������p�!.�:���?�N7�,S�<#��|�U<B9�J��O���Ձx�*!�ąH�qٖ��	�F7���U��F��ؕ��6�өI� 9ILۙt)0�@ ��Bۗ;kj�x�%����=M�i�m�,�ӞԊRf8�9J �
2���Zչ����p���Q��}o^����P�R�5	x���<���r�׊�� �O8ɂ>��?e^z�֕L%A��;�cN�#S:5-�l����؝��ɡ�u���K]��:�:TDm�oT���1�՛"�hT��tV����y���>n��'S��rGO��YSv��W!;ܛm_�~o��N�r�8�IUܜօD��W� �
�=�`�+�*1�mމG��
n�#_��|FAS{$��WB��d��0��FP%M̿^�O�Ja�~���P"�����U���sc���Ԭzm�[�v�e���gh���ɩ�+�_�*ٝ�
Yc�aW���*�C��aC��Z�RhDb �pȂyP ��T�͹�l�T2u����h2������ޔ<�)$[6X�!�O��Q�'J�J�#�.��A��9	^x�s��>.�h��avl�k�	��w;��ꤐȱ���d\3�201��UzF�:Xʟ�g���vV�fo�xg='HV�� �N�[�C/grH�����x��)��/%e����C,g�����ܸW�,\9��]�*�J�դh��Մ�>�HJ��+�fcu�ЁZ@i��!=�^�gP��/�q,�1���j�D�S��mǻ�����\��K6�l)�K3B3)��<W5� H��Tۚ����&ĚY�Sn���G�-23���O�'g�qӮ�}�#P�0����݇L�7�hR�=وX��ͫ��nl3�w�T�B��}�<8L�q�,TO�E�Mկ*Ȍ�xj�k��|�� ����9�Z�b��-�����i&+�2�!���$��0g�O�C�߸��k�_��nf;O�����;��W�4r���,�E�y0'���]ZL��s�[���]�1��9 ��~V12���аAEV	���/mK�%��jQڥk�z���UK��������ɝ�D:�G5�_������yM2�Oj�sGA�kV��%�P3R��׮L`}_g7v���M�H4�7Ƃ+�Mp�6qw�]WG~*`K!������1&�ɭuz]ж�/�߽��Ⱦ�JK�A��Q0^�l�� %�SѤ&bg�ń��8���C����t����.Eh�9sa�?�� e��>j~�ɗ;h\���h��2Ba�4�"j�w@)�|Z1wTU�֎OA���l�޿``�gh�#�����=uؘ�U
F/S��?<~�j��N��j.¦1�	�_�	�@ X0�������Aq�}�N9��S���W�h<�t�������z ��#��=�t�
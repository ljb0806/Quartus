-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UDapoWBq6HZtVZoiNEpOMArzUG7HE9FNdeSvYX1zJ6ohTTSDxi66hFMBhisOp83d1/JQQUxEoGgk
CcWp53/+pjjzQbqTcvYf7ntmut/tGP9JEEaORPhGle2yEc+GmGchCTCBzXqNAeamWcxj4/SuSzvj
wgEg55l9PxbfrnD4i24eBvwet2y8N04nDjy0ybC3VXnceMrgIbLGA+psr/Mv1OooWXQ9hd8o2XNh
0+CBaXGwYQl1QU0EZWqSo+1KIjq7aBnxp74mX+ptgkH3Ho4Bg6mwzrXp1iNbzxjFRjIcYJQJhLIK
Xz4QI2gHbv7H37QGxK0YbWdJ3SBRw1PZDb/GKg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
6qNM2mYmpOp/KPLHnFEfvhKVrh5R3IrFGRHtl27jGrIB9wx+Go2JEJ/3R4a7XsLkSsyWQGcenop/
Ps90vX/pSmb8bqEaKuINoWWbHIa2emfUgYU6oEGgGLHS6IyHatwsXSc40M2fhc6Ufsf6REMtl84l
akwgRa2YWILSnLSaYSCIIi3g1aqxSxBwFcLRiuQj+dAcOpZ0i0HqvdirHlPurE0bjs4XHQlAy2cw
MqI6bjxw5OrvWn11pUsIlbHqRHlWabh/N+iSvt61J796v9dUJcm5irKpd7U1Gh1vW/Jyc4Zp4grv
tsG48K/3Bh9HPT72XUydw7jIfNVwdVrxMiOq2Y9aEJGWqcwXQb+D+CcmSCPS62DUuko4MBi1xUXN
kiZReBPQJTkCmQH7yT04AoyeGIIF1HZpS54NItQG1q6Kq9h/Ybf2udqr8nxBOJBmfpoNISI6OHwm
WjqoAxOvrNBaVQ4NNu4Oy4pzQV2/r6Sw/VmW+NhHrkC9VmcSUcS0oRJBtUYZCXyDVy9CKl9AsDo6
gzcdovzlkm2iuuZy4V4PeF3gx/kz0qU8WZVlstH2A8tioWLtGyOqzVnr8U25wBfJugEilIwAsnJc
IOAqLhTAP8RkQMQlT+qm0Dfd9xc7sO+Nq+NkXtE7dsFuBbFqi187YQ+nzM/XSSPiQRcyc1W8aEta
oODi83V3wNkGVZeIcYsStpP9hhtU0E9pFKdTKDsk5sTz2h+pJNksF3bYKDbFUV8exbuqUeTRsUci
4yqwGIDGc2FgwnQGpyvbu7QsCnABMted7fgQ1UHRt6U169nF0mELLDWleXHsR5QoQ2UAf1foQn4L
WOnKMYUGxM7DRbvG6APsyj+HrGbg/2fghyTzLEQsMS0OctiCwGxLjTgA87jQ50VYCxQw+B/NbT64
D/fKQahSe314vJB5cCeQUYGy0niJuXaXoVaqLDMliZQ1kJ604wtYPFDQCt1LOxCs0NssrhHk+dOV
eokhEppLMEY0sytRTOAY6kD7qAU7QW//css/Od6B2F9Q7oeFjKsigsH3G6RbKzRLD2viDpKv0c0I
dKHPqjQTEisx4nhufbABurey6m7S+LAGfNKbqR0/yn4EEaFU5mwhbQGU+eF8srv6U2igYB/bTNRC
2x+09361lDY5Beeea/kkJqQ5LH0KdfYcI8MK/6e923VRsAPfM0c+DAIGdOJx3OVe3wEfDtCHkdLc
mkqVCmJ0mPoSHRt7ITNuI2BNczDr0zTADH4zn2Ot5GSBfWyC6z43n3bgCU2a/FY4jNgVyVwZY+17
/16ZrRAt+xrzBcPUo+WdBegRRYIT8USRlQ42falSjpDn9JZgUcUwYGX6kHhyLuply2ZqQWFZxT9T
cE70abuXwCNPmgtOtuHlVsKPNdOg3b/AB1qX+s6tH5asgECGlL8NpEhBkzD4Ce2TwA55P4alDoGR
WXVtKYpgSIrz7vjKeK5jpBgASXLZWseB7OGIri3O24oSoIHGVkL85sK6kPmstmWKutqIBDFOhqW6
NNWWl4GEIVMsneEC5zeuKceiN2eKk6PjnjQ6oB/xTz/SP20A3kcBOeEYMrDYLDr8fZG9xitNZ91A
1iwY9EhQRSRIk5gTRfyGZ+ZpMOy09olDyrifgW0wEHmArH1UIP8Qp4Me4wDyX67Ne/+6+K+SoE8N
UimoyLy5+dJKeJY77Jl774csnXgAyjk7JRlh9zyge0pB+RjmKJn2qfSzdC68bQbUnSSSf69aUq/6
U1++OjZM7rV08sXufMFFfGFbHWkdkwDzgr7eK1IwgRjucPJpErrnLtuel4y3NAt9IXBDELffb5dN
712PbZrjl09a/hWHLPA0ImJdlCDvwTv+ORfX1HSMtb1t4RNr/4sJVnFhmB94GZReHpc+kxZWw+9y
meOcjPr9HC9TiRZy3nNhA+5gtb63mofV5/qfrTmo+72LU74unYR+/+yaBWAfBDzbh3curx43+6tY
kYvVfLLkQ3bjPb6msylNr1SoKm+dBWPp6r5oR+HJThiCsR9DCuEJdFTw+HA+ufh8/4tiRPiY5Z7z
HWgMn+XVX4acUwTeRMmJoqwdKXXyi5K4fMl99vpTrWtqaqyPZ1sm1BhGmAniEjVs1sIwrw2VRVCm
tY9iTZKwXw5nlySIOqggufQiCEMTMT8obE3GW8GWtjaMawUSqx+aXrFqqlod3j7TEGjCaO3dQl+j
sELt3d5H31H8aPxMSx2Kr/0uvn70PFlCh/bTgKAvOIjmJpWNNBphGlyuJK9VBbVLZVQJ5giub6Ie
pifk95GKNG2b6Wzc14k6PIMb0VWw3TXFdY6VfcOuTPLhOqad+C2oWTYZVP4P8llTcZBy9CAuV1BA
LlsZ73iPLPeueBpBt+pd9CvII2DDWi5UpiaL/B/MH1Soak8G48Nty/3ihrj8ff6M+j+OCLLjpIyq
hffyTZkmN58NIKU08jOCoMMj+TR6eunVNnWnneDz0tn8tm96BBbO5wqoP/wNGVaqGAOXhJ+1apAK
Iq/2hGU2AwQcS3cvObzXWtKeJBQ6vSNCZyIL4dHektKV9/Y0rb6h9iTxZI1fp1Uc8g6ESsojg8jD
j45zXrL7GpAyHZ7Z9gj+tVB3W0PrMyrWpIAGvOyKP0Yal7UOk/id6UUXIZrSKqProa21lqCALj2C
Z7yT36JjZyZWPqGcmuMZASPxqX/huEKvdd/Oa5tUR3zPePdQx2eNRFiYWBg6XyDSdOCFC6Pc8Frv
porV72C7hl4zCuYmYfAj1dsxUzqLEB8i0SfiafDY2FxhLCwIzKquTDYyMw3lHX7YlQiBtfI9G5fg
/7gO67cJVvc7ojuY3gz8NOJpZ/luEY5D5qQ3c7t2Ma6pDk7Xee34CTIBSzkFIm6rERqWg03VosNF
1jsf9DKh//z54QLlbNfjo78ttr8niTyec6v5r2OqeW0Z2lPV8IYvgF34DmC7ujl7CTmcAiBeYsoi
BLnFTOvm0xr85zGcNWEVj04ljN7Om3tkytATZABcQONuLul7x7pSX/98Uu0KsZNoEjGVroA0c7vJ
eP+pBeyhcG7vuzREGabrycmADLBeXRobtgeh8FOheqpaB92zHQAFMGS0IhOgEGhtq2tiPtam8RTt
ZzP/oj0qZC5WBKF1y+MVq5f4c31+9bXw3YuGdHAjHF/fUYv3EqE7IikB0yYPXimcMC6+8IMjPBXK
/vKq52ywTKY/SSoqAbeB6iIGx5p8lVNMKAvD/GNFd0kPlU76PAymKWCSIXMekSBqiXk2DdQXfJT3
ruqdd9ZyHp4ajbPAuidZlCLFr+vFpVmNI03ZImtjEeJyYZSPeosNVes8IA1bXqFUUBZPsm14xrZT
hm9Bus7M+Nf4lPMqpk1LNDu3djFEyhoyb/AxPYjLjG5AaUcmawEplKpMTy6pwn8S0mk9YpPq6SYb
pZNwVcEgCldW54j1hN84T9/WwFZmA+/xmZF3Pqm5Sb3EcV4QFy0U/n0ga0q1GL1WDZ0RywEtBb23
rWsdSCX9SXmN7iDBvsx71ve9gsx5axWs0HvaCWfLMcXJIEieVIuTYSM+G/peUX1/gn90KnnSjLWz
DyvGsYc5VykP2iUImNapvy/M883mwnaeGuZrsvgEmAvV2AVPj9z85poLjg/hBEqvdQuZ7nrn87aq
ez/rfj9/GALCnplnS4i+fpQ6kNNbRZJn6ApFup+yTMsv6YtFLEnzAiz8sgED/9V0Lz7AMrnRLUBb
SmgkzYHn3bT44r9nCsWbkg8zkxsXfFt+SkLWqjUVR3N/1Zgnc/QSyQ0vpTFswKGZ97iiqoARjhv+
uqznYJ6c4Oe1xyPkC8aRCCrqcMLA98fMhbz8F9KhAu0o1cBS1KXq3lbmqgoncNWwxeJlD4JBtvId
8G+GnM4c5mzqFxPFzGCbuhELLlLtGUi62IzULfDagP+HQRjoHX9JzkF7NbS+DDwyFJTev9kwbn8I
Rzc5GLrlherfZ0lfj7DgxWiwCEyo9Ft4F1L7+k/Pzzg7ndAj+YZBj+MQ36kq2bDhHcG7RyGPBtT3
3Wn3Lp4fUNmE56RhPqLFrsu9ofCb3iH+7jadP1vPBfIPz++/P0Hy67dljfZKnqtpGG6WNo8IvxPV
/+Vas8n8bXIlpSm0HQKx+wOJEDx9kPNxECtOq67+gheeFgvZ5nUe/9tZFgRrDWKWMQmBmRUa7SGP
q1waR4f6CzQ9UlzX4der+zOW46wbUeMTBMpCyZslguUNP6ishTjHxFw0xDyztDZYm6bHNR9Vc3Ku
wj7+lDKZxlK0Xq7TMqmv1ZlmZUMKg4T9DIHYdNnkVaSNNoj1eW6jei2jug4FQzUdB6n0dDJe2WYc
PjAEMLtDuvUue4HWLzBQbidWjRQiygHGt2IcGsOC11IjkSNBqxnB1qz5uPX9PlCCMJvZuLkQLcGs
YxVVxHts4hdzRx0LbF1eJszhWKsevN73g4tV6smCjOWqiwb32e6l0tafZZSIThG7lbVhFdyMJLTh
1jow0GipYoPMp++cTy9xJr0Rnqa+I96l0LlhNkm7RqfTKpeZ5f3jRqZA+QprTXX5kttD1E+FhId/
vTEM260VHzMs90gpBwR4lyTW+U2DFp7DIGgK7DalJPxQ8knIrLwuFzCexUTl81yeedcw6oSeHr9L
+LTRBrocKw7sy1n2UAN8v9F1FrhcXXqFluNswtteEp5nQL1RplDIl9WQaTWPPhMrA5CQwYn3SH+V
/4soJ3zQ6H+bphK+ZDmV7Ct1fbWuV67BTG5uMWrjjml7+wVKx95neWnI4T4f3fzMM+aQO2G79RjN
L1PA8aGLXZFPGYNd6gOzBs6VaSCuUANXo574JXbowS629MmsiIROElD0q63ozAJaioT7o7H+eQZu
62kYcQBnvhpt0uutitIIFqKdb6lmspzctg6rLe3GHzvmPIqHwJEyALgTSQY9fNI9c0v31Sxk+eY8
SrAvyFq/aiWjLaV3ASaRbzmCjAECoBTNmN65KfDIaIn+YImcc2+A/Oc7T8e8GUotCBziTDAQQOro
x2x/mGWBclG05AQs7Jj9s4QHAveC6lY4lpN1DcAH2djgQ059aSJHQcdvTkwCOuHZ/kVPxb7SBrD8
c3Bvh1bnWac0z4gxoS3VP953kfuhSShQjGizlvJf2Z7lG/NzsC0vAVznD4bfr4wm69SekYAeUxMr
ELpTqczX+iTpbSgk7Er9MJEvC5S9tnnLheipgRvsKQIG0WDnxM3o+maswy8n0JvFPEn997nzcNvM
mgoAkv60xzWsX88VBhJTgRncrUjjI6pprdWkZMcq1/G/O/i35HjxdOZvU1gPTgrbiM/M7T3jcyon
crCIRw+Glx7J4SOCyOG73zclb2sCzSfEeqdx+z/1QUhcjdiiC0WyTbDMTN3mK4p9rZbY/yGo4uyq
n0wwumZIKoJgDQmrCumOABqA0Bw6BvqzJw3iD9fg2wovYJyuYHXdVPGd6fXEhvFZ/eZABnkhQrvv
US3VJE0M7/UQ36Cx0+1wTm8rjrx+Uek1gxpVfIIy9Zz7nNEUaB0lz9DdT8uOobO70qVLiFnbSVWY
+mjAqbUIQSKa41eXyIkkWRveQ+T8Yk9QNFWaoyysIslYg7nKKvif+MFDOt9P6jOOCxGriAi/Zv4h
KUawdS/Zrn0D+ubepWq0Y/5yWQ5ugRWXRN6TsRXgXDRKBP7K3zD83xN2t6+wX4U0PJi2b46+cqpb
ngmVx8lFrN4ggkpNnPYlqXorelfFTw4yi1dc7N8iwYqkcXwunl7oitpdatByIsiZKtgwLNKn5+7G
jR80rkzgAmxg0jKpXXEdd+EL13aKVAf5jEqu+0oUL+VwceMMO0umf9GglRQfWWsyyAqmhe4UEnw+
Mjruu5Z2rC2WH/n5oLskmA140KeAJ6BgzvF9OhA+Swil4jKuC2TrhQXLzfNmf71OfFGrcLoKGxhU
gdE2zaVSMhcOnNAIYASDWVDbpruKhAt4/TXvXf2EoypYLF5/NM4vjkIM4fDY/z2lCAyoobf5KyGX
Y567LrxDNDlu+ZdirqUvGC9Z3ph5beIQjGzbH1pf0Rc4hE4abgR9TO+yjNY/88sL8oZs68WdKkQV
KKv8JGgN2ZrsVi8+9TuwsyMG8tTwyGoN5FJ2jSyY1BJxDMnfLsDr16rwVkyqwUPk0EJLm2iRX2EA
70+34mSY6ihinT1NI4olBBWwwL5SQIYbgfsRgcNDs21isZis9AbVYvLCTByaJZz5xavCvwL5fBkh
8655sDfH84LnUeeiPClLFIUvgoM+Yq8DWN3uEUb1V5qWe777VYqsJ3QHPlADcgAtrxX2CDnGxbKX
oqjGYRJg+XlI/yHvA8WxS/Sno4Hw31xFhjqW+psKZjAjze16CrdJvMY7KNEI/AaAeOF4ZRMY0P/V
xSq1Gs1xhBz1uBoF0HXpRUsjatvzLElrMfAZ9FEvD3VJ03hff516pP/D+IbOa/RsuxqmmjbCx1B6
409x2TzAeyvSVvMyOyiTnce5ZVgMapZrQ8wgW/Yl1fc09aJUg4OEwWOfInrTyfyBJgMPk6f1OWR/
ArKW3w04RqdJFI7q14T3IP3qnJq7nZVM9G/j3QxesXq+rXP4nMdX46gj7Ls6Ys4DahzsPZcMt9fc
6GIjbuLadDGozhdKNlbocI+s1rZUE8nfWWBWqkQ+OD6K/F3Di1LAO/Ewn83oMfa2rbMa5/vx+GHB
rhNZVhB+lKfm/MqK73vHUlPOHHZwEBeIlAhZoue0PdiTg5+ot9eDr7w+V2NKZ89dI4ESHcyy69T8
9GEEMo4Xlhsq+fA3pz0sOkyWrG+x5lnr25kaBVVAx4qQ4t9Np0LMNJlUCpjlZpgA4mezX7uZIlpy
UBghIJiG6jDqzuXUG1GM/r3+yMioLS7oDFxuKbh6cxpXgmrvioxOCBGgi1pt4b4W9LciFLiM8sbB
MOoVmHGg/ZKGwFtfe/g9JSOai8CsehPDHxULx23AQKppJYf3mnpKOFSuMMSF7fvMqsEILWPplQw8
DHpqcGJ1oOt5wNG3qqZuR5O9Xpe/DGfbilOuNaiEJ2/9ZgAAFiXJY9rvSoDZVehwctwvth7OcPBG
ZqX1AeEE1XNxiKGF2WwAsLfB098dmvrfzfYbQOaY1PnZiDJ+OXnJHos0S7DpMwEcb4wi1ResqdYR
8+8pjOB8XIGbWilUC+JMZH3x3Fa0UafW4T1uSxEISjLt7EYeHFst2xeRNdWvflzUl6R2tPooQwSF
mlZwife7JSg2KLFTNDUR7uqSNVf7kikzPGu8z6pbWZqlyUcgkUY1zMxwnHqxENz6XixbqDzD368C
AkJi7/NVg8Iy4VzXVIgqWjjHgd8CfflJK41hECcHzDDn75HkOIJ0TEt5MMV+0ZVRvkWe1Q4eehRy
ugBuYDtvzOPb45KBlqrW9UyKsJimTfawJTb2/PMaOOi+WWC2DOVGkis5tVLXZX0+MvzYl2QhO+R5
MYjDt9edMINyPnmOQq+xGgv0JduC8IgorNF65CjMXGz0iINwT3lr6G5L7xMtXobxJWgaSYJGBt0K
EiSDbt9sNjbwP8KTMsZoTQIbtMctoUDBoOsT2rU0MhlT7v5i8CrmMOGFux1A87O8wg748TK55QWR
/qcmjR4JBq0eJfCtkH/WQq2mcxDFhnaRsVZ2IYepat9GqrscR/JcHC14KAFUxWIWxMwyEVxiPakx
NH2wRC8aPwmLp3ZzG+FXJeYBqa3FOVHe9U3ISypWvOFIFykA/hdfdJTWFz1iGArB0CgihGFqnaBa
ZXVIZ2fKDYar/Uvv4uE4IpJ/lsCBNmq3D6m/pmPYnIWO/8ufO+e9/oqPUoUE1kZStRFOaOMan0Kk
5SdIKUrEvtBvdDz1mAyM1+Hy0Qkx8FNQY63n9xp9CvWFyqZCANMgYL+4LFO2zQUz0KzhhC6XCOKv
GnzAWY+51iqszciAppL4aiCffqlz0n32lpSGFEljmQUXYurnbkeLfVCznrq2ghLTQPx0mIdK17AX
hOA+nfVqO0pGUbshJXEwNVazhFDPl8cgiPJaY0aE9Yh6vvD74dknJvPDGEUEs3v0DvCEa1gom9Vx
9k62Dsn/B/OlPJ7c+7AHXcToXrsiEnGgdp78tb6MkUKenPrpc/WXEcDmA/Yln9gAtH1N6Rjh5D4m
B7fvpi8dFDioqNzzPej+dszzVrzYmks+/3KfZKHj+orM01Opf4Wlc+lvi85jIkM3lFv4OuwJxXcU
cdvxqR8Wfdnhu40oJWwQZGvdTMIK65zBY0ANwB1U2nSPwLxs4SdFRBz5Cwn6QyujJj2cyIJKbj/C
PbONxhrx7SZZhlu+CcT4lfQ93O1v8LWKDd7E2wq9XtUQmtDXgzk3QwjYceyMr/zLIkg7RwAe/Njw
ffvdismJwhcVPWqgY9hEic7N8QoWsgoqor26kfW6vnD3m/vux7VcniFyJ2NhJZUYFNojgKh9VnWB
um8mTI+jxynahDwOt5gXygFWaJijLIM2LVjEGTWZ8Sm5lalf2rlv+a1n5ru2nTvkNLxGslUFCuRG
dKTzQPJpiOLI1UtsJwBi27zt//KYNDTcP4rBO+7Q6HwFljgsg0jxhBd+aE5Iwd+InmFC09PsisjW
BByEbVIjaOE2vfAmNlX1c4T2QQbZqTWJjrQDpdziYGxJ7PpvMde9xGeRuidNaW4yRvnMvnEE3gbg
rXNycQ9U/6bCkUMFzBag4hBjUHZnd8azG0HI73VDn8YWztpUitilYazmwHFQi5T/fiFiuXU63V79
YYlK0FIURI7W57N/BUB0POBFkzvwJNzn8Ck8jGsuNR/d2WMpc5D98wEwWceUDzsr2VmW7NkmNDbe
hY8vICaI+94qa9yU0+gXzGGKBwQBDZ+LyTeeaturE9PuAKAzp6ImbqJ8thpBGSZS28H7NRQwvnoE
1349Q+L+W0Suka8eczUUs8BO5Wc6AZ2kI3LOC6G3xiMhJ6oRuKoUxyQmTm0Bq6mtYqfqOgNmvgoo
LOU0KNlkqXai18NjPkf8a7nPERE1+2AgIk8KwRpDo5d43E0Ynqu/3K7quvJKbs14tWUqG3JW+9KG
CEaMGPNOs/QvJf+yjEMlJzsb6XpZ9s7Ib7A6h/4HF9Fzv948Ssozg8jVr2uDxr7cdOmehBNC3Rqk
pFJMaJSKw6U4LjLpdPEcOJ0UnjDQcbbfo6Ye56Nd4fHjeKW7kN2U6rh5YpN7f/7aaZg2eFnjI047
R7D6mXbkmlEdrv+k+deHzPpTd6CgYfiP7RV0NRNBUrbocpYJITtg76owZzbNpSqerSa1GpoZw0+T
CFqsgitHQFb5Atl6cHLZiTS7of0wGQuXOvbSfdQ6zShnt6DhlNZhbaFJmBAVrv/kF2YHanBCmPeG
NWU7dHkOEinLIiyZhMdrmgr3PD7o1M8d6K4bFg60dVjWURAJLQTXBrOKBck9W+KnK6vvVxGy3bpb
Lrn4sibg7J2jp+xt0SM/7DmIO9/v50ZsCj6+2TWYQv4Uko3cibA4UnkPszTJyeEqrhoQ54UvAlw8
j0807tNiepApffdiavfaTeL7mBRA8PSU4i8mmArgE9G+FVFvRlmoUQezSlgnx97kVbsfyUYuMe++
UMZuzPZoOJ361HBNL5KfmFbkJ/e854S0WsoU/Vod6V1IhQxTDogOfUSYdKCJbaNMWOZqx5sJRNtW
jzOsDN379CyyfvOtGta5pjP27HVvuGbbDVRTgP/kukDtQPlvCUZrQZjnzyt9e8HdiKbWkMVm1jmY
/O3OT3ix2H3L4apkxqCqozqW8YN3JzJHBQ2/jlukZj8SlmDbsRJ8QYOHuwY62m/YmUfhxds1nhY/
xBqPTJswU0r4+x9Js5dbfR98BUv4M5+otAlyZrRagHYMgXVbm9P4XW/21kE+8ADWKP9fxrbansYZ
BaEpIAySZIqI+k2emfAtvzR902MBmTATtesFbdJzBmwQjkn8drB6gfgbhrq+usbWiNgLNiteyn+n
9gLdt148Oeby4mf6P1OyLqPGE93Pcjz7nyEWHV57DMk0bNGWu3V0la9kEAOQZCsBWFjZluHCH8oz
MJLyoG0G2JZUODxKkqp/qZUmKDn4/6uZarxszzZd5p6eS9vju55IYVrJVb3z1L7ZuSUEEzFYpn+1
N23qE6DuPODC0topMED79VukcWXOFJ7wmsXbpi+iEGf5oLOkiFWLqrwyathwqFhWvuz9oyaJPOZY
NrdQNjdW/fBl0FQaphsrYwqxgh56FnJDoUNhC1hksqVjFoBS+7u+SGAFBmwH5KoG0erYKVH4L3qz
wwW2K+JJcO5Uhv5yVFSqm4H6w1754FZjTfFSXlULQP8XPx3HavFR2nvtlTNkiAiaYbmWAFZJ/HNc
ZdWiKiRHRsc167Q9X+lklDMtB5z9QayNMXhgLJGoys5MHNG0bdVFP5/RBP4JocDVe3FtBqWB+FVB
fKymbcmnaZrAlEc63+xHdIceCv7QByJDPxlp75E2HGUXwGm5ZpffRtyteDacYdZtbwJOOxhcN6uG
VwvJoWJ2h5P5kyR9iLDDk//SEBW8GZocrHMS+OXsMEFgjwwdfuidzsssJUGMtOrfDZPG6ryMtQSO
jEOVaVeWNPqtGmkp0C5kgtyxiyu5/PzcjUWfzcYzG6sYZGilDqGVi2JQfRc12kYVw2q29BWAGGmT
jtFGaQTETn/xykDIARp8O1K/e0goAjNGt32uzVuzf0DTjzsV/BghTVvke8pGQKwAJzgSzeQBLBtx
1LcLvWGA2b6p40iRNh4gIFZRS13g9QoEioMwq9m6hUX+Tro38eXXOWDjCLTpUaW5VcOu4MhuKW7r
n5NsWjBDf8VmqAHblVqxGRJ/Q5GnmaQL2CB5ZoWlJlYOJJrKUSXCxd+27nM7w3j39yi9XLUdNwHQ
q4USTXM7jWCvFb6mFs5ScSjpmpbbqZXeU7f13CtVkahmT0/rrzJkfQONL20v1Ifj9Ffsb796nnZq
rHxyd6rQi2TNMYG00qFroBHLQcT5Gwbr/q3BhleMrLPcEazP7ZwiunvJBw0UlarhyfQBb2wE0jpM
Bb06zAzNzLBzVd20xHOpFD4LdrgzTphFs44alyVFSKeNry+SepJ1QeBDTE4rX1OTA4Do4OLF21Wa
Jf+0apXc39bVok932vNb/piKkSpAuDX4iwl2B16i3OKf3B7sK00OKP5jh4hXrICZXnDIHqgwoMMU
mdJNNXiFaa+nTZZP+oeyNdFqNrjl/McYCvTvv+vZhKmz/ZiLzf7kkwNIcA15G8yHXIqtuylq+gPt
EAwvKjTeZgws5Buc3RmAA6UvtOS9R3Ym+Z4tzYA1WuKwd8TFqQwy24gpiwisyiN560gM9efIMCWd
I3OA2Lt+EZRN+pei+xnTzrs7Svb0ROQ3C0hhTvAI+kCgBSJa8TOJSSfdmRQJ7O0LTnmggvLa10GG
AZ0GGejzvOjINYYrmrwprZFgyfK9T1fPK3xlzaSBTBsM06j20qV1Gu/mwlkeKHXsaWmlfc9U+67q
D6lGMa2+O2ACNq6Hg79NZeDoKbRuAlhXk+ViGOFBxW3WxiFZVAH8kAluihbDNeinTUSGp9ee7s+Y
Fw+GWuPsvG7yFwWDAbXTXogt0Ei1zB6cLWCrkqQg76IzC7Cp3c1qwX/ntGPkQXwDjk4JGQ5JfMER
nBVfP5Lx1HwkWRPibhi+jqm3jerJThpYo1pBQ+R5GUbgDE0Rn4ERSqsfw2yhsimLi9squQ6CCHSQ
b8WfSa9Swr9u9tQK1kxWjKWcaHDSz/tF0ggZpiXwSH+5PEeP16jeu6Zc4oWfIkwaqb7JgLkBnr4h
K1BLpOCHQka/T5W+/BjLvgKfk0CXUHCfMnY/sbbvsY453dc+Bbd9BoVLHiFwPdcFi27zpuw8d8kd
qsEZ0MaUwMm6YfLq+Tr/Od0KNREi8BdhsL/FAAhqj8zc0vxUZk/e5BZDFlGBfu3dV2aW7NLjAAmE
Ot0LoTOlVUx/cMjFj9NWxJqdQMiLNSGJc/23k+kcYxYWPxNgyzXnxMGqQ/CoVIDzih8FfMfkeZ7C
ToJ7wBDItfW26nD0RbD29cJ6RdMbj0sLqt89vOV/bkGqfp6Xvyf0I5Paw2LHn0/AEjAvTjpISHS5
0E0KsYQ9KNerPK+9RiyCo/k0oR7yZAt8TiGx/5/gSOqB7BBA2b8Kx4Sd4sV6YJGkQZTdATenymuv
op/sUFJQS8DjsHaltp8/av0uBWNwlMWfTPM9Tza/iFUbZOnCiLOac4JEDyEhQU3csaqTmAOME8Oi
bhhkbmqQ1+X+cqNxt+VgrK6qDpeqVgNhaSoavcb7esvA3Eg95Fln+MUpYw+EP+34u1MY0geyoKE3
iXZtjYjjVIqHnEypy/c/QqExUGQ2gYq7/Hsg+KYSTIf0CGRazgqShK0dJ02KtYChRGoNX7nntnX9
YO7aT6PyUZY8fLQrVBHx09IujCzbcq0oKYpjUKPGk6ZTXswgjTEJDhtyZFw3rCoS7LB3gSKRVM+9
+PmOgkIrJNdFjqeOxZt3RFTWQoz35RICFEcKDT27Tk8VQN0RaPKXS0i1k214aZn0R71sSmC7W6GU
jAK0HeST7JzoXuWCgAi9N+eromL8qRQcjAX1pOXaN5j0pREYJTgWX98ORE775QCLw8cWX1KCEtpI
1QvT1dc3jCHKw45MpW81LmG9RRxtVQznf0bKeV5oTV4T8Dkeoy/eO6RwdFMQmuGVC8fmUVpmsFlT
QehCE7KqN/DjhexNhzoQSYJZiYFeqvNu82clVKa5w7Wz1MVM+ktJaPYel7sWL8dC9ntAcev7TfYh
QAYB1IhHzue0FxTVN+r9WffL/FFwy2J8tex3htq04w5kyyp8U4oTNs58J6cHbt7yQgbaYEUSd+pp
i8CXM+GXXIHQBB2M6wuCKrSJUu5LIVD/OS6azqPlNFU+sZQ7cw4h8sMQzTynyak6eQx7Y6L6otSh
J2M4fmqP+FL2S1ElN17QyKkut+AC+AKo+D+CQchLaYhpI4ddoknEgw1jjUav2Xtr4Z6Fg0eD2YQL
f0arhUprY9xJ/na9dUaR8n8R7F26KhHLDI6MzzZzKB+Rdf1LU07dfi6+f1Hfmzf8tNdk05X8jdDO
htUHHvBpFW+9NGqNmwXnHhLdmPvZLyK12I7c2dkRfrZTHy79mVBKzgLrsTQ14NOOt+/Vr1gIkP41
GTN3JgBeToZJwO9DNOLmGyeWs1flnBigzn0X5jJuJiVKkmCfP6MPH5qS24kzTBG6UpaxLXnr6+vl
8KGTH/RvCTcdqFiNhYXxAsBlEeCH6qxlxKldL021o/hKIGGlmI5lmH+gGCBlFcM4B30jTtrCSHwN
BTYFf/9HehiRaLKulRF31eV7JWOKODwzUVu2u92aOnjqP+kq1LZB9mxcYEB97nAM0KiJeFqjkEJR
nZjqgA8HLt+uZS1IhbgcPBDmil5JCZCjkikNvMgxvK3YV35CqktJbBJsJA9qM/9/josqNsxGQU+E
/ElCcm8e6Ig4X6rbzi1IbN77C1/e0GT8Nsn0vozXDeiQuKNegBTWWhnBBo1PF/JC08Ch8k14d+Hu
dAxlSXfykZYwlWF0GGwHLPX8BtHOLzIcCojLrQQliUbqC4qfFsjEaccnTJzG1gg5+lvBjsftEgue
Q3RvZClqkKcMINRPwnNH/34OU7EA1hhjcQGrnPDLfzMtiCY4gHJF6pAC/ugTBD9mdvpiJJg=
`protect end_protected

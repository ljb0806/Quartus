��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��n�Md0u��"�ܖ+���T��	C㭘�c|��UX��at��il
��f��{m�B)z��LL�����{⾝4���Ro~��i��5~(=z�5��{x�I��]�O����G�(\�!�N����ё>�o���^cĴ�q�G�b��tLo���3�������%�FU��-��`�x:(D��M�)CC?�!��<	������g�Ċ�|U
Mo�F�[

-O�}��z��c������d\�1�U�5�� 1�bHw@����p�g3Ú��s��
�v-Gt�q�6����M [�B�4� ����,{�7kҶ�w�¾����3������Ƥy^if��⾜n��@0�p:Ӑ�N�"L�����r���̣�>��8!*�z�"q��Y�뎋���=Ƈ1E|wo��@�%�O�[g���c�='r�>G�:DYn�s�]��|��<��S"��s���s�D�j�}xdI�g&L/#щ����$�?��f\]}a�>�R:�5��EOO'�"M�-�������E�XD�6>|��vC�`SA(���bj����hW1��L>��I}�����vt�@K�����8��]��N�. ���=���-�S�c[o.u�p�R��[ʎ5{�\{.���%wTE�ި=5��fg#�9��TsЈ�0��$�"₝~{�ڕ�a����`ZJ��(1_�y�@/��uG�䓠�~��3�)��͘�I�D�C�3?�l�*8�*�|�[K��>�g"k�]�]�hv�c�#��� ы��%a��a��g4:�+�������V�������[�d�UD��){]��n�neŎ��
���W���ȩ�����8�w���sַ՚�}������ǧ�r�)r<u5N�Z���v/�FM�Y�Fe���;c�C�?`=������/8xn���G�'�;�:���<��J�~����qp��w �Ɍ�I^U�>��^ �61�ӽ�a�E��+�\���*DGϿPx�WBKV.� a$����J����P�*��Lr�Sv��K�T�El�u��|��1��C�A�͋��ӑ�L��k` �t$wי�������j"eɹ�x�{��p�9�?�OJD��۹}��6�%QA ����,Eș�d���4g���%�!X�Ж���l���C�5���o��\�oꉝP��N��d�O��etzl� �ZT�!�=0��+�qZ�Ly�GѥÇj�f��*�2[t�S�,�O�e6���_*���� �p[�	zL�|!��C]f�z��D[y8zw��W�-� Q�E�E��������	�U%�~��T�[���:�d"���a�S��87�v���B����H���4Ikq:�+�=�	�4N#SJD��oi��<c��"��Cg�jS�l��*����
�"čN޹!���[.e�d��ua��Қл@&�s�G��9vnC��5/Un�oU'*�y�zr0�`~�w���ş���?��N�>�=�a�׶����!�� c���f�BC�uoa�GtVXqM��8������
$X��i���x���	��'>�Y �1{�<.�1AR�۽���x�U�?vz�fuh50�lI�>>���*��涐�@��K:7ϯ�}
U�-��P�f�.�U�3D�&)�ǉ3�����ŀ�:�Ak%�SV��X�� m�r?D�3�V�\��J�o�u$Jvc�_7�f����6����:��h�MŤ�uD���Z�����Q=�y�a�ʇ"�$�94}5�/��Ԡ��d=��Q��Ў���^����&~2��1�Z�L�@m�9�B�en��4���I�=z³S�\:E^l��TV_H6ti늽e������4��=�=q��%�jā٩���ݡ`�
�zq%��s�I'�S�:�B���'2-�e�Hs۲)�t��J7�F�U��<7���iÙ�W��ܲ�N�f���e"����RM�	��Za��S��V#:}�*�/�9y@��3㓊��;����Ŏ�������� ��t9�
`����1���l�	��R~f�%j`�X��;���qI�����g��f%� 5NҸ��$�OJ4��/'�j�l+B'Z7,��j��gx���5ҏ1I�á����&�fq�x����k�,x���PB��|[�Y�|k�gЙ���P�k���,i�x<�r�N�3�: ���rE5l��M��0�Df�Hl�V���"@��k�*>G
+o�U���� �����F�OF+z=tf�w�C��@�v5ϱ�P��{w���6�w�S�i�+V��XW��_��E�d^BP!>��U-��U۫aDf<�K�M�t�w5M_w�R��}�=��G �����U2���zNs��>ݩ����.q��Ǻ���jEWi��-��s�� Y����̯}�Ύ�@}��S*�W_I@�h�˗U4x�Wx�$�!�ݐ�©��#ޭIj`�
���[5��M͊��l{/)
G�~�����
��N�
��A{#<y��@쌳��Job�i�mdm�C0/�̀�C�6�V�4�o.���~�� <Rz���=��/�^�r�(�HM�\颇���7��?�L��*�k��!�#�NѶ�ӕY��=�i¬���B|~�$$Z=�-���G������@���iP\L�8�(��w� r�?��{V�TY��R��A��9��l�8+�e.v<�Aơ9.��sJ�gVI����F�9����i�d6���̓�B�Q�8���"<r\�+=y�B���5�!���,n��ť�f�,E���r^��
n�@�u�6�,9�=]�RD�:җ�j훺 ~��R���ٛ�b(�7��(�h�l?�5������V%��ϵR�����U�ɤ�������nd�i�xO��d�����ڠ�zB�c��C�.Z��E�ʄ�{`&9�%Vœj��#T{
�頖؃��a�c�З�בU���Z�-cC�MLz��2-6%��N�/#�,S=Vӽh$�E��~�>����9��������IL�%%���2u7� ��,��#S��ET�/IeP*��-op��L����D[䄅�� a�y��֜�H�����<��Eu �vd~�X����mt��Kδ0�;~�B�&�x����/jL0����~�o��$9��=T���ɞ�Oc�`�^�F8Dr₍�ʓ��p���#wS\�pڕ*���M����Dp%���ůL��������N���~��͓'H�ϩUM8�����5<� �3���i��Q���+s��h�6ǧ*�����,<>�f禮!�YV.]�;����<�'*��A��ş�-��*��lϟ&1�_Xi�dw��L)�O�0���˹>���=Rj�T�7'jk�I~�G��g�Qǈ:�&���/�f*��������P���-N�8�p3aݭ������఑�3��8k��e���ۘ�G+�H�^�R�I�������-���C�MP	�\�1ֿ�j�C_��6�~��Ҁ��F��f|e��r�c>5�dj2h�.��A�M��._P��� W�f�����ͪ�N��݅��>��JT*�����S���mF]mMNy�%ITڱI�@Vs��8:�W�B΢�x��������V���I-��Se�v�ǨMr������;Qg��^3
��&IvoJa}�r���?��!�K��um5�p"�/�( � �`��^m})�y%���;����ǁ���Ii���Ƒ�yd�%����Dq��9�6̳��|����&C*��M�rWG���6:;{q�?߰γ^<����JM�5_�8����+�W�p<�˙�d{qm��h��j?U�p��CA��V^�St����`i�2*J��Ll���� V�}����u�o)������_fK��>O%J��Fl�U�+��	��N x���O�ԗ�@7f�ɝid��T��E�49N�4E �(�f`J�v�/W3��N<��T��[]d�T�1��đh+$��M��k�N�<��~8�N'5X�z3����!'4HALR�NfE�����C�v�cfi4��c�)a�k��q�� xR�eIz��i(�����U�F��ĕ[�4�Ғ��L��9y�O��1=D]�5a�:�ǜ�y��{ P�5{HI`�`� ��Sk�ߤh$�P��������CFSֻCc[����t��\�\�{�B��KZd-��ɧ(�F��;a�!p�``W�$��Bs2M��=���֮<^���yu�C1��3�7 z�z�L�vd�ȩ���V\S(�`p���_?��-�r�ߕ�Q_5�u���%�q�������k6�㦽̿�#w�6��]-5 ����]<u�����Fn���~�#���]�7X������ao�q�z9@��$�DX���dz���ue,�ļ4�dwQ�u�5oRkPE�?ٜ]Q$a��`̑<b���?�@p�n�F�Rc�׌�$'�,�L�#Ln����g�>	�MX־%+u����e���x��E�.���˯��7u(%��a��ې�DG[ʽ�whA�C`�)��m�p��5���vb��'�2�H���Y��ޢG8 ����=)���'��G��� u�C�X$�\Cu�F�оl$��)��6������~��d���/2shl~U��)�����B�w�o�Sl��N���KS_}�3w���n$A�����w��b|�1D p�l*�����2��F5q�"i��wpY�M�H��Ĕ�$�,�H�L���i��US�T��d���18���O9��_V(MS4�����ӽ D�?�NA�IY��bW͟=��������VW�dҖc���R}��B�2v:����r��P�m�:}w���ˠy��}
�!�:�d/�{�II���TA�P3�8vN��q�]["�Fzބ�̌�}��h{�6tL$�x��;c/��3�^�#;S�Z.fL�����:���u�1osM���/��ϟ"vU��~�t�`]�}�V��÷��ω���=���lj��1���.z��i��j�B���H+AX_�J�<z�S*]`Y3|�WZN�������<.�\�z�X�� B���_�c���+��l�.�1^"J�$Uh�e��\��Ւa�����d��՞v��=�ɋd:R������(l��!�'߀w�zL����;j����X@�J�A!�z����ܸ�i3��t܄�G���8+\��҅� ��+>��Z���ٳg>�$��Eϥ�pEja��?W����{�7��
���9��J�k�2�E5E�*���pG�M������rt�Q*���	�Tti�@8���@�`uT��X�:r�-5݄+e�~R��AB��g�<q,����_��Q'g/ƒj����׀��	#];�'�"I�0�<L�R�����V��*�7$���;��0�e�J����[��,>U-������t]KOm��8�
6֝z@�����E�v&t�yO�E��|$�V	����[�����>q�!��L���I�շ"���6X)�3�A��j.������>��Wl��B�x�\<䱄��hZ������=��b����i��Z~���һ��1#B�<�C1�'8k��1�	Rt�2�%���wrS�1/!9�� v�K���y�v��״7݃�JP����'�m� ��µ�P;�)_t�,��+������4�BLro��+�3��J�[��*�$�$�Z���k�h��|э.���p�'�z!�����qK>U�;C��Iz�ϳ�F�������J��OT$/9���^8����͚��E"���mo��W�ai���S����΀��?�-m�͋Px�nJ�΋Y�qN׸��d�&^�n;O��Cת��M,I��H�5X��}��vc���X� ��Fou ��2�:t�A6����Zz�L��Fe!oL�5�q�*Eް|؏�S����|�{
��E��h�Ys �Kb�e��C�`������9ԺS��G?��.��1Zն�sr�����U�m�����S+��xrQ�"���H�� Ds�s�>3��><Li��W+=Ŭ����D3�@�r�$�%h�|����Az�}��>�f���j^�f�$�K ,��g��X��s]�{П�v�����Jf"��Ȉn�L�~�E�����k,�e�����������(Ԁ��U�\�s9k׊k�S3����v9e2Q��g�-	���XS��r~\�oV@��L[K7�\�J��wY���%�X��vnds(�o��=�.omdn<Q�����XH|1e&�3�G�)U�V8��i��P�I�6|Zh�F]�xˌ���@���4Ⱥ�,#�޳�+�'�E-�� �V�s�ӇX0��$��} � ����gߕ;��q��o㮈����!R�Xϳ6/�|����k��Б����� ;$=��L�{r���Kn
�t�`6�o.��vK��C�,^G �+���T��D��H������>2Z�Q�(����^�^�ֺ�Fʡq���&m%�:��l�NM��Er�)Kٻ^R�rb�7:%bKK�1O����>�q�-�1�d����$�)���)r:^��kW�-�{~��!�߷h;ƈM�A�y�%	9"�碚;ՠ{�>�4.���AU��qd<~5����T�2R�c�߽���N
!E�z�d������ں�~ ����T��7j6�w��X�C�,��⠲��}�����`B�,༭�3n��ŉҨ�;eZ�������d�gO"��*��E����I�f�����>��Y1��K'���$��Dϩ��/!��"��>[��N,V6��������q
^=�Gw])�k!�%1��/�I��}����$/��8^�u�k�����1�*x�����x����(9:]j]6c~
��.k��;h��Ϩc��(ǘ�G�v�\��o�6�MI=���;��d4�D3���7��s��i�;;o͊Ypʈ���kh�AL����`;�]$�z���5<z �p��>þ���Aai�6ɢ�9�P��	���}���9�7���H��R�A��E���h�i�)�t���ǚ��о׈���yͥ����2��?�0c���Tp1@�,�9��G��LN%�ۄ^^/��L'�I ��
� B���T��Т�fu��ͺ�57}�� ��@�e7��m��Êͽ�| �4�7����>k�D%���T�3�L��N�?O1�y�C��햦㾳�Ur��<�og/�oţު�ʎzJREI�R!V�E�G�]�̶�<e��ć�{pA�2%��̘X�8W�QX�^�²�4Cf\8c��&�Լx�9o�WW��K*9,	�Z�_T��D��}�ƿS;��8�f�`��	^gf5K��ɑ�G��|��Ǟ슁4KX�|�����n��|Fޒ����������x�f��sP�>f�9y�ȧ��>��x*z���}9�j߀���8?F���x[D���mc0��G��(z��86��C��K���`O�閚�~V7Bύ�"G���%�&@Kv��-������7�����G23/���{;`^�p��i[�V�|���<��z7б5�-�[6�yHS$��-�_�c�F�{䴨,��Tvd������V[�eH2�þq�si����'��䋎�����=2 mS�����
WА�֘d���ɏ�c�$�Ԫ����*�+�׼�E�0��k�ccT.c�]���D,��qޠ�4����#P,���N��,DӼ��]�I�`��k;�ޒT����ȧ�nT������Y	ܷw�n�͵X3O��ӂtUV��G���(�
�c��<�E�z9��Ì ����j/5#\�%j ��2��g�&�*�ׄ� L����.kJ�z
�u�s�����s�@�F��:�5�sq�+�HY2շ�Ap�n�g`'�,��I�ֈ�{�|�G7�k�	�/�c��J
v�����k��z���o" ��F�O�3:��L<���.6 T,9t��+&�O��uF�������e�Vvh�+N`GYFa_K��ƘD̫�nW��������~��K�:� q*���FFo))RH�W1��������lau�2�dͬM���B�;]VX��2��(�̫\9Π���B{V�w�+=O`�=#��Qq�>F�t�7Gvxz��d���|y�o)!@�Oˠ-w2�(6y������!#�v���۠�P0N2}�r�7!�����Ǹ)W�-G�d�@�4��;x�b���6��������X��y����`c��x+)������&��	��2vM�\�v��z2�� ��ph�7��;�����v��p� 鬴�Kw?��3D�Q��E�׋���Gl!<���I�b:ۤn�ԊD�߂zЂVQ8��b�Z.� ?���B�>�d%��k����hN,[%-U5��֜��"%���Ϙ'�0��O��׍ �5Ra'��i�}���N2�q��d����'��=8M0�B�h-w',��5Q$iưm';�17��48`#lc�ׄ�\l=r��Cq�,�E�LԈx��i�O���Hg �Q��5|b{��T6$v�zK�V����
z�[=��;6��R:�>sn�_��w�����N�_�:C	�w�Ȣw��d4l�Z:�0��}�;��"�*I뜍�����{)�'p������Ɓ�Cy��e��h��YgS3�Z*=it8Z��6%x��DUsP����T�3��H4�T�+eTf������k��F��V(7x�H.����xu0�$��ɒNT�I]'Kb��6���3�V�Ȑ���}D�t���=�^�9�f���3�o��T���[�.ǫ���K;���E1d[�b�����v�V>>:YÉ�&	(#��vp2�����Z,W�ɲ0��M�lw�~a8)9ϚCWÄMW�EĴ��$K�?mZ)�N�|>wC��)�����R@A�u�7wT���)�DZ���h�6�p?�o1l��łQ�àl��An�x�ty���k�p��Z��X��o���:QfH�� �x9����D{;q[��Ɓ�(������!�~�j�t���]�s���`p�D�/�"�z-!"�5_G
-y�6�0���zHT��)J��(MQ������2����[i�0^~�ȧ+�7���VVTX��Ar���PG���D�q�i����g"˃G|Dm�'f7��龹�]���#��%;���N��0�m���l�[�څ�����Q#�)R��yl����&~�+۱,��K�������.�M������0����
L}��� kݻ���L
7<n��:���ҿ�H��X�%�v���c^ʁ�3�0�~����f��1�*8S�\�(n=s����&\�y�>2#�uf�%��?����@�ZLc�ґ��ŪX*�䲵p�u�R�V�B�b��Uq�I�w^o�:�f=(�!sK]wdF��3��ug�no����g6������Di,��q6�!�J�Qg+�������k�]
O(}��vT��M�7Q}�F�E��	[4Ԑ�X��[bD��8B�"_�1�l�L���[Z�׀1C�NB�I��DX��Af)�ꇸry��Ō���v�'X���o0���#'÷:%F��1��;7S
�Ę0����Mru����hm3�-n�?}?�Vq^�o��8m�S��w���7�{����sd��A�XF���s��^�X��Í���/� y��`��b����K�����嫛�קCy���O�n�'l`�OPo���3	��FS��`�T�.�AHr�ӚU�-R���5�g-*p�/� n�~v�����>�}�{�ȝK�y/)+���f.Ʃ���8�؊�����<y�E��M�ǋ/fG.B/��Z�<X��2�p!7����B\1���sv�P�wt��W}����P��sͧ��"�@�r�w9�<	�
MM��A��$ҽ{����^��B�S������c�e���N�Sԩ,� ���l�C�Ԅ�R�#�5�c��e�v�K�i �9�
�Ař��Fa��Kq�Ռ�g�>��9ǝ7Q/D����94���#���/��~��� ��~rDpv�5�F� @�T7��� �WDMi��d>���F�3�b���鸰,��n9S�����Q籷G B����B&�{Ž	�F)mA\�;/�K�����\�.��'P
�n�bZ4A�`˯�D�J�k>�Cֈ�yԂ �U�PMJ�hD�k��c=���p=��k�j�Q=�\A���d������W�B���,��[}A������OT́D�{�SajA(���}�S�	�$9�+��T�U��'ê�S�E:r0W^�q������N����M���T������Mar܄��8�)+5�p�=m��5��{k�v+d����@���y����U�����V([�jxb��_��־������_�QJ��@�Ǩ�2U
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uYU1MpH8QneX+0WbpacBBp3SB3A8s1drPrW8ccCvwVAqleDaio0rNL+rWM/I/i+uWM/FvUjgHp5Y
po6GlvrjnZbf/8AWlebcR1ZgBkVc0ZU/4i3Af6C1Qck8zfcdAxJgwXb33H8OTOqB0VCHHXAAY9W7
hcNpMWChK2LgFHL7l+PJW7+e68granDdsXqVyP5FJJr3yMQ1Z+jaT5RYtmsIPg9NSjAaMdRLVvaL
cXnDqEj9vcWD8LYuxmoH5UGCJNwQ/TEdafaFG+be0bLc5AfTadyGmKxQqZSq4yBJ1E/wsymLYcPa
rvmBmdlJWKcZ4PyaHbNHBdXGHLw75MQP9V089w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7664)
`protect data_block
JlzE4xWd06aUM5+0edCM42TgCvmw8mXnlhTv3zZsryyD+jKT0FSNpGkWlIuF7wYXDmDXehEx57cJ
Fm8tzBYR8/LQL7U1RufISpZVuDqkmrRyCRgt9AnwHmvaG8+Cfr+KoTz0IHvR7dS8V0wy1y5SVint
2L87xycIkEACIEYOYY6zOwLCGpTB+Fwaa674fIBhGWY1yUzWeSH1zgqy5o1eBx/lfzCGmV+Vw2zG
Xyb8AD0Qa1TfsLvwujcelW6jrfLfBtmjkPClFYnu0cnbWzVEdwUD2EhHbjgsfIqFaX2patppl+kQ
bIR98/f8lha6/KZuQStjPlLzUy+DPR7r6oZkHeZXJWqf0bAbzLNrAqBDppPYrTIGKHIhXCc++jka
KNKhA3gfje6700L7xNrZnBQnXeLO6TjBBWZZO9mHXIYES8joRd75dRj/X+AyiWmLYGVMGg1OihFn
uIzAzfxMM1Q6vWEIEiCmTvPdeY5/0TZmKoEAyXb5hG0rCBQcVpqVM0gwt3H5RqwC4KaMfEZhU1f7
jDrFtWBbKIyDAN5Z+AKs4eicJTgCNoRn68URw7IUG3r4NB4x9VB5wGM7v37vEpybGQo0N3C1AtVV
q1vYrxKO2hetLou8wsOwYUdzduiKhuKwMrnMyF7Vz6FQaYdz4CX+GN2X7JjU8LKO2OoTfC5pYFUQ
E9IHUjRWBJek+Noh60pa08gOUrB8z07dPJB/TKbWBYEFGRB0usH5TYCoWTNF6FUrtoAysFFSXQI5
LllwupJlx3wWygxUdHPwfPoNoiC9OjXBa4btIZAZ3H2Us9pR71YPjvR3lSMjGTWvQ9lsCzqiDZQO
i8+Gm9CJh4R8IU9xSKbTV+lFOO2FP6Nm/XF+np3mGZyoonQTLFwKznmovNmzH7BjgghH3Xaqog6M
va88ZBM2m+EgamBJ4+OjGX8EMDfdc7bVIup82oU8ktcg5UChPcuMMW1SIWQ7iQ3vZVZEiThqzYE1
Fq7wyAx+fjIs3VeiaDUObPGFbOdlAWPFrCmrRFchoiTKM4XdYLfL+ElKF4tmQ4hclDd9KRJXmkkX
82YWYP2086FkEiLT3qlAF7g/bfWm6ups3HBvzzh5awbEQyzBCFzJkti8JesItqTitN+wHM8ldttY
Bz4s41Dl6JMjKJsrI9hdYDykLLBioTFVbgB6Kp+ZddJ9wZXg5cTA7sUL4BMjTJs9cxzYXu3n6Anl
/ynqgtzs0lA2vtIzXbgkl8fKklbGN8AGvNEfdDDWkx2nR/8xX9otO3OhlaxqadEA7pKIDdn7s4/l
4Z1BEQS+LHFGMXL8bGLTivUKBA6f03yT/WW5cqoXOhZT+CPePcW9sJG8oncEBBQVi66v4/+4jvTE
sy5IaG0Kp9aBU+UdFiXR8pR6WHRlxvPnbA8YLdhPvS+1QoZzda22+DClUhmdd2LLgfc+BP70+riC
2iLfQz3jQIaQjm/9t7NqKpLi868wLF3c9Rn9qA1uxTa1Z3zK3YLf18YGV6NrlMzxhluu47MuyRq/
uPnO54S2zg/K9E7Gjy5Q/uy/JUZzBO0Gyg5BznHHaQ0S3li0yCQYI1e2Cw0uHZlhd8yfTx0c53qk
DKx5ixJX2SM6Jil6KqF/Ua14xOIdgHz9IEfDtPoOQmFnU0E20i+Kmv3US1/HXl42Fytj1Xhqko3H
/tY57Gy9OAl6452LWmyOaHZmEzyWDIl91hBIUUkxDT1FlhZCMrCpvZlRQXoWEfM++/9l1bxjRaTS
amuCP46hEthzuuYOsShh6Gs8MR3L1bLGBnsVdrPi0tNlSuTZrVkbR7o8FH8fzhFPXBRH+oZQ8LCP
uD0gJ3soMqgtGYRz0z77Udsguw9ylQh9DdhNgKyilXtBLwAaNfwjfNJwLxEEgJ8RvkGd8YzpMRp8
HgB62EJyO6ABUCpsNH7ZydPGDJCuGhIUEKJmKBTHn1plpbftX52tojF8R6dx2CXyMuUPih/9pL2w
Y7LTu9rFqYlBLg//uLAhN5bNDNbXacMMaKTU8VX0PvXwVTWYTUw1iBiBO0TjjYL6zA+G/d5BldaE
8WrALNAEVx/VsmfaFREe6dGbZoarqqqzrLFkAUft9XQ+XxyoPnRIqa8MQDwvHiHHehT9dL1M0wkz
tBFgW9rXiNQ8bcQfnbl4XrX/kLHevc9DxtVPz/LWTl1IesBNARSQ0GVvGlJ3sb0IUsrrALDM+iUn
YsljypNl7ZkQ7M8O5LUwc7HEkTGq4d8+Uvaucm6EV1s4ivcUx7dwAPNnfqRXE/jtSKDj4i5cuSPD
N/UwyBWWLFm7ftJ5FGERxkwwdr0VjZLcvnBWl7XX5DHraVtRiY3ijOAj65QHKex5OAkFt8Pda264
Id2EIFgAxdh5vYWijaxEId0TqLN/1LE2aOv2Y9qWDbsU76HGLweOUZHEyMXRDf0IOAz/m76Rpy3P
JuwzYouCP4xXOgXm5qG9r7wR6j3P7uW4Nd6JHwVgw6zA5a6n5YXC0Zsz5hTcWqFOJnvCqd8rGGF5
ltfMyPhwm8sUcq3z17hBbvUzHQZSvYb7FaljQ7cs6zd2tiGYFqlMWQ/sRPpQ5LW35EMvOoV9GR3s
YsDYlqEj74ANTQ6Y1YNk8JwNowsDho3S6pSJvz8RBHvIKVwJ6CgBVpDniU+PwpktFG2zKF9A7s8y
HGIffe99D/7s1fEnswKCsRwggwO4Q0lqKRqw8LVVu0zmh3mWW7uyEVmDPN7vvutahsKPeOJl+jcF
kcG7MQ6pVUpOAS8SApV25J48jpAUKPEEckWPwq+PqnqKrQdfuprHbACbGThOltQFsfsPqH9JpgOQ
iNdTxtdufNchD3aHQBw0PFsWbRjilx4KMLq39wZcbVRsw6Ph7DFoIfuiIxUADi5dGXpAsM1c3cI8
nO4VPI1wwgqYJE68MseQPwCfKX1UfXS8tZskoOklnTROTKUoDeLQ0fXx0Op/JSjIUrP2+P9b9gzY
RRxL58UlrFVOrCr2j22OJXmCtVBusdxdgmvhD2lfy57RTk2uo4Li82PDx0FDPnz1KiVjCw9NJ4L9
c7CCZbQQ9X5xDRS/62f2Nj3XgIpGrw9ir1l9+Fuqm6xdnNA/tDeZMurdq/C44zHHgKSMxr8v5RKY
8TBO05uAXmr3GIG1u2Zmk0V0glECqZx6h94dLOVCi/UvUkQxP4ZoCqXuA9LWTTrtEvEvuGNaAj6x
n7S+MC9bubLvrEYUFjFtnFSmFknBKRFQrygM8XLzPJGoVxgixPVHWklAWOTpMq4FOptaHOlRA/fR
jY/yqW57TsAlqE53U9tMNctN2+1GVr7vceGge2Ed/BLRR+Ck/rtVX8rVRNoUYDaiD/i2871IQY4V
Hy9cLyAWILDNb2Eip0/dLWfuts8QDeLj7eE9/CXD+jJVDy5B+JMqtqhHqkzbXDM4YG4VpUIWQdq8
JDN9QM+jcx27I7Xo/Q1fVGhdgr7qwCDoQQkbQ2sAaBv2bYvvzSvAvi8Zt+gyUjh4CpvfjsVqdUim
h6ehktLnUQLtpqxXgFFaxY7NCrDgWsD9XRpXfd0qCRFkeIFkM4AOvPSaiDxtQ6xbFsq3j+CK7pQg
z+JIjfvPrBZnh7sQDMDkrUjFK5fKJlPqO4roKVqoLCytt4IMz24R/ep0oGln+/pd6gtf2CN9FbjB
DXiPYJeHwup6djaShfpBTHfCHoZ+EoXC6WX8JM38g/oq8npbFFchNUoZWnoZrZUkfChgiUN+sDZ3
gr4Tl469gO2uJ1ut86YeQ8NIAeFnXICoXEYNz2gR2KMaIAqfgBhTme0a7dpGb4de+4zZTNRBM7AX
1P2gi6fgAKuoDba4H1fIDitbIc5FPu+KgeBrNZNgafkCByLqJh9rALk4ztbwxpRBZpdR8cwDIj0W
BxFBmNnFThjNsKfAW3mcKmHLwgDWFGIqbC7GHjFSOTtmasBGux4QFflqp3xa8Q8a2y/oqfxgDUH8
AkxRMemVmITRR5+lmX7UDGH1oMB6+LnnnGEyWnBsg4KweDa4+CmV4/VlkJozacAnmqa6tIPMuBJr
3RwvDCEVlNOs+u1zvK0ag40UY9XlE3EYnYmoLbg2b9mRhgB3x8qlz6yzlxIZLEr8XYrjbZbiYvWo
vXrQuUGuubbZn1szOsKPBNUCI2LlIfIe4K3sMTZp1zkRMWzdyWup3prp6ByGteySnf+COL/BEtEM
YRHns8ml34QTgMr7y/reOUF/LcX+RhuzcPCCzsqnxYmw+0a/yF7lnnn+bmbbOq9Aev5xMUcRbEWK
z+01SuLp3nkdmnAfvLl8e6U/ogZnMr4G2/OL3ZLIK+WvH9ApJtPPnSutQUHftDp/tQAgYFaeSF7j
onPL+wDA6PF2AdFH1KSosSqGD8Pzt0H3eFW4AOcpImNAtEeT/juyyZJh8VgoJdY7MLC2uu+PT8iI
rd1Q+KHczPic118ZKdc7WFs+QkLSt78avkAj/Wj6E8+flmylfSMdPLBpOn8LUYRwq9XFwqClliNs
tRBznzHkpcuoFBjZpMzlUSixcf5WZEA9PjnJXfhIUQhD2yvoZSoumsnQ2HhA5Ql1mpbSrMfO+8b8
DFXHWgggLPFnYlH0/oWPaCOOD4YILPj3ilvoMGC3D0D+D79NJH8xEel18Wqb8tfvuL3bolwEpflT
Mz9/NFnFiOFiKi3tuejG1rDKihGdNJRFmBHtFdJQcYbVdwF9ODbDnbedXwjmgcMDbjIACkuXqdM3
qM4hZDw9dpL/Lj+VwA8eNOEpX3glpG1COTNWe7VsQ8zrvHInIZALL+a5g35RqhVoJ2aQs/TJ36uk
Ak5ukI80AAheYUQB+d+OxM5f0RdJ/9rCzntnZrSrjIWJC3wD6XRHSuABpo9YCeLHtsIJSLpGzdwd
R1uSHwdpgjp7DQNu+DLbQrtvZO/pXpTAZ/itiV7yOOOvHN6kZ1zPXBIYWC6sAj95nep3oeNzAFe3
lU3BKz466A9IoQGUDzuorRfONRhJHNzdzx9w28zzSwuzGPi14yrMKgJNSmr0s9GaF0SS1gaWQ8t7
1XLApUCu9zo+iWs2mBjInGgoV3lUEePyfWw/ZbnltOqjV+CiD3pjGdpadx7DNOwZhZvYyjuwon/b
6zbVFIAlfq7BmmCvgYiwTTj6tYZVi+sX9Q4YBa5dB98fC100qRZfSf5YbhCB1ekZ4ZqSA3nJGsuk
LAzncdrTka8FU9sz9aSbqNOYeOdwPDgTMxAh27tW32cB1qqZ1wRCJ97KdneOKivABee8JZTh+tVi
gh2jxuBtW7PiDFjFudgfcex9tMExv2miPBNixppltCYKzGLov3oRDqdwuPorveObQm89JGXWqS+W
sXWb1fiC3MuTIWsWQwWqVWte82BjQtMwD5LcLnl2GE0eevRirmpgnJZppWYVj4pHFNjY7mS+M0JZ
MFQ2i0Dz905bi0j/IJudHtYhoyCbX9O0HeHGfqKjw6FtsZFMCGlYRN2u3kkRlv6nQHKx6FEhHTB3
qM7wo63L2TvfAnq46RKelf3QNF8GBXv5FJ5me4jHWRUg78qDeuATBkOLRjB8JHpvtGbpd3upc5Qi
XYanPzdK5Wt6q+CEd4WZw+lyGauJuYvsTXsz1wrW5qD6k0ZhdfcSGtHAXLkpZfRX4zTpMYOnrxGN
eSVoA/AadbbEuzUmU0tzxH/gMgrK1Gg0A+QpwGBXvZpeYsrkPGqfcBv55St0IFiiim5Yr+tDRDaR
V/vnYo4k66Z0baUp2sSBmx8VEd5a5ZaUGoWt4DhtisB+y3icsyqVBXFM1LlaOGr1HLEptMdOBZeO
aCi3AT31AzF72WDAqajQNY1Sa36B6N6wcTdpVZdqvrZhTmxpVkHW/RbNnRQi6PQXqSnviKh1VTwz
UjckMrmrFPxPksDgDOnJ+e70F+Wcsoy1CDTAiCATLfjLeTcL/AHTsPw+znbjSPHYuzZY37WXcWji
y4Q4O9t9vXxrzSnmFSJlq8HKe4MOegB5XzbJycwIvShMcunHancanV4SCnjKmlOgXYUtv5MMwAdd
wlCeNLzHpe6mszEjAjWHCk5gHsw4Xpu06aNq276ow/B7l351k6CqgwMESSfxhkSuzafVAW/w8/Ql
DggJ11OsZSKXjImZXqT0JQe+HN4PB+DfsLEa/mOGFHqevYSCgyIKSUDEqCx+xX5LSIHgROmNU3sP
DtCLlrf0yn0Llt8bE3o8mTl9kAQPuA8AFj+B8rjMxMdw1bHN/vQusgus5SjmTr0845JRRIAkwXzs
aAj8QOECPnO3RlTP75Jd2lBXTKhaCeFMVkvSK1zA1XAbsIuxwlq6t4LtRISIDm9cDBPFsUMZJQjt
k0sdeqM++ecAodTZPru31Iy3UvwlBkjtTFBJEXR6fRBBlbJYoYYjYJ5+4WmjKc63Cicw9S6fTXyX
0viKMA5W3ZFGk90TwPSUrq8xVI9kT3FGUfuZp1sNp6n43AWMrmd5wP/oFrg60rNA2A+mRxzmsGDM
CgsVcJfItpP7eBY+9+gDmY4vFweLuf0fdGV+TCw470PvGWAWct7nYLEQ9GSS9e5sczouyzQP9S60
0cJ1F/qaYbHWJPtIof6HOvpH0vhe2aUUHdSA4gPANYo1yoOC2qy7E7547L3TnTnO++SduZIE2AVm
z/4hdAOWnLCGzUhuJSlvZeTNFkCg592uZz8A72iKzJsKp9qnJql7twuFKXIEtw608kwTTSFWnETF
rSoOtsmitst5s3TX1X1UNL+HpK4/iAtd49/NDiaPPgXBG+WEAZ6nRx6mUZwO2lJ4/+ob6FnB6uiF
M541uoD6mfWOBZHjT3bqnMaPUFJzxCptvAzRTvxbsDTGkAHe/MGEac2+NDtYt0UYLNMB7mUB18es
FkmxbKNyWaVV7qQNQeiZUO9MhpHIOSRPA4am+AMfUN0o//Npb/9t0fH0kHONBe+EbanyiWLo58Bj
L9cf6De8ScgfZh9OfAedK1zRMSJMI/yb3Kuq2FA/KlukrYFeDaeC9AagoiN3cWBE/NrbDcb1GPjC
0/HvFQLYT38S5Fukw1JNl4CwsLn99hE6GU01whQ39SQ00NigCCUJzEuEIJIOc0O+GLdfiqSEi4MH
3oEZRFLjDBBugZmsOKcuheFq6OSdvivc1ljBBb+Q3wi4CORIEjcuFG1I+MktzXmbJQILi1Owr8WO
qrGXFmxPoYUmkT+ifsDeIVZJ+MN0PKYSoowAX995P800gdh93XVcwpZtfmOXdoJS29XRNbvX7oVW
MxZT6evWSGRvRV9VWpzsEXW3BI1MxC43Sy6MCKe7AsJHe/FS24DPjDtYP+1IJokx5wYAfHo/HVm1
Z4VgxHTBFg/k8LDT4UaimN3zx4fFWkJOfTxucVL0jmXCBpn5iDn7jtLN3iXCD8WYidI+GGJhTXQm
RLFzoKi8UDl5526o7/pxLzzgdnGgdBYHqotTsQ692/Q+JUybXnqyQBrcI9NV881SidE2GK/Reuyh
eaET8dlCMc1srpykZRpSdaX0apab6PY7JC5d+reigR4dmXzETGwESLxUjKtmVsvCq7wcLkNfGflk
cFwY+GYq7Wmu8bdBNiwfAj5MbYTJmCaffVrvP1UPc6I7+FBNeixRn+1omogrOjqeqvZSegbR4tOX
CSM/OpiycgZuNPo2Nn5p1qDoK8kORXY+9BnSzFKBcvYBhkiZk1bunjeQD4h+NVH/cV/OxZ/Ho5n7
SRywj4RxlwAx7BNoira9F4McN1vTfijFfdvYV1ftdcHuVwbNWHkDWv9mliX/YEUYIbEJH7BORo07
WrlyayJvk0q8okOjtMMK0JlcPjW3npheac7sQ9SSbN0MqeElr1Yvxcwtfkgw4rbwQISrGwfL1FUQ
8ipy1xu+G3NbuqnryaihU33FQy6cf8k1uxWW0qVNIZVmdZT1um5TtCpkmx0JK+3nQhDNHQDuHlxp
CLZM0fnaWF1e6B3oHgBoRmFl9YugM5SGg7oD4waP/bxz7bVxVVEFbJ2O3CUGBwJ0U3b6rFRdsKZD
KtmwCccD+ejUZRMuFstYpQnGIBWzYAmzjcOW55gBHMT8y22sWYTzZXg71luiqRjSjBVfhyW7R8N6
LDG72QRcxgKh1lPwyxenvgORGH1tdhAcX4simjXpxolDw+gAFJNAjojNce8zjh8EwDampDol5JU+
pDbHRCzCj9n3DMVLKeVh0sXJlS+3skzvNdjgiSLD1bYqi+fJFIlqeKA7+1vTdT8m94M6m7HsPKTg
ou2+p8Bu8oeG+pSJTSSO0RlIzf60IyIlthnSPjc1AaktLndwM3F2Qxa1/pReVRBrd6l5XW9kS+9D
20XWcJBURUrUqVvZP+7vJisnSADlXFBzygJB40jBCjiRMfh5c4vLyKESqxKwrornC5YlPUcb1gDQ
xlpcADW6pwX31YWsemxX9XjAuAV4R/5b0zBYLYsRgY2cx60zuzhpqhWE23wRQA9OGNv4NX1eJZ/R
bAXtPQruhQ2fgkOS7Ni3eRX71ioO8ziyRrsXFPEVk9PWrt1E7n+xrc8bKggd+bHo612AgttWLado
q8DewwgQpCmpnkT92dt141MtDxA4/pyNUkS4q/SvSvzO7ty0laOprDptHplSC+XaybuEzBFpmaOV
SImRKBukv3sP81FjfmsQQwtiF0CbrEEYU/ZKXnXcBSfsxM8O7KmZpsX4jmye3l0mdbyBNv2b6orN
SgENFYltbE1BBBzNCFolJEnz855m06S5jrwHO1vwUtdQCj84V2eF6SBLKV+pijUY4NtxZxHOhKRw
RBDQDU+zaRjQaSi9LjHdPWtw5C6ziZiJ50FbnUoEo5HNu5NR2q2VTzK+krzADufb+10CiOnr9wB9
f6tab3qEyI0N/QeQnzYq4PmQK7sfWcLbIbUc7g+N5YwuEluVmS+IvtD6VsJmQymW5CXB3Ybupbeq
YcLP5nBQ3YDhhmMAfmANpeICRmqhUUGIubQaZAQ6PmhPms+0WOMROwyHo4ZtMU/kUpv0FYnyaetR
RTb0fGW3qoKIx3bznVK6Ra9RzG+pkeJWNoHJBJeW4FHIRxYzlAL6EhlA/Vmrs5uvyGp9vTD7vVln
dAue++/g0a3HT6WGEx5BXyEP3sbOzF3uwPRx+IgvGQEva61VLSYxgw+kLsjc7gCgtBpwhUmcMG6+
pYEtZXgpL4tCFlV4oVfcAl9yUSJmpebq1TrtvO/5gpt4PerLvSV/5mvjbiOl8ENfAJt1s31/Moxg
yyKcvWTOiqlqzhYVufE+Pqqs/oh+p3F95OOh5Ix7CYyHo3l6p7FCbmdpfUsFY+ycwrZ8WhawQX4a
+TcJ4D+MJmiJCppVsahc3hlvIdbiJI7ZZjNdCUnPBSyRddGAoaxJlcNq8d+hv13Cm9sGyEhKrYF8
8CowBBQEEU3OTDbJi5FwWIw6zt9UgmXmw+eAi6PsnLjCrpSSeOCXydiqwh4v7CMWGNTxSjX3kCFN
82ByFo4uM53x743vAo4C8pOPlk740vCUWE/WaFOx05C9OBR3rAJPt2AW6OdSlDIwgVLja1dSQvQ/
LZKgCKMD5ivYZlamf0QBt9LbidiUXdpNiGtvZskrTiTqMw7tf+MRijWrK4BXDhCqH8HniomWZ9HG
yNN4I24gvD1wHO33E6P05FZkcr4/CMOd9d0KGAL3ajK1FiqyOqdGAQKzskIQqn88VRYoXLj+yULX
pTgRUopLtGWhEsGneKOLSdVejyc8gXpMUuE74xH50VvQwbZyj3y0BHbXQHGK/a5yACYBmXLq3bL9
L/Jq7i9hZRXRFf1PB6yG70ONdSEAfshhH/KeSkzVzHWfCuJNcUUNTP0Ru3e0E/nbCI7A0ewmhsdw
URu0rv2oSAzgLvZ+3WAOeEyN+JSiJBj4LvVmVAbz9ulAFM1ying71+Yum9leVsNVuUJM1xDoXELj
KFDu4IsvoaR/C6Fvwtc4uG82HwKO6soJfOp4fqAfgpcrEyxbMw13KfOPpxrDK4adkDdhrAl1GUYg
1fv+IZ0McHopv/08anv46QpW+tbyfxiMTx7iHEPSBQ1SqvtobVtucExuUA/KJxilFkB/erBASGe2
uZvOryfvkpgAeBVTEGNk7vYWNOtY0Nm0/Q9+DKwJYSyERgp7luU7RGWIJZPoqT8GiJZOzHIg1FVK
deb9uCLw5HRxemAYbctX9dlLSMbacf6jvrBQgRPkFKh5JXHAGLhMHXddrl2iD+nmT7UK5KQAgKsP
n6EkOZ0LkZUtqwGfxAMOVklgiNzSMnwdb0w=
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
z40P0vUdLIa8Nez1Orejx6KPdZxZZmKQehasq96zTRKGa4mlDX0EUHfGgvgiINgiVLRhvUy8znB6
oSIZqTJZ5cukn5YBUsxLuw8zmhQoJtqPwzYgR6cCzq6ShhtcR8TjquCblNElZNXb+n7++7qBMlUE
qynN8EWWXwgcd5cqMBtrPsmHib8gaFM+RWx64FGFXdiTGVboMumKz5DDSq26Y10gjlMcr6rpXOEK
jkuZwQ1f2uk2duH8d45qbbz37hKQA55/imp8C1mXl8gk0oHRRaL2d3Yb898qKCZCYcbERnMwCAN4
LGUhQxNyD3qqPJgPQvxOOByuXv30h5rmynbofA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9600)
`protect data_block
royb8c3jbAFhx7eahpvdQc6FH0J3xagrrno9kynExmQzSJfsd9aCfOn0fvPJdpL+tnqvk8mYvM61
vPGKP3pFPSA/+fL6yBSPK2FivnqkYHe0dp9SrVBXera+nFsMkKMg8eqD5U9Sy/9WRP9nlCG/BeFf
ZkNWl+M6JljzXcmmlUPRgLXCc45dHDxNfjbWF6TjNJJLXpC8MvZvTJffRoaRUjsKMxNJAZlA9wEK
5jw48c+6qNuxMeMz4nKMCR4T9rMVp5BKUiHFUgWJ58i/vwLIUHNg0K20ZCjwVxzPeG5H7EPQgttT
iGD2KdSWVIVl2rlXToSkl5FZNAGKqqZy1GF0+O5fLETSX8MgUDxp7GZORJw4o++3fd6WlIBAKTl0
ahjPSfFVNoG9admbYb2hRZ6STD+mNd9Q+4fBqAolTq1H+QIGcJn59qJul2gRi0iBnZkaoPiQZi20
5Rt3HDo/AJqyK6xCIdQXMj0NGwsYlSTrBG1cxKAIC867JeQnvmKQvVGGZe9sO40T7EjvIEQWjyLs
X0M2Dmvd6VVPzTXVH3vcJLT20dP64cE4mEsV+WDXyZLwpKTzmNwZkZGCr7/u+NNbCfj6SAF6I502
pii1xlDJuZkuZIxY5khaRHd5w9WiZe9i9tpuO6n6qhg6R2SzDSbQOeqxHArVmseZ5RZcZR2lId0x
bzGf+XDArW0pCzJLQiZbzKKpXeZTOTIjNpeIk9REzRfBRDZnKyHrHX2UYTuLzvhcXoDD7p6+DCWp
29ioN7iEjZsVL6Eu5/G1G15pT7JlFMR1UGDwXUjrYS8nIFPeATz4ztvj9B2xv1izQSs9MxMuOs0t
bhQWiMi4wGQsEdlbNKvp2+Gvfdr8+H6DCW5xtoCqAkMunL/lJEyKp2AxLCf7WrBiYPXsXeAKg8yN
SvAuUyo32D3MisEmdZZtYtht2/juXUVgYU766Qw3wngVXRVjrSZac43F8PwPnZspNLNwGSoNo0Rj
TTBn0B6GgbwT3DvWriY+0kCMLUJOc4YGWg5eJNJZ182Dd7+DrYCgDKKwNQRHFEi3pgTktBcQZAO2
dS+JszhayYBxcZKxkyAYOHuUKkq++w9dGWoxb7b29hLwuZIZXLwHB/HsT4EXD46VS8vOu7ci4095
vOgRk1WuDS/xRuKCt2+o0jkDp0m+N8OoK1c7cUzk1BORn4uHW6KXY6EYwXAfi8cuIIkl3q/VO7IN
1VFypmJ4PBRZLtsx6QilniC3Z1KmggwNdKx4kUTyrQDRk0QjcaNA8f/T0VaxAe+nm+d8y6xMSSSB
u4OqdJVWoRRUhuQ0MnzZALrkeDiu+0F6BNCsSskz2LZWSx+YPTAXdKODBW69LpLNeFuYruJr3N3u
gT1GhsT1YEuu9Iz/Fhh3lCcaGiLSgrO1V0YHijl4oyOyLdOCK1pzAB5lRM9e8ifRvCl+t7P4kouh
6WcvqDFWuUyeavVkf2Sgp/KEokmDZXXTknyBKswwMHM74pn8ev4MO1+3yHdd5iPruND6O2H3PFqB
tWrGQSaNWSJjynlQU9py5GblH4+vsa5vzRmTlEKr0rw5vYk+Xv4uEtFSlAYGV5plrr8O8jXgx4Ro
/DiWLjubWtQGzTRhIVpDYTBgEpxlX2wX0cpBDvhuX3kKqNiOOK2iw+N4BVgGA0QfcznkWhvqagHn
mk143MyysCs6S0cHBnxOwnBxqPqEOMMw6kvBLp/zFPUAtFe+42xjKB9tWSV67WASRvLKo/aY0pyC
q4IvQYFMmsekCNZQUu2hIV8QJX4tC4I90k8LEosE6IkMnpkSNvCwYFPAIfKX+gOnwBmaTzUeWJD9
h5QbtMZlR8K3kS+j62CetV2V223Cp9Gj5Z3LZnPssFPEh/xok7UIfj1TEaILF9/T2JdBCBDkwIg8
8wqALEeLDH3ZKguzoDgWGF5nniBPovz2uvbExqgGGk4wz7GLuwzE6JyFyG8NCqa5U7qbs5dnnI2N
d0qXQkIk6WNBna2XeJMHhy+nOW/0cgbCnJ6bdk/NWQy8eDJ1gDvA5cgPVID5J1rAy+SedVUEmwYG
mawwGuW8rs35UlecSAeYZEmujh6OSror5kHoHsMZgb3QImjbpdpCPj3I2xJogSjEd4bH6+1R0gS8
2Qs6EG6COJCNFYQ66n6aEpPjC7qqsw3gjx61w7gSmUE0R3aazqusYtmvRsag3WfUBOwfsCnwa+jL
0oCG6fy4qaPDV+2Fsy5JZxL2RvXTZaOqca/A3VwQgJgbUGibipWDBB5g/CkEadGGETebE6YzdQ7j
Ei1IZSK+ms6DPfbwU1GR0RHYbIvm4E+O+umRpVfSjO2OPe8jNNSdB60/7C0Gx1DB/EsoxE1P3HD5
95SOFCGTL6qIcBGySQT0mCRwS6NcTcIofB6JuBnuyKdIunfsZ96YDpTUnrlJEh/lkiE8TC3BPR9m
9P4hWrX8FB+w+7b2uuihI1EL4XmaHuzfAva9ZeKY27OLJ5nzEpgRjHAZdnsmqNnasA02y2Z2EBSz
CsoK53HYIlSDrJ5CSm/6IRUGvMe9nxQ5E9rwB11FxkKqWjHC7A6BeMH8XN0I46aBz6ojAMLIPoAc
dHORAnWuFq9pnrFVdB/7gDCAnWxhrEWdjKJToXHDC0z6CS3j42D/HAykdPO2J6TVoWyLFbnHHcnF
ByAfSLauVktymZ6gp+WzL+Nm5sNnCfxNCoQjv+3x60GUgppMmePTStpS1lRdvLuqbL76Z75HFzYp
fJJu2ogp1OT3sR9FmIHeohlkEnfjRcE31bgrXGH38jjSbhOb3l3ywdd1/JUkSF2OzjIZLA5aZ4zU
GyFVMelpZXsegdfP2WNNJVctNoTeJKLHfv6sLdPZFsLbkfZTD8KaWT9CztvthHe4aodYcxJd2kTL
mAlCjQB9b4OQ7VDOi72WJYc2dOnXG3h6P3KASFD9l9ByQaCOi/FDrTOKIE4e2roOBWDNFRSnx7xR
Aq++oOPOgz+avtFz57BezHHAD3+eClTNJVAeymL8N5C4ic4JaCN70MdccODxDdpz5Ucnq6f7toJN
Y/DrVvC5zwCEBV93ORNeLHXPtQiyIYmyvWjfBCHplREZvYN+0lJ4EjmVAiPAXSS6QYrwtTD1YkNG
6SNWuWDF/1Fa1Ate5tZpiLmCTPj6THC1sFJS3kJQrj1u2tlDoSEYdZDAL1CIfLbECKFuuDYE238G
6FiKocuaWBgBEObuve7Ahk71yHXkg1COYM4PWqNG22B2JoaYeuzUXgjpbS0uGPspJdo7VvH9UACt
xs7iJhbGeOFPVAWZdl8f4/ZLWOQK7FvLufL1sut302nlAKrZnCkE1CO5pV5gcjzfbnBKcOhotyJK
ZklLa10xIQDDnH+baiPmCTwAc1UcrkxIxd4KDbrpy1zzDZkMNP1VnKYL6D8oOCe4SKfE5qPJ/9nb
n3+MR7vnxMTamwlX+cM5allkCT6KVFhTNg1ukKdzZC7kVAeNSzcD+YE3kRW3flQTkmSusIJElRdp
hYWKdwraPG6H1clemjusihohwJ1Jpnvwx3R/he4pdCGJMqbx0y3ik061H2FbuJ7RsKo/4FyZiDd2
H+GEd7AJIosT49W2N0KPMWczHl1xM4/k6Q0xGxhqQewSLZeOHP6NKAlaMgebGVxo2KuoSoOxQr44
unjA/ig0NRYzdbIHqL1nLXBls3wEFfSZwvK8CRVo/xA3xRqG3ifzkdzwjC4DKZ80kL3uzBzjeML1
5tKvs5QkjnxkYDTF/oRF1LXkVfjwhPoBIxdh3GkC2DiwiRTbJieOeXoc6kcgZOVGuBu7lXyJJV3C
e4PwCzxkbAPRvZGQzBSnngZ0PaHgv6TtMIBb1m5DRqsTh88EM+bpqkAGU8hJYDJCDk67+J+R3omE
kHINcelwoL0YkLVydHBuhZrA2wBbmhR1UwKnO6b/Du3nV+FDmxfEksz5kVONxmnCziUWzNHqZpHX
718TxHaQ/NY4/wxmshtZmGS5Uw1XgFMgLNUCDMGxhfxIdXwDlrNCwoKPq+QAChyIXlSxp1CWkDAA
xPyK9+9UGVnz/IM/51nkcset8b6l/3sRiLyjU+wzwHOJJ+OzFzHk8XEHbc4lG2f8BxKy+FF77hhM
Ul/VRBoZO/C0PNcUhkX+F4VtsGG2BFYCxbI0xYhXBowgLqU/Gvd/kcaoD0nCUB6kcGKPi1iEhzxv
YQ8C3/VVZan84V39AnHr/H46ZtUuVgZ+6QJgjFA0DSS4iqw800FxvtckbiIGMXigMb7AGLqdRWnG
XYFyR+GvzY7fGC0mhXJJJvrx1/frXegCaNZoIh/YnK3EYGd6aMvuZldIXooiqsXiluNxsX2Vztwv
pazw9SPyYt68qQB9aiarfOyD2HUoC2xf16j6BmwZZfa8q5Xheiq64cQqe2JTW1TzjPA+h07rVP5G
Oxdr6lfb/lY8gctdYxXleIcIpafUKboFLJTZJIYWG1S4NTzoJ0YUzyFl2gOYtiRFVPxjpWjhS3Sh
0JOi7ba23nsIEKe/wIWOKUEF/Ec2GSIFaAD1NeCMXwfwD+Nc3toGraFSlqb8piRhYQUR7mukgCJC
cOcocFoQSOCm40kBR5m+e9aj41zpcMelv9Ysp+kb4Jj5Ys8oDaHBK++L+C4tnEPraRJjY9Y7iIfv
wTtMjYfkY8KqMuyKS9PtPzk7qXEV2dbDciE4+KpvUZPWkrKgmqmpbBaBEF11edH/9FehrsDj02PJ
lJA9lQuAELZBXdCXLcWZhzzHONhSx9jsMuAOJn7X47pbWghbVEAI6nm/7q0CHqbfpl24prISGCR+
oP15pe8WSs/KtTCXYsmfUaTEXrrnbaQJv9v/X5tQOLjrmkGfhp5flMVPyNu50dj1QGgMkq956bZ5
4m/D00sRvEu44lMx3lUx32DEINScpALVCSxrAo6mzfbGMAkuzpDrxqXmy/Z2xQAJMdYO6NBuRDYH
kza72CY+PFBKzgZhIAjs+L9bycKLNebq1CtxiD7AuOa+oR63tN/XZYwsfMm0dv7MAkAOzCtiodNo
pH6W+WXzjUaLoRXYBbFfwDP0wuiXn5T1yH3gssg8sI+/InQcCK5cUKVflb2R5kiW8+ZdaWlvxGyN
pDNunTnGDSRqTSdbvQXKPo96yrviNsHlWHbSeJDOvGdhfqvUTxc+wmCZqShUdm17WsTXYB6gkZmA
Z5IJjj7z+jZ66RMXYftQhXWIBLv0usA+o2++3wMhREPEhNmBNoZvF+hOufHHxHyxTnfvPH0DgS4+
CGdukkHMBAWQvCnwsGTZX5pXTKQ34yrAGjv9HlkjmWBBq9h6D0PseLvYlI+9A2Ie4g5Tq9qKs8jG
vEj2YEo1Q2r3Wk/fi2E+nqAdHlnL4QsgXaA5L6/3KbxIzlbB3eoNdZGJrfrIlC8DAK3AcfckewPc
8XCFfOrtFY3VrQ7nm4x3QiRfjR9BmF8H5MmimMtT4gIRjcc1Oz2ilnbcF0U1kvFw/X+VshIAN4/l
LBiFMmXwJiuEOJTmmsID/8mO1StdQw+0ZaBcPBo0IiSJRKdjAWWw51MAbNqPFt9oOGMpOuaKzCYb
qxwLl/EExqU3QtfErfu8y85kJDI7hkNc1iuuMM564K/k7Nkn1fHp4Ztd9yRMr8wl6j863LdjwU3L
oZW6hxmP/LrBCn4Alw2swFQBUrQsq0qZspS/6bLtPaHdsKFNYGYgU3cImuLJG3Xm23yVMYRhkGkb
+Jdc4i+DYCETOb4eMsGohvWLn066V6jM25HE5QcA4FXS6VnAgO30tsiRuXtm9dkB9Mj0NOftS7xW
cb2i86yuZ8Jgnriz1FFreVIGPamcCdphLGZjr7MHgrviEYMMit1s9j1eFHphHwO7k+u0O0SNOUYh
FWCSSnVzjaejYqvG0Uk6Ttr8gVxEj5u+sffPGWmQuy82wZqASo/S+yT50AcRzjkV3+IewhkBgE9/
pbtxJNlGcM4yf7Tgu/xuj2O+aeGLLlAKIizj6ccrBYgQAeVmioJZcAwn4govCiNGVTOz6twqBaTa
KBT1y/VV2vLonOdj2FwHDWZpmmDKJE2GHyFrjCbnxoaL559ZoTxVnOPYzqgbFgKfztter7MNozeB
vMes2yatOtohhxqTlRbYU7SQkFJzRvMgVLIg0cshzLbsN6zF4KQfuyw5Uak5hXJnLruibjJfKLt+
hRbSFQWb845FQd8xCfaOgp3kETZbu2yZBcCEEpE1Jw8eP/K2c0orS7TaMhdkVNYB1dxR/HiYXMmx
npAP+y3SNGds/APaEWkLynrK5tdJi+aUyxNe9hUZHBNGuwAXvFODyJRoK55KJ9Pn1TL7kH/5uge9
KKfeWeLw+rZxJd90c51FOBSDDcU7oT/YhxUjPTl++eonOOXRmj322weaWDCo0q8EJbuOq3R8G3hL
VjQroWhXa0Nx0sOeAiEG5a+yWAA7jTPW91upOd3IvSKshWnZu7/xBk/mLuVlMhJejS/hoDhyEscZ
gw6lzBf3HBpCId+eADcpq1Sq+Ch7nyt9h8ObraEpDqtcsULwTkwowhTxJFSKeMiLTok1d1iYTFwt
kCrbIjLV3ayPnB6V/HYr1m/xOpBW2f8zeei7sA1MihByQzhKTFqbSgPO/j1mn/VmGOfE64JwBXeN
xUzjB8Qzc1umbwJ2y7VyDaaA1CDDVy5m5v0sCoftRC0Eb9bmYyMVwc+HLmYzkd1YfAZn7mNKpEr4
xXvKV2XXUvnWRIcpfLnPpx66n88e8ki727E2Re3LQogGlPrWI2s2cAuoqcBn0ITGTNWDpAErC/Hi
JsjubvXqEsI95/V1PpgDy4ueW5VBoUJItr0CTdVqF6PxnHrupKFRf1e+KKH3ccyskjzqAL92xRNr
ze8eHZN0f8kC/+5+tG5/xDb2TMRmC99VgqaUJCeHQvXC04LezRfcqnxOKprX++bBjN01IV08b060
2ZlUh6B+4dri8nxxIIIajl+TcIN6DUb44LFLnkabBCheu0CIcH/s0ZK7+gRAhPIdp6ZKrLYRgb/a
2q0BBw9Ft/JM0Y1KOOouDhuP2v8P2IRlt6dwK6+W3Uba3EUAy7JNdDZxexWpZystHHJ39qqldqN0
qj52KtlcI31CVVUrnRuqoysTEM1kQ3ekg8hK9Xzm9mU9wIQrk4qOaQxmMYwK1Qpp9FJVOVtiUvAV
/lbtRh7hx3rWAuwac7j4pdqe8CFY4KuAOX4UaaNGo+4tHrz4aao7pFykk4n43r+NZL8q/11j3lmI
UE2a6B6VaGXv1R00E5YDEA2FyG2mJlL0iNNqBGsAJEFmH3MsPtOnQjGGYuJQQ6XCafA46xC+SrRE
BozM6vWV4D50QQu590uOUBf6Ah7sxc7Sb34cod+TvX8a88zb5oxRBfLtgrGCOIoRQMhdfaZX7dqb
jvua5oi+v1xzUMvyQnXJ+hPGctr57twR2l1i/n4uvB3ta+anCxmVnrAlbve1u1kbdP4STfoA66B/
ST1OWFUOV2JaujWp88HAICbUXRDlElooN9R13uB+ZzUWOK0Hm9SDg1dGCoek9mtWI6HqebaHZtPf
nbRclkcBnzBpl+wfMerWGVHQRfMgCc+Id5aDpHaNlbkErTu0jJFC1ndfOBQQ4os7iR4qf6dhAQUx
CjVgLC3y4/ZefjzWpPxZc92w+NnecdizhwyerfC5Bl1UF1Pu/zZWXj1VXG1/m5DBbo/pg41B5elg
M4t4G7Z5QEyONZVsne8CDaBLc8kP6p0yNu9L/I0GBZwaVkH0/4HCu+/q+/IJ1dnesj93JSQmwuhq
rkXgcUjevjU/ur6H7GkkNU857nBg1NysllKS5OtXm2S/5O5keuWrhTG+EP3ByCwc7BajQUjMwooy
rIOM20uu5gu6jyXAZz/Bk10CPC7oFJKcMya9TqYJi/jfAWGnqZLFoQhYi0oUOMPryqJxXV3HDDVV
d/Ej0gmB6oKFQh3V0xtXPMtgvo9rn96FprDlo9evJkwN0nLP6q4hP2JrCqRLxMxSKnTW7NvmR3hq
7yQyP9zPPBz5T//Ho8FKY5yVvFmbmKwPpi6NceSc0h/XXFbODkaiNfq7P4TJqidWr6mK/dvey/nA
3bjQgg5NksyBYgAG0NqwpCQetfLwYy39VIJI03Wc96M2lZjhOB9cv9iJfK8TguRmebOktmOvL6kr
/4sc3nnNHMMAda+JANLl4anWEVU2u9c9arLCmoUKTenn301S9talpNt8eS2ZjnEjxjEqrOjvhuBX
19/kgjYw2ndfs+maFFAsiOtSQY/ZugjU+5q49zBQfqcOnQHQWYZ7ZFXz3aUNRVZj1pXeBz8vZdum
SeA99vMJNSA96G5p+WzDnY5QYRH2sbe2uO7rcmKSd6EUaJUGbQw+qOqutxa53003O86Xr2UytvBl
8kGq7ubh9AgjRhB/Pkcn8HcJ1arMzBkl0lhQwfMiElJA3wEuIg3Qx27hb7eiP7b6kI7T0AaHn3ZP
6tIFBZBN8uGUGK058i1hs6aejBgQcxpARFTm/M1h4V7CCrUGbftnUJ7BLQW3gilE+iEInlKwc8Y7
XYxf7O1eAlBoXdpjo5qmQZRjf77r8/Ps+SxsLpxRd5u5lbH9y3sfZVCDaoxOhJstJrH56CTYm/vU
zQFEozGbqN9u1IscMRNsLlFarM8DE12y7xJ5zXU9OM2nNAxg1ZdYl/7nlaBWnVcL44kVN/VUHsdG
eU5mqct9caZzEhVibCD+RDTEOkckSFwR5yqMq91ieOZhsEM+4gIxxGB0gT8rR3M073m3Xwcknmrc
gGDDSzflC0Y02xd8PpbSI/E+hfvJJWOLIWodVcdWsK15tgdKvUjGcAM87CoplJ7M0kaz8596n4MX
kZd7sZtZNW1n03DNqN//e03Wdyb7hn9NY59LEdzkAcqxQf+o6gDrVb5vRYH+Q6xPOR6xhmFwYYBh
zkcbsI87P+zpCvXsdYICAHTsXtD08YzvVFVQULAdnVttK0Hh/0utrh0PJ/4tFk/ysu9mnKmtSxSm
fA3GuDwBOk8f8et7NkOIodtUfm2am9kpjGJF7YQKZpfnU4utsgSTqfQyd0ssPC32GaCnP80otTrj
pjPFexl2xi87UbI/LDVtQeHHLV2HS/JA9OnjuqxyPGTZVNNATNw1T3VQqT8RCN+IGXSH+tU/mjnY
Yji/5wx0XbGA/2Hi1jI4gqC6qFieycqCl1m+rpddwAXszMZN1I7fKwqxnsQaTryV5k/j9VJeGRQC
yUw5ZYN8F/JoYgnuvRJJHkchQK7fAlncgIQYqYj5iU8M8Azmf5MtzRe8gGcXZI2COh2GL0X32yXs
J2ugJGss2Fvegf31IvweEG0ki1ifu8qC2cPT6sud1LlHt7UsCp+mmm01wcGsWWgddSguHZGJv94M
JErvyu8Tzs7AIT59Buh1NeCHlMR7IpuvDErZ8osZC4KW1ODAxFWVmXZke1rIOQl9onxoBbzzkO1P
W5YuqdKWIl+sldAK3JpcLne8N7zNwltefyIEC3TCF6KGHkI0BGHCutXAOXBUC2CTPUkDehhMdlPd
4m4KI85sbEFZhSWsPdqnITHQYOOF9mTEinfg/Po9MskcrNADPeyktWD3X+fTLs5rVQ9N6xGUuQan
Zo9VOclHEkmyuqIreavA29cRw0I1H6EwP2N8IG0ITx8ehikg0KvStLTdkQEGtNKuJfEDrL+zlMUG
ibz3Mry4OMHrxU1D40O1aIVrVLDPptF56DYF9SNNPJ2Jrfh6SH76AWq/mbrYpUm4B/oGDyLPeGpr
jgYzoEvImr62ZY3x7joXCjVDRJhRLwthmprTa0g/cs9MDz/kA6FJkQhnU40GcmVgLCSRcQd9citl
0oe7qG5SA9CkRSi7pVMpD4Pv7Wht30dD3ZXISSjvsSr4VYt1DF6lLDJxXEeOGP1l6LEN3hFrqFmh
HhEFjt/edPrR9vZQ85FsYHNsjqX7Xs5d4IXfKbUr9ASUGJ8B43hlmndbRYNV3L+vzEoouPRPcYMQ
DAXMm02k4s8jSuJ6wRha/1u6zqSgDwuBiE6HGvciXuUhSl7JJc6U+GghauaDsTTyH6Kq/0TJy0Pn
n3vJGSJ+ZQ4x+tIp12YfrcDQmMa7SSCsngQ+xlyjjOTsl1WCHXRDzvgzGs5ys0epSQgRBMFNhRqf
xTtOpvoIWlycp+f8IP7bhrWMP5mMtkkcPLbrT7IYAPfNS61DJU6I8SYAn9npQaIoYyC4NE+ZEsgq
WI+G1UxNoonBNaLbvZY3H8fVYpQ5GR1NOwdmN89e8ZCaLxWoHyRtywh7s5eMKdNOivP9HK7fqfNO
Ci8YoKkolcc39qM+u8QpzFZHWSFnQdfQGIXN7idjBq/x9j+eRPvMBcCPPeMAta/Mx04OQ/f9SAGK
EtbN/V0gLaIkWfNZ+W93vb1wLuVOXkN47a8pAJai1tL9s6NcGJQEErTk/InoyyMIVp0wlwaiQNp3
nYz64W4QzPY7SCVQr6NbcpuTcicAwfMFW5JatqL/ZWGhar5oaZofwD+41QiTLpo2tEKMfVUCWeAf
XyQ6U4CqzWmjVkNJF6yLaRh5BGn7btUI7+xLxwVNkv0BVjuvgTKocvkVyWj4EAHNDamzG9ZFQ/m2
lLeoEvi4kFVhFJMLSvuTbc71F/Msvl2t2pLY1nz19k9t64by3YQoVGw+oPuZl5GICjf4MPhGHe+0
sXFefMUyqX+0i5S0WsXpWargLlXQzb3ruvvicgmHD2jnOfjK5de/cUgXMAHvoc7ya9Np3GQM1Ec7
Pv5mWw941idvyIfnra8rH2kHy95+qqSAdQ24nsxPFwjUyCob7lGa4jjF+KtGRQGWOWsJX/H6yz87
BLgQmN3Nc9bdC5MNGwHTe5J2q5y/O13Ea/ZXD9K2Sr8HIM0w/LAbmt7GfuTtK3U2PzCzTR8FFVEJ
R/p9g6Kd7/OyfBBcecF3KZqkFL6c3p3rG+K4FqdmBJc7nbtDnnYy6ONU+IcgQ07SqqG3ZD5kJkuL
roXeIDBrXcO6QdtPf5w+QKFEEoip/8m0CqEUidfMYDKcOyjz3pV234QLivFc8s3BAm3yrWoctf/d
Xi6NqHccm/79TiYTLhGcKqk+cE6so4UI5QdtnnfLB4Xmetaj54gEUPnTPpObZVUQ9MapZLVQzXXB
/4diau1QqViFjTOKaZALcH7lZCHWfLhklCQ1zsGfb2Gmj4xp/vf5bWZs0CSIz80oEO1tS4VBykHD
EWzN1zKmT3CGwzz+DXohs0OvtRf2rm3IDQoljJhGQqK42qcmw2Tn40IeTv9RMTfhnmjJgZ6PYaLQ
EEPlAlKN+FHDxq9V9hBn/V+oB7jY4QFzR+YRbzsqFcrfGtfogMStOV3Z1kRGZIsvBK162w392sHg
FLatOWEyXp/HKdrENTkHErGn0W5IJxe+WGWTK3LF32KTBioTrw2ETk/ctqTRORqDxH5uYfYNu3m0
gpUw6mMJ2V1k/5qAwoYA3zmweW/qdsN4sv6AKMaCBIvDLg+Tit+SCWfVwVWmPim9bAwQRhKg1frz
iEGKXrQFyUCWXaPIDsv4lhB/saV2376w/Srtf71VEZvhHtVLTNIP5bsS/JmUFGJ/mSoo/BByuBBo
WiihLVY+JetLOjulbKRZo6t/d5Xack9GABc0HQoq/bmt5g1z02fBfFkMdwfQT2IB8ZjuoIas4KSg
e3quoQCwGUpWx74kmQCWXvZYd8sW6TDG4WCyLn3ku1CsoaLSTexd9GLfNUTEwL/NF6kVtALqZx78
YbJoXB1fI6nT7JhutnIfhHIhWwPKu8vCjOCt003FGxastSFyr8QDN2Wh3wKTOUh/R9ieceR3WjXG
qakpAJvTiMcC11zGXTs3E4yQkIQU+bYbRVryqlpEdSgsZNEJmwfLgZiEw7Y1OngXexxRX7GI8o2W
O+cPQLUpxx4dpMxoixhZbOyd+3d8f8sEHklEbPHdKHPp9hjbj66y4788QnADFvSSvFVgfC+O0oRC
WGwdui4siPJqCaBYs+oFmn2KM2L+EBLMrxKuD0FmtRTPRJftH2ChY08car0upcUfY19JNQB+8ORn
zIwV87rTJB0beEEfV/ZwjCTMt9jmZc6zylS+i+495mY700O9+dSD0M+Scea6rsPIN6dxc9CySpnx
mFj1SA89FakngdT3TBuHSlYe4RK37rjOv7ftgc8OuIOASKD/W4aMi4WF30SHufo3/mPtDFTWMJjE
8asXcvb8cKzL4IjEjgDctVOu+uMxJgww3OCGT2gVbLRIzzvp+eenPaui44jdudl4U+EpXUiLMr0F
8popEM6hoijXZM7p4xGc+cVp1+UscDqR2upMAY45WvM6o0IMWhxxwYVez3X7+SiirS+O2+wI0fuh
rWaNUXUzM/NAsMShdpFGPvtxq9i5whwhiHGYpQfPXtEusfY3ODjvyFkGSf/mGswoDepcMN30nZlZ
5BoLovg23UA9GPl+Sa2lruay0CwXTFUtPQZVSbykfc2fad8N/7pCpvu6euGgMQj1g5o+Ni2djovy
dwfxWQz4+bgZgr2gvC8JsjW7jkxlFGAs+woUsdD9p+iYPAOqcckq22Gn7vA/Lcz/gJQSB2f5Q7Tz
hjzW8hV9baluhQwrkVLWSLnlz8U9YiRxaIl+klC0IN/XuLMSWzr1oU48Eb6DTnKEA7hMbMJkx6e0
XvhrVsBM0v4pDDe2LxB1Wh97lWto+h+7I7XaFl7XJS/uGnJa2cdNF0Ui1m7l7e3oNsxykwGWJ73K
UAy6SADyq2ZPJjiKNu7tONunaZvUwIergNVbCdHiGsr35RtzBivYKcJyJYa2cFOcbfd9N8CkXh/h
IPX91O3FduoaKb8wLCwXlEihNbQeLjtU
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qOJ+kKfsp3jrMDNmMskaJy7e6tpzEca5maxgRWeJQUvlW5BC6ePs9U2JZ/s3t9RdSvLLg3bgriaz
ZhXFzHwOonJV7cIoNhroTKvErNf2+E7MaErfoBK8KXX5C5I8ud8tONVD2lveddYFSTKv4giaRfr9
Sj4uUi8k9dYmOMILE64WtKizQ68Oyxd/sak5wB1gui10hjt9tYjUvizUzsQ5pU1/BYMvdtNkhXVJ
k1pr5LfBGxTAicOV+98QgwBHUQ3q1V4bP+K8yCHMZlcyByE1hlMuGNseD7cceamJN1SjxWyEa3Rj
akg9I+Om0Wyyf4F3kqJ47KmAQ+HXxQY2z3ZV3g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
huIH/kWEMR+RWFFLlde55g4qsqPIz9Dtak7Dm8gEvQq0zltifuOSsQtcaCaHq0qraL9n+thpJ/bv
C8T8uiXB+OvgIJAY7aAWrfLVICr358tg+gUaikd6UfHkzl5t9LKEjXSWlBrxTfH0MImxE8PT+eS4
laCCtsLIKf7fJDCVb8yaixQCeL2J2ftu+m6nYxx9490hVI93uOtCF9Q5nTsUNPsC1K4k3UFosKRQ
7zB4GIXD5wzpoIM9wiCldL3W/zPgc4aIn1L5JOdUu9RFXzE662PuaMnCo2g3N3KtKdKFOgcCiPYF
bZVSEw14cjzHgPpmEVpQqplZWxdhnA71N/naeibZUmF6cOmdCN11Yu9m54e8/YEt/dn+0VLiliMd
N95FLLiD7nDfTI87ZauHj0fF0/yL/VuguZGXzuQsu4FiZdmyi+16EOZuxejrem35Hc70cUJycNqT
WbSoJu8bASQmNgPgaNFVq0ehF2ofThE0s6blOAxcoJazjghgrnMkg+m9ojCARtiJ4Yka2KuG1Y85
S3BdVHpmN0eP1pVBmiUpmrsej7lV+sn56W/0pNZZTGZBALdYqmOGnApnaIrVjaV3J2de2kxewWJC
kJJ+SMMUFJaFDn91IQfBzep2EzN2bMOkWpgFdJpcH6MVcVF7wLc7ZYKy+0lbs3nwIhfna0k5CChP
l7bKnEydm2pSaLQ3NeV8AwH2KRUPhjXJ3KZ915XP0DziNbemUf0bkdPSb1U3q9DDhKsx1nFGGppE
9kLxqE1Zz4WoNjE5cNWAkUf45SMvB7M22ptfpnXC6IojFsir7viCJrKmH41iRHKS5ifr/Ksetg/S
wch00bN22t1St75mBjHI4jbK+LFn2vDusImWCpao5mRlMwNr7oMJvjGTuBrm5FBuqMvTFnXx4nph
fNlHY3jhmdoZXeE034j/IzY62BDuLCGXeCTVZamrLtkFPsD/QqIpFZi8NPP45FTSNA7hPvLwuRR0
6g6Q/EScupIJRhVZtnm97kIuQca8i2g/AFSA2UxiEQTdBIjQ2CF+j0MkK36zoSRxS9OrRarmqE5P
5fiZYkjq4Jn5R3kFUNUm+IW27WsT+yi9lNEVb0Ckoo5v9ElHxX6X0YgDUHQGxwrvWqXjWfZxY3mX
lgNqU/TGQDO/h6QbdNfZPmjw6BVgpuOXX6eMT+N6tyNVWes+9B9sCwxnjDpGzP19mFMQESe46VKO
w+jPhxLzCwJuXQFk8f/Ie+3lxfl1aiT27gk6TUac2lhvhTQbIWil0scslshuxwj2H6KiYKsXzYrG
9DPmNDg76H0GuEUeoHSom76EwTgAqVEhgCKZjXUckA2k17YZd7Lx2q3JZqsKDGYwPNxtJqkQyvAc
/4bFjlJJu/r9b5rNDn3MhgwGNKUdZRfsN/UsseT2JWW3tyZEgMT1Od8Q36Tmw7I0w4Z7lvJeQIz6
mplYkK371FqQIDajsKngStVScybiHMkVaVmor0UFXhI3JJ6cN8bVf52LhnUInbkK3ifX12fuYn1N
MhrUhbfUAXKhxltKNwkStC96HIOV6pUuYXsRyx/O4YcczyF9oawF9zm9BhHUMI/COFgmGsS8BXJ3
zGlzitKJ/k4FeEi7VVSVX4EyQ93C8HV9iuRbJVlxGWqXum9VbIExfMPx8wOYTP8ZlSLeMqJnjzNa
+KuN7sWgjBAUW5866qAmrKPPucJy95GNff64Da8wL/d2sqJgSGkqIEgw+eliFAudNCXa6BuQUR3c
qBIM2jMZIkaHRPLYbpB6EmjeqS5l2VHZtkHJV1boR6DJIoU8iV7zFjnmNWqbpiM7BoWCmmZzJHIo
RHGOKFn7QNkmUx5yAZ8EPFJjMQoUOMSaMd7F2rMkwT6KiTDVP75qDJ4468S3DuCEmdN++KbGBCBp
W1m5z9oK8vT9Uz+3w2DU+SIpfPKlFWQi7CjJkFDQbfNsUrHTSWsgylY8Zj8i0pE5nIMZAQs4DvXW
saEB62Nu35Z29t+wuUj0x+mugA29A0IlrxXvQ65aE+1JpdHRXRamEtyJlGcEArh56VLmf7SXiLJv
u05+k/JCrJTz5v0kHtCxq0rVrZjJodvrEuGLVl/9GdF8oko03vMZ2LkDlJpo79BbuiJaENILxkUu
awhc94VbDC890/tnLYBt/sErE5CCedAZzpwsLw2f1Q5gA/j3nMsmZlI+lxkd7mCMOjIlxczXcdGT
KGY0rVg7RpX9KR+G2UefnEeNqzHS3/yVEYhD53x6ykkqSeVrMsXs44x1Uyn2qDfvDClIE3Cyz259
vf+a8oVqhXGY7V67cufAA7e7MjVVjdNF4Jhyqzs82Tzy0FJc1ZHdbJ53D/HONgwP7PAbwn7lkJaF
tHZKjzsLvBVXPTUQHu8cEYlZYm08oUVeOk+qtR/nqYmIK/ShBDF+Hy4mv0KUmRvphF+Ja8jxc5xb
KkVdGmSTZIxiCG8XlApD62fxIcIlnjETsUPQKo6LzDPnKp59nLxBVqEmUNM0vFimcQE5I7ZBfx4t
Ic8J+JgFjx5c0YNrabl7NrWMG7kRpuDr+DDNcUBHKbaCM+ZULQ3BgSVAPtqO7TMFYnvOr+F7zHyF
wHUJoiNZgYv57ZS+cfOAfenezkIBJBN1afqQnYLgjpZOwlEWWc5tiw9+H6Iblu2Z+Lt4lrtMDtC4
t+iR7DNoY7K2vodLD8MbCFVEFZ3rse7Ctp97zaWlRtHLB51UBLH+XXdOAZ+0Vg9hhLDEO71/b8PD
Y2LgBX9VQyIloSu+Yhh/VEgKjvYUNt/uHDzY1bE6Hfyz9OE2qM9fvE8SWjpFVGvPWF6aGb0mw8Hd
r+jOfPoNbA6AzmUj3njoNzuB5LK3+Y0R5FxP24KDD/Hd8ltXOZCrdctMnuLPpTYHuI536mEeSPRz
bVJiuIjuvaM0qxsgzmWzvR1hYBKVxw4i8FCKSluuIRU3Zt7YfDfU+4QWDOG+jHzXcwKpIY14QtJQ
q7waK3sA//Evn4npB4q1bcMSN9Fvmixzav8sJZdtz5RoyecmKRmQOtMa1MJIxpVI15jd5iqxyOOM
MiZtDHEjGzWdOgVq6rJ6qdqgK9WNuInUaX68cwl9LAipbSjb3OgdxQ/5cnybl2FYuID+4zUJJV0P
9xPSiDqvKBScdwHsXVijlHZ+UD9WKj5r1JZ7Cz4mnnNPfJfMBZwywz/vtqH4MylousiPI9asHErd
a6yr2oM4yGbUonSUcv5ujr0pAmPCyUASFwmXXqXKekK/JlU5gjdP9JOi13JqHfKhrRRG0hspbagG
N5P+hR5Tc1m+TT9LGBdkmvzpKM+bGfHTmqEZO029A6E9KOdTL6ftCYypn4RKmYYdD6G7YcbxmPo/
yH3LfqPnVEGxlo8sBG03cdgxxax7Nw75/b6xa3G9Y4GVeZE7hVtE/oaORlRHmDxY+do0s5qawTN7
3x84KoEqgCiYOmQHctIJ2QpTURSeiDgeLKwT+8dqEtoZvSlI32feg32CKEFGrrmvW1MOcdTCHe37
uA43WWt8jQY3y1exjiPPBHU/o/1a+bQ4sJ4bPYjhRhDOMINUnmKjJPWqDNLK8A59w8BinYNSrnQW
mLzOljbTmVk/qWanrAeykPiaAcvpYD+eu2547vQIwh8QR3e9M+FgRFILwNx0zlVJ4Job0K+ofGto
M8gaLS5alxEYe+gTS4qdNPxla5faIgIZvzWy3+2fHUZu/k4xn9puRDndfT1zjKtntSAoKDBsXfYD
NM8u2UrGvF36jIm0Wkwu6Fpn5KpBAZrjaNEDrWxcqqxK/hj+dV8mAfLGwyIe3WI3NZZvef5graNZ
FFCbJ95+MqyXtkps2mfdOXntw+ruDYr/yI8BSwK0y7i0QwMm/lhTRJLLfF5OmXpuTGt5PKAfq88v
ldjnyk4PUsVynmHwQvs8EV07BtLol6JlmLK+0FIh77F+/HyLvXw7xZoF1aM2/MYoPVuEwP8cE8QL
X1rxU6Ouu4+p3lYBc/e0CwcjXT2Cm+iA6KBNHv2KxZVguZMpLdAG1NTTMtlxpGgRfnYRAv6JU5T9
+LhJS4Q7pOsETJ1gx1Q5I1OiJNSgKadEOQnCmROWfOY9OOWJKapcBhQBqEHfJaeSX40sGZL0uk/s
4eXgR7V4GruDS9Pczu7gSVcUfVNwRnVX/HaRjK8ewskP3VXRdzJh2EaBDE2D6yGQ0JKnO91+dMI+
RVPl5o2GfXjYHvLAMDnK7nZXEnF3BAPI3/NZzPWmqSns8h/jw+9S9Aapvhu5nxGFNmunue3bmzVY
OAOS7DVL+vy05sR0ZcbkMcq0nhkumg2uzh4NfG1SwSXy9VDGjVNgq1hiQP0PU8/CnLv0XrCiDMyn
aio1CwlCvSFBdRkqNWw9VKsoOY+n71isUihWYtZIrnvb2/UhS+75cQrITWCeDygH79r0U8FouFDT
h8HDwOVuW/hiXdbd8j1DNsBySgHU2uz3S7anGF5ItI6WRZugwSoxJ0IsqqZGa1b97fFuAUGofVOV
NaPbKr6HFYmAB6G2wMg4xEl1bC7UiDbYLpB3QDvaYXdKyQKaFrRhurgV7P4h08v6dJ2GoVwFnWl5
L0/z2CZA3hoGU3H60vXQz5wJV9gYDx4hjbZN94fNtLMx9E944jdoto4nJnvsrutvqsMNxJHD+b0W
hWAouEMrJCUdKoG56b1ZxYY6Xj/yzzTZN1yMM/mGLIOUeVEzgBugrOI2XDo22kSV9NgYlmaXJnOW
lsGdI/YYN1nm+3sGJr8cddHVj2N1DR/BcqdvscIUTDWedfJ7CdoLlCLuQ2Ha9OvlsqbUgndSTgWi
UEHRAbmd1hVcf9oKqEjH4VGHlWK60HwjZOK5lcPza3QScGHHolxriGKURNHyMvNO3X9PrJwtD5e8
MUogSc827Uphr1NiKr8HZBO0xEsh2jI6LjO3pgkRyMbHg1TCij88SCBtayB3xCixScZEiLUED7Iu
OigLHn30oRyZcWQKZpjtEI1S9i2qIj1PHYDMZS/Fx2gLoZ/kEK2+PVHCmAX8mmNwsRhufWlROsXt
9RaW9hCl+Zt1twVz1Ecv5UBz23MhGhsaPSmbRkeoqRjEEkZlQMrCeqg2v1Or7WxT1It0au0AwV6b
6OALgybXgXEMaBkym5KcAlBN4HD4RXYs90aIKrnsJkcSgpLk9x3Pq0TTfvOz9zYzvAZRD8pRQrat
1SmUpreR+CMlr/dhNZobXPaQF23p47/ByfwvSXOSOR5yihQUBR7u736VrpQEGC9dBri6hKpa3VxV
2xFPbs748Wk1MOidtPdMQOcPOD+pyJmkrcgrDeH+mUdkJFIaq9moTAUubFlmIUTDO4qzXiPJbxse
29jIkO0j/uzf76TAA2nNB9bAZfqfgoST87a0POJkLQPp13emkMdNaNLTGTPt7AdoCXzJZLekalGO
5Ajr2eeZf1ISzOp3FcLb4BsOJuUy5fli1aIWDeXypL3W4i426wX0DAZuxsnqUCZNSGMV/BET5vs3
PFz34KLKoM5CPywMCrFUOrUJWs7XMDKQaMGpt2KcxCqhW/S55mfmTQ43NuNRCnyWXJsDRekOsYfu
Ydr5Bgk7rM+GE2S8W6HHff7vo57Fl5Og4V71yx5VJprdHzVOYTsVPXhxqSgTTSLPwg9eGCSWosv9
0eeDK4rJijGwsS8TXlO3jzWRXOP3TPLYbWXj7cPKv0mBKD7XNl4lPF2JCSZqDHvqY4TXSJqAGAdP
tw8HnVIrv7zu4n77Q+EaxrrpE+DpKTv18t4Ggx6WyhLZghAc+RkRIB7v1iOFxjwpikdEywSuG4TN
yWVODjVA3e+pUs/4IptSeM81n4P6LWyql6/L9K+tyaIytfmffZ8yL4PiiE6rEuqSg856Pt0yN+bd
esQgKhuv70xQexjNxGeeWQOSIWx15fhFrPJWFWEdTWk8vJaer35aZxcwMHt7MwnDQzn0A4EAjMzb
N+uvH0/ZsgCszaDjwW7elyUaxXVV21JxH2k06aR/3Pv862jGnjd49kLR/a7kBTcbIyqfkT2481uq
iFDsTfMCB4UmvyZIDIAIQ4on8YTYoZ3CiZMVCLWmmhU9SMt58s7a/g3sWdD8sQM/6FRs0SqSfzq7
fpOhGzPENW/7MRXwzUpF3MsdY4P7kNR2MbqoVV/c8Kbvent1YsrnFIg35wfwuXZOA0l9t9S/yAZb
40O2SlJmYAFoQHgxvAPmOU/+EvqLe1p50i25YWoTs5YFNSr2MvXcxZ3qJL90VSAxrryRA7e6XG8y
c9gVqAWxztB9FDZSirk0xFO/ue6EuLWqr1oirivexpjhvCJk0E7s8UsERZ4FLmHq3JLgu+/mt9Fo
li5Au2OgA9jhb01rW+CvHrkpy9eqgLWc5BiD6vWNXJvwMduZH8fmp0snLi7mVahOB2/nv36e/fo4
58Huos2jzOilrflCjeFaapA7f4881/2D1ZR3ubHKuCzMNtdw/3OLOFwyViqMr+GJp51IbtBB0LAA
Cpm9/XtvRqUwp+6C0yd00TW4yZ3BM5wv8vFFVcI6Qv3g/tE31meKSpuw/pKdrnVvm5BvZQvApoiz
k2wuf1W1emkdSyqGEvHF8B2vJPQNMlNCN/uoDqWSsnp9T0LGE0Wqi9uBmJ9ksSVbzxVKParnKp52
SWM00Z6pXFJIE9Jn7X18JIXFaLGuAQiPHygO3oeWsLYsPT1xFPrzAti3rPOgd2mRQ/AL4f/mDbQG
YBu/JBk1wux/++4vigTR5cf5F8O7+3+Xin3ryY7zQoR4qHbNk88oT+TrUDVW7tvq5z3NO+3vbe07
JCI7Nz39AVH+GO1gS3CNOgICoEQBsiTuW8gPiA0RYycaTrtoprbux3cCvE228p5bYhkZd3Pzff46
ch5auL2e36zwO+72BJdfUbzVrwymkVcb8FGDiG7Z0a5sT+22pq5cFdGTqWM5KDWfc+gCJyawRRGl
Cv5zhNfPbsFap0OoE2KIB3TuXrKF07NrTdzRXgEhIvx/ndOVrNyz4z0Y0eXYujoyCdwJ9p8pfjY6
GU4Tu/mZt4+dz0O5QH4Q0BuT6Mxps0aRJR4UGee0x/2oJT3UW2TOztOZbhiPkmZopSBiHvvvzwEZ
wylmjREgFW7TtsunMLKNKzaoknJe8ra+Jwi1bDwY1VQTMeiEs4kGFVK87aTOKilVM5vYGJR+n0pO
SB0RDSi1Y6Yy1OOpSILKc4F9/obRzcBJzJHLYmcUjrxNqUVtHxz4Gu6JmknkUD46KdM/rIMZP1th
ijGp3WtlC97yuxaXoufxLcJNTUQTpMm/kon97e5897js+AeCIwv7iw8LKfA9XdwOwUY+WP3dTsUq
D0FNi4dd3Rgacrk9ID/8ttQBQ6mlb6+6k6lz/hHUsAvtzTyaPfHmNhwhgycp5IE6IigupNe6uenT
Rbi1sTehJiIBskXvxUWi6ssVVtPpvRtflFwO8/W2C5IVKqyf6EHGARhwhITxz/+vOnopdqt7bzhF
nx7KLOgY0YktGLn0bDt2utCfAfjUXOt4jV2+p0x59VSpjgzGqH/X6t1cV2FdZGsfIYefX7p4v0ZG
6IiyFTZrqSMdnq8nygxBh0T9NrTgCTu3cwg/KFbCq3o76LdT+q5jb7J/zNBsBAVydE0/1DRCCzBH
9Rv2GGukeCAFdnQIzRxfaphTdNn0zTGLxAYeuxOhStGTF3g2YUtckiqF2FEpBM/5si3WIjN/PCLA
KTnby9RuUkL9KvcA0WllOUyMreuyf1T3JEGgAjQXLtQhB8PyOUCAeHooOjNvDM9uuObBCx/DyS9Y
eVFVk6Fob1DeL4x7/euPICYGOQDMtUuDXPy/9lS13WwqffgcYKVFYcAlZKFGw0vUNfhAVC/8l1uj
byK8XrHIomSc9FM5QI1i7Tp3z4aJoPKMrsdLVdyexKDuv3Tql1zKc6BufPI5F6k6Da8GEYKRl4w8
SHAAs19icquSPaQvCTg9yMNyTe8wD4UpPWZ+UwMh5nJhK1VSmuX+HQmuiTXTAADyA6OSksymuG7W
8Oeny/hLA8XQ/Ao62JetzW303l8FfWQIdyRxLlSSUBdQ47H6fZWcR+9eW8qJovgYhOxFB0AXE2VQ
iyPGvv5U3PzTm4vyfkdrKgTfbiX839zdMOImaW0NFgOUog6wBeqro5jYKAuKy/YBQeuFjgsp2H6q
THiEz5+ovw/UahjFzrNcFKsMjReqUN+BNib8Q2A3DY3U2TXGuadYQpP5tVrN2zSBMGRE2ylx1pgf
Dtw/8g1szN801S7ZRV3aL34qjJCNy2RkxQ2cckcxL6UviBPNy/ceWte5ddUGh4Z+urHO5nYbuUBt
0TKbY3GF3FvYczEiaXhcTYqOELvoMD9gckusHCC2ByNlLBPeFcr6sXgdOGIsEOOJclhR03QEHil/
Oj/lRoElC2BK5FS9UM/IfEKTXbWVvjaIwBitE5r4rxgsFRIwjr+SXXIMHljyjwkOjuA6Br+RUKUA
BGXW181Z77UrbSIZn6AsOXOrkdTO+B4VEbNapQ4Tu9twB9lm2jtFYl2DFfru2/K22lYjn6Ba5Fd7
xpEFzu+PPQ9TG8YwyN+mgV3bo33p5CBGEUnW2MaT1tbxD7uoC8NiZg1eDByXH5+hi6aq1fgITVQG
2syn44XbQz8yvCvF59oP6jOPmM21afyFfeuvdyVyLMiSZYk5oDv7h3mOzQO4jTx/NhZ73WrJkEJ0
FxhySICH8GWZCvNkHguuvHSPyfvbfmisB/3tyNeQGTf9E80Vfj0Vaoyx9P3IYHjH2XOMOuIGK+Cg
zYnNcmPgErvuQkp9EQ4ZchazJjNlNMMOl2jGs/3Zo0QS9iCkedh31EW5zEZk768ergS8GOfrz7A8
VGUHT2wih2GUaayprf3urBrzaqUPkEACFTgcoRGUErLw8bsSg2tJ3sk4eCrn+zV8keQKui/3Q7T4
lYq8tU7YOslHel00RoAAAzfkcU1Iskc9RB5XJWJHOgAmAC3iH592WrSXTyt3zpxnfKR4IG8eG8wD
Je9kfCJYfZCBSTiirnRrUMl7UwDZscjv6znJFf60+q7kDB53JNKCeW5Jfu9Vtxd4G9XYLuh5v7OM
Oep/+OzB0MLcL3KxhgguFyk4j2Le8O0yJ6QGwIH/RPKLxGaVt5yGQw8NEaasSUU18GHC+qdmhlvT
vXIDYtXCfGS97F0yw/LGDFnmdGey8C4aT99XW0Jn///fyWsEit46R1DZoXojvif0pCf8qIEUHTAl
+yaN/3ip4S4LoA3ve3/DYFBwIzctbEai/60sBz/+oILD0O6p2qQWSNsp+l6vbNu8Oj+hmnrf/O+1
fAjssr6h3RA+lwVDvE70sUpLMUYMMa3H2Si1co1U44oXSPIsYfh0p3aC1s9N3NTtO0FOshEFE2JA
owGok8CxyZfQQRqzKS+M0wBipe4bGtHtLzaiiQYl8nqdWpPMZYDGrHyixxBkC//L7WScgcnG43nV
NHE8WW9oT+pL0hUW7cXRr/AgnSB5vzB+Quq8UNAiE5TUDhtkCWdexfxuuWEwQwuB6oDOOKhgogxu
emqMDV9S7/snXql/iAPtAq81VwyHfS/N8JOwCYValGZYVvaFDXu4Kuhi4EhBhLrOTo4nsv+9dgNl
E+d7ysyghG0TPCDJOPzL66O3moVVKN0q9yX7IURdI2KNqVsuxXUtmMgQ2lQdDVMxzRAZo4qn/ZLm
ospEdJ0jRybf99gfPgaBxOHO30jZY/5KNcCR71uH6ZuFTDBdTBbXEkOcYK25tRqvXTp3UVii+Adh
EpUUL8csFeqz7ymX1paPOC3XOYGtUZamGezov3CDfqI4jyMg89CfMWqmPtqU5BejJxLaOyuUWTej
id8Ze203xVMOP79nc3cPN12aUvZk6m5veovMKrtS+LOy7Pd9AunA6P7OwuUajCEGK+fJiNmvSxXl
JAlajTuf5+lOb8YV8JVdKID0vy5710mky5k+yV9Ik30hZ+R5PxDVCXtUKo8MNEEx+mk/wl3yK+Me
voHOwzImBO7LmxC7KAki7rNai6jw/vfO+1ervE7KCJtboq3q8Vvq5cNloAqFDfWDjH2uuauWhL/w
DMRfS/1aB37jZwQ2jO99Ht+wXXTMr1WeEAIN1X7yyvYEXeb/Gqtu00rTr7uL/ebw/rMTWPKRSB6F
OoF6q2eeB/Zaa7B61vOrucN9Z9vbOKryjxAEvrThn1MCwXb33+zJJk6o0hGFPmC2ca6PmMzTHV5F
XSm8w7lx27417Fr070/ovkXsfoWjHQJP9BE+q6PUGMaEdIuwSqP3cq9Ke1zfJ0UbvvGQ0/MoSxrh
ojIzYE4DQmxNsZWuPyXpcapESmAwDptbAOEbO9qKTpwzoYV21NSP7tCsZXifgt4CZTFIZ+O3Z8M+
GDOOSCOWSJDGoQD6jzsqz4keqPyThzBjDZDMcy3jSbo3FU3P6pj7PDbe9S6GFqeNUcAUWd21M8E5
cV1q5azOK1oXqjVzSulEdLhUkHyJr+W3wI/BBp2lLt8VJxLzJ++VvzU0KeC48BqGmNOlsxi1bBkq
roB5yP9itxWIIXYFCrgn4puBSuERva3Hzq9eGaaKENXFERBfmqmYo6YsTuaCb5Zgo8IO4IzIyXO5
q1bhJlQ1ayK+PndufND1mERGKIlJdpxy0c77wDl+/p/dkKS3e4ziggzdF6C59+HFWX+FAshYUwG4
pt/nvZ11HAJyaqAtmqodYWklgZ+g623JkTvTOAQ/kHUqZ0wuC3ES4A3WcSVpb+9rbqdcccjDjVwD
CIid4COS+SZtyRloxSZH1Zk2kkl3KXOGXsRyftGe7FTEMB94FkdTIimOmZOGAI7M9wIEUA4xlOpY
+OKBsEWXcgl7wd+seaduoMWgSIeR4r+xj8e6LUBkcc9jptSx0QarcP/xzDJ1FjKpXQa/H6HmESDL
F2iAF+tRHjdJSP7mVngYBM3asw7H0XX0ksFfJIps34Y7PofC8cSRA90itL64h0VzekdrDPe1v4k7
KQ8PwCuQdE8YDQ47acinH++xX3L5pHpieyzn1WqxCiBmS1G9OAYvR01PEmRU7tVgF5LicQk9rWhy
s5H0Y4LuMgOM1bA7fqWlS313uZDxFu4JhCcovaufEBiniBK9Kvb+rqL4rpA7iRRjbyw8SwLLg4SV
WXK4v8wpIyZ4k8F+Tpam99IjdMHycQJpifOvElv33RpdndB1vkMK3DXKNDKPlvdeH48mvq/beP7K
IUfDrFfxl+JrllbRgb0ybyCBX3K8WkSic+EHEzQsDzKLczqbDOLOVhPzS9Ct+D62UBQniOZTNmDV
mMOZ7nxOVTu7LGJgEYGOy4A9KtVsoxe5I9mIYKxKhhGR22C/omAg04SXe2cntBUa+Q4qv7wzaVhQ
k1zbGfE7/Z072Nab3gehirKHKhzn9aV3yUphLJxFX0DMHkBl2+KfiBfyTU3fmQXxfEbVLTk3Pct+
Ab845fcATO51SIfO6vFAOcWqJBh4XHyfj5JB5hlXgI4vfhIql6bR3RxwFLHthS0PZn1BXIFSnClh
CZPB+NohxDnhYNg0TJ1q6xnsczAk7Vqa+oqikPKncGfDufOgBnbvFOkktP3x8GSf1tHa644qX7Wk
CZoDENA45brsjmUKY04sofqm4F1OJTziQGXDbfLOYbxl4CDH4RULPs+nV8+l8eJkIf6MEAGF0ZSn
a8iBYlImbjXvqNjHwUwmyOEm65+oTkVL2HfUlPxvGR5nfTIYsNB4IYUGrv/qDAfIIAlTnxDTImc2
RlPudEf+F6q1LKCRxVO5pFXqjJfogRfomJqlJBZfqx6fThjSiop4v4SxQ24IjQ5xH74QAgt97CrR
oyPqPIaG9bPvJwdOHL4UupFjSKcEEIERI41u8wVxXAn02Zu/Fx9n0cESF3LT8fXkjBT4U0WVHeHi
L6hHAMxc/2JZXtoXt45VWl6FbwSBh59eOfFocJPDGryN5beodYKbCJNMMohIPhbk67oAbX2a5kXQ
/SlFV4xgEy807nxVVTuKiaI4BJ4NuvA1J9X+kGgtdImg9YHAAMDTsTkKUH1oED5O0ziG6iO/Bf2k
oBX1YQf3GMaetenra52YEWAtMaaYjKyJB1dsbfPFUQZmgllyyc3BOMlvmKRBez3aqKJzTOTTHAAk
I9n9ikn2azs5pzW4too1+bB3bfoEjuJXD2Sy8s5Xn1+PV+2rMiUXicW1tpWQDC2fzP06e4NftrhL
GOINtHKd33MHFc1uB+P4yI3Gwc/jCp/0hpsVuB6yH+/hQhsDZ8IVxJNRsUweNADDfYPA2kA3hbQK
91jTk486hJp3yU8UK2ifmCZMXnoiBkdoTbyn8IJ1bAgyvyvYLb8L5E9FDtO/903BTmybtHw3WMA2
WCI3EOSHgZYoAVx/uQeXA3E8ZZ3oQpen54c/erHg/6QDTlXYiLe7d9hwhojTp4hvYGHgV03UQz2g
F1sMqIWc3+Uo3YU6an5eZOVDVM7taZdj15nmZfydymuwJ1awEplPSeULPemf+g20NQ2WPywiDVRm
e7VcEczuzPpfVJO9qSXJxVuvocRuhMsaoarp98uqza3Rc+JXHynHYSg/i6Dl8/SPwotJkIEnIQzO
K818DDbi3qJ7vPYSRjU83040sKNtbaNhnNbcJ/jXxKP9KER6nF8zR8U9fBM8/X6i+bIW//XfBJma
gR9IgFCH6KWKbQsVRtpQObbkTaEWWERQk7ke7qb9yaGzEOTFngAIJnIf0JV+RbQnWxfn7w8fpue3
hWhqwFREC/pXF7jwuKzBFt3RQBvtQm6D6IjI4ziXCK8vzRVROzzSpRP6NfEMJWfV7r9SLjTLh6dM
JuA3PcX/4V0rbs5aXBxnhHUDVfFnGLtDis5LxkXgxPtGp4ZYEY1ep0RMsCHz0H38vVDGxF4fcjiB
ob34ifubsl+qCQ+UBwVOyh7vanmz+SASDTK/2EU4HzQ3nJeyn1DC3mVjMh2Zu/hoVrKhTKGl37ap
fKOlDxdM+xSxnAz5pT2pOzwjWIWzxO+LmCLScke0y7M1sh8S8OFIrLMwIjBY+2zAiXWkYZFWFndk
cos4CxiJeCpxSqMgDeui4E7LRQmots+tGEn/S2uudmNzKpTPsvQV8ryBjb7zoQ72ZTrUJ9KFdxxU
wyKqjK3DgNFQBTtZv9VvfFMbiC+eX4i1Zv1xEhtkdjUrAEW4IdBjf2LQCIwbxNk85QjoX/HvXGxp
Cs14S3ppeVaPags01b4FPzQnnoWGDwEBBdQ4MpURWZslIgRi04tTS0AaAeI9KqigWc4hx88AFiht
ippy9WrHWHNPDkfQA/dSKW1JFRD6aN8653w9qj+9/9+X1eUCFQtGuVGXbQ4q9EsWdZio1NTQLGvx
cv34jFSlxJGq53A9oRIDSOXOXVlvpYyRnwuYPdSRXRlL4MhafSpNhJMazMNBdTyGT5nW6vJE5abN
tS6vFU1aZl0Ww2sXGwDS38GFdPYktnoy52ScnDJt94WnbLfqJGheB1jZDBA4fi//RtDosoKnI0kq
ayB7vlooUkL2/bgfueg6mmP1vO+PCAIdJ/Jd4J6VSeh1UO18XuMjpirgN5agChXeUpzCUk4olxVG
8HmPrzZBYssQrfAJjj1gipgNiJBadB1igrYps/8x31CylZmxU1SC+zQIJlqlZoNL/kE8ZvO+Qz8Z
cXsyVSgBzBRBRB76298R1nc9pyWf7sDBCMQzitAXYjDrO6L0LgzQW5eanh6aY7aY9/QFOh3WbpPk
bhMRETfeLAeVanGB+e+Pr/sU4UpXjNK3s93I6hhIXdAQ1uyzE1zSLsl1L+KMTzG0ADKJ5wrFs84D
jTxB0JkN1YrBzw+fp4U19TMkVqwn9xvKFUe/p09lCoQiBP5ww3m46LSUj997Rnit94pCdu/R7+Z/
T9dMYjZ+xBX79PoNxsYwoy4Y/6Cd+9UBBFtvNXCi3zeIAlPS8tsual4rERo8lFtukSmuc5Rbytsv
KC8lK5T96Fp7sLhtVgagXOmBmmoJiDwv3jA0PzCqAqaYDBp4UetLL//R4b1a9FIXhyjLNnUCRDVT
T5HnRvxCYneusHhdhbWOKSbQruvVaZrTAsQhhjlHwPvgggMesU2mFlOjoTgPNLnzyMd0RG7F3YxB
gFWDWkyN/czgipMH7G0U979GPbMplimw4zixsD5eQ/Gg21Kr4PXX4E4SJyZc3Io=
`protect end_protected

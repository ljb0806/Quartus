-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mV/OIxL5/j1f4NzRyTNqZfp0eH/NKE9mu0xj9OmGiOUKKgE7B0fPErHfTKDCafYGoOWBXOdNLZ8L
PtwzutcZ0ti4bGEKD3UMCpLBFGHwm8ALXy5KvlKSy6K98EK7/wTshJ3W9JuyBmsDhmkZOethSl6E
Mkwn0x94Jx8T/v8M/D5BBhYWlJa+SAzrmNuAAN33I6exXL81nezLBOwk1uU5miOq81ChoLdl3UJu
C2xCTLvM62gqEUKCTzQ1rT0wZIfsmjkJA1yEb1jVvNA1oGNAIB0QlNCIyZIJsrM0BIHhgUsaodqy
AHzNFtG3nilPodY8fFjyvPGlZ3jgLnKeL+pbLw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30288)
`protect data_block
JxMDN60PRKKi5+rU5at/jhezAVJffcVgxO0D7WmDLPNkJwWfmuD9RS+jJp9K/ANcqFqXnnFCuRg3
MgfxrCwwsQy/FRg3tEuJeoKTQ8UTO1m2bXJNyxDV6Z4ZefjOdS/9alGkxFoPsPI6g2Jvf7uzW4U8
smQAcW5kwqEw2R3t/QfvYRE2qfoEUN6Dau+kJUTklg2vATqVgh7k+ijrx2mwuB8OOn2IR1KDBrEV
fj+gBPD9Z4f/7k/DYI8HgCg1mH4phUIdUn94BlY3wE4RjVhSDo4WX7IR/Z/bLZ6wmRT3nkiXFZoI
YMc/7nPcAtKfn3y1IGWwlU+2kna4MVtArP9ToWN6ISVW8cKwJxp39Jj54X6T9JWuxiWXYKXP2dA/
UmoB4ehNsCzp+PbkDNYY/Q2M8nhA08WvUl7hGE6OjCyIvFUeY1KmLmVGbj7AvQiIdzjVShq0zwZU
OE8jA51oGTo/dutE6QY7f2dntHv4Ftc1WEBMRMmJADaGtezWOUltx2GoUY4hOrbQHZaED5ZoIQtF
RvtCOf/rhcJbD/vk449vK96iJpYLKWROecXumWYZlEWMXYWTxy1fBJXqG7ocJvvdgexfSM36fOjZ
TYDdqLYARL+Sip3xjCHuKIMe2uZWwRyv26FjC0ThfDCIAMn8XsDu26oaUy8VwAaQtlR8d+QWXehl
6kXlLpM1AysNhc8TxdkRD6qPqjC331CmEtjDn9R3PNjO3KpB9090DCCiaP02iaJPjNH5X4WE7dTF
Il1JCRDaFMr/SHFKA96w8P0+6o/YWcqr+stgF5s9WjXM4E4BaPXMQzhHeqaMyrIl/FOh4jgCrjLc
Yvhgi/8C5n9v7JdpmbPKYXTJl+im3ooP6mYfh3a0E5DgVFQzwKCoGqyZU51o742re1YVHFtk82zu
/oLSgB/AHyJCtkvqHHszGu74G5OpVmIq6g3+6v1+jkyhBmMKW2H1iqF2XFl+J1kcq2P52A/CUMTR
+Z1XKqD2nluJSybuFZcCsV8H9U7ebr0dzRrJigi24XUgHjY42Tegl4m/ZCf3XBmF2kvTL1sUJsD/
nNWloSV8VSGtT1TT/EP94qclZcDA6opfGV0L/Myp2mZ2EeZMOe9b8KjkpQU4bAcCZVPKw5ssYtF+
PygTUDs27pa7kdSiiIIrEXl0/n4cYLQR31ucL7BdqIaRIRJYgLh5LS+MAfE15H/gGT60y5jppru7
bd+0bZU1AShcth05v3gmMz0La4KdsCUtj9Ts54eurBNl4d7nOraHPqRcrCJ3Cid3K+Nq2fSPi+3v
ypGRY0p5hW6loe5p8AfP0pg56x8gc5RwjA1QhwXAqOnH7J3iX/Fra6CSkHgWkdDAZzQ5etjiOXBE
scQL8NQrnlY8tmPAbX5bk64oaERgKukaT4S/dzDIgcxAVxXEkRHy2ds7VoQmwayfcFbjT1vlLlTp
ULYtBNRMy9JBASAyzusUFn/dM6XepdXvQTfBm9kmY3744B+74813TEk7sL191ZxcPsSb1iPuYNRR
mk2SnZNyGasVTzWq/7JYruoPknnLsU+R+fzPjhYwoE/TXYcQnU5iL5MCZvymFRU7dQ5PTtLDGgRC
lHkVUgbuKQqHWsfrKUlqGC1zpM/VD+ehjthnVpcYwQRGEYqXTHk4J9QmzhJ4y13rQ3oFpa2fGMAN
UJk6TS8/X2HUGITVjJbRx412Z4prMkw8Bi6+trx9ZKDw4lazqoG/xYnM4+RxzbK9QOxFLJf12Ob+
0G8jhLmoh81GRdq5Qw9qi2jCO/pRHF9sGRrnDAZY4CT99tqND4Ez6qYeAqDyUJYz/1c0hxu6Pr0M
In8dogpTgbD4JbGv/+WCFGieSkSvJwm1aFwFco5Zu2ZNPh2FalSADP/8/iO1jDlk5ozPw6cZTQRu
f9bhww+dAf8a1k3Gn6NLFZ+Jy7SfhL4QMBmBb1FfRFQTvgykTHiqd5YmTxYcB6ivf7LjMIZGXoI/
cijv7tQr7U9nagEKtxmi/DmxpyhZsngt6IoUL4GTvAsjZd5nxaSMbXmC/ImeLCcns1+KDkPMx5uE
iQIutkVBKO/Cug7/AwNVvkc3kxE93/wkEgVnkdPhw7tkjNevi6Bpu0Z+gqvBiGZxRGeLZOMowVjo
ZFyxV5nmX0KCWHSTPQL23G7OqgNM3B8c+3WY4phHm/Cbs3J4YUlW9s1dkvC1sRFzqsSeFENwEfBv
cNGY6/wFUTYxdmofg5IJNr/hiXWT0+LDrOKD7rKmOk+F00YVY3CMByQfynf5CMK1JQ1GR4uVTPAe
KDQm+VMUXC0WI/6g9MJiD5mi/z3MOUVndcDWmtJLusjPSWeby9ZnYd2qsjCN/9fzxIYkedJz4w0T
xGWbcs9XOtT6d9tW1ASRDKFolDRai+wZx7jM/L48F8NS9qP7uoqLtEsKdWjTHXnMOQY1CAP5Z3ml
yQev45/RbEa9NYztsG8bXkQw3jEg43gHhXm51ZLvH6D8Qk+x1GsEEJ+UyIKKuWmm0bsgP6z+VHSE
WQhTb7ye6w2nhJMmbdOHUJbl6wBxWmEnPzeDo4nkGXK5vYt1B6ATlio1kGysiHS79ts9FQnWJFww
VUs8drItIAOUtMnr1vHiTaIYK4juaSjr2KtpftHigCilrKsL6dDDPvtwxFgs2dmYuoHUTTCCg+IC
ap0h0UGDgzgvrIZ4BngPqKkaJ6Em/+RCbHcve4lAhNR+fpQ1bLjVmwKZqjbyVLF+dk0dZWuuz54o
ulJJL1n+oyGFlcOkl4tPRP3nt5SZmc4wW+V1tKYzFFSMVO2YhvI1kYUCVHDWClWjpoQXo/2uAX7w
k3iMMd3m8jsR4GcpO+s61ciFwtYWG0ic1U0q/40m/ci+8QzijcXs21Bhvobj/QJcPvBKImmEL/sy
aJmdR6C8NGLPONwvwdXA3suZcrZeDRjeriN87ARoyMdGJVbkjT3dkGwJyzBGXOj9ZbzEVU9qlkYk
Xi2CYz6HTaWqc8nBxuSuawFSpzeyfH/OKauQgjqX0rDZdkHTtfT017mqHoyF7Dv0TTXtK2FLDYGJ
joQFg1mlM1D84VWtiThKjKeSXyvFTiT4NGuk/Tg9Pyi/CkmH982KW6DiTGUIAQK2Bo7zejB5q3vx
LSfe6sxH5qJaTXTB02iJ9mKB0fu89rwmU4bxykPQdiN3RdR5IiTDgke2Qm05t6GnjovwSGQryzTK
hopTZZc4uQXxo0f4rCRKx8m7bFW/kD743MivLF/2OXPGUeWkUh+AVxbA1gH/7SrDAJ0PTeYWRtps
YJBS/kll4j9aO+semKcm5eOIVEpv6mMTn5qg3jvN2CJU/9MDENdE6g9DfDRx/rU7N3lLDolenjPC
kUuE76q/s43C0zbXEY9R4Y6qLNmoOMwLjj4ShqJgnySxTPoafYVPCeqEQfwuOlP8qW4ZEmU06/Ra
ufwWTrrVON9Ad0x7BLhbsRhXD789ZkzegenlrUJxv88ezUMshY2mmXMF4wRxhUqO1qQpPJ7SPthj
tx+fs0NAXk+DRiCG1TsWc2v3vgd3cVQsGDR62UiInYgmOAGr8mbT0MO/GYT4bD7TBaZCyOmXRpU0
aVwYDhp1A+UjQpnmpaCrve6n3FL/06RtWCAcgoq+/9j5/jmWrfSOacUrJ1KOgyY80PjF/EWdCff1
z/OJT5S81gf6KNhbqbLbWwkeuQV04RzhobpM+N0xUQZnR14R620w7LDhIX32qBMX/8O/Ez5X1iUD
D3F30Iis1brFahzt7gMZ6uOIIt8iuSKauaLI7HGCPWEn04O/KIkRbxGIdaKQOQ+Q4we1lGYX+PWU
BXARgMmgQpM4BH6dm0J9reBdG5e5aKyKglv59ofvE2niWeqIvKH3lIHLy14IloLD+Y47xdaaAZjI
l0wgoLWgbdFwQzAGWniKQsTuwRYfU+n7k0MbPD9pKPQcl996u+Eh95CKkCH7KzEQ8SdS7HdLDaIh
UohyInyDeeYWAMRP3Dc+HN5T4ciszrLECUlMfPBGKQLmSu0ouelYhXZaKuw1EkoWyt/yVnHVng8/
hkHtE9ai4RCQ4bpVdCtsDXX9jOepD2dCvl3QrrisI305Qt5myWmhY2L/awQWCIm6QXp3FpuLrxLa
fQrE4D0B/kTOknyUwPZRzTyx04ZlbVSVVVj3fG6kSQRTewgYm2IU2Pv6WouOpgeAbijzrCwxqzaY
JG0yxs24jkkj/OSBgGmxnLz+uX8yItPGL6lm4kim3eAswaiH50QjvAwsCyV7h9IQ2lJLqrGdC1ak
5t5e7wuz+fzOs/8HU9/LKAp+Ex2PIQBXHm2yd0Wdmo8JusOQQyluwejokS6yqkpJMa9sk+bnfLE4
lZKFRpnCByPSjFgLYmhoObL8gs+Z83nUBMYA7JAVpPuFUA03y39OUdvFtzgPCzXu7eSGIbDVtPS7
FGcyCLZNMNFQZpA4TxUeEc/2ABmfPtYEwskSoFFDiUHhJe9OviGA2PQhIOa8rf5PUcCKYNiHXoeP
LNbPOxnqe1cOGzPDHSh9BDrQTI611NRJNfL//Ny+obKFBPYaZ3SfKyg3AKmunH2FfYXwBAGOWZn6
4S1Eaf0BYBhHTy8wS+T//pJb5eVREdhq0bMBSzaEWu9c2qs1tM8y7AOg4wR0YDwQGSmY65EW5JUB
r4qIIEP/PtkM4yDeRt8Qpf7kjF1voplWqlrm3ksyi3lJ/vPrcvbcKY953uWzgmIp3GQz9iMRCkfr
TA4D6ak5TuqRSSPM2/wdiVfVeohg6EEPpKcWYkvdrLWlnX8i9fCQQ10svYTsqIn/lPSplsNsnofq
JG23O7r2GKObeDuPrDNfnfoPDppeoOZvUaRpVwH31flz0C1Y6u5mKlgtBDEz2p2pv0J7xp5Jk7E5
M6Tivmb82NS2+Mqpd6F/5MtC5stxs6/tm/PwFIUH7oeK9Fl4AklXV/B8gL2REtgn5WBtczHTtYnp
UP8QOecGVc6LUIZpCswpdIps2k1Xta72dpbjbK2sMn8qA4on2/mSeaKi43L7+uP/DiXUpH8iaQsJ
vHsXJfA2p7W0I2ERmQbLchvqfFYzhqUDM1ZGtbO6N5JROS+jRp+NFGBlcYYwi8ScJ8EQVM8ApsJW
ac0gaQngB+FIAvCb4boWBtK47BYyRgw/sFVhBT1eaLZYJJbE4w+1YCMDD44NU4tjfFN7q2nXkYqI
5x1ZdWG0sixBww23AiaLrv+4qYSjQnYYztrdDB5uGVjzJb/dgduLBgczYrbY6eV3fU09EMvY6t8R
2UEuK8tGwAN/e5mu9CXaNJ+cBvseZ2MC5XLKW9E0K099yFfJKR8X3XjtKep8AHr7fDQ/Trevs3af
GcCvftEowff/VEJYP3vhdZVcn8Lzy4V/NhBlZUax590Yx0D05CADf88/akbWzkk4VlsNfPN08c/H
S3jr/Q3pSdLFaR4d4KhV99SnhxLF3HBiWU8glIvWhuP6ZRCJwWovcU2Hm2x+CBC0/CmM59dUWJZ4
OUt/Ec8c5GvQ+xH0IuWsGLAPHsbyKRXHMLaZ6z/xUq1X5dQ6rI11oHzepiOo+e7nXB6eSdDDaZ+v
s16Pli4nUt0TrP1H5IeE34e/UZQHyLDp81nWiklIKYBujkMbw2FHMfpkSMHeCqKcV3kwaGzaALkM
QS1ME7AAVc2e+iaBju/bM6OH3cXTpRWYcFJAnlZlbure3IAy25vKI4BHJNjiflrklVQ92DEQSWKd
sou8IdXA6zvGQQHXC92jFiD0sOgjdbB2RUxMyQZxGQG0hCQIoe5kj4+S0RlbIVSc107tsQr0jlEL
deNSH3DhDKKppGvEtnK4Q3ILa3DASLP1XVQthmG0TVmWtxT4d64aNQoPxqicnd7KJ2AexomM26Ux
9FDYWW/pp2XRdY55eBTJ60pWWXLRPKXKx5pxmHq4gKDm4mVcOfO2mktwwTShalXjMKOsyGZm6AAd
ZtKsIt/8Mtfo2HZr9XoDj0ZFCoDLMnGHuUnm10nlz1vTw8vUjvEzG+Khb5aBC0OyPWpB1pLmjp9H
pz8QcNqFzzghMyystRwic8ENOyIJgTIDgrWxWLhXKv0VJonFCli3wGL3TXUv/udGj0z1Lf3pZWaz
gU5wk4PXrjueXUPdq3AYKL5Z4nk2ZRTHv0EX+7XcDi7HAviSmVIrrYVb92GTZNUnbjaH0K3DgRov
ydShbUJ10yO91lFxIecl9xLohM1GpEmAiz98lJcqF8Xz6miWU65l0QLDTinaxKwykoVvMZGDUxFl
HLHsmG3Rie4IVqkmMa9fFHQQEJqEu8TJVEHYzxvWvLf6J8yj3DVjNV9mohUSbbS7h2VXRjulJoaO
XopLWMuZr0vSUmfidp6qqe6pgkrkN9IUUX/MuQR79AEKWEWpqhedy3UjpaKbRHwCL05SVMuCc46S
xEehsa/Fq72PiKznV2sP5vzmrtGOn8xsShnQcG8foorHlkFXXR6bKWPn1oIa3fqhurdueMEkuY25
5t+A4QR3O7k8JPYLusIflO5j5c1aAIhu2YatcBAJPq4kHZNQZXUvB+eYyMNb8CSStjLKoUvrdmZH
1Kwx/9ov7HnThBg7J+/3Cv8FaLuecK0S/ZIUrH1V3kk8JThBdU24flaicvrSpmRJPjXlNxT+UJKn
5RQ6xgvyAy/kXDI6exTCtn89X4adkk5ttJ/rN09KijgW4OnGrxmahI89VHos7msOOQrEft5Uqj13
HihCE71fCQgXaKrui3mfCE8uZ6trKaJXV4Bx7KytrOrqnAn4h6k0UR9pKRngl6UQl9w6Ha7lwrHb
xAry3fQDzB6WVkie35r4DhC+26Jsf0Ee0kp0VHSe8rwKrKFM1+1i80m528NCZ4EbWkrb+pqjhorR
YoKIPuyXn4ujm/Ul/ToIXev1/O/HU3DzIyVGwWAGQJZU4H3WvxKBh+dMxTSEvzgED6YOZPmLGXGM
m+BTjRKjetR7wUhFPFdO3LLKG38sXy1hb4GeReMc8lrgxnaDPJ0RvVnzYyVpof18aac7vudUe/f0
It9wKuM5gBMcGO9BWfQ7z24yA4HtgRQ9CKVvGVF//pQfvxwcKRCRHrzloyFKUtWpdKZUyvdc5CxN
4d1CwjevuX1kKtSQu4QNUE+LeqdBJmaOCGBzRufC9rtTR5QQx7Ok8TSKK5chIzaBXa27UCZvJgbT
J68Qa8+YxqxOPXkk87Efl+4uHZ5tNsg8qkxl4klokjWToykMLgdILuSs3UN9euvN8a+NRv4CML3+
7GYyuVPje6D/HkjAmRfFEY2uYcWcsSWDo+OWpHI1eoEGXF8mPa3fqp9A074huObB5FwF5hGsZ0u6
Gqq+7TOxQUfh6asmigemTgbo4g9YPUan0tMF96PlmSQE12WAjBM6ihCui5Nu5Ja1T89UgXxCk8Jk
ZhNHq0ZvTZxENG2hi3BCsqA+utMg0BVRjeGYFQUEoirJ5hsP5uyph78TD3/o8Z40VWYE+uLK6MXg
uLQufAoFWt4nlA8I6WcmxYZ7AWVxqyZN+hGMfNN5bdEslMfqihUZYFykLWMpmAQsZOEIPmDa6prb
R3R7E1rEMpj1vqTBW7A3XCkz0eXJJ3BjeFbeEKyo91gYPdpGSZqheE5dC+vYobusxFRUpBXGOtj4
j3FMmYkN+06AF9qAM/HLQ8pw2BrU54O9FKwOqlnG8MnswCqDi+K2uayvZ8GybUwZaDy/d1N5dlmm
2waPZjs2jAxC9y2pENi1o4lzTrANOb5aZUhwBt5JNtlv1GbrsPIIXK/ynrdZUeK653kHcRpHMlm7
UaG0Gmc4ZeEqYG97jz6tMjQKaJI6OtV1S/Y4c7SKaX3/fry72jB6Knfdi6FgteoKDKNasTXl8Hd/
dzDMmzn7cRqb8QF8NUJXDQn0b8cCPF228MEv8KRaEEV5gagxg5KzZ7/OqyNPX0f7PkfOgkUdBVb0
fLPJdrlQ+X8L+8KzYy0BEq6onozKY0Nu65qLFCf8S2gOYzpZ2gwv+gP13PA7HFaNSnKbqzZb+7TZ
hu/SUiY0buQEBER5ExWCqH1GnN0ZwKk3gV04skAUvjio1Z2W7UEOyf//yHHaf0VpPkIRy2dWKLvM
+qpOCM4VD3KdoXTzEe0rIbZJ4uE4DeFYT+AIylGoIm7p3P54HZI+diN/LmvRRJ6H2eGAG7MXvqOF
d60cxGyXZ0DTcWGKnd+urLCAQLlCTw7/M6icc2rP0++MmudnQ6bJ+OqH4YMdGhP0f7S2tFJncD43
UvMFYCAFUfqxzgNidCgUfBb+U8MIzU+8+mT0UTBoGhfhMG3k6M6HQOaPVcgA/IuX8i937ESl+Goo
ZhEGMU9l7SvLYqYwa3dDhvYqoBmsFSNNN/ftmE4liTu+Ph1u4t6NvC/8KE4D7f6K1sj+8cJq9g5T
jSlfCQUcbhUn1wzRBoaoJ+zO97wLfBA92S/P7oDX3jvrujtC3xRyTjevWWSgzvy+81+CE9GnhmwG
XBdXKCGv/8DNCNljchl9TWGNfOCfbxD8FrO4N+O5ixbtGGQtBFHprLUIlcyTVKZacR1er5eHqTYO
ZReQWkcFHjnkHbfLCrDhyxFC8m49nD++LRtJyH/yRUslrox45ln5zcdEC6JgAGXS8801m/Q6o4Yz
SXXVtcsRJvPjdFz+pbKvj4igIqxLkWs1rg1axsfiGLfgPe0YwKPBq2NT35Z3Qga6okS2VXK8UK+7
QVmbVf0Y7hVaZ0qxxceOr8/zp+8Ue802sluW+w1u23UqccESKXBm32R2ejK4AJF3OBpmEP/4bJf7
6QcCuozcXgc+N9th7ck1zMDu89QI8VjoVauy+0pWchUFWccjYOOPOZCsiK6S+pRFFY1eFz5bK9Y3
xQ1rBIELBVa6Z+L0N5ypE4U9+xLT5OqHLjj3DXWah1EByWXigvG6Gbj2cXSgsOj3GXDpY5rwOEuT
c0ZYcY0txAcPoq4gWfQtmwRSrUD7CLoYV1ym1ZaGKwGnl9Bk8IntZYBOpvq/3gWqtBvIrjQsegBs
C5x7NKG5icurYRgWUrH2oiFfU56jjB2EKym63XfiijPmTjaKOL2rqDIUGKPbx+mv1SZVupah7JzF
O9g3oX6WFxQirHr96jIaspq9Qp5EIv6DOgYEmG9Rao2OXiNSAqxo3nHoBQONgRxjjA5Pi9Lp8CZJ
rx4sIFfI6k021JbA5uKdWHz+2WMTh6Kkem+Cif+Koyx9dKmG9frNoCFYO3sls6VxVBjgSSEBZ8Y3
q6z6dyz9O14MyOYwiH7xBZ1UhztWc617L+YJG73IoUkh+PAO79K36hNH1Qh/M+O5TF4kGeygDOTX
Ru00wzIIXNrksMoe8mL3E3H82uDFaQpal2PaqUHGwjzg2L/EjbPdUf/BiIN2tzcENCVcESIZS2Kl
NYI6Ut3IXbFBKwfeRVS/dSp0Wyo39lOaYz3fzrjOupNVdWKVjHxrZa6AhkYpnYAS6OQTHyatD4gP
NLNu9peN2gZd8uud7eAJob6hptLFs2NVj1dYjZmSrdfY3SFMoR7J4ng44n7XLtBEFq9yLVKvmVtp
wKyCN5hgYbvWOp6E0nMsDgrU+ggxAOuJLHjonBnojXDosf8KbcNqok47n4d5foYXM60GSZfh4GUo
7u+iayYIvFvayIHzjL1+TKZYMbw86HnbPvEx73P4Vjg1mn0kRwPUANvCccjs9QFXsNukQR90sDeK
1CAmpGBaPmg+X1oEvqzkTPE9bVJrq5afkx5SndwDGfWbZXfa4nVCh19C94jaqTyIpGt+FShHNtmb
aToYr6fuYatJDb/TZQeoFDp6AKhggyr85ifseOXnb9WKkh9j1yXSTwuuR9/fjOlKeLWcYz26e+hm
mL3qyjLFgPDQUkav9VVRX0xBNLfqMpd1hP0X5SJUKh8eNCAIw2uLGAllrAcQfEfGRjDonRs3/4b3
tXO11cYpyAWl0drFsOYZ5JaMeYPSRPRFD66U40ogbJylgYul+7Bz0BQKvvrNS9hK1lq2oY4LxnNs
lJJZXmeFGpeuJOMK37Vt/1Qwg+EIBvY6ZtmZLIJpjN//DutIKyo/r5R79344TRyMIk2Pl/rQv3jQ
yLk+BLu3HXihNrhL8ofNuhdW+oVtQwl+V/52ljpo20FDWPBDXI0E+ft1y0MZewg2vJjz3u079dQZ
9BZ4AijPU+xhsyVbRU8zzfLo5F5grORP1BovAv1HGdJzfPVrtHzSoKIp5ley3RTAlrRLz0mNya3D
+jCM9kuO7i1OeTox8Kyhwuqytueekc6a2jxc+ID6U/lpgR7V8mF0I8xeQU6KY7MjtvWMzP9sGs4d
KYh0TPqEugJGRo6D139EHNjbS017M55xk+jkkPES68mzy1PxtTeW8MVQZ8cdhAyni+w7eLbbOfOs
ia88sUyBpbTg6pu5LjEdWyrLsC0MgZJy9EoZ1jURm08G4ngLqdfLwf1DQfl7u5AQVDcB0KTv6cI6
Jrg2gzhtdJykeivCHqe6899oAg5ecwVF+m8f64oZodH23zQngcLRQZ7ebiHzXQEsv7SO0QbGN1WG
/5xASc6mVFIqDOQC13ZJZDF5oJlYS0zbdGGS+sCNPoziPEttd7xR96opVwE5dYlECIiyHPz+cX85
cIXnDPD037t6HMg56ekoMVqK9zGYHzUrUhs1w7uBA1RLFoIW7UoUuCWr/Tp7N3+dbTfEvvZGVxHa
yq3Z/0LJbg8wFIxB88fox9zgSdzW6LlBCjGkZGuiYbcD56rHpw6ybNCbYCj2bHUQkf9FwUi/hQJy
EnnG7+GGGu8M3OUa8SuwWY9D3CJ2IdAfgpOFFPGM0XeJv6UMksLKC8G73e5DIDYa6uZKcBfINA4H
f06DOi/kZeUh4UZgOSwTMoY2/KSnG37jlKu3hwiFFUBsCKSDC4UgDumunA/0MOHvqSnQ1QLF3ckK
IUTjZ3EYm879RrzdTlEshlsLbKiwvUzVugarl7Sa9jQhPET0WkaU58UJhxG98/NBAKql+OLzMp6E
ByQDxKHMuf7jqZDWVI95PpTCzQNHhSZcsFzxkr6vSoEKE9W9ggDSBWNNuogB/8hERyLE1CqTJ02J
XLUHrL2V8MQJ1Uet4rkinJEQFMzeO6KhJiVWpUsHltEXNuvjuuAWIdHkEpxtxCJM5lsRWU/s5z8J
4ENtDs/WLOhTMFVN4uZx+SXMWJ8A7KabmJFQtAgHAXt4xSGaEHM6xIw3QFqjFU79ciGEWFEXgypa
5rIrVe1c7W79G+FTXQI2jLQc9aNbHUR9FONsaXidJmJYPH6ZkxFdjhoDbRCVcOJ0Cm29FtutcBRy
/IKQxD3EpHZkjxgmoLbLC3ako3/8Q1pxY2hbgnoa3taLi/UObpjqxiO6UiKtz1+PPjxFKKqDHuB9
+wU/MKheJXSkTM9oRlnkRnaWexwqbkvyAl6Ns4JOkKyJBjR/pMPHk7HBxTWFU4a3OXFJEVZqob8m
4puH+5fefnJdADOcxBgSQhgIOo1Rzy257RuG+0hXyZMwGgf+FLwNm8R6+jW8CfC5UlJS1xhasefi
1V8U3LJ2BJb464eDeDSWlnh7/L/RYjPhHKrJAdi9U7804q+mz2DSnng1jhU42k6y9+GfzlY3BEdJ
Uxr/uO+b74Tyf+5QrRqIh76CmrFRrXFvEQVKz3w5gYhnsapKsds5KO9eLGCPsX1c+PVugC7m2eXB
mcuiSYkX+9CxDtQyompL+72rmPGryDRFTujqti/6Wy6C6GA/FY9KKxKY6e1oYEvtTRTMQAP10vo0
iAqlIlq+Jhss6vERYdOZ4MVj/chQnVDmc9RaaP8vVjSEoHRMY01TPN3Vx0/GGY7Uy4czaCMchtGY
Vr/cCQLdszuZOGG9+tga7ECashpksOA/Zi0EBwnNgcqLKekBTkQcyja8OwAMR7G00eMXAa8GaZE4
oO6/Ml1vT0vQXJCprJMhIq5b4VdTsW5B+uBb6f13BwnDM95YwTgV1PNVhOlZflctVyEobnFfZcpP
Do7CiJe5LYghGIz0Ur4ly3GV+d1KT40sikNhlIHAAFNOkcoLWn2qFWBTkyou7PsIpTLqtv+VnuFH
CChPlIahMYVOKT5RK86rZU/SQAVYoSnww3lalLTgVsCoT+Q+ELbjoJMa9HVzgxHMrIQWOvu9uoMM
NlFcTJXFjxX8Kmpi2iKzyBVNiYAKBb5WAy2Lmuj/qzNnpHY20gqPxhwqPERBisubn4e+hA2ADiL9
l4x0X6GiNKGZ2O5BEsYs1zM61KLxv5RoKBBnA6gHWz2cbFyo+LqIsQbqtVpsSu74QnJWRnqKRA39
Kpcceu+m2MqpJaFys1nFdbt/ieoHqgnWXvf0Me7bYf2/ab60UexHrahHnsjyQQ7ghllRXpMDZhY0
6xMscnD9dtAdqCJkAPUay0kpjGLcHTVqarKCAmdKeDXDIqFEUo8wA6uWMdJJeVQotiT2AhfbTbuU
NBYu9E0zsde2uv4KLRoM78/a6D0Q5WFx+JzSQML6YVfBHb1eEr74Npc6i0d+PP3SMXhh6CVmZ79D
p5URXQ3/1bnbErImxEinXqzny6WX61jpOjwDHdkeafEVjv+dg2ZigL8jP3PGWF17iSQ3F2R8APbO
o7H8DLqS0sDRnljrtWs7mkKxgQXD9LQKHBlUuF51hpBNoOOcTDlpv2AW670B/iU5btf6p2nnYxiG
x+dlAfT7It3X/+8Q+HFrAsb+H1NLICKWPLZQlU9MOAct/NbLCHm8mKEdaNlCGZ6TO5ab7UHlyU8+
6pB6pzRNJIw3LENqzsG3b+Nw6mZTMnhSkGLme7Z0vndodaYmLTuoeLMWTb4wS+W2nURMt1uwUwkV
88U7fwTRZreOqzohDwg1oJfwfI9QiFXQ5s92sjE/TuzUd2eDSmjZubajlhawUkcukuYy//1yontR
sbhPf5/fQfVxbV3UillvJc/dZ6fXVWA5OLMDoD5Sjjhq2SVQlCcrffs0qPC9sJtQ2xUz1c0EgAFd
XOguw48zlFHJAfoLUBTIwSX2ibZG5crQAOVJIZHO9OZqaDLTPqQhcpI4imPwBDmuFbzHFmRbAUG+
j4gROK9cb0r8rrKKktkM7QpgyFrDzoNCqeDWaECXCfn5ku1KdLdX8SOilAU1I94AWkSJF+4hlUoR
21huc03yDLLP5ifTP6+xoJzGojKmVqRQzTBOsSBtD2KjaVbuKQPIj85QAcTC3rw5Ch8ge7sTjgac
n3fMgRCqBKix6rFlIDEgDEr6zY2Uop5r8TvcJI19NHfc2UxAHbVV+ArhXw0iczrSqAl+rHqAA0zo
tCAFjbNlDU+Y0NnPY8w68q30RnancOLl4bMK8pY3QOaAhSoMROK+uGR7f+EioguPQLAYwVPILx1v
laAorLf8Vf2iM2pwvLaL/je+PxeuFhN369fXK4jEPvSCtdZPJ1eVCmfu6leqy9SIPQUMyImaMHTT
aloxonm0WglHC63WZstxzGt2z3Z492RArtjHQzKFS8W0zDiwg4FmW8XCUZXQkaQ85k4YDWP8ob0y
SMOj5jrzRluQ+tqnhfEbdJo7y30J90G93Ejys2AwiOP7vdLckMWWl/V0c+52QdYiM1G/wZPiy66/
AyYs5VoReAwj2hFgJ+D0ZpDGa6C6hB/GOLirgXuQqaDi58ZiQrMxCFstT3zMkh8q5vUWQNWZRHhZ
2dC8ixB8cJ8Q4uqFjO6ysFsmy41d+B+p0kbtKEV22ljnN3URGxaBTQQC9dPTxXp9x3ipFN9SEs81
RuDMk9FHw8XO+NpGr2efIVY3aMDcEJRCM4gpWwShrRBCHAjAN5tAu8tZpG49I5lbNS88w7D2+9/l
W/61VBQYzY0zywXUxLiZdMM35ppXijQLaxJ/MSjwBUYhu3iXPBUjuJIFb41thakOdmdwTSAlzKI8
dl0F500uu3dhS2AhmUMXekrI73kLQkuFMeoZ1oC/JYSZ7WjlYBdlMIY2KAXh2uzqh0zpqidaDXjS
0TaUt1OimZ89WuOP2t5fWHiDUP44ludPp/IMNCyEWmma/WVd8adCvVHErUcTcy2BsWu749kAIsfD
KECpcgftmiLyQIRhthV4NTsELnsmtMUet6FR05gAf/53nFvbwwCmDEaxtCKAmPR5JbDu21IxGnEV
W6ftwP9PW+B2Gi0kh/jJQ6DJXe2d8dh8KE9SG1Nz8yVVPvvtWqPugN1sRkCEC/VjxzQOsDmTE9JX
CCHHhCpKJkgyZpvbQ5oh9A8XFj2uHYqpFO8Fxg5w/oqXMX14is5P0Ho7AYR7OV2oTuAKlOr6hlVt
shjjMCZskRvo/ra8xngB91f7eee/AomWqFyhhXH6wXq0F6Qj0ydEFaXrEgTUF3pQnAGBnn/V9Tsk
l6ld/t4TbImffpJV1PjAFYlulLQDnAq2nptRXuZQ5RSa/TjM5hstChJGeyOeDJaV7iLP+F1yKAVK
blc9TOOjReaYy8tuWvy/liqxehcbURr4Gc2s1j0kmKw99TCzxCXuI4CN9dnE6F48yT4F/DDxVUuq
/nlzXzqQi3QsJ5NCg5kLXK+cFIWJ8uImZmBymxuggWXwhM3o9+5ZUnWg4hxMlBZ5lRdo6ZUC0JTx
kzbx2+J864RuLyrNtrILl+d8LpJuUeelJWXYyEmYBruowlz/FznQH8+oDsJ27KqSeq0Lf1OCL0M0
Q6Zjx38zbu8gWQ9DHWfQsWdghWprygsXRoOEcX6xuroGj2O/aD7ZnSGINy1hYkxxzS/dThExOrYP
61k0Z5WSiVByIfdKJfIiZ3+5ApU43oHxcIduXlHUBJwIxb6afn2O5qtuwqGRuNs7fyVtuMjg4N+e
hxRNew6Vt0r3LfYH94B/DXyzCzLs89XK8XgEGnvYJXkL0Od6QPKNSm472ch7eAkjU0kM77N6gRPw
7vWT1unjcoh4Oziwd9ZLZj6jRS7v+ny2AjEZUlEtvAYFGMk41j3QJ8QgzUBWC86Yp1AeQFkD9JFz
45CsVjmzjsj/76bNsn1TVPV6dEa57lycEj2mOzm/VIFkjea5DzxHbxOlLUIYVOfAYrN123Nx/0HH
RURc9Gntj/HS4v9Txk7DycX4GAh0UorX7ZQFU+/dkksxcOYhLa3SKDzatICWWRFkR2l4i/WfRQ1/
FhL8OeY4ehkzlnO7j4OtKnpXmCvQcl+paQ8JIvtjUeBGCG9OmHFRtvTRv0+fDlfBL6Aggb3YGsbe
ACvaJqvWORrAySgsMxe55oKrPR7gbvjJ/+iCsuhHviF25OirkOP9FxbRD1zgU/+9SOHtd6Zp+jBh
Y6frJawrj+qGZgGyYkPGMC5b+x2O+K38yBpLTC2tnTRpS63htSWIrxjlS9dDTBIbK0A5vpjmjCKA
ElDfkY5nVuiSljqGY2BEf1HOpBQ/B/pBseufZ2g7sYsfK6PEQEocxjJJeUzUqaWjNycYvy1Yl4bT
F8T8xprhkwZ6RzQkKDhQuusS0CVJqJfCIEmbbHodP+20okwAogjktbG2hXDlRAS1VYfkHTW/VXJH
F1cDh9XQvb5ZrMVHIdyt2bIc7xmNFXU9nEFbyvs/k679fac2MsJVaG12jZQ0f0+iYhX6pmin2LiD
Oag6Cxyw9O28J3h271sgCjt7fLkFc95qpaQL4sjn0zjtKhhJBlru4WC7lp2EjVdtxnTzMrYsJ8aJ
qva0EYBC8Yl5O0RHueKQLce7wXNX0TVSYT5YkV+P6Ymw1WTEbkiVhT1kHhaAwJJfASW+4sXG0zOF
5dBeLv6slFvl9/Ci7nRd26NvVEWyCG0L7hRvNZoN6UO7A7WEumQFQzJV0LCjfRRxoyIHTrMePQkn
weGpQ2VISHok+Hx2QE45MIm0kkG9DuENSUtIJ8v55snWiMi0tCn/sJJo9TLZ88Aw9tpjxLTdB9qL
s3fC/qVpJvm2Um82K6ce4BgEVgjK5COn/rKiLD0J/1u6Jx5UbumfWfT+Oj9uqydZFMktZEiVUG1a
0FNCZl7ybOu+xYt+46v/YuosVtYpjpV5xhitVH3+miCrDkRrZMG+e94tUVVyLnvU6oqRt3ErcGOV
cImEBNvtm7klXe0UT5ugGU6E5Z8dMKsPQM2tI1gssgBJNp3NbG5Xxq88JGM2/tgGH+Fl6s3iTHTH
pQO1xYLA56fORF3bzguAsPAMpDWyCGUNELiImLs/UfYx3FeOhP+x+JQT5O6qd8ULpp8el3AQb8Dh
QQnX+UN0Ys3i3QMa0mdg0bGnyPoxf8V/t0j1PFI3WZ5XenJ7wXU+p+LO2cyinTBVvmMsw2HSGI17
xFXGIr2HlvGXqLmwsU9rqMJRVVA4EPQvgA1UHs5ohFwbIUIF5Fu5nMD9VsqOlNpZi8J/cOy41+nj
7nsIkLCc+XWEisOzJ2xu0aQfPXBC6zeS4Nhj0porvcplQNR7OsStD0I4+pMQBSmjva0PzKc3ucsp
cUrUiFqRstmiPXvT6wZKZ/F1ncvzwTBwDcgd3LymNqfJCnH3lJdxBm6gPDTxD+sUoM1YxqO0qvee
eedKa0oVHI4rMVs3Db28hoin5p+OPVXEa7Ub5dzKm+WeBOvw3swfIQHgOkGPONJMBbJxsTxBYHjz
EsJKxYH46IF8euKSQ5XNe59aF5VnBxHnPMWSwdz6N0nKeuumnLCl0PzUCg4kXM64gkHvIo/YFnmg
stCRIBpTH0lxR3H7N+Zo1Vy6ZEEPIxe4i3KUuFNzE7vHI75Iq6mVDd/GwfQTe8O/9QbHvqifoc5T
/iPwJPtMI1RlaI6m9gD6yYA8OhagBUeeU/FltQzn+5sDo0/cIEkQZI/CdZS3kvVujQ2v5owkKeqD
y2/IxdiY1aj0dlWe2XtHVg+G0ejena7ESn7BRSurNEOX+qC0iOf6H5ICNSWv+S4EvSbQV1h3A/t5
9iSFS5xCMYrqQCl4QbgBJVyBwDhjyDrZwxlG3mqQb+5q17xkxJjJF/csevadiUE9agcYE/o24NlM
OXuZog8Zd89mbGTMMJCc0UXy+Eb2JRE2jN3bvbp0ancpQ/aBS2ie4DAqyzRdConGR3lvvT/74ijd
LAPEzKefGyxe4HptVXfL4JgMF4Z0zkruukMPEGN1KoULSSalLq2JevMbeOAvvIwGsUeVN0IcqXUm
21iQ1JRyxl6d5HuWtLjq0VbiulX2FZk8X0AlVBSiPtMYileHjAFFT2jG0VVR+WzcJ2huQ9SDN1r8
JH8vmDJ/87BfucEmHaPxq7SxvuSVS12Jhmlwg3uc2upxfQjFaDSp7Pmx8c+ztg8iszlJx2uEIqyF
+e7dTX8/kqU18WbzPnnb4d76iv9ArK76QgsWlvM3OEezBfY1m8r+Ton1WCUBSemiQqXXAM6PafqH
8mgYA3kH5Z7DlU753sy8FMWoLApv4+2+2ixG3KCe7NIYF55tl9QyF0zTEZTysnUbEtylyrXnkXbK
X3Jl+5ZzLjGYjaYSUb6mC1Jogg4gICBIgt74tC/W7gCMtxIZYY/37wzebQWQV3z4i6xQutI8x9BL
y/x5FuH2hnSylp/gIfxDH3OrkLghUehztReXpxcK2HUYBqcDsRT4oG71ywflcVaN+lcby5QQQdnM
+KGnJE/7k1jnYUhbrRY/a2s3FTVckG1QPDPUCi/0nONEND8KXtv2ud/VlFoxN6b3jI9GZwFP3R+W
OdNLkF+AiiGJcCEwPiM1qh0JdSMAkuZLVhLIJJBdTnpRUgPGzPzwwuaOwqPNWSQ/ilBN0C9e1GBh
7lwUoVqpHxEH7XrT9wPlAu4cAQp/PxdgTRjYUPCwfLBUM7kd/+JCsFNGWZiMCKY1zbKBxI2zMlJH
U8Db+DOMPcrmRRotLpf3+4S4M5uc8ATH9PKtSRr2zkeHa06vivIT0zJhcaIqroqhwx7duqa96wFu
L59T79TQ+Zv2YGbaSA1rl6LWKuu6nYv+uh+4UcBzJGoqmioSUgAb4OUeGK1lGSRRTYh19vnAJ1NA
UhPW9lV94KQPQxsZgBC6G5mgonDCdcBACSEj5GWgwLqWokRrGUq3Q1x+vCAZa4Q4CzCYo+ea8roK
ts72GbzDN/01x09YCVe4jHA212hpsKyRKsWKqYRe6ZS9DGvFxThz0raE9v5XlDSGYkQ+NloI+vGQ
4OKfVdJaHo1yEEKWpWhK9pR5jVWcoXLjgKXOFzuqHS1z5NeyTDUvdg8S4+CbLdJXt7z/tkRHX2Hj
+1ScicJ2bP2mICIu4P3+gvjI4QJqAZTIadOT1expVY0T5C+Af+dDeSO0xNFc+uuwIe3GCgacAg2c
Zg490HJsvrGekhiZbSheXoUnd64h2JQOAl+d780eBEoF1Lrq6paPMqy4dxco+OTO4SPT3+VN6YNA
PLkyoYRyFuB8O+MzCsRBrskkw9HPJU2JibJ7C+DS38xyBD6uDNxUMwWC8rQrJ69m/A9MtG2QHH9A
Cr6/wkSku4wXnQFhbp/uaccrXUjli/LOCbSlm+ImAhw3coP3CKtZhD7X94RqKBCCKjJTSSnGogS4
7UPH1wmiH3V4Id5crHa1KZXJwuzT2dZLGNxXkf4hbexuONuE2zjonD9d1VVBqs9gHe0wUbdIE8J1
gWjIS3OX+XujbJXowxHa685y5xF2/GKcPEFnzF1HI7M5MaGPJRt8PfRBdXm9Qc1NcOeG5s52iRxZ
Dakzn2GEkLqmWmxfbfOVhg145FLoeW8v5a4Lexg98vWIxulzzOrqjapVuhEsy9OvJ/tk9lqCnUL7
DE3hLvyOE7PIMB7HQI78d8D1JTuXFQeX5ky1iRYi2nQCa/JNnknhY2+0CV80M8ijw5XKv32m1cvV
izhRTXkFxSl+t8NY6kNNKJWCZVbEYs9LR+2J7be1cqFcicT4SiPKjmHV7lleH6/mPE/VuKPNVmoQ
KZl+F5pNf7Az/UAEJssrhIHOPnnXUAZUSfX5icIPhzTgvsDL95s9okLxTG/iJPU7GfRKt1Rt2Rhb
RnMmLw31t9zX5BecqF9egMay7JSiMMbOtk81V8z5jrthAUryVAQAtBoHHB7/qxv/nAPLBxnCqVC2
QiaWb76tbhCmartHK9riXmNAuvB95vISU3ZpoL3wMG+wL2akdsWrMHxZpjt6XebllZ14fnU0nodu
2aIaMNaI34jLEg3zIGWDTSTuMRxtbJEUcO9hWocTZyRuzVrnk/lY/InsQG+FzOxVDsU26zsNT3oR
N3pqOK1QwbGIUtV8dP5AYKoKqL8tbsmX1Esvc0C1hXkQ2qsWLgjwgHovfOcgNjUrxUR3L3sPD0Uw
S6I9apynID4zBlDZNkduGmGF/pKgQ4x1WSDRjYLASBC26Z+bExw0MfbhIkRsN/nRPA5S/UNrNguE
HRZypWNloGN7YXRAJedmPvLDhecNTvnSxLZpkbjUFO+BJemhVWWYJl1zVVKMsMIwUOE7UI+y+rb6
d+YQXHvM2MMOKCEcBwk3VpSlqiX3E2by7/CDQy0xfmy5Catnepaa8Wtnll+DteK4GutKjUlVHh5/
5ITDCtGXPeN7TlZRvjZpb3vdvl7HYvKWm08REIpXdgnH4jqVd+8O8yKRUg+twQw2oera/t7IRVXf
VkEqKfpHxVkPOPCv2vqKVGEHY3pOF3dqwQEJz2D7tVVvG+c1J6wh9adLgRNhfA70H5gF+AgC/f1s
6rblRuqVSXpIzJ5SjJ/zFb2RQj1mJbRUij1ob++ggz6uG6gxXbY+vRn/ZivDg27Kkse4zUxWauE6
fq26ysMV4US79zCN8MbItm5cSwcY4r495ngSDGooYMnyIWXueYf9OsRtoE5eDWQsRIRypGsghQwX
33bxnl9oNUk7nZTCNBE4ljJg+VWJygrQxSmqsk4eDHQrVfBzRSgND8kvwUoaB+6znihwe4N6YjqC
pmKKKmpVrjpxyMoc2t4LVlR4djuExgSbP6Y7LRPZhlY1XTT1BxRoG3kkkfd2BdJLVnIDJrYXd1wV
G3DB1m3ylMbl92r8i6R4hlHzBBHLs8Al5MlBWv3gid26hu0Ujd5wkd9mF9wGrLmEpEwYx0PNPL7K
Svt9zYlmapkoh3iqiK1IGtbZx4zqf3tB9TGt9JkOeKQJ2k5VJB+iGSJX3AfNpe5Ea/AmkPl00p/9
MV8iZYKpciQ7KQpGTobDFUw99uYKaoQsMyVOJJ/hPzIpkdrIr2vp00WbOw4EHd3YApehGLyYEcIM
wBWoaW1uG0fmZ5ewFwKjkvdjWzTRuLtRNjMGpsRxcfK88Kqva4L1VbZ4zAFwa2FS/UgV/mEOtXvp
WyeU4hr0BXTHgMFBvn+TfxbxjBqchA8DRwYhExP0hLa6Tu6ZFweBm2zItPabNCDbg5oFA6VirvCK
+s9eRUmf5dQQQphZ3qHN6xsZ3gVk0aFKToG2tPjpBF3x0ldW2+7gHv5uT8ncHMS7vCqBT8e4RABz
mgNuoZZ3PoMqYu7oSEJARV1ulPQOCCvMJ1PFX6fgFkTxd5abhrsg9zDfTpiwmfJQwA46BKlGWorq
/+4CFIOjw75kNpdrI4Z3+f1Wy5LBeyfXecLAkHzZk759IBCDEKBJpYN63Nw3dh87rQD6P97G89WP
PC1E5VRFFc5aAcabxcCgbt4QgaYGGVNFmb7lTZ6Q2XvR42NdcKW3jsRErSdko1JWebJ4oNxr5YlO
ROynXThKp3cq3mp7tvgfIuLn2uQHh2Sw7nlcm9Ixa063u6fYCCv/DJKG1GrBCvmjhk2wDeOQ8QsI
1SHtc77eWN2lVmhgg2PWUnaszk2G9nKUiwQNkYKfBgaXwpEhZqRkm7D7y7Fjgon/affgHhR1UuPN
6NKw03tQ/QA5X5X0kPcb1XzOUjTPt0wVF2D4Itl/TIUXzNOvPm3Ukxmy1RtnWjZwbXRUpJMhNnc4
Gp17OrAyVEPQJ6xLeBdNeiI8JCSGiPsepA6ns+p6HFFAKnZ11MTj7/+yaNhdb9+ZbkeLDy+DNEOE
65aeSQI5PJ+HX70yKDtF/IZuHT0Hl+pGqwWMTKoeG6x5RW1OIFiRj57Vz2EXWTB/9FyShRBZbz+R
1mthYai12RDZzWipXdYM6akH8VYbqizKry0M+OX9W/2I1qyfY3/UjhlslLKWON233FuY+5AdYqyy
QUgTXE7BcL9pCMuLfukl81RKyTESmx+Xpg96SPU7LejrHoyX4nJfXwMEyavFwfWWKEuDji08BLdW
SP+K9joj6UZbav5UObWbR3n4BsubuCMd1i7DTByhLpjyTxc/gCwNxxDRG/BZTMSXfUd0yvN2uEYh
blDXV7j4GYZExIcuwGR+3rlAipNvHGHi9Rxlj+quFauungIdtRT3RBjsIAVIsJteYRsYt/Q9YKfn
x4EAgbXuCXO3sa+91OkBm+wc92CVjtADhuuLj2acYG5KqcgMvNPsOQNnekVLsGCXSvl+nUcX5Cv0
Ms0qXi2UO0T3W5xiIPhKlkvqaIF4gnEQONLnUNCN6F7ths/gAaEHLTFfIQF9hX3OBA5nBnkyyDLE
7N8g4WBSwfo2tLOBbUaTZwCUycgrmiRY4tVdEeULU5sZ7VFy3V2/oEXJg8kH2hfAD3ijQv+X/NWF
a6TA3BeowECI46h0qly2T4+3hVcv+78YFSd5t40TJI8U6/m8oGhPTq5Qm/p7JU8SlBtvSrBvjj6i
DWFCisoRmIUxRAHP2Je/Rlh0br/DXyL1qnHevvHgRQdvNt6QoVzd5vEujlji6N5wKQl+N7D8fd11
COZ0e8OHq0CRnF8DdOoXqdhYXwfPUhNPStFLc+FIvUTqVQJcO+xtO4wjMvfl09lt50rNWPGW2+hu
Zyncg6tQ74n5pXWTzzHwVjHeHPSbmWFfFteNAPAI2xflXibV3SbRx/mbUw+fGhVgvT7nAQOPmJVi
rzN87AR9Mfo7NBxPMlJ7PyN/ayNw8VDN4DqUYChzzQy0EoCOZ72xK35K0gthZB1jFyjRFP13tn4c
fHFPDrpQlVDVHZabphOWcpsnVPbaYpg/EZFPD3sz7GrNyMHo5KmTneiqr/sNMBR4U5KSvOYpOUyA
gEZTY1s5GjqvA8XqBeEZKsIyUE5yLfF3YnSBNY09/VTjh7dPXBD5wwTwSwvvq72HbUwngZdXpSRa
R6K3qqHWRUUM+diSG/5znmtU/6H5fy6CB6y/g1uAHOQZDWNmaOFmMLGlJxMAGFRJz0bK/V+j0qIg
+rYRnIGuFE3XouQpmDvwO+6l4O2hVniQwqd0J36mU1twNH2BEvIl7eyR9GFS56hiG9WIV8yUQpGK
DBMLWwQq3w0cyxUxxk4zDBwVuoX93yjJT5JV7iNP4T6pKxwG9NBcvrMYZ58H0XjPyjma4BdzvyzT
LTkTuh+ZyoLHEk0U1K/QDqBy7kHtIQ+w8tT3Gpp24BTeQaT5wBIctNse34aaDpMeDxMZnbA7nVkm
cQ/6Wo+3BU+D1mdLTPBerFGevYgcwqn3K+3DACIqBV9KApPnCAfUrVK30ZK8l49Sg/9D9G6wEBfD
3y2XJDWjNEeuLRgp0A66kYG+JjIGM7wo4QYBidIa8la5U7gBLWlOPgVw13CG1lS6L1TLW+2M+R4o
f6c9qMU6kAvu4H8Si0pR4/sp8ASt4ctygkQC4aDQ6xlTvIZ1P7t+xR1rdsDtDwBGeZA9pt1V8lmv
XAn0CNCR68gqFWGQSqRlBT14f08EtB/SEDbnjkMRKklKKSQgzRJavYgr3JkQTwOWBaV1ni/1ZDXi
x58fnfuW7QOI0yS2UwSJX6QozXmyJXgz99GrC01l3YZkhWWsx7fbm00LeClmyosgAJkJuesuLXK+
q5YjT2k2j2NuATQdnpXl/URRdKCgSBD0AIIoWeJytJjHmQTgn9V8cHqYMxGZIfojZPy+YApGMmmB
7Q6EZva7TSdGBpsj/A5Zlb9YKhXBJAQQmGUeY1FpPRCi89HSpKewUbp3BkjMyiFdqw3YB2z3A2nE
lMvuXUv+rTycuLTNX1whG6SEfjFEnKLaiIDugEPuhJP/W+Imk8GRilIrU4i9Spub1NRy0ZiATqW5
IGqHR+fQpXgMtzI+8sm5HumY7gQY4UP36lyPPCankFpG4/lnWdi2MOFe9SG/QFapJon9q5mJvjUL
DOXnDgI1+STDU3Z7f8vg+BezJpcqLa22fjN+sOXYsRWp4j5u+Wml5jgc3+oMJQE2GlFpo8qq2boR
S0qbRVoFCOObzpXDI5GcpAmeTlCpgK1SJtrcGXB3N8NdIE9aNdDdbSbHAb6qD8xdoIAItJ3lFtnk
EPz7ErDVWtlEuf6UUNVTgGPIf5fUUUOlt0IH7lFWNV3SHSbB2baHJGIH7rSuifDzdKbKBgy7A2r/
JQ5ALs77l417CwanSuwA+qpj4BK/IhICaCI0DQ0meqMS7zgfUJRKGJHqRfZKcIdcJ/sBiDWswtdD
Fm4AfeZfVvXmhbBhTthtwYCYiDH1Ap1TfkqRc2md2KuFsOU7nLzwD8zdqtHrYKB2LZiXsYsb7lhc
b/U1REV6pPTGLgglyBOj3bL92cLLGQPuidOvFWunzs7nJA6JzCia5C+pZgOvP2FNEsxD1FQ5s7Vc
cd6qpbwzjWOqczceMaq4cQAXO1MsINulb+DwUkFYUVA7ImFuhE2V1d1is+zsSafqbFmSQNWGNBdw
JBf7tzdqut5BmAqw4cypVVK/KO4UFMfTd70ulLMgNMJAh1eAPUVzeT6CncEr4xq5qbSRAKcIrN0b
RbOCXj1U4cMnaokGCGIrap1mKLdbyIrW3Xqcr9Yk6hPusZvfQ3R5N1tEqaKAGtTvLPH2i1ArxlAe
4zfv/WBDSX49jguHYWEy4Ji0na0reRVEfU4gno96jcukJrohVOuK8VPnY/NdmuRNpwhp2Jcn6yxP
TEomVMxVlSlE0ysgerNwFwsV5gZjqv26NKYpxxEjk5oplD57AxjJsQ7ixFzU78KmHoJ02eXgenkW
ME7PmTlNsVv5FTvBSA87m0p4Ee89hkIXnT5qybFA5lRcl+GVjoq6uHfRxlgwPjiQcT+UgF6cZzwA
yUIPCSp0E5lOAqDSH/3UI/DH0EzHglnbfPNqKXeQPRYcGVweFlslqdUMTUmJsb/wFsbGdFJRjGk3
arYIS3Ew6TP4gUGP+21SFDMCw2G6+AeFZGF6IZhWL+pEnY+k4OuEws8DidMN9mVXbAEPpqp9fzYl
Hewn1MnOrGdFuHdI6QJXzHnjOtK/4yRM+LHj7Iy7A0t3s8ycfr/jZOziSoQqbOW9ac/GFjnhGR2N
txg60LvoRyI0kp+xEfR+nRGrEGBqJtq/mLIS476j9t7veSp5WJfQs4ICr8pAlXlpf01Mw/yD7iPH
MJkvyy0h9NTOaDjQsuy5B473msjwfTW0rSFCg0/uQ/Yx1HZnqP41pUuakYpUMU5w4TrTH1QE7gtX
pOVn3MOkDCLmQND/k9cFQZNgzf2xZMxBip31pEMcxiurO0pvYZWHoqaDXxQNHqv+M9aNMc+UVfj/
kJbLpFHxYLLDXyVJnceep42g9bXc0fIpuTeDhG/0RyOdJMmd0Jh9ma9lgaQVpXbPY4sWKR3Nxa+P
bo90JCLiUD/KBJ2xV1DTy890kX6237gbUZezWrH++thkUK2Oy/O+wDSXhGQ0+VX4hEGI6EmdATX/
CQ8B+sJmHwjn7j+w263zk3jzTabj7q5YApFF8XlBYZMLHcDXnobJzjK0oqSEmOv3OFKzt/iAFoAA
FW/m6ebXGXalqrblZfkDTdOXm7VEs4Vc7Au72QjPIvMMgGrLk0fWJpmSKxl/PmGg9uTpyL66Xd9/
ULtdxjwysYB/LSX7SZYAyYgeEtmLp9DgJ1ZLFFwibyelCgdpML+FXOFg1MSfgX9oW30/NptThs4x
sGGjcpEFu9d7855+w0AkfHYvrZ/GQ6lCNoHZOeGyrEwLFVOVNYHLAM1ebxTSFglXRBlEPc3h/KB5
WaD86fV6vTIcgA1x4Q0PJZTw3LB6WHcB94CpSLup4ur7YKkPFdBbOKR9g6VJckVC0FFraXx7IcS8
u1uJHnIypffjHEjjNdZwOyKduDBzlbXUQR3/XwZVIbsKWmjJdWeM3Ra1iW54OxJo7PfOoCQXxTkG
Xq5hOJsaSTEbgahE2Rxg9taG79zJCsSd1SICAOkyIjj2LA7vcaiOMqK7SDba0qIa5JNkNhznrDBF
7+OLyg3DrlcN5NSAav09xtAQ9oAt8xGkFPYv92oK/0UoFP4QKiXP7dCKcDdNHx0HkQ/fZpLXflCd
KxfTKAgRuegn2pQP0nJQ9akHM4Ut4EJXR1xdiyBRW2ajXxOknZ6xwPtpSOAUdS5DpLe+pfPlErlM
hgRzFvUKapCxdHstR26hgMLLKW6SSzqlGVniA+nEgIlt7EUrlJ/U+VsJDfwc1FoO/80UZD8h0vEI
tvSAX9Ni9f73KsvFvlz36LqCiTyq+mHvWH8korANEGfmz5sebBSfGCvng+h+efY35PQDDcsmOFiB
v5EV8qo7nD2s/fqbuFDlVjfXjFxTTFMWrOZ3ONjHh1jNhD6uGR422JvoJ94K4hyO87BTUBrmLLRj
4Ln/G4uc+qN5lPoDaFckaU31emSWt76lJDeQuD9Q/0xDpCswfa6bswqnpoc9C6inzjl9w0bGlhDi
SL0RJah+sxlM7XoDPJC2+cKMW23nyzggAWIfIZurdc8vBojy3oDlaGHUNzU2WbrzSbjAouf+8vl/
MLQD40EE6jdN2RBU4bEGOgfSMeR041vGmmuJN73vanes7MnDz2EpQPR8VrYoPM9zcQxv84WzgBwP
2ap2I6WkrZCUV/aecHLIfak7LLiPm7Cou8UfipcYEPyk4y10L9XQxk9Avu5SlGK7YokCEJgLWzR+
+zBeNQGDvXjrOYwfiSVGoVWHstRDgiAYYq16tirXG2nhczug30edTPjV38czaciV5ZGSrSW2J3Lw
GMN3QzRe37aeMpjDfRNhzm+IK2U6pM9zgC/mwvXOVBdjFZYrli20Fple8MyoId8quIVEbNoKd7DC
5QSMgwzXbW6G+UnZLB1ivYKdESta4m06iiA6XDIfkvLIvvBWGj62eJEyzmpT/SmqjrywYNpo5EuF
s+FCFJNjQLX53jUglr47lv+Bb1+EfCTn25NaQn054n0AiWVe1AYZFOiQap9TGiIaIcMNBh51jEtf
Rto989vZHhz2gwl2OPDdmF76QJvqHyRrQmOS7T/mmtFFYqZimq+erGFonQeESKynSFTXwZOR+LHz
Ca/iqYikcDn83/StNbWKVsyH2ayGLGI3FWr4MANtkBt2VnpZ9o5v3LIlv2r9hr6yHlnrN9jRvm7e
g5JiB25rtIEYFoP6YP3AQs1HBWJZ4tRaVzbXKAquf6PfzXkX1foUrwxsQhBTgiMJSA74QP58dMNR
bst44SAnp86S8URkvHoJmcHLWxRjyt83Ndh3I7s+SjSFyliMSb3eH4Ua5JHdycK+Ps4ZWR7Bn59t
Yd1UE+4Tp//5uQqL9CXt1uP3bqSnr41tB2DouQsVzWBo0BZ8UW5HSMopUlhaFhYwurJnZxw8vCKh
vRbwa2PxarxaKkp4jqTYLh2x4x6EFqR0XybnNqGVP0OzEKEO2VciCQFMyubC4eS3En+fbNjh9W8s
uepmS1m7YQ5kd0xvvQyA/UW2ER1MDlEYfzL88lQCTrdr5bVB1NhamuKRBfzQ1ZQo7jLe9kU2wm6b
Zxjp+suqMCkg+qXtGn/AT/XcI8ArHSuT0c4dWUy5KipaZQIDpUxKvcsmDUc2ljqJHd6dZeVQaFoJ
adR/Sc7hqE5xAozCIkCD1WVz5EtDaVrz0Xmud+y9MUBPgHZ9Uw+G+MnYHARUMyiwQqo63gZsRahS
CKmoDAqCIfcdaBQ1jUdPPSMZx0F8O/Pt/fyU7i21l3SPFt0GQpROUoDsSyeWiypVuX16Nt+DTQ6k
GLNoicDQiuwBE/M6LaTBDODjiKlNt5o2mngE+S23gbQnxxKoFoMCbKtS2e/CJfy/f86PhdEd5on8
yi5SIz1H9B9eC5sqPtE7rU6ExWRhBhdXWHJBX6UAHjvtlE7cRMHYNYxecG6uKlAmqBMf6EEaHf+a
0KE8u84MRWuv4Y03y520JSdNalZ/FVL8H9SYHJVb6IrYhO4HRMlrdYOLKR+ttr/N9Aq34cugnXnk
GWpGMJNYTrn3CnHyq02fMoQAEFg94CxAD/26sD0f7kImXEs3ndpnesDyGPWm1S+5gcUzBk3xkIgx
Ega+a0LZj073EL2pcbVWIC8n+PIQmGYT/Bl9V30wEKoOg5LmdSweNtMl6Y+3s1uNAFR3qn/i2TX5
OUW+qNG3hY8t6y77PypiACbp2fsMf6W5mgnhAe+KCEc4ic5AFhX2Y9VTWbIJq4opeqj3PjeW7XMU
2T7pLyaumvRPVmm3k/boixc/nS8HP4se4jE9ubVCdyEfnBzT0iNDoekT7nfb8GMF0BI9AkfYz28S
lScpeGvPgxn+VODFH3EHCMPTFhM2EX+nqkGoTgrhxdCr50k19XRadCo+HHWWK8qrUUlPnzLmt4J0
mP+XgqdIi19ARVzID+pdcCqVx02W4lt9LQkvXZbS5SAQNHyrkEEap9QaCLHMPfDX3Cv3qhJ4aPFn
bwY0f8RBrbCg9smF5wehkebaSqUC3a3MyQ1ihlqIHCxmEdOPgilyPYkRBAbM7mnwTVCVZ8nZ6yLX
karJVVBy5FwnrNuzsPKsmioyVR6O1oET83y6h5Wm8Gn9yL30PWb0ZckP41eoo0ITomIVJyScoCEC
L2ya8ygcTHHCvneYssUqs79Udx8LhrlrHVAUUmnOruxHN0C79SrF81GL7AU8Dq+0fqNYqGSB2fDh
kO1ApkD1F6VWB2VpOd9OZP2c2q571lOzoNEZMiE5gr+hAqSgywI1eAWN4hnNBPVmHvKk+gR9oHj1
x8CSzNeU1Gho2zLtJfI3H3thH+DR2tuj9b1dvKQ8Xc5vjeKi6196vut+Ecz5wKFaKudHJCXzx0XH
lrew4AzpU3UIN49tzz6f1MYNOzRq1Ag/qD0GEw+Hck61a494+BYFc48xPuPXzFVagxSb1U2HOH/B
f0k2YUYPWxvxFtvh5YCfa0eA7Voz1K+viz6JxhtnkCJZ03qSBN64i3gHcDl7kROey9mdfQb51yM6
r9PxCDEr4pUtnUJi6oTh2OQA0c0XLoNyV1vaaNyFxBO9ORQ/RrFUXjndk1aSfSFl+JfQHIQ4OEjb
CpfxkQde4cb1t4PwUAhiVxMjupEg5pZQ3A/BLvXH71qAhtZ2eAyJFpl4hApU418h79YuFLL0KzxZ
647ajBzAAZBUNWDkBT+q2bChgH3oR+o3tnQGM4qcSAtUhntLrCnJVGQqCoarf0odifsklaLVeajQ
gdXF3Eoj1OVcw7uwcz3uXKnLiLmmmRWtZQAW+/4b52mGIGjHRMWtJd8LY9cdh8nVE8kogCIWYI2X
9nBuH45ZH4iARUUQMQ8XWGRt9hdAa0xMeOce80GYYjsUcQr15yqGqyfH2d6YVvBT/PUDY+36kdNP
TUmXH/AicOPx3FJPGyoJYHNGs4vbMXW3nr/Oi53BbXME6peXG3LfjfcUsub8d3eJDG1oUwX4P9wh
RCCiQu3nP9iU2+pVpbhnWAZlhVmnmF2Y0pVAPnx+wkNH4CKbhaxzAwYBWC9Ji4A3ET2pNIEOsu0Y
0xsGavOet92sa9Cy4TFTo26vdfM9vUNtSv38W5B/32HmNLIStmmQ3TNUwynQIxg+eiCJczfS/HOL
DZA/546CcnpgEa8Tj8lFy5HqfRJKZPnWb4+gZZZ+lesRlc3kU2OW9XBgTO85mEIBTIhjjaSZt8fk
nPKTRDTnuvZuF+iZm8ZSsdRmSIGprSvhYpjYhxDxPkiEPH5XlSpObSCS9EMSk7j/JeTQAuwQvKvg
v8cAaKWGS8IwUlwzqOhiY7kVXSFi0dYWo3eBN1JjcbjTV1Hh9Hm0FxH4AbFtPyU/QefDa/ysvvpG
FElhOZOxQ+yitrqvjFztkVYDTCc1sy11lczNxgF04EKT9vdYxgR+QIsI/uJ7pSeT+UbnUJRSl/5g
EZ5fJKF/P/ZNRXWAOiJEAoQVpVNaepuTGf/WFci+E3B0nLRep+6yCl74Qn6lf1JKQI0LtWb0Y4H1
h/ACYuD5OJmloKRi7FT40jazDCU9CLl8creUfgknyUwvLFfDWjbgMdO0NVrHezHMEal8KCJ1KDHX
H2htXI27i+EImF/sls2UpdC2RJF3i9awp0fXAAW3Cnwa0afPC53liMZm+qiCnupzpvQ1i6apXnIn
tVfRLIchIuWXPaOF5KrcUh2cmORx+xAF9B1QvyOH6UBlGR6zocw62tSvHEd7HvAMuj3jXd/sq/ny
HOwVsbwAQvIL8sAWKHD6neoyP+aNT0J+b6q9vZg9WOCL2WObFEO/gnFpG/x13sXzZoUlqbTKNjyd
YYeHeeIFPpCHucajOlkkhjKKicTwZgBB8bpz2aoX7oI6CJxN+jChmx+gkQJjLtRmd2/aHdgJ2BXG
syjV2NRO30ejHSPKw2JiFhINWrMamQQDF3g0jx3NBexnDiC0NLNtxY3TRDSQjBTRC50s1oaPDL+/
qtH9blqjumhH4e6L1JlTV15dqHmgQunk5k7SHOWB1HgZH0c1HTkvQjQgLJ81A+g3HPOUZSU+0N76
EGjSNFkv7puMTMctMpymLTrY+dvcrI8qz0mzgvyWhPVxOrjYt4cYWyQjU8e2aUpD3171mBKV785F
iH8LpVpu4eEH8RHVHCXiIl6u9AIQMLLORx3H6Y896iXU1joBkzZ2Arvq5f3QmFp+kIZ8458KX3kK
Y9oFNDWzATT9vFNwFXk5Bo4SxzdhKCgS1mHx2stzIg8T99gCh77Jka8wscL3N1H3GTV2ay3lHwUX
c0VYSQLaBm8RIIze0JToLOrF1fWAlwxTmNl1+ep5Kk8AL7wyW/BMpUIEu00PVXDgycV1MpnqjSEI
gkzS2zJ8wCCBaVP8IFzpaYVRqWDENqfF7W5gC+9thyWcq1xsq73RTlukv1b4zMkW+03LnrUuQMOh
DZWHyYBt0UXVu+R6YjVqBfCqDrwCFGacSlQTrpvro3ZjrF+YwLkqtx5pDgE1OMNgZpbE2nbqjllj
oNXr98aHrfvhkF0nBsdPq+8rhXIOqShFE1+baBThTnGZxyuIVy9/REQRY8dKD6C+gJEFoH/uDOjr
tAFya0NQxT+VEN8aSKjbXJq69tECQaWCbtUzilFnFzEnnCxX/D36dEwjDJhoCvK11mN6Ze6oddIm
EsDcd3eVZi6lZ8+2Yh732LqFQk/jREW7Yj6qdNx5NPWNYLDnGwQOpU7CpwrDl7FB9PnI6Uc6ZReb
wtjQMWORsnYbkif+n7bg4Lqu2H7Is3kAQYm7o5/I58XH65JU5eOFh4YAHjrxCxhPR2vortc6QNdb
UfrtUeIuRokWQoMXilF6aKGQdRVlLqzLzYuoluQSo9srcpr/9e2A+tyB6CjFQgiyzzFfjHDUixtA
PzETjOE5gB2m9mPNaAIpLy4O9Ar5t5+UpaqtLX+d6TPlAzdnaFK4/B3gDR98RsyMVTuMjS+bP+Vq
V590xwKaqxAvmJuNFMrDkNjWZTl7uvA35EE1UjlvAgloU1VLpszIggtIZEgMjQLiZCyRFX/u4bUJ
n76Ix3vZ1Kin6GylO4gGgfLRN57pMuTabRwOaWWU0A5V7QHKTqq5hq9Oz1JWaFlZ6ustuTYshR4e
WTIcxfE9HInakNI4mfqYRqXORRKViQwcilarfV1z/P99x3DBygntBsDb3crUli6vVLJWSbK6VozC
iJAHcU9bnGOzsg6+RroNpBU5/sTCr/EGK449mOfk+DR+6KOMlzHxorHCVd4gInOw0Z3hlhuSenXc
gNI91+wp0y0b4Qyg3iW5elI4fdWB2MB4rhLVyRDhud3/0lNgxFsggUKl987Ut3cbMqrTrYZLASI6
NotELNcLcUwIUR41R0LCL1doiAp/+4yJAwb9GUwj8rugAR5OufNQI+PIVcojVESrfFLwnEg1xbeZ
GLJEfaFlDGWUNr/g22DYMPYjS8frWiH1+voj724s3Hy9zGsKRaCIF0JNvHp8UsU1RM7jHhg0AcfE
pr7rc6+3YU4/lJxWkWhlJ6uay2VoqDd1KSNC2CHUr+eO9tONJ583rrvRLhfiPmxhr4ja2pkeLJ9d
tPkicqe4HrQlma6LqaQPCyAKrKlybeA6xDS+IFUgpvWdr5VR3sDEBsELPoWjD8e/ZWIpstHYRZt6
25Xbz+DHqQy01ddryrh6B5oOQpgh7jRW+fKHtq787OJweebtwVeooQCyKZ5DDs678mcT8fFoUiU/
HLLMjhZf4ogy5eur+7NjjEt/v3UEOcS3NWCVEAI7B2PhXl08oIXn412ByAQkLFAegnJyi71uQde2
E939tDohXXVfUeH/537CjWrm6XRTgGOmfWU2u30uKrQ1r3OC6PYyystXj9ofPeAZJVoacbMo7aHc
NpQVNxAoQ7QO42qoJzWxuAonCQsqts88gAxLk/Ef9o2KgDrdYfovhLgHhnHAc+fGPun8Be8PYg61
uqjlqDhnw0v/SXKjJham5SVkh34PMRbwR7hVPbHEjyh+M33+SVgQOIPLIwm8SUL0dB0UQC1PRsHF
TiCSgMwbvABCYRahF3hKWs+366hJHatahprBELHHJ3SgX8FB1BCBqO+oBtBAGRnYzgnRizNP3+9S
Z9bcjIbOZUhJTPUBGEkbgbF7fh25Pdfc+N5RWZGjqcd9m3i8FZwhIlu4c0oAc5azKePxP9+YS/ti
iH20TJG++8HDheYfXXte3RolgQPaSeWkDORDK1k8P6JYpLcpVsZi5OPw3kitKNgkQLSO9sUQjLIc
zUm1c7KZ3mhfdYEcIQNjO2BnVX02pRpiKwMdHrlWLUt12UXJer+4+Ed+gUsoHf/4U1GgoRx9/RXH
kjTZTHykjFylSDhGP/OkZeQOzw9ZptAsK4siIrJng+7jVDPXYfmOntGCmrAK8G+Ki4Zb4f2nNmWL
o4Pp5hcAUfJqinRHLZ6sm3faZEZZIc9cXIbAfVmIkafmovX3vqqnzCJuqxz9f5/mGLsRRBDGdl/h
9ZsLEJ9MhSw2CXR35oE+jh5eFWhYYjfhCbhIkdjq1VhSowwhhHirnrDMyzRBLC7spIlSg8zCAXq+
02n/27vLIPdS9SZq/2UDrS3OZLvbTvdbL8df6hPvUZhmgpiq+gqSv29FnoAKwarx8mQLxlh/SMoS
85mkr3NwFqunJiSpBFOf7yjGIghFAWRoTU86w5bpjYM0+3Q+c+jZOgOfU8TceBwsQNxgjLNdNLc9
a0bQQTtQUAQuhPO/pRn/OVw9LYgLlDolZ4geaeT/ug17lgOPZ2JO31vDAmuUfOQkKrpoBGUi4RAz
59HaNF9KD6G/tbsP5mU11wTvJwkzsDq6zUsByopg+fCofKXFPpHoAdX02y9xv5qnKuP69N+sS6S6
DBH0XFdppOkh5bdRn/WeI3BL+9cJ3SJbInQNL1KtZUQtdCwYeCna7yUdybnTL6jkJFATXXgPhNtN
dU2KeLGovC77+5To8hVHbLL/JaSmn3+oclB+Pw1yUprXWjWfGSJwXygt39IATtjrmX375pcHUKdy
G1AznUqfjncnQd7OKTq/BIQ5dvmKSzXZopObuQsgthP64Xu/MsYLoi8BPFfhWy+dtsXSgouKSsC1
Xaa1QDfJzA4M8kHrt4juSAiac+mlUbfSayQOH2IV9djJW+6Oj70uUqtPHRprbC+1hZuAg/Nne/7z
f8cub867P2ZJ0hydH1YvTDun5UlQ93+DwGUOBgLbnY67WXErHoW5t8LdfG4MEFCK17Dv650BRP2o
iR4c0vg24CghpmdO/mq2UIRY9FNg5rE5RRSar//8XsNq0SAT3y0k3wDljFWtCadpocpL0cnZOv+h
35tfcxOitdV2Rz2ZO9EiXj4RzND2hTzb77qTHkJVNXNVS93wCRu4Fm/1bLMqu2PnO1e5i43eEcJE
O8/7rcJSb3a5+oXDhLwWMw1IKwIEqyA5H2zQJaYU/y0mWvCkMK7ZSUDzAR6oA3g0mjh0YFZK89rA
zEEE2DlxEhDhJ0SFJM2vgbZ8UoUTU05jyISf2W3h1PcY7zAu44jtEYmhDw7t3F1eGAx4tnnVIcGa
ABdgF2epgZVM+RcGTfoKJYwz+sr3LLWbpkHMdnBfLLLwZvvAU4+2P94UkpnRj+s5iZ6I4N9qGsvO
2hXhsvjQcO/zO3B7hni7SaxquS25ltMLFdurxFFhFXddm0TKJMoFhity+ZUqCUjhwUGAaZcpE0kg
xI4IbhIMuJfexqt3sRiEj3aBmkCMNmX8lXYmZ4a7R9s5h7+P32XytfUc5iVtmyF0H7GgtoL5L5YS
0gCCBOyruqkjY8QZeNjimNmvrqpBkbr9pdaF3AZ2NPYeqHz+cQPDBe31ExKCDh+QxQs+elnbgzq5
DuNy1NmRbBbXcQghTWFlYhplaAzTvPmOyNupZX6hF5yDY9eui5COUoN0fwtcxarojKDhESKuTHZx
pwOt5m1nfs5UHeCxZBmGxaFFHF9O7k7nmmLu5SyR+lAImAgeGdFdUINBzlc6FO8lCEsyHI1RtFrS
T51ZP81ncw8ivokOiAIEfV0NiOAdQ108/UndTol/CcPtUjI8A+ZAZ+C9WTR7ZFoIM9ZpreLRzoSJ
oalOLm/57tIc6VhhMGXUozghBVIiV2rzz3Qv6h1YDUzepPb6BmjY7uFP6WtB9WdW1DLsmM7wSGt6
KmOnK2ziB/RE2/RfqF90xh6aJuo2sGHlPW2G16oecRVgoM57qldOJZWrOJ4ADkVUzlmIkjoUyCAO
ejE/QUPQZyYgxo7yZfrWJ3ppd6zPfgiVxPMcpCpA2nnQhufK1ySjndXX2V0ul3GVma1DbNcbTmOi
VWC95E0NX0U03bM9wBI/+JWU+qORDd+VSUIt7o92o0RsclDdlxTkgKmS7ckO/vObTZaBM4SpYKwa
mzxiWWVjN/e7cUVXT02ULVyg4Y485N4pCJ5F42flIlS4OCmsdInh4/iKU8GI9xNbDV8KmRnXMAxb
rmkV4rFiVLsalCuPdaMVDlpVn1OgzoL+TA3Y9BVLxhu492KMSri+zgLJHPkadvhENas7CD4+ji9J
u4GfCeXNPCkApTzsbherVpDeXWGsf17fOIB8S+9im8sYon/mtP+jPwGkuQwnd8sARWq/IpRm4UAo
mubdnWsng2vS/5AdOImeE7u+132i986c5Zkad/ZJdZBgEh6lu1mH4x95LWpDQH9W9LAprBu+Ullk
BAHuKkAja+1Ub/UGDoGCNg1xUhkMlZNESpfH3JzwDkrsiShfL1Kc9/2SlLkYNiGskUn4XxCUKXQn
Ma8kIB4pBeLcRZyoxnGppFVxWRfGVfRhQy5BuCe5+r3GMK4HJ1PqA5TXsV9MEbLO+tDCFC6Hr9Jj
yPuZdqPOGfIa8QkVVqi6IZ0Jyl0/zdkPCn/B6gbSmNJ8cyUIzsPYTY2uxGBZYYGf4itmTPFnd4SH
P+fzEFYk6WZe/+SzfPUF9sXJTP1gQoyEpHD2tOA+SfG36zXuHaUrLEIyN+ie0uS17KNIXD33jfYw
RBBRdQVtmw9HWEMRZFbfjX2Wq+JF/A/6SuPk8YT4N72wkjqgbij/7MmclOndUJHwGjIYdb5p05ov
IiTmonHGYF181s10xiT08FQwotgJIPMEjZl7L2A0Zp0LFk1vmjQgLHsJkNVOwODvEXEydWdhher/
6YBuDq51m7AZVC1Op9U1JxikSrPryda42QIfiHt2ODfwIJYa84F+N6H+gFKIGQrH3tFhDceFnqoM
alfh58zMVtdoYWzXRV9bNmdFX3x1fmdRMTFYf0/+q6SBvcB38zgBbb1aKU6udmIUlYNLtUl0I6Ff
Es6bM/Oo0dxwAAvvYcrVVtbyb/FDX9RQT0pkUjAgVXVlevHgqo0z1Z32H5cFcyFlX7nlbXdCi1Yq
CjPhFbdKDEBCZxs57sdlrjqShwydHUq9EUbSFgPW//t1Lw1P/wS0VzrA4CzDVs2Ew6+OxWgml5Jw
QnqhAX0SWAGQV65ibRsh8DAF2VhzxR4Y1qxlaqdkVMLAkXEUcsvwN7thYq6QpTy8fsV8yWbIXkzq
leIHyWLaii4fbJcxuvpoVXBRsFam3pnHkPQ9bowmpBLJmwToA7K9vAtGqgRl8WMe2ql8m/mgv9fO
hloV5Mud9yZUOrGnBwT4JMUw+zTmHn5TYvN8Xadko+CpQQwIKOrfAxHOMxNDoG1M8+s0bGqzn25z
9hr0gxDPNIEvyTkAs+qh5Ya5sjz0wlfNztrJDSDwwSzklbqQ6zWcO/ZzgxjPHrzWxjc9PeMTmi74
sLMegpVhaLHSUlc2HwpX9ri3/DvGBnCl8VC7fl7bzAN1GxHbQAx1AF6SovP3LfJCd512WNWOkn02
KH66qjKfKqfAiaB9wODMtQUSK+QnpHC3VeDWOQ51iVnnjZ/8dxufJbgeOIc2Vw18mTRZ85O8Gt78
dcJMYdIdeR8wNEInOmbGOeJDlqV9roF9cFYjMu8RlLqESoQ27nvxxksCrH/030PzEI9MI8NuNm2D
EXnTFdMJ1ICCVfhOOUCt4wyhxmo2mLBlUUtJ0wJI5MOrpUfxveC2FuKO/gW3ja6H7aWJJSFC6jzK
fhM+kTTjiksigU8MAcLGNNeHTG7vYJCSkD4MB98O4v0U4/39A0zmL/peKA+EKRi+h6R6OfPOVtgC
kM6liuEJ658lU0E0w1a5XG3q/BDeqOocIAzYwGlIjoCyKFp9UbOXMXymeh+2rI0iLx387rZlUuZI
3FTzfm7JqX51Ib9zW2stOtOXPmwDJNUZ5e2tD07fyQyoNp6qJLnN0HrUehFdznGIjDTu0q59FtvI
el0dwx9HWvTjdGc8CrJmGzR9lFawKlfKPGlqW+OTIwcgQ3Suqhq8mfc2DJPUuQUNmWzTpqN8qB3F
Bz4OHIIj9CglSHMkZ31pLRGTf9UEyWQlXIDpPSpZxmhzJsx2tIbqHGtN+I7Z3W/jWqj7934fkV0u
51BJ5KshhQe3kdLjCr4QMfwiKrApU8Taf7e7fGsBx+C27+UFXzQK7a3ZN1b+mpSx2TeI7O9RtU6O
NkohIpYDpmRsb8Qc1VCyx/+HzrNJUkccVEtMrjH1ZW5y30z+P6MmHReqcP/fttOUAlqQjkyqS3Ij
d2xR/dxfyRK6K7zYeqgJhJkN1Rouo273UKDL8WqmOBsA9oJrW2RIfJMsCbsg6hBDyLkrSg6kD01M
TPlhQCfdFeTMhIQZsRgpE3Ij9ES3EjlaxKv3ikimD+4d/pKof6ih6PcgVWLkA5jyQRa8Cp8dQNIj
Z0gcswialpXu2DuUDffrA5ba/nQoEqVsaren1x7QxqYMVIOnD0DFuuHba7fFNbFB2asXIS1l2tA6
7xQYuyOo5etFvAoyEgyNqzW+wZ3wgRhJ6hUGW0lYSe6JikHrj982Yqr4GTQrocAooGp3BIA9ZeIg
xpqnJ4zOHmKPap9JBL6xPQ9xB9mS03xX8eNV2L5yRh1Z71mG/1wTLHgBUCjJm5MBWnQ4YG5WQ7DX
dJhIh89ps5PYjULYToNsB9KvOVj6T8pGzryUcnc6AoCnN8UQjnMIGLj0SfnPWyTi3VLJ0/ga3YcT
Eq11Bk3w3qntANjodQvrABnrLTZxGiBFEfxLDt57xPLXdkV8rxVd/KqYPaEsr24AFdIAU5c1640o
KfUBtAN3YNrVuL2qWcoUe/XMQKaitA7OwHSivUSMd7PY5WNDDE4NxCdnIhLG5T2//I/6WIIrbo9v
LrXsUvfAPiK/MWzFVHdoJpwYSSdjeC8bBapxi+0DneCZiTe7wMgkT7PJFv+oHmbr3sYG1EC4o01h
r+N/6lPTdn/RYzqdUySFznNWO1IA7r7yKj+maLombzHeGryPWQVRvcAGRItVgcE5j82wwZtaALoz
cCKvPMMEBuqBcH1A+hHtVkIQsBIVXYa0TT+AsJLTDISXKkvaRPFfy2gjZsj0zpjU3BaBqgOHHCZr
T3UwlNzHlZD4mlAM5Nb3BR3930w8vny0BNrqa92VbTzQWnsICjBuCQv63NVlJ3rsLqD4TuQ8V5+6
JFbcQTS/5V7lMVEpBFNLcKSC8DBb2AP7EUEBs0uevvF5FHjwvqXdZ1JA+BFVAn6UqpBZeTrDENJX
dpslew8iOzu4QxkRjcPCOqK3DpNMp8LW/6/W3dRyOnCtzQFFf+yiPF82XYAesFeN/8Fed3QspE0n
6IJgKkJ1cOHtgUnZklV7HSyLSyUFWaLBc7Graiodq4FJc4/lEa5+ou3gSxikyzU2+qMrrp+UT5w2
MDwR+ojTJYF8jvQouE8Fb10MKOx9M1KvNnTuDwEykWLNTFyz5U1b5J67cwx0FF4X8kuh3KSgx7zi
i6sZGeCddwJ+DYkQGUTrz4VfpHoqQmHXf+jAUXA8eQMiIod+nmIXbb2B5u1GGgWUvYqcPlC/8r0X
I+A+LedXOTnGWs70lEDYOmsldDRudghXaPBQSWBYcpZwMEEac1iAoY7GCF/2Mt0MCgurs7QIiJlw
mihz1r1d/62md6cBzYgqgg5HqxJnBAxxg7ywwBmanyBw+JlI1HbSdtlkOt3mg2SQyy8tm6cYuS4N
Jh94QKE0LMjJCzMOGKJEAcP/VySv4dFJU2UcbY/ekJPfmh9Sm5zat/N4jX0FVLWS4UMsKSGNdX/F
h0PGRyC7KYHegtkuiiViFJSKJtvmwdEiZY4cj2ZKHl9kPtd0IruJEB3Y4cip+e1v7+CbG+ya3qNT
DRwa5Y1xqPdaLcl3b+W4OxuowisPhcyPGwAr/pwYxuaRQ915aR91d9nT0yqyCdnc5WLU2C5svwwS
UylVEGPUqRY8uqGhKbTd4AOAec7Gjl0x6SSjlAyy05JOS6rNI4CgCTHpa2fXAfR+jHmBpZZz6fe8
DjvLoWCiSYXO1R8BYIMnNR4VOinWCBZ0bj49biG92D9hKpNrH3MnxBgi63r3SbRlLhfbY9CRl2Jv
pVXPnHjO13Til0LUIYr/lTQb8LUlIy/Qv//kqwidVfL509oN/PovpwxntuI36YXdvje19Jk8H2aV
PFNfkJjmGq38JMO2ASUlo25SQBbJgCSY8FFiRsdXKNCBe6/cA+526gyzcc2kz+Eavx5cocbOpMCs
POVnMKw/SRFS4UWdvVg7zM+lnez9Hp3hHkXspaVyMLCe3wcqKWIV3pdv89w0Q7QbJQ6zMnbIedeR
OQaNzsavg46a5qSUp6Y/s/ucodHzVVJffP/L2Ah1IJjY7dlj/LdCRVk3UFEM+bezb8uUJQiyyJrb
CkaWJH9pGXflc8VNcd7OhsiVjQ6iBAv8QYqpQ41mZpiui8xkPTwmmWfy+dq0pSWD0K6xFesSxllZ
9jnScaC7z4oPz/MIGPLpmahzteLG26Fu3ADJ/OYaAqpprF+8rSImZfUYwVET64AkNeTOT0TSrA8w
YHowCnzCSCkfMzUAbdoWTYI+XrRETmFEUauMOgVE9ecEPinFBEP7tx59nRhLYhcqM706seV+pi9V
glkHz0Fw7yb7TQtpDb9AdPl5eH0l/Uyd9VCeCwalk7RNHUHBt/LR0S/6iWVTeqTT0pITyOIH4bdm
GkRIA50BI4cLIYMRRWRBzWvCJclX0x66i44TCZsWMVrF2NfTf1QstZI/AOPhckzkoQS72C4fPr9+
/zvZQjOe/fEKPP0lRn4rjfzAZkU+mGdSg4Xbp3ZGAEn14Qqw+7Sgr4eC6l2vNoD6QbpTZGBQwEc6
5JMavG8248h5X1SR0rYF0pP+/e/GF4Y3WlBtLKnKYIC5iy62/0I2vb7Jqlc+teKHDai3mNA40+ga
ZOTIXdyGnhN+l5QhqB+EuA+RSQic+FtiHPUq34pBSXn4J3R2m83WZ4q6oODPRjm71o+v319stATx
xIvxa2r5K8MzZpoE0u+cF+Y8uAiuDUUbSlzRgxTSOY5YMswWoinnJNoXTYHNqZbXDX6GEldJv0d/
/QIkcQSX7uHkyYLqpnP5zxajlo8CWo07OqfPFg47n9F+WofU3ROGK8XWmTF89d9C7gE/eVKK5eDI
O7ooVggiDCDMFN65LrIWVHSPo6g1kQEozRF98FU5+PbDp15UoQKPWa+IL5IKuJICA/vDABhQu8d/
Td40+SYfAzBDaJzbLyC8Db19L4hXzbKhq+QKdj/XCTDV6/+mCndJXRdK1dfgFxJtGj4pZ5JgTodz
aoq9yisFt9JfIsrWgSm4j/5HjvCoZvFA5R2FO3JUNQrjnOrGyNmzylyzFtB6kJke3doolS1iJbav
9oCg4OivbuZVwUh8BTu3sqv40lyKP/0X0rEaNsmA0zK8rffVOcJ8x+pdNsO+1MdQxBIvZzdf7k3/
LMO0V1pj3eO/q862o1aVNKxt4djuAVfB3qdyK+AlyEiRG6Qm+jeQMtirvIocLXjztnEG5VGiaIwl
hNbVsY4VyB2fT27OCcLfSDQjyQhyk9O1kBJzmEqmGmWQ+3fV1KChh7oh/W7B9Fw2UbTxViyYfjcx
fgrMY8dsQUEhMpcDPNeQ/s9ITXSamym5UN8Un2MVtBHLgXKbyz3MQzbvRwBkYkipLE+vtnZ4K+OB
QnS9n3nx+KEUy40SRTMRWs5wYqrn2LoPCaZm4ikfUY63N5sR7fzjxH+3/VbOiXjRF2B2DJVfrIV3
ss466cS19btSH2CHURkEX8Y2tVwJEIFcIo+/l6B0q1Af0IhtucLdHnikb4Xh/rYUxvVGUIpfxan2
E/XZKSuV4GjelVA8XSwBzRedbjxr2npv81aEfusOoaOyMVopFOhv49w833SeBl3LpvUHiXtByv8K
XOk6facc2+L5rWLUpkIN1wlKrMRPnY7bIpv5xBRomI7KYv88eBzQ3Id3lCUoJ2aNnDlRDGxiDW90
rw9nXeYB1Pz+3bbw5wRG0z6jnM3cxnl3YZgHZb44vyw3RJptTuipRBUp/lawwjWrDUgP7+3l0BIz
1Xj5qUDa5eG3SZlkLqLckHLgR2GphKstl2SOhLaF3px9pfp2E3uLxkeqbmxD6+RjQ98auTDJC9nP
MwtWARbib3pCphKeM2rV+RGYkA6Ukp9m2RBF1AnPq0SqQCw7hdQi9vPTiHMyzhEyoo4PRaoUGj6F
z66c4YVH/nWun50Pa1VqIpPR+VHNo995V3reyGN3/bAr8sP3WdzAjFuE0ZWrwodecBHOH5ib1Dz2
oFE5EH4vRil3q2xKAeXpKt+Lj84L5HmQP6jOnH5Ob1iBqP8YxDH/CBKbKAyo6bir1EM+G6MIhJmT
yCy9qSi4Ysf677mWas8eyNy17XE/iCUcOD0WVhmBKGv8dDs2sBOlae58Zd/YnvzibmvotD9otqhr
zn+YtvCGPbomEG9LhtUkKvXNoBZuzqXtzeEBnGgq11OhxrnR2Tz4UCfN3WN3T3N9GX+r2G0Ax87W
9A19U4scjefGko7Z01anKSFf+TqPKpzscUXov3QcKcu8Xa65Z+Oc3V1mFH4ZmuNtKxzckS+zrBZw
U6JBrl5vNzfOykWJftRxkuEfxtWq
`protect end_protected

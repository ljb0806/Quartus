��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�%qV|i:��r�1˲i���sd��P4x��y�����˂x��ۈ��ȷ���P�{�G�mp�T��Kz69�ע�q�l�p�ѡ��n�$�Z�H
M��q��@���	� ���
�����'��-��؀J��a&�ŭ}���Rpտ��Ġ�=�	5O ����5�h4gf&��tn͛��x�զ�wu����?ƴ���\��b��R�w�5;m��P��{�d�n��5N]7��S��t*P�Mۡ1� �[����G�AN$M���P�����O 4�5��08�'�7^�$B�r�;�e��e��H�4'�D)��e?��Z�H�j3��18A2��ti����ե�^l���v5��z�|�3��+�m�v'�:]?3��I<�$$0xnO�p��l&���M��^R�06��X�V�i�^�uwT���Y�N[T�f����]]V�B�4p4u�0F��2��!o��@\��WMy�t,��'IP��1�?�����h�T���J�L�v���1�ן���m����7�"��~�؊�\
/{%^9�ض���H#G(���-�1gs��ݵr]�����:C�XC�#ƀ�3^B��?CHW�%�r1��Y"p�ڞ\0��:G�!���_��`2��)ﴂ�c��&�nH)呹��Jpv��T>�ɹK����/���~�3"�%in�@�N�����\<�^q��h��t������M�о��}�� �K��|���%�9���
��)Z�s�����_4��	�c�Qo��yvv7�P`�#�$j$�Azv��3��&��Z�&kswe�i����V4�ߑ�P�������1@�쏫���=|1cG�q���#(7�M�I�p(Ǡ��s؋����w�L�ť���,OB8�<J�2#AT�W
4SLo��H�+����̲1SY�jUe�|0�5{�۩!��hI���b{���]�|�j�Ӭ�z$,3��NtQ��ʞ�#Ru��i��uHT)X2E@���ѥ�/�3���:%�� �,�J� �q8�vZ25f���ud~�}R�6Ņ�2���o�{���H����"�V�m����Y *�us{>�G������ 7�\�C�F0QZO5�s-�⡔���b*󋾣��h�h���\������."T]����|�h�7MA��D�Gkr���81� a���_�a�
[�a"�g�x��_Pn],MYզb�P#Y��S�cw�OyF�V��Ғ��莦�s��w�Ш��}ý�R���F䠯�P�o������#�f�[ �p��<7�g%�\4$����(��f�@u�]�}^��r��V�`�R)Jg={r���˘���Q~5B����9��Z;,��L����G��fϗ|m���k"m����7�$sb]��!J�޻8�a������f`�@ijy�TB�e"�1|�.�����}�܌�����F���vM��N�S
9x�H';7����o�(��}�nD��M�����1b�o�aLy���Ø%�vau�r7��a��ک p�����uM���+d��q���)i'�Tq�᳭��@ y.5��ۥ��V��,	�W��A�@|z�ʰ��He�/x������]3�	�D]��J�C��c2�%:g��ON6Y�;�<�+d��ⴉ�\�Ƹ�K��P���d틑��|�㷃\4V��2�,L�4ܔՆ�o��2��
���H��H��Z�ua��-�(�I�i�C��0�#$TȴA��3։ĝ=�DƁ�u����cq��u��p����'焱Gj�e�ת���?j��;JK�J?H��E�(�5�wo�(��e��x݂��!Y�~��xh~�V�|4ud�8Ƒߖ+� O5ܷQ����@�V-j8D�6F�������Έ<�Ie��k\��*V��p�U�hF��_T6�C���0�v/?=Z�Ѭ$_m�t7G��[��;!!����H?q�����&�<�Hk�4W�fsYǭ�̮4%��q��M���LNq,;���?�Q
c�yҼS)Xhv��W�O��O"�C.�v�"�Q-�g��zn3t�����ɷ瓲 �k�r�a���RZ����x�o�)���\�16�kq���W~m�R=����6t�\ar(��"6�j���;\��qΖ��qȺλ�D�n>S�x����LR�xg���VO����f�9�G��<�Z;+���)�߆�IM0Y�dΘПQp�� ��
i��5�J�ԭa����뇔��}C�m�g��%DǼ.��лM�c��L�z� �wξ����0�Tt�4�n@��O4w�y�i��B�NG��T�bR<T��������n&�~�W���?��/��Dmq��$j�4&Tgz׻�����W٠u�Ưw�����2�{�@���W�R\��N�a�F���	�;�,��8?.6D�`�Mt�+��!`�o1G^�
���F~ʜ&¶Q+�y��U��	�9�w���z?<��x�T�/w��wjT��
���5m�S��u���3��H3��N��L�P�=����8�I�	'�(��1�Ly9���#u�T�^�Hl��K�����6~�h�;�&ں�} ��"ȵ�j��/���"�Ľa�3ҿ�3���[6,h�4N@EOH��1��|JtԒ�u��YR%b� ��n0{}�f�y&�B�ρ�� ����б܈do�^�K�L��+�#���Z�%��`ǖY$v���;�7�|�l�?��:h��ӓ���A��kQ3�R��Uks�-^���unZ�ks-�7�q��h"��(�̮#�r� ���<�����o���z�ށ;�-�Px�r�
�=�Pc�&y{N��&�0��zL=;A'��l���]�:�`�_��y��"o�q�\��]�G<����V_l��pHKQul{jc�����{�Ô�>΅���+�y #QAK�g����p�U�yw� �n?�u:d@k��8�-�a&�_a|PO�d���I.1��_8����F�^Va��5y:ľL�V~��)+7�\�>`������#_�RY�u�6�Cwý�pvQ^��,�.W��Is.B��`���Yr�Y7 ���S�l��r�m�B�oF�jf"�&7�.G���l�B�B�Ժ���2Ĕ�mk�8���
�������U(䊼	�@GzSg/կ��>:�%j���;:�=�}1��>��$�="�B.]�N��K�b z>�� Dop�Ӹ>>��g��V�hty��艜t�Ër�/0k3�)h�C�?�������t���{��xi%�@�P�N\X���'	�&7lsc+�e��NDͣJp~�+�}�'��º��.C%��d��<��䒬}./��I�W�r��"R'ч�p4ۋ�(�W�A6�Y&2$��N[o�b��2� ����~�ը��`��%б�韨�F`��9@ �'�,�Q�+��BE��{ܒ����A�u�*��:�4�a&(|)�F�	�ͨD<[�e��!pƴ� ��.�D�I�
<v�N�RM�g�l��o���A�ՙ\��.B����J%.2�x�6>a��7ߤX� Qh���ͼ���Y� ii��a�x�O=��K��+�>>(r������w�R���ol^����s
2l��Ll����.�5c0��4�ۦW�Q1��w�֐�Q!�����YW������P^07�g���ڞ�
���X�R�l�ݒ>(��:j+���Sl?���q_̣�r�zeG.ƞ��$:�t'��hJ�OriR8�}y�7xmN��]~���}�����D#��|��q�U�,�/E5q�Jұ|�Q�&��@��ͱ���B%%��q.�5y~r�����O�)���qW)o�'-ھ�-�-����z�C䰾����pD"72e��/��ZR�@Q�31�##���ܳ�� �l[����� �|gP��>�G��b!ԁ��{� :+���?I��w���4��.��z|�;���,�H�Z��� ����ʷ��l���\������B�ڒV�V�X��h;W����2�[���X��p���Â�!�Z^� ��n��e����K�kx�w����t�V��� ���Q<����4����A�*�{(�?q�X8qԧ�08��z�:�.q{'��͞v�UN-,�e>1�Ŷ��|�����1��������k&ZZy��_B[��R���`���#���G%��	q��J��:����R�
�i��8{�۶��k��>�!n��@�0�ٯ��jJ��ݒ���`��i%79�z�~R��UN9�+����-�)�lP����SS"Xq"":��<l��hxw��̣��y��~�A������Q��|2֞	pL�ǔpX�����=M��8�SR�Z4h& �W�<�.�Kz#e306�W��1�h��۞
~�z��:7[=�W���h��dc4^�{8kQ��jb: �2?�T:�1X��ԁ�{�9M�F�7<ӝ���8�WU��Ͽ�[�Μe��I�[{힃�����S�꟪GU?����HUi#Tg��< D��b�E�EN��6�f��Mqe��n-����Ps ��p:a��WS��N����:,Q[��[��3,B<`���^&�{VIpS�o��]!�}"'G�}F=\�P5��{�l&�e�_3H���iJ�Ӿm)Uc� o�k���?_��v�#�=�,+�ɓ[A��$?ߎ3-��,l�4��s�^�ML�)��<�oº��xv��^�1A$��X��+.��N�QQ-��@�%1�J�����m6�ߩ=kl�/�y�`.��cz��� �%%v#5�ɡ�:��u��D����^�l{Q��9+�K���0/�"&����SRo�+������ ;�Q����(���< ���D���R^G��2�3v�ބ�'c�>��)�$9\	�����v1-M��[~5M�f��G�q����2�iP���23������k=��$����4��p��[W�:G���
ى{6�)i��Gj����= Bb���Y�1�m��h���,��|���|{N�@�Ev#[�RV���lQ�p=�]���p�G��2�
�g��{ZG;��N�	#E�B,
d�@R���lw������Z�B$vp��je�m��֨��|�(Ҳ沶w���ɑ9hք��v��O�{ �o�L���"�3g]њ��Tp��~G0�Z�ή�)�v� MA�i?kY>���@h�d�M�3f����>T�^ ��wÎ�P��C8����e�(G0�?��a4��	����<eY�{/,�WF�G$�@ݓ䴝8�IDUx���%iP�6۾L�|*��.�-�8}���OU��d�tg�������5c���;o��"�3jM�0ڒJS�;$�LENTX�����(�F;}��rH���5V��
�b��*�3�m\���h�A>�C 
Z��i�GזX�?����!LMN�<YN��ׂζ�ߝx�9/4�M���T|��Q\">�͙���:�'�^���}5�.�l"� � �Ӂ�V�@���O�~ ��IK��|ؤ�^µ�y�+���N���}��<�XMl(�|:�4��:nr&)ٷe�*�^�_�w	�r�?	L#@�
��Ѹ���c�h����`�W)Q�e����hZ=d7JsrT� �r��>M3:����S���El&�7 ��Z�v��{����:�z��a�V�r|�(���|���QA����ߝ����6i!�����E�M��F|l�ݘ��Y�O���Z!�Ҡ?�po4u����: u��R5���ZUdR�j�����O�7e}$��&w���x�n��~r"6p�_Y�^��5C�Oq�
j�lW�{�A���X�r}�I+���.�L�
�EjNE���#c��%�-V���R��䙪�?�'���P��U'/O����3�����M�p"�DD�w�[CZN�����U�x�������߁_F�9��@Htsv?_a˛;=�o����E$|���X8C���E�C�kl��.�y��V��}���1X���8?�ȴ1)���Y�n�|�D��x�ĀWQ��I2���Ji49^�p'@�8�g���~P��s��&�u �>m/s:6��Y��9`9_����������@#����1���@S�o�Kg�:~^�gh�/����LTx�Nb_��!Y���O}�T�Plz�l��g� @��)=[�����Ĝ*�i���"�Nc��>Җ 3|Ƕ>��lĢ���l��>3�\�r�mV��̨q���mw�bDB�7W�"`6nK���s����y|�t>��%3岒J�b�����^����Ҵ�(C�3̈́���̐ R��9e_Z0���iǜ��o53�%�;��|ʘ�z�6�r��ٱ�*E7{Zl��	�B�8�5pU�l����?ٹ��`�+���d��V��������}�6����n3w���G�1Nk.��˛�M����)�b��Q�d��N��j�7!���=��hbb��]�Pc�jl�+�pc6l�-�n���!��߯o
�s�D�v��u6Ze/��SFF�0�40Ջ��f�����+���j�;$��J����ծŽ37�]�r
�H��Ծ�CM��y�����~֓��G��b��P����D�K��S�� m��c6O��k����lކ{7�2�c�4�qD�7R��m�fo�`�Q������w�����x�"TX^�r4�yN�c�a�u�7 �I17]bV�A5��R�n��C$���oCRQ�=�RQ��u��3s�9��½�yЃ9( cn����w�5��jIg:�Ԝ�ͦ������"� ^%�������XF��ܟQ�En��{y(^��,��M!�$�T�@<�S7Ϯ��_�L�pSa��m%߶�~��#BAe��K4��z�Im�b�ǀ���b�5���lX��s����B�!#�����/EL�g��8gbnM6"Pb�49K���ϧ��<s}��9*`�Z㺪�Yx�_e�܇�)���_��Q�t�wJS�J�����N�[g�B�ʤ��t�9ӱ��5��ƫ���T^=�˜)�W�k� �'���th��A.v���I�k�#����G��9�8M��BI[2[%$e�y�ay��1g�Y����ޫ��dgukS�q����g�����}c
2#Ʀ�f�~���(�y�W��	�8jj:]lq^�f^���s�z�� ��d?��$��p��-T0�M�O�?E���D�B�k��NXlž��B��;u�/�U�*)q5���m@�>��#�X����-���;uh{�?d��([O�= �0s'��G^�c��������h��s��n�1�Qg�KB��;���M:躓����d�Q��8/ݘ!b����	��������gα��#ޤ���'2 ��#��U����is�jt��$&M!�t�'�>P�r�|�/�t�: �M�r;�����N�Ϛ��E�y�߭�$���8��i_�|"���tL�s���n{@q���m�b7�`�q-���;��Y�`ay�`�AH
����d㏲3�yU��˾�$�:~�sx�WuZY\�Z��ge�kBn���F֚0�^o�����F|�"?*�Y��@�����6K@�������Цիvn��KG4����V
�4Q�X��nz.hxb�e_�E�w!���x���e�B��Dj��~jR�̟��ᔉ�#�7맫I��:�\��|��2E��wW�B�4=��%)J��^Kv;g7١�h����d٘�'�\4�n�PZ�C��Cv����U(V�3ӱ$Ͻ� �B����25�rl\y��*b>৷\4o>����� dA�Y�q���%�o&���q�ŝ���<�Q�OGmؗ��<���ƴE��m��+��5���M���[�~���c��{U���FKa\gd�
HG��}�맑�ߖE�G�d�2��������F�v�C#2���'�JMJ��Sqt�$�Z����4��q�����}q�����`
Ћ�ֲ:��� L˧�<�BxJ�F�c���x8�=w�k1�ӕr��H�}n(��v"c�{PfP|�o� � �!�*=?��"EZ:C���ЮxZ�ˋi�w�ɪs�r^u�c� �VM�Ϥ*
;M���`C��u;�<+	�&l���&�_����������׻��ҕ�l�[.��*���N�#��b(�j
����+��V�8�[�v�*��(�Z��fn�.�,�٫s)�,(Xy'3�Ux�%4׮�B�`J���Γ�<B:�3��7Jk�-K�=5<���I=S�C �������dt)�W~}5QE8/��dZ)�)�L�s岻p.��� �w�0A0��Ad{�Gi��9�W�Y��s\�c=a@�4�2�\���9\��ϭ �6���P���K�P��^�H
q���1�����bi�"/Iԭ��=�n׉�T�u����0�{� U2�Z�����/�'�d��W>�`����G�d'!�W�v�O��:��p�v��#�;�#��Gk��8���'�nj��:�پ�|�|�IB���;����| ;4XbhHp%g���ʗ� E,͝b~m�jq�b��H]�(�lԍz�;����uT}f���"����7c?��&����^C%.�t$��B(&�����E`�0��v�:��]{��NFV�Y@j���f���_]��=h���Һ�4��ۚ�C���:5��w{\�b�+�c.���}�����X�{gDysa�q���ϝ�搋�
L��=���t���_��M��,REk�Ɂ�ye22�g�'��g�;F�I����?<6G�n���^�jܱU:h�t�f�>*��2�-��5��d�+E@�]M�ʯ��ܶ�>��n[�< �;`�Ml^��zֆ���V<���"uNȦ2щ���XH�u��#E l)D���)��^D� Բʹa�Q�^t�JqS7�-��\h�Kc��H�7�s�g|V�������\K_�lc��e-��Iɠ��������~ɂz��NvP&=0LǶ�DA�6��eA�����O��K�o�m���KH|BN�t́��
J��p@�	&_� �_�̙1�+K���}���+���s�#J�MuS�b��+ʪ����wy��A�����P�)��������7�^�J��QΕݱ�w�����*��Ui꾯-gjW(��������o&���ŊG%�#L��j��A�w�:��6��儴"~��Ǜ1(�-��Ma��#(�I�/�BG�x��H�P
=[��V|d��p߃ʝ k_y�e�ė�^�o��.�>)_�ҧ#�������l��,�m�e��2֏S�9!�(���l
eS��' � ���u8�mڻ�p r�E���f�w�<y�s����;8�������ؾ����m��r�Ě���p���9D�F�̌E��ŸE5v��C*�x�8�� .��S��7S�q�3F���#��`4�6�~�� T{Z��j�
]N���Ûkȟ7��Y��>���T}6�����JդWW�|V�<l@R�NG/1$�Z6>us�x��2��( ��)�jm)��sT�:aB ܿy2�s��!�=j�ũ�@"���gk�n���3��չ
��},y?��} P�9���Te��Dn`��S��ug�WoҸ�{j�Y;�z�h����j��/�&򼜭F��y��D^&c+"�cg���Vr'��|t�rC�,��(R)欁8���@:� �FR�
��q6��N�Nz��x�B��g�C��g�]�<?�B�^F�B�;܇��హ�Xs�K�>7T`J��ġH�	��,���B�r}t�#S~�?���&��4��}j�k��q������0�g'3'�B�S���֏�܂{�"p@�B2섉h�i�PpQc9����뤥��s¤Û����~�v��~��}��x��;u��M��~_~����"l�U�m���8�.���2�.A��c��m'��!�wOaQ�թk"�_�keӚ�2Y7
"�R2�{�����:ƕ@D����o�a�{m�
X�0�8�� ,�&V�Ë�:�l䈀�=�t��KS�Q���-:":��}���:rnm�'M�S� ������Ą*|޼(��$ֲr���Ƨm��D;�~X���i$�y�5��84�����{�z�-\[�	&�Q��������9G~
����}��3���`ѭ�Y+��s�U�]R��c@�2!9�21V�\�ĐT�3��~#Y��9�y�k[2�'��y^����M�|=[�j��s���`���a Bl��V/�|��.c��Fz��'$�Ԟlם��w�_@衫��j��|����w«��bZ0R1[JZ|*�����*� 	q��_����������*�^_D�¦��&���b?��	=�2kE�Q�A�oQP��^_�+�ћCfm4�(I��ǥg�dz0�1���Y�H3{	�K�-�Y�(Jv�=]���t�$p�&=t+g��JS�dMH]��:��5`������9�m�  ����5�=����H[�\�_R�6��y�(�}�K��� �*#/HF/�6c�$ʃ��e�ƵV���a�U�2�o���ME��8��d)��`���>���:���v�5���"��)zz� 15L�s��M�n-$��HfBO����ـ��EC�Uo���6 ��幬y����q������:Q����'޺����s��0܄~O4v�����������O�H���a���05����du3��T�Ϋ�=**Z��o��7* ��Yh�Vl�q:Z5l��<��.;����R�Fa��L��>�8=�_��#6!p�9�q�4}����@G�q<��-�TR��)!�d �ߏ%��TM���x� �Zc$�[W��y���"Z��������ީ���V��Rv�>�]Ip+]����?��Xc�򢁝"��׮Ȧs1H� ^�V�\�_Ckuu��.?ľ���i[u��!�0P�����*�,V����!��a.u��9�P�O&S�8-���\حCB����G�I�5�O�����̺�/0��^��g{_cvL_�����BJ��l�ﰘZL��?eY�Z��V�]�/'�>
j�h&�2�T��ծ�]S�yh5� :��î����릐���XBul�Gs}m�st)�/ M�$�Q�r+��6��Yafҳ`w?~�<{"�h�ɝ�2���7h��(j#(�'N\��,���@h�L�r��BE*b�is��Q��?��n��ro '��G3�>���ԓ��cqJ���g"��i��ť�q�²�xI�A�i�G?����O�2���5 !�
�V���qKZ�M\�T	p��\.�&�������[�����ei��Rh׵�{� *4��5�E�G��=��>����9��-2�)*\�g7�-y�����0=?�H<��;��8�$4���N�FQ+5�re����*�wA��*�*YL�f�R�W%{�$��l�������5]�3m�Ph�p:A߳L3d��S�r�KF�?d2�g�t9Ċ���)�QN�&�q#����:*a�gN;���M�p��|�d01����S� ��?�.���yT�
x����^9��}��!���8� ����Rq�b� �OhW)�#g�ş�uO?�l;�Tt�j�u�5�����A��S����~:T
K�c�	�Żp�����LpK�Q�4���ǜ�Di.Ne9}R�׶���o��G�/�x3P½�E�s�8E�-'OG� 4�O�V���xX�p�C��	5�����2V�Jj����	��h��N�)4r�n�R{�$'h��me�C�0��8���#k 0��Кi9��-F�ϴ�T�f��%�_N_-���Y��� /�rr�!^�S��R�ܬp�BTL덢f?
��Wԁ���h��=E�x�P:���B��o����v#e
�9dN�~���f�yD�|#Vv���9��~ē�	�K�.������޳��w׻v��|R�o&PMe���Z� /�TF_��D�'�<���"7C��o������Ã޺�S��l7�Ѱ,��9x$��, O�f��a�&i}p,!8
@��0Y�V����?�nH�[�(�2x���Q�t0�ʌF�zy�!'C�ekt���.˲��:�B�!��h�į��_�W�ѻ��ʍ?���r,������2�������v�-})�.�"]�8�+F8{4v��F��L��(���	,;e/�j����.�T�`ip�;RZL	�����T���vO"�"��U)B.��� ��a�H6A���H�}|M¶���Z����yN��h�4�y���m�1�>;�aW���������e���7Ͽ�p�an��{��_k�=<�w
P%1�2��L�ox��z]�R&��9��(q�s9�1B��ZF�̌�;�=U��L�K􇋙���:k����e5KC<!e���UH����LN�7R	|ĕcڟ����£�1�u�0��Jo�/Fc�����9WQ ԍ���J�a���D2��+�8���@�D?U-!���`sgr:Ҫ�4s�C�����X�8�i����f����m�'�%��o�ٮSS�Jd����w��m���Y��i�]גq�),H���GA�[;�s�L�ʰ*L��.�%��ٹ�.j�b���A��A����l�j��mX�{A��+c[w� m�6/��ً(�R�.k���+QdkR$>z|f�O=��sc����S;�-���||5��F��4����j���Į�UrM�_����ͣ���$�F{` ��0N5��2P���i��ׁ�+�� p���yPd�q�#����􀬌X��q}�9��s�ߡ��7j��)�K̜�J�����)i�P�4��z$M9�(����:�����3gJ'[-Y�Tp��N��r	11�ߞ��j�r�L�m��@��M�_?ݣ�Ɉ��
K8] Ph%r��Pn*/`H*v��:�@��q~ �J�ԥ֙"M��B1kLH�D�9��/U� k�训Ϛ}Y|��_�d��c�*x]�ہ_�;_Ӽ]�q�d�U���˼���tS�������j���F )�`�����$��dG���@����ѓ=��'$a�4ʦ�4!�;�~a�e�}x�Mc�#��*�I- hR�uXzf�O���莅�
��R�2y�sސ�B���mL��~]=���X�����'vc8c�qw��gL]x�?���3q�8>Q�a�!X��Q塧0m]۔�������d�����D��((�`��` Z���I�\�Gog��$�������&�!�֑�p��@��^z��>�ȥ�ȼH�h�8�
�j����ѓ���0��Ny%,���c�<�� ���҅����H�2,��WY�d�������y���{tqq� �<��$��s\��x�5�N1ٜ��tՐ�)ԇɇ�~hY��WOv�
�b�&����0�F���4
O*�=���:�w���1����~;��fV��B�M�@�^���
bo+UjDfzQ���M�������(�,��2Dw�tZ��~rY�V"n�\������t�	�2���_ ��"��a�J�\�)dGnz�Ia����]ك�O��zRD�]�C�v�}����05�,u�.�kM>�&�r,>i3e��]5���\IxT��n��
^�E�x��ߔ?��O����Xu��ޕ�EԺ������e��3J!��X�^������?m8W6v�ǥ��gג�
4�����z!�S]m
P��,�S�T��:���f�{=�V�i{�1RN��lg�"�Ŏ:8J��<B�b��0�5���Q���e�$${��M�ߥ.U�U�x���S��6�SN���s����GP��-�/�N�9��ƀ���*}���;G�����|fAs����T��\�W�$J�9��Q�ri������<���gw��5��6Z�^��aS1�$98@(Ŭms�}wc�h �'�mw�0��?8��i��5��n��N��Ѿ>������?����~���ϢiY�dM�-ɓ��=a�b��)
���9���V^Ad�Dd����`p�fXFM�?�"� �Gu,q�1�gY���'��Ě~K�E��|��et���<0$�-�K�
�qƵ�X��K�ܺ:�I�/}ֶ9ȱ�5�`�Y��v�4��X����,�`�o���8Jw��P���I�l�ޥ$ݗ��6_eޘ�31q#�J}W�#ê�ern�j9R*���S �Y�Y�H���o5tyօ��:\
�i�,7�-�(����:̥��sR��$�@�cF4�9d�1\��j��B6���/E��n8�%�<����Ⱦ`�0�*3�o��^UsٟnWO}�B<�6I�灌���������a����M��;���������˫����ε�0��2i�a �<j������������u��buo���^D�y+�p.#�ȑ��}�J�*��=<�2j���U�%��l��&@`������T`�*�<�bPd��RM�3�����ݽ��3z����l��yG�(�dyI��)���r��O)Q�n.��B�d�����{��.���(�猪$�؟�&�T�n*f6~pbs<b��~�����CU����y5�7��ʫc�Ek�`r��莬9NV�@�Y��B3�إsڽ��˷d��v H I�!KX7�;�!�3���1���zEuq:���Xpzq]������t�u�	S�%dw���@���<� �3	w�{A�s�+�i�ePq������X���p�Ś\�Lԟy��y�%N�t"i�"�-��'2�d��+�!��^$�Lxf��Շh��Z�~4N,�g��8��0��C�P�I�����)�]]��Ŀϧ��y�خ�(��DcI�әV�Uj��|J�_3&��K�Ni�A}@�䩠���H�������
�M����͈rd�I�OqI_�:�4�F"'�<b�Ϸ����S�sJ�(체��j��_��Y�o�"�C���x���P��o%H���wܺ�:���6�ˉ|����l��L�������Ehg`�"�f��חT������D|��y����CLs@1*e�U�R�v�|>�2E��루Go��L	qSد:���Ō+�]W�-�'��s�fi�r�1h�p�p���Y_+�R��==f
���=T�a�r^�*�,�y�mv�M���V��N"n�Fo0�8���v��0��+��]0�!c&�8~�0���Zb^�y�q����`ò����y��`VJW.�ǲ��»�|���V�~�'�E��f���j���m�E����Km+/�t����hYWirO��* y�x<r�-�/7�G&=�E���{����I7M����	�oX���&��&��:�����ه��5}G�8Mm�w#���rǣ�@�P�vO�B�p1q6����ҙ����(�o9�Y�F��Y�ق2eA+��A;�b�wEy���)~w����gL_���])�Kr���\�B	A.���F��2�Eo.'G����������_��>��v��	�(�|��H�E���T���#�}�إ�.�:"8�r�VT{V�Z�
DT{A����9a ^��*��Pc�"�;��m�Ϊ <�<H�����V[���XV��֥F��M�mo��i�Ϻ�{�e��ve���Z�!�߬��#y�g�B��~g�{im���	�v!X`��q2*������1�T��a7�z���:c�'|.no��|���|9���viD�a.�A#��;�6#��	x!��:f,�N�ݷ\�*@!�h�ؕN+�l�o��51�{���W��%�0�7.>E��0H'�����؍����tt����S��x3��/%%6 5�Y�:�yEŖ.�§/����Ν�e2���Ԧ����,D՝�秄��6-<n�4��d0����Kli0�䄪e�Z���I���$qb�Q�&d����p�s����P9kW]��"�d���;�M8�塉�δ�Ϥ/�`�F�����c�h� BN���^�)Z�����v��7��>�jRo"$��XU@��|>�='_���Eh�Ce!�p���'N��a7��������ѯ<��~�.�cz�����"^L5�.���jV�PR���L�=\�D��at��M�Dh5�t��V �v����`w,�s�KL�d�ڂwvtS�����J��[��i��mxIu+���ҹ��_aڒ�fjj"�'��O�[��*�y-�M6�؊�T�8���Pd��% Zi+�e��v��K!����Ew�_�����Ng���t����� C����C��jo�P펲6�<��LVY����%���n���9ZȪ3�0������f�s��<�`e���̕�*�`�'�T�5M�ށC�Q��f4� �"~�F�ţ���,��Ȁ���:`�R &���6�X[?���9���[e3�ck'�%e��_Q���R�6q7v���B��Z����=+�h�����C���Ϯ�2��o�YG���=I�MnN�zG����k��9;����,�n�~�($0ϫb�@�/��=¿�T�MC�;x�Ձ�a�'�[�"��,�
��t,�դ�,SNڕ�=��S�F�O�3$
�@����s�Ǌ�r3;��������o�<?w�H������b	c@�$OZ�r�W.�l�g4���������f�5��W��l¯|B��^�9��%��~���O�mó��JؿG�"�Q��=o �V��e�T>ȆU+����4_�؆�ʦ?T4�#��ѡ?6\�c��
�>1v9w[m�>��E���ъ�8���H�K�*1�=�ޭ����5�:&�HRe��	� Y��@ڵ_>۞����F�^*9Z1�S�������X&�������۩���.�<>���tK�m��`l�~��ٕlr��=�|�֡t}��C��x�C�ٚ�tnb�M�D[-y���B�g��J#�#t���?�VәJ>������ ճ*��I��:q�`��e��Y��zT1Y����w���|�� 7�d�2�!=�;Cl����u�)ҷ��Z��?`�f���7�D��H F#5��ya5DՏ�g�_{���z��Մ��{#�Z+YL:T�:X��H������������~O���)�����ɍ�����AN4���x|��IC^*�9..5`��v�t���qP]I��&�u���ë��|Ct	��_b� �s�^�����i�^>JJ���k*��M�N�t�����7�J��ch�a���	��`�B�ۃ=��B���k�ܫ�Cm%����Z@��@B6S�)Aa'#�����n��G�_cLt��qn
�����Ǫn�M��a�e���7�n�\j��n�bK�$����)~Ր �q�!�`��U�3A�f�	�C���H��<9���:ݤ�*C��e�;3K����4��;O-���taΛrx�~�+�^'�}��#�ȍ��4�����h';o����s�w�-V&Z���$B>�����hbp���4�n>��(ߧ��f��
zf��<߲�Uq�E����ܷf��`v�x����[4I�^�9�C�$',�L���&ns���!e^��j	�Vg�����D�R̐�3�t��A��?�<{M�)�>65��@-C�f�ae�Ghu[��oh�D�d�i?V�U��Я����t�l�Z���d@��?N%ĄT 	��� Ч�`�&($Ļ��fk@-�zb2�ط� j�x�{�jS+!2�)<>���3+U$�x@項���[���֧�7�m�����z�gS.���Q5V�FF����P�m�
��n�x����4_5D�`0,;x�q�$�#m�0@f�����b}��&���hXhd�������W�*�![ϒ�'�9���!��E�ys�6~p.��S��[�$��Ƞ���P�^��z�p� ����q��QG
~*W���v�������s(Tf���� [-q��(A������4c��Ӵ)�?�a��AE����i�3}���`���Xe����Xȭ�LczF��`�ǆ� ŭ��P����қ)`�yQ���X��a��<����l����2�p1��y4wfTV��f�XG�<�l�����=V�����l`�t.A�����S'='��]�6���j"�2T6a��FO\����*�r�~җQ^{�-V)"�E��4�p'�}�,8U�h�5#�<E3&�PjV3��Y�L�џD���8,�K���t(}n���{)�jI��k������b+�9uIZI���=<����f���U�ိ�*�a��G�H����6{'�)����|�U[��4u����,H5�I<�'/w�Z����b��� �&��\#�"��f��ɥ/i�T�W��c^ܔ����ȷ�Rx0Kh��[��UqF��R*��t.�p�%�� �$!����D�#U��~s�Cl����r\�\z��*p5�އ��}��Ӧ�N/%`:їA�+��I�ěS!6�c�+_.>��l�܏M���ۓ��˪����5�X��L<HJwi�z-�kcA|i�qI��oɾ2L_�G�u�Y�!ڋV\�3Y$�Y6�6��a�)<ߥ��]?��Vu�ș�4�������)���[+Sj�ܹy�/Œ��+D �#kAYC���.$������ZSA��[s�~'�D?�6�Lk����,}�bRwu�U`)�h��P��tM�-�2��1���������G ��Y��=�ܮ� ��kٰ4m���J6|#��07���B-0��}�g������DԱ�o���o��=6��j�� 	��"�RyX���n�����B��^]�i�[�ʒ��U�zܖ&�J� �ڰv�=�92ԦB=z]c�a�uܚTM1�MK������J���x=dfe�\�,]j��ta�jFN0�pK_a.W&Xf�}fS�}!����a쳲��$��Y.C��ڌ�
�jp�S���5�cB26�qO ��mIr~VF��Wel$"���L��/>������w�O((�.�k�Y?h����Y�56!PA��[VR��ά�zO�V��1����<����]ƌy>���[��d��y�c�{�����F΍-�D3��T��&f�9���X�U��O����s��A���e_v�n���s�a39�s�,E�@p䗋{հ+&P�ײ�P���R$�@7j�,��x��y�P�ff�VT�k�"�Z��|0��/�U��ȿ5�2:|�=��<����-�P�X��f��&��D�h��BpPu�e��^a�!c>@ƗSnRN���x�8CnYWE|"� Ԟ�td���-�g*X�ECvxKv2T�'U��֌K�]��R�Lc�,i�r@*�1~4��M_�����ܕ����n/�ْ����n�T�t)L���y�-^�GI}8��.=�Dɺ��PL�Uɭt.�]A����z�1�A�Z � ����f�*U�G� �
*@��jl�s�Ѱ(�z\�Oy[8,x�F�Gy���-l����G��|��U�Bp�8]��dl&���"8����3}x5ٕ�I@��X�$r��*��>��'���Rߥ*~����!®�H�o68U�s�����j8T�������x�T� k.:�Te�|��\���A]�B,��gI�{i�p!�`�;S*�j	�X�!R��(���M$lW��x��@��Y�3�Y�Z?��I5�9��� u?g���d޺'��-��7H3%�ZA�6��a��ڸ��psV@����1�� `��C��&��l�Fy�MZ1��zEaOU�|5��ޜ@��X"2f�+El�*�������n"�
���Gi��da�c��g��ɴs[b�}�}�М���$	���I^v�9����=(b���Y��:%��L�L���h��
Qtշ��q
��M{�����U?'����9k��R�\���{�#@�-��Ó�5�'EUYE:��|�V2�|[��ӑ�Ycy�b�����j�&�
�@D�'����䝨.5q�n�37���L]�xQ��%��B�F�`xS� `��hr�.>s�hb���`�9/�e�hS�,��*��."��1�6ݤ\��N���D�+fĚ�;�Tl�⻈�Hn}/I�q��D���I	�Og��n$7@Y��4�3|�
VS.�R
`�ϼT��y)��l�;z{])�H��u�Y���ٟ�^^����=A��~lE����R���6 ����4moV�(��ղ�n����(h�&��F���:N�����?�Mf����jO�Wt�_��ƀT�|�^���ww�a*��Q�����]7E�p�Idc
�7�ʊfG����Q�b�4���Էv"�'��E�W����Լ \�)�%&pT�Ӝ���eO�e�C6 �W�0��єf�!ve ӗ~��NFa͊>����Y�T�'Y!���맡�3<���0۴��B*��4�o�4R$���Yg��,y���VTX��A� ��.z�Z�D��p�ɺ2K�I�$�/7Qy%2����2�ul%�������恟'C���=���cLZQ�����#��H=��tp��eIr�*$|Y�Yy�w��0u �~�3{�<��dR6R����Sj�&ZYL)�?-�!9ֽKΕH7��(�F��#��Ȩ��0���/	�׍b'ƫ�;Іh��"Q��%� p���/d��������k������H��S�d���Ʊ��v؂@�q�#ۺ���X�-���K脕���W+�&L�0SL!�ृB:F(M:�/z �/7���	�a���r�h}Sb'����Lށ�Grl���H�v0����-��	���5"��(��w�l�{QE���^e7oU+�^�׬����Q�]GH^�H	z{��j����!Q� y ��݇aW��7E��*�G]�V-�\���>��b�M�^8
�j��On%Q%!�2�pZ��i�`f4������{�q8d��>5���k�E�
�������\�t���w?��P �+�&���	h��	w��p�7�Ɋe`&�t�w��@�A��[�����D�i
�T���M�o:�2{�À�[�!Ӣ���E�/i�%��H�O�&[�)e�� ���f�`�P,L 
���|���BC�x��%x��x
VC	���-s#��
��'<7����Jo������=�2&s#��6/NI����2���TB�|[S���[���n�����nh�3٭�r��"���r�s�@L��u'��r���J(ʚ(v��(U�n>���] 1�Y��)3��	Z��k�$�+�-k���.��'&{�Vvaf�q��-��#�1�ӎ�l\��'Q�`I�9�uxѾr~.���P��c}c��?u�j9A��|9�壽�,Ϊ,�����ʩ��������wC�S�*���d����qt}Pq�/i�~сl3z�{:zW|�E&���'��ѕ�������3%��0{ӛ��9����أGr�`����DƠ�W5"jD��
"��2����}�A:��<�y����#a��Ќ�W\�+�1��o|Ȯ�F�O��}\��Y��Y(�����K�C����`Y� lZs�k'�%�������i�jv~���ÑA��6�{�(��H��׈�7r�AQ�4NX�e>wRCmpCnGN�
�p�0h[���U��kź�����
/ n�I���K�\��[�YH�����������э�x�2�P������;p֝�Z!ᰆ���v���|]O��_y�����B�`�,iBI[cQܸ$��&���߯��|�iG�m2?�w8�w5��l1�Ҽ��K�2Z/�+Mz�DM(^R��+!���&.wL�.�s{�ë��w��7�&��(V��Z���j<6x	b�,wR�Vr���^�hA���z�%�p~����~����;�:E���C��Ȅ&C�BLθ��NF�أ�r�i�����p�\�����Hh���F�Ə-�CԜ*V�}�l�.zo�҉-N��DO�r{��tf�Q(_j��C�����,gο�S%4���rU�)�n���#�#G��j�H����>��}��]���r˩�Q�`Bꄙ�g���^��c����d�,�JBsE���G���Юָ��n�7�5ŵE����;�\5Ѓ�� !h���s������M�h��`Un���r��p=�^V�U�Uk�*�L��sXh�+ՃuG���=�{��"ߦ8����5�@��}DQ,ǁ������g�M��L���C
��B��Z���Rg�F���4Z����yQ�ma���2uaW>�C�K�<-�'/
2h�h���m�&��H̢�8#�Q�9
��꒍�;�� �2"�ІTf6��yE�TY�\F^�#��32(J@��*v�����~�a�
m~�/�'�&^��-.p^vE(�b�, ����| ����"��o�ܙ�')JB�v�~�>�J��/�_�@7�Swr��0au��^�v�0�N#9BT�se�W_訶��k��iِrW��ɱ��}�,��{��7�8r��;�L�{��R!Z�2@�ﾗ-XÀ����w=\�5�aGA�!�
lal���XuÇ�3�Ck��u�Mޖ�][��VL���URY����o��`�/!�&��u[z}9��j������<bDh,�ޙ��C$-�s�����ǒ��e�U�^�!�����sM< X�bw���rU~�>��%������D�SbE�2�v�5Ǘ�w�^T�f&)��#�_�1�����Gd��X�x7Pn �T� ��Y��0�STu��;�͘(���o���(�</L椣�mKȄ�c�3�Vٕ~�J]|1�[����Q�z}	@�fS��_ɰ�)�1ݾ-����~4��I�XV����� .|�v�_�q�^������N�o<σ��b/���1��K/���*\^Ih�X>X�h�b	�3\��EZ#��#�Iro2���&!s��O�u�6�J,�� ��081�oEC���f�a%}R��(����z����qC�2w Jn��A�J�]!*���>*��l�0�$(�k��\U�%�h��8}��SF3���������ǂj1�6�@�˞N��6*���N.�z�����)��fte~%R����P��y�z������$%[����7Hͦ����@`�Յ`��vi��ٲ2>]�'���Re��忡n��7����P9��xP�H��T �̖�bx&�����]#K�鰴�.�$�12M���b	��R%�~؄��	�VD�g������ѯ�m���6��H�Pl� 9��U���Hj�15ɇ��)7�����؂��{|j.f�Kr����,n"�f�dj�On�lx����:�r+�f���r0pY��颚���GZD]��!�G�R��V�1��ro�	�w��豫�@t��O�O��(��e��K��!�uh}��Q�k�YĹw~tf/�;~���+���4挺?�c�\o�hK�a���bS��f�`���=V�;3'U\y��cl�e����x{���?�o�CBcd�����5�I3b���L��뭉A����1%��y�iX��v)5���et`��z�Ļ�}�ü�J�\���]s�(�B��r�6"�����y��O�c��m��V�G�U�h�RId�ǍQ��{�y��$��Ҿ��_��2ci���d�����#��Ǥ}�L�w�R�N�����w|�L��q�B��`�w�'��k"��sx��
،8�E�w�
����1ko��B\a$��'���w=��#�#j>2����E�N43XO��Ń�@>�J���wM��)�l���.
Ms��$K1��� �%f�3�l�u.�*1(ڡ�����,������9��Z�C�%�M��b�] �.��iM��5F��$��jO�f��wJ�-���z����V�5`u��}�����a٩�;�2t��=	(j
Y�����"x�@��ז܀1|'���d?2#���awߓ�^���=���Cm&��j���i��o'?pCw���p6�Nrht ܽ��S�/gr��$$�`���M=%�@	��÷tˍ�Lu?�\���	�.�>�f���`�c߮�gѺ��U8h	#C�M2l�W�{t@���9��"@�J��۲��t�?�������F��c����%C� :e1̵�ǰ�"�5-۩RZ��whp��[
@�&L7�Iɶٶ�XOq�t�;��(����!�����W�HE$I�Ѱ�
b�
����Ю��:��L`�!��sv�|�c��	v���d�H~����w�C.�b����$�6�^����#��~�#���]�.6щ�L��|�%^#O�L*	v7r�(�lm����T9�J�R)v����m��3@����R��Ć�\��y�N�_D5�?46Erՠ��E�D��C��ң����ʲ��p�dS�@+�O�X�ڛ���M��q�j�tLc8n�]�w��&Ĥ�N��9b��g�l�l�R�!���}����K5����[Hh�%)Ov'���J���YR����$�%���ʹ,p�y�Q��{�t�8��L���M
2�z���x/3�G(�c�_���Ўx0:��N,`iB[�]���n�t}���e�|I�U����{q�� �>�sA���Ʋ���2S�Oӷkl��x�X֘[�aI��2��8NţD�����r�e�kxf����Ǒ$܂ل����`��ɾ*U�����_������kVő��#�\e�Z.�vs��,��$z
)G�S�����n�Ti�6f�'y���=�+��|�!���KY�{|
�4��Lo,lޫ� v�R�!�t��]���x�w쭦
��N�X�`�p2���%!����N^��sn�S�Vg�#\�����r��l�A����j��^q���?�-̉�[�'�C��㚾?��%�wf�)�p���:�"eh�&7Y�)�\���c��.U��d��1��r�-Iމ�Euii��X��BY�ҳ咇6J#�d�C.a����:��A�:�KT��xR�\�3O�ն-P�ӑ@4
�0;�xc�W��Z��|��nP���?�b��jA\�3],�{���$�0ne�dsC�M��;�{Ĥ< 34�$ዾ<@�,m��L[6�Wbi<����_�~_B��uM^�y����IN�����}m�y���g���Il�/�*C;��qmo&�k�G�rM5��,O�:N8�t�����#�X�Bςv��M��q��cX1���5�s���\�D=�,��/��%����Ys�5Ƀ �mԥ�z�v���d�H�ՙ��e�>6P��>�K�Kӑ�܏�֞)�{�(�'���2G.SN�-zE�V������급�����N@W��iǥU�>&�c���+���4�鰳�钖������ҋr�eA���}����a����4Z������^��,��VN <�8������u�@pB?�,�x�����d�[�C���c?K
��y�ڸ�=Ij�}��pcDp�)�$͹�䖒6b46�Yv�����	o�	z,�	M�|)�`��܃6����0��2R���b ���F=Z�d�C�F: �,M1Fs.?0�7���nZ�b?���ު�P;4�����hϫ
�x�iu�&T�F�{N�N�c���)sRO�Oړ�DY;�#�6�����J� A�H݃f�d��4g�Ttf9�+�7�o�<v�S��B��Js7�p3��.N�U?f�5��������]*�Wѵ"z�-��(t��sU���h�	�˭$�I�\Pc�v�=2d���X�_�~{���]ѓ�F{n�-����x(vu�QNp�S���q}�`��_��RWt��*Ω8j����8�`�S���)wH�qJ���c(���vت���,� S�΃t��_��#�!c6I��d�ME��$��`�>��Cp;ha��)S?؆�M%�ċ�3:�h?�I�)�eU1z��������0�n`�/,���/r"j�7d�\�KK=�SDp����%�q�l���ǿ8�1��tL|H��S�*`v_�)��	����`a�_uOD�~���EV�$��Y-3Xsd�. �p������Ӓ����	( U�U���B� 	��	C��� K4����H���S�P��HEAQ�V�|��uMTޛV�i0Jdo����T���:�tg>}��c�䩘��$�_V�3�eb{t�&tg)�l%�5c��(AΛ�H�`�#��I%��0ӷ8D����|4�/0�Gu�;h洦9�d��C#j���ay�Q�����%;�s��B8�����XH�� L̈�s�shGBPA�Y�e�6��%��CBkb˝2J<�A����6^�ڟ�Cd��W���@AY;(L�Ӛbԗ���*�l�#g�A����j]��lL��Gс�>V���$��^�{����ڄ@�ڬdO?m�Ҩ܇v:����jP��=s�eb+�:I��f����RD���C�	��j/O���Z9�h8�@�
�������=������d_��b7��ՙ./S^t:
0�F�r��[�Y6�L|��Et�?�s7W�h��Ʀ��[g��b>E�S=�5e�9<�g.� �4��V�Q�8�r_M4����Xu<.��Kk�F���(h׌T$A!��pZ�HA�5��X +O���e�0\;���.A��"���T%�`��'O݌Z	�����92�.P�gxe��3�
-����I�lQ���߻G�M�0��sT
M	ac�6�d���J]C�_5�~6����K��{{Ƚ��Z��ex�˾c�sb�OA��ށ)�ΘC�߀ t�w�4M���Jq�)��"W��nJ,},$�^q��#�ڻ�4~j�uD?q�f���f�<���Z�v]��R�⨣�<�遹��q���|�'�-�������Ҫn��⿟UA�I�~+�9�6�a�]	\Vn.3֗?��9|��%��%�4U�>I�F�{��]�B	*�T��V#�
7�i�����G��(`��ȧ�V�8M��]�J�ʰ��wڌ�oD��J ���&_n��hF�bm�uw���|���K��7���kc8
ǃ�|Ö���dB����cX�򊐛���u �19*h*F�%�Y��A��|�ם�V1d�B���3������K����ָ|v�c�b�S��M�<�D܆�GH��9�P���Ւl���j���}0��� ����q�سc�Pc-��Ęk)�Wa��?�-�.�]"e	��8����� }�s���,5�������hb#FЭS�f1n����G�s~�e��9m|Մ�mad�G�-i��+�g5����1i��;�����l��������Bk�{ư)�� -4Ԫ{eʂ�O�ƻ����;PZ�kw+�2c�]4G�4{���@y4K;�y���d/�)��)�!��T�/��r�L�h�-��U���%����A�Ԫlc9o���x���e�Xxɱp�pjS�1f�Ɏ�L�S�N�b>�����˘�wWw�1�w����m'ܑ�}�ϕe��<�O_3�W���Ү�z�3:� ��d2�&�
I�۾�p�Aw��S���Y��U���mgg��8��\�+�j�K����QՔ\����8s&����n�ߍ����Y����NX&�:4���&�8H��6�)����߽(?���� �½G:qρN%:��z��q:��<ts�B�Ճ]j���:��iR���>��c�1&�r�c�� ��-J��;�V��0h���������) I�n���+l@�t��<Z�-.�\�����A����:�\� �>�l��Ħ���΂�G�
�+U+̥�l�P�TvY�L:�ؠf�:���;�j�k����2�b��9�H&�S��9_�:�S"�o�WPk�e2���F�!җ��b+Vi��ܺ��4��2���0�4�#��}�=[��O B���(���ԧ���\t�e����cԻ6�mjEG�}�kM�,���C�zm9���\[ǭ�A�X7K���$���|tSx��*=>��/>���0��^'����sy���8�ME^�U�T�����4π�eS��E8�=L8�u��г�,��-Ry�Q��4�h�n�o�_!��w�+�2�P
և5�����`�E���`6�b��'���1pa,?�*��2dX{Cb������o`9ҶG�Bt���2�'����@p��ԀO��c��ŕ�L|A����|�=��X%�wg����"��TP��?)��f&�����S8����F�x�/�l�GK����0��a�+���;RB�+1��w�~^h�ڿ��ޑё�� �����p�����>�ާ�	��'�x�>Y$]
�)����7J`m?�k�M�D���` ��ͭ����ʥ�p�����c��D	��=/'��hO����!��h�b�̂v�����A������^���"6[�Nr�L�
�V (�S$`$4�ݬX���������� ���kq�+"-J�g�ە��V�y�h+?~6~r}�$n�8�{~��A�.F��"�:��ܹ5�==e��v�Q)��{ֈ�M*Z�T_�z~�m�%�`
��?��� c�xhO��An�ƬY�+��.B
�f���9�>���L�r�����\��vǐ��W0T���D�A-h��p B�����a�H6ddU��#�^�Xmg*�c�jʀW�P�Z�(_��t�:��ǽ[2R{� �C�X��S�o3��=K�
��c�;���T�s�q"f���w�#�Ts>.��x��ً)��Y>��X��-pb��џ�j|K*�"�,ǯ�m����B�h��HFE��JA���O��pҊ���T�
�Z	�%Z�l{�x��'�+`�s�t�{}3HK�2^T������?~3���(���E
yXnPK���j�V�h���t��h5��
��:&dK�6����A������B�Q:���&��v���@�'ؚM�|NG�u�g_¬8JA�fK`*ܸ,�ݞSD��U���T@�;��^ll������	>����JGB�j7*��C����[oI��g�&`��P��'w��r�*�B���h��dӕ7��n��-�k�J|�X����>`��� IGr��5�	�4L4����
KyS�o���*�?;t�w��B�5	��@� �{�t�%����5YYx�e�L���є��ϱ{��17�w8���B�t���)�gұ�m8}'`����X;���	�?�m�_�f�N���N�s����^;�C��]:Z��RR���0�9$��J�}��fU􌃠.��n��ʟ�)k;Q6E�X�E�O�#\�[��M.�_����H���%�c�]�V��_�(7V�������Ʃ�,��	b�5����o���4u����s;�ڗ��=n-D<�p��g3���w��c#>�t͢�d`mpʜ�I]�3��QrU�B�ջ�q�n��v-�9���V4�8H����	T(ηXM5��Ɛ�'��+��M�у��R,"qtH���--nK�xU����w��A�A��#X�{�kB(��sZ�P��%sp. V1�4�p���LN�����
NP�2��(�7)҂�sع&ǻ�ҵ�����.F�U2���z��*"RiH��� {|��^C*4A6|��!�c�D�U�Q��%u�9�L/����Y7�9Q�r��U�3�ʏ �R���5)��
z��aŵ�!I� �/��de1�C��BV�0C�qX�����V�w�С��9�7��Wt8j�����V��Pl�	tP��#�:�n�N�6�v%@g���IC�f��o%AϏ�4�P�.g,�o&x%���K�@�[��yd����㖺��g�	����Ֆ�K�dH�h���~�v8�@��S�ջ�uKF��PE̪oyM�7�/q�K.C�_�'�^�rD$��ܼXP�οX��s�Y9�G�w�L]�����D��-���O��i-R�a��Q�n+�H_-��V�e�
IN-ڼF8ah#��`��~aO/�)�te�У#>�7@&����Law���c0qwr�ޡ}3W�N��lB�Դ~�`&�27y
bd�7���}��<�ͤ�%��7 c_�	>��SA>���e��ǔ��q�R�w��H�!Y�R?̺+v��(*<]�MK:C5�?F=�5�@�'�^��=x��WtR�<l����),U���� ͌�Q!>ӵqA����?Ŏ>��g-�����H�ZR�Nn�����D���@��\���P>�ۏ��)����-��̾+�[�ܱev+��s[f�.�@Ŝ�s�F	�)1i�4S���~�b4�_�n�柳�C��L�+_�4�F�cx�/i�c
��mJ���b�#�Ћ��|f�tIsx�gW�W�Pg~h�R��%p�97��9�DyaUZ��c0ۖ��P2��7�.�z.�E��T��v#���k+�@����4bA�<��l�C���)�����wZg�{�~���G�>]�
��o����U�pRJ�<yC���t� [�L|,@�U�}��r3�Z��c������O�Z��s�zx�-8s�/�0-z�=����S�Y6����O�t���H������M�l�ኟq~j����kg�K��L�܃L�}��Q$�g��W�I2U�]�g�+�E���д`��+|���Pݭ�3+�TZ�b�5�\_;S"'�}�b(({�kH�!O#X���溯?�WE]��&�Z���B/�W��(,
��J��������G,��:�i�YX��'dL4~�3���6��Y��O��{H��Sڟ3�����
:#�cjD��w]��v*��J����5&�	 	F�����3�:�7�U�'8��`�Qh���ڞN�I�fi�ǐ���=�>����~�[��*�Z��,��4K�!k�Y��SRC�%�yGd�����#f,�}�dex���4�Z� �[	l��;ӂk,����a���M�5�*ѕ��,C?��קځ�����? l6�׳��M�ನ�=̄�S��n&o��:��L
�v�+̎�I���V�%��du���^QT�Vl���|Kg��`���֢ץ	�~��T���D��IY�F[@��WAs���뼨 b<�
�,�����	;�h��;v��V�Q�y�o�?��]s'�EV���+��"�h�+~�^[�ˌĚ�Cd�����>3O]��	�n�(;��|/��&�H&�:�]�Lv�-��tt>�a����_n���S�gf�}M���fX��W�N%J���}ך�É��RK�X���J<N��?��&�ʞ���z�~��-60Vu|�H8aŒj�p.�}��Y.H���ѻ(4Y䗪-S��F���h~]�.J�Wd��)���e0>x`���!=�T���ɯ]�GZ�lp[���68����M6�w�?��%2U��,�y ����{S�
o<	�/�_�n�f]�I����:~�W&E��,��J�j��BH���[�7e�ʍ����;�#ɪ�R%g���О����3d���*�)��������mak�w��ȟk�Dc	�I�ћ_�k ј]�~�̐Kъ��Ųr+u�̄��g��,�c.�y��cq{V,��Yj�T��c<H?T���U��Z�M��ߧ���!Mh��1�zɎ.� ���p�ƛ �a���p*i߅W;&6z����W0!Y�F�T���b��g��l߰d:xN&-j����̎PAaF9���h�%Z?�J���:&�);}��c4Z�}���<Q��S/�!K���L��SY��ƝK��k����n�����"6/���!�i3�������؞��G
��?��l���/��1�h�	��y��	J�.���D�]��2	�W{>�@'ĳL��<t�6D�������Bb�lw�5p4��x�Zc�/D(E���2ͷ�i#���뽃��0���\E�7���0��n�Q�ܹ��U'�� y
>aB�N�4�#-��-$Fx����b���E��f8i
�0�]���6�i[U'y���,u=J�ӕ��U���	��Ȭ%MNZ��%�Ǒ��{�)O���3i�W�2?3M�B�Y�����ws�G$�K�|���k݇}�^�~{�� �A?K��dY%�
�Ӆ&��0?��#WPX����Ja�z����[�J6����a|���E�P��	��$u�#�#8 H)�?�DؓH�->�����#A��U�Ģ���R)�vƪ��d�xM���e�(�P�/�J�87�^#������� t���w`�1�5)�����g\�k�(�s�� �9氱�艬���9�\k��Cg_������*�S��)��d-�.�M��x{���IX��"��a���ەWĺR��Okt)k�l���d@�@	5o5Q⟊D�IJR�W��=�k�o��p�o{"�ao�r�7�r�05o�^G�٣w��C�#�u�{��c2b��'��>t���z[V3k>��QV��<�2��dI�h���)����-2���O;G }��F�@�����9��d�h�-��������R;��b~Z�ŖgL�D��`�^��K���+�_�X�@����-��Dd���S���-f:\\t���ń��������9{;�H�]��c�xF���֬�!��x�<D`_�B��ȱu��K����0�0M��BC� ��]�;�T�J�]�F�|��`Q�hb��]S�dٕɩv��][�~ѿ�2�7�q�ү�bA�3��;��k�g-�ߦ0���L0��f���d�Q�/��|H^E����A�/�+Y��j�P͢�ɷ�ylF��d�~�"���J��]�C<�w�Af#��(M�eB�TX�"{%�Q� �{	I��	��:���j%�=���T����Y��Ũe��Q�i*"2UH��n�|�X�B�%��Ěz�gx��[Ԋ���9���D/�/׹+��Q>}.�"�C�ZWP�3�����e��M�`h�Z�v�>��b+��t?�'��/���U0Ҫ⭧�4��2���'a:������I�q��G_(e���J���XQ�D��l��Ege�X0%Ey�a��k�QaD��Lȣ�z�p��0w���&m�E�"q�#��^�
�fy\��r�X�:^��4�M7��3(53��Rڞ\()t2�*ڶ1�Us����a���[�W�+���w�u�D.��~� A	=UzLZ����,>��Ft����Z5��}F[T���]��k%��ٚ�"%$pW	�?������� ,��F�j��W��������E���I차i�]F����_�K1����jgiQ�ȳ�4+��o�s�ι�ōO��Ц����]0�3��ų���+a�u&S�!	��[�+�u���j_2�rҘ]T޿�c�|�Z���G��wYP��}�9f���HCǬt��r����VC����������b��-��}J̣'}����'-����E��g��𼳸�{Sl���]�؎��m��#Ap��aK;޾=��;�<�t���Вv�C8��r*�&�a��/P9�����&� ����~>�����O��zi��*!�v��/�x �l���ɻ��V�4������ ����&��g��3����!f��s�2�5�>!����ʃ��
�h���#j��d�[�D��V>��^ښ�O�?͑������>'R����*�^ ��XԄp0�v�B���U���-Boa��x����K�k��yUBX�re���~+gH��������)mYH����]Sj�� Zf
Jk��o@U�hƠY�0#��p���L�N�LH�������b-!���J�gP����O�{���W,ʎ�7��[�S`�g�U#E@ј��F.xZ^Jr6���Xq&�`���}\�6OX����B����@���D�P�����n�|vV����d'��������N,x�s�g�ǃ$P�7�m�T�!�t�I����]x����CQp�a�/$�\��s��EoD���t���-đ�:Z(?�7ԭ'�/?ˍ3�a�2�jr�A�W�\�۵>y_�I�q�<�i�.'^�Fl�����\6�$G���{��S�T�Җ��8#��h��-%{���ڷbm[�x�\b샗�e�'Ǖ�I�dKU�uET� ��<`q���o��lQ������n2�I��]�#�8�2���h����sJ�|�_�	��K-��*���":ۊG7�� P�ۧ�G,�4�c��Ԟ�P��la�H�f�ȃ���Y�v����s��H�)���/z �:+�L�����W�؇T���rw��x��It�b���v3�"u�4����IsiSecY f��%2���f��w�� �ޞ�">ZD�t�܉oA¯0�5�)�*~�9I�� ~�hث{��d��`��Q�)_�tq�꺭��˒s����<���2�%ն���V	'�H����N�d�`b�����b�0a�TTX�!� �5�7�*�_$�е�� �~����JM�9��4�+r���=�������2�H�D�2D<���(��5R����?�w���͏�:0�%�_����(*�K���֮�noǕ2�5�#-�|��ե�uJs�L?���(��/��N_�Ioi4�Snܶ0d���yot7����m�0���B�����WC�,>-1� 
ګ<Hư�M�����9g�a
��~�_������RD;Q�@ e���������˽˅�*�>��[�k�MJ��� w��A����*I�5-'b��3z��
X���*Qt\�ID<{���I��B�����
|�fJ~ZZ�S�{�dvRv/Z�K#Id?5F�h�a�ל��a��Ҝ�Z�E� �v����A���"�͔�~�: ATDR87�	�D�L��_G��@�:~�[�ΈX��UK��$9�Emr�$v����������=���q�S�h&�E�F	�c�)�3��ş*��ק�⫝�Wq�<�F���W@�I������ㅒ�2�����?4¯�wB���c��D�:*��k����_^t�ݮ���g�;o%X�Y��W��&��
����҂�95*�W`O�kO�x�m��E{�.�؃V�'k̴�]㊹-Ұ8^z�w�JG*gs1NzHкa'��O8#��ѳI ��m��+�{�����F���H��!� V�s�n1*ќ׀���n)遅z�}w8�k�^t��+�|	Ug�i���Fɵ>I|�����F����n娀��V�����N�1��7�TJÔGGD!�ύ�k8��-�2 uvT�P|�/n�	��$���ū�1'��c���-,�
C8�څ.D$�px8�Z����%��?4(UF� �,�=E��	�e��L"����=��e�1K���k�m��lF�y�À��Z���3~<�b��6pv�5t�{m
�ƀx�(�>��۴�����H@� ��S\T�xV�C10�ލ.Nx�N�o��b�a�<�,��C�Pnf�b/�2�K)���#�R&f�6N��P����qk�\G7 �]~SŖ�$�l�4>+������ʝ���9O%�خI�~��;>������g�0�wScEsȿ�<�-���!����Vg����@A�t95]IfyC��-������3��gT�5-J�����=�*U��HӘaw}N�O���8�gy�Z"�0�}Ί�b���Ҫ�䫚�DW���������z����V� �(pb��F����+�g�)�fK���h��Ie�^@m!��.�N�0�"�ܒئl5���$�:���Ѱ��Eݠ�(o���CW�vˎ��g>QiK6��\$`*'-nXCi�����m%���١��0����_�����ĺ`(���7T�\L\
��<z*C�����Y�ȭ����
�����u�q@z���6�7��~7��0t�n,RP�J�`�c���fQB-�mCVY��w]B��e��-o]���]?g�6��y
J�I4��F�x�@�-Q���`�ع7��QR�ց]���H㮽[�i6M �pӂ���8h��r�Ԏ�(Ո�����`�C��)x=����L:�Sؗ
gc�w������K�U�.���G�a��D��_+�xA���*�1�?G�l���ޒ�i/7�T�X,����о�P�2}�ٜ�`��I��,&�wY0l�^Q�2��{���b�ˋ�cɮK�r Iv�y@L����8����W}K�5�U�i��!������f"�P��~­�-
 75]���eٴF֜m$��n��MKt@��Sʚ�T�"u�2w�L�7@X{/׀n�,�_�-"������mߥ���7q��1c�k�N�UL+��r����D������W,��D�~Q�΋r��1}�9eA^j�dv��i��Kb�'ߴ�,����h4�C��\ƎŬ�ܬU��Wf}�W�c�*������s[tsP㟟���S������c����2�)�^M͇��_���q!�|K<�DS�|��V�6�������[�>���_�(� L%�|y����P�
��v YO��j�\D� �C��v)�P��0�^�|�D�C֞�̉Gi��yT�am��NN]�!L�̪�a#�(̮��ĩ^�+�e���3zQ�v
��>9��Q���'�3��(k,���m�����E�b4
�$�h�L�#�������}(�t��LYv ���{S����t�	���X���3ca���6_�t�2"&;&�(����s�q�|����M,['v�=��EB��F|*lKSཧe��K����i`�Q�߸3L3x�VHe/�X����Z����sj��������h�`�4��=gIQ&\�l^�W�!����C����'{�g�t��2�מAT��,[oI�,��5-_�ˈ����é���tM�?N�oɭ�m+|�n���qG��C�хl����I7����[5����8�<�+��ϖ`l��BT�:1���U_�J/�%l
��S���Of	b���n��捿�L�m�ש���țyz��!�F?l��Y��z��A%o�XO3��v��%a��5jM�m���n�n��F?%��T�H钞x�ӥ�lt󉤣�S�n��Z�1����{�M���Ϩ���yp-X����.*ѷ{ � +#���ޟ���+(8�ت���X�9�ϸ�/��i��ZG٤�ZZ�Gɓ�W��d�K#�+ό-�#�k,��^�[w��^3�@&%�؛����I��24��n�<��S�'�M�"���X�8�#c�Gnu=񓗳DA)��t���'�k=ƪ=�51����4�����j�o_o���c���፞��{���1�����G;R�'j��奸����엲Ԭim�ӱ�+|˱|�9��a�I�¦����7g����!]�|7���+�C��NDF&G.����*}��J�g֘5jCVE-�t��P��'�A,���ذU���S)�{��:�n�4áǷ�it+�������٠WUe������}"N�p��Ӿ�x
�v�e�����kz������B��-{� N�F�v�6u��EbGLmJo��1�h��G9�%�Еy����ӂ�)��C�4�"�R|6$���F;�ZCL��f�O��o�4A�Y��c�2�_lN��uzY�r҆l�y)յ,¥;a
��:p��c�R�p��Y3��쪲}����(h#���m<�E�tj�9W%=���=ݮ�P0���X��+���v�´K�L����7ؿm�$9?�\"�J���~�>�ף���b�L�1ߟ�aZ�#e~y��Գh
�D>�Ɗ�-v��mO�~9S7Т��"�+]���S��A�on�<\�2��(�`}l�x�	/�×�� �[c���PӍ�^|
�+���~�L���/`�F*<�ؽi����(�3��R����k�8�Y�)i�c�K&��<�!��I�ZTS!V��}���ٖ�D�lz �֛c�KOճv�p&]S�%�|xe8�4q�*����xEX��U��]�%h;cܵ�)��Tz����x��r׃�ۨ���%�F��;l3�g��s�tzfut�@L�$�f�]վ�I�(��q�v�\F�0w��.��?�Ū�6N��6��f9�FALܿ
"�Pc�r���%�P��E	�hQ��0�_!��較KY�� ��I�O7,�d�\H���3���d��Z�PX$ku)�����2\t_2�{�#�sSg���L�j�ĺ�qRB��,B�v?
����҈��*�>d��Qa��km�G�h(�)<�����B�}K}9$'��,s�_�w������O���γ��Ge���"O����̂�� 3�D�.�V)I�b�&�#���h�bM��(�X�9���#�b���gym����X|��Tz�|���ؑ,����m�Ŧg,K V:n5�)W��1n���k��F�Krt�x/jͷU�ܑ������l�6�w��*�mcSA�v�&pj�<�$��oͲO�I�v�"w��Vr��\!�k�r+Q����]�ܝ�o���X���#�c�@#/P6)�v���̈�mײ�I�v�G'#"���uj5������b�%Y�_19��������+�P�27{���V�Ld�=�֖nk0y_�W.r����#�gM��
|���M}.0�y����C���$�o�d/	ޑY�~	��Ȉ��Փ��g��[D�i.��S��k�iҙ���;M|�������h߁G���B�E�%�7�J�f7
l'<��?�cYw��`bF��9!2�{�Z��Si؉=���ɿ����F�ُ(6���u�
Yl��Y�Xq��W���i-��^��=Gi��w�]�[��̮�ʭt�U)U�7�)��t�F6�b9�D�$���T�D�K�/7��1KR���`C\f���ƭ�JFZ���ԷYeD�z���	/��37:Z{챸�XJx##f������~r��$�v�C?��͜�F����`v��C$���ۥ����i��ae�>%*��H�k6�%���S�2�� =�d�_b��ī�*5�i�1D�l�Y,�<X&6KL�_y���gw�$�&5�蟵5[AF��5 ��W/3�B�]��s�F��m�H1�6R1�X�u��N�ߒ@r�֝z��
ۻ�����0�HLc*�.����2Ve��r�/�:��k��r��gm�u��5�ӈ�=�#y���To�عwlY�e7j�aG�T�0���ʇݑh��5,��o�H����t��}\���m�uy��?�/�f3v"���րgǽ����pά�4��G.����Qx�Y֧")��E��u��iœtrd�����T90��M�7�
�V/q"�Wpʫ�'@�`h��4�=��$� ڣ�?y�#�K������n��,i߄��W/��)IV쎆!0\}ɭ���Ztޕ�\i�3 z�x�>[-�#�DB�K�O�>JA�������qd�+�pn�����m��F�Q�!�h��H�Ĭ��fn/��< �	p�Z�[�����ʏmpgߓ���$�5�V�{r����
î��B����������2P�q!Z�D��V�����ش�}��K)�m�iF�+�Obj'���WT�T�t
GVW�{/���G�F�*I+����W��B�q��q�}�:��2�	��+�F�~�a�i>��T�?t��o��9Nβ�+�O�UAi�e�X�zP~��]��ዖ�$!
�;Bh�mF\ϛ��TY�j��2ӰP�c����0:)�g�
&��V��p��Y��zᑛ�#0W>d1����꛼�]T �*�c�����}lbآ���w`���G@�ód^
�.��γ�ް��:N�Bܩ%�x�#�SvVDRz�<��"^��>l��|�Uumw7���Rvd�o��.�9��,;�0	���^�� BZ���G¼�|ozEf}��L�2��Fu<<1�L�I�4�(���s�#k\h�ǻ���$����+��R�Hx�Q#+k�R�46wj�I�1RR�&��2�?cxQ��Rj�pf�����k���`Z@6vȁ����7;�+}��Ԣjze��'!�~
$��5BF�+3f�opM5@�������9��St\��[K�ʚ޽kR���H�Ū�<��L�d~Ȋ�,_J��ܢ���;�eԦv[�����M��tu�U�9X��ExZ߭�3�C녝�e�?P�ꓱ_@�J㐸
��TH��;"O���N۞��ҼeEe��#�����;�S&40&�t��+1���j��R@�cw�uq�\�|4n���3?�S��xDL��@ρ!Ze�t����pc*8����iҒ{�׿@)1z���$3��Kzz���D���!.=wB��JO;vJ��k�Bo�"O|�L���
y�m��m������	��4���2�����a�D8³6>����ĎZ��[������gWѱ(�g��vh����K�˝Rp<�iQ�K�$C���	Q��m$��ܟ�M&�d�ʋʑ���,�B$q"XA?�&-_�-.��mp70�K�����[��.�(�ByR=v��� ��k��>� ӎ
Ь�(���˧��1򒧜g��/c*� ��s��Xv]�G���;26X�"�0!�f�W��C�nG���
+��y�(�[0��'���{�M6����0bC�n���r���-h6'�f'����t����X~��Ė�\&�y2Kc{�v.\����\dd��g4���#��fڷk����id�M,N�p�ɍm�١��a��ۏ&�����3
,[���D�9���j/>���b2�3xzv��)��~7m��WA `JGe�����3���:K�6Z�mu�/Y��,LGy)��w(�
��
~���W>�b@(Ф�4T��)t�R�:F!g�3��{Jz�+��:S�p����9|�\}9��l�e-<"�??צ
�$J�v���{>�6ּ����::�2��8�@Z߆�1�5Ҵ��������%��\4w�"4g&���(sDWL��X�	�f��[z�,mPe�u�����*��Ip�#��8��]�\�k<2	5�����u�=�����-�޺�|�R� b��%Vj�64_��F�+�:T�2_Ʈ�9j��mԝ.�r\P���Y�"������%�v�v� ��I�ʦګ�R�[r�i���1Z6I���B��u6������H��|j&M,�f��u�F� !�e.�Ӄ�e�u�VB-�)Ĉkf��aZ�Jz���m@�$Qfc��L����m�Qp�&$��+0^,ot9[)�N�D��0��@���=�l��?�"�j���{K2�Y�P��j���]��r�d��"��e��g�AEw#G)��i+52�6�kWiUvP$"��g�F|�Cd3���]�@/�y{�}�Z����о�������&:� �����0��Ay!�b�c�b�H��B#���oЉ�����U3��̨6���/`�y��N+5#��<3e��?�=ol�F#QM�P�0�z*�m� w����lf����I��z��A]a��:�C�ȋ���dJ?Di�����l���,������3"���$�\ΰ�"ll����Kv!J� ��h�1~�xs�T0$j?�� ���[ l.�F���%ᷥ$-���Vq8ǩt�9Я��tz2����8V���同D�nskEP4��s����?�8�W�0��\��qq�t� s����\%28� �������R���Pr�d�o�C��u<�$�|�)j�.�%��U��Ӽg�`��#����"`b�(l�'ӿT-w��YCw�Z)�y��d��2%	<����?�Ae��be�p�:��"}/6�&$B`�!��*�_)��"�� ����3f_���t8pT�J�*A�, h�?�+�h��M�����#��b}�<�>�l�>@>сK���� 0��c��)�C�\�'ǳڡ��zI���ea�1�^Nx�s��p��I�g�Ă3t�h���$�gy챡`��9��W3RǦ�3��x^�ap�X��q�	k/�L�\����^��;na��ʳ�!XGc�T:��I�w��Hp͟s�V"ɚ�Y2H���v{�e���� �6~�~9�.*��v����6�B.-�l�@�5��*��ʰ�*d+kEhpN��M\�IX�`�-�i�R�T�|R��/h�Vı� �|�Y�vo��̙t�TS�����H����"LNPzw�[��nb�ڈ!�� L� ��՛/�gKp �r���� U���W�ˣC�̞�y�	���&��I�I��*��4g1�I7�����?v�Q�� ���(�zY��.Χm�Y�"�w[��U���`��E���g����I�p��iv ��P�}���p�&xQ����z����JNsG��M[�]̣�dG���j&�6=�tp��L�<t?�P铯�HjݮȆ�՗�4�!���H��C�9��>g�}{�VULV����5H�fS&���c"�d�Dtb��	�*u&������d�����3qҟ�p���~�Y
�0p�Q�>x4�uǓ�JY�n|��Ԇn ����Ѣ%���.Mں5D�n#z����������d�ճqs����I#����S��;;�>��%�]E[/R��KX�p�b#%�<~C���S�� o�B�V��/���VSr����`��L�����:�}����̽�4}ljp���^49o%G�F�q�9ah�[�on���=	lKu�1��j�o��sG�t&o&`�9-Έ�$\	����q�?��#�H%ܽ��,�G��C�ڊeh���`M����r���fx	gK�ס#��cR�P�	#w^-���P�F姥�b����bT�f���S��?C���r?���� ���6���ԣ��X���RR���a�zO�LN�yI|����;���?8p�nJeg�3Sӌ��,T�����EU�=�/�h�J/G=ϙ>]Y�4У�1�D�M��g�ʯ��rs����W��ǃQPM�Gҙ�=E�c����v4cq�m��s
��"��j�c��xzA �XW��QVڍ��|}�-/��X�%�@-ׁ�jli�x�����>���0������E�E�����ut���z0��Oר�?[ �ez)�F�����	�h60����&扻�k/�������w��w�(�@)�m��6��fF|���3V�ֽ�ƼZ�� x�������TL���H�c[��O�a�"ic!ӱ����z��f�[[@>�+�;�'����O�����Q��9;{ �'\[P�;�� k�S(
Hfъ���.	"�֟B�l9�B�R=[g�z��y��A���Ϝ��x��^@�{>4���E�Kύ�a����	pnw��\�d�R�`�w,U>g,��CC8�A$w���j�|;(IU�m7�#�����S
� Џ��a4�yI_f��� +/�,�n.O��&�����r�"��M��0Ȇy�P���LD04X��چ�)<�5uvѭA�3�C�~����F,�$�qJWȲ�����K�y���u0��AfPXNwP�B,��S�\�wa
P%��5�:���P,O(W]�N�u��ݹF�I�v1���RH�\`X
���4��\���!C �Тg.���@؊��o�u��7o���ڊ~�GbO4�E=�� .'�ɥYs����cb��-�]�����S��!��VKR��ߨC���"���X�"�8����Q2�---GEi����*�r��ÓR����E���~�qԚ=J\�������Y�o�14����߁�f+4B˂��Ŭ�M���������hb�ģ�=X�Q,�,�ʤ�x�#���((��ؓ�)���}h���ￒV0#�"���J���M
 ��l���f��G�M-@�\�u��V��z>�:$[fa�n*���ȭ_�4�=f��a��¿^���'r�94AƟ)�y��7Lʥ���s�Di�ܱn�i��9������0}*�,wή�t8�� ��H��M��-��A�d�Bu���\TD�*/���(����D�����zz�s���~Ȅd�r:����m����
_�qycF�����@jb��˱l�$�P�p�$�����R^@r���+����U���j�T�5�O�#�b� ���;9h�3s�,Lj��`7�c��c� u�v��6fP�j���E+n� ��E�}��g�1~����S�n����b��o8
���KI�S_��پmE[��0�$`p�ۆ�#Rxʮ�Х�<�`��>���K��)U���W38	�n�kѦi�89�0涖4G���s�����,���ₜ0�x�lz��;�"����ջ@�͡�T��I��3Jg�V�̰��f�%7��?	�1�M�j�
�^��'��.����Iq_)�BdR�cw��z��!L ����"a��Wy^�vJ���3$�K�bq��_��C�X���ڐRoe��~{j���ބ]��7�9�]z�₱$��e�ޣT�=+sB(�!��[��f�op&��<��Հ�s�iv��/>�����8+�RZ��68��C)�śơ����e�2ǝ��/�$*.31��/���	�<wL�&�k%��^�
W�c_�X�Va3����t=���� `�X�	�~t��!�a��� k�׭s���5����C���j��5"� ��4�{ޫdyuZV<�p�~�[:����`P���ī�oG�F�a��jM_��7�{B���
R0��P�:�X��U�ƶ�=�F��WEk8�*0QSY�@�af��!���O*k�ʘ���N�qD��ش�j��RJ[�Bny>��Z�-n�<� ��W\a3����><8��w�G(��A�T��Yio�*�[�.��ȸ�2S�r�]"�'�� �����9FY��j�����CVy���h�C��,H?�?�$���w��P���|_9c\�a!�a�Դ��>Ӻ�%v
g6m�q��!�TO��k�{��ٷ��� �x[N�<`�Q��4��U��R�M�yΆE����j�5C1Aؚ ޟ�
Nܩi�V��������5�%a���Ik˘�^'�J���`�������&��Ñ';�V����q��PK�e�:y7�k*ư��|Y���C�7'��_�jO����x�@Uml�+]�+У�` �z�Q����ib�ҩ�7��������\��èL>k��ϲ��pnFA�����b�/a�;G��.��.ĿSF�c��&��S�ޜLH�>1i>�X���kkG�'��&JE6�������e	�O'��n�ʌ<F�ɺ7�cl7��mm�8�b=��U�0&(�2��b�h���о�d%��[�w�ގ1�v�v�}���X�H�hL���(:�H,Z��
2<`�L�|H���VɯeC��)�,[�T� ��8��6���M2]�y�7}�q,��S�3gd�㩖��D����!�g��Eƕ ϓjǧ�0^��yؽ�M�E�Y�d��)�u
�r�45@�姝Sq�V�[P%֤#�Ό�[�6*k��/�?Fw����##���F�[�}a2?��ɨ�gH f�u��i����o�e�Cn�����+�jZ�G����a3��|��(I�ʢ�˚�޽��B��鹡D�2��⥝���8��Ձ�3�~C�ܥ�@�	,�=�3���[������%�V�Gl�=0$��Ѣ���N�^Kf��<�כ�-���9��U��/��Tρw��kp]oQڬ��@�N��7��AJ�΍���r����Vu�%r�	�7�\�O�tN��,�ц�^�5�����V��d-P�;��m���e$��@��/�P#��:�����Nbv�<�M.@�x����mG�1�J7������^�ƕ��b��ޏ�YA8�'�E��-�'?_F_��ً+��>c?�Q�?+����ë%y}�K������Z�W�_�NUղ��z�T�G'�]���kR9%��o������9�3o�Rݵ;�`�u�[Kr�[��T����>"z@���,\�<�@[z�� �J���w澶�О(4�\��_-bD�w3�r-U ��lD�`�/�F�ʓ2t�fU/��7��T5��5�z4����F�Խ�)�&�>�5���P��L�;�/Qz�Ѫj$�Ua�����G�o�rg�����0'�L����
�m�}�2U-6��S��	@tX.�v`]��N���Q �k@⛥��;N���^0�0�yy��׉J1��ƝZ]J_�[q��'�*"�cv����B���W�hb=g��^U��O�J���G�H��A���c�n~,h-Q)��aö��V�M���3(8�(�����A��I� �L_�\���-i�0��2�p��;��D<��y���̀po߽����HBn#B��B.l�e��y;y>��EC��g���S?ȍã�#���:�e�ۡi��p}��
Gͤ��'b�.�&=�.�:��X�)�@�^�Q��T3S>�������a�WL��C�,�=�GħT��=�@����1�
˪�|���e8��I+�8+ǉ���� 6I��x:b�_w���ěGmp�8�9(�d� ���Y+�����tIa�'<W�)�L'!\��|��b>j�7��t��h�ΓA����L�Y���/�"��BK��V�$OU�P4Ôz�J����/|3�OI�a��#��	M��iGX���'���R�xx��n�fbu��j��Y�%�i�r\C�ڮR���1J�X\'�E��HŘ�����~���&���U��C>���f��fN��xf��W���[|�'Ȯ@x�E��W��/�����br��v&,�'���/�+)<w�:�ݯU���
�	*�7>��Uhh�,���I��	�b��]�������Yʏ��g��ur�lz���}͙YI*�tA�z�Q��7��)�So)qЍ�q�EB"B��q�tc����(ǈ������Q��Za�7�ͩN2���K����i&k�8�jd:4������4�!R�0����m�W�F�v��7Lv莁��<��K�i�}P��i��%}Ψp��u3��^.��Ђ���Eu���h> �U�ΏI��K>ު�O�#ԊY�eͤ�jk���R�u�T���Ɯ{�r���c1G%����7�p¥3C�Ev�����Tѡ�s4�&�T�k	���%pWĮ(b�)������_��z#2�9Sԅ�l8p���P�~-�їd|�G�4�+*���]��'b֠q�ٛ��HXTNK<��z=��I�b����YǜM��C���)�վq�0@BV
G;��'ߌ���y_$�	��Z窸�"��Y�p'�F5� �|�C�k*ڼ7���ŧ�7~c���W�1��-����4l��j%X{�oqi���댧�k�!9[��(�{�p���h#72E���c~B� nVS^�\n���"�s�>���{.��u$���![�>�"8�ì|X|u��Wz&�����
g�EOJ/�r;3�����W����@u/���c�����H^���N��rAJ���Z���asHM�ÛX��Z�� $c��'<mef�m��!��϶Ԉ�i��g�l�����Y��,�y�3#���D};^��J�`:v �U�e�"���!���R�:V��un�S��&�gU���.�ٚ�>gx�joz��q� Ud;Q�b�B��cB��1��{��Sϔ�<��a���06��'��P��[V��ЏU��?��"@�b��[ j�@�-Pz+�9� �����ߐGzhL�H�8v8+�D���.>�r��1��:�؇��ճ2�a�9L}��Q�jd(�˙wYnb��ᤡ����'"5|�<���3L��?G$ܿ-uBg�9�]�"Be��[���&$;b�n~��V��h~��ɬ��q7��J��I�('f?�5D��sC��=���&����D��𵏾��l���n6�����k����F�gw���r�~|1O�J��n�S�^�uvkQ����u�K�l�79m��;Ղ}.�=�'Y��]��q����%���*��t3DM�Fj~<��B4�S��L��������p�v{�+�����3�Oׅ��;E��?ҳ��rQ<4�F�D����TϧX"q����b���Ů�.��6��ͺ\1]��qb�Rxi����RZ[w��1[��]�۸������\�7�!k��{Jm$���� 뜄�Wh�17�#m'�7ψ?6k�	��W�c�� �ȃocr�'�j�&O����32�k���\k*QL����<�h�j���:3��CZZ��s�2ڝ�\*Ub_����
4%Ť\KԀƖ7-�� �U��ڈ��v5�M�fF�� ����v� ���V��9�+���Q���HH��:��4d
y��5t`���$��V���5����7W(�g�4�#Mlأ^�c�*�uB�]!2�V%_��x��
�;a���l������Cf��1��������{Y��>��t~Մy�I��;D�y���v����;�]�b/)��Q8��bJ�j`��<��)��i���5\�.T>u��n��3wԪ�O�W��5�/X�C�ض��L�in\�A����	iA�L�����R	�m�\�V�iIdot5l����]ͺ�"���4U-��%k�Q�BȀ9[��n��V���]��E
1��9���=:�At����=��+�ډ�15�
E|ђ�{����q�'3����yZ1oN�^ G��
����7.Q��t�	N9��Z� ���v���8w�@��	��í�^�6����E��-���K(W*M�c"�qQ��/2����'��?"��1ML)8�R�����P����<��&؁�ۍ��HBN@nJhٕ�d"M,z�JU�O���4���Sj�9K6�	�!&�9q�N1���dk�q�����I-��ˣ���R��?". 5��1+�:�9$G�EEK�,;��eW~KV:R�,��q������Vh�e�s6��aK��2�щTm#EH��tn�B��}O��LUn��(�y@���Zr�����"��W䤥^�4�����W�#lLJ���6���j��!Bۣ/Pf������GrE%����!*Y�ֽ�1	��=��y>�@��.�|���[Y�g&A2S(��P���kq���%��7�[|�ӟ�����	��"$ȭ#h��w��Jda���5��깘K����B34^ZR�d4Dj�Ѭ
�A�z���э(o���Jj�5�)�1'<X���<�!/�(�5�¶G��S�;�4c�B,�<f���ꪞG!��To�F��=V��v�s�A�mGj�׋��nO�ȀMG�������*$����� `nJnn���-��hu���f:�d��|	��h!�.䟫�,�g|������R}�lה
{F��	�9�:��������l�(�.�*�r�].������8%�� ��w��̡7� �	άFW�/\����>���
��}G���<�X���/� �"�`|y(����>�U�b�.�	F��[�F2�k�����-����]A�/�{^�N�6O���;C�Q��A1Z��/��əD &�#U �e�����%9�Z�ǉYV�����R�do�;[����ņ���׹C4�瀹�M�0H�_Jݲ/����K��<z�뿗]�*���9h�������uH�8E�V��\�<�#�� �NZ�P�}��P	'
���1��!�w�+��Hq��3>�� �Gd�&��:��d�|����8r5�?5�D��(�@�8�:���tW��iߐ�dD
Uv�4"���{��B 5ئp���N$2�e@<M{�xD��R�Kw��*���N�ѹ�R� x��)��1�#=���\9;0���'�>�������+���H��-����-O�%�:�Y�cҢ���N0i��suZ�ceղs��!H�y��� b!#����#M�Հ�3����b����D���y��^R�
z^O��"��ð;f�ї�/���Q�
��>k�6_����a������C��T�2U�>�����u3	���G�J�b��
�;�ѣ�\�N�$�����	��"�/;4N�z,�;�w"��=��@�/X5�%'W(���a�24�nE~_N�҂3#(2��I
DGe;E��̣� Tp�[hϖ��b��Ww���ֺxW����m���[��%��2E�ˀo�5k�F#k��q�?E��
��	r֋$Y�<�U��ՙ�N�����2�R~|3��k�PTy��BPV�z�'	�V5[��;�
����j+���DhC�y�C��_�B��sz���y�{'`�Qc��7�X?��X�E����p�
��+(W���#�|s(C�v����t�����P�_�|�m�cDn���Q4n�rb��%�.7Ͷlc�>' �x4 =`�VL�4�:g{<$!-��}�� K�%0�a��B�cy	��|"B�z�i߶鰧}�K
���'���F���aq�-�ƙ��}�L��n2PV���*��R���fJ�D���d�R�,Z���e-�x��@�y3����A�թ�E�o�8�l��B�˗�����A�`��g=̲yݠ�����!�G�$��L�HP%����0淐�+[�@��|��jo~?>�A�Z��q~5a��&��u��*�_���,oM���$��d��g��׻��w]�s�/D���ݟ+|���7��7��	a^�Z��[��_d[�2Nr��e�)�Ϊ �큑��+-��-�N����is>` ����ªs]ħ6��B�C̵�ϰ�K��m��J��?O�W�dj^��&�H�@X�PR��u�oN���da��H�LkNx<����k
D�M�T|x̯����,��>�>i	%�B�t�ړj��G���m'�����*ld����5�H�?��ħ�j�U�
T���5���Ɏ8.(��8�A7o�qo��l�L�H���y�p�@���HHV�'ؑ�n�F�s�l��ryX�D�;�թp�x�^��P�,5:��8s�鳗N�v����g��I�Բ�|,Dj'��t׆���H�bC!��g=Ua�?��l|7w��B�ѕ�n�_T5�.�dS�d�v�����L>%���'������> �g򏢰��R��e���ލ��	�qp�{z��J6�E�P�-f�C��?
�q_2I��ݔ�Uı��/,}���)�\e|���D{kE�-*G���PQG鍮utrn��Kޫ��5�	X1��k9c��t�`<k��jB���k� &kb�|`X�"�_��Ffx�k�y8��1���ߝ��t���fJ��	ɗ�dzs��p�~�z�����?'Y�m��~�N�)x�����`�5m�8B�]�/=�Pf�cX>�&H���^���X[�	�G�[��SS��o~
���^t�ֱأ�Q7���;��zy�b�r��;P�
���}Ɏ})��&$�z^���U�i��?b�c����w:A$��Z� 8
YiǤi�ʊk#����T��mt:�+S�)T�g��X5���՚.�#i�Q�>��;kZ�����˵(`>	��������qͼrj֢�d�Y��� jW���n^����(�:���=��<����'����n�u��0���1]�W�ub�X@�����e�jg����k���v$Rv]��d�|���<�Γ=)�j�4f~ɀ��e�C���4*���ס6'��=/f��!^�TMN�Ԛ�X�\��e5�^�#<'iekqn^�D��b�W��k�Ы}��7κ�f���'l�'��?K?`�;�����kG�l�=���9�~�~��Z��4�G�J\�>�J��ߐ7�D���K�m�I��Pu�O�����uL�����*��E�;^�e�����G(�Fڡ�� \pʹ�/���S�ʹƪ�e��g� A�9[a屷��~�D|���t\4��%�+_�!j(���� @�+�WU9����kq�`�t��M益o�	i����o?�^��Ϻo��,�9�F�Z���<�����X�V2e����3��T�f>�4A�y�b��x���Ƣ��Y��\�l�3]4��W.�U�u��ʕ[��z1j!3���_�¶'������~rA�.�	��P��Z�9�g�ݸ/�@���V ���1�Dw�f9E@��̵�% �4��^!�^�.��}]���ȵ)'"���1
�d������؎S���A���js��>/m����YLSA;C���x���U��
�l���3���d\�Y�#%$�������a�������I��%u��(B�����$@F���P=lZИP8�S��		48JiN�n
��:��`kl0ʱ�m���Ar����B�NW��*?��^ϻ�"�h�����k����1y�ie7-��6At��#|E`t�Xz�����*Ru��E�N5&?�Ȣ�(��Ч�_��?`P4a��Y�ҫ����e�h0�
��B�S��6��ر��H��[�=��.����;���:Hi��J����$���zLVD�mO.#0TJJ0%�A�u"����,��?�@�-�#GG�;�3��5#G��cڭ��tq]k+r�ɕ����$�ͬQ���ƛ�<���P�޺�T3�Co*����N��9B�i	�]�"\š�y<�H�J���l���:`ㅴ#����n��Я��w�e��c���@:ˆ
4'��hW%f��8tu�ߐ�f��� ����ُ寽��3�-�����Nȿ
1]k� ��WV�;��9����s�x<'�+S}T/�y91�y�ZW�phJx�����]��*A�"�C1,�����<a��ү��*Q"�!��Oifa.Fx,�D����x]b族ٚ
�نԅv��������ǽ��9h�^��n��w�_P� �I�jL��8nd��,���g�Nd-�w��b�\�洽 ����bvڔ����V5���h�;\kn�w�0L�'���`��DNICQ�;��l]��:Y��f���,�|���z�:E���ǔfN�}f�5|�r6R�)����oF�Dʫg���a�S�EY6�&��uD-�52���Dxs���M��h�h�v����A��f,C�>p���+B�E\X%�)���zG�ôH<�C�\g�{�i���d_�@��L�yݕ�<�}=o���ge#Ӿ_������i��ǑN;��~v���Ia�_KW�<���I#ho]pv[>�=
�!� .$~?�rΰ�B���_����n}xK~�)�[f�5RV�ۋ5�&8^�k���jw���	z�Tq|��}T,MA|%�G����_�4_�(�ݢ;�r��>nG�lP|�ef�N�^��}����C�tt��^�}��xBn�C<B��0+��'B����Z$ �3k.�5�G�>��x���T-Qj-P��������=ۼxmt#�������e�h���9��(>��U�D�i�0�S*�6�����P�g2��Z!F�G<�� �x�FT�b��$�澑�u��<��\!]��1'"�ΏҮEL�j���O�X�IQ���X�7����H��v��śĄl2�t/���o��e� �P#����Z����{s��b�����/�>��}�񡏘3�
&Z�g���^����m3z֥h�s�����(Ģ���� I�P)�#B�CƜ�:%_���l��P��l+��R9�NO��)��ܟ�p)�I6�[������X1f��;�/��?�����c~ƻ�$�!T�Z���G^	}��y�-�:���w,��=�aW�C���oI��1��� {���Yjʝָ�
�<��*f����W��.?~��Уpw�=a7�p�) �j���|�6�z:�����C���w/�I�g����OJf�è�"�생��W>��S��Ց��WEc�q&��]y���t��`ץH���*Q
	U5�i��w(��0�7_��M�Z���W�N�3oX@xZ`�v �~�[ç�n!�~�S���hjP��g�}���,D?{�����k:*xk���Àˍ�d��۵���I��p���3=zT���cqU��yy�9��Nl��p���,aca���P��#	���&�e+@՛2����� �A��i��ࠀx�{Xni��zo0r�
�ݡ�h2��R!g���)kp�<�A]�"�9���i�:!����]"�=�i˔�OV, ]����|V6���]'>��%��Cߛ����NI���$����w�A��v��@�ҧΔ�j��`D�: ��Ilz����$ß�l]�F?��[��Iπ� Nā�`	B��j���Ӏ��Zמ��n�,z�Hڼ��B�|�`�&Д��s�u_J{���g�8����眛�
Y����0�C;��Άuc�.��(�N��8r�#�4�/E;YT /�oa�2:�"<5��뿖',���������SO�J����i����bn��.,,fH��Zg-	�\>J�n�A5���S:ш҅y=�����!�/�� ��ۈ~G��̷	3�x���a��t��n�i��2"f��"~�!>�q7�tªz+����A���z5x��p�����[d\�=z#�-}w*ŽR5� �1�;u+����-*�νA���}_�Jp9��`��G7M��I��D��!}�����獽4�IZ���u9j����W�B��s:~{�%�ӹeK��@�'&���z5
��z2&���~3��7��XMIeݪ�wmt�Þ:�c���[S������=����83_��{��q��D�Ԭa�pR�]��{���S�V��78�<�.��������__�HQ�mݱQ=�=���������9��m�C�X3�u�͗r�bOĭ���M=1`˭]f&�@�cT�^�,�~�`-1N�2n%F����|����P���b���?(�awMاF����.h����-�ޫ�C�������s���^���kXH��4q���{���9�3O�����Dm��xo�ꯉ�PM$�>�s�d�jӘ'aZ�5��/v�ݱ��F�,e�6�\��[0*�����:�ݎ�:�/�j���NU`@h��<��&���6D�#h��w�EC��S�t���|�Y���P&g�i��axuJ�du߬x�c~�X�?H�V��q
4ұ���äoz����n��7�wg�(�e'�D�_>Ǥ� �����e�pK�,7�.�������0) �ؼnX�օfN�@rh�D�v��p�����G:�ͺx�ӈ�Qѝ���+낞;ߡ���!%RK�����0�(��/Gj�1�.�(�Ϥ(K�/<���W���|ni%�ݍv�2=�μ�'���]<�c�	ח�\Rr7�XQ`�O��FdDϵ�ҁ\qQ5��6WU��%�|̓[�3�N1,�J��섍Lݩ���Ѯ�w�BRy������#|��E�y�7�K��� �d	t3Oqo�
�z��re�,��M�Ս¨�!�����/��pb�	-�Ni�������桄:�p�$�:��c�T��]��2�\5�:�uVR�A^��A���D�V;|Mŏ.ۙU�Wge>�m\���<n�k��:m-�2j\�[|k����=�+�%����5�3`. ʹi��K�.P��g%Kˡ��(��Z�Hpy�C�Y��$�!�m�$�S04����pa��	��*}%����O�A'�#pGQ��,�!&rQ�Z���o_���3��J��v`���3R ����ݰ�Q����w.����.�CB4ޯS����PTWO�D����.�������6�����{_����p��`��ǡV��U� ��m�g��/Ȭ8;Xځjz���C��w���g6H<�abB;�3��<�a��b�ш!�	��#�!��5I�F�wq� �d$���Z��n&丳��s|�<�t���1���lql�ѯ��=A����&��ZQ���v��i�Qe	�\�e��^�)�"q���^@&ȩ1����K�]�]��ڂ��M�����\��pS-뽡-�e���	'�[h���:�ٻ�͏pj��rCKR��T�`�j��OR�����d���˼�8��5�^; ��-��T�a�`M�Q: Hɻ�샗|^�Z<�/2��f�|�@�õTP�����<�@^�k�����7�G���э���c�+�W5��H���j��N9�;�˔ʓb�X�GMlAjsd�&�|��"�	n�-�:Mc�7��*=o�N�ȑ���X�
�#���+����,����"�oHi���V� �a-������X#�Ʀ�Ze�Qy4]����#�`g�a��?q��J{��N�Ք�զ���P���xZ��[U�!Z��|&��Q�3eٓ��A�A�5�T���瓤,���-=�
u��ɞ+}�[2A��u3��8S����7}���d��,���O�wщ��S3\c2#� G���Q).�r�]J#��s�D]��� g�������K���6PJ隫������}P���#�Q�Gx��BM'R����5�z���e�5n�>�t�K.���I���ڙ�-eRzd�Do�V�>D�qB���a��;��V�VH�[�a~�L��?M �L��tz�I��-�X���O�r���A��;H�n�_Obbi5�����&G�7�ˣ�V��s��_�F�uM��� �V3��`~U���9R���i����WY� #��B�hB��C����\��^b��DrO�R�w�������b�wĶlFn~����Nl��vm~HF�j;�$��Sk�["+�0,�̛µ�$�3�g�,v]c��յ/6Zd���6m&�DAy�\���1K��#�c�f��:2B�-�Liz�b�����L�>^�QX�"�X���'7�w3|MH��*��#0E` �VHZ""ݡ�d0C��F(} �7�g{۫�Ӝ>�a�yc7�槨��H[��@���tV��tD�B�[�oֆ+�R��]�(F'ӫ�=�0uf�|񐷜�PS%��s���}a<����nmVA��(��[s�[�3����[	��y�4Ԝ5��M�!"�
�O|.����}#�����z(aD�w�������׫�O6]FD��]�۴y�	G�_q`�/��fE�t�Ƙ�I�h���� nېm\ǀ�{u�$�޿H3��W�]E��E�+�T1r��U=&9���H��7�=�Wl���_�4���������g�*�-~��@��&)s�������-�5	%�M"�!��m��ғ�k�#?[�BX�eS�e���d���)0�)�b��O�72F���D�9(]^�FMK���Tj�)J !�����H6�<e�e�ZFV�8���c���$�������5��uH�Z0k_7y��L��>����Xw��y�Lc�6�P��?L���`��F|�j���a%N�Wپ��/��y+�'VʿT&�4��$�ۉ�(.�Ϻ�rֻV5���3�54z��tn�"w��ËqĆR_����D���~:�y�^��%[��z�����R3�b���j��3�I�_S&���J���,8Pۻw�ҳi$:��g||�Y�e+rc"��6l�iOb6����Q��	+��$+p[S�_ЃN;���`���4��B���]噛HU�f���#Ύ1�p��a���qa*���*����~��l��j�^�����}�>�c�K�� �>rP��)$'��q'�#����U���ڻ�\Q�0<��>�eP���הB
�s����>Td�� ����h�
@ R�Y5�K��[M	@� d׋G_�Pel	���>�F.륗��p5O�K�R
�7Vi�e���ĕ�ޣa`ȬA ���lp�Υ���k�u�
4��y_��h.Zz̏��O�Qth��|*��j������<�旿t����C�� ;���_ś���#�S�0-�s�G�2�Ծ��leXj�����c  pK�D����̖Q�S�7��0���,��*T7���4eI�˶���%�:�e�s_�=�g`|���ۃ;�:���
V����`S�ԗo �Y#U��F��7�o7��I�;�~��ӆJ�Ʌ!O8EL
!��8�01�5�<�%����imB���D�V��8:A�'�qh��l�Q%)�#�J��(�ODQy&��^e�,��ʬ �q%��_��X����!@5W?ԏr&&����)0(X�~���~�R}A��z�$-$�9��@�,�:���Q�Q;gejt� �[ɾ��.�k�
6�ح��H�U��mM�	Y�.}̢0�����ik���(�}&�&b��{�|@��a� �Jtp6��2�����r1T��@E�԰��x�X�ڔ����'B\�V8>��0��g:��s67�+B让��Si�Hs�]���,�a��ME<ڢ�%�-����������C��2#Mr#*�<�4�鎜%�Jf�`�1�NP�C�^�@�W��Q%@��i�C�Q�.j�X9�3�"��Fq'qz�����f��2�}�%M阙ȚsE���F���is҉=3��J����{H�Ȋ�w	k��ښY3�	��[ίV�NXg��JrS����ޝ�%���E�-<����˨�ЂN��O7�;��Z�o�E�F���%����@����sK��>g-z�(N-8��7�e���7gT�w�ƭP����4-ى��7�xf�W�t;7��A}B>@~�idʢ�?��	Yh�Cs9p�ˀ`l
˹0���!���(d)p�\�J���CC�x��f�!<�h�Q|)bU��>B�˝�Nm�8��G��Ic_Q�\'�7�P�W��L��p�j�"���!��h�����X��+��}�b���/>�S��>�7����?�4XI��.��}r¢�������^��,i@R�����1'\��0S���T�����L�F��9R���C�d
�� ׈�fmN0�r��Ц%��a���e��YLY�263&@2�Ĝ$�8:�\�k��dؐ�mt!{�p2��	P�5�wf��J4�ϓ�,���<DM�"h��R���.�դ}�J"s4�M
�n�#��_�6��<����|��-\P�!��E��~`�'�?{!6K[����#����rhu d~��W��1��aQ�Ԓ'�q���&p��ˍ�wQ�V| ��6k�c4���+8��%"���k��<��j��3����Y�}G0fy��x�U���x{�Y��N�ퟶ�b��d��0�Ε���X�����W&,�L�ad�ި�y���+���;B|�뜖e��2fU�T��)p�v��*O�
Dt"���"�� �V<���_lS��J\uH-�P�2G�+���6��x4�awL��a��!�#7�KE-�@��٨:2��lc|-}{��߾3~�ؠ}@����T����"�g	����ݬ�Ԃ9�~�o��N���O�}�(�;��Op[w��A�[�S�[�#59���Q&��I��ƍ ;Nĵcw���D3����H�#�Ԑ��հǼKT}���v��a���.�Ut[_�,�]p{S�n��eyM���U�৹k��uI��� ^����]��nO���3�9ի2� �(�'�ȯ����*I��#�|!2��W|��,&���`1ߏ�t[��4��~��]G�K�ޮ}z��p��k�`���T�{�(�SE�$.�2h��&`�/H�3�޶�����aKr�����ȗ+����W��U����|������	�z.��r'D]��3��V�!�tn�D��bw�
\���f37�@5'��@�Y�����}ڢ�g�(��b���X����eZ�ޮW��͌�;���S�J�[V�K˔
����3��	��2�KN�a�2�����։Z���3	���"Y��\��H '= �3�_lߌf��_�!�o�*��MSt)�^��hOpC���q:���_��C���ל�z�h���Y�1�����D z+�=�;k���T��j����/׊��#��o����Y�V-]�G
�?��J�$��o!h�����m@�V�?���g�g������Z��� ��0&H'E(k��R��4��
�;�#A�P[g�:��k�"��.�*��O����W������b�\B	��[kY�:>t�
�+�J7�g�5dqe�Re,
�&FX���ܻt�$�>�m��� �]1����*���~D��*�Es_��33���{�É��\6�'#4�C���:BY'��Ψ���N{��
�j����a����x�kD����Ĭ��e���9j�����ب�?v�O�^]�=֓ϙ��@�d�7�/�3H���.X�N^b�JdB�rOk�<�l�n"ǲ!v�E?���U-ջsG���hS�Tc����V۬n�g���F@B���w7� G��+���阝 �.}y#i!��_�%<B�r�/�^�
:J2MJu0��E�=����aG�	��S�l"��s�*k�vJ�V�y�m;�<�$�X��pRL�j��e�$��(ŬgF�|�@�З[�4O��Y�,`�
�{S���;9���	6ҫQ���Eo�G��R��ů@QD����=(�i��\aC��{�=C��3�(���uV���'��\����ՊRrQ$GLR���
���S�O"-7�P�@ ������yzHQ�me�r����h��J!i{g��7���/3-z���@�!���>1�ee\����7.����ǵT(�$��I2����� ���=uv���s�R�����`�J��T<�a�=]��:i�uYm;w�W�!�e�'�Ȝ�Pl���5x���駝��������-=�gR�x�*Œ+qE��G�fQKa2k���)�������������uG1��2Q�YB�r2�0")D��@�㵌Y(�$�w��nK�2[����Y��=YH��96�|��1:��J4�}&(����nd�f�&Y��@��_��2�!c�w?L&�6%�Ag�,} ��H&f;`��f�f��/m�M�񧁿��lR�w�l���똍���7��Y`y���^�L{Z�)�a��%��}�R��X�Ezlq;��
�B�]�n2���[c��6]sCJ�!�g��P��� �r�e�/�½E�,�h��B�Wr%)*E�Dć� �T�~A7{xX�4������iz�η?m����/.]�9��6RZ�>��H��*4�����ɕ��\�vݒ1��\?<F���
g��T�y���n�$W��������X�b>0����^�+r��M��8 I���6�����n�����Pqh��8���`�ّm���L�ƥ�
�˥�� F��l�
�uO������/|*P�rIl�t*����S��7�����E�$�[`)i׿d}�J���l�~�Dg)jԑ�7�9���v�'$O�%�u��2���=���̲����b��S����V�l_����_g�;9ðZ�	b���?
b`Uu|�h������+�TxpzQ:�oWޜ�!z�����\2���)Tz�c8�{~Gk�ߍ���*����`þ���Q�s�@U9�XkP��鈚��un�4T������~r���&��(�)SG�UF_�\�ۏ�+��枻b_3�ޭҽ�N���h����yl�(��* y{��L��=����=w��<.���KO�<U�9�߇5�P��ɨ�m:��&���I���t��Ҙ�����`|��flÚ��{GFT쭐����2��39*-�)BZ���1n�*����4{4���L�99܍�޳P�V��
ӆ��	HQ�J@8�jP��̑��/-�|u�|_K!��h����%��òl��Ƿ|E�]��צ�Mu�1��Z?RH��̓�CS�O���->\"#o���B�ta?�T�7v��1��_E2G�/���S���s�H��S���q��4�I�q�Gޝ���bFZO�E�0#'�/�r�����j)I�T���a{���6�<c�;�a\�_�vh���jY	0=�!ɸ��,���y3�$�>�0�N�Jp� �J5��q�ա�C�S�%��r��gf�kI�������π�+���?�)6�3�E��J���E���B��X�g]�Dn��d�F�����jC�\M�n�V�9����t8��n�<�MGu�
��d�
�|S퉾��c�.@x�_O����`շ`Y���.`�X��Rѽ?�l�(E���>�P�
]�Ȉc5�[��E�R�̷7�Zi��b��-�g%��/�RZg-��vɷ�ԐT4ݾ$�;�Z{Й��d,��eJ|�K|��Y��W���3��5.�m�=&9!�Z6�F�~<��!A��*?��%��yS9),O�њ�TID=�]��>�#�������s˻���Ѱd�B?�x����0[í/+$�W�k�O���(�8��K�6�*D�T��)J�|�T�Ay�:�$��4L��e��.���2�L{�P�)�%��4O\��0�xh��v���<�xT�Qo�}@~��~��t嵤BoO�ܱ#�1W��5^@[/!��Hq�*�"�8��Zy��;"W'�J;��gA럿v����٢>�"���8��YnMmp�z��������H9�ƨM)2��r�jK��'S�Vdѹyق,vX�p��W}��+OXq�B��32Z["�\3���3_jU�v6��ZG#�*�2��9VC����p[�4J��UB��p��4,�+i������mv���:Jdj_�e`5�q���tЍ9@����N�Ik����V�Mw�hȁÂSް�L��
'��DY�����>��K|8�/Ut.��S��b#vW�R[5�]Ƚ���7٧�N�/��H��V��4h|�bd���y�]*�]�BH"�O{�2�y�!\�.۲��+���>���-���x�5��-3�o�H�y��m|�	��$��k��?k�`r&�	h���ѐQ��?���RR0��sX�uJtC0�~�kv�d$OVJ�]���"�pzY�B�կ���N&�au�S���6�s&�A�fS�̦/�3+t*�泣�co=��-�����Ư���� bH*�	�p���H�	"���ٱ/�0<D���,�+C_"n���:ٜ�75�f!eo�!�� ʱ#W�8��iBl�Lr�#$,������lh*�b�����b�:e@��$�Xe9�T0:��?IT�6��P�XI��xe�� �M7�6v3?YZ
ԑ�8g��b�d�6(��p�\;�T�,:�s���`v1�e�V��S3"�h5����t�<=hĩӷ��=����|<yz&���>��4�yv�c3cA���0)��S[&b�S�]�])�ץ������o�S9�ć��r���J��vunΰ��|��R���ٶ�gDS��R�����F�R��5�Ҳ ����9i�$��AR��RJ̜4�su�w#H��~<�Z�w�5si�S[gp�e�0��7������9���|t��A��h�t�h������O���d���x�0���^">陃LJ���ę�ϛgI�+n��A�؄fS�q-��kS��.GN�1gKܲm���q�x���)�r(�lVGK�$��M�6�Et��E1��5��'�&SD E��/t�7��B���xS�C�.o�_߸x�U�z�\R��{��#n&�7�F�E}7���5gm�6�������4K7=����\�"�3�D9����1�]�ȥ��2#��G1�34��yF��8����i�Q��tY����I���-f9Gq1u�l+>
�N��Y ����KK>��1�ZUg�f�12�Kq���D�+�ܟ9��g����2�7Eg�����u�^ôP��M��^G�j[Q�}M&�i�g��y:�ػ��W!�q�]���p�[9����d�}�V���#��Ȼ�;V��̟��_��g�v��A�L��je�_{L�I1Ay|%�`y��E�[,�7���-�������sDYs�ÛD.Uȱl��)�U(�k�!��,Cr;p.���)ˡmW�Y��\���yE��d�]/����O���0v�����:�׿���)�j��^�[���w�2�dew���8�����>�-=S	7(�6Ȣ&F*�c���>��&�h����c�3�PzZ6&�m�;��T���x��_�.To�h�PC�8J,�|U�K:�C`�Z/���D5��8AN������B7Kv�1OTe,#c�9��>���ʌug���E��X���$Ruzy
>���T��B>�߬G<_��4o�`�|�v�i�Wm��پ�(U�3r!o9XiV�.����¾1ǋ!���_�#3ҭ���B	��ܵv�k����%A4�+�	��'B�'�c�d�g�q�zh���H�7 �i�x�8�ڦ �``Mך+ ��S$�x����x��U����]n��Ϸ(��{ᛜ!��ٰ�}����(�4���)��)�}P6O�3����`ò�Y�u J�Y��'��S��
	]�7���K�)�
kEm�}��;�o^�7�k��&�=��ϰ-�}
(0��E�jG��G����Hm��v����0e�є�?/^��>���&iub��{�_U5�k�xzc�nI cEC'%pD�(��r����x�����]�r  #C0���m��d����RD�>G�&��Q����ެ��G�j� �Jᬨ�0i#J����sK��\J�l���27H��R������k @x�ܯ�!�v�h-zz����^Y\�9h��I�էsN��u������d�t�ەcw�~@�^� �y˲��:������a�
���f7�~���cp@���j/L~KH-�L�(��bV��QÛ��v\���A3;��1+��n��'���1q����¾��h��R:il�"2vC�D����`<{5/=֏���*(�o6���-&���M1�d�5�?�@y`T����}�_�
�X9I=w�eۭ�t��]Ɣi��ŗI�ëC���7��l=g�y-�j\۬����7�����R���W���_�T�7>�|�� ���L���~Q٧��mt��v^1f7�jg<���8ʢGd��nک���B���T���J��3�
 ������٥��TV@��2��_�d^��7+@����=��cJ7�����eI�K|,2�S�6:��PP���y�~?d��|a!Hi i��i휗B�T�5 ͩ᷼vYw��j���s�GA��k!SN�>^O`�+4����V�E^h���MLTAW�~'>K�$!.4)��	+؆�� Mr^��.y�*A����32Ǟs�)���J��Sf`�ՠVm=@��Ӣ�$���iO8>Fv�qF4o�����J���gs~����� �h�m��W��<㞲w:��QyxH
,# ���/Qn<�1�7J��b]��jR	������ik�[	�:�E��V#*���|�����"��1{�	�Z����z��+9�C���|��Ӊl�0-�\ƌ��5��JO9�k($�%�իQ�>�fw�
�0P;��< ��8M�]YV-x��70	O��u���s��7���KͰ9��J�XBJ�>
X��j�x�r��2�KIC��KQj������ Iޛ ~�N�np�нZ���
��i��ȷ)�v[[ǔ�t�a�_@D��"�}�.�4���;}
V��0�`��,���殞�]z�]*`0����
B*�m���ܪ�Lsy��F��c�(yԓp\L������Y�&�nf�Mͻ�3�m7c�?�T�}�����/zb��O��|B�b��<�h����3[V��'�p9.3�s�)��)ͯ=0����$z�I����g�|�/y�\k��z���xX�F���L`��PG���:�(�l�?��'�
�x�l�:
~c�f!(���ʮ�{�d*�fm�A·��A����Ѿ!�u5�5�(ic�ϥ��������13Π�F�����,�����o�P|5L~�ag[����Y9�X��6�FA�`3O#��/Ni(P��殗y��¸�����X�NN�������/��gM�umrl�!ô��@6X7q:��V3�t$82��UJ��U־IBP���i�I��������FJf���Jr?�9�!����
g^�s�0F�tw-5��~����2�q)l�Y�vVX�8��I����@�\7~Q�0[�Ai���86�%����i4�e�|J2UQ6j\�}�;���͙�}[����(�*\���D���s�<D���+C�=���oסi�(l�i�Y���WA�/Mo5�G�eB�6�����<��%��'k�A��!�=+�u�}�Ӫ��w �^(�}|��_�А_47��l�f�d§;�9�i�����tr0�A�En��k����­6�C'�pB�W������R�J^@��GvIb��R�p�o�EH����2�|d�Å��	Yv� x2&D�k6�t���!���S�n�ʰ����9��8pYC�8�`tٲ�yؾ��XE9���]�:+d���1�+y~���y99��	v�Cq�$oX�/�`��y|�ֲ��bE�4F�v���g8K֏�i��؁�Ϲ����L�Zq���B�8ן��i��p��vb���z6A�[��p�.&{ � ʝ�<��N����w'=0;���U\�k�v.P�7�	�{Ӹ��<e
�t˛d��@��+G��	O�w_k5�-g��6�h�>���������zk�#J�=bWjG���#ηNUFTüG�gh=�j���L����.�LpK�I��3"L��(|c� h�R�:T*r�Ƅd�ea.�v �������U��>a�6�䏷V�u�_`�������r�t<B�5�=����xyhS�_2.]��id+������6K�D%���h�t� H��s�@�*!�lG~-:1���Fms��j�>Ǆ>L`�c_���nJ!A���()���W�'e���%�X��M�9���KD�j���t���
�D!��w��쀡��Ī�w���	K�=%.�_dz���%�G�����R���+#�c�TBj�O��U�~����7�C���^���"kWg�t�>���e���0�	�Dd��MR<�.����"[�DF,�)}X��Ryʒ�.xFr3���y���Ȳ
�\����z���? �� 	ޒ1��,I�;���:X�\�~U�)�������N,����~ �A�i����m��VJ���q+@�[�s\�k�6��W����O�5���(,�7�C{�c����]���=�C�:���V齭���щ���O���jYoN����=���������K���C�3�we��������7�mHѩ����u$�Y��3�h5Ѣ�a9�Ɨ\ys����|j	n�R��o#J�y2�"T�W���1��g�	cMog=���N�Y�NM�Zk(�i0��&e��~{+FEź��#0C�ipjI�������#O&ď�)� 2��v�O����`�'֬��8s��U��vG[��[׻�<�AmC0��ۈ?�d�Z�C����D�z+&��8J��GV��솠
x�/{/�f�s�>꽦����elC�W:n�#���!��,5b�S��f��+Ʉ��X,�0+m}>��T�Rg�����d�g_@I�)N�;S6Ȭ�gr�,��#\��7�LFۊM,��U��o�0>v>�TĴ�
U��F�kc�<-"��O�0��%-���:s�F���q�{�n�Ƈ�_�\{���'���J�Rkj:��"ɧ_�="�p�*�D垾ֱ:�|
N�3�Y���*|�i0��	�kg�`��uR��̇����Oir�3�1����˵��:�����nʪ��3����n/�Q���
z��;Y��.����hh����K)E�#�osV�KE���,��4�׏S�e��4�x���������F'*Ьp��j1ؖp��&g%�2��+.D�I ��c����q�ew�C�h���7�^W�=��@ 1ƻf�񹀂ds��_͸�4ubUq &�MP׍=�#��h�:�z�I�*�V_m�m�Q.#�3@wP�bTvqd��8ގL���[�0�h_����2�L*6���D�����=��Vnc��<�:h�a��C!��S���'Rv	Ӊ�o_�&R�G6I.f�]�:�KSh�':ҫ��
�>*��I7ì�B��\���@< ��e�#_�`�0B�*���k�v���(C���<�y���ކ���B�6���G��_�3����</sS�r�w.r;n�x,==d� �p���L�)?�荈o��1��DsP�Eu!��b"���Vݬ80r�����]8R��o������]3�\��(ଈ��Oᠸ7x��2�hX˭�ݫ+{a�� D6�6��*9
���`K�����\����Ss�>/T���h�� @Y�U�Y^�g,��|M��-�����	�x��=]����&�䪋u�����!计�����k$�#G�9C��9��X^�����y��;���0��r�Ch@���'�س[����[uC#Fn�=UΊ�WR=��)���ud�:ML� ���:��_^�X 㬷 `t�pMi���`�Q�D|(�F��*��*���qɇ��
ݱ�wb�nh!����Nǲ����U���&p��o�m�{^>�s�G���->a�Z�4sc"�ZQ�Q%�AY]��:��~巬o6��a�BN;}]ZH�HXC����j�E�g�v����(��V��@�E���O��$Q��2)V&@c��U��xcm��
bJ��dϐP�3��:p�.~c�ų�ω6�>�������Y�HOi8����/nh
x�h����/���^�u�����ƒ�\������@�4�8��rw�����$�-#�oZɽ�M.��~9�m��ޘWS_�y_��v�o�8��誂ؑqI�uS����yD�k�3?n>}hO&5�vVzf�\U,��HU�+�\���p1��lI�NL�YESC�Ɏ���Zs��aR@��[���a�e6�`����+gt	�wB9]����I�C�������W�##[��ս�T����]@�!�Ipa�X\$�2�r��X*�-�M�#��1tP���!�>�UQ~O]�?�~ۦ.�\3KE_'�N5�n��BBNvUt����ۇ���4[�͒��B��ȴM�Pv(��'H��K�<��G��?�?�L@h�Osv��S�nm��0�J3�ʬ���q��V�N>�L�w� .�OԻ�Wh0��5�ɻ���0������MW��1�x�%I����(S�P��7g���t����9)�}A�ʫ�^�E�w)-7�S2Z?T�[_.},j�����1����,�\n>�dz�Ų�k�#>�&�������xzs��Z'�7�#I�xU���O��{�u0��@�ĳ��:l#挖�-�L��ۺS�媡б���>w)�w���Ĝz����7䀲�l�����wo�>G4�78�:���X�%���?���=���QBoP�^�)q��=D�We{���/��DxE��׵��[?ތĢ#�*�-~������ƿkB��g��Cfr+Y�7�`���h8.;o{Z6�:q3�Gy�QK�wvK3K:5��4e���x� �-��*�#Qa��&���LN�����T���	%��9�������?Hz-���NqJ�x}b	 U ���C�K��#��-�]U���o��Q���k!��`��/[��y]��� �	I�]�y�U���\�V!E(�lA�y��,'�ae���Q(	��+��%�\_�Sj�&=G���?=�	2]�����ёHV!�ʡ; �䏷�DHa�]J�Y�>���Y���d��|c�����ū_��hE�z2��_�O�=h��L�!`2�q������U����8��c����:x���4��,Sg@"��g��7��V�\�\y�Zx'm�+riXnD�wm�?��L��)4�G�}G���L���x]�{6�����#�!���yByQ��qz��F�.*�ʈna���3�[�3�Z���qyE��d^��!�x�؀6��>^�Q��k��%Luٲ��A�|��2�6�>��%�#�+wQ9~	0k��Hdتi�8�˖�Y�vqg-l��q���Q,�}6T-�BXK�"p��B��" ��f�J���q�ԍt��K5���5�øC
Ch��=/��ʞHg%k/QL��
�L=6H#�gH6(�S-�M�n��Q�%]��b�k�N�8pi��ʋ��z��{��g���"b�;�`�(ھk�oX�22p�ҥ:�`f�գrP6�����%J}K����Q���2r/�+��,�O�.jc�*�$�l��q�?�N+l��D���c��S�Hz$��~�=�@9K�N���>_:Q�BF�P@��E���l��4g���1wW�|�dx�
�.�,Ϛ�EJ�S|�� �P�J ��N[�X�yʊ����`߯:Z�˙�8����������P�@P�L��l�b���H�*�$��w���1	\���[�z�'4/=��8��߼,X��w$1�-D�Di�$6<TZ[FߚO��P�/��cP�� �6]�a��Y����I�Mp~S�vx��)��� ��<]`g��}���IJq0���-8�3�͹D'�Wm���E%n��U���U���B��P#��Z�zĢHi�կ�!�[��;�0n=��������NO�X\1CI-P$��xդ���GC��@j��,̾��ӈ+��1�ֽG���U�:�4��G#ybǳ@�YI|\��=�v��Cs�۳`��\�O�v����<�����Ol�59�O7i��֮"�\Ɂ9Υ,0i��;��o� ���(��K%��'IR��ٝ�YG3��L}���#ؠ��!�ca���������A�t�n�,)���c ����Ju���h�� �����9��h<��� W���K��y�2y�E#��Y+:��睤\�q��
�Q֐��@7}X���������F$O2�ܻ!���)w#����"ޑ�%������Ь-뤁�M`�ѝЪ|ydc��0���<;*��9�]�1����.-"O"2�J_#��ǝ�z�B�����H���?��C���θ���1Z������.����p%е:^)���d�?�_颮&�LV����#�L��bS��6�1FN��'+�H�1���Ee+a�O���tn}� ^����ܵ����_jC����&q+��3����{�?�K�˛�[8�	Y���U[^�JXF1��=j���~M>�����P�8��sŭ��{��$=Ix�WI�F�<ʝ�ğj��-(��RZ�s��K4T@�J�L��;�{��Q��}{d���������hX��$��0�^3e���4O{
A���E7���6"���P]u���&��)�L����WP��=�'y~hA�v��L\����
���k&8|��|�t ��߿
�{Rl�8l��K�dS>��PwiQ0���~.�����Z���o=a��V7C��hT&���c��W����6��cr_�qG���ɕ�,��\ŊT��_�[�a/5{`C?MlP�/�#���o�t���:6�9�ݞ�+��BmJ�K��6:#��2����
/ؚ���a?�YV���{^�x����o��i�5h���[.F0���#'��`�U<�!�gW�]�	����|�B��`1V73��lq&��f�U���N7���C�|��FD�.eOL2Q&¶���ľ7��0�L>!?L�d�n�J.��Qj�Ρ��I<��iz��q����D`���mg�}疳�zeQ��f�bL�ˑa؍|dϥ�X�W���a����;�E��B=�a�X_)���5��X��JDz���Hl�~\y�zkew�xȩ5IFex&@�(�K2��p�a�����{0�W���o�J=����W�Ǐ�����%�%��HF��Ҥ�9+Pv��dq���ʙVd��u�ڀ�����ϫ1�{C=�RL�!j�l�i�{:�Ǖ��
�1�DhJ�!h��؈:���6pV؋��'	Rq�	��2i+�Oע�q����R��vE�K�s������/��F��=�j�Rr8�q�DK�%2�P��R�"`���{�	i$�I��#e�U��HoH�Q�;�J mxy$���0�Z�*���`8+������]3�&�N�OV�>�`��׶W�����ҫ���w�<��m�bIÄ���b+� �YĆn8G@itj!�3P�#�s����`j�Z3�;Y?DAѭ�<6�g6��q�!�Ė��|E�z'�_l�9ޭ����tb{)�O�S�;��!P�����ٙw�����8�dp��(D�(nDm;�3�^U4�S;�px�~z��-ܛ��#O���gA?����:DG"�c��Ō9{�&��SL�U�q1'��+spg����!����ݽ�B��:n�Ե#p�D.�R?�)�t~q�1�8�z�խ�P������wpHT�I-~�q�5�#(*��>h�e�!	#(ay����Ԝ�i�҇���� ���\�d9:���&/�_ /xó1�I�[���B���F��F(L���ݨ-p�� �8hh�Z0zk� ��T�=b#z�]��š�<#���.z<9�36{ɱ	�bA��ؼ("�X�%������r��N����[�xn��Q�'R~�9_-˥=YD'O����u�;<�yޫ����[�@���0\PZ9�S�=ߝ��6���IUĆ�9��p=�2o� ���&��΂g�aC��.�j6��oVط��W��Y_�����t��
����c3������0��^����	T���tΘH���݀�+�V���t��X+���i}ܼ�F�s�p�R��>w��W�Xk��Lv���'��.�g��ۅR���I^,����{��B��o���*�6}���K=����v�/��<uc�5��ڈrb�2�����r��&%i�1�tz[�$��@מLʔ�ۉ�H�q�F��l߃L��ɇE��73�q�I�Ҝ�=k���sd 
.x�oK����7�9�O.����q�A�\��w��x����µ��ވ!��<�@����NWY�ܩßh;��ׯ'�;T�֊��%�1֙d�@ӭ�4Ha�����1�o�60Q����AL�5	E�l����v��k	�@�+SwZ9�~��Ls���s�50����R�°�19����Z̙��Y�:Ht�=SuH
�$�D \_���穩����YL����閴q$j ش%���Z��K��S�D�D����6̜<��� ʥ��K�4�"X^��m�CJa�J"l�JD��GY�v�l����@�ܹ�O�#���!�O��R�EJ��j���À���?'�S퀛��]�L�9@��Ù���KN؁��Μf��8���8Y�\C����õB��{��𼉛A�[���п�K�y8Z3e�}q/6g�+��� �pj㰽w��kXk�8sC��W������ܱs��Se�/�G92Й!�����ruVW���=�Z�S�V��%l�f�����ݥYK�;�c����<��6��K��=4'\�K��m��t;	�u3Q����Ə��<"��@o�:u��U�L���$�|t�<y�+���w����\:�z-�5�RGv������9P��	����Y/3���:����ԡ����A�q*5�V�F�����oZƁŶ!��� q�UC9xi��t��H�1�Ⱦ�m�J�i����3��8�B^��u����6T�M�f40.��l��&�/ �����1�<T|��܇�/s5�0
�]:��݅3җ�ظG��hk���z�����(�;j6+�g��9dv{�8~�S�Β.m�n�+�=�b�������Cߟ|2!d/p���8Ԋ�,�m�}�Xٕ7@mY��̭�<1�6�=;$�1��6z�A�8�~��j���I��Ynz�d{`��/'����>�$��bkǇ2���Z��6�kb�Uj+���k1��JH� ��¸3lk�o672�����H/q/b2y�1h�-xn��/I�y��Rݹ$LB������Np[AC�rW��'<v�� *�ls��BѤt6���!��&���m�قK9-��i�&v��{}�긯�O� ���t�t�~Y�L\"P��J�_q3,R��\B��eA1���u!cǚoK!X��UA�Z�C�e��{��.���Z�@�`7�te������x9�1�A\�Ah�/U� +�B��9�Sg��E%��D�J$7�L�9�C�
�kͳvi�!��	�'����Z��2��ң��=��(G&̬rWo�O�+�w�O��\��M[su4+��q�qk��jg�;s6���՞A���ݙ��]���?���� !K���B� �j�`��9j��l���U���m������� ��vˮ��{�����4��vۢ�,h�w^qr�cH��'yk6�"�G�B6[i3�g��So�mk���L��C��2�D���3�.;��ph�-����<V��	��Ӡ6��O&����]\��ư�ғ,�/���H}A�'p��J����B:��8�Q�'f=��LѰ�r�Q�1��b�>�u��9����CÖ {+��5��RU��I��m��y�qV���a��{^����B0�n*);�h�=G�1�6��R۵��ʒ������Dg�8ޣ��>:�N;�[���n�[�yE+�H^�����a����#k�)=��J�h���O�g���!nl4���gɭV�ƌ�UgL�a{s\����y�U�m�5���\�5��"�D-��l���ƦH������/!N�����ѻ��^ͦ?g�3���F����U@I�Xl��x��o
���bY�S�jm��!���)��x�����3T��8��=se���!�e@F�..'��e�cIc��I�ٽ����(i��� ~���YI�F�Z��tZN*�0{�}��.�����1R��{��	`4�f d���D{3�>rT��S����&?��^b+���4*-ļ�A�R� �����`8��Q�Is&f�=�p����<F��u���zOz�GՖ������B0K�C��C�]�4��;;4+�n������?�@%�z�ܩ������ֽ�u�#Mrso���$W�9�m��ViU�co��r�D֦u8�����q?9�dAA1�<&���rT�g:P���k����Vz=�#ԩW�� �����f���,]c�o�>%��<
�]{vQ��d�:��}�<�E%�;��nn�D��9���f|�c�`��ct'�7�"y7�����W���?q��m��� ]��� ?����>�G�_��y��N ��	�\�)(ZYZr��3c��>
�O����^qX�$����w9���։�<����N�Exg�(2GX2$S$v9A��EHe���&%!�Ϝ� ��d a�zpr�����U�kS��F�y�@�R��<�=,���+lɝ&��A%ew�p��h�S�u�su���1�rl~ɲ���~��U�! ��2�T��Q�����oP���k�A��"�|���`̡���{D&H
�㇃`[���)��AL�*]-�.[W����D�]- �F9��M�����Y�	xe�\�^�ê�o,��\Uy41������Zz����������Y���s<z�3S�Q�	Vbq��	HE�N4|U��ļ+L��>�'��`9N. �l��y�r���'�W�Ҳ����SFR�<���&�%X�O���2�;2�Ǜ[�~v��	����(��|ݸ7��{z�� LH0��U~{���Y��/�5$-�F��;E�Q��@���*�;���c�' 1F�l|\^��"�G-+Sea���t�<�I���,��&y�N��٣��r�2CGvz��]���q����i��(v"g<ǹ:������>��*����h,�Z�iy����fm��sߓ�kU�^~/�.�Y����%i�z�D�T�%kW?p�_��!_!w"h����5/w[Go���
_��W�H}!�I���K���Н� �p��IJ�_{v�m�M��5��%@zV^���mO�����]ӌDU`xkpS�]�0�^�4&�{�pF[;��g�&�"��1���Xf dQyP��}p�Yh;���	Q�]�m��V�����	b4n��0x~q�O���jA���EЮP���y^�N؊��*3�h�1�ж��*0�Ae~��Ic�2�8��RYuw�˜]���-	�^h�X�Ɉ��72��Jf\QGޙ��4��SB�Xg�^R  ����Z�z����.�e��E���p@I�P�G΍��x>�=�|oQ6�R�g�X�zxO�hSJ����ӿ޾�V;,g��{nI���kn��.��Y��	�X܄���n�G�؜��Lz�M�̝ �����j���8�<Y)͕h�I��Z��K�d��K�I����LԠ�y�������i��$���b&_%"�t)�V�q�Z8�be8nҸ;.m]�c����*l���X�rqo�l��ӐQ�V��SK,Kd]��IVd�����x�6��Um}��M>�;�t��Г���dNĬ�������[-�^ĸ��-�pG,�Dǝu�oW�!��B��D��I�S�@�-�E;�ee����6C�r`�ʏ��N$6Fmh�;�	�J�k=�=Ϋ/���"B�[.D���L�A����;JVE���e�\/�ǘ�VN=�v�8D�1��d���;*�7��No�+4r���l�}ho�{�4c�c�Uzٖ�A�X�b�������Y��FM��EFt�����2�I��T�����i{Jl$�Ӻ��Ohmf����G�L���$���i47�1�����7x��>��ȃt�|L� ұF+��6Lv,d�
{S�nB6q�k��@�k�F�w'���~��=�L7��C:�9�зW�,XW�m0\���D�����~]@x�Z�ȯ%��L�Bh�$���%#��S�-�	ɏ��>����K��Ƿh�D���?�S��<x��b��#���@|�ΟxX�ŵ��a��y���˦���uH��2�T��K����a���)*S~r	ů0-��e�#���>���d�x�%�L3g��Q]�db���*cdP��G>�U����Q~���E��d�ٝE,4p7�
Q#�ظ�z�y�>�8bS�ȉ	�iJ{���nf��#~(;eۺ����X:���)�ya�����@�b����4��,�߽���'d��E���Jٴ^�����Ӧ�d.P�y��H�Rw�Nn��7R���2P mD��B�4T4�,^��0#�R�����H�&������!�&��;�؂f��A��tR�:&@�������Z���|��N��j5��:���tr�氀#-��l��j�ɳ��P��F�_	�09�Z�5��G�,�o]٦D%�)u���p��`+���i]��g�ZQm�X��� #\򮈧QoEט�8�:ŅD���ru=��Q6?���k�.���F*,����/��c��ڬK�� L�P�W���8�ࠄ�U����r
�np�Ϣ�z��%�ذ(��|E&+�фK/�V�����?'T�(���1>�KjV�;��vQ�sVڵ�.�@���$����F�����|Һ��L���5I /�o���z�~�q-�e���H���a�����%!�Y���V�0Lbx���W$��o��l+�z�ѵ��K\Y)!&�!P�1[uU@ͨ��t��qq��T�1z�����GoY{��'�֙�h��*ѐ=�}K����RܦJÑ����׷��6a|�E�"�y'7�f��xI][98Q���8�nAL��A��XX�=��ׄN"�'���2H�tS���=lq��D�7�/�] �� �I���pQ# l鲽��@t�H"F��Sg�iPиI�B�h��&�#��C�ج����t���@&�Ӥ�}��?s��24*qͳL����4�`.�o�r���,'��/�ӡ�֤����DM#��Ax�"ȱ�V�H���&"N~KN�\61��tC4���V��65��9}&trk9��f��t1B����v�&���X��:g��E��k)�V���U�6����fF��g]���\i�D�{[�}��سM��_�2�_�G��Y���JN����_|Z�$ vh�+ی��x��|J �Uw���] �{��C� F�Sw�V�ө�4�o�(�=��d���8��������bi�G�.�ߙϾz��]����/@u+6,x���JW�s\�j��6���c�޹څ���8\D;���>6�aj:��4b�����R�Sa�p��"�p(������u�e�7���~�K�q:
���'�A�Fo1�_[|tt�<\,�}Q��7'�d��ElH)M87���QFE	�)tbP?aj�F��戨�6%����w�i�a⊷��(%�Mӎ�L�Yݕ�>h�{�c�����e�������4,�������)���=����+ޕ����!s��}~R�ќ��L_4*�E�Q��^:�l�������9່�Z֒���vV(�VE���%�9�r�K���rA�. ���t��^�['8K]S]��s��9�y��j��h#�L�7�?4|o!.��9Q�zvL#���SM�[}y���3��������2|]�;����TЯ�m�W����r�H�Mj�p�:ϻ��qX1�w����O���r�9�+i�2vt	�n�JTV��i�ƌ{��>��ۋ=:��n,�]��vZ�4.,3�]�����`��ds{F�V2\��S7��9�ގhAL�U��p�3JrZ�xm�52��{�?�㝇�&yB>WZ��3Y�e�@��V&6�G�s�o�v�0� �_���rT��|F���z�x�@8m).�Cے���J8�c�����rV��C^��AAliՑ��I�����@���u��f��b��=�hWCy/p&~�����А'����Ajre�&Cr�8����J'�$��ĚG:�QT���x
�O!�\�T/^T�n��t���L�ۍ�`x�[�*�*�C��w|�k�7楶i�����[#��cr��r��zg�j���>�v_ټ�~�(���FS)'	��n��LѿB�x܅Dj+�@eش��#K�#���`j��1 %~1�M�H��Јe�=�,����'@�r��<u�ڇX��ծ�3�瑴n��1p��XA� ccX//���`�o���̖Ō���jl����T�q����=V�м� �A�"4�#������Y2۹�Ne��4�W}jD*She1p���zSz��
���o��?_]g��BkՊ=�n�7�|[�d�W���@��:_5�;?袍:��Gs��R�|�8�ұ�SS�-�'3����#&`X��c�}_���Y����1���1��>Q�ֳʾo�O��rh��N@x�v��X��1��E�5�I<R6�R(��v�v�~5�t�g�� #)h'��[D��L#�QW�8���'�6��-�P�����'?�J��^4*����ke�d��GPI�)ةr`= (-8�z��o�F�n�����Y|����Yg�yqa�=�F�x��eh�;��T;�8���H�6�}'���?t�/���掤�o`w�2��ol���z�5��d�p����ď�]T9�3G�r��&n$5�8R]f�v�v�̥{�%G��\�	�j���jD��WV Y� PG�u�_���`$�����e!y�7d."&Zʇ��Ҵ�����a�=�\�3yݫ��O�~	����� T�X`!u�HC�Q�G?*����b���z���VA��x+U���{����0d��-�t�����\�|��x�@�cB'٩�A�nao1(@_6&mp%s��]:�&���M�w�B�O7�����5��]h�B4k��E7d�� t���2���od�s�Y�'���#�	��$ʮ@���L ���g���8����� 6�'c�e�����TO
�.|�JGr-�x��nriM�����p0�d�D&���/�b���q9eG��k�J��	�y����m������kʼ�c�I�1T���A����3��2�y�*w��d�F�e'p�o��c��7 �:���R�%@�|���K��F���!Q�ޥ~5p탯���O��=ɴ��=��U�]v$���7	P��Jk�L}�c��U�>�/_�y� �%Pu��}�=�\%T�96B�5o��������S�nJ�;��P�L�,ɩ����`�j��Ӡ�]:�EhPR0܀�TOG?K��1ց�6�(E?��c����X~9P��`ͨ��Kq$���)���U+idA����̄�Nz4f��>V��r���a?�L�s�S*��e�x��ŗ��lbV^gFIB2g��fۧp���Ym�ů�Eȯ���2��+\��h��VF"B�S@�ӣF�>'IɵHG�G9�|�5��٤E&����_
+��mȰ����`$���'ueA��yBQL|�_b^�N[J��زi�dC"!��dcS�����BbZp#��r�ϫ#
�%�\�t	��pX�zH�!N<���6��t��j��2�r�� ��ܸ�9��,�KU�XwDS/��0A�_M�O@eo��C� ґ��!����*8,�q��%�&��;�^�ߕ>_Q �.#ᘳ�RGgP1� ���}�h�תc�3�e��7Z�
)�5��	����*��i-����
��D����i��� �p��~��9C�����d�g������zP��|���L�N쑓9���ڋH�c���ײ�$��D�h������L��)�3Ecq���(mO�}%���X�����(4��o����)w�%�����;Ɏ�ꐴ�{�=�$&���;"N����8oh���aq�����f����p���D`��m�ɳ��=�zǏ,�j�\�W��W^�g��9���͹�>�;ݽ��N!�(>��+��`_^o!/��'����E�%x�oNh��A2���{����-F�)�⌲�#��02�x\�I�	2�Rk}n��ى������Q�)n�[Ԕ��\�f��'�|�T�eMi���q�h�
v��f�Ahh���L	���G�s+-_��myV�$��E�:���g�@���������@aZ���������U���~ԝ8�;O0�*���4P�P�sd eZU��c��E	��Ì7CZ
�w���7֓ �33ȗ��6�,t��2��RF��1���8H�8���?��N���\]�e���ӷ-!H��e�8>�j(�#Md
7��DG�3?P�À�����R��GOjņ�.o�ѱpD�&0�KZ�@9�я�#;�}x]��jD��7��A��@��(�q� v�]G4R��e
���@.~��[�@�>O� �:�c]��ɸ����'�B;Sy�ѹ�&pG4����-[S�K�]�u��G
W������)	%�t�RnԇЏ��a�ooz�S�������w��nߩa|�n�X%�8�OS��������b��rW̋�D�*�7D���
�mb�����6���]�h��P(d���j.����e�;U~����(r3�O@��r8w�K�|#V8�ﰉis��tb�9eM��� I�U�J�v��C#k�i�z?*��ٹm�G�����i߯�)ļ�b��w�Uq��9��\�O �rp�T������@��>R�&����f�Cek$m: �}�*FV��R]H��&z@��֛��m�Q��J�4��P�n �%Y�f�:�������)�y�	 �kt���S�-YL�u�����WZ�M�2���u������"��i��n��BotҞ��zj�Ud�� D�䉸���9d2�\��hGG�� ���f�p���E��e4\\����C��R�1	#O#?;AԳ���kQ6@;4�Ġ�cQ��";���(��7'˷��R����������LYg�Guʵ��A�ǉ��&�6�{�m\ �ȭ�Gq���c��x0���t�Y-���ր֑E��Dd=a�#i7�D����@����9��N������?�S��jG͏�����T�����q���c݃�d�td=R�/)=��T�t��O,~�(Iq�k��� ���
�
�cz`Iyf ��ٛJl����HzP��O#.y�����ɨ�Ҽ!���Ä��r��^��uod"�䦱��7U@��:`)�����cB(E]�+u��_���7㎧�F���ߌ��c�7�W�}� B"V| �?��~�2Yj�|t#�Fl�*@��U5�<�9UZ =����Al�g��b-�I�D���I���g?s�?����yd�@�F�ikD'l(�ɇ^Xh8��la��H��B e;��o���I�3u��ٖ�B��vġ�A�4���$Z�PL�~�,�o��W�C;ᨤ��q�N��'�X#��R�BWM�KYMNtą@�X Z�&�7i�jzi�/<��h�9W-(�B��wl;?9��[~p�Z��.�6@���Vj����t`p��ƃڛ_o��s�.�Pع϶�A��/��4"k0����Dq䪮���h�9c�ǜ�"��?�<ׅ�Z'��fC]�c>C_#4�i�`P,`��I�Ǔ��4X���q�)���e3��̺�b�Dn�3��-o��K�oY�b�tB�NC�q�+����2^��:Xb���oBj1x���C�F��Si�)��������q�����O��^�]a�z*�;��@��/ݵ^�����¿-/f�6��P"ϡ�3|�C��K��8��:�����i㌅r�uE�׈;ab&��\�^�NBtqi�sO�=ϥ��h�ϫO3|����4e�w��s}�UZ�O�Zv�� ������F���ڐ�fd*�)-�Y9a�r ���ķgX���5e�Qj�u�lص�:�[��*-T��,� \��؊)D�S�S)�{����V���c�/�
nz����
8K ������r��A�.�Ġ�M��F}h�$q@y��G�h��f������h�ה$Y��:/����H×�eB�9}�X@lV.x�DVZ�i�h���FN���E��6/"���,l��6`�^�?5þ���d?D3�E���ݫ�H��7$��#]�� �r��+%�S/��	a��|�yؿu�1��P�����s�q�mK
]w	&H�´g47�,�#��~_������\<g,n���V�Q\����
���w)
�"�c�;��ʌ��B�]y6%"���J���ɰعo ���1�6�v��z���f�9됡�׳c����i8�
I�E^�h��,[p��>���ܤ��j�I��m�}��!�ά�%��xS�CD4�bK܌(x]������D3���52S���p�A�P�e��>t�}��J݄W���Yv��8�I�7�%��2��O�BI[�7Y]+eQ�9�W�V�yG��떾�2D 'F��h뚜O�������S�u�Z�&�>f�.��$�֩.��Qf�.��9'�4WO׭/}$;�f��*x[�ڀ�9��:�3��O����NIǡ�12� ZNvT	~�;�X�k����`�1�nĜۘh>��^��DR�jp<��{zh�7�4�(|;i��dd�6���t9����������nRVP�{^EwE8���Ȼ�׃�s�=�7L N����n`!������;庌#Xn�������� �=Q��S�����yc"+|8�ņ�W�t[ɹD���?N�
@Њ�ǟ�`�9H��FK�$$V�I�����`�Q��0� .Xq[B�I�}�����F���':����r���.��&�C�T�4���y:(l<CӜB���x�<���ǳR����y �%�Y���-��y��R�؞�fȹqWۿ�Q�;蘂1ZY!$9��T鋷m4\�q?����vE�B��w�����zߨ�"'#�N)n�l�x���=F��R%*�A�jJP�y��}��\:ĩ9?.��ć*�Z>��^�I�/j�d)f߃�7�ȭ�j�!�� ����U���E1��,/m>C�ha*B�wTM�ڃ?�0�'$k�\v�M�χl���ˑ��o��@�KB:x���M2��o�Ob����I��A���__z�)tL>'��G�W�"wc�V�N�T:���`h��?�չɆ3���Th.���u�ʵ��o����z�ԎQ*���ذ�Y��Z����cŜ4�����eFBv����:��ɏ(�h1���99�H������3�}Z�G�eő/%��gCĽ� ��1��s�T�]�'�!8l�D��m���R~h=�w8_,�o<�7����~���mk&@�|I:H�;����mG�ئz4��	���́~V�C��,�k�x����h�"� X�o�X���k�\X$ey�$T�.[�d�"��苬"������L��E��T���b	̳��>&�^ɓ��ǜ�P�fBA/��[U��jb�UU����Q�SN0��o�R���jsx(��V�,��ܗ���h�u��6
�?D��/.�^u�oK���� i�'�k��qx����N�h���x��K��* �g=|~�ߴ�O�W�`7�7npP=:nvd�&/j��)�o�����o�X����獬���2�ϰ ���IPg0E�Ǣ�jb��F�����d��^X� ��s���
�|�� �.,Rzi����:-[�����G;hM4�0�vnF�ږ��������d�`/��XO���q;�|)��ףIE������;�m�E�+�	0�7歺C$����-��(g�kypvS���kԑ�A�0׈X�Zf�D�aw|.����N��T-U��t���OM����2�RKo��}K���Z��@K�%���D3E��A#2\?�.݇3��'�ì��fA�+t�4��΃�a�Bx�܊����f�U�~��M��X��P�py�]I�Z��Z�
6�5��i�
 ��X��;����������>�C�^�����܋�BHw͓�k�W��xA'�*�AD����J�hVP-��s��=�6=-�Q/�F��Īȕ%�k���V��b��;��Y�r��|��^~��0�sM��A#Ug<L�٪w�oJ5��c�~�&}���)��`�S��q��&<x��g��>~���t6ڮv1����_�[hFע��tpK���O<ψ���9���Oh��@��֣ڂv���`~����t�@GK��$ �	��G0r���bա�L���~@4DT��y�]D��n�c�OV��@����\�q5l9{}
,z)��,�	��6o���;I�T\nѷ�c�jԣ@W�[0��<V,�W���jlo���*Ү���8)m�8S� Pv�+���9A! �b��1A1&ӉI����S��pq8Z97�<�w�G�B��.�� 8�/��^§W��6&��ٚXliV}��v�'�i��z�4��Sz�\r��>k3��d��zeG�z�mCJ�{u�m4U{�������䇾W�������#�|�hIjW+��8����E�e����H�MSݒ�+�O&����p�����xd�4k�};�w0�f������
�4־E�� LO�l���t
�q��*��2������\�6�f��j�8���?��Ë#xH��EݱUܞ���8�7��R�����@6x[@j�+���� ��X�*L�7����E�����n��4�옌�m�����}Q*@�	t��qYS�9Q�8�v�A��d�A����7�u��3��\P����0g�=�gh �A�� q��u_0xw\*�����P�̿K4�n��>���i�s>'��p��� �����W�s��d���T���F��S�'�3r�#U�/�Hb���cG&�B$���潳/�bG=����I�u�iN��#�cL��D�t˰���?䍤��ې1ok��<
&a~P����/C��y2έS�]��-����U�������n����R�<�:�������&��t�����
v��א�e�5����&�"�KE�����Zz�&���sT�6���S���F#ǌ��9_�9�[�кlݰ��"C6ih���)�U��NrT�P�R�ζ���:��SAe o�]���V[�en��cSiN�,�͞7�֯���9Ɓ�N0�;\�!���.��7mx	j�)7ҭ��%� �	�l�i�v3(ls}g/�6w���).˼�kF���>@���cb�n�J3u�]Y7C�N%���׽��2�����0�|�1��c����+��W9����1�qh��XyH%u�ғ�^���HM7�l9hwk���K�i�)~(mb�w�dG��9��z���r��?c&t<J[�8�R�>6z��/�Zl1_���("����;>u4K��Jd&������Q�x�{U@�q���>�jǣT�jXq�MpbM�94�'H�m3�=]�~�Ź�X��m#\r�X�~�'3��QL�����!<;Ϻ�)������H5��0/���A����&b�@����Vmv���޼]k�#Bfd>�'��C���D��;]��gX?��v-�9W}�"�ih=������÷������@s���{��-ώ�v���ѽƟX�]��0>>��K�,�^q��@4�a]_<í�"�4{�8@�(��x��j�3�-���{P:��gv�������ZSs��[SӖR�V��.��ѱs��Ja�wz�I�3'���]�7�6FU��eVyҠ��Y��'�zֆ_`���N���A��v߉Uu��g���.�3�~���c����{��j����^��S��:�P������I $WI=�߄'��L!O�q����.)"a��0R�gd�?�w�\w`<O��oSIqK�w�v0E�ъ��#^m6�h-D`��%�|/������Nq�G���^9�<{l�ۑo�
��;E�r 4��o�'܄�w'�xs�47k��y�->�򪴵�:���v�ϡ�w�G?�Fq�5������ݼ�E�1�4�}��o\���w�V�ѐ��9�m�,�Ě�O�߀�{0A晖��_5�T��������f� �)��~��Qt�o�3�|����0���n��[aԆ#T��u%͸�Xn��4�Ç��mL��UM�o�aR�U��D8���=�	\���3�7��NlI���/g����n�:��Ѫf�kF!.�"R��!�[\��fW������H�Ѥx&�IZh�|������ڡ/�[�WQ��w����p�mW�]E��AًR���:u�7��jG�ns�sy��@���ύP�P�;���v�bғ��[C)��_ ?0=���)v��I��UK{���7�(Nـ�~��|@�51T��Y
<����Rͮ�с4�%Y*t �j<�q�"����v6���k�`�$��O�[�D[j�W�v;��ߺ$���{|�+y2��.�[4D����	R�l���"��R�$�+B���<�> �oL���F��-�(��)ПMjn�i�Z�(q;��.g�j��\�x=[��z�28��f���8�@�@z��&��~y�h�F	ⷸ�+EW{^bX������we���}�E+���]��j��k��'@���^f�~ ��f���nݶ�J<�+�+���6$�h��{��AV �q����^��r�ZH�_%��y����E��HOv'�� ��x�y���,�=$�5�mj*A�J8�5A�K�*�����ݖO�	":���Z6V����9|�E�f�u
��# ��&��'��T&�IQ�"\Q�ӹ��(!"J����l�DQ���#��(�?t��@�#�WÖe���&	Xjd���z�t��i8�}��E6:�k ���ks�����%A6������QXE;<��6��ovU;Y���5����� r����1�'|�7(����Pn�x��6+'�&���]��-~b߂�E�I��Ŭ��{����i���-���������Ʊ��4���c=�a,�����~��G�o�F�A�S��3����FF��ӌ�n!���1�TX�kOF.K)�� ���\��ڋR^�Zh�x�3k �q��;�����1WΛw ��QVq�O�\��Q}�':qǻx9�E�=�^��u�.O����(ɳ�F���h�,&胜"� �4�t
�tB���2��}�J&�owR`�F
����F*��̗���L�V`����kyJ83��KV�V��阇��/�v�F*Ӫ#d|ř[�\�%�;�j�<�l�,B�������.]2��0H{���jt���6g�}]|t+#Lt�v�N@��W�me���BͿ�a�/.g��g�/�<�;�#��w�3��K\{�v
x�	A�� w����~q�s�S\a����������_CG��&9\�H%���ls���RUBq2�$4��~&�Sz��F�$�1��|�Y%�ihU?�c��	t��@zy�n��T��~�5��~P�>�Ď�}�[����0v9�H�eŢ�
�<K�g�`I��rFk�᫞_��LU��+Ŀ �[��̸�����L� �Q�!S\�iPvb�X+��:G��p̛*�3��r�:��� M�ۖ��4x�	�E�[��0�
��|�fL�w!�#���S��[��"[�i9�)���ff@`*��kĆ�@t�"_��3�(rr�Q�(���oǓ�V����T�(�'�.u�������U[�r�b��>��@߰�Z���+��G�6Q qUA_�ĳ	�ߚ3J���8ŧ�;"?����]�^�!d�+�D�h��ؠ�bz8��%Ze�Ɓ��i�!�����z�'�Y�*�8�.���W)3�}��̘����lT�(�<�?����#��8x�C.Ls�/s�����
�3M@ɝ؇��m1t?2�[�
r]�a&W�cu�T��=����J�v����7�+�^ʒ4��dt�8k�U�:X���}%�����D�3�&�#��ʖ�`ϙ�R!�3�|���!�8\��D�ƨeh����v��|�F�����r��7��D���X�kPK�Hy�� bd.XSPҼK�#@�|�Q�a���˄���A}�I���������Y�_�Ģ���m�=(.Gv�5Y�8��ڨ��0pD���
I_�o^׊�� �%��Ue�Qo��Ƈ�pO9k��o%��b�#�� Ŧa/�����\M�%wnbO����s���(�]cPG%�v�w�@c~f��M�>#��b-�-�Z��ZfN �pF��j��ɖ����o��ۊ��2��6��V�w�W��v�� �zX�����h���#�miR��:�sͼ�z��� ����DO�x����.7�/+�x[h�E���$:4k�9�+p&�XAax<R�+Y�i'����i;��w� �-R`�3�� %ʨ'2C���� ���Z�@���؎�=A�+��l|��r�=Q�?�D%��#ܮ�]��1���<�'��8�=Gc���f`#�!496�\_�t춽u��Pۮ�I}A�\|���� ��_D�Ski����P.�!WJ����*r����F�&���_��Q4κ�Y��|άW�ԝ�ǵj��g]��%D������]�x�R׃a1N������"��U6�6ᒘ��0K�����^�XA�>]��p551�
��K�V����H��˚;=d:���˶��7#��":�|�Ou c[��w���|s�h�{�4��Ʈ�r��0U>G�;�F��cE:�����T�� u'�L�@��7�<�ur ��m��V۷��K��g�&�7�2p]Q�خ�~�t�O,��l�t�E2��t8�^����	 ��K��P,f�bh��QVA�_(B����yX.q/(_�z��DeEY�>��S�!-�,���pG[���O}O{Yj�#�T�u�V/����_bx&��� CQk̸��\؋�c��V�b��YRy�&}��8 ��H�;}a[���j�]d�>�/L1ǌ�VR�qɃ�(O���'w�&�\�f� 3��J-N���\�:`F��_#���
�,�	2LgN�9f��H�(ͦ����� �X\�d-t|�t�8ѱ��$R��iGVm��;|��i,����@�uk�a[�I�d ���\O䴳��X:���f�B�4@�����z�R@�r�/�3̷[�|����T;Wv[-o O�3�@�&�?��D!Y��
y�@�T�r��A���W'.�
c Bơ����<Nc�HD�3�uaTD6�vh�KW��ť) ��W����N���ԱV6b��j)����H	2}�Ð����e�7  �}8�b ڥG=�X���/0V�pYv���L%��lvN�L��P��MG�� %����u4x>l�;���8;Tp�8�WE�a�^�;��R����
�wL	��`�"2:��ڔ7�P~� �����7*5?\p&�1�����)ޖ�K�)�
��^
ro��C������նյ�ㄤ0<�<��Q���"�*[�?��o��4�w��՜#e�_�jz�� !(�����w��}1��ō�9v�^rڨW�|G�VF\�;r1�/��n��U����Ի���70֣��k��I�r~c�9:�V*O��`��O�����+�R����Ȳ���y%"���Cr1d&�ۑ��ٮh6�F�73r�I\#�_�vw%f��j�:oYڗ-�g'�����`��С���?�^�QC��{���8q���+���
��hF+8828�����Ϧȯӝ���u�u��|�w4n ��M*e�؀@|�Ǥ�g�`�<`آd��'7�L��y]?L��r�4�$��ˊ�6X���0��
c*��� �S��ر`�d��fz�?�i��a���S�$��Iݛ��E $����ύ�!�z����p�"�*�9	����E��� ��r���p{̕I�e�ʭ����V�˸5�t�q�����e1�C�d��>+Ǝ��0�O�ƾ��C��3�g@w�:BP�d#$d,*%���/�FzB���J
���h���,lscY�5H����� y�'A�\���hc��eC:B���r�9�Ɔu;��+rx��b�%ǒ0.�Ύ��:@,�*�q��0z��7��Ӑ�Y� ��Uj(C�&E7h4���d=��wLG����P8��49_�ȄN-��;
�u�0�Z����-)B)[�`տbl'fM��ey��%x|���j^ \n��x�\�9����rp�3�6�9 �O����á���^M�m��J�(X��kպ(��x����bh� Û��B^욍 ���h��1�)�#��i�#	��&h�[w��⻐� 9�;uI�n�5%.Ah��PY���^`�F�OiQ�jB����H��2�[� WL�|�L�_��xſ�F�z1HP�Z�TP!���Fl������_�k��j19g�sm��zU���I�nmԟ��KR�[�(ݩW7BNwҳ��yk����s�x�V��@���d/�T�Faa:%$�v�.�2���:-�Y�^n'z�0��d�|n��T���s�8�#��rx��[K��-t_�wr��i�GT���8	�#&s2#�6ʦ���e��bI����D��G����B����"�QȆɾB�[q��)�Ic�i��w�L�gTLz��em��X�&�?�N���S�׾�H��Y{6�2�g��[�L�.N[��Y�z$`>�����ؕ��U{�
���ϖ�s;�����5�Ƶ|�k��4W���s`-_���e�|q�]�<�{t���^���[�e��K�ؽ���A��r�r^��kp�7͙�`�E)��+d�/,��0j�@���=�$�`�-��q�����g��~�S�.�g��ɮ���6��"huc΀J�׍�_�^5S�q�;����e}��u�qa�`�9��G�T����_�wV�:�OrO�_ـ�?�{��������S��M0#J�d4��%̔̀8��{P=�H��h�(�$s�Nɕ�Q$�)��p������#�И
�,�_t��M���ῤ"zPk'S��L3$>ht��y��9I���j,��,��^�&#�~c�W�B�Q�?��
��忻�E�l�T�>�~�O�ǥ��V=n�o�iЎ����A����wI��o�@K�uz�)���麦VuD�	˜�9���қY��������A�K�x	�OB�/��{*ԕC�L2�t}�?�
ΒN�­	��i���9�y($'���,�~�J�n�������xy��8�|A���a�@9�O����yE�T/�a���� ��o�I��N�vR:�c5QnTtx��j���ʖL�*_q�wh�q�y��1�N2�!E٥_�� s��T^9c�%�.(ؿA�:��c�g^�=ez�7�H��B{b	8
�QQB�649�@j)	ש��l����NQy�Sl\[z����1"۲�f[��k�N<�e�TIآ��\��v%��*�\�aY�����߱��7!b0ӌe�[�uyL�Z���n3�^*��?�냭̗�Hn|Q��$��J�����^� ݢ�mڟ�,щ�S0��ZFT@)����%��t'�=���,���K>^TMl�f�B�&;~�!�� y�9@츺��F��䨽C���t��y�L6M;+T�}�\�Q�-�ORKm�ϰh���"J�H�X��?Yg��B8��XfAT ��(���VFjn���&�X&@F�Ҁ�V�G��
�y�ۃV�$���㳩AY\�Q4S�Vuzg�ַp�%8�`��H���L����k(�'�Ɯ���>gSf��&���
�W�[�ʷm1��#֏ʧ��@-�v�>��Yɟ)�,`��<��S;��"��]I��=r�nq��u뷬�/�w�Y��6���=��T�O���������i�ɾ*k����St�Sz��w�B�NB;��p9�C��������Z4��q�����6�~�tZڶ��!�萚�!Y��q��x�>�]#^�-��GA��|��U��q�ʙ�JfE~�����	�;px�mq��^�ߝ
���kp�_�o�d��"@�J�KB!g����iZq���m��PԺc]A�Y��R6W?���������;�q)�*.)޿D�Ӣ	�H����ؿ��XSRs�1��D2,�D�jҋV�E3�~3�i�6��{�;�c<qߕ��U��#"8�6o���XiƏ]��B��҂h@#����E�~�#r��� 2HڿfJ��z[g9�E��m1ˣ��R�~�a,�Ӡ�z���U8E�{�'�Ĥn�&$���ޢ'���J�~�?q�Q���<ag�
����R���kذ���i�� �Y�b`u}�g��X-����k��k�gaX&BQ,��;W���h��拐9���M-v�J��1�Ԫ�2�:4�qn���G��W{hf	o�f&��X�:lB|[;A��-��ݜ�Ӽ�Ԍ��$�IN[%Y�aG肬<��l��B��Q;���l��ɢN�ko��N��HbhX?2M^�ME,�C%��g?!rH��O��w�J�<���e���v���$��No교������1���'�r �!�J�f�G��Q(D�n���C�����N x�[��q	S�)�uRc~S�%�ˀ'��%P,��Y��
�e��\Fu�+�"��pP�k?.b+Q��N8��5=`�๐���A�x�<|j4��feGA�!�T��3�=Y5�]c��b�[~�|��;�Q'�
6&�T��c�0�D�*�`a?�<�Ν�`+�1�,��։�u��!+(�x��@��q�*��Z�h��^Qv�l���5JX��������(-����Hܖo�陼O���p��O����'��\�jf5M<��y:\�X���HiįC,k+�1 ݺsv�x��Ǟ�y
#2=t}
o�D�`ɒw#ڼ����	����k>C�E�N�d�U+<G�߯f��.��/~`��7��a[1Z��b�)�lS�刄�5�Kǒ�
��Y�u%�x~�ZAv1�Ȋ6kܾ��!��'����$���t>8&U
 �Ф�
P�/�XP��1��Q�h�կ-�ר��
*�����	r��4|T�.�Lu��cfd3��7�#�b�-�ta��$��A����C�`�H���^sf�O�*:���6L���b%����{�9,T����4�>gQx��aW�ǘ9����q��yOo�t��P7"	4��y��p���$8�v�*lɾu��w�}	��0�EN-�|�R��6�"$�pKw��-6}/�O�B�R�+_(p7�8&�%f3�[�Y�|U�4Q�*,�a���6�����ԡeU���X����8VY?�<��u
k?�p�Z��o���l��'S�⛐��]�iN(�8�mr�2A��@�{BO�*_���
�=�����X@,�0�'W��bJ_����	�N�����]�|���AUp]v`F�DW��-�z&8�N�(�y'�p�ԓ�v�r������[�N���~iM���H�'̵�b� n��'1�4�;0T�gy_���we�
�:��-�Yu�8��Ҩ�X@\ވ�d��e#��<���k�~�6�^G��/X���JLDc��w��I���ɀS�1e���҂Y��Gdd��N�;�EL�G񋭹XA��ID��~��ʣ�]qJ)~����!b��G�M�-����6���Ă�Ce=�P
��O,�#�p4�F��<#˕��qF�K�7�����'��4��=�#�Y�30l����4��x�::�	��s�j}p�ٖ`����t�x+5�fk+
�!��/�7�4vi�.�<�5���D01zБ�V� �k�4���6I|��l8�Zv����j^��uk��S4R�X 	�(�2ԝI���Ȭ��H�L�E��a�H�!Q�����qT�PO!| i�5#�^�Q���6�bG(�趔�;���I9��H�1�Q�ڤkQ��9N�NM��ڤھֲ������*rA�r%�*�c��T�4�t�IwJ��aB���5��$Yǡvc��k��m���|�T[.a~���S�<Uo����U������U�v���%��tSh��3�ȮmKS�ѫ!��7�y��[�j����.T�/Bi�dF���l0lG�7܏��^SD�Psu�i��%�&�Aғ{�?��=�O���X�ӈ�+y����NKeBr!�^ñ�xs��:t|���a͒��;22;�%�.��6F&$����� d%��ϸ���������|�;.�`� ��0?X &��0�6�x����A� �,�.�8��q�[P����y���rÌ9���g�C�	C��B��#W�V���F=�u4����E�D��9j�9{Ȥ���8���2�)ŎVFAњ���]�#�٫�7#�'�\���ӈ
D�Z[�:���T`z�7�z�NMq�r��+9�,@�d��g��+D?1��2QJ�fݨd�48�$db�ؚ3�{!���h`�	,�ϕ�pϘV�"��m ���<��	vw�ݘzG�	����6��I;>�pe�I�>��C_,P7h����g�6�]��b�K�4@V��KKjU��q�T��WV�Kf霠�𘮦�Y�%�X\6�Q�DT�� ׳���t��Y_��/1���.2�q
�9���>�}ĦX!U�N̆/�ʇ�PUo�ݚ�-i8��jY�v]Q��L��?���M���rĭU��⚦�Bx�� )h���偐�KGt���P���x��}>�v���d~�5S�ݖ�2� h�ye/�
�5nVw��GCtW*�3f��?B��s�����B��@d�R����,KC�Rf�t��͍�f���N�_��#��@
��zïs�D��U�[��I������d&%�_!A�Zm�	��=��䉎J����As�]Na1S����!�%Ӡ�	G,��}o�7h]=�H�m�촄-��H���9�<�Am҃���[ ������VD2�$Jߦ���X��J�`߸e6m<~
�����t���IIT��V���>���
}�2#��Gf������J<3/����hDS�Xf,�n|
!f�t��֖��h!^����'�E癈�׫ x���*�5�G ��*�#���S��y K��&D7ǴZ�Y�v̪m�B�
"�u�u\H�t���$d�1Ba����6	��@BVn��][��R�AeA>t�p?�|l�Ν��bMÄ"���@	���Pg(����Y~Q��p]Y{l32&N=
~8��x���VFH�-
��@U(�d*"�3V��ۑ��E�
��ǜu攜U"I�DӞ��6�z��<�K�O��S��uAB<�Xi�	!�m�:�h��޹)Om�=�m�ʼb�ٞC��4Mj�y�
�\ɚ������jkl�kg)����S���栂$��X(��[��~����P�>}]��]v8��mW�;�tw͡�w�4�����K��e;TiN'�D�#`<Z�Y��E�����օS����3�ml�5����\���oT��R�		��(��O��Sc�m���j��Sq�	��t8)�'A	����_��-I\�+�@N��M*/@H�����a���v����Vtt��������O��&U��"�\��}�f����9%�Q�4���$v̻Sa$��/�BvVG<� �+o~5�>����&ʟ�iE������0oOā��<2�i�=[ۢ(�F���>�ނ�Fy׹2�)�;7�(�-�6+�nF�w;���#Ƣ���$�Wv)����<ؾ���׾-�Qt�7�Ę|�0��Wx�I}�鲱�-���m�c�F긂���x�j��x���Pm l��=T:�Hv����0���ڽ�f+&�Q,R
�o�Nm����$�g'z�a�t�z܊ J��I�
/��X�?M�RO��oϪ�	��cM9������'�F���.3��f������!�V� C_	�����}������ީ�H^O�!)�h��+>h�Y��;��ھep�b區�g�ފ��.���S� ǫ]�F<aȤ��;�;$�Q��J�>��v�z!Z����nP0����d�!�*�Ij�/�b��#X��M�0�4�H���6f6۠���390'�ul���xb�S�7;Y�dvB�l��E�����I~����\���u;�_N�m�M�t���alN�t�8�N���kKj싚%�k�",�U���r���ǧC�\Kޥ>�6������.0�oc�Ϲ�~!!8ͪ���RTPr���%�'�(̩K!T��w����-��!�f����D�BO�q�㜫�/Y��^��;�{(�-�en�zQ�)q��Pfhuv �vQ7*bA<t!#�Ԉ"��2	���p��t��N��Jf|o�Q����Bn�����19�#R�72���Je����� r��X᳸9�ot#�ڐ�I���d�XG	7�8��訟� �t�:ۊRI���Ff��v���!�����L���T�yA��#���p��Y���
"LU���R/�)z�7�.�2W����o6�2�<e��9㽠�]09b�~��mZ�W�]	Zk�]����'�z�?�Q�.*�;z���cx��y��[�Zy[�\�����%������D���w������퍨�P�R���|��e�`�x���[����m���O|pr�.��J6v�����ۨ���]TFQ��_w�h�VG��ډΐ�*�q���؃�q&v�\j���*J����2j�ڢ��/҉��r9oA��H����s��O�)����r���E�xx/ϕ]z��Sc��,��W��{�=5zDk��:�&�d�ȱp�B~;S�/��5`�~8:Y"o|w�J:�p��i�\����0�Z$�`y��ef����� �]��8�r��J�cV��%���Z���q�7�*s��b+�-�0�N�s�v}��$�q�br�D(�HI�~O��8.���J�̀C��v�g�o�x2�ka�I��7��bqbx�B9����a���5U�0�U�d���;�STA�l��"�q R)T�L٨s�#	7����hj�^�-��B�J}q�
��e���.��E�F��q;l�)5���И�}M-��]s���K�����@���ߛ�Hժ��`������Z��1rLE`X�����HG�������d�R��V����8ҧ�PA�&����Z@�̵ⅴ����c��"�a����`03翐}~��w�g����s���-Օm�->_�LðO/^��(�n��6�l�vX/��N\�O�>�`$�r �m�\�c�]�䞚!�!�ŷ�_="�,+�^=R�ۭ�y;~�u�����kb��u��E�or890<T�=�3��;�/�H`?u9\�Gk�<%�,@�<|%s��[�u-��u����T%��4mY��Gq�\;_�K`I����0WT��A���������Z4���H�>��G�r�\��6[5=U֥�%ϼL�E	����]�	�
������!2��>/2*��B�泊��u"(�r��ps���DZ�4ϖ��4��i��6}��{��?�`b��5�b���.QE�v9t��Fi�ʶ�d8
��R�QFw�!П<������CK��tO��+�y�>�d�ZZ�������$�����;�ҵ��V�O���C�4�ưO"��]�Y���FV��!��f�,|���TH�)�к�M���ׯ�E�v�Ɩ����,Ȥ���Ǻ��d���%u�I�J��]��{�
�_��u��+nN�ɜz ̝_�!pxH�<>#�����N�e�Ԍ
{�ݷ=�-yY��h��r�{���$����YI}��V��@Ȍ԰�ܫ�p�Бr��+H<��.�FW�G�]+š�;[���}E+���O�m�2&6ȴkm�f=I"Ǒc���}>u,]q�ׅ����Vh������u4�I8���#��
����;�Xb4���O�I^E}	�r��2�������|/fy�l2���.�S�Q����{��van$A��`Q�H�mܑp��_5Gmu��.r��FGv	�+l���ċk�$�1���ă�_��'L���l��D�ѝ��e�I�oڼW�d�cd-�؇/�C��|���i�0���*�%L������z4lh����J���	>��\H�i4�(n���x�`2�W	0�Hu}y*G�90;՝��%dq�*6�༨�
0�t3�: D�s�o� 7q������u�zB���+���ͬ�y`��U��l�-������S�=p���$�d�r��D�B���)%
���#�X��cZ���G�9���8w����b���'_.��'7���q6Ga<�|�KϏ[��,`[�kȅ��}-�0s��Lf(��}�/��3�ϴ�Naͱ�Ր�gq���am��h{(���yO���	��e�?i��J]-7�@ӽR2�K�?����jn�:�֬����� H�<i	mb�C���sP<x1R?giOp=�p^X���C�O��a�?� Ӽ�Vj�`��T9�d\��C�~�P7�����B�V#�Κ���8RGs!��G���Ų�
��ʆ� �{���s>wx<�b�����������\Ɂ��r�,.�x�2E2�I<Ķ��	�g��?�V��>!̇_��J啬=� �B�4]%D��.5m�؉lM�d��ޛ��,�δs���1Ə��-4f���Rq5��8�Mc
�3v�ή�����$��Oz�hJݗ�t`g%�=	8�v|�zR&��:;�8&�:����G~�NèN��e��,)����o�
R�U������yU���#��$�]�q$�P1Ɋ:ߤū\�	
�\��)]�0�!O6R�.mE$��A�4`z�4�wke���_3.2Y�c���WMwzw��To"4��]���M��X��皅�������rL��?�2�s�zQC�r���S$^a�����N�7�5�cs4<4�@�%�k�C_s�-�cZ���s�R��e1��ˢ3?U�@]�R�_w�4E|]��vx��ux&TV�%�
�ٍF�,,����_o���A"�g_�_��n|�5��Ra�㭱�G̩���0��C`{���xA$�a�p)Ki=ʞ�Ga� �a�H����a�ӳ>Q��t9�x��e�p�Sx?��~4fzH)D���v����T%�����~3�V }�Y�5�����h��}�X�fJZ��2��#s��cwP�l�zӏ�`̒
c��6I(��K8%]`M�eW�z����V��P�GZ-E�W���h$y vT��C�*U��Z�c��	����܌�n�Y�9����Vj��Aߜ%G`��cM�5��psL,��>]�\��_��dt�m�r���kvMG�a@���:tG�cY���5�����n��b�p����ɯ�ĈV����N�*���E�v�3���C�ؙ�])9+K����o��?�ܦ1.R�����m��@�l�)�Τ5�>v�+�� �6�C3��,���g@ ��ߑ���p�S���ò��^�S*$���-��!N\r%0T;����F�뗤��P������֌V�i��NB��b�a�'�cw�ii���?r���QK,=��<��=�}����E732x��`�`��(�����~E��@��p���	qBE9z����U�@���E�6i-Lh�H��t�����QS|%��e���F`�"ju<�̕g�}���)*~5J��&�Y�?-�q��'��C��AW�u�L_H뗧���m�=$���p؝�GR��64(Rʾ,FW��a� y7���PGB�| ����t;�h_��JLU5�-ɰ��k�	��P%�p��+�/����BU5N��^p�Ej�M<g�rR;��=�T�	�NE�|`DH�<=��8}�VaA~�Y61�(�S�k�������siR�������*IL���䭳1�o

���3 �C�����(�O�
��_V߅rH��3e9BQSy�<!-*�����H��@LN;Y���*:r�6�ob}\l�A	'=�v����{���
���o�r��Z�'_�VJ��V��1������,!��
�o?�U�~������'��k��s2�VV�)����(�DvM����k}k��wg��<��W��"�M�v�e�AWY��a0z�3;)Hߩ��=x��8&)>�#��[�C�Ě����ne�B�*%��]p?z�H�A�����h
�L�<���0i���C�g
5��mf�YC��aT��mX(�¢��ޖ��1lx]H'+�u�!������g �G؃W�<�f�8�e�J�t��%��n�zJYr�~f�kpˑ&>9%7_���v]�r��f[7*N�=��[(���.&����`�-�H�'r�4��2Cf4E7�N��`��a��ǂ*���(��VjCF>��;�> *�)W<�X�J��T��u�V1L��t˪'i�/.�k����(�j��� ��b�'F�.`B��h�UN��9��|���tP��ܤz}0l6qz���1��y�:Q1�|�ay�y�d���FR�V��#�(u���g{�J�=T\B�rd9�,I��5�af&�Ϭ2��>#ݫt5/��ͨ�Y�����x�]�i5�Nd�r�5H�$&��i����p^��ЅH�P����ɚ��~���)�X���D�t���A���֕]�v�Ḽ�e��m��S��Qɹ�!�
��/�m�5eN��̖ș:m����#ՋWC|,m0��������0�z��P|�� >e���;�nƍ�c��\{�]�QDA��b������D�0N6������A�� N�Id�L�7(d�(�N?#N����?��^��>�����]�e�ջx����J�Y����cM��l&	���Y ��u0u��9�A�,����I�s�:��j����z:�S�� a��z�9x).g�e����y���iҼo#� ��n�����s`B�>�[�5�O�1�����C�7��}����r	t�]׸H������-��A|�tk~���I1Qğ�VR5q5�f��o4L���5A�*E���N�0��Ѥ��# �1�H1�Z�W�L`׆���Y�����+�}�����B3D۰^0෯fUM�QCꈟ��6� ���J��yx��L�m�l�rȿ=o�H�c�^m��ȋ�)�wТb���`�7W|B�?�y[,�<��,�m��̵X��<J��f���#��jx7�z �(D�L�L�>+��G�k��QWS�A��]�6^sG�S_m������,	"�a�)�TC��R�ucN��dĳu��Y�vЍ���(	��(��jg0���f�p@P^�}�^Av��ꌴ"]p5�#ϵ�D]/���hvb/s��z�a"�:g�5t��.����=�D]3��o�D��|��ڶ�N�S�ݭ�� űz'�H�Y ��,���gۻ���lQ9�-?�A� ��'�y�g���x�W	�ѻ_ɉ��i �	��/���8�Se鏧�bY�z�� �N>�1�N�^P�[���r���n1|XN��dH�|Gc�B����(�~�� ��ȯ�p���Xo��؈0�PK'j��b��J���*-����6���jܓTm�V$�`KR�X�4��b�3������0�_��9Lz��1n׍�#B=gYq7�zU<��8���9���|B���S��=�q8�����-�?è�p���C���0־��K仑�/'ۊ#��t����1}�<H�-�|X��]�|���+VRV<���
`Z6�Ls��3��H���IU]�V}D��cW����l*�?���xDf2��@~�ܐ��a?񚔙��K���G�QR��Z/^�5W�0��"m��}��M��m�`��M�؁�J~�Vmx�#��؜����@<A i���G;�U<�Oz�]q��������46���/eu��l����-������-�=��q0�L�u��}�$T�����]��d�,�>��}�k���*��?��àr�~0͛7��ķ`����ɂ��[�Y���>;���;�(�q�7M������/��٭W\|�\����ˮ�Z�K�W20D�7�p6��B�$S/ɯ5l�7L�k���3a)�2"G�y���
m���2����H������N	\�y�ъy�_,T63��k{��hM���>t`+���hD [��_2�J�)<���Ka�Q�ې|����u&�7�r����i�:?�o�!$�^B�z·-�m��zշ�-v�d��ŝSW_gGn�(-��B�Q���Wΰq	��~3�>>��F�T�����ߕ&��%�=IV�Ҍ�J��٠�_T+4	+��?�9�y�=�o�!@%e��;�j��N= 1�A8�u�>3�J�|�f�R���C���z�=���0aɚCo�m�z�t]�q����_�ӱ_���d
]�!�	-�Vԛ�����8鐺?�T��Q>�b#�Y�CA���sotl�z�U^ą�^̫�9e:�͒�h���i����(��� ����6}�_mW��c��*� ^V(r:tȁ)Ż(��BPKD2cN�F���x�q��m�|�|j��"����J2w�e��R���ī��*��]��Ը����!�(������X�۲dK8���V�� ��\j���{��O�O��ۧ>^�z�D��kL����n����RD�`ÚZ�&_�����X��ǖwT�0
7�%b������[�46g;_;N;������"L��jI�Ĳ�io'���p�"_�މ\(���{$0Bħ��KA����u�~M�3b13}��&$͈���$��6�� �\122>��s��2����i��#S@�PL�KN�i�UCZMgSѣ��I���$%��J1�����c�,�,��W��Aq;c`�_2d3�';��p2���:���_�{
������G�f��W���!Hԕ�� �R[L�`��I���z鎑Wy�GU� 3f�+A��n�A��#2��)�+����>���a�S������u�Nk�9��,t8h�`WO��]���5�?����ߟ	�~B����-G���3�_���6AC���7{��l���[����E�T3�kr�M��b�M-�J�O/�N2i��h�Hݴ����Az9+�!�(�1G�{�����?p_��\���#�[o�����Ԓ2�� 1�[��b�h�b��Kd�ϗ�dU!aԻ	��K^%5���<�ވ��!��8��/�* �ZAɱ]y�?�>±po?�<3�}�N�W,T�Ҋ�&��F�p�"�͵r���ܐl�È�/p����Z�y��3�T�3�}"�z *�cXw(�"���nQ��d���O^�@��e0����WgV=��,
1Ȅ�\��@0�ḑ�5Њ�VQ�n+VN�B"x|�Y����Oe��wf�Os�W��^*��\�pn�\�=�]|�66�jU�QP�j��˓B>���Fy���"��v��B8�x�^�p� ��3ei�3��Ft��H���r�T��{|�����^E��_�,w�m>Ս�L�1t:		r���5<��9���Rt�I��x�S�T�D� �}��TWM	�9(E�gE%���2�U�
���,�W8ۥB�9d{QoBa��{NP/$`}��0ษ�w�7p}������?�EE��D��:�Dx���O����$Z���TWeQ��vx��[8��[���mtZݔm0��N�5�i����5z�9�Z�2*bv�8q����t���ͯn_�%Iǎp��s���0��c>�P��s't�R}Zȯ|DP�$$#7����y�{Z_}����L �R^�h���"CB��:!�F�9cS�곕����_9�(������
1��1�;.m�,)d���"!`���d���gpX�E�,;2��܃Q����'CE%n�3 �`�'$��a��4�RCu��BĤ�Vo@�t�uJia�J�p>Ń��)���6��)����mƈ�WL���VQ߁H���0(7.��'�����Q# As�2g��7gqa�D�{�U;H.=J5����ZA�.��&m��:��\�8o�BFj��[��Eq|�x`�=0��𵓞�' F������\	M��Z�1����nH��K�B��]�W�9��Hۋh+�[Ѕ�R|&/6c���9�0Զ����PP*sy�M�,�~�P��9/�6Y���@dA�S��+�K�H4�R��e����sfW�">�R�fw��)}EYK��"_���~�(���P���ग=	l���Q����*v^�f�g @ � i��˅�d2��m�+;t�m��$Lg�a��Zv;U�� ��bm<^��d}�(�۱v�o��6k��I���#���hd�؏Խ��k�}��%̓r($mS�!�������[-��y���S.��,��?� p�Ճd1� OI&Ku�`ԁ`�U�, FDx��j16Z��A�9����l��/�9NӾ{���"�X3���!�?/z��T��D��� YM�h��O���`������Ǫ5��\ Fp*\��~|x�Q��zd5�����Y�9���W�c����K�YR�m��H՛��~�։3v�WY��Yr�zx\�uQ����Qg]���"V)������Q(�/�&�b��;{�+s�p~z�i����v��Bl���K�
�����V���s�ѥ�t�n�m�U�E�~& C_|��4,�4�~�J���o�d��E|�=�+W���|�_jb�=�0I�nD�������Ab�Ӈ�'����p�W`/�͙h"����J\�|�(t!e
��`-�
Ƈ]>+k�Mֿ���p�֪`���@`'�q$�'� 5��%$��:��Ҵ(�')������ �]������0�q-kmyRE��r"e#)�E�	]~�5���6�Ί�H;;�,�<�� ��]��\�L#�C��<oU�Jh�].��u2T��~��k��+�!e�m����xq
�����q�A8�~}�b����EC��-IV�-��,`�r3�^�����4%<Y~W�'Z��֠elB?
�����75�1���	���a����WI����r��"a.�Ư�A(�X�L����\�K;>bu6:dM����V�Ii�G��\�n=G��Cc?.�c�L̽�o���|��QA4�&y�az 8��RlW$Hut��m�JU|��z
���JՑ�7Q��'��IP���+{��)��b��3��e�8�����@u� vrf\/�?͛�n��� 3q��4���[���Cf�΅��/��M��=Sm��	L��̊�^�i��s邬[���J�3����]�	ƷiHd'&�n��i�S����|"���1q���j�´�cU6�x����a��D��tGx�������BN|F��2�6��dں6��1����Q���k��f\ȷ�� �|����2=7�1���V��vrM���fХ���<G�h��ΐ�!�:�,߉�1�u��g\��N��tR;
�+���-�e'��2���4�YB��Hcq��ll�l�E�,^��.�G
6}`�.+�>;�U>K�_�[L��\���;� h�Ԩ����[��\�xhA���N�P_/�:�`�t�~ �F��)X/B:O�s���3����mi>qv���.�D/x��`X��e�����1Y�2Ē������1��ރ��,N��Y
�""T���9�"A(*�0�"�����q��9�q�+6hA��5�xـ�E�-� ��e�FV�s�`�.~̙���R��i�
w���j%������Ia#�P��{�M��R9�::ha�3+���G�y�C��E`ؑ�'�l�T����@UA5ݐ��l1]ZQ��:�N�Ğ�\I��c���,�����Yj*w���E_���hԐ`@c�n@ٴ���6Z*z�/�3;>V?J��/W��C�䧓��?���� �+ypg��ܙه�a�ه��*w���g���5�\KYA�T���G�(ۓpo'`��V�1R�����W�bKǣ�͙���Pu8B�B�,,�~ul.O )Ev+%E�$=�'�m��i��?�E鴣g��RIﾟ�@Z�-�6��KYh����f��k][�5�.4C8�����	'�$�	zB"Hv9������u�A��U�ơ�Cd�(�nܬJ7��5w��I�A�ZM쀊e�>p��Ӱhɮ
��s����a����ƛ[-x�2����-4C5_ Z'!��=����e�H��jY;�Bj�K����?�D>֫b�ev�O�^�B�X���5���HZ��VfJP�/���J�F�7��Q���[� ZK��K9d�-^e�Z�O�#b4;5ɲ�q����g�q���h���%�U|~--�����L�Ψ�\�cI�_��}�g�п`��ww3�(qk����c�G �Y͍��9�a<*8!a9�_�A��2��ƈ��lLj�=z�" `�+r7�e��)�T�]sٕ���Z���%�ʽhO[�`J��L,�vxI�yz}�=8\����iz�v�CZ,R��!x6]� ���ɲ�Ϙ�D|{���z_�Wn����4l����5u�0`��_�*���S$ ��̒��f�
H��]n0xWC>�z��-lD/P� 4󗓚Cj���!�-��MX];7�%�U_�y�������%�H`f���!9��V/>��عE;.����#	3Ѝ���",ӌ����'-�� �`
�Q�>k�O���߇�aA7�uN�J��S������#����O�]A7��('h��֔����y2<sE�xE�������r�P�v>6spL���r;"NZe��"N���=��H�El��c��Fs�M�� eq���h�L��J��)��w.ו�Dń)s�3u�9���l�B�T$΁#�����&Z�T1�¬���sVm�@��1�T�&=�^1E�
]i�k$C�	ܕ:���aM,
�kD��r8��[��W����^s�1�H��'��(�>6KR���ݏe�L��ލ��09KH�D���\i�,Е�t{aS�y�)\������(�S�5A���p�"|��z֤53���t�_ܶ*�iC�{VeFmxn�'t�~Ǹ,1</.C�O��{D ���!��À9]z)��Q8�R��d �����а�x�*�ϋ=�+�y�m�bF�J��"�+�f&l���K�p��k6���i�v�Oh�A�Ay25�	��?�NyP��a��hr��J ��&�Fd�S�8���{%��^�?~a��P{=��᭍�i��I���\���Tsf�c5���M�{ٷ�| ݵ�E� P~�8;�MX�i�F��d��^z���R�
��F�%��B�ŭA�d�'g�ߍC3��`����%2N�do4�DB���2~�l�y����I�㉨XJ!�XD�s],/�'[v�o᦭�����}���O��p�0���7���r2�n�#e 8���������"��J
��B�Mb$>��{n���#�늟#z?��Qذ���.�E�W�>��D&�60��O��T�-]�l�0��%=�B��#x���Ѻ�=���F�Q���a:�� � )` �F/�������CBߐ�Ɛ�z����x���?K6���
Ʒ�<�K��qpQc<���2�S�v=_����a��͒��@:&]MT��]ǲ��2d�A�|^,^�w�!��L�����?������81�E��1WVyV���BN&4�X�¥'͆����DfO��]&��&"�#k������V�X�pD ���K��e�[�o���tr���91vM]��fQ��i���3K�3P���|9�$���AC҃��
([%n��f�jB� p�-�&���`5�;���������wg��ڳږ�:Z)P��� ް� L�73<�=5Ӕ���8�ܻ���T��BY-��顳"�1��}�w��D�;j��>����7�Yx�ODȧ8.��棞��!�%W��~oB��͟��8v�4gL b�����ɇ
����Y�bI,o��W
i�1s{j~E���4W�Z�@5ӏ��E�=E��V�*c��K�s�s�%{��(��)�[e�����p���}�����B��Ǒ��������sx����`����{bM�\�..0b/���V�� ħq
|�,썉�&qM,"s4c>�����u�٥��f���̤�g��F�[�>|�<kd'�,8?f�FƑ����A���3��+ab��k�����E�c��+2����@���k�i���}� gʳ9�;���X�À�s{3�ܖr'\�*��~�C$��%d�ߟ�&&���x�v��ďd�1�ٔ�s]V9I�����%�I��59OoÚ����]'\�u�!3���Z���-�-����;�lU��N�oLm�i@*k��	��AK.�ɢ��W*GƝڪ�,��I��g�����<����rډ�D\h���$�e ��k �p�2ws2)��uQ�	!����E	��7�P7��`�"|Rz�]��O��o2���&�
K�� -��������Wn�����N�=��ƖCX�})ZӇ+LcwpN�>����p�*T5G5G#Tv�)(Ͽ�*r��k%�@-�_dY�
��qU�j/
r�$�Z'�l@iگ��Ȗl���_���ق�|ې�t��̽�8��� �1�X =||�e�i��G�1�Bg���,5�E�%�ٮ�Ԣ�&���+��e�U�+��0K#�PP�$�8L-o?D��C�c5[��u�ar1(�H�0up�����M�jR�M��9�:�-4�'��	�����:x�_��֨�n�	`M�C���҄�%f$��]]u��'��Sr�p�_i�������x�A��G�+�4>��#Ck��` ���z�$<Jtâ�'x��-��� ��~'��  ����vSZ�36�xģ0s#E@B��O+���e{�&���s��Vbu�*,�q���t��=]63���������'��s/�-�>���ǵz�A �wց~�M<�b�����r�V��b��w��L���8�����β;����~h��n�b� J$��(/��4b4��i߬]�{��X�'r$>�RM��6�G�$dU��V�@��:Ș�y�	�ۯ��P��s���</J�WXc�H�l�y.:['��뿀XJ�|L���`�o>�s&m���2���.�a�F�SAGߜ�ȿ���#����S��gP� �L��-�tm!
b"��)}�߽���D����"d��:�'��7��-���!�%�|�ɡշ%2bm�?CWB{܆��.G�W�1ke��f�Ř��2�P�m{����-�~��Ƶ�6wɔ:3����?�]������
�$a��������*uͿ�(H��VQW?c��� �Gnל����@!��#U1pA>�f���@�-�,W�=��@�2�H���I��Z���9(uͺ`H!;��N�q����쓝z�7�:GS>r!�3%��~��1aL(�
��*�X�Pj6����6F`O�� ��vd�7:�:�s�f��K���\{��$��؝y������jn��1��E�U\��b���hԕ?�J�>Aᙼjh����K�Xl��*[*g��k���2D����=k��q���2��A�o}�Ҏ��+��X9�jɠE�<��n�p�lQ�y	�Z<�LC�I�xV~j�I/���d�.S���ڇ���4��1�֍�U��Ó���sBG�|7&û�`��:$%�v&	j��X�o͌�8�é�1�}���8�VjԎ��sc��?���8�z���#(eG�?�v��|Vatq(Ң7
�W�;'�� "�����mO�D
/�e�!^�>W�#��f����SϤ\��|Y;5͠��l)��L��;�;�ؐ�����
*�0HX�G1��ET�t���|�b7�9#�+���7R�٢�@n�@���,�0������*:	�]h�� 1̭���JT,:��DyP��<@���v%��x�������� ��o	��Z"UU���gԨ�ܙ��V�$�:���!f��F˽ h�פPZP��Һ�����=)������"�F= �2��Nt@ꬄ�Q1��!@ǳ�����j��_�H7��Ө�*Fz��X�</�gH%g�SB�Xؐk(��#H��PBsGh�8��n�m')����<�m��,!�uY�"C�`w>�GW}�/�-X�MF���Y��D+�Zm�
�:��Ԑq�,؀�Cr��{���Ѡ�?Q7�{��'s�4k5�
�7�9��0��{�-�D2�7�r�=w�g����������c���I�����X�7��':�A���g��Q�E�a�	۔g�����*�;�~�H���=c�NZx�EL,��`��.�=�7����Pk��a$ ��911�N��dȴ��!�OJ/�
t��26	Q A��X���?�*KȏB�:=�^Ӣ5F.���T��F�T��J�BzD�8�����E.L]�I8J������#�KR�G���P�W#ќ��y��1�r����Ac��
�ϊ�V\� �P)B����&���wLr=l��Y����C�_������de�c�o���_V�w�jZ*4QgY�T��M�]~Gp�}�� �\��VF$�30����n�16�Cq��\�ݗ�����#RЈ�H�����M�ǟ�9
�!u������&&92��rG���6���U��p����� �S���GL���������8��v��[ԏi��[�@��P !H�n<&{2�$t�i��/�;�I� ��(I*�㠥A#�z a��W�j�M���e��ٵj������k+����U�(u�N�bf�� 5��MH�7�b�A��U]p���=�=�0����46 �]=k�0��e����o~�v��z �_��!b�����:�����Ni���\�G��FZ�gD`*@_��K�C'h��]Aqw-؏`���Y���^����]�~�*����&Ypcg��Q�C*d�#�,	�wA�~<j�v��B�ߖq'�N�-���K?{��>0S�Vu!6}���>�q<�%�tÀ�w�u ֮���u�Z��W�������2�uzQ�ݳ���I����dE��i�P�i�h�k�5%f�m�I_b���^<��d�\�]v�%ըA�
�/�3�D��o���b����@j5N��
&*K�m���9���r����ս8�\\�\JAW�*����}w�԰�@.�d�����'��)�u&�LgP��D������W�Cɦi��A ׉�>�x5Yc ڼ��FTa���(��Pl�;��U/����d�_�ֱǜ���3|C���N������m�{�G@#Tw��qzE�4C��Pܨ󍹻����xzϱ�B?���ݩm8g½��
w ]GWڷ�����!�_ �4��M�gԇ.�H�'�~��r�=�����[)`k����aNӟjP��K�4j'�C̛��Zgj�A�y�KgTpi���e
�4����=Z��g���&�?K�U3�J�ɥ���(�v��ַxԂZ_N"~=�`Q���+��8HA �?pD�WNǦ��'�(ii�n�z����(���՜Wr�ń���\l��cM�b�I!x��
�$^�b�p���CeL.�6\ꥊ/�0�n�/��.�� ǋ�q�nGWeY��4Un�he��yɊD��v�eb䂲۷�j��ױq���\m��� ����C0g�u���Y�k1���޴؅�Ҟ��h�.ˆluIZ��{LJv�|w5�M*��7`�j���JD��_�x����[�_m?�G��+5���G ��1Ʒ5(F��q�M�R]�o�)��ы�,��zL�Zg��>d��18E��(�HG�4k ��|����Zd`�_9��9΍K|5;15M�XY�Z4U;Pk�΂�G���N~D���[��T#MO�Wec��M�d�=�v���G�{���g�$Ę>'�@K��0���m��Srf�c���A߷N��ɘ
���q!�v^����T��'>W����h�ɛ�]4�$�Gd&�'�-�3�񧺷����=�a>�p���v�A�L�er��w�k�1ۛt���g�u�6�VE IR./h���9]h]Ԓ�C�e'��x�-0������=������م�����ܔzW�[D������Z��� 3?W�,VIL�1Ù06K͗�Kr��A=Gd)����֫y��zU����0�d,�r��a����sG2��� ���	��=�����k�)��*�0HR/�̚��;���9��Iu@������vZ�{P;ͳE,���EL���3{��3��f(�-��#j�����u�]����G�P�1�*��^��,�۪p�m�Th�
U!�B(�.�d���9��ˆ�(��8���AV��]��nd�A¦��M��A�EݶȀ�r��hg�r1*a���0P�!�
C1ڌ���$���-�\�g���\�[�g�鍘��3
����w�p�ȀƷj�䨔_�ػT��W@H=X�<���H��ն��H��_�.i�����^�#I�B��W"n7	_h.o��r�=��p�~�$��dIIq[��ahN�VB3@)>�6�X׵<_>�ڞ�Lۚ����C3�5�P�F/����q���2��65ߴ����8�4�(�J��q���=����M"�fC��i�)x���҂�������Bg=|�/R3�Kˇ��=�O���_ޮ̟ὄ��*&��:�ز z(�(և03w�!��7Z�}�ңˤ��۷k#7�b��}v��L.��pW��ՆiV�*��w����`"��JdeR}�����uL�{���e���Vɧ���;�T��ߦ�q!xcI1RN5@|[g����]S��w�#���n\?^����vA�@%�S�.�Q��*�΁�~]�+�Q����%�si~��bK���5���~�i2��BRC�P����O�<�����	��)FJ�}��=�?�d�'A���v	Z<R�.��:V �R��W�0I˵EH���@�R�qH̎hCv���Vo.�=�����pj�R52�r�ta|����ʦ���ϯ(/��e�D�0E@Ď�2Q#�k�h�~��A�!k ��	Q��l�eʽ���Gu�\ x��Mt�����@��*��H����$�Ϻ��r�������x,r�~�\h���M��ň7�%YHo4ۦ�����G%*tS�@�AjE�f;H��/��瘙���������	�dկ��)h�K�,�\��C��v#Ml3��H� �JL5�aT�j�J��=��V[aҝi�����8�'��N�KhA���^T��b��0�&q��,an�,>ahYTRfZb�����o{Uꎿ	:%Y�ן/E��_Za�x���UQ�O���f�2ƨ��i?�4�Ze����E{_�XW�>�.R�����ar �`�C^~0�^�x��fa�];�>��A���A&{�$캼3���(�)ݔ7���ސ���$+��u�dz�����A	wG4�$� ~�����[?�h�$��2�M��R^'Q���t]�U�7F���C[��Շqz�jOtٴŕ�`!({�(�<�����/���L�A�W\*�^�����D_�N��SO	F�e��d�4܉�jlt:8k��A�v&����:oy�4�#j3�xeo|Lgh"&l�'�aꎪ_dy�2��������S iA߉PS=�-w��+
G&�DT��(��3�7{��D���}�l�~�φ���4��O���L���[x'����i�A�;v�N:�W�(�b��9�.�DCfV��,�:5�(�#e�M!��.�YoX\��>�[A�r26�r�^
��59X�,��k����z�Z"�\��j��8L���w!��eeC���؎Y�RG��׿H2E,�-^�� ���w~}�S'�	�X��y�@@�&��aS0����{��y����+�8E8�P�91 n��覉H	��
�K��Q���V�*�S]�����5����=��&��Q�C��D��ʵ���~�t� :ƺLl-��5�=J0i!F� N��й\�`����ɯ2��V3��Ix��'���aE�H�`)	/ �J�����y3���{��%[�99�IP���e���O����
Y�Ⱥ����ſ&�8��̲�ˇ��yϷ�DM���ma$X�7�ǟ@���4c��܅
MN^��V&Ҁ�'��k	��?�'����㰗Ї[�{�!���ֱꍟ7��Ѝ�����FY�����|�a�k�����p�fu�:)9�.��)�
Nf�BSv�VQ��Nu�e�U|�]���AQ!�}�(z?X�*ک�<�N�v$�-�B���B��4b�t�u�b/�Z7.�w�zcU���7���d�o����V�kJ�k�)��PZIf��_l����g��mθ��p�l��b6�7�&L73�vv��x���/��^��j��!��!;z�^l��[#};�k�z���}A�k��܎=bl`2H��i�gҡZ?w��WH�27q�k���
�R�[3��F>!��PSC ��R.j�3�8�tO|-�LN��!��;e�P�~���4E��;�&���VФt1�*���
�'�."c��`�V��N�h��0��5�qY������G�1�w���9�f��;4����������"�ϛ�,����	�����,z��^�`�
M	����	���~�Ju�>U�z3 �Ȏ�.�_n\�����-��%
Ro0P׃�:}[6����.�F���Q,�dP���󐟆��e�B��CG^��L)^9���w���rg��%&"�!�2\Tm?���'h4~}&����:Y���M��A����\�rC��0R��k����^��8�����1	���lQ���օ��z�,>(�'fIP8�D�!�Pw�lns֙�1>6��̨2�sℝQ�K	��p<I���SK�:�v
�ŹՐ��K��WY̡�xY�������!�^]-�	ɓ�Չ�TLZZ3*>ir�J�^Q9�e�.C�h/&q���2��Ơ�� m�"��҅�X�NR{^:�������xF)��3y���7�X��~��Z�%���^��I?�Vel9(Q����J5�n�"����,90�q����|, 5+�*����sQs�b_������y�p`�5�fAU�3��!��1�?��#�Z����5+[vp;a�~"��e�+����שּ�7-���(�2�Vcu�z�S܉�6zn��J�̀�����́�sS���<�Sd���J�E��i�� GU��O����>�ǈ�!�ԅ�C/�`��H�K�0�rg�x�d�<���Vg-���8n��h���wMAu߄=qH��v��K�b���+ڵr����7E�ܵ�"7CJ�*��O񞕀��		�a���;�R8��=�_=�®�'џ���:󌂃qW �э�9�C4��)�m{����S0�ך�T;
�F��NJ����R�_�n#��rdBas�ʌ���r��Zn�l�ln��x� 3�%�QsS����X��j)�*�6 ��|�H�.WuD��K�.?\I��K������;�Z�u��\�G6q�	П��!�!CuOo\�B�@��{����>SVx�t��G�M�V�ؿ0/��C�>)��O���(�M�!f�˰@����k�P> ��6�etb�0��"��w�����ڍ�#x��|���(�|}����,�N�	�cBk�(�r��i���nV�+�z�n��Us������?�8К�&V;�e���p�W�ً���j~�M��w��drHN�P�ҧ�Z�n;Ѳ�Όݷ��!d���T��g�`���c��1kbO�MS}���X��+Qep�q�.�Д�3#ع"�,u�2���璫8ө��Sr �ᖦL�cvc���)��l����-m��Շ'�Q;Q�7�$�}�y�uȖ^'l���6y&�>�r��Շ��@��F��3�#��h�N̓�ۓ"���+�n�]F��1�20��&���g�L�Ao�6`ȃ��ٖ3���q���8yk���W@X�V�D�ݗOP��(��f�����4�W�߹�`!���v�O�mɠ����z�(1�R��dg�����r% �����o�D�6^���p/w�B�� �G
c�Q��mE�Q���Λ��Gsۧ�yl������WS��77Q���.�u�Pv��bM'���'�Oݗ��'^�}e{U�O���A�S�#M |�	{��J����`m�M�2pE���������BMȖX� ���c���C���W6_Ueb�Qw���Dg��Cp����W������p�9u}����&F#n�e��aT0�0�H��!]3���$��ӳ	�"��3+5-�i�ge���cvY�㰻�HK�"�h�v�>7-�_
�0�)@V�pω@�_���a)Â�2���P�Ȟ�D���e�`�G�7��OZ�E�@(~��?�!w�&����e�F�t��Q��P����e����l�~�����o�%��D��������Y�JM���+�
���zI��4vrҒdo�cn��cD��;�+.j��g`_�0�vT��x�[_�.�|�~jZS8��T�n1�.���Z���ʈs/�a	-��Y@z��IʷS!��k�e��G۲Sdf�A��)h���=p�g�PJ:+�C�I,-��ɶ0�F~1��
?��טB"wn$����gP�����,�Ug�զ�$.1wF�j�ϥ�����y��W��S����Ua�[�i����&Ȟ�YD^��ok'D�wܥ�9³��$"q�y%��E��٣Ⱦ�;�g�T!v�G��ĺܔ���E�7���^��*a-zn��)�X��*���?T';�9^c�>�1d�g�)j	o��F
|񦲫\`���G�N?<a�����h�Wtp#(��f���*La�A/�3����_l ��d���;�����~����� b+�6�b9 u>5��'i��orE��lͦ�����4�QA���N�!nY�W�ט㠆��LucD_�X�d��F̓+5�]iHVGpʣ �R�Ti���`m,;q73
�8����5WS|��2�#�6V{/K˾�`�+�!Zo��:��!�0�����z�0feb��=Y�u��=��<�MYŎk?IXQڶ��Y�^-O�5��K�*_~�6R9����`�s�|���P��v�J�Wr����X8��Y��lO���<�ch�-_UƎ�\ו��s�VCJvK\�.I#�W�������a5ΜY�*H� 9�܇3�~��B��Z�-jk�l�PB��Ϫ0��0�3|n-8�sk*���
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
y0H/ZtY/Xi1SWF1w1QnDhbElDB/r+D12CFz0IRg9jYB3ktN8UeUc+3DrYJYUBQ2SDzVFqkLtN0ph
350H7Q7d6BYfgjcQaZil7Wj7cOLV3qu15nnqfvJVldrzyzER5zao7CHJYdQow75fb0JXFQ+u4VQo
Djjx/S1DjxCnzeHz/y/mdZCWEn+aOJw7cNeazpt1o5DjLYqxq4x8rISu5AmgO9zsVrGf0nWAw5M0
+UQ52yzegfGzk4JZw5Ez9Do/4uKRz8+jtuu1rKvGMKeYwpYK7qyOywUNrqC0HUIcQo0havI3U8om
Her9gjeKMTe4hpYcwTI2V+xL0FbUkUoJLitnig==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14528)
`protect data_block
RCGMLEMjTyKk9kIbMnJMO8q/CMifeXTjw6ZwXTMOxvwpHjIg/46piAh6xlmC38FUZFU88+7mgGAO
3vjrBc7NOmKVLAm3D5eWBbzga354VLwpVScs9+nhOor1uBlf0W1SVQKMmVtq8TU+yNnuL1GcRU16
cwmpEEGOBxbs1AlSwFIJ0HAWRcuPlvtBNasGxfZyJKUvRqZUxg76FvJ3ZF1+I0enyh/TgwzAbuOP
iAj9DRjBh8yYU1zSKC5purJZqOFMplK5hoPtEI6pdX0vYX+KereGv1G9eNhJAg5PpKYTwHdozvV8
LBkRtQW/QpAfwbxTEnGvJyGHngmt30QbxJP3mShBUcZZaIoiPM9gxixniXPwASLEDpjWFpBevh15
M2jBs28WWTDX7FgEjqgIviy1RcRVCt447i/Jxj24rx+ouyX8gRh9O4D4L0La6mi8DuSGx4v6LEe1
LMyBloVENIOnFVonV5w/YHZ2sJ8Xk9LWEltrKsh/ZUdp7N6W09Z0gv5MI2w3dWBiPAktyD/ECuNB
24tTOAhdOEYH7zwYjmiKEbmOBlZ9irT4NbsDqxjtHRfKFJWs+mngqh/9b/0V9di6HFUcD2GACg4O
qYpawTHK3lZNqGoGqdasfnGcZ1VCNryF+uvGk5yC4R0VS7hs9GCRVfNOCzZHFBM6W404ld3ZBDFV
Gy9nEX9MsMELX0j2SEfzhHYsD0LFEwoxTkRow0/p7zaGfWbNhBu6Fw5gBYT2Ja2sGUSUkKQiExPT
GREaBEhePuOryll1lWwD3PP0+NSy9txXHthxNrJnkfxaHwhj6p+dZSD7ZmNMhs92unGI4dZ3Jzez
Ai0J8qQPOxL5pfL9JcPOAOKmyR2l3d14o+dJkP2DLEX80bwbOa3M11mem4mqhYLw83I41VN/zine
Yu4D3we+UVYuQAyxRyuRYgbF0OI6LGajZfwx3U+8Xhsmm7MlIIkjEdcrd/EVf/fIcn76v+1pEVe6
xoPSan3yo/gyD+10AZyUdTKJeelC8fbo/pVu4/R3Avc6ags0rv7Et9my0nZbNBqr0BAzDQaXDShe
d9zcbG86Rc44S6WFJHWnAp3hi1dbjxxLTbyHvOvg/COdlkRh58AAwZbREZ1XmJDJ8ksNDfgI0+Yy
SqZgXYpsVe4z4WYc7LCm+2fzGo3A/KlEsc96kWCF09+B1UU1mf3dFUn4zJHecK7ziVQiv2Po5rHp
a8Qwmmz3P1mHqomEQ91RT33UpNBr1e+mkgUMNPWMyvD+TFdTXwsKT8yKoXv/nVbPqdgkgd4MySbZ
rzmuzQi7gB9tFNBF1fWX6VLlKgHjWYvL6uFkhLuqvM+KmYjyarnTttkbYsqUpr1CeKI5muB3iHQr
YqECrOcT8nUIVFn5dtJnKnCiCgW+FgDoqT5eZY/lJ5cr67rTVQr4QsG4RBnEZCQMyhN2mKt8UCWh
R80SAp426AAPlfGA/NXSFL9iBX9nRiJELzwx7WQmDqajZyIfZfIP/xDXyXWzwnXPCwD8qK7YtCxf
FzcF4bXUGSsudxTguADB3+1NlXkOQgLDejoQGjjgAjt/iK8ARIVgegFX1J/nz1wgkvB2/fnUuMc8
o8IhC4D3EGnirTgYt8j/ct/tYLzPB92CTY1rytcYL3BwmkBK6+kaQ8TPqr0HysbaCl8el4n70hmO
WvaeMfAbHHIxcjfo0NdYdQ2bpKkOyfluPSBIktsUkOXVAD4mcSLwqtM5wy4GApXAXkhIIae+VEgt
QX5OBiS7D/B6y4YmsqbUMx9B1WkKrgXCW6cTcm2NS7B9dO9rV41M01WZG74IyArxFrG7Atelz+LC
znYy5skFcoR6lPr0OYnNJeNSKo6l1Ds9Yh3HBwSF5Gw6B7vgcdpMGO2b02q2fSjjhZP/GbBMBZir
H4HHb7N4jEIHN3ooCSDE7VSCxedJtI76Qo/WEgGo31MGu203QtfLtVUwm8Jtw6lesLTirvxYr3n1
fZTXzf9g32B6eBOdf9dSeKoCVWHlchsurZGpp8pCO/q0L+VPj5xKLppr+/WKRufN+MsOgliy2Ml1
Y/GD+yT7q52zNbXGD759v1xO4hVnHU3ZPB5Plmo0tDSmvEN10TuJWYHQ5ZRRJ1DMbaDoBfj+9xjw
B9f2hZxhB3brfEGka1GuOESD8KMmCHSruZTJPVTD11qzR/NlBHDy62sStKUSDI9Q4kVxP3dnc9Co
oree8w06gll5MCDskLvwSS//NygnDqQo084xf2JsPSkwGq9b92A49fILT45f5YIs0NYt4thMiPWw
Ebkp35WBNJJBQOV0rukbyBkdQw/j4H1DzIhLqAexAg9NZF+rZ67x/i40UOq5CSAQMihXip7Mespk
1+fdGsubzpCvuKDPm4ziZZe5Gf+CPmyt2K4zILccb5VUUULR8GY75GGyRpLL3M57AXcNeam7syfp
hMqIfnai3O9nzWizQ1r+7odh9gtgZMdUHnpe0uzlieEFet6X5JGU8tZ0vptEaClIM12asoyta/sa
XiLb/qMI3kQZy4Cq4g8n8Qx7rTnlCP4mJbDUPxYaO5ZdnGejgjUbnB6XeGf9sMvKNfIAxkCrdC1c
LR4MtUGdk1p4aLLMnUIToemKSHGJH2QUNO4gmp+fDYGCLZCe8oMcoyG3JdVlSCYOiz0y7NhcLF1O
aohDDUUax5MWobjaDNHf5APcRR85+JcYTpcX2MoaG05i2reTGF9Zt7Y5yt5ggmxAgB3uh64309aU
wexHzxfKL/KW9cW+qqDbFJW0ts55cX2AfD6lNiUhn0rnMVOPR6YtRxKzsc95kQCYOaSiVGt3rXCS
2bEJTbxO5ovbbAiQ+xEM03ZdcjOvc2qo44PUBoIOUbHd6+vFldWjISs9mgOXf6MPNccTw+e+A38e
ufLhLNcw0KsaGnE+Mp4SbO7wiqsQt1cwY/4Wv4qm/cwSTNB1wV+oLUGxCXLakMcgD8R2hwEPjrMf
G0iLHGW2ZKOIhPchNlU61PMLznoA9bHx0ptGcFJXFICoptVQedznX6J038kVLgyl7ZlvQvaifU9s
499MVAbKjx3YlVPd7jPXCmYGyRgccbdp1q5L0sl9lrAsZE7U/q6eSfjBbm/BEYNb0xWHOtWYFnKo
L5QEOd2YzJHCXFLXKQpqWrlAtx7B7BeRNIDKhRZRghAYrRd51Ygy8g3H+qjTMsoBj3EGImLUARUF
X3nNPgZSk9qIeX+hzHXch4okM74pRpVwor3ZahbcgSSb8OyQCQ60t+zE9wPCtt7BD7fqFLs2dx+K
EA9lyqdX8wr6XVVS3Ex5HBz8eZOYcK2J8AlogaRQoyLV2TzwY3RZwQcQe5NtBHEzbtM4vkc5edxY
c0w173O0WEl+i800gXyZuN72LDljar4uORclJMLqrkWSXn7BoaJDeeVNyVFAF4x4j82cvZoP4ZmM
WVSnYlDZ1yoPWLvS2u2iSACmj/vQoflG87PajRlh3HySDVuhFI355nyQRszDFEaW+7Lbo3VuLVq5
YlobzoPlScZ+ogDn+4caTwqQJRgFDwW1dbHErC3Y2Hi/20cUWFsHmlo2s1yc3RHmGM9HoAN2EFCe
6g5UqUF1E30ibYYH9FBvEZ9riMyvm6kJy7jWL9edIR+dJRzyi0s9GQNARBqT+RpZdGfunorTznHq
TZojnzMK7/k8ujoph80jrPuNdrvFlIfCeDN0S6gnJjZJIxS6xkBhXuHTEXRxESbzxlNKmtN21AMX
8/EbFBrQSeAzXoU7qkLn8wTEr/gCoeR0y2utVTQ+tbJLrjn9B0yg6jLRWQMD7rpM8auDn1zImwE8
FFC0QsB2x2qLuvLoiuNqtRI2SZxw2IGpl+KUkyaZtCIAmMkMqS9yRwmCdEYKux/ZPYLBF/e+LHnq
XbcazXviU8FL87mEPp3V0zeLgZbi5b0MEA7ytBN9qP2E7X2lAE77ocr5YowhuXJWcJzLvh+udrUU
C0Mk2x+G6O23bzJz/P2ADKbREUMXhtEU9zVc8GPyjlYt11KTinz0m7m+mAHPhYlUTsuEt2pcb4hi
WQxFwvlIjWaBcKwxiwW1Ur1M37kXHUu9dkY1t2XqBSdQKNEJn9e/0I08mAJblCWFgn/vRZfzuCEX
ayrP2AV2jByF1p5xW7XapuMpvADImxQn+DtpPX80v25cySla0dWUV9SeXm+czYUAJxxq9J/TcMFb
sBpGzScWPIgB86S3gQKjuRPmJcf1qLAsqmAOuJHojoAyxBduQAJbFeb/j7FwWzbl69KSESzaoXMg
pFqrHN4XTz782gvEjlmrk1wxHYRc7l10lWX6Y0yGGFGyj+gkyEkZeilPLA/aJ4L9DYwP7LrVGHrY
oE19evklcZC3EBD8WQdblnwZ6whigDlXezWDcMRpY/BXKqITG9hSuzxI5/hc0uYRcE7cMBxAOp8U
GLtGFeM16Wf/p9fT7x0717Qsn6bGah2+FZDAn+ZFW0jS8i6sfpBxfmPaHzDNjVLkhCgTTTsJcLNZ
7gxdy7F66wZxxrmRt9VATLfl5yWVWylSnSJpoaj70grpzPZ/mvlpqABl+oH95ssPXFkD7FbzC3yp
TSeLA4P0R8EE46S/6x+FllxInnXlSDpiJcAIrMvagvnqacy7p6dztq1WmGDnO6JewhKep1WBu8nw
H3By20/iNywilxr/+dYGkkzcM4nGGWWiObtILtNkpTVv/hE50riBkYnQudhqyqAvJIPay2wHLtXt
wtjb4xXP1LzOkVQou6vTAWAzIcK1xV0nEOgB/Y7QdF7bHalhAcSPM7zDxIKxs5/ced6el4IIFuAK
0F3DCh4oAemowK2JB8hH8xmpkq0QjZeZR3gkxJ+7qiTwDGiDS8sLWTC/KbK3qorhFTg/S5YVafSP
YocYFe+yZt44IEkkx3R3uwn3iOYU/rG/fyyqtTUkdyBGA0Va+CxcwPZhGH2QsBdbng8yTBi6XyV9
gYzlk71NjcYm0KW/5erpCpGJL9nNP7DG/Aq6QdqNbe/mwyCsWRDQatDw3ys3s2C6/tSItiEDdFD0
LFxw5Je2Mx9/6dnPHCMGKF8Ya0fwCfPEE+lXhoj8s2KDJF/xtClTVxdbaEfEOP7MsH0Ot+k7+4/L
6AnMzORX91TAPyui8hZPK2C9nqJWO47hP125WmEX/lCGKcjdnyRoTu3036vJ8nLxu/t99F1SGdN4
3Lts1ipeh/hrQ2L1msSANxa/1QgIjNSOibGqsYzi2ccBsURwnQiMTcus1uKDrOgOHL/ydznwOgO6
j3sRlzxCEsUWLcRyv1FkvlTskwRY//XuiqLR0ZBqun7cXzXM/oyBBP0BxoH1rXj/mdiOLGiPKIxi
Wa96uAcm+SFt4E9jsxFBhyQUkrvMs64iu0qG55mxlArvOTVjPrwaBTGuz7La2hNqvNgp9noFwvTR
vfZVWbAKOX9ix+68mBWeBPcfVAM9j9P16OcR6i3PSMGD7d8a6owKmXUDWasr4PxnHOgs6ar2WzDy
IgMJlw8eV9PXx9JwmAP+J/5fP0K1+4V+0TJdbFgku7jq0iu7Xko1M4UrgSSdT4eF6PftGDKqYoQW
GSOmXKqBeoqH3jtLsUVh3lz8OdGwAEc7IBM5hcDxme5A2cSGO2O8OYQ+3tYq7DPHlfVfIqBdFLHq
n0ivdEXxxeb2NtYVmFBpCX3h4L1N9cb1skUOAZuGXgjrFFdF/bGt2T37HMNUsBDlkRYxNjHtsDBw
GyBwBNZadike+8cJ9R7tv6Nbk5R1LsEdYaxCrf+zZFNHaaHQQVqTHVTBxFPIuGDNMmYK/n5y4xpw
e/vsepeHTd/XaJQeJlnCoAhMd9/3YgLf4w7xuxRU6z0ziC9DUIPJXubi4hTqR0WCYWL3BA4Yh5tF
FvG/B504uMBbxZ/1ClAbTq6wec00X2acO2l1RlPF1J0l+g7cYtYpJ4M0LIY4rYU8rLWDZVuBF3Md
Xm7fzPvO5fFGFcaxF/MpcAXn2lg8OlO2413kS8/8KAYMUa9I34aApFfryqck+ieoMSlPNR/FW1Nh
olPALUK9AGygyt4qsP16E3smoGWAel3uEYUhw9U0bBz+Sa7iibRlPD61ulQe2z+Ol3+DcH+6Y7t3
yAiO97XXQtD3AmFvqHNHsGDUUB5eUx60OD9AewmWnqenE3DnXcDDtmnEu81M/jTe22LB9o8q6F5h
soE2M2Js7NpR2uHgSu6OilrPD/9K51rl0GTa9zUp56Ix5Y+wDt43RmvBKBF2HXLq59XPvdIfEWGS
top2mAXcY/rqVGpjFaM1pMqvnJfOkJRxEhTKYML1B0EL/+vscrVP+6xVcl2dagLRwyC6RKx3s1sB
7qI6ZW24T1No36L4xwa6ImAsLk+xuXA4yG0Ej2TYjxjomCNRtJupIVM1ZcwvhVze7ql7FQLRNOPg
Q30+9ezOQ4+bNZ2jGJNhYZcS0NOJ2We4LpMxr0810Ng1gY/bHSRV87C/B4Z6KqnhXNqFHdZx+9FH
ir7TkjQAiAYCMgBMPmkbO8IhjVJjwa0hx9yp3LIJHigJ/8YUMzX37OdBZUsVVoEPFsg3cQJW/2TF
p+lNuoG1fr9g1/kOX80X8snmvpbjQKiJuwQUHwTR2A6rd/nKHqf6rpDLDG1OBATfS4iZvET9Qi9F
HY2LVZTGSaFEClrRRfqNwa5ppHYUZw/b5cXX7uiHR1C/ig9K/iMIRM9m8+FIAySlazWKq0s/lleE
AxVo4oR4EKkMBSKbqS4xqgLNlPQ8UzpQ5v31RKVZ+CTbNLQruj1CgfLxJiKJ5fHwQwkOBo9E2fuL
HlEipfsdyoDPEnzRQzXOAE5Z6kx2+XA7WHT6KcZsJIG3JdfWm9TqJsMy7GWEJBSxUy6G+TfcEC7R
iEQ/ZApz3V5rpQ83cCYLpPLjpPEr63AcOCEVV7fBgKP2DidvnabrQ2lVTWi5ZC7RScaSn9IIaJ0W
0murrqVrDGSUZNVhQ8S8s5k5cD8vuxSgnj54vCfcYE8vWRVHaMleiWMzpm0jlh4T6D1RXHHGhaOp
fzdRENXxoTwh7izcg46wrCLHKdANpLhHhQ3K/Az4//DUzrhkDBz52upMB5dD5a5LmjPJtAFpKiZ5
PhyTBPwHJhAz7d7Z/i2K240rGoch0ZlnVOGvGQG4v6NZArWh8NIhkdSv9VrTCkjtF4L3qCz686d1
hwe714gaIZntX4qf6uU+8KcvQHk4Qv5WlP5VyXXSpviYyyCukVxx0jhPZIK0qt6I8T/j8iGRFcUw
fuK8Cz98ln9keW2WbABxq3mxsATaoYLqwAO94Ct289eruUzsT0jJZXlFz9QF+BAcwmfSFDvAskkv
VXQ05S8Eah3QiH7OAh6g1QG/2ROykJE+SRMDe9CfX+IQq4UACRRmEe/is1uOZVxUdjeZXAd6nClU
nTPnxkiJtzx9tj83/3Ifkr3tLuIDU7GOVt5WEvKm4eo3sF6aInaxNLmzI3lzgZ3rN32+6vpfgIca
9dXUpT3SYb+ClfEhRyEG4XtwKLhSx/0ERpjIzNx5DpOrpBgvy+1jivRrnVPQGpT7qce4R9B/wf+z
xOWPgUiPT4Xx3TGUrCGRPb9Or9b/hj8O020sIPQ7bioLRmBMgV/qk+2KSHJdLGFdJ0iSzDR51Taa
gJ+Bg9IMS3RBlNLmANCdWL0h8NlHdHtZwibuAmD70i/Zb3omihkZtKQxL/s6nGGFtTNtyjaMzlKK
8QQ8p4YqgvZkMqHrz5H0Ao88CuOafFbzvTre1HlBzimV54INQVL9Dl/nJCmb7khSlLBhu6BCoUI3
+ELI+Edq1Mgx9yOM3uqSZgHFegGxV7fKbH6xcPj/TqFdkYDpYH+ZKnQlRORPA85OqpyM9LVZ8/UO
3W6ZmO/Zu0Dti4gMvPtQe7mYVa4FFjcomFSsoSxDSgWUr+iOAFxfRkzxwgCRHFAYKWs+I8i4iBNo
OdRC47SuccIVITn6PFxbb0Gq0npwj+s1pwYV1SNvn77+I+Lpl8+FNfPhT5I5hg55HgZnWJcg+a66
As5/vPvDegKqGdVtUxOsi+97B70i3CDQDqN9ctxO2DnwzJvelKKdzIi9hKlDTj+RuiZhqCXMVIyJ
jQKGHX7rUzWpHisEbxYCcmpQ6Mq9zBTjBYMRyE9VbIAYsDYw7NTZpfs88Qp5RrO3c5Z++vcEex/E
WCloW+o1TG/9lIUtNW6GSyX/DuzV6I5jCr4VBeyxF3bSiay13oHY/UNBOvW9VbsPbHlrd8RyRKRz
jbWE3/uTJuOKsEEXopMotaEeHF/1p5L1I9OSiE2k/Kp7EA6C4mdle83IchNev3Ee06s50LitDewo
LLA0pe1b3wZpxq85xg4S4M41LKoYIdptTOjWwTA5IMbNM8RpuXIT0I//v1QIL2aD5HwmXt9nIHvd
ZXdFkkBTXJekLqH9G7ZERt91dhSaaDo7874bLqY4O9d5kEuoH24+conZF3kt9r3wjmen82FhRuhy
6UaAr2lGrsPVKiZyKmFips+lH4HfAQ6QVg/3/DOEcMxKwGUZmYGIMvuXLnd9zJTF0MjEDS0aqulC
bVeybDKuLAH4+TCq+MaJHqGptH8n97M1scGLryiQrLUVymXqu8pHU7g+7AohqIdW6vjiajDh4SGM
FRdOHIoe9td7ew6xOk73Vv2dtBPWdwOxwMjHzvR7x28N6/CfxGlIjuTLSR1cRloLKBGD1Jt8WHm1
7ORMMO6iuNKhJIqBlKmVDjwkx4zyWPG9FwZOmwPOzyyhVONyjPtII54YAOXthnkY8O5CJnmPSs7s
vpfZI5+eeLS0em6bbYfzCpwWpg1GhwcSxzef8C+Zq0KuA+5c/mDxEAnLtYzYfqiW9oY54kD6txQT
hLgQspdMsDLjbuCx/qrA5bAZEFctwuTZaPMu+JxkuwuitBUCxi+qtDSBJvF562Hq1OXJodvAzpxy
y4ze/ohYAKZJ6tTLqm5+NCV1pAaF5Vqph2pEpSpoz7NNAyLjx016ASpUNO/jxk/5/ax7QI48upvH
5w5d+sx7riCTerL+PagDMy8Gw1uAT8U+RMXmi5lNaMb2vyOXxlqOzfAoFFJDdlejPCsnjiPiMB34
uSwE988L3yRdPZTkkpa7Aj4u7FAa+JCyN+5BdKtoE8pbaj6/HoTtXtlIYcYRuGY7gIrhLTX5nOSn
qcjk1VdDi5b+DAT4c+sxKgRyVxMjDTiQ8KNXGoQFDCPgBe/jW1E1mWOnuPmAHy5red4IqWah4dcp
BvhNl/DfIFkotyWuR1LdUM0sZHM+WSWtelh8fKbElDQqDWVWfNuJiekUvl2JDS5VHocgeLSi8goD
BgLgTY54q2EdCYRDYn5aeLhoKCgk2v5X/kITaTotHfFufsc3mLN0ERmBr5OCbBLhhJ2A25P9J/Ov
UX7oz8YgqJzcv5InUkBhCO02s+8RXYZU4EioW1ejvagkkVAA9wkmjwOrckhqRrGa1aFH3eWOmZwu
cZIFI8gKsDvHisemZH1ndnUyTGU9PdsyzHpg6o0ok+ShyM6JrKMoNTCMXvgnaCLa92VW0BEAhnbT
G5MElcGbsEDuA9OpcU12NukKn+ArktV6JncJZMil9jEVVM9XlsvUHmasqlwOqXVJyqxT73xQL5XK
m0M7jO4XqEpMqZcko51VGJCAThVqN1OJBGIv/o+gt7lG3LYIvKzH1NsgsCWhaDhIz9Iu7NOkYLUq
84OsmXybtU16xcCURwTomw05hp73PStRQDPh1rFGmhWIv0bIUZCKb6tcOf+hk+l9pcRKj62doDJP
Idi2MtxbTI0chgkgzkWj+W7pGaPe8HR9nScybMY7oI8U9KrnQCgNyHyzvF1IsYMUCBKHFUcvOBRW
Fy1j0S6RVjHSSPD5CMiwwr32C+gLah/JxaOfgHtagy8A4wvMbceqQ1hFmtq+NDrKPV+l3fdQXcKG
AVKGERCijZAZV44fJvnchapyB1BxG2NfP4OghvnNZFyY1G9YqlOzsf7RieU8I+KmrQ1s3sB0m5FD
HgjTvPv5niOzRfVqLVyL10L7X1Y2ChgwhjZfiadPH7mvmH8MAUWY8+EYroxOAUq+c4/cj93zCaAp
W9dRDxVFvQgT1ZEqChVn1sDrpdXSA5YPHPEAjeR2XVkq6SfwkrhHt2aOKW8HtxwX3IFXQrGqwEgU
W6hPfT3SajJEOYKBbaSLypQA+6HntTy/84Uv3I9OhHNcQuNmAP9xMxQCflx/LKU2o8b2Xu2hsqyE
KX0ZFesXp9mZBxqYQLzULsymr4g7ms5WCU0UNnySjYVZ4HieJMxGiU0uG+ggyvvaNCSie9T1IR/m
+bT0gwxCWzEyxP3cR5tElYqMgcqLvhsoNr8SjcnBAnTS6LSr5NP/iyjCo+/z/t+HTDTl5RPyJi4m
+Na4+BthmGjOFFaCOX/zWoepzoVcJyWd2LnObGPYDh++zhfZ4g8+yTtItpx6F/7K6E0A/93+qGvo
O0Wqwo4nXpBC0cSjAD6Yf31+8Lt8M2Ez4c2CUHwU9TehRp29/B9CnpcMTUoD55lzOfG1TM81jkwb
IIlT4x+ygkyaKj3yZRRg5YrhfKUcOza2Kg/Yp/WpaIs8J4goBgrVfn7CxJVzCawOqHsyvYoaa9jI
NUgBT2zNEY0ix5opL2l7Ic7MH+gNRKudviparjM98bhRs9bXRTmW2oPGfWifp+FIq3xZfCTGgy6N
PcGNXrmDHS8htBRa4eFZBxMOXCFDgacbll2ELpOPHAJKtMkOiZniFZJOJAud23XEUmN0Rb+D45VR
1CjB5ZLtm0hr9Ps7AaEl1/R9oBxktlxIOalX3OayxtA1Hn1zZ7+J4+eb6b+qv46NigQ2aPNJUzD/
Lch+sru8WoHoLbK/fnRbhIO51mLaj5cf8EYXNkhGizIAUIzJoRwzUJf3UOeMi0idKB7X8P3BCbBP
3/5hK/wPqhgRK16PJk1jGGFGwR6PnDUQhIvjErZtNqLU5I3WvIgWUiPMKyJDvC2hKEH6NjMRZshv
Wwt5XeP3UvLabiRcoZ3yWQXhaQZJQQJePAD8zRLCWXPEvgCuBF4al7lFGMTbxFinZUCTLHjktmTp
WGzGNLjNjKNQHidg6StlWxiLGRIoJP6jE5McdjfCPQh/MmO4D7zQ8uhkFim0Lg/s8HaleQke+pxU
xKilUXZJA3B8t2j7CbQ2tFlC36C9p9Muh26m0xbIr9csoSbI7+ZmzeW6yMMv1Vu+ncxkG5ft0V03
o58aPCOo7QeUCkYtCiGESZBqvzSqmu6OL7kNon2q1NyEC46RE+AIJUYKEGicARjmB6LGdcLyO+v5
5FRLZkf1TCUt69ihKTKOhsVdFeK4Gt7N7cH1wTPT0W3aSdUX7AK5dg8kvFV1tVQYsFP78rKYvfQd
SHev/OhumRmEC/bPefquHkC5GzNkWoYCK/bErS4R3Ug0vT73B0WS5lJgYgHfGcVsWqFRE3p4Waat
Ks/OGPzXadqxVXY5MKafBxSnL8mHibUpu6V7r+S0f4vdf+KWNoLI1J6dieqLdYz1HyzLjDyOgR9U
tiF5GlyvEDnfbnTF5X/e9+Zk7GQ0m4L+b+XFMgR6sBKvSritPUqCV2rNfeFDBw19TnOFj16T0/wJ
JPT/Rcqp6VhyLZKHNzUDAaRcdEuWi1exs2eA7Q2xDsBT10rJb/AFAu/OJMT2myqFHJuMzk3cW+Vu
A1uSqoEl+E7eK/kwO92x89SUn6OQJpJC4VgQshlWuSsm43p5Asms5kfasHikfGNDmKdnOEGuZ+v5
VZCINw4m9CCoxD+zKZ9O5RbXRH+zfFY0wvxNkq7KWKqCkwSrrvwgGjb/AtMg8PxCQSq/4yK18YXn
LdFvUX3pNNdJDeH16HHwdCwvkmOBESkKQ1E0lDWHIzDEPA7ByfKaBrZX6M+XJfJW5949wpDaglyB
Xgh34lKi9E6k3+blqiXiE8ez26nCERm69w7EPO2jWzC+80+q+66FsE3o2d/JDC9y4Mn1im8zKfaS
LBmppjvJrtp16q3Kvyri11gCeIIJyLz+G9830NFF0/A7X3osGlkO+kUkeFdj59EEZ7TJBULKKZgJ
KhC22Iopk0QdFGja7VG35hOGMQKoo7Ynei33yfNj50exaUgcEVRkxdOYT1qX2q+ccOSHrb3ZLfQ8
gGcMQ1HdSG76giRa3gnZvzp/0hiGb1mO9AlxI/3AWCP8PfjsUV5dwrKvopZN7DtWs8zoA4L7fpky
j4u4o4gMu8ipxaaEaKdP9bYsRfzpOrMBNuIjx42kVGsQ8P1J5Lry93ySACGgjWbQsP7B0uQ2scLs
MdeBDA6REYrNFB8YGZhrh2qS2KT8V8bYDzDcrfFh87DHraI4tsEubq6wBIeV4prAVHALMOv8zwuC
DiVKa9IXFNe4VCsmAJmhexiLFApxszSngYcuPTB5ICFjbtUBsR15aKAlV775PMEucH896kiEfSsV
TZxVeNTkrcF2u6phYI04KXvqazxMlJC/RYT6m0JiRNFZSWxkVVRMv/BU9mH+AzPK3xnoQkQ1H6PS
atGRhKBJcwNIMO5ZpPygaGsfCC8tmnkEw15CG8Y5Dgn5JksoJlH1dZkCKfiH5OWGadukzTvS9sOD
2Kqqgerw5xH5UeY4WI68qvM0/VSphQrF3HYCn8WU4jSAik5XJN+PDsagL7DRCkkv7jZarpj9aTjV
oO8nFhaoDzW8w1MLG+QEkqUvKsOPqojo/RaSmaKvE3RlAhkbutGgucIpxQr6hf8avBsWqp2eaDxJ
BIzz/W5prHpYciDUzxGWRpYkVufhdoCM87Ge5zEr8oPIQe+f8ytGA9j0T8/llnW8b81vSRhoN2Fs
atS2uSEo9u7ZODKmAB60ctVW4AFCfO9GWJo4F31AGOyD1ezs33oAC3X9PfxpUZkl+pK/o9Z8gIij
OpLj+6HMztf2JNG4F8bLp32KGsCY92j+aYAYTuuVQNook6SUCNg7/FF6AZp1tUH9CdfKA+FrUx0D
/vkcxVSFFOYeS+CgNtecCZluB8lZR6XmzpC8XPKMOcMSe/o9a/UqGH4McCMe0+KQMSmsDNXSDidw
VgnUIFd50zFGpSr1pP9ESmmhTjOFjD6Cp7OJJoIaJml7/x63JjGehltYwErSIOg56EcfNuGeX4Kt
+YE33XsByfLYCAdSz5hCHuVpIN4Qur8fnL59FYwG3f5AXYoCBRZ8Zq5OGvqRjoqp+7jaE8bumPgB
fDH++iudlQFU6Zk0l+yJocmXIbZPoZiZbGMsO0x6PDwKvpXgZEkoGwIfnq1HKl0ylpSxUqaME2iL
9AMtznuZUITFImcelBL3jklyKlwOaXRPQJSopAoZTTjCpNzgSjZnYymZhtvpt/TYQtQwFtGCT+Mo
j1t5uufSJ+jjq5G8cimHmCGcmnbvLK+3Cf3iO0Sqim9TZjUiQvfJYs0KtB1V4qdRiz/FnejccF19
kVgU6miSzyimT6n6ahAZGJ8YsxINC7Y8fdP+o8oKJqz0x/Tbz56rwMFEIgf8W4JVMMq1bbzlJnk7
jKIrgtjfVyExiN3K23zHbfFkXD3nQWhHjJ1fDYIqc9bsLSkD1lIgG6y20DvMaH3s5KI12g8sZ4/m
Wk4BV0V8v6MCO+v6FZP9sVy/h9pKMfFnQedTKpuaOCjj0ErYPXeQi5gK61gah4c7RJsEnuBbUuYX
Q7x+JjNVuEVWng21CgdVP9fhzC99nrXWmxD9JqLrWx0n+MFnrka72l73SK/or3mSU/VQ5DjqWxuh
BTE7N6uFuaqd1NPZTO6i64DOih437nnqkHRTzWRutlNB6xU0SDJL3b1E+oim/ZnLGpO0FeBK2XYF
l0L5bKs+LI2Gphe+lpEaFSvMuTYkiDgasTf/q1Pq/YfOuWgvbu27IWJn+oK7CU1g1zbTWuTUhpqY
1+ETwvu46XnOWtwFncwV9rWD+CkAVfONQh5cN6O7+ZPjWYTsflMSfcTgZ33vssOhXfLfBU+o1UUk
NHwvc4kP956XjOGuLbFq4hK2xYw1gEMI12gPC9xf53DTKILLyTfTxeh47COOMU77sJOX0AxDGZYm
TnLNGpFgQNN46xluV5wKl2p708YPiCPIBA+BBADAYS+0GlxNuUzZqBZ2YQJAyN1OZ+2uymRLXDnH
4KBfT86FP0XwMtGFxJUP/iSgcS68/CAF4e2iMlfZ2F7jIGPJ2I4zhuIbDHkhNm73uSpbWq1lFlHC
K1kfGkIhPI0kKVv+0p6S9ubY3wVoLD71F7IOfg55bqa2oeXLdohbYnXBWETpvU4gP6rcpM35D59N
lsvDD+G6oWO1nf+4JFCxuJqhXM8H5KjnHGMGJMc6OchKuO7j8iLQrvkKp9b9a1U46CRTcrbQHd7F
K5HgyMXI1z+JC0cgNDMcV+y/LI6Y5cA9ZHG9m3MNk3Y9XOiu5hDW0fIYOZYDWx7ObpR20u0Liz4o
pul0t4FDr/oFaQ8eZi3EjWt8xgdPGNxnwMZ5HhJW+4CwWH5qHamtwSRBj/unHSqwGYNBLFOIxwsj
nXCYkuBzrgqPthPjbSwssA0HS15tWeMCBwNO5zuyAlNjH6NeLvwqAE0CvffGuDitiyMMqButlawQ
nhjaJJ/UH5YlHV+6oUEZzwtS6yjmPQ+uA+4+LD+GeygC8ZVJUneY6iFpypCfn0tmkyS17FG9ThXm
dCJi5MB+/Z1/BbcGtGZkWx/fd60PN169iILIA+F2xNmpbQuvuEHXOb7nYAtIBv/gYWrqFhiSPOLf
rrg2ydZFhS5xpL6Awt4PcXxc6yXL7lnGjJ+mFTHPRrerAaGN3c1htsDuWwztIv1KbDK5P2e27akV
a58AmNlokDVFjlHDh4JKRxud3KYSFTNM8lMUj8TVkRqFCBR/IfSL4C/dgnSMl/sUc7F2kTJwEUX5
ZOaTad1zyZgrmmSfXzR2h1PYha3UeY4DWIg7iIIG4sOeNP0FA9OkVOfWmKiCN/A76sLTLmL+qGHh
lj+7JaNAZ5EqWI0uKv+Wvdm4uHr6i1NKdr+7JuXTUn4IqPrPHyceQOXFbmXPErXTRjYWFm4b3/T4
5n0eN7hOCqEnDX7Vt7Ii9r+FYSgOXaSx6Z9Ad+V5S+7VA1x2DOpU/UvhTvOSS+0GET594xMQE1M7
qv1/TpaPbSfK8Vt72P85+mPfye2NlSGjW7XdewWNnXNvNXlUvJGAasBMcoD2kS3Mrc2ODqoiv+KZ
vAHqBzbEYGW8wyGGRs4HidmzF4F2t6b7ltV94kfSyXGVUVdWJzjIwEdqvsh1nCkRiQ7r4CSZCxQQ
1lfsQVbk8PBx+flwNqDcGYyStVqNhrnUZoKH7Z3tScB12ClGkISsvCaQH2DbYzeEDd49/pEHixHD
EpPeQkGO1pa9zEQFhbtvMo1JqQEEhAebaGZSujxno9A64UDFRxQB/MQ0uDIevzBrpXhK/96Sh65d
SOOpdXJXQqHGWhcCFyuGC9h0atlX05Wcav/O4lFsCTiD+brB/2uRcg9yXOUb93wj3BS1d4/rroeH
tCe1+BuvYm8ukHbr+vLID24guMM5mx+lkHTS7w6sUDHZdmHJQocGr/EtCin1/scThCEG6CBhHwi1
f2QE356eWOhePASJmTJdmPSmclQ4TbqjkdQEmylwJ4vtjvk+SqsUjHIdxEehLYCLqTmAwBgK4cfR
pXe1rO/jK8J0rPr4sogI0nNH6O7buV0ppWKfEq5YyoJV3DmQcvmHezkIzXj5CQAhI6sMkGxwEPmk
W2JgxrNuoF9iw/4b1juVKpIZrMU2lQnsd90eEk2fbON2f4BkznlbWHqx8G6L0zAq9uB2KztKXwJQ
3UQ2CxtlxATnFIESmR+QrpSRtN99QJQTc6Oib02Wl4P4Z1INWqYqiKwjgFXK8fVEU7BSjtx4uWmF
a4qljRnBZh9/rul5I/jS9XtCmGt9E+eWPCLmKFmeFz8sB/0jvlgkBKEexvmXakQr4gAcazN3FQcE
kNo+HaKU/ofKeBaw3F0w3CQBQTrXdQb2iTyaqJfYyJMJlmyFQsS8KxjuntdcIr7IvEgAMDMMi69G
h4bDKBq3k4ZSPw81wBcZNQnhk6UrxmaStqbgV1QP9oJo2Icg5wAUXDrQlFGEBVXNPE+CdMe8Z55C
5eQ36od8Ks3iT8sGN1nY0mAQm5MJaeOx3/CuciZA7lj7//7Z7AkuffDR9Q63FGirYPVlpSPFYx3c
F5r4ro7Fd9AQiqJ+4jHXrGetphagYX1GOwlr4JXiSn71wlK1xdZYtnNg/2hHugejaI4OyjUgQqjF
MwKSnqBw0iZVdpfTpDvD94wKlTkha7+4b4yfQ6pwQEZuxJZ4+mzrma1s2XYnH7iYLC1l/17qNgVU
WvlCjxQcar8QfbRCqY7XbluZYrresCxcDwO2aChZSGR/aCJeZ7Urzn2dviGD2/Wi/3DgMXtr7Rfk
OUcZpwfE5ocKXFHWAjo6eSA/S7ICbN3NoNfZYysoGYWQ7JUffdibPS6ssdmWFEF4eEQj/mQQ5JhH
x/VqxJxFYVmrVm/Lu28HvqbeAVwYdVmlJLUMoGlPeHiT4UAOGs+ZJN1k72XhE3nWwsTS6x2sHyOw
Z2b2HdiFY71pNPP6r9U++bEokB5FIfp8Q3Xc7lz9WuEdBUITwpNxa06ngDg7E1wpSzaTBroLWNj3
mCInIs1fswXpdsDwyWYd2zI8soNGdStndKp+ehwd/VDKxOdLoaiP1GQr5CW+8ASdtgFWjJ6mgPCc
pHVV0pjtpE/8MzF1sK0JW9u6lJ9XXA2i6ggHiKI23sxxQdJXFdGyPhSLlo+tJd+4HYr5JRWbGqu5
H7BJLR4nnPQrcTrQn2YagXEB84PQTLb2ZcGdBgWB25u5zS6aWIlbC3Y2Y0E7uJ/7QI5oJkcQDlte
ZKyI1tJAIr4P9Iw68OUW3IAlqSWtvHcrNNbCLCUK/DZkXQ7j6a//1SXto1/FWSQwp93cu572Oy7l
vRKHQfU3Mpv6RTmxA7ioxqtf6m4xUJ9VSZdbSuyTglQW9WXSNg6YbWYyY5jebzofWjAeb9akI4o7
XMODvZ3QshLG0QQuyJ1zZvLuhmHrkDIQSkKac6yc/nHryFz02Vpy/7N4uBcqNI6w3Mb6+zh9cOBv
JDRcrsrPa3g/Qi6IwE7OM2Ql+ZpsNOI1XpiB6wMYwCSJf8/mS8dGXdaJu+7VHR8NAOd8f4iV4sWa
HjRwZxxe2Bdd44/dgWR7qhM7XRLHYGZy7WSG+oH9P2i7i2K+8UL64gPDPZQzZK9hC/4PFU9LPuue
Os6UR+6zoo2evWEiCuV/mytL+m+1rsaNaoCSS0ICobGEPO7oZPB0Fs0RrDQ33fm54uCdBx6oNTEH
aKtanPWtpNowKmUSmBO3q+Mc2djnf6dgMYu0ZDPe70f1NSqym1VU2qeEqtlEMrCtS6NaEfwfEemy
/R8ntmxt6i0EJ0Qfslfre1NYVJCk206S/VqlrC/e24/QD2zNT4EjCeoR1ZpHVqzmLgKvQHqOliMG
Spnjcir6H0ASkVpPCNdeX33KfnCxbC1OBIiWBTWK8te8mtNoe13Y/nHP91kctyzAY+flVB1LnwYl
SwxrqtiQMSnpX3JIiOIXypV/F7E5ydXdQMXprtQdbNUL7BSeH2ckY5xnIPxO/FR7hzyClCXWCj2+
Q2TIwKnAkggfNGeuLyIXacCPdx04LQZKFEvs384H7v6knfbCYBl4aEUSe2U2YHIfJ8QPputCdaY9
I1wQIZGckroqAkljF2Z/DK+BBLa8unfr6iHYL6xjNjvpRz4sCxCjFgK0lEAIWULq46EMpcKTRfhI
Zugiw/QdKTyVhVqs/X0lOORIzJBMUsbNzzHfP8zAynJmzX+fKw767NBtJ1cFS6f7E26yho4hxLG9
3TirteopAqMI4XbyJoIZSLV1C2EN+CT5Iv8sZGCZW1ZneF+pTHOa3tHlq5NdfFzimzJu9jE6u0lL
8v7GQ05HMVun1V0kkYkE4x3Yyk5UZPI6MFEe2StoOriIV04iw2i8ohwcH98onlRDn5nTg0kEJM2N
9NCaYkww4P8mlzMixy58YkNqT2CgrhaSrq5yTgu0UEbHi+U4ltMCLyYXIGNcDfYCZWfRkS8VWY0B
DbH/hpA5LZJLKatazxtTYWu8WZ8TeZXqq/hnuUH3/D6dcHcLc6iFVSgxA8i/tcdv/yTM2PDv7yIi
O64/HtmpDDsh4fs2krpiM9A/CyoVWtNk03Bs3enyi4+rLIX+fEkQ7S7//GrTrXyTLSeorQtMynbX
IF5udIqsK/vWnaJSTUrxWuOwfhrz7q0WHvpDvMTc3PiqBmhF78H+j4Lh5BSiUqf+5Qc963Dm/uyu
rMAk9lg+lgexlI4oQRT5JXqS3Y45quMDTMMLtnCXB8BlZSpEHMJQK0uqTRZJzX/X6IhjGR6oEhOF
FesBDy2a/n7jwXYtUQt2CZFlJ5h/1a5Xl/F1J3+6jhdyeFgQd2ZN2B0ZZJyBGtqkpjZN2nM+Mvey
d77Sm8faV6s+VG5ecBC5Ke2f8RNy7wuLq5WedBkYSB9TT5LeM+GQZimX8ori4bQ1adrrQu1I5AHY
zFH65WQ3s1rVaU0nO2FMVNPN6u8TbtgM78D6rR56GPiJ9lQYfBZSqdqd0nLPo4530lwzeNdyO8Kf
6viU7xBnd8VN6n0k6oNHgR1JWq9JueIjDqAa7GRgO331EMftavnCuRM6Jf9dnYT6RqpYQvtc0MYR
Mm2YGpYt2evvzhSWq1UOJIUUU01X9o4eIw9yAzwImUBpV3htMg9nhRu8EA3o9FnVvbIP0AUe5ZVQ
Z1NegFty5sk/mO0hGBVElMem1QzSOXOGcGRlMZTpgaSRJ5a8wBlZYTCYUhPdfry+nTfZ+D2sfYDS
Ytxx1izWwDiNyYqXXYnLnsnfAFyM5VG4ECzriRz9CWdpziXo7X7gA/fNEUFwgLcn17IUrdTAtBVV
qRpH36OhPMbQLfBCAyelG/ZxV60UDSzw7IAu0Rso102/aIKbItz9/XGYEJVju1x39KaaC9AxX7P/
ZPAWoxGYmiNfWQpjLQEOQLt9KHqv5cgC6Z8SLll9+u7vGHspcrKuHuA/7zYficzgyGHqbgCUAJYr
Eyz56OOIKBEGRFXh8MAerosuIy1r8FMiKxv/kpQ0zZlana/+fq8ZFXcPel7SU4RSAdcIT5lAN37U
+BpRM7G7DPO3bMPgks7OAIHNrJSllL8Ruo5bPsoubGZfRSHiw5NVivfWWSlkOhOELxvQj4/Rw0zQ
QL/5Ukjg3N7JlSy0kgPkgvL8MSvjaxOyRkgCLqgyrAWzQq88jIB5Jmcyb6Ya5V/nsUigMgY/xb0F
nneM0Qxb1hdkMOnXFAzyRtGoOlJfqLs4+/ZmbptFCtGFT5b6J4Q5cJikRU/Qr1keROLpaTWb0UK0
V5Qq0WFHenGybYCS5XbqT+dHuPSYQi2DKsM9dBU1VOkPaz+x+qnaBXNbp2qtDM7MJuw=
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y-=^��l�yN�����(D�p�B��uY2��H����s�X����� /`��:Q������bs��(��s�$-�i|��jS�d������ Ү�)��s�(Ȧh��N���Y-5_tݝ
�Z��_�Y��U����yn}����ٍ����GGS��~�1Et-����^�o�Vb۞��{w���R�п6����VH�(����^�'$��NՁ4��`���<5�C�q�s��$����[?�J���M����Q�J�|��24�g����Eǖ��T_Y`�O�/��6���ə��?�)�9�&>@�I*v�}kF�D"E��� �h5A��rh��P8x��5��-��j�]�͍�K��ґ�߶���i��a��U��s��������x=��3d3��G=�R��NYΨi��B��
�i�m���'����z��Ы[�Zt��q��̄���lds�	ėʃ�뵟��J'��K���Gjq��R�eq��bB�����/�G�p�ң1����G��ߌ��lWt�FJ�����K�խ�b����!�g��u�>��i�~p�L�"y���������x�KD짰��V��u{��,k��s��?g�Y� ���韹G���e��x�~B�2gd����[�gɛCO����O��f�?y���֎[G	h���%O��/|SN��*n#2!h��J��>��f>�<�&�!ct���K�7d5���S�&���]O>�{ޞ��k���+/ b�Ɗ�n��Y2�t���;������Hz\�E���3���NPn;,.�[�f�J}��R��e������_�a{).� C����(�\}�7hFZ�X=b8ao���mڗɺԹI
2Xʴb(��k�k��ˆ����E���vI''`�T�8(���E�U�v��A���k/=º��7d��S����Ψ\�*��_�D���Mm�L����b���B�Z�j�.��?���Kd���!=�c�GOX�${H�.&Vj�'e���w0�n����)w�H���f.�c��eU�o�K[���څDr�V�����4#�ɢ�����A��M5��'�p%q�mM���6^�ZF%�v��[����[�)�����P�nr9<9�J�0�
�ۤ��:�z����˴^l���R�j*Sp+2��O���Y��(��۵�^��[������kᅿ�<���?EX�L3ڐg��hVn_<x5kZ����]�$�粩����,c��]�rڪDj
�K5�����L�)B�<~�p�����l���(��"ˉ񧅱��Iٗ/�g�*����Z��+ݺ#�VG����RT ����u�_���� ����K��5qƭȣo<iLA�P�=9uZP#�뒿�|�j�6@~+@.�	����$�z�\{���yC���z���x|+Z�О��-������+�x�z\��h+��J�b�7��U�x�b1�q9Oڠ�#Iͷ��N�T��U{k�?"Q��a9�0�zc�-�wb�6|V^����-����O{ب#�M�4p��%6P�k���%�=��&��9� �H����u :h^���	z�!�v�9�x9,�����#盳,��=���Q�π���W�J�:��c��(��gTwN�X�6�6H^@��H헣��	�t�i1:�j-*e��o���QK� pLA�=��^(ji�M��v;a�e���/Jg�iaXA�/��jׯ���Y��E�b�=���;)�$�Ab<���X��8�t�L���N�{X��L�S���T�9����̀pg��.bbwRY��I?��hK��ï�Kh��#8W�ލPm�e�).��|�s�#�b��d-��~�R�G��ish����a��N�8�w!������i�d�9f|IH�果�v���|U֥����}��R�pA�� ������S~��=@f'$;U���'��m��@$�U�d�u�B���`Q��}�G�({�Jy�YC��!C2m���Xa �Ƀ�i8��:qn��}�y"�d4�F����%���r����)���eWj� �.��N�a��n�S�ۛ́>��*��̙2�S����wv]D2�䰄dUk���r��͵PK6��ȏ=�e��:�n4�=�=/�o
��9'F�d�������8��� ԶA�D��w]GHԎ�t��U����]��#�
�(5g@A_�_����8�YӰn0uN�1�g��O3�CC�MK��l��GY���Tm����q�0T��Pw��"B1� ��Ѿ����HG+ҤL�\�T�k��P���r�/L<��gOko�����+��*h�z�1��J�_�D�L�$����6k5�=K捴�� �u@W��E*!��lP_�>\���`��������u�.da�J(5x�Y@�N:��_/��)�ld��4Y�s?.�����;2�W$���æ+�=Ekݐ�+cש2�=�������zކ��d9B����C�U��RK{�Pm��T��,X,~���Orc
y�?�˯F����w���X�B��`(���\9WC#�3kO�#�Q�xP���,���[������I�T����tzX���r#���,&�����;�#B@��C�ܻ~�q<F�=��]ψ��w��IV�T����)���s���&`�ɇ�^ީ6�۳>G�Xn7y£��"z�^k���M��	'�c]�Y�U%�w�IZ��Mk	�����Q�4e�{�o��KpR�]�pvq~�]HG�X���i��0zH�:G�@)��Eې�[W���P+4Z��(�t`|��Os���U��z;{?Ԅ�w��UL�rTD��c<�C������(+�A���",��sc�����3��8�w$zr��UI�=��^�	w��p.{��ԖN#�4Y+�~���D��pDB�Pp wJ�q�N�0�3)����
s��I@sl�Z����>�ۯ-���������«�CB��o���y��7ja�S��s�G1����#(4Q2�5Z�{��
r�8�;L��}=����J��T��/� ��H�+�����1�*fzԯ�~�x�O��\H�\e�\ @g�p��rn�TS�h�S
IȮu��T��1�d�-� �)���D,���iIYn�7ˬy�[�yQ��X�����n�Se\ؾ~�^C]��d3��W݂�W	�́_'����0��^Ū3((^�I&ϼ����i�>�,3W�u�6�'ڬ�>���ΐ��Y*'2vW�P>$2j�J�f��re�x}6>��HZ�5=P)�Ղ0"q�4����G T$�W�f1j n���Zy��XM��9 =;k�g�!Ĥ:�#x�m�����A"��4�T�9��mN|�+L�����
Vx���Iû� f~����/�*:�{�)>�ƃ����3�MB� l���V-�6̡3�j��I}�Ո���1�'�)aŲ��'f~�VM��H}�_U�4���!��iIG߉�a�[�?�Y�~��K�8??���5C�$�r[�e �9���i�Cͮ��gh���F�ڮa d�9�ؗ�Y�� �����"l5ͱq�����w>�ו16f�Ͻ\@���
Z��
�z�R��I�΂�Y��#-�x��/6>���`<x���!'�3/Ytq5̦��h
^�	t��o��g���u!H�Hb7�r���w+���@�#���P>��+��S�TFѝ����ӨVg��N�6qL�,E�BE��4���ܶ�+�&he�Q�m�"?Z����.FƵܭI���+.#7�f-���1�/&��� ��9rH���������sU�u�� ��Bȡ0n;��R`��%���UDAi�A�V
�R�����	U�u���+�����#��+s���b�j)y��t�d�C�R�a��p�/²����&��r
jX��邐������v���Y�����f��Pq|�T�\�(קy\�֪���zU֜�O�j�]�]V�x@+A�ETr��b�D�x>��x`ʷ�[�V�_�k����(e[��;�Y� k7|c �:_�3��<Q2��� ��e�fB(O�l�)5%�ÑͧSqH=�R�@�˻蕑�+�o�>[������+���;'�Vr���>��0�^҅�0`�����L�E}dj,�?�	����gr�cS�6�/��%�_�kL�[_��v�Y�H�T�!3�pNH
6�����F�����G�}�55�.;����~3JJ��#�0���܂��6�AvNu���:�y�Z,���J�7C{�31�R0��C�)���z��U�k�~(G���a"�L� �.������d���3J�w�mg�K�>A��Q��X�o��j�awJqn�:����ޠw:�	>˱���� lu�G���M��S�g �Gw�>4@�:t��D�[ܘP�MÄDf�i��M&V�XWz:0:��2����]H���47�݆/��P���{i����N�Y2l?��ʥ�w��GV�^�c��ߴpy�]��$; �h Oi�ۨZ"�z6/�K�כ�\��H$$$Z�E�ƞX �5��8�f��!�zz��LoǓ ����2$�[�_�����!�׃���\{�w�:a���/�.b�]���-���H�UxK�d��#
���6�~�.L\)�ǥS�Fv� �Ęy���D5C����?ܰI�3��M�n�*M��|��{��)&Y%�-�~�%�����F$�5w�J%��}�!�nI�������#(��h*ċ\:r\��lc�g�֚���ch]o4����巗FԪp������
Z	�W�o�oKl�|�l�[W�<�G�^`���PP�0��/ ����=b��n��ڐ_4DP5d\Ѥw��	_�8
v{�4>3=Tpg�Ţ>L�(;K�9��ԙĔ�B:��������|�Z�	�;,�u+���8�\ˆaj�X�g�2�.�c)�Pn�L΂5����AO�l}��4�m>*�h�w�P���Τ*@%��c����C�
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rlFR5WYmegv1ILOmBDbE6SM79OheJHO4xErGOEffhyAPWMSvX/QYnvZ8lAelWraAzBwPbzKh47dO
sCXwIpOTLYqrtGd5c0yRLsfW2niAXB/Zz9xeQNpuUcZiXs5LPjUmWF4UJ8jNhFoTvuI92Qg3O9AR
cNlrHZUIvd71tpwzNVJfn/EBII7tBXQip3R9Nv9RvFjFZsnh3lY77A57gAABnqzVMTppN37EVfff
g/KWZI5/Yvt7n+0Dsz2lwDzY7XOSUp/hdAFJJruKRbgdkROw4/vf8uiEQE5W40wVmWBxEXlL/Q/6
rkjk/46RKrqf/UEVH4EIPuWIgNZUbYNvoh+nDA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12848)
`protect data_block
lzRuHhdRCh+/9fna8NcKgif4Q2+kvcfiaQotVjoyJa9IgZ0U8+dV7yPeIQTR7zeGt+dJ4IysgHSE
1TYcyhSTIeEBxsWOD2/VjGA5PdYMOaSjOaDGfNLV81We1uiKRPUp3XGNNvnErtaAahyya27CC3LR
QgYwLZmzm58BJS61ZzamVyI+pMtCzVYgKkIJJcrpyd3FnTpFg7caig4sihHIGRA0M96APSohiAEY
p7lsG0/SXgjheK3AaxvUIrIDsZxsxj4vhOe1rVNdYniMhJB3yGYBVW2QaNBAYUZMvuXM1qvfykfP
LxZgGygoty3AZaYJG0VDWLHzBsIfWYBrjrNJrIHoUW9OSx8Hf+xynChCrk4CXPdcSxp475m1v8bK
0xc8MPjLJel56YLxzIf/x0BH95UKNglURkU+BGk191Znl7iI5wI2yVfAxlNHlS7r8ZBafjO1l6ev
NkuwwIRR36UZdetCK84xnme02Za4XXltSOI+x9rDVuOpdTUYibEncHLqIkRvion4siuebYxYkHu8
ituvYGRpqImWACXbfd/3lsKpwdfo4ZQFD42arxoislt/fSkB4RJ11ni6Ic+2ynIAjwJCH1gPXzib
4cpmAKkvrsmhrnummKMzzmke/L2/+0MKhmSNi01eQVyanea82KkZN/i+CljmELcijA5um5R/CZfw
v4IK2WmnAwXotExhs7YCpsW8nEXOu+GnnFn088e92mZoX9dmOs07cFiaa3lrxPUMuADEUZyG4Ve8
Diq0CYuouLJ4fMYRMsLHWiCs6WJAA/BE3Xxt0NotKhjjreoEKJSw0nXM8pdZaxMoMp+lSTEbs75n
TejQKqPvBFE1RDI1UMOuBceLejTP1iUZuy1Ip7mffUKRTlyGZnHsEh9orTYZitc1stWz2y4mWXEh
J+L4xwT+krWHQuD6nTDkJu4rn9CHxUA2KVTV4YjELYbGt+vhxwWzCkww0iykxd3Wg15+5vKIIFPe
yo0hRk0syFBjaBdaF1RUG0t38zVJE2+bp1cYROMZbI7hQTGouieiIdWV6k5OI4AfrBKdFBZF4D5T
IuQdP22xcvJNvJs1yGZ/GJm1ubd+pBscynVpMsXUTSHYWFr6/XxiCpz0ZaL0SHvPt6YbqbFe16hZ
FChWOcChC/84lVYNDCRnGwTVIu/sPIrNPhAMugEdR93ZysorWnBA/1g8OQZji68fvPef5J9CFMhP
AXrvhwIy5O8Jge4WTyS5ICKeEMwnwV7wLpVBCDS3GbeTKLBIVJAfolnj6cRuKhPa+s7cwwnWocsj
BnaEbvRFPnYsPq42HhtHwwnvgRbpDNvqUNhPotZOQQrVN1QmLYMYOBM6zOjk/cy9iZpiE0Dv+h9M
ddVyDqNqGNUXO1UFea7d4HrCnye0FZgxhzveY72/R2AUrOsBVcBWZyA8f3XC1mLIelUNqCWYKofE
l6pqsjh1u1Ngpb0YYSCR52sj3c0Z+WC8MxPK7csHheCT5KalWonXzCXE5PIKoaJQ1repcxSLV5hj
0M1qphhsO7gza4B6Ao5rvnBphJ64Yl7LOom6MHhNKWzEoQgaXE+PaSrmLd46fzo6MNEYf7BWZ74M
4TO2LF7Tebvnmhj1B1ki+++XA8QprReLD9lTZ83fCL2HX1THEeChs8i7P+7EWdIWAsuxNQ+9iA2m
SNRD1cKvWUmQ9nK66dgVTTkEEsqE7Nwy4geBTBjheid/lEtdQb4BomJii2CkJkqjAAljp+U40kJU
2fbek3Vg0b7DQetXY4MLFs5lmWGEZ7FwkFmVYVGocOwFWW6coaQ+gqpw287e0YqQKVUTaSKrV2r+
T5+sYa28vKXOVww7sneycrgO7H6ro3YlVi9rRZ7FzfwN5jC8FPVF2sEEZPAOAzp9pk9dqtLAIwXU
zi2wk0ObDBYkMPjcrI9L5mWQKgJ9lBry3oMOfXoBE1/W8+UWcrwFUM55BPX/fXvGtFk9g9Lv8bDw
WTF9mNtapRqQ2VoF5jMEQrrNeXzxvCQ7seRw3h0v8G45N8UjVCEal6dfWPLrOsv5mxB3ZrLuoivW
e4Ud+LTpaRdO/ctWiTpWFglKcd3sPO4fW9aZ8LB72lbVRJ+kGmaVPjG9fnwQCHN0BM87NfkDpsTn
2y4gWcFOIFfnsPODj5jUQ7rdw5oEgdsXXDBbMzoRJJXzREeH4veP7Aas2z+69o19HZDxgjx6q8K3
FJxohOO9GXQlkSTY6n4YXMtARL8yOwB1oPcL4JIOZvn8mygiIGR/mICCX4SKucwVjMJqX88YEr+7
3pFHBRTaxbm4CT99S/R8fWwDSHgxoOWQ9fvH2mUbt+xBR8sN8MzMNwp7mdaajQipp2fitvW8B4GI
K6UqxnMEuSkndoWAOeM5u0dMlFejYmSoIPVwFDVF/BzXqHwqZpbfIzaK0K6VGRJ0+76QjaHdkv+j
vlhc4kaA5EUncyLJkBzQ6bejSM2JU3Fz7XEMR430FsO+nlVL2RvCVksZAtqoCPjmpya09RIslPB0
FaP7bGKFKvNg3epKXdc9QECD0ik1AbGUlNpe7gcj5hkedXp7XY7Kfh4yl8jIjMRkMVj4jGuY7Zlv
hW0e/1KR0S5/Fl3FyTjWT5dKbgGpq62ab2+Ak9tJCandbLq9SNPb+jDCCD4/dqPbkaLjj2b+NtiB
3zdnPB89UxwVDaWBf8KUbt46kAIEL3qNtEBO6SYxkn4lTMZ5Of6JJQ7vK1sfUIFwUQvTthrbNOax
8RXiPYcqiZG1TN7APcdBvHL4hVYcLpyCaDHxGkUNvitQ7/hwcBV9j0/J0EOoyukkrGt5B3aNGeUs
+2XuZW3tnAGqr3XOfUkJLB4EBE6fiALDxjp9NyuudhWyOsX3rokqDsnbQ8w8gZ3608IZdPnpebaR
tkWYrgFdVeBFKE7tW4mHbhQwxbxD6nzphZd+5fsstEPHuZ2yd/+fk3pMJwwnNpXQ8/m9F9poR/c3
E8Kl6eaO8lpbh08lYGFCX4q3PLSQW7v6fAri0G5SAyb6QmE0jiyiLBw6cwVwouQXjpT2Y3HOFq6f
62dYDeSRF4AIdzR69CinX+5AVfttak5jOU0KratpW8ytMZ72+skT+LNiQSYNpc0avNln+QvyDxA+
6tTDJ2IMDf9wGMI99RTqVreYkH55MSbKKmsh0Omtugah2yINeJoqmgdbxNJM3iXsZOik4OU0iSF6
rX1jGLwsprq/tcG9FOw/0NbPrd8EZm2jBiZW9eLxWO05cxROa16l0BTZVkuuIdf2Qb+Yb+KU3gKY
qqKGjTBbIh2J5Z2k8+Cpw6IEaZh7zSPoLsI3W4oJ/PzpK3hIpWrhf1dCUhRcuczI10wRt101zrbI
H1pF7tVrpRNa72KKWI3rGrma6BWAQrO249g3EBSrTvUNleK2JMSNZvbeUsw2ZB5SZDYJzMNvZ/Gq
7+9FDj4lEuG/WZKfRoLsXZjQPIOW9a33/2jLfsoB2d0qJv1vgYBRy785fbH9Wn8F/p7Ugey/vZlg
omwDih9NRM6joGujmjf5C7wshbCai8bc9xl0m/Wup9y3cZ6BnGHz2OHgkijebcFWw19F8cK5gar1
IaX8E4EIEv/3RfqcE8q650lqldabzc1p+GfFvcIJr814FkocZV7xSMCt24jpXyngr23qYNQAOEFs
zKr2nSbevgXe6oRjVAnUh0nATJ/igq/MISGQSLZrEEJ6onW3UbylRepq3CHe2jxVbU75NZ8Oh3yV
nfWLkAiQFIBqzjSzOrigGb8kyLBcRWKvS/hKiEdMa3Ud8IfueJOFh+4QYm8Et++0LeJ5pnxEM0eP
KxCq5ilrUbbv7RE2waKZEgBOqQJbEyv1GFsPLvRvsIHpkwBQIXt7bXkZSGlEQbh0fS4dKA0niEDi
IohBfUIlDdHz9yWfQge7Yo3FXbdFc+D/tTVPjKn2YBLQIMs8A70YUikjGj3vpjyg6UGj0vU5qyKW
L4mX1S/TB9D+/eIOxujp6uHVO5hK1oR5LYl50h2XtpfHIZW9xkZqcwpoVE7gNacHlHUTtbWRnNDm
ilLqOUHLFTcf0oC0gmQUZreH/FAa/Hg0j0TEPaD8EkPLvh4KWQegTyvGN7ahJ12s6wXGdq63pQ3J
aU7nIYRaMdcWzjs/5T3QP+Nv+e3hhmHqu6SienfBwm8lURw2sK/LK+IiJqjuQKFG5UsVmhbVmbSV
OUpdD6YaQoXhzjkT0YK6F7ueJzoLOQE/QvzHOpPGYisG+XWIdacobvmSnYwbiWkHtPmB9E+8qZLN
eYnu0x6YRFgsKZ6tBSVwTe7477eO2F4yFOTkVmkwRo+JNMMHzqTAAnndeCTnhsppwjitXcQR4cz0
5AKvzmkWWNFqx+dRN2q5bjChB3mqu4vz6odBYmqqFe6849QvyE12++ewWQTahRP4ULqovtFnofWZ
FMhr1hr+ceiepwdKnJYXCKgO5P80Y/R4CzjA38J7j8AeLNrBmtcZSlxZm16xI59B3CuH4YOyTDmq
ho5LMSPVNFCmm2gJX0eO1k6JLPkjF8VpYZ91hxIXGmIhioxoT2ic52//lvMevxwk/UyWZDYJuT3a
+ZZ/TtCZiqAIZC4+MJWNlBDBZlGK9YI+GFhu+kvJOS2LRc4EWOabbwjl7REb/fbo5u19IwJPQT2n
oW0O/xFEOzOLexeWIKQpwHNDXArX7cToEUX2y4hmD9iRe9G0kcUbp2kN8w4/zfHzxxBSJbqLrez5
aZH27lcM28CZqEG1PZ/aWZpSKs6P0Nz8A+vjpPuaS6P6ru3XSbweCQOa346V5IukdsSGaVgFxNVs
KqS08AQAWU8LBOuLFPlR4nRNR50COAJHRt1+c8yxDlFjQdIvCjVG5Wh4WcIPuOjkD9WsUHO4NZ+5
YzSXdCXhFk34K1xbLMRwg3077QFS5iBfd099OixiG3P++ieZ+zeKwxNG5e7kdxJtPKdQI/ieMeb3
pieGbcKp+NDJnJPmOQxgGMIt+Du1bQ8UPThlTyVV+qKkEAqCx8/wPh773dGXIFwq3eOMl0YIlJLl
pbFzThTfj3w8JqJ781zv0tDu2jWlBZti95wK5yznP5DZ0bsVIin4CSvdhAeccu7EXic6cHgbIrK0
PblGmFtpRtWyPEabiAfQxuKt48dpg2sPzb/SryrKAnjMlso8Z/glsMqTnxJDJ1Ohjq5p6TdXWNPi
6LzlE4bWUJzQRc/P9tWd6BCxkYm8e1eyd27RsZ7VEU8F3jJ1CrFshc3JBEUOkh3u+LRqkte1GRB3
/ovkZypNam5X90VZAtJYCJy6hl0qlONty0GWV0rVdGiI9dmt9u/pOQGx64AYrjQ7Un1cXH6X8G6l
OfH0EqCLSpnPr9yjUgLOGkZBoE53pziKslqKkR95H79XDZOFYHj5N9qRVXw+AImDyEX3BwYlsnzD
/7hdeZf5fFfBsCX405JRLfaE38VfF7o/by2lNKfXIt7mp/szvc7EY/eJnreBZ+bzWurN9QT8j/U1
30pi9lVofEKKdn9HlJ8sEWt7pias4kvSznPwKrWWHPowiY1V7po51gSRYZCCWNwmFWuJKhamTJoJ
TyPKk5jWp0nsUkXA7zmzL/O7/OqvUOl/VHIML2lsIxofd0TSwcZK2QhCWpCFnFjZm8vmsKm50cTl
8SiFqwlXcW8jVAR4Le3bF9GNk86ES34+sSHJkp5DVOHYOY83dZUn4Vuv2zFTqH696nszssAw4iWO
3ERoebvx5KAwcjIeavfm8MSyJJILgr8wAQt16dBha2iR3mupnnFysn5B3/bsEHLGAb5YTenAecYG
ybRuieMNBf1pihuIWUMJ92zr/8I60Alc7m93wXV2Vw9Pfqjxwx+UQ3Cb1JZL42GZaCDQIGu2xuLR
CrJt3aavff9cHuSs9kgiLRFmteUZeMt1SLNT98S6JM4dKa+vvdyouN/b3r214a06dqBEWPLLt0Zs
kORqpBvyrnkKo8ciek6q9/R6THw7/6SZmd7mDsdiF3lTrfBOGfgvkUO30aEjvSZzeRT6PcgZAAQK
ysp+6DWQth5QbbYwhjNk/A90NZ7yuBQxD77kJIHrpTIOEUBquA12NABvSQ5P1LngHm0SFyhrtSos
OHITI4J+IgEML6B87WZEiuCM9s17ZcH421RLAF1MBRAHe+5GB+seucf3ayh3T4CGNoTpLpLcSY2O
33jGzvqjJHsIAlR35ByRaHEVuop4u13bP0TId9rhScAsTgSKfkZHYPfbaeqqulJhUUIkvkae4MYZ
jWE6OnOe7gFdZnqgo3nDt4BXzAT3f8DZQv6KEqup/cdhVC5NszTwYgN3Kf41ZZkZw/3HN1dbFqEl
CwRt//R14215FnvpRpNprhS2yVjIdRMGByKDbHu3LiC19O9UUciqBV3IxFTWxwkfV5E+8WoeNoh8
NxGbtjZug8ne6c95zrNxQ5RDAhKoLMvGsEpORCY8dq62Tcc2S+uE5BLhfvzdGerFokBfnzfdozmG
HUJZNunZu4m13QclYpTjMq2U9yIhCCUhPc6pFRAAWoglTUK8gTeg5qxOlxSe9LCQB6k8rwsTstGx
WkMyYSU042OoYFfTOB0A4DjcpEiq3RdT9oMgxtsfiuRnKKUbHXujSKlKrO0J9ccZq7H6kEM2+UiU
koDrUiqNjNNOQr9yUixeqj3AoxoHSWHY3cJDINRZ6bKoO7m8oLFlX6o7NoF4WB4eehJMtXzwpjGp
k3L90yW40Dz9xB9zhoSwB3OC/GQOsvYRNrApQnPdzt+yh2iLnWY6q+b09T0QKEbWubFjD5vKglFM
WdZlINL3FAiPIn1dQDSx9hJ2Zp8JjgHtzm8ucJSUSEaf2MuLHMnKvC9kkzMO67SM6tSp5HR1m4h2
DmLcUn01zUkY8TZ9DmG5NsbFAY1cm8F/l2eLA1+sf8lb3GGVqqWGno3KFkANi9zBky1h21TLKFJT
bC/va8bTtShzk22gAOyIBXTPMPiGr+fuPjgkuWAPYOpX84YdihTNXM+LAW1ziJGhu0IvKlGYATxI
0YVvrdmsDsAF/3iKc4xUC4u84+Ecrb13pN/kvyU5LDjTgm12r8gh6cC4tO5aXeBwD0FAOfIOcu/J
73kF+oGrKzJmcNwoxHfFSk19lr+tWx0931pzQZUM97o5+lDppGEgkh9jT58QmJ/S/wqSG0SfcIHt
yu3S8E+vV6El7/qBPAKvzAtpljoEN58AiHvCOctYD8oI9tneznow6jdCUCoO8MIpIs0jp+vauLic
aT/3bSdBToIyyDnV+feSfYEEjVOXXqVJtuINfaZqR9HvUuesXTQZIA6LgZuVTkVGoTzdUwcN7Fy5
t3dW/ykgWX0XZrDaCOVOs3AUTbc+yjCrQZa1I6rtps5xaT+lxw4ocCTOdHGwC/pd/H3OFidO+qn3
h5abYFARgOwLzT/PajLIY8/eaOfSp7b7E11imTYxZdtkkUWRc0RD7swbKs7+fGPfU3pMBzSgZLKt
goAHS2jWe9nbtjhzY030A2SUYUXLIbfDeaPMZjgC5nJzU7wq0Ho6N9CPHoHnhMxCnRO0KOV9Y450
y4tnvSDFjnkyE+TaEwbSjj+2RiW8ER++P4AZZwGVWeM1RTrQUpnAPHV4eedm9i0kYRLh4qGVD/eT
8GQfIJvzaatfOWoHNY7jBfpgMh5z51bBivMAK19XOnvfeo7SKbwxW7Rtw1VnhwcRfvHU0xNAJ0Fv
8K8qT6VXm1jjdY2WRinWExLF0eAebFuDKyBLPzkmc8oql0Kdxud7Lz5dpJ2o3FEY+thr9m0Uxc3x
RD0gYewrWfmUSqBTvzBmBOsmnDzvH0Nob2OdHej2xRakv+Uzx4PYw26N4gzpj/4fYT9Mw2WT5F/4
XstZiuMGWR2VN+3iZbqF2MYfYEuFfbXXSVWSIu6vheLPmms6SFM0xK+GZFZqWWtqjfZpMo5NpvL9
l6wyR5ShRtpidfxH9dxS2j1ewT1mPiv5NQ7r3CjFrr37b91Ap0PE8zfYSqhT3pRhtHo14RzR1P2y
QQfwxjSoh7stozOo6B9Jy+Pj3NM7YcldAm9BRhTe9wg/Vc0ZZqVZW5veplECE2y/rjMI5ur8fXhl
px6OzBNBCJU7P5e98mcscrhDe4X4im+anDpXl70t6mWcD9x8Pfv3leqRFiFdXYSs+1/gjNNyZU/H
WcUNU+WOpjYw1O4hkiali/RCH2k5YppRL/MKJoDAtJ3kQW75q5lyb0S0p1+nMvgrE4zrNRva59xA
AQNO7k3rrqAzs55AjQxc20Wz21Nvhtyd6qDnh0p8szlNgo7LZldo85h/CBTLNBzgC3DQG5syogDm
hoyfDBmuTqFpLf2BiA0yzyUTlqYv7zO+ptVmyTgdsY4Tv0sRltaM87UQWAe53gaTqElKvQIcMoN/
kOFywWM9IQWP9aomOlLqHhGCM9/efd/qA/lMdecPrDSWTaKkg8t7FfSq/DLS2PW+ctvWnmb5SOCW
OxZR1+IKNjhgwR2P6xbywNLy7FghE/UrRm3/oqStxdrFIKh0lyzmAlpQ436DBL7zULDNROsiOkVK
omO8iJ3oXz0PpeM0pCL7tcsW99BADOmM68Or4FkcrzliJZHIqnVv6kpIsLwUsLq2zP5spAQsc7/1
h+LrLpe7TOWw0HjoHgXX0B4B/YQJ5HtluzkLS/339Hk3ZzZxM3T6WDks0ZW81m48c9xxekXFRlXW
AYK+sjuNKr0WSuludYKOY0HVTZNSaKQjhNRVI05zt2HdzWrXKlPTf8KTlvgnsedQhZcd3NC48o2d
u3Tom6qVhxsHkNZL8zN2JWlRjU1mxGxfWYAsnjCWl6CH/NP6tywsKIICy7F+P2jRPe1Wb0IJMRU6
54jE64z4ximCms6Sb8IUN5RMHGhd3Ss/hMhqivBaChrPsK58f3DK0nRjNVe9C30pXX3zCm+p4ZOZ
2UAEG+NosN3h3OJ/rCHwo191lanAFLbyUFNf2Zm7vT21wYJ18WXQPMyUdvdpAJuiMhLE82FA0naZ
4jrSUVtEyFD2ORbCdwvIL9yfv9yArL+5k+gODpiOMnSK8yWhIHC2YjJbfUtTnHykSrSjcuGNlWd2
OovCk0zaI1Xqx9yk+OjrK8mKETm5knMTLSmhtgmiPH5JouByuK2qbkl2wiXY13SxXyM59DUugHzH
5+D/IEBoE3IuyqLwPUKzR9y+ZyRq/pIGtSyzheb+E8I5Fn6qptbbr9nNjk6aVOMRZRkPP181aL0P
/bBZCFZJmuf+F64VlnA71QBrBzj9jdIMbhHUtJ3b78CgOBWhK0TKWR7Brs9P0js5zWfOq1a5YHqY
kztdf/N5D0mY6Jity9JZNnetdPdoaI0k72u2sZzv9gR05ZXjSBQROQK6sj79Vq7eJVc5BUPS1Vt1
YU3kE+t4NuVldmM5SvnsG3mK1ywQ6JiIBctODT1X9vgYqMWl/X2sHkBjglwSXkYOPTNsYTHsB0AL
ZV/wFbb2ISLlFlCIq4vC3SNYD79t5rKkTiFI6MjSKOnijHaFRlIj6At/Lbh3ZQA6SiPr6urd4qSS
dWRGOXHZs97JIrYa+qY97WPSA5jDIOh5vKyKHxzW/rWBoGJ1SeSXi7YDco/x4Y41oObHPzXPHu8b
21Swr4NSVuu1wKgKQxfislvDJWRVzr6w3TbeSgzlRY2Yejg0PrDUhThNsd6Fh5P8UCB4+d37bKvr
Xmqh6yu5y278HfSgfANspUagp9v7DILY1mv9mA+xnyYmuNlLg4FlsD4mmvCDGkhaJLDSkQvwSFce
LQJaQCEluitNg87sXLQsvCjCiIOjKhXHqpxJrJATUwh0tXjw9l89hgCluzo+3m6shSDbKL6Xii3/
YoP4Z+ZkVX4XfI4IlwYXz6PeqIxmTIUZvOX0j3CHgISm0wsSkGAO1iv4BMCBJR2S1g4FApDbyx+6
xMUqYCfntS3HavZwmiS5GAyljSU+CyniUvBc2lkXu0XMv57gNUpthwi5zWQRsLzS1ija9dAsy4bQ
6iBosT6kv51g07IUVulCxdNHrzJZ8DeVda51ORjWZr2MlJaMAln2qKM4e3VSUERTRzzBi96CXkxy
RI9sONGA2fA6SPqHqtehIvhOAsmN3b1PQiOA2C5PKCB59ADeCcsD5zoxMKzL0twS1Fpwr5xgIozg
MQ/TKUQqTUcv3iDNzbUfT+iVTIIrkqe4yhh3Kvmr6TYCuk9biFT91Ldr9d+tliq73slR7i1sI1dL
QadpCIrIcGSeXdkdNvqafzGX8gfT8dD2diIIjC5sMELA9z7KreWcvjH8vZL9vEuuHnR8ftOJ8SXJ
UGc+NzG7TjMlT2xysYoVuyRuYNL41weTn0xER03IK2GYPKMTjDtmm6xZ48ts8KxpYhLo/BxJKFb/
l05lXZOm9iPgVkdhrtdzoZm/AH8okRYW/O2oE0QEMXaDNlTxmItK5WglnIxGN+EU1O62GJJ83teh
ZYFRi/8nLHsLqM3YdghQ5QC603XKuyBy3AmeGnRKzq9Ba+iT5m8AlKq1HddxIbzXNCqaos7xNljl
REgOPBk6aAwq8/37HEs9h/qbDvmRClq0rmoZPHahHD19PdzRdR9GDyZ9hEcOAodn1YwiFcNe3U1N
Gyn1NByLUA4+LpMdpGzrWpLdia4IIDv3B37r30UMv0t4YoAQdiAAPTcaxIxIvx7GxDVrg41e2p6a
BNoFLq5I916Z53QCLngr+Emz7nxz0aeDWDJzquq0+vXkm96afgcNHyMQuVg7oeWUa2fZTTtzkt2k
Y8HgYzEbeL0VBaqc/LKGOZjq/JkW6rdcq1Om4SkA8ssRMaQ13OlOP6wnOu1u+aSZ9cKDc4rjRBBd
O5k/9YN9KMU9TFy2JKNz2mRClLaV3Lr6Z3Qw4+TFV5OKR4pKjU9hQaJ4R9vQr95LKxA0xi2Efz9t
Erwbmv2l5XvG3pwsdercU8DDDGT87+y3ePbHFUzfy44qCLja5wWsa0McDV/FRXdOiGKNy6zy/Peo
bylramqYPYqkThD/eQwzsH72SL65dkZJ/6W65cqitIlTEiZdu54c5O3Uza/5ZF9VPxBhzFp0H5Rr
0+74PtHfGFTN40KYqiuQ0NAIT/Zc+1RZ3uPj091uiqqmE3xLKWdpCQ6d37nVoojjlOPWlr7mhrP3
7C/JUS4ENEOmWqIPjAUaTg1vnwaPFDcJ7LQWVMg9oJiTmvxNvHGXc+0J8p11VUQ8v6qSNkVWh+Ag
1OP0hv8ll0WrnekqL0tzGjxQM1FxM3npqhHGJkbAeNYG2hjrwHn6Xa2v+utgo7IS0WWSn0lVbZSo
yBOQt8l1J33ruIp7nBBqTHqfIhIHK4ivbx1BTFcp+N+qX34YWXvQ0IK/RGQFxS/a829TMP4phNks
Dm2zpJvESTy2acT5dhRHgkMiGPDPHe56qQjgDoVu6JFsKAn08zJrps1zXj/HTNm/5D0gi4VU1/hD
/tO/4URCqp4WZdsfgjEEBbHkQgfOW7DcWz5didi9rH+gvtxUaucbEybk6VNY8+V+HBiPe8I7oB1C
i4mB6ioQL2DW1oZ4Kpp4Dk/xpniByCgYUBNaSGfwc2sN2/67x4EsGVshO3OW3vYDnOCJAprW1vgo
LgzIioPDBc1W5FyollK60tJUd3gwr7DIuP6wRnx8XgkX7lX6HrM9kzD/l2Q1U4Yk5pgUFB76ETk8
FXTeOh3+rIXdMNPcni5wq6exvu1HKpWSxeCBl1p71ZNyMTlyFx6xwwK9A+0Jtq1AOt3HBqZvPSJI
3iJXZZkrrcJ7TBDNZSwVb2bH9tVFNaTukj/gQrf5AsGP/3zPq31BPhvOQ8lKEfl5Avd61JayOGx2
CGRPUQzx9WpE5UHhW9DGcVXvkvqv9ANsZIuYng7Hh+6dYxxd7zprq2/FGWB/Qbew6nu/JUrt7XwU
9VCqedlMMmU2MsFAIPRbphpKIWbi4pYreEuH+Tngc7DMzzdaNmARayy8JjOtwKqTLYpAJ/SVINhV
gzwbBOq8lutsVVscSc1EMIVYRYuZNdPPPiuOuC6iOXhyQnk8UZp3NADt9ezFxJuiojTpz6bB0JLS
gvemHigiXv/OoyrwrJRcaFQ3FqKLoI3LUoZvVLCD/3Tm8X3+EtA1LMADv+TsMXTiS+2UWR1jP4pa
lRCjM7BgsNhKWBGoVDxnMmlpuw7wMZFtLrr5bOveym046ftyzsOZz+s3b4CT5ghDQUcGUnX6K/+e
s4GtbMbj/VcF/lTo9HC4ccoFPz2+72KnEm68TiEm9ofoX3d8x0qiLj7HQYyxDH+hNW2aj4ylRX/S
PkQKvYq+hUbzk1qt5NeQW0o8eG00Ojp+LHi6uaivlI+AJQJ0qZjEosuKA9SF8WZFvZFgJPJUokR+
P4DvCKFsFlGBgZQE5j+r76AjUaMpZyhHJdDFyy8fFJ7P4s2Gp5xyfyOEmrNpXdBfyMhxZNXodkdv
bI5HBfnEIT8T41Ueb+25reeF2wA/3Kg//Ur5vLXdDosEbGrZ6wW8wOfEuoVAt6JLzl41c7t6fuD3
YoCuS6yqY990JCqEwMjKJfZEi9GSS3nWlUDzn/Nu9vF+YeCfiJ7TciWfo1a6yK2BSJCJK4WDtlsa
CSiqO6VYS47TLm8cXh3xwFosTbDZiohvElS9pnj+rTWXUlYCJVFkPYuBzSwFDrrpxlZTsjsfciFi
Oo1NvnTEuntsgkQkYXvMs1xjSCL88ZYhhALh3v4nwVwCq1axjB3huO/d6aR1uhbI4HXwgyB/Aa9P
GqKGtMngyuiU6CPyjv6OuFvaaYHiS8iKDCNUASu8HIU9sgeXvTuTcryEM7k46KZVjo9FofgYmur4
eJctqqziASiGTNBqW/+Zga76zgy+gVS7NkpLPpYsZaQ90mvAq3TMK0MuRvZ6HT4rsXURMO6Jk4MQ
6uEpDwYbBwGBhQcF0/BYGt8sQHcZS1/yp9OpbbnYHhulLXoaYGDRQuRINCc9KgvwFwRiKTTy/O9i
dw2gzgWt2eJwP1B2fugV4HFnWgcR+nXhAKQPOe5UeL8ISaFxcBs+0aWoMJe88dtDcAZtum/u79KW
xvWVLqIZoFQ3OwPtKNvqQfT9vrodqIJRSl24/ncMctZ+xGcB4rTRDsHO/gQsAwUWsQo3X9hJP45L
Lna9yQByAZdnv8LFoJvTq1p9brYNAC7DY0wmgi6SwJs0gzJizblyrEp9A1SlOShil1RhTUryZmz6
NsJp5QEsCrJQxHFKMU/BXENzuHGOP4QRFeia2XxY1r/47eJWoU4IPFwQYrYDLg/2f3/sCAmcnAnu
Uicpn9qkex3pvdnQ68ruxyhynLE8XGzrucdktMjhjm0vPFpy0NKRNWsZ035TJecXd3XHQewvZJOw
v4WU2sik3E+pxlzw4AVIWD63wopuEcxd+jVWA/bGlhUKzmChHM20bIEwdEbjOX4gZ1ExnxWcvgU0
iOSTqo/C/p2uIDjUln70fIpsIfI5UXwrY0d9XQESc6DV3uXLPQEu8VeGy73UCoRFFkjCBLOratcv
VL3THaAol92u9s1oPDOc+3YVnAyXLCh+hIKFbQ/3Pd6r7CnCgsFO3J/f8yqRfKqaPhDk3iGCXhnx
iOZ0tM+wbyNQy82xLKv/0jA5XMqB0QyqlytEgmMjUhR2+xY+1pjd6Ke0qsGGegABQPwCQ4wtXs/v
Jnh552AaRHLxSxAa2QxPMTjuYA0eC8PZwTQHd13vltikbCIkeYLfiXUY6+EdpETfZlvG5237WUUv
q4BvZ72vTX8MVlc7RMMGNIUK+6/Yt4hong1FYnyvEyexeUCvbzu0h8cGJKMp/WS9SuJVaG7wNldn
iYjX4qzHODYJ3idBbldWH23A+/Ffm93pKL+YwCEFKTgMpul5RT9939Z8AnARaciMbr9eKlQ7gFLl
9f6zngXkgqmsWaJzjmAvMPU9shoSyXtD1GB0E/K+6PoWWgYmgCNHyutwH4ssGYgQc1fbxcvHSfj4
SnP7S4raYmDgZA578SzZnlk/MUOodkBkMC4UCxsTU4tv1yjb9589iBcPzCXi2MtspK8E+yym0TAO
IXlSIorEamauuRVR9zHdSoLs7TB8iDPI58B+88WMaD+jI7IW4yEkN2OtkPInSs0tVhWh1PEF3C8v
cPhhc1iHHMvsOl3syD8uqsR6FNo8j5rhBJ63wwxZ1qfOuLM+QjdwzwVgGPDPptGuOmYzGKBm4V6p
xAMu23VYYLR+0XgoGt1v+1ItLKqJX7bh2o9oe7c7CjPD/yovB3QdRH6xrWAJBQ+tMTUKRN1McYRE
Gzqd1HHszKWJj11Tfmo2HoM1/8lyJzXH1L5Lj7JZ59mRkUu9dW6me+9eLHcAmZtxC1vSESU6OlkF
k5dupmDzf+NEriHjr9cy+EJYLwpqACxLm/Ai9HGYQDfy/X8XjpWZzBGQ6ZxuYpsnZbRfumbdqUih
JUPqg31Ui4AQKTStBGA3MCM6SvL0b5fU4H8GHuqwsAGqdp1ZrMCykB4RL4DUMIrheoLle1Pt3Fdo
aKG5o24DhuqYow/43u6+5BbI4Rgt40Xj4QnihZrQwVchFklH9VGKNQE4R8q18TXJUS3AJq6rrFYB
PyJJsmbvo55SX63F5Agz8/qlLh4VWZPuruuFP/LW9beB4aYvnszuEAhV/+SD6KuFhhixKx3OkhlL
ZU/pvjpZ8U4zyX2GU3YtptOWk2rVBhmoA2nphFriE6WhxyKbioBcdbGp89gmJAW/es9w6+mgmNPE
4z4FrTrvZMMbJglGGQlde/41o3in9Y2zwRx1D6Ez/AFrwl//o1OrLQd4byq26P3+z+CA1XhPCxyR
mrrqxViB+WEq1cMRAsWyC0HwuqEyoLv+Ew/CArrm3CL+7WccpiN2p5+a9etfP4buo6N2hshjgfiA
/wgM+7yx7inqgnAg3F5/oKW3d3sUqoI4nZdm9C+T0JLf9tw+3SdaA1RA9Yu0EtjY09WdAA9HNtbs
LwGcDRwfZkgEgjwt9ab6MdoJLmBV/6tXvVik/JYF/k4owFROuv1AbspFQPR7l74gTKjNcqJFnovR
IWcm38Ds4AZlWXNqZevWFMV//6jGBFlmHNJT6g0XKMHb2tXpl1+bMljj1qz8xhAgTVfrIoy5bzZF
5JtSx1dUxogmpmcfmfbDF/EooWwNGxugm/ys0A7GZDL7h6/I1yXLRWqaKG9h/rzmBDXXRP19B1JL
nxsOkb+XWiu6BvH0j1jr7c70tRlfLE3rfvuiQeG5C017rqqOS64MSuNF/V6nacmOYjSbKcJOtaLy
empvFQvkvUqa8UK1dH949jvd9CXraGAyagDcV49LAcWewuwqSzKX+CbpJjrlsLJn+W2/LRHYiXZV
+Ou2xT83y+dfuVf3mC9JgWWTJUKLk+UPr+9HpWrXPMzkZprUSZWEPcG/zpHg1V7jgLt/f9HbObRB
vpkwBFhUxgxyarwrTaHQUf8i/d4/VUnl0GfgkayF9yWt7soCIINjlomDGK9j0luL2u3hlYSGHAwt
3BuFp9tfkUlQnqzFPQAmVK5K0jDEbu9RQPisSyOWAg+zzCyahELOZBtFsqw6Y7IzCdrjoXwCZ5vL
S5OpCWDSbSw7Jq+OtAd+ZjC+hHA9NqB/aegyk+vW5IwYav1vizmTkooLyYG3rF6lYdvpGbqGTFAn
66smJt2s4kdNGYFWKvOna4iF9yMoIWDEUtJ1gKHIosjjX+eqahpRxUpra0kEv1akqk+wR9yqp/3L
g/PorCem+FdQFMnS+BqMweDADHD8LBumjBrOt/JtwEv1cgCbBXYFbSkwPwx6z5Ujm3jE+5kk5MAl
IZBiklrN48yCkt2BTXaMpTIrAbgLiX3p3NRPIsXeH5Y4iq16z+plIy6j1M+W33R15kRytzlg06Su
tnNBNcHt5k5WkrxOJ+Fc1n8HNwr1C+MCQsOiw3AXPCArFZVNN/UiBDPg1ork4z89+0fT4iOyVFhQ
2avFxyCwnVwg7taoYlTcf//yFsWqhXnEp2+3YXVwsep09k6ScrT2NESTs+2vElIhzC0KvG7ajFhX
QM0Kei/RTD8cB+p6j5CIBKri6LIbOsxS0K6b4slTur1WSSHukdEvcD/mknOEXEamhyeDxYsWp9C1
4YzEKqUWDtbrQendLcl/ysD2RqxnOrugSUAg/mngoY1aXAXqY+VyKrGIFYK+p5nwZAbLCNx0IBNT
OdUT7OWFzLOc6ocZlh7+R3sWAD53rDFNaPPp4H/3lqKKa8RM7JONN4QV6ZwqBdUbXQb4m8/KDWLQ
Q24BRpgdqdjKlJBkQaXtBxydllHar8QIwe+QhqUPFVdWITtxwcNcT4WsDhM//D/jQx0ajoyHSerP
DfzZCgfFyGcuYL5AfhjHybBPiGOq71NvpVVnBDzf/WaWGddBcWWHLYdDl3VA9xLNq6ghh9K0N7Z1
L4baMAKo7DMTCmWCOBpiAym0Qf3tueZaUCeiBkrG94pw6XaBWpmcFsyvgkt1GEpg45K/q+FURqch
/+ZAKJaguW2RaD4OtsxEaBvV0GM2ff/6ItcRm9ylJjgwTC0yY0ldqWOU8fGxPV1oQDx813vU+S6i
f4BSF5mpk5Ik/0LRKaYIbTIW2Q3jSnhuv+Rn0BQOYM3W+udUreR3GjSwCFS0XIBqVaBnCGcprcEO
uCE21OGqL6Xd6My8vy1LEvMJTJULiyyI6Bz8JT3IXrW+M5BX5DfYLJCoWjbucLUeGxyqxJLZ5Cnb
UXpgPEbxQ0TNefGuhx1mjeGh1J7PHLMQOechVTJprJgIQvGjagzhXtjbODfjgOlpX7QVUzvKQQE7
EZWJXGeplSxA5Fbbv0M5iOtS41DpxoumHKYnJidzt2pALQfAUkjJgouh8FjkD7R+TPRUT33pWRsd
0P+MFVYwUM0yY6XxCu5M/6n06euB9WOP7+Oa6bYAtvkthmSxX2nI3Gr+JzoRl8IqKTF2/Ujq4dnU
TspRfU6NCj6AgJkrWlW80vrpTe+5F41WD+ifgPi4Bl8V0KmN8qUafkFGsuCk+YpkCJRNjMzsK0oV
XSpxUGQbZaTCO/3TZd+90M1Hc5ggbtbQo/KP2sxWhjns5McgdHEcEdorMavtIvD/PWs0TT6tTxdn
Cj+JBk1BJYMtu+gINsokOj6uhlECrr9s6TKhzTwHF9GXufPH+374fb8ICRqsOfs9nTANPzOyWIhw
77XjjX8U5ZI9iwGFd1/1/xeDt5oslqg=
`protect end_protected

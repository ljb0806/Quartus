-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XzU7iTzUJwChQgtHG5qm5N9/DF3FY42r/5fQJmQ7iRCVQiN1HJ6XBSSXg8KjXYDa4sT6mU8X2oSp
Iw4sIyRnX6pLoQv6sTfiRsbJiRWLBOEBzvghdw6EFz90w+e6+bjYHWXxy1Ip+7GUfooWO2/9HRAp
6QS6JbMkPNoxX5ObyVhLS4umkNc7rXugzFgFj2RLLCvPXfabQ+o3r7PMXcQWZYghW+U7SrX0ry0V
8ubIWQKU9OBbuPKh1+CL+05OHU2Y/DzVDDIMb4E4Qw5Hk/kMZ6CnhOMzMtx8JQnJSFHpQy07WLKb
c7rG7xJCqY2QNDzqaYmD+cM9g8k1xbBjfd2f1A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25136)
`protect data_block
DnzLw0k7ZQwqR+igQIzB6laNINwp/3HH3833Q0LvnSsExHdSY3HjET8NzfzBz8EMWNZeab8h41uu
YVp62DtI76jn26UVSEptQnEYT9g608GaNdSNYO3w5yV4Zoor563yMF7cyIdoAOCIxG4AKPD+gOhv
1u+oN3NqPFlODbjyfcS2UOUk4APeeHx2vEpNXk+0Pge+LcmaU969YfpKZbN8NP5uGrSV0UeawKRs
LMS3O1BXhaHVqfBoxlC7tUWO8WfC/hasJhS2ZtdFaRkeDk7inr+lC0YBAJr/PNH65n0TT5qgXsv8
8or2A5NcBRRFig1DQd23l7oyuQ4PeQTZDraCuHZDcCaG1EMHRHtLjaYJAyccZdfLHaTYCJcCNDIF
tpzgT8IEY5JsXd6oxlwYstDPElRqVcOZmNabTlZNaKx8QSIyTYFjW9u1jg7uQp68y0RgrOSn6Mid
Rqp7Sou/UxFiHg5LHjDu8Xfqkd82aGloQM705seePiqCVZkLBbN3pcHJvF84S9v06z4YIBSe/q6E
/fcUuRXlKcdoGreZuRNcenyU8BIXdljgbkY80UArDdfjBgWBDHwfHiCwlj9k6g7tzjLtUDeBDX76
/zEqSUpzej7SjGmTbf8mfxqRYtYz7hIc3z9fJfimRRrSdQ/6WRWofP2BIR7/au+ZDM1jwrhAPq3K
b/EtNBliEURgsDs/yNDsx3vkIMGxzXholFaTURduParCF3fhETNrMszyouS9RRAYg7MV+xpzn7iT
nMuhdnZVGWJ/GH1RtsHVQRosaby7aEPbHVkkyRKnNz78QNZNn+LmrwvoDeG6NT77AESDOuSE49Yp
PLnlb+QEF43bpBEWFNPuvHg9wEIPJdZkPRIUOyw3wTS7b2qG7mQU5znitBmXcbGZWru+e+xssBxX
vDCCyCgaf2ybhPD9fbF8kiB47eEN9p/DggU7uy1zjs+zhJsgVCXXI1dYbuNSYdjPazKjXEoc2XXs
AxffEKoJX7E8T0BqvzA61sJqVdlGDuqS9A+NcuiQSxNNk+qfYo6Gdk7X0iMC0C9/MSS3Gx+2N5me
5vNupNvR+KoR4mMBRfBSTYyUmfKx3OMdLAMmRidHWTH6LRx8ht507gHS8EUCabj+9Ichvt7Az2EH
Z6BHzWiBBuTUkxSaqDsW5F7zN2eBOMqyOM6+6hSlELeKAjs0qsXs2rT6dQxlfLFhfWe0VJpz+Wc+
11NqhG0BuyeOFmjPiSJFjtBuqNXnYZxuA7vuqYb5WS+0qVBUnWCZC+BhMuWV7R1YaoXmFc2Z282J
pteD0P4MkwvOE1Df2fMkicuuMHXdQUyfgf0sF3kyJJZrmzM05voaAPoKDnox8vCQXI/xSVxyixq+
G8cENEss4bh/tN4/zbJFm4/Hr8K+INa9bWguqrOwzEuYInjjXjPp7Yvl8+lkEuu67OeVjeF3mf8t
KzMWrtCgNsYfUgbnMlQFTP2l3qIxiypf/JeMgiZE2nfmv2SpD/n6FcCPy+TM9ZKG/J/2Qyg6/nXa
fgOVh1wZj5zqZznK0GD7l5JfyhJ4dOEj6fkn6NfownpvSataaXqakprEAqvRj3aZFxfHiREpaVKn
ubuz2rB/msiyHZ1wkY0uI07daTE/emO+lOFhK1+dFbhrRr01GQt31q+EeTI3prp4syx7As+cdVrk
tbFp3lmevTguQvwo9EWv+mw20NVFfZSSE9PS89Ltg52glXwry4MBV1S2F2oICNBT+PCYfzxRG/VH
+kWdM9GEat2Os0C36OsGmg/Cyz8N7Ot1bMUTPel/YNJUvDWlzxcGtHcvnjUc1IT9Mb7RvXEXYCc1
C8DfpxFyFcJWqjDKDW1d6F59K2+Je3eMHsgZB1TiPkRc5C3HnrUp7jP2I7tfheG8yBAZrQiMitiC
DSXg/sQ2Bxat6Iwl9FgdMxFB/rHGxfCABjqdot56z71cy5kGdrYu+zcTuyBTW7Uq4pPXcOnzMeLl
EMMQcoFl/kFmVi7pqmFHo4TX+HbhmJ5txrF1sfeXUIr4q/LApAszpM6FMd+z2qwdJFMX5qC4TjdC
SoMMKfk1nqpTENF9e16GXmInd+WNWvpFn4NvJRtsL/Q7WiQLZ2EUhgV894gqAYg/+8FXH8hpw+B6
qvKDnPeQHUQmTfS4SrbM8FsCVA2ehYu8Nc/zGUm0IGkAfLYBzA8OPKxmQXcBrLkTQqtxRgFQW52X
B595Vw7bMepOIg+bJvl8ioFK8PlXnfSqVGDzi/rIEPq1O4XiuOBbkO3/4yc+/ecNkcnpk5YABxvL
Ieo5KsQW1K09/yGNRzmgR7CEXK2t0Qd7S3jbYS/EBgFQD70joFq78lkjZZLTX1coMrfL0sd5t4cy
TO21sMpKdyfLhThjokS/+a/HIRutqkc1aymRUTFW3OkJ/MIc+NeuVFypBiawUxkJFFl8mV46Llx6
pkVgOCtE4H0rXa/xS4j+8n73ZCVqpI3AG1Bduh9hQP0erO+s8XB6i05PxyGdsc5OweManpZNMx3a
KlLBB47+zBmRIcw7UP10j7kYkZe6iLNf6fn6vWEkpgFGjAeE+ToMRCUveXhAckthIlXhOtzGhKcq
lFwMjpYXWI99tlXRgMR/pyewk4mi+GwUwp52Jlc4RmI9dCnjiLuqYpbwVDteUqadfKE6ARtpw6Sv
lkrqb+RXaLtB020eP8MtIiIlgsz9WUOJbvfQv3v4EIrjdk42kMj1joqWsbpBN41LZR9gTkz1scjX
ScqKyVETeX1751cIlG88se4gnFYnyimNDtRLOjFCI4R0tej+BPGNDL1VNlf9h+rJc+bl3keJQEFL
dHwHrvcVjyDuSqpmU5fZWJhcVOP1rUNJ/ci6xjTHOyYqaumaw+DBHi6Oh1Gs3cYOQr9oPQcFu4tz
0WnmlyCk/mf5q8ZLGg4DEeprSMHj5GmiJyo7tkMCjPlqLvdPZEITAkSmetaN8lVoo1jfereickQU
0dk7s+bN+xWhIUG0WhMhjiSL4ArbLlYszvCCSycfZDgmtYHwCE+Uqjb0GQhFpW7YWav34AH7vQbM
VYajeOpK9LyCV3xHjBES5mKsFBFlHX6o8iOWt52AULUmg4TTTa2TOGJTKckG7U7KWs+fAYst8BlF
nMuXDP/pwSaUSS7AZMX/0xTkypCJxuNY6eU+u3f3atKklFU2F1hDE9/yIm+lKnnaYVXKtYDgYvMR
AXteQrlTodk74e3kbBEwYWmvBaXmkD4FLGyd85yt3Rs944M/C95o6mTjWW5U9C6RhJNn8nADyC3x
3z3ReUNW7PBhaXnqi297DyjqkYoVP+r1p28i7GBU8OpgLmBLYO2tVWkQnMB+ynvIL/UqaygcbD1R
yXmUWDdKuzVxJZtMNiTEUM/DIX6EpQuIUmvyYzei1b74ZC4U/WoSmrogo2QRdV/uptq2c0ZbzfnV
ylOSn22oHW3hqYXwBrIrwNOggDM+Fc5kGF5RpUnKwHiHQYM/DPIvVneOf65hCp/Chu5m8n+gciO4
p3KT0cgNvtI2H0g8lncToYfWz9s7f4yrLUxn3kLIRURp00ff0T6HUfUIHIw0MR2rvTK7MaPo1Kdv
WI3rlF2akE2cf6Gfhz4dNqOCQmDhVhqvP6x3Fr7fmWQ3XI0euY3jVPSVXjrybbRF2A3ixxDzlKpJ
O0NqABNPND+xBWPYTp6ki6iQy/dZ0O8taiEgo5dDEzdc0zDONbTRCZMR9nFWX6simI7iMFa3OHYE
RHilvGwoYDqPEifcH55Qrs4uU6dcG0GwzJ9Zce06TSLQvZbPAXn6YvfdlzLcX2aHBHCYi6vkwXDM
0IdYDHu+dkEdKJJXaGYb3BCJ3gTWmj9/lqMf+QsN8s7Zi3Hd69d5ECXrw0pijKzJiiqiDDntBq/9
meWCeY2TUuHvy9K6l5lvHDrUrzNfK+VuhIHXZdjh88/bPIUN8PudR0MTFgSj1srshIYM6oOoJxPv
3SjkaZyM1pyHLqGJXosNjUq55TMxN1+cPWBXlj912qUA/bfjjMRjHu1Kc2QiW5HajnXRJDRXWHLR
uKTy0+vAus2oqPeQYIf6bSzDbf8uAOvPnVslQPcw4OzB5RmKrmRGr7Gt1paKSBqVytpyshV3MjFc
WVSO0Ww/T8s8/JEqLLYCKgT2ZAG+nnrspH3KFYrcvuVoc3UqhzREE0Ju7BA6MLImILKgv3BVeFAF
ElNFlsZdOe/98HbWlnj/aVhQmIhAR0FkilaJVp6GIcsquLmrwqOE9BdgST19Fo2YmJ11XJWakg4G
xubigPa27bhY0UN/OOOZdOs5yYPcB2wxHmswHz+CogZe1eQB0jW8x226xdC9FvZ6G4/TkzkOSsoc
ETHVTilk5nEo5jy+cZMlDO5JYJ3Mij79ocbCuZ4kMEQkMMHQWeGOxV6Gr5eZgPZBZrMfRBMDg7Zt
sGy0NOAdjSrw39PEk170xFmBr11E5/GUzFJiSxcG78KXjuuS/Iy/1SwQXBcP1wBEyQZ16X7oSvYT
eCOATSiEPq0av16WdFqkWrVGzYAn8Z/p8PdxYYBWwSxxPtwIb9MOK8f6INv4px6KLarRBLgTJ1NN
MciIk4T2UQhhGFcWTQCyBKDNX2q2lvxb3E/52yK49Mp0d2mlJ7cx1Rcw8+Vtwr6yurB8RWS514HM
96UxFg3PRav0iOxOR9sRY2XXWK34Q6tseJh4sNlG5rteMUnoOfC3snqDoAqg4uy4Sf2ZR8WNbEX2
d9iOnP4jYUTwQ3IOiNhe2AdcNJ4eeNk9cL5yk1G30Yrf+Gcc07cGCBn2XxHhiaRBqDFxURgqrJjm
gBTKpSJ15ZMgoYyKcUMMbVcogwprtl8s/X1xH0tBatSv79K7P5iDVxkxIc+UgWsf97gZp4aqsDjI
9l8hJonp0SEjA15c7Vh3VrBkKKWwAVEkp3YVwuklga4Vs/IdIW4v9fPWn40LJdf1T5SqYdM9hZSg
EM0dpXy4HM8SCeb1cyLfvL/d2P+f5gu3yBM3WIPpfljwfpL0xuWpe9MtKY8tWIdsTMb7yvH3IFHg
/Zu7FOLi0wBttjqdkxb3MSsqxzA++/CmStj21fZPLC90W7bI6H6wOZ27f2UVsNvGPBRn8Ihn5VtZ
zTK5FmCZSPoYi+AN4bdarHWKbtLA31QK8k3ulQhPpw1ZtLThwZQIUVQdmxLYU6Jc41lxlMF5p3ki
En7uQjOgo1GsFJZ+O5WWbrSUmq262FCzZHT9JIEby+vb2/BZ+FemDh9Ww5jwvF/Nmuq6PP+/HMDD
UcHDy6i6DNMfzDKeCVSL+YroJ0UbP3dZ+axc05xvM3qiqdhRyEzR2snVAAFFuIFQLCp60Pt4DONs
3mawfGil8aM34J2pUVEaqEafKcm73+J/rQgHCMc7Csd+2ynbLh0XF8zpkYvXkXhd1asb32azrFcE
ZiDyPj3/3io1Bmk0XEzGtsW8/GILnx5msDSdheZfyLa+L+AUUY4lgc97Wh95Kr85oAaD6UUX9vzX
mx2beRKsot3UUjySIoBvZQLhlk5eUXEDhBRo4IBQe5HwYbvCBNj25dkINfskN9eWdWFuE2XYpmpd
xC83e6FAXaVGMQWXN9VyrYbPHuD6a9WM2MD4t9yzlcLwfx+EKB3Xgp9QeXO5wdSloo9pGZfRIlfz
ykW1Fh4f1XX9oBLGJShbTXMgZeSK36UKQqqfDHKeN3eU135PiyYrbZey4mY2zB7W08Q4gEDfCFjR
MJ7ESJuMl5oNZdoKI/rFtUoXE/+frs7Y6Jp7MjZJXfjBa1i4bXsE08py80L1boiJ98AU1ygtefXt
88vhF3/t5mruW/PR2u0MSvSBsBdQe3D/F6cX5xMR6WbDx4YADWuczyo7asRUY0O+JAOIXvIwbpMN
b/ftsXkgEbs75qlbfumosyIsS7hOoVjPXEw4SZG+VbzwDfXxJu8+/QosH7yIXMPH1lH8Pdt83VSf
cYb9BoA61oUXyWfwG3zbbUbCLMVll5P15bVjvZuMrv0TQJG2tnC+Qt9tsKYtrj0wTUgojLOFptcO
hm5C2azUTfe/hYMNLdiy6dnM0JRrgILQYhOYgp5XVb7YrXzog6+osV9Bq5n9fSP1Ao3h1Y9UQ9ZH
CIlhRKL0g4wxgxeBA47Hn++7+bPI4kyDnTGwC6j7kRzUYvmvLDEQuRef7dlOwws4t9J+IebnWTEs
sS8L8ZZu+7dkH55pigyV6epD1v5B/gmxuLCIAXv3o2WJ6u7oknAIo4X7VUjWSkttyRulaKdU0SJC
AcVe7//ghQxjnt8LYaBN4jG6K7IbS8VCHa4PpO1RU0EnFrw9TC+tKA6yDW/qm9gw7lb5PkJ3/rng
OWnj4OAxElKy/DN5TxZkorHf4iaIR0iJ8AMKBlEvOV+f0Elitwd20g2+p885+YHF40L2bPF+mZL5
xa8wtaXwjjsjEu3iXz45ENG8qXBW2XzK26DP0mqjQh8UcPDQ1n+CCqdxYpGeC8W3z++NMtKgOqUQ
yeRWTla4zzCTjmmrTm7Jv4zbu3cWENAOvovtinU2cqn71g3Okby1TDVYmhDUz/EXcvKlDDskSpwl
Bb8n7tGEo05yUHJfg5vGcggLwUiaEo7QeGWrbugQ320TOp0Lx/8AVjedHOpE6VzZHyRBQ6jg+54f
qfcc+PN1bZeGMncKLLZS2nbVF7CCr22hWIW0kOeoagxJ/g3TvlreLIZGLHzcJkYuUyK9cT7tB1la
aUOAJlRyJZ4V/tU0wymnjeP2LpkbbAnrqh+XNwcEtQ0NXMp/s8ZTio/XzO4DQ7MH0fxEbdDRpVNq
XmYXWGRa7gcieCh2Z4SINxaq7aBasesbj0yo5ECVCqKmvvMtftjvUPrTUBntLH28bWrU2mP7Zi0o
wYRFNFz0M73Mp5qm9idLzp71jK9fuWE1vd3xrUFfMLLkwEJvpAVBe2bf6TX0y84LQSPxckHB8PH6
eEBNbCH2LVQj7K4bh6ihUepvH1RTpEOStWTfh/CgdmwLvwmceOzPbfasBPHmGemlfnoRaNKRPt6z
SpmusRzo1IA7s/cUyghwFtb55OKMfYeavkJ6yVeQxG2BClbzeV0CmORogk5iAkrbzirP/9y9gN6Z
3G5zB8kH0k+cRhYbduWXpNJe05HR8H3WtiQtDbLa4YyS4XqUEVLS7hFnW91ECqmkSJTnIUoM+oo4
ZH5H33wenip7Kl3Rv4HHQ6UdhZQr6imsfvv4FxH1fttvFe3SfxAu6x/N0v5yWjMljpW6leEWx1ea
C2b4nyg4pEVzSo/ANpjDrxsQ/ZN6qnxtCyageftDAqjJ4LJX0Rvnw9a+rnulm9wAJw2NPVWAZdmk
AoBCBu73YQuM0kXlrjRfNgERsOxFYE6RvGrk3XzzCOGjmrrktRV+OGS2sJfz5t7Y3Xio0tg39dp4
CXrgQFLh0whXjNDDpFhuewraWZu3Zu3QIDX0bHxiGz904/mQXMF178ee3gKYlFxy2riSEJMKxnQx
QZIO//GUNkLmLUtNcbvmkFE4sqkX6ZB7OVJ4rtwtA4eCc9HKCpWyuW7kEVR/h+5yhQJmCpWf8oE/
IN2PYUTzto49i3t3vpBjWhnF22gyYi9tlUOrCalzWlR4uRyMD11ZwrCizAmB3i7lUbaWqckU/MWj
NYni5JHO8IvxyXkNhdj6I9MUW9O0qvygzTZmQp2epVzbzODUt9fAeEOowlxNEHn3Zf0E9ULqpb7s
2uMVlLBmD7jb3e2sLlVXa8t76v54nWvZ0UuKWSkEhW2qectU0/FCcHoB/gE7LNy8HoRe1n3avCk8
E0VI041BQ65y7l5P4uWc6SlttHxmTVouE9KQbg6tew1LXDaElW4VrTyP6Qqa4FwhUUlXF1J6U0mS
v04Wkkd89HJgrYzu/frbR5/eYmjxndvEuFwzFk9LIjYbFSUH2RzAZrtW8UJwyTIZeoQNJNc1N2Ls
usl4AUEBeL4Pb03lJsSmK9mG6y+S0BGnCMSwLnvMojeZ3DMTLPrWam3YKujqHjqDUBdfHfkCr//u
8C3egI9xlnFpCkVqq6PO5n/csbuKHqWNG/hG1KRr4cmYJWM/jP4vv58+d3HzH3l+w+ZY1bUjMrLj
neYayJ2upT2bI3kuOW9N6nsj9DDhHO64SJEAh2/tTT7wWL0fzFCNIEVI4FGbg9QmDfdVsvdk1Gx3
G+gscAgO1fZkGX1RWyo86gyj+JV/53+ULnWZEmGXdEeOrSzMdxcvmuwJSd3H52mUzzDTPu/yJ7WZ
31QzPluEhIzR8Hu6aocJgyNG/EJHDH4HGXazg2w/JJnd7E0+37dKwEWLaS2QN0bhXBGXCDnz3Lvg
+p8u3KqorKZaSX8hX/CPM6SPQ/DJxPzXWUkUo/2xFv+bpf/KrMNHXH4/ziy46Vy91MPjA1lvphgS
cxTwaPMkkP7vs5UI+tSoOF4axpeBtZtLBS9CX7a/t7HSCeMyPrjzxXEdbiPu/FmStSf/qVG5Z6jf
EMfulgmA81V9m9j82NPaVLYJsvr8LD5xMM8OFEau4k6ydXmXaciFp/3i/675pgbalHPoGUtBUrbH
1MPTNKO5+gnedV7cfL9e0di+qMF6MJFBTPbklcW3knoAQisf0Jpudl+FgZjgcEgISW4MFuypzJOu
GK5WnJwcMNqV1MHMgC37bU6/SYJIYRzYJSazlhSZinyNNlv8BPlkN024TBFfidGe3BfHbsbQerHB
H7pK8sVh75Z3rFy0SoOkYCvOIDO/P644xjU2ciDkV1jgpwL/ePIUWq3nN9PTsxlORaggzl6tIZR4
cOuxua6eoPGJzyDZ4qPHiOon+oLsjSLt+su/l61xaHQYDVTuEKUlTP0WhknIkHGCJeFPrg9Hahlu
6/gHnitIPSq2fVeuzFeaDWNT0UC8QTk5m8rzd9kloHB5Oz/Cy9LFtp0UnQZcCwCDpPxWA59P71Mc
qhDFWbWZG8aXsXmjGT2V4XB38xrEJzGtlxhaA02q/l10epiEIq0STzZadkjdgyMSyJKsQQ+mXsBZ
YtY89OZfhAkDG7cIEJIDqW6lpm3N8UaaEdV4xSCcl6cdeMTI1hPam/O2lYxamtzq/VG/eueazXHF
LTR5J4bXrwY1bdLvYhKHnIry10wKVYZSJzDbrOUFA/7Nnr5EUFJTU/aguuWCcXmCFXkwH9m2XKRr
+Gvxvc9Bnx+Vzdc0KX1u1rpU1yoNvHJu7hhUdRFrFoCewAeKdm382U3ROM99EoMkwXW8aSanfDeg
YS5l4eBpzmbI1DT0UvGPwW1rWAf6KwvxhGCcZui0Q8qrFDzmCAKXCW+qUXN0wmTWoV5jTeScdOLy
bMWmQMRnlYTsJix6+FBnH7YF4WaZ0HlZt+xfdsfxz92KyKfAaGH0Qx7+PWFW5tmaiWhCnQsXsY9y
ec91mnT27n0nc8NC/IQ4e4XeesB7h4TyHOkp+9r6FkBopM05m6+TA/s49kDGXXBmQrWtzXB81lLq
TkYz/Ccg5kWvQ1mzH7dwTJKT9lUfAXCtZH7eEfMWEik/7vsILdE4Xn1ezNRA4WXOHBCaeNWPMK+z
DMd0AvMEL5kG6HFIYOBiFIMyRziFBNRL0JereHQCo5X/vxjKkjxjjemAHA5UANTqAdZfj1cI3qUX
lNe2vH17v0YuYex+aZ5fDu9BrJyf7kJbPfZ1pKFug1lZuuK1WkkruuCskkmCa4V5qmJUt8r3O50r
WhvAsbBRphM6K7KeqWvK9IZcQbop5dPkGJdCU9YKvygo2pR80Wu9zK1gepta1Fc0NQhABuOFmT22
5SS/FV/aQINOnHW/hVx/X5WrHUFyGzgHvo27/KnXin3ko3ODMburTtke3iNwe+9JUdjPueQ2JsWW
ChGQKW83TPqyf5P5qQ6QVQ57VHLeXgqB9wGbpqxNd8gbHHjNQruOdiJOnnUsVxcLmIy4FaRAAfoD
WyrXirorCN1zGKMRPVuhvD3IZBv+YThiR4oTTrIUUsMiaGO4Z6QFBttIj3KhhZOAVM4MUXKAeXfc
h2UaOlKaw9WLmCQdrL8bQE8G/3GJVGVzdAoHcdgS3NzE5YrwdSHxrqLnZrtC31VR/qjpQQUAK94Z
e6peiwvARvR+svfr6OP5sf4MwKvAp5LBWcY/W6UdqswaiYITvDZuCqzV1YQBFIQcbtO1e//0btfM
w+kNWrYd2otaf81ySo1FAnvbUS1UFADjhoV8fpF9UobssC6p9V1R37xiY/l67Ywwc9G0Htm7cYCh
FBxIfHf99JWkHcUI192hQkbqDwu1MjnbF81hSmYb8TA0I9F9c8kX22XkCnWtrCZNgPbZfosTTSfS
/JbmdkVRrMUQCru6Fh9DuW8Wo9HcR8YHXkV+XP5A1VA8yPJ+t3ivvrrNLT0m6hL7uvEhfoZ/I8E5
dmEAmxmSp+1cnlxK1iQHQG7scvEhcVToib7OeLs+temK1QYWiQhFREAigLz/7ll0coEGiYOadJRu
zmLW6BTBRTRn0byr/sgRGtVvBb82g0ifpUeq3uMoZM6HP9Z6SzZMV+SF8COpRrMAqFzXvW/HKhW8
DH/5kEfpCygkJmYkXwIqz0w2LiQLrNOc6vPqKnyIHlA1Z5MJdBlszE5RSphzXSlOc8U7yZmVXJjX
/dGexTSBAhgYdX04eg/1xx7KhRE/HxzvjMV6ffdqfB6+6a2zlZUl0+SnR3YBevh097VClkTFkga5
l7ndO1B6j0FMTktU7wTQUI7XKDFq/ef8eFD2z7ZSPPclcFlHRY2QxMSd6H3uZbRWqhIr1KFu6jHr
xXc0Je2TZC9s6Z36ztpiLmqWlnxU2XxwCslI9tsPs22TvIeGPuZd4n2WwTiOWnMTIpvgtjduD03X
w7vqQbSooYjdUoGlNYb1MBt/WxBsaDjvF80eEhMf2OT5caTg3spcJC91LLOgUAcjmFydUjtrdPkF
0rE4dKYgmaCEHr294dHidYHo4kMSzppAKOvVvwX0ilV17rIsJoqRsv7YgwtbQYyLMKuTh+zB2BIH
BPmMEsBiwzbFNaFCL5eYIBJTjGdKajuj0FWViZA1z/nMeJMs3i3c0krnyn39CYJfEidS5Wudc1zD
SJcosiL1OrM3Lx/ora/p7ICjRyzgnSy11EkIz83A1aLR7OBdJkPm3Mt8fyhUpunmRkZ1D1yxaYAo
swMSy1E4kDR59chl2v5XL1SoJZNjg3svNYvvp8SHMzxddAn98J0/j8ucKZZNyYfQL6LN0suEQfez
k+uHZsN9PpA2t5poZhnUgX17WxNa1r0sx6JC4W9bdUQ7fbCWZ+6oMBeBat/T3ci9Acj/xDliwW3/
UOIuY6qEb6wIJMG0ToLCXCXrZ+qB/d3ZiQnyik0DcDadoMaOgy1Y9TNcnTdsgSOMGjJSX23Zpvdv
+8ja/Yypxog2TpdQCftlmTPr+Eo8qmvEILK1NC9JWQni3C0fCtoHHDxnDTRwPm4T7gaG+lBSYeTV
ykMLfmDzOS9yIU86eWwrNagcNaYM8rHFOlMqER800/HZD9V9dSfg4DKsBmwskdL2B6NxAidELj22
lPBZOMkClV7PSeZE1ZAT8QLIVw/3+Xe7w8796OzYcjUyo8vQcAIodNJ4n/yWe9EAG0I/lRdxnf1Y
9EuSFbul3YmW2qWwpj+ROkIAChjFHFjFUndlzrhfPW7gbcTD6/Er0tZ7kA9jZO/m70d9m2K5pOiE
aFRkAvDPU9t6sQx38FtPEhXdvxqRcfXaAjJnJCXVH0gh8B96guOQtExEko5QMHTPAhm2/btyRPqf
cv0B9oAOTp6fdV5R+NEFC0tWeg4oPfWPM7EW1001iAFaCqJEKL5ga1OMWJ8othQ8OjOBZt6Y9+IC
8VZHUU+ZaqOGec8CrlvynIjeDNTcTmjoLMdXApk3Pd7H44oXjDY8zPN+QE8TbSfpqwaDmyKFMcaP
I8t+TU/i/USZ0oij/mRiG4xVPlnKiJe7gbNLZ14RQ48+UOTHXiViLopaHRAamLBec8GPhBG5V1/3
QdnfPEfzerC22lmHvzkO0OKbgyP9s8Pv/POWOhAFeL84ffwyujCuXWzurTWxO1Aqcb1ckB/vSXI8
IuIHfnE403hyqi9P97lRTJXjuclrMFUzo8hgMoBMC3VQBd8lKyTO7GQsMKuEvfGvXj8OtY4ITs9F
MdJZjqK4DgmWbV4SDU1pE81YHpBaXf2OSuc/nKO3xGcHSlEZCwE8EoDTacMucrjo/IRe8jY79ojr
2ei9qBKmzV9+9QDZISPwE7mAtiFKsLgl+xPd1hWxs/pUpEkaSoiYMXS02COLwWtEMcY/5k0AaoAo
6CGOvckPfxBhgLV4BRNRJm4tMVxB4Vfi7pTc1gBrKAAdgYI81tnLrbq2aWJIdyNuECNA/D+2dnkw
7k3bI2/0noxqhDZzfqbVHeeCSg4M+E1Wkcv0kAyX5hK61+qKv2zTOb8M/NDyCU8WNu6QffIkqRKm
P87/oCBBad0xUvz31nGH2iFljfOkgp0zdqs1ml1dhDp2HktZUK3EhUnXH6uoipChuSzVs6d5PJ3J
e4ROG8SydmfEubJpwRc1LXefhDK+Q3nXvH8TWFvgV7vgJ97X29c+BTIJIA/ZC1DGHnCFFph6ddZi
qAMCXTxkRaDkJAUaWI91MWRfP8UyTMUwlJJ9XCMZ63bQX3WxEEl51rLb7FcDjcT9hyrHbLXBC82+
t1x3Fz4hUc+5Mi6G4Oe0akAXUerjgPzaskdmH8twLMMfulFegVGkgUJjqoXCh219c0vLfPDNaNM2
0iAd6FdhUCnJJCOcyQfNgihq4qx2eRTe56X8UY1HqdcWHIrj8mtLAvTqjrE6nfZTfoB2wLG1sLzj
2c5KKMWarxn28Zh7WiSRNdnMdBfIp4ztrceHZNkTos9CGOrw2F9WbGCYh2fgsu6vp3nYGu2N0ebx
komk+UWIut/LK6D4Qpz51OHYNpnimJPBbE62kgmXJNgzsorFOLYqXqQadeBn+at4PTw87zk3YXVL
Jvx4sKeQiK+w7md43QP3QoXR8qX+/RnWxadq+9GrRuPeVqu3cSUXdV+pKPeKHAkhOE2hLPYQkosP
/3dFy46rE0MVt2w+lfaFEW78jdqNSF8Ez/RF9Z9ZZa3o+7CihGSgSikJIKDFo2OBvOwRmL2tYmG8
xDRkExtlN3vWZAHLAty0HUCjoQFW0S6h6+3vxvvixPnmLZ6J8nLIz1gx5/UMXKT5rd+Ec5uyGLBN
CXSDqUVaedA68Fz13haI+qxiwb+eeFtmhPEh35+oRBA54SecbnN3UcoyKl4Q2hFGVfVFMXQEDdnD
b9vKWiGvrpZYPOk8D7bfPU5QAD07Cw6cYz8hJrzSOhsnjudPlYTdMKGACWhlzyqMgt+iKIbME3g+
8FMgbmFbpFgCm+AIxTfsFJvtEUoG7kqS40rjpFmaiiplYpyCrlXsETP3IL+XY1h84t/QLzUsGvAH
iFChM9qFxS/QbdDrnn2KU/edrMZNutvJSyQOOW6goaxH1+qNrN/jahQkJEYYncILxJBY4oXr9e0p
dh5bVtQ1663YaB4a5ZgOmxPlO5+uhW242NiqoH+klBVzy+cLKMoOBcq0aHgaWbzaBQ/C+t3CJAWz
89vMzjDpsO1KbGLAWDpG6V0oEfeYxwkBJzVjsOAaTZz3tqJwiXJAwOkXgR+onduNUqaoFw5w55jw
JZx6+I3jKU6bK17wQWBYPCweZVlUoVvh+pyk+pLuk3d9BCabXIR2I3xsRNlQP/mJ8C2MgQm9O8WL
eNGUdhKmLPN8KhvjZw41o8f6aaUIpgKpv7y8jb0zHTzEizgUUPssZs7iGrfRYU82La6UxoQMljUF
5IKm1NUy7a7/1JR/bwcHpyV1TCZ1JN40bSooAci19q8TRgWIxl6lx56Dvm58LIjnlRGQkSJ5pJgN
hymmkf1J87QqNMvM3zxM/A3Vp+ZvcWoAjmWOp9aQ651MH/Qqen5oX5Ti+GYXbIEjptFZnng/RCQ+
mKRKXlfJ0QV79/DyNOv3Y0cro39TfczagnNXqglq5qTVscYXC+P7TRW4Cltkgvu0wGnc07Nkv12K
VezFHZVWtaJB2BQpaZgHL91uplbwl75KFCup3QipcENDAVJXNFXWHW77uMEjxmq1mRDQUrBrXvgS
J4wNA6l29cZIWH2Pt9ZIuSb54qEhEvhE+8YCrvjWxdk0JAS65spAhrNnx+p9gbqNU1e1tmczNuZr
WREjXuf3bbNw56FazoHtH/aXrAFdn4A75WOH2CoeQz0BLzKRbMu4QI1DcY2YYmMLxmJ7F9MLO+nS
u43x9JhcmkZ/5+r8OAgrkoqIXPukwpGDjq2CtuQTeURD16LE1iBlmoeLIJEv3UXLog1FDM1SC90b
TgG0QUPAN1gC3XV8cAzgJ5NYIfCr9DnBm3MWRb0sP2qWXefUJyXcQhXgFdm77xV+kQWZILTfAJU1
pyoVEmjy5DwO650ISdmTWRnFV3+BxkfSycaEsJjD9WAGVmjNr1xJDCbAByq9Bedu3YR/MeDgiCMZ
A62bpXolb7yKW6IcA+M9AloP0TfyO0F5Bqudc1TP2IyHXlZmoBVxXcK0R5/D7ts5NET0IdJb1lQC
TjDsmz5Kee4d/dKNQlD8MAiTr/CaLNl0CTTC+N8F+oyTMBom+H2XoUhd9fj9Diz9R5GFrRFcbPDY
DH1jYlpq9CXt6o+BnzbD+Zrxq9mIbv6bglVowvDJ/a/uYbDOFFPrfGWglcUKd5tpZhIhab7B/WyN
9Pxixyvbk8VchH1beQlBSxvUZ0U3ZVtGg7Dcl3fAzRmCjzrQT3GNIjp2ER65VCHbugAdY660HD9p
0yTspokskISgsKhjHKJ3m02F4lVxirVBRz40E2jH6k6jI0Ij/DLPlbJALNUYB2fMV70Qx3CD0ukB
imEIsOwEX8HNhKUtEKSgNzncwJLe+29BQ1SRMHxBZdjsO7FahGSZAozinYbmifw9WGBRu+5N1wlN
1fgrqlDTnJI5lskFvCST7RaDqkkT3lnR8jviwwhCSuFX5DRYaGhlD6uhTmQRg8FEQyTGIR6/9c/3
UUOQ88BG8bLbO0CnZHVtM8b1kGv4RsQE7qRuQ06mTyxXcEJCAB4tAr7JAe+kr7Iq5ippR6aOZbME
Rf78wPrtijOz+bwyqGinFqLrQi0UivB5mm/p+kCoY/7UvQtLHqgn4UF5wbnCKHkJxn8BlmE9yMrf
VW+VsHJPQ4PK2FPGH+Bo6IJuEprll7M3u+333UA63rqAcxTKa97pdD6HeNYZQgzHiI1NSQuXzkwr
ErEImPfYNhdW14snvb8l3X7DAoNIAnW9qO1MYg/l6mSOYQlbC8+y+U/My4UI0f3GqW2wIjUrXX7l
xLZhXB4R6UyI9d+rVBjY0oguHyRxXQiwsQvvSllbZavekcyOhvYapZ8iYwXroJqGM8LzlhavU722
kPaCa22ZnJzEqyxlBQ4DGajS48iXg5TzbieyyhE1rxzNYN6nABy0+NLWyuUb9Ckcmx+ISJ2kl9C0
sA3x4ZvWq/tZJa+b836es3qmadbpBlHh8XJsRCgouzn2w2da409tHKl90mO+3uBqEo+Z6w1Wdtk+
c7k15kHuEaXiObbHqb/cTXYgMm1d5n55guV6At+Cg4GrEu3QoPBS8nysgB0/gCOLKGVKWd0pecfo
fc/M8+ZBFlpwVAkmrThkM3iiG8LC70wMbMwX6wrqGstprj7pvbIuNCqQaByTiAP1o8zZ8num3krW
HpHhJ/6/dhBTefbPskSadNkBHIi+1xE+abm1Vd8Zye8xCz0AsEuIfEN/FT8hwQpLnxJ5NBQL4h6n
jlHatwzC/2QU7ge3biKOMxBzcK39L/x5P2j9WrtXxDyLUuyOD1VfWqqZ0zsI7MdHMs6/UlRuxR0y
Mw2FF/tyhh7pl/HbTkHDYBXTa27hL4WsbCoISj9B72TfFrXz2d88cek0g40zqZnno5+LLbVa3QCv
3IdGNrFQssoAX6qBRtWJaPe6QuOOsuaRSke0yW8r6dSWnMJj9xe7Nrc9Rb+MWt2FifTNjvvNeAfd
j9IOYO6Ef3ysFU+6JfMhLMh9/0TbzrRgHv1sa4Dha4WU51xVxROTz2+QSnybPQz5PVNxBaai18Sd
fm21sYWcsE9MojaVgqEnKLuvYXQzv4ecCT+4P8q/8txREOMfs0jije1Hxk4jZjkvKL0s+IZciTt/
/jZ3qldJINxrhw0Cm+0WMn6UneplX1853x1ZXRCfaF/X+REKlop8VGtY5DCxRnDDe7V6vafGmBaZ
B4gPy/WO6sidDTgr2glGUCIFkcB3uEdhktOlhl3I3fV6jc04D55Mjw2SLR4dg2Vp90Dr/7hSuTm1
hjY2UoY8f2xuYweMB5wVPV+plMx7tQCAevTrHv/hFNud8iFv4g0coujvSz3OjhXgG2RXlLd8QU6d
6F7oqNA85WU6WeuNHMvoOZ8O+MMSCAC+hUfPtHpF3dE8QeMyJEAgI5S3SIGD5jRaufx5pa5Be3P9
yMTgj+9gpMVetcWqg8qGqbTMfYG/QTLvCHdLdpbRd6/kEOYSY/9s2jknukEVnarWsehapatJ5LIu
J4efamCQKVZM75O+KAmeuKF52ca3SGV43YFPH1bD8miZp1HU6RRuZgn4GjGllSZGpHWrRkFoxOP+
m1zBIUfnb74o4FSjj5aVr3t1VgiMHgAXexv5XWB355YQMu9wEgRmJlPJZUYegeaZ9ITpClUKSNew
oFRzBbNldnPuDrDPYzq1LLlu0pMDGRFT622+H/H3Pp+aqOfpWF0ChvrT6wElKWBaiqEyQi7jgQlP
FR21l4/91BhRkJWu6Mgiki9N6l3qA/2jR7Adg7tccpcfRpFvSx9bKr4ffTjHvPnEUKTGVVKT45E/
xfyARQtPGu6nEg0PqjkRl3KnjlvxkRLLGYrmXvzRZcY9hAuZejT4HQMY6sgDO+EYotAKp0LVVl/v
OjwF87Ci1Vi8h8ulfxfWK0xMKeeseripoYtCDsErRolnDqrVu6iVRUh0gMkHSVsADkJNZhqE7sX9
ykrWqOywZASM3ReksIVFOx3oRDaM48S+FH1aOijyVXn5m0SI7yJCHomitd0luE1zxtk73Q8d10Do
bYt1Nb1kkca2ZxlgLrOS7leSznjtECMuRFeJz8qzPGxZN8UzmnwEaauZrOP0dMaCcGBYHRJKo14/
mPQAnLbnOqkSHYOVg4ePHP4OyxgwhhEQufPzRM7JR1A3SWIs7S/ohqs8AfzD5TcYaA0NAGmslWfj
GIDDVKUHTNsE9T6mZosIlzvUlAjenCKP61SMn6fjEHCOg1RVKtjsF5Gm3JK6EsEl83JAQi5h1EnL
FF2UVyiJPHmcuYqGNBZWG9D/zAhQbx9Bikhc753l6Mxko1CcF1bE7mBZLjpP+zaBZRcN6cgzCBba
m1Xa62bgliIG4XRsU1S22h+JYEoG3T5Z1UobxlAK780YiM5bNa4CkzYmFynVi20jZaK92t9piAzU
ImMNsD835TFCM9y0gERbjK0bPeY0HlzLuouzrlw39qot8adYKQntDFFCftJhbbDtK3pdawSfcdj8
eImoNpOram1RobHgUEoP3LwIcl8Ra4RJh/jgMkafPP/EICUbotFroqM9aQmL5/Ptd3aDnMbOv/Du
TsV1zNhT5h6nSZSzMoynEptwRrYsrRv9p/3rckZ2yatoqvEoJZfF+3lytcXneyeByyAMO2jhbQEO
VqNM4ShBywggV4efPtM0Mg3xT6/SZ9W6o8WkUitB6eZYxJTrL5r17jn6q80SWZvV5wPNhXZEP4z3
s6MprWnuJSEmFtG1wnl8sa0fTLW5/Vm060AcM2Nq6VkWB/eBdZiJm6csT2G4jBtnsJ7mOg+SJk5I
Yes9QUBLhbeco/ygtgLcvhnD0lWJVpv97BZer6Fxebo4O3qwjfAOYzSlZ35nsHI8sqNE1K6I1DPl
YrA88YZdzCYAvIAOp3IBVVOxYMKlcZRLWnL6Nz/c7MQa2HY2rgIvIf/eoI0AIAcS0Ffl6I4vzw5o
9APnnqxglVnlbVR8mt+mQOrp5wwEmLssU17VefvDDG3Iuk2PAc/Drp1/xpHZAmiLNHIBAe1x8q7q
m9iyAnN3I4igdkmsTScblPIFTMoL142siNVUulCxIYBMu5r3U87JLs9JpkaEihs9/fad4Bd0GFy9
xcYPwFgyZFriFvPKWk1Yl+D78g1qrPAoej4z2swhiKLOgd9zjpmVdREhB4l/ofSklXdmJVeYEmvU
P6KMZvPYJMIlJ45OGKiVGJBKHopLRlKwxM2/agDvnMmmjcbzMYXKfVbaGHxHNvJ/JDUwrkgzhKl7
XE4avYaLO3MlYuKKlO9ael69i0LcUVLcnl7MvfK/Uf2Vple/8RuVFU/72ryjKsOyFvYpk+w2EdEV
74+YYCnVXLS9TsKxTdQUEdnOdcGirXyvGcHME9B69aGGn3siJEIf1NffZ0Gat9s58kg2zAfIgs8u
rZXbP4xoFcJdnYyAB1SSdScjly3RmPDiV1azLm69Fko7m+yt9bMNRjvqS30WOBI4TxNrTAahUtCR
/IBEOZA9ia6wCRr9RPEIYGqY5Cb8pDLpZY0tQ0p1LlfObV9Zsq5JfvrofRxUdBNvfECyu6Hcz4xG
xFPrWGFwQ7k8hl4eROHWfFVjFPtI/hy0XlmyaGQ1YypZjgGTihDpISKM7eveTD/DHsk1MSjQ2lHw
f95ZFNBR2TEOd4Gh1AsQFBFcbC3cY6YYBfftaFtcXrBbDuzchgSb15HngbqPF3K66hXDvRFG8r1I
eG+YkCc29T+hZzQuV3zcXsGbxpUmQToCSo6+GiBZdr+EHOVXqTT8r/PhgkKRaqYheyZiRJt8s/eJ
ohEFYVXtWXwKYNCt60owm5koFvcsJgKoOpd0dXnhWphzVFuxx6JEzXVD6iIJ2RiXHPZYuU6d7SAs
hyCpCxFUcG9gPmWJs7njiqMl79BRInGtkldyuhxyRoOwyaThCeoF4VJuBMnTZp6hBOp2rd+FuUli
n1e4hOR09yHftUpmMIivC3W6CB+M2Damrkyp8ESMNOjFaRAtzSGw3gamjHgZdIjALVxH2S2OZIYz
cdJnnCS07hI7BazIdF4X5xYuAl+nTrm1pYjjSM6synwvJmOkdvtsNG/bmkv8J59SKKBAA4HCniGf
HHwrWy9cikW2UO2laFG3Se09+oy/wuW9E1J6sy74tAZMdH/u3dHdhE8FOXkRVfcP0tu6YInVf5Yk
J3hjNgLOb5g3QbvcMgVH8c8vEECdjKA/75Fxu4mhpOYYXghLYCJWBN+dmGW45EHlcpLn3Cgwv758
nVs7J3kqdpR4qqTeL6Jf1na8Q6uFde4A6pVPyf4sWSUMSWPixWcG0tbjXQh/mtzMrOwV5rwOR1+X
ZsmpLrWv+jc7MT/RBn/YLVYB08p7PHtWkotM7o5my0lTg83CDz8BCgk8MCxdSwr4jxieXeN6V2rV
XyExvY8gVgP6fSOpxBKpHCxrl8wD88V1ORtGjjA2u/xLnXzLDte9KS0XF+ol+M3tG9mIoprlI8yX
RA1qPGN/BX63oGYKj0pm4HgpPrPO2HcEgTmfUTQp2JHGhctA0DHybJYqI1SKG0FsMr+BwaCbBRsQ
BLMTgEhUJSsCHr1s4V1ei4WGBMHfknPEW4uoMqu0UyMAqcahA/6tLD2py0X0eEkdaYF4eu+E7Rsl
jldx1Yg4P2VTSf1o/rLyEAUjKMyXJsRZukh2qlIX0Ij/GgVOqi9X2n7uAMf1tCB37POcId+GNbKE
2UChfuSO7Nczvy33EIUHeYA5JH3DsDk1rgWvqhglWUrtou6qHAZU6NeH2x0MT+mCQuj+SgbRLk9n
1pnexape7zgPPWem9LZfxJuyhOVte7Gajju05GZT/Wbhml+ut8nihTfxtKoR6koZUZ+DtQOstYJ1
ZENckJGa99RQesTI4U3OKK/F6GSCDwoJDKoSyRXgmIrhJahWMZR4KfMSkO5lCEzIuImVU55yyViD
p04jtlNgpdVFtgfOcvrxHQuc09TnNhR2ntiwHQdfV+VlrMO0wz1CNlbqh5y0TKPNjSgUkwftw+tS
88Rxp8CKC1mTcUt2drH9bNijwcOjzLmb2prZ/TFoC9YA8SwjHWJinWhkqb4VMxnoaMJlJsYTedH5
w/tJXyE8TU7EbwQPCfwau2HE3NbsP9xMB9MfLEDUZlVb6Mr9sdJQVLML+NJmECkVNSk6Quk2ywDt
OzXSZviwC/ZfYLyJPsamiU8LmjmAClLiz5B3semQgVw4gRGfyBrkheT6asCOfA88hFRsix8kRrxJ
g+kc+lh5qkmc/JB2Ms7wne7oH1xYD9mq7GhziXa12hDGAKvKfk1hwq8v0dntoR5HQ8UChCapqLB1
5sglX7BtRh2G1In/TLuLYu/TDqe24d5zmPPzQCyoJRE46CJ+gpiDZ4cx/fo8UTgJqcYGRhm1nvtz
2OZG8ijv4f2FQ4iTsxVwD5kMGobNqSpBW762UlDoxdHLLBXbhz7k/Cl+rN1FnAH63TM4pxjbm2G5
DG6fDR43x23aCdHjtddVzlP9i8ZwQWIbOopcxuA5f476IC+g8rFipY1f1HSijnKDNqlIZNlts8jR
j2WEC96Ns21CpO3PEGR+mr55yTd4FzUAaOO5TnKGjT0L9BeDdEQX1z0dmeIyW+zTy2q6RCmAdj8C
jsTzhwLKrMKBvJten7UwPvqEK6urHn6RxBhpr2LkPGJUywA0YAcr5HjWXGUTl38jojIF9rD8TGWy
JXgFDvj9Q4Q53CxT3Kx4gbwI2ONoNTtMoM3H8HpDUhIzelhMk7p6VySdIF+YLIYoTcAJ3gObTQV/
1Ir3cSHK+pTnWxiYJJ46u3PR+gK0Mkh4JeHTmBI/4Nf4pVMyMEYhzUGIbMVAWl2Z1F5NQQWxCad4
5Mk0irDfNyDgQSk26U7JISe1axgBw7bLNSAq1Nq+q3UqpXWJGEiKKv4S2FYXAHQ4MfV47LTxQQv/
+6iRVV2B0J0y53+YHtR8v+Ldc+ppAkMvsfkq6X7Rj5T4EqKsbgJwWVMbjidxCHQXaBqgFs3gsHIO
YmJHeWa60oOx1E3PqDpUGRPiLu/WIIGNNWw6a+fldZJUuyECb/sbUcX9oERHem0EF0fSnnoiW4+R
Mswc0F2D7UG8zSwV1yxDfri92ZPldWDXEQtzbYCQkiVollPUkCo/o6mdtuLQfHoGMI9ucO+dECe+
Emav4roXbsxlqSVgxT9T+93Sa5/Z5LF/mXs2EwNjhFNTQqW2297t025Xj4tjCqksjhVmW1gq+uqU
6otJs4m/EV4hDwgiBuUWZug31p6KDFyGPZ/noQoRKuLnZy0fsjI6kd6lVMkSC7AW1PzMvE53kn/Y
nQycxdzT7BSBJsucZFUiP47P+aJ563/UpsTt+Z0J1QF/4vjvYzRuCakUSxxrFqxbpCRuvTxov5+b
wZddEkD0RtuD1zsSDTM1Nm0oSdbSJ/HaUn6umY2wqwr79nGFiHF8RryzFTz2sqzB14gqqtpfs6me
/7eh6yTbxidbX/pgqcRdTsxu8gInQ9i71oO73KNjNMw9RaAVa6Iu2wRK0caFMHM3tMvGmmIN8tya
xLNKxS5QymvtH/l0orpFrz4EECdGKz3auJoP5RVGEwU7OnQHvVvtgQ3irYbj7tKnRpgqdidNyJ0h
kB4wLg8rAGapwN3FxQ4N4TGus3b7btQU7s2jFH35VMoDyAukS/zU1rw3DEznRvpsR2vHtxPaG86w
QNCDlVVoH4MKNRaGkkufUmCjH1jiEwJ4vqgOAJ7LmvzhtKNJ9AeV/q2IsY7WV0JmgzBoiYyAfXFA
N4UCafj7IbhwUXjboCasDEZ+jdEtDUQAZgCmRxqW7F6Wk9em739R7jIcluTsA8RSk7lexv2YkNms
ihoF/wAZifDJfzXx7WayDGxx/l74kdYnSJNeOthGWOZC2ZprSvh+KoaU05Rl8wH+tnMdhJ3+sQqH
uxc/YzwbC8kQsk+BZGzyoMv/XUjPXDECl8IzXzd2XDq6ZbNZRlFn24/GmR0/4AB0snOa8fxi/gQn
ZlimngdPQUhLdxbJBjCtabDsEWuF5ZAUZijomUmD/fK6hq5Xmff/1jb/RIvS3qXuNctDEQTfNRov
n8I1BSrh1ZBfxNKG58lp1rOYncXSQv+UHZcsA1uXp1A2rJD4Wb44e26G1rh8EznRBjb36KIw4FSi
Y2gXKJa9HzpCnEBB7lQ0+DNRxI4jLL5K18kuLmfMxT1+TjqGTdywQ2M6L+9w4TVmZdLpZIK7VLd5
hWRXj3nNysh4xYGt7sN63EkOyfvekuvge/it8kLd4kdK2y5swimdQFTQ+uARRAZ253ZKwUBKGpa/
BIymf2UsvgVVreuECXFeqVSa4pswlPI4qNOcAh+z65y/1XetXZoBdYE6fVbNbgJI4OrvGBOUhbmW
G5jZCHmY3Y+guT4QMMmhoFegXP0Xz/61ARR6tg5ibgbIexhZ33DGnYOmORKxhbVqAn/sBRrwJR+o
H0SXBGn+xuPVBoMCYFw0JCTFSPpAX5Xc5NI6ozryY8PvHj2ZiiB17wKCrhDxPbSIXjGrc6veEiIL
5+67Q74TZBmISODUapZuC/AHA3CFb+P+rAk/VUQYG+8NG2i9MeSNAWiJFcO7Y3HP0EcWgghzGXQr
I6HqrSc02LUjffWnr25te9Bf1Z+6eebvtJj1Ag+Mlfmxl30ctKlneodOZkgzhXw3m0WuMkqqEM1/
KC0dMwOXLUIXxPBQ2V3qwA3MTUCwtRtvtWpvG9A++RBeZXZz1lbVP7JMq2cBoa8P+PYw8NA8PucU
D54HXZSvrPtuAgPPsSa9C0OXwOCATx62X1GJF9BolqgBsX2RoYoHMU6baIOpg4AXcW6w6p9cF1s1
KlYTtzqYccb9nuNPAxf0Y5wn/u8/FtreaWlZe5k1kBjy+Nr3DH+pex3VKELie6hjH/ngdgPgZfXl
VRxfaLDmDQt9iuaRBhWu1otrrM6DXDH30q3MGqXIzphFM8C05XqTE5ZkZCVTIHcx47eUdJ5nDG9u
DiMrmwMQCvm2HiCO479IOHucVKmlMyUAqbV2wOobhZ5kKpOGjz02zhsiTOGy78IwW8WcduycXkDG
tHZu8pGqIDI81PSyuC6TDNO7SlS23uVhLPLyP3zBefk7HkQkV90XHVpicVn+fDmzPjA7gnKtH1ld
9rxl0YhGziTywkOLa0huuDnoA0nwkcZuTJgcoDAwmbxM8lVWjR2umohKZA5HviDhwmAibzKAL10W
qGX8NJkf0I4/yC2sWfjugIlX0cRwhxchFYe64TUumJIWOqaEBCwixaKk8a8tsDmuiXPLVd3zgdp0
uR65Je+v1H1MNgtRwqyr8Ov8n+0Nv3cmLYtgWJW96+bJmf1z3CV0TnOz9xeqA1GXtTblc27Vu59Z
quUAokj834iT6lKjvVGHAqBofa9K7OMWCMBqCXv9sn0/Bx8QVVP67ckG+6Pm45hd3I85NdtVj2jz
hvwS+2xaXVwZpCWTWdjt3XfSCD76zoyxg8bxCuhbKJbwcsuPjEo4RcuweHsyk8cTxJtcseJPi8rF
xMXCHvG+qf6XTpkz6F4z8uzuFooLu2D0c2+OHARahKLkx8qqFBKbqmBin7f0qrvkmR+1DhqBKaqE
3aYh6aV9J/YScWIskFCmxARhHrdDsSzQg6VWQzs5wYVvtpz2BMG6WRGH4JB2KswB5B1G7K77bjd9
CyfSpxiloUU9BvQEwi8ZtyQLvHIM09RRET2W4TS7PuaunbeOtn1iHIJINer4esIAVj+GePqZleJM
7y8yUxbELXrFWqMZwPzs4gaPei7kcW+UhAyBVJufE4IPA5m8oTd74MLSkWrEUd4FYumOUEj3pb44
pM0fPZEDeCgRuJr14d/O1vo0nJLY8NC+jpLteW0zGv2MTSSyhVAhzLuz6qtgJ0kr4CibmnqLkOxY
mH6cZgHlREyeguKD9FBIHGFTPJmoeEXhybdivbMscB7Zk639I4gGgETLFunk/EK2A38ZecRHFCAh
6DZTccVGtJUe4gFC1GECQxE08MAbVmiDvUQReq6LaGfYGNZtF1kwXVpDd87U38n0WpK1CDzZKn2S
7i8Ru5v7E7HgSMi0E7jfce7iua5clVp1cRoc3AMGkaeEfWO67HWfSHE9YI9Ct/HCX5UkGt+q0Oz/
izBY58x7ci4aTKwot6g04EwfpYxDM1RpH10ym0bB+DCLzNlem8Vxg0/J6lFzCJShOYiQV6crf3vt
yPc9GEj4VEgXiGEcNyOO/jgspwsP5pfK6AhebCQibvOxLvr6toyMjIX3WC4YbhBjHhwGL0pEbFzZ
sD+amPXHv2B695DPrjtUSJGf9PKzC/KA23tDTMjuHGhyIooGHYozEiB94oW2pKtrTTSk7x1SzNr9
ntWlIeE3EwSaySYoHSOS5Wwy4K/K7f8T0N4KkiuXAxfnfIkTAo+eOm8+RA+5LMkfRwKxavCmCATs
BYKWEryZCQa5HBiz3VqVSTa9JlSeUNZSH5IkSl8mdC+7iWPmfhnk3/qRCADS6sZgNe1kF7Sn6bJt
ekZb9uqrdVjDJfSwcPAZmYXTq3kGboTkL48dju5mXF8Oid4KAQwFtIiAU+H2vqNYpOqUBReddu33
XCqhDeCZuMMR+O0jkOEjivZLYg2Jk+adr0HULRTRGwTMpsQQLpsl1R99gk1d0XuUhaLCc6qAqZ+K
+oZnrQ85loG4ooAA+q9yh2XgRbjSRC/TtWgU63pH47Kgxpe7whLzbvCQhCcB7Veah8YB616t2PjK
wUQVaTwmWMY58nVTT4sPIJlrV0C9poXyzhhSBIB2tu0gnDTaBkaN+ODfQ3cH0B94Q9oU2MdlhR+g
B/0DPPM70IVMKu1uzRumQzQjHSo6wjANkKLztjJ1Kz5LWfdXLjTE2RnBkV7FIFK2mSGAjCZ2T+bc
cizv6lRbFx/AaZpjKTwVLudWBrKcmOURd66NuPKxIshqXB400g42xfJelUwZJUFajeyeIylCoVi7
W5xedTFpfdMnNJIVUS3iY8liyGCdZngugrvXtHeUUseNQRsjxhA3dnYHu3EPM0jCUKm8YRApbPJL
jvA/BivRkf810v5UvIgFAL5SZ0hxYrNRrNX9BO3cqVh8GLFfOdaa0ogqirCp9mKIKuDeNWjiKQLH
HxmKE3QdKArI0VqJOme2Omn5bgUWRfF3ysGC4254HNPobc+buboOFj8LI5eLlkZFOew3jxEJUpHQ
jOAK79fWxZMLKORyfqNqDkmiJth5MJJ8oaVBq9SobjUbjMbJYU0o2MER3T+OdiVsQeveJWn714tL
JMq8SIDwkeiNh1Db3K7hupkLB/IZoamQaMpuqDW0z/onxj+vFYXpJSD8ihMPNshy0gyFH/sjTKa9
L/HCQwiUh8n15AAUAS5LMoykEruFmO/NSE0A84WGJAHKh6RVbgaHsdS9BJ6Pk+TcSCsGojQ1iMtK
F/SgYxacxVvyCeL9xheszC1niQ0uIyYWopLVraWnA0QpFzpgrnDH/MYhxyHUMIlXg+9O2eKry6tK
OLlhfFFfIPvv/Qzq7f92hmWV84vhdUu2pDPp9MZNv6VX2OTdP4+XH4lVYfkRl8b9N8VW1GwZE8IQ
IvWoP0yZO1nPljezENi3RZwo/riwPEqI/jZjWkm9clshvM/MSAkg/NSn8gtBeaCWM+tgTIWOTDhC
hAJGN8B2ft7aJfIbD7zjXyrtNYVndEwLSU2dMsklEQilkfrMoLda6jPAHE4Eu1g09OsGv3wk1CSw
Tx6yQN9NIPGCJ6a+8UV80I9m+0E/Oylb9YYC40Gm+1m5srGfgPMm0lBR0IZwGyXoVsqLGMNEPzHl
BaHOhrYq5znZooqiIEG36wHiQk7WSn+x0xP6KiiNYDpleUG43LJ3rk9+1Xbe3zE2O14gynhjEWAK
f7BfY2A9XwtPTXNSf5OyYKutAZVqSqw5wHNYk/qURHPmGyJ7enTy6YzimZWztO7d5/ZI1Lq0xg06
HSsVOWtGbWXif5Uc3RVDBdoFELKVMgKXavM5Hs2vt1V6DDWjBeUok2qgnGHmAitVG/OR2EDE67iy
D0iWNnYFwRFFpeEkAQ0pFqWTTvuZFKxxAYsP4QYBkIw2jKS3/fr2ALS1HAFFTbhqFWi6nBnAI83e
LeH7fhw1mYG6Mb/riY7wAlETRmWCn9Hrpl3Pqev2OkNS7wcL7tng9I9j7cyLsBfv42rig7y85dmU
NTR1qI1YgartqKSaRpyBtoaxunbpqPTCnIe5K/5yUglFFvQy9Uct8IWlex9NsCpOBWAh9hqq2ZW6
+S2QPEuQHSmwYW3CPyPPNpIf+VSSu4Bsj5WIjTRARag4lzjjOtEOqwNhQDTx3wi+3sJyoLSzH4yN
r+ajClg58WAKc+YzwKntXkZTANGgo8kPi/V9vf6z8+vxyReDmtnX9J88vbnF1SDSn3BS9Ce8D3+Z
edELzkewM1xMsTyyAQTByda1tjcBQL+U3H6NSt9CYcXrq21mXJj+9sf+tHcPrBE3vITmb50/VUA5
S/wzCinNF/p4zRzFyV53rFdRTg92wJitjxr44Cq742zR5JFVHFBgh3xvF/kO8XLzYK/B9uyWXzPQ
Kl+SxfLsQuXBmbwzm68WT5NS5TPMWFD2PkakDHcolprsl01xBTkTEUsSZNNIwAkUrrhCdHxgPr3e
JNnftbKbIicGTNZJEtbUO2bD0JwjVtem9+ryiFajU5rxQi42zxaWZQna8ThJF1445EKHiEhhT8Vn
89mccZK/AGuaBEGsWhVyKHmSMfyUWoKNew8FitrQBW60h5B5DPGSxwLx1IyNsyGsWRBFCWZLNdTz
4Iy/xiaBJgT9L9EpXj/hUqRtwmh2q6jY3HO8vD9wHjLzw44sbD/L9Ge2brShajzQKCj36w7DHnmf
LfntGpGjasDawFdqyPoUfWUd79syK5SR2gyI/nAXazPDfkFrFTvZeGbgnVtRKtNFcInb4/8jqwYv
yxbICYXsur5UaAg4NF3PQ0DhvfDOQak5RBXJ1RFK6fGduDdhiQNf9Kv8nBeSBbaeDsGspaY3tLEW
8kZUCbGoCd+v5BjvA6G2RJmUFhjoSDoHaf+GOAqAsV/07iw9tQ+uUQI4PgU+5meAI9Axgp8Azdxm
NuQTvMQNsXPT/rEb6Yrcx8hKRSTtSVUjqXsYYy2rR41ID935GRo3LpIznmPmHVWs6gNzVuCEeSJm
u1IqA/cYroHaHtXxdLW/0dVTYA2A7APO4Zm/YHezWFWimRn8hoCCfj39sAYsJHSBy4uEPzNSw4T9
fT2PHahH1rpSUKpT6oQd9tAJzMnBzdAaHVLq9PX2YwGsTixgwDcV1Qxw8pV08wulzQHz9KRn0jeV
88FR65dQy4PuIS6wW+ktam3fUxeNQZ2vlRZxX2Na+ZPdPzYVfVv7JQjDXB6mmwoEOQR1xNy8soRV
AZLFj/JPcgePhAZcFllv5NzwJG+OycmMPm6rwJywb4ozl6IjsxpHYbpPzuEnVk/wjaU8rqR9QFSG
OKWZpL6qyCHLoGnz32ucWp1pMp3YQkfqs185iWguDWjtQm6VyUA/+VsVUfgfBcSCshBiXEVOFJ2G
V4nOoaAB9lrmN8aUExkI5WYkce5P+wSVZbO7t0NvadsjxazrjzFHm7egMd+razAUD+uk5Pg82hjf
21MSqy5EM1goxMRUJyReXVTnvK+hdtSX3SgjdruR7O1o6cZ5fBBnPSYlZDRIFT6Nk5laRjTmNIzu
PrWusFgAgnVR8Gy90VBKG2gI9G/2BUkFYdDu5AdIjHjGAPt+XY4Xn2RlGzAY+pN78RbiL8kXQngF
H2p9Jriv8Eovfk+CFIlQw80jot2HREbF5MkmArU7SkhWCAt2ELUpzfxXyki8vQLCkfY9b1fGuh4C
yZP2b7WxCDNcmfPzRIZhPTOzkcSqcYI2iqaoZQFsgoHAYRwdIbUl1p0y30v1XxWNJFuodbh5uqeN
dsa/sMjoKZkcMq9b5+veO2dWS6yOWVPw0QJe9ZPJqX5tggEH5k/MeR2UgJ7p2XymwhDW2E7OjvT3
aMR+AadBg4mzsqGKsj7A7Gms0r9tFXiWz5sH8je4FPSSLHNHPjmy0VlfdTGMBJ3oBi4vd99LmLrn
yhTVHWkCXP1MqlNRnh0Z6PJnQnmFI//Qgp2NzDyvfHp0dc6ZlmRwnPoBjOvfnEMqc0IrlNobuWA2
MYaTr6KP9t9nH6x5hsrqnIMWVLP7WUYnPN6pxqIc+cZU93dehhAGSNL+zs9ZUhTUu9OLuOpEcUFH
uFx0JcZkBDKBrBe1IKYq+tNZmsVnJFvzVe93zPP746GeEHisTIZBi4ow7PkMgiHQQaIEMujKzmvx
yQ62qHNUB6thOhos2JVRQ0Y8IzII+O22EmVRoF1N1xbGK8O+aeijdpCQGvBlaw7XVJsvE1GuBT4o
FGrLzeqmmBgzYQ8dnSCFTH73ppmDwWGnTRs7S+SUAXevxrV8O/nM8na15Ml8WVadUCMOCgMMEiNY
Di+nJ9MdmiueKsUj0CmPh0pqAxO91qObDTH11MMPd9ZzmmAzPh3Cfm6IWyVlbLSaqSgDxkIHza9a
B3iws5Hugo3Ig32n7dYW5WsWiYQ4vNAjlxj6y8tShprO3AjIgcox2sWMCmTubn5dQ4aoSvvEuZ2W
/zZyP17ImVBoFFfPFStX9/LG0NPEFwhMnpRkZAkv41iIrOrPsJHeH7hAa6qVUXzLUY6+rM5OZEvv
g0j1OANN9LKIzkl7XIMEg2Gu3Bq/mccH6GK6cEOih9iPD1hLzIQYrPapGv2wtyenZKCxy1EY2buj
LDu0brZ5HeDbLhpQNMHE7/iP1vYyyM4Ww0cdzwiBrV+oUfrkog0tIJpeDLT2/ArVNVKizzVeMW/D
/v8S0vq/8M+1NnWOTLCW3+clox8+mx5EP8pGCXFh1gEnU3FRAkqvqZ8Zi6fMin47TutNS/nLn0oM
E10AgqnKSDoPY/7neNFwP2XK9xzsOonf+EH44hHTaNKRF25J6FVPfEM2DIjff0d+Y2n3HWQyxhJG
sn7kzNETapM/30599JjSIxJXoV8ih4V0yevZyfUcBpmXIrJWrq5BaIsH69chd9v+lvtIB99p5WdF
dJ1ioWf5nk3pvZn7P+GsyKKvulS0wmKu5YsP89MoG4bQ+PHDnGQqeKaiQhP6GYYH+qoNW1W9vB58
Gv8bhYVfaOjLWfBmWxy6ikuA7AV1Rs8VBevqEuDuijMJ1gOFkD1no3V9RhqEs7W82e6m68JD4cRO
cEeDqOZTBQgZ4ArP8QQE4St5M9sgMvEPAyPqvORebI8dvYjb8Gjo8+s07X7E5WHoOGJOzkmy3qNl
KZEt8AcfPq0Ugar4+9IzojG7MXcRt61zHCIM+DO1L4s60dz5H3IHQFHb324aB92yWfGYR6P0VJ6S
MQ3qP4hWD04BVdUbut5mtRDN1esCOOjlITQT6FdcG7dRCcni/sakmdY/P6y9cpTIs5RfU07EFMkb
Jw3sOjTUGzBI6/R4HwZe62P8TK/UMD5D9EBl8GLzquOmxFQoSoiZ8PHXENpr+RUC9XGwGhY1UG6c
t1GWrGFvvuibVQGQqKcg5C71OowhEFCAjFQ7mRtZuMSGQfVhndhngBxQaVvHfsG2sH88E91maPXW
o4yTr4as9ldeLO1qByxOb9ON+RDQqhUpiLrLeggPzJdPwmlmxJfpJSbrGGP70VeoZd283AYIdFaA
XWF9JGlCOYw9QfddYn+7Z0Lln/wgEm70riVvlNwo78lP+937Pe66lhWO8ce19/StGOjxWKVZ6szL
JzUvnwkvP1l9PhDzqpcTxOKzRLjHa0b88pV6vNI/TMdYUKGQEn2MOac4l+KYZaP/x1zyqUsTO9MP
cEmRUIdlh2h+fKS2iuInoY4MkoL6JSPBC7loEFr0WWzdTNyDb/qqDBgstlO02XvngkxFQLw4QlU4
7Vqri83vscYVwj3gmoWykwfaMfDbOyAQiuY7HgYkR9Cppkafy4g2Slfs4+zPHN1hLCfCjadE9kEz
Uk+n+ZZ1sK+m7rc5GeE1rP8HeWBAuAGGDf6UoY1AZj8KIh7E0/iwDoxVr/DgzV0uZi6lvFvR854f
Mhrsz4rPtoK4WnNdWduLNdFKMWI9SCOLUaPSbrKXd0FErIqiuNI/cKG0Ez8ordoqhnhmf0UrbGrE
MOgY9vXrbO9tLXDl5zlPbqA8CRXV5gXG9/6g732kTVdZL1u7Htsq20/HB4lrZrTgEdIBsHRKBdCX
iOy0jyTHZ6A12HOi7WynHfrpeTcMR/tmZEeD4x1CZUm2VJTPNIWqis9VoNQFU96ltcCWjYZi+Qit
5OTwnQY4E2uQaP3QC2jeRtpob8EnStCnIxzVGK/YOS3ECXPkXBGAcC2XrJdAKf8kEsuuX5arlW1f
vgBkHX0EE8VA5YB21HQ4GHxhoreIoATVGlGc/rPdrsSr04pNNPVOkvDUB7Z0W60kF8hj+kAZmU2h
bGkO7RGOtTDwH1wPPHdJXvnSyimy9QzziHLl9q9r1sSv6qutv3bG+pG4JVpXamcL3ghpjnXAxEhC
K4a3O3w4WVtJhfXznH4qDvgkFi8G4ZyMS3mMuGT82l9ftwtHRhdGlLcJOsCb9YkJ4TpcH3EFdJJp
YAdo6Eg2zmY1SJ1Qeqn7Iu/JCJ55n3uUdCEQW+8Vw2AulDYkYwdfaivYt2xv7tpnwJsdMT5uJLuH
1F5yCS0WufkRvMO32ItiiYlbUHJ9qqfTFrh60USQMfHkocDIsG8IQmrvpbvcr7Sj0bZTTPXZnNjd
hdptrw4KaWFZ2ePweJpxCVIOhBEaZa0mJQRNATvCXz0trrOm77x0FaDynFfTQq2Tlp4o2NpD0InH
yiE2CguZSR+mpAKrGQuYcyx9we9IqSlSIZAuZYEDXbnJgQUpizHlgOq1XLGfnGYahxkpV9s2h/YD
tOWkeSB87Zd4OQZpYpVuFJu4TagIk1K0cSWIzrz7aYgf/TjRYsAWTILGLrrigA7uYi5PAKuQAyJh
8A/Vm+5YR18llb1WcriExAiekhsAb5Sc2t5JIBWSfvgbmjYfWs3Ar/PIcV/jmQv3t/HsAiGfbtoZ
d+3ZjSSBIFLdKmpsX7CJpVih8142p46b+DMi87Njj4ZVGPSN9u/kYx9yYhqLpj9c9IVNS/peL5kL
zOwoyO/h9Jfl+0quzVFPhzHuQeegU6ZWPA/IE+tJ4z/DIfC+DD7sB0NmMcsXy4crwoEMLsATOXZ3
GQjHCbfaruDr0a5AQZ62ZjC4A47kCZx/Bcnu6beSuDmQ9bHJnkgzHL/i7RkHtGlMYeqci9X7ZyJU
k0VuepUjT9oMvfHB2PS8x89ORIPeDm9OyGR71MuPOmrNQDP/7bJjYWcPP6vu/8pSfnVp6LQc1KRN
iHiRZbOWMTv7lJcKHoKe39ZnsYEspbonbkSXHShlNHfa3i+2NUe0bW5CO4CKI7SlwlpoJ3AybeuT
FZNx4YjWsBbeg1A9uhaubJYoF5UxCIC3G9vGYW7Dry1Xlx47TKMjF0zD2xPa0MYHk77fi/7+0GQ8
Cc6MPiH0SjJanniAceEaZExC5PUrwiUAwrF1g0CmgNT58wcp+9sGuC/7JVSnfkOvMDy/+3X30Wiw
PCPRITljIfSF1q8f985ggN1q9QSni/kp8tYa8TjxV0+btYf13SkTi1Vf8SzAj5Xk9HGKfBeBXGxq
Gq5EozuZmI+81fFH87ATPjIe+h689jlbj8PjK2FNLi0gM9zD+IlIjbtAFsyMmGs3znqrasUpRD9N
MJv4PoZBwKfpVlZl2vqUMgxM1yYZf0VkVHZ+eEZRH9AftXnrg8IQJMRqTH2sNB1OqqsHFCRpkQNG
oq1hs7s9h28gNi6msQl5tKQKOnLvZZQ4tIBfmSfkI0iw09Wi2+wjUwF7wtC1j2MQUR/di6B0IjPc
1kb4suLqSvwtxpb53dKswRLgTTSS4lUtmIF11D8gj2ftDSgp/m7BP8C3aajtQcypf13s9gS8DK8y
a4F9n+4rXJjsRqz0PKTLHLJbF+g/goVwThw9HHql6kNQNn/l8aCF9XLdLuVh8+2myjfnw7OFX/sU
GkYHtdLuMIuTH1H/Qylg80EGVpogUKqP2qubfmMQuQf/yvTTBlvP1/Yr/U3Rl+QzRCfY4FVamaHP
3DXVQtSZlTlRtJRyAfpkSd5+JWd1QGS63FbVOIYHqIgrDXmuWvSIj2jLCqitBJwkNZqLM6Zvyqgb
QQSfRRwh2NbFMBHCTCO+SVxPObriGYOYh0oG5UCkAyt0gb7RofA7pibmq5kIOezo5yYjpvnL/vQg
DFmsdiQm+RAc1dT0rDovwQEPVKmlMKTkgkWPoHF6gEiFYlFGYNuYJtxPcThUCzUrR8/pXQpGDh6L
oW8L9nldMi7l5Sp8yKGtnWRLolMKcFY0OZO+kdfKrgyTDdpXo6Z0w/Dr3FprEzmiUfubayS2Gwno
ZuJapxFVUEofSkqm0+ASbOSauKpQUNXJbIBdyS5uRnGTOZiPMYTFOBIkBJXc7xN1rXJ0gxQ3F3tf
h79FdwvTO8uPw4lYvxGMmW09kE5o/OWwpGUKmKCpjfnEyXdMK01oFqhTCnu6gi3QTF1JpqPk0ZEw
JuBFsZRuNzY0f5ZQZ4iyd4tkR9LCGPmJpHegwBeTJJuZcBJDZVbNqD+wumkpcvObevCggo0LtCWt
9cvuvirUHTjA2Q4BaRPNxAn3SPAPADRp1VwoI28rctm2lPqQ3nDyrFCChZ1ImOC81HdfYkwB7Kti
NPNHMMbZikn+JY37Rdm3k9VjnSFvVW3/4FLO6coLDrIE1/oHv3ISZ22fYbO1pv60iWMCbfme4bon
wLgkcksoxOFQ0+PnzxAfB7vbLgwXPlgby6LnUUaMf5g/BlWKcqehj4bPjXjx1G/w/hJj5uJI8EtT
4I3HDw8aIsm5zmd0XLV+r6FrACRKrYwWH+0DO28YVqhLJ2no3sCRN1hGpqLbXCUT7rcGBCY1HXDb
YLZZDVGZlIzqsFp9PzNXeSafclo27cUrKVqSXviXVbapvdEvNg+6BGz2KzyGqamQ+s6VdXaT3qib
XrRJEbn1cZoBi57W2iu4e5yoZOuINHD0XnPrMdRVPNkiHD1jEtKSK9iNYraB+GA7eJpMxjcZioUm
IuTQ3raNdCPJ8LZMZzqRinSlsBsMfQePNvcyhK/VZ2etxZMA2V9jIONfLS05WeDGd2CyCPd+NKjp
1vLyyk7F0rKJoF2AxVs0OI51H1aM/AN7zxvn4eVdQsA8upr0J2XZGZUENfQNmQvF8bGd05JSLIjx
cusYNmFLx1sURI5jpEV9qIX4bf9RWDrsEOqMcu0F0n6+2SsZ2DseJck+xN3oC/XD3qaMv4Y0ZlTw
vvga2AOhmhgLCk7yK9wGdGoZxxJ2VlT7X6iy3zS4rC8zTth/3vyz5f4kIirtabg1rWgZV0pYFreG
VqZgMTzYdqo5eQiFG6yalh9UTGicGcCVuavuHpSKwmaZJgFwZPKxxwyml9L+ColojpZjluFu8pTK
v0WBjReoPh3zjN6cYD/YO32JfjafpQYa4bgX2dVQLIv71nMqH7DAkN65MMDY9R3jph7EQq/w8WM=
`protect end_protected

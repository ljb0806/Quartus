��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�P�)Bs|mH%j�w뿲��[Y��,�Nl[�$�M��]9`��\ﱭ%/��q]���}?���������aB��;�L�34�_��]�ڒ�謽�`�VZn���9" h�@kKJ�p�jk�G��^9"y�U�`���/����N��hi_ɥE?�"z.���5-�о=I����R��
C��Bc�y5&-Q�UM綾/�[��?����1n��Xa�Mx<�����-�*����:}2�|�Ͼ[`-F~�c�?x�,��'K��b�+����*~Ս�-�ǟ�Y&�ۚ��}�Z���I��?�P S���-�`����S�u_J�D�|��-�\-ӊƞ-K��M��	E��R<�9����L�a�����"�%�!������>�o�f�Q-<ǵe]�_FؾE�bJީ���m����:�Қ-/iX�+�_����J� jcp�6�.p�<�!j-&�����4�(��DB��� ��1�'��䊄y72�T(rS�%�
�l�1�{먃�nW<��fJ��Z^3�#U�U%�n0�"�54��XK���������4���w�c�I,f'?������*B�ߒ�p���x4��c��C�*���E
b�̍d)���{����>?��z;M�i�W�4���A�(<P�;�����[I��[��w��N����,�J�:�?g��Ʀ$+gu�� ����簚oVZ��!��V�ݚu����l�i>&̓���-�
Eb`�ّ��[����n�آ�Χ�C�&;c�(��Z���sg�Z-�\�*m�E�X�y�\��hr)�;^��ܖ�Ǖ���B��(5��*��ȷ7�%_2W��T�J��@i��ʜ��2Rz���Mj�|�h���1H�H�n�ꑩ���&���4U ~��v�[���cr��'��Y�n!2p������*@ѕ��W���,�e�=$���08�j��^9��0�������*�z�w�QO�(R�.�n����Ku4MGsS��A�9���<��:�kɕ>�U�iK)�<����Je'��r� U%��
���r���C.��d��pQ)O���Ӫ-=�vq��0J�C��ހ .�NS3{���xJlcL11m���s�\�;2�����"Ac���iMgw���W|o}ëoOӡeN|?*��LĞZe�8~`��QƇ�b��Y�>O�	@�1�H:�+�?�7���q`E+,hq��`��*0�~cGYN���v{xPm���a��&��Ð�kBb_)_����8E�s��V<�@޶�qF�$<�Nl@Y��~���:�2�ЕG����o�fZԱi9ܕѸ^���y.�{�.����3�x7ޠ���3��k3r�H�<�r��ѓ��z��H!����,���v�����d� {P�W=��b��0D=@���v@���LQG��C[Bg��:����mI�����ĭkҹ�(?�ZI���G��z�����z+�As
��G1��@R)�6O �{aE�}�J�:�x2�h����~q!.1�Y�j��$*>�HO6�����7AOJ~�Xb�c6�ڎ��ύ��q}y��K�KU�븗�VgKa��6�У�%�!��Mi��)�QK3+t�{ԳjN]�r	��IǶJwP�)��I7������/�O��η��(�_ �Z~�������Pd��b�����X�ꝋ��ƈ�_al�y������g2�m(�z\{�����3(h�
m:`d)1R{w���]DXR�h��tۮBV���[}���� �
�;�ި��r�R���3����(��0F�o��E����ˀ��Oԕ�F�dP����'4�R&�~;�.��e�(2F$�Y�!�%�R�?��M�[�- V�r!�m�qтGCb�4c��>i�Χ�A��&�1g�@h,Ȁֈ\��C��_H���U�MG�����P�]��N~�I�[����n��]1��j��(T�Q&3�������d����}/���`d'��բ�Pt*b��ݓ���EM�J֬�n�p$[����W�!��ߡ�/�G����񢒞 [�xɩ�[��������h��c�`4�9O
M�\kyD�0.���Wd�Ga)�M�9�y���6��{��!B��ɑy���R*dt�߰���
K��pG�Ӣߗ�҃�ͬ�il[o���"洉�ee�*_�()���z�����t�7� �__G2�4�/mՖ�1�W�Vb���C���L�]H��z5bK�6�f����g��쏉�Ta�aT�ƂJ�� o���3͊{|�['�č+m%.j�H[cCp�L���f�h�%*�߻"\s�]��2�o��1'�� �~�g����������B�VY�6ئxY�0c��>Kn����F�hE���Z�Z�{t��T�-I�dR��mZ��Y:M�P�'����Gd6N��Lr�/�q�c�<) �2���UӮ{L�� ��]���k.R����o�v14�_)S{�P���<`_�� n����A����6Z� ���/��C+5��_�����E��,�.h���i=����4�{�]��κrI �u��w�/R�Rr2�۫,��N9�4�l%��ݒ��"��,�K���x���ʾ�- �]`p�3@uu��O�6�;6Y���&w�S��m3	l��e`Kh}ڲ�}�:ʅ�+����e�S�y����4���o	DטVqj�G@�R;֨t&Pܯ�IE�L�ht/�k����J=�>1�pf��/e��{ Έu��2r_�(V\Ǔ�!V���~�|8�j63R���u�7�;V엛]e̶ؐ3<��;2Z�۲�Ů�� ���NQ���9��{�'��s���.��X�b��l��Ař�e����a�U��`��ܒ0�;��%]�2��y8�'�����I�Þ���	��Ȃ�l��h$��$o�	�x�4bՏ���8�ȋg̩��z���ZQ��:�C�X��l�9�O�J���
���j�ז�<,e��%���V�o�>`�ZY6w��� \9û�U<fi�7D�\e�!J�7Jy֣��W��E�9/�4��W�,�GT�yr�#|[�ɔ yT������L���T�f�r����FZ��:R���W�g�ϨQ�[�z�7��]�"��-��A�F �f�'�x�Ho��C{�Ob8�a���K
����|�oڶ	�가\�CN�|		�v�H"Q?3}�&c����Wu\V�p_9��(t��d��T�J���v�
��>/A��������eet9�J,n�٢�c�7�@��"=V*�,w���~��-�)�
�� ��gL�d��9L�#8�?7iљa�&f�]!�}�kئ��˟T]ņ������6�7�����+763ϑ��t�90>����sV'��ūn|�4���)I��%��I�Q�2�'��Â�������ZP �o�Х#g��R�|m��p�n�"�B|����;+��m�MrY��*�9i�ٓ߁>��C5����Ϋ��ƾ���R���,Y��9�I�v�+E���k�?n��gs��Y�[Ԁ��A\ 4�YJ��Bf�lF��d�����/�U�M���;`��a=�Ǉ<�e�s�.���?��H2�(��&��F�c(��;�LH�������~jk�O.����fX�<�sً��CJ���?�t�o�M���Ac���J�DZ�{u�z<[o!��?X�My�o?ID�zY��/do�Bw@�� sx��.cRJ����Ȗ�c�7�
��2u�Wɕכa4��G��A���Ao�`Y�m]�-�b���9+\g-��� ��n
���C�N<�C��`4��|׷���"���ߐ7��� �1V��t��]��͙��{�)�i�Q9�p���F�l�$�(E��C`����6p���Wu�ș�6ۿ���H�a�
M��[�SK�$�(�GG|��v ��K��ywL��/���r�j#���h�+0����,yLOZ� �ҍ�Op�Ã�;�ǀ��g�;O����Zۨ�i���>wޛo;U��kr�]��v�#PT��o`XH����d��g&$��9�(�0NG�aQ�3�M�����; S�&����e|��Z8��S��6WLt���f�k�\d���FC�PV[����bY�@�i�,��ulsG�Z�q��BDj�pRilZ����Ml�V|)�Q .
�e$І�mW��ra�L����V��o��&h�����g}��Sہ0��;r+~կy�Q���^�y�2q�7�j�#����?X��pr��Hu�ы�#dr�JM���B׎i}�:�_�4�o���egl$�3��8���Z�����!�a����(�! �؊z	���轳��#I�~>�G�C��A�~����R��~��.:;w��U��t���`��Z	�杵�#,V�b��igy
�Nt�g�m�d�B�AOȊ�c<=z��:=B/~���`>�J���!��WQ�P�*��&�M&ݏ���k�f��>�eٙd�U��&Y-r��Kb��F�_��{�벵P�yG� Q��X�j��/������i��L�;ȿU�U�?�G]o�_���t�����~����#?g< �R�dQ�w�����Q����w��43˔���i.�Re��=�[��T��d(������U�\m��g��m����t�><m�31-��J�t����ː��t1�ހ$�n�ѿ���%/_�H|tow��V��^״&E�M��`-m�!���q��7��%�JOB�E�t0�U�ZT������������{�!������`�\�3��p7rR��;<k����KS��� c��	��ܴ���СFr��'ԓ'����IH�����-�Z,��h�;�3�֞�]ˉ;�TTsi$�tbXD��5be7:�cds�u(3�5qW�����:�.1�8����0�"�rC `�h�=���@R��Ko5q<�gKQ`J��A���%�<W��Y[���Bώ����b�(.Ԁ���-��v�6�z"�m@uj�r�a`�e������s is��w���e�?n2k��s�z���ּ�56�۔b�1T��f���� �gB��_TM(VL�N&��I	w� x����7<��	ϞnT�}�`T��%"���g�螢n��'m�j���q��Ad,��0��#WeA�
T �*y`x���k*�k���D�����2.b@e�~����i�K�M�X4�6tߔ�1-�ᑢ�������u��b>}��4��٧⪝���������@D�y��/V�e�j�u&������t#��\��g��
���"��A�_��<�oA���s�D-��G:�2Mmܟ���Z?�=��W��c;�粢���
���Jt��/��F�� ��4K�����<�����N\tr��@��k�Ig��ҍ�t,.���MÌ�7�7��	v:��EϽ�W(7�T3��[6U�/z"���\H˭⣉���	�m��mJ�;��Ϳ'�Z��-���XZؐBuF_���8>e5��!�y��;�LV��qS}�e��N%�v��e�|�PF�����ǈ��V{�S޲�J��;����d"%��,��ᳰJ((�5g�ԁ1��O����̭-&����HA���+�4͓�r';%��7���������if��|�\E���Mx��Sd�ė�o�)5W��7u�" �w�w��A�u��Y���#�O�n:rP�d�a�n�g?�
b���q���Ų���[C�o�!��J�%���h�j�S8�#����--�֣�]}�8�1�3�0�����^��3�+���w�+�i/��8`���_���Z?��5?Iha�3#aTLt�M�G���^a{|p���^0.���K^����Y����c�l�û��q��To߯��?��q �h*���!Nn��)��I����t�77�Sq���D&��mܧ6s�-����
��͟�% 9X�=��4k�|T5�$�H�P��d��)��6��1���6���E�[vB��<YK��<��n�B�<�䩿�7��	f�񎷭;��#�s�d������ee�n�"E}q�栟�8�)�E�x�[	������P�}�#��܀����z[a!H��)PF�����c��UYOpn�� Ņ���\��7�෱��S�Kz��*k3f�����0f�5�쉊�� ,H#h��j�2��9�P����VY�pK1�G<��N�G9�<F�e�ռ��z+c�����z�vsD�8��9Q�<��g��nی���w�p�q����-��n�G��-�_+/D�������(�	��9��-�M_X"�?������N<&�>s����;nL��2�A��#��B�J���������/l���%ׇ�K�T�g�Rʞ{��9M-��-�SG�W�XP�pF���L~4��_4�z�REX(ҹ�K(%Q����i���3ͺ�5���M��9�D�������+�T��,��[}f�7I�N�\	y��>�z����}�a��n����}�'X`��jn����~r�F.^���Б.��|c����3<��
��v�;�����ær��1ctf�W̶��kz�B�����{%�j�B���o"��'��n��>D�*���4M￱ ���(s{eث��-^�3�c��6Uz�N���z�5F�w�b��Y9)l9/Q���'����1l'�>��PaN�V�oh6�͍�-r]X-�a|YO	'��-��� ��1�(��J�E
Bjմ���h!���+�]��B���8�ZSj�^{Y�x�G�j�zY���S��:��G%-�v�(�����P21Tz^�(�(^W�s8��A�[GSy�e�h�*(-�X��21(�2�,%��Q3������8��i��p�aTȸE�7��W�W��Z���.����|�21v?���<���@�%�&f_�˞�b��زx>��)[!�p?�'7���F ��E��v~C�*��膿�������'�� �ve����m0����	�D���{D<��X9�����1��ޞ$We����=t�_L%�A[s$�3�4HL�����()�^��٘@���J)*.��e�	�����0^u4`3Ad+n�I���KG��I�6����(�A� .
���*u��,}��A�e���YOf�b^�
Gt�����`�*I��0��]f�k���������b��锄�&����������. ���ڒ=���؜��Έ<D>�Թ�pV	��%�}Ng)-]0�F�r�u(�a�C-�ΰ���*@��}��v����.�
��Ȩ��=��<+�
��Wu�I��@�b`	�)�.�o�ڹFDx�2iK�f�K槷�Y%n�)�׮�I���{䤿j߄ϲ����N7��vb�D�3#�.`�ɦ��˾�ۤ���H�~�E
B�MF���;st��H6yXo�ڋ�&hW�pK����2UqRj.�e�ϧ�x��J0����S�5�6_C20�y06�"�
�1�t�4�g�bK�s�ʽ����.�+����o|�Q�w��އ��$��ΝU�o-�܈�T��f ��'����Pa�RY�jI�om��#����s5z�O^�X���Pjg�E^�?�o����=�8&v��#�<��K[�al�(^��3W\"�$�T��O��b��v�*8Α`�@��^^�MN�tG"���4��>�;��@�+t��ɸ��0!MK���`WZ���B�Ŏ�|C��m�̨9�!�Q�Q3���"�*
�:�ǀ�>E�^wMy��:��dVҞh1�D��Au���,F�2�ۻ�o�BT�x��#�	4W�y@�2�#��Ά``c�%�/^Ͱ��"��e�Ub�2T	b�����;��܊�����?kLD|���2�f7W�������4�S6/d������� ��1yu����Q�q�|�Z�h����EV�.��B�X�龟7�<];�� |����M���xbaw����S�.����f2A�S�3�^�]����swUۓ��0�礧��a#"��A*c;��I�"+u9�i����V͗{�/~���6�FH�.{�'2��Ӝ���z`�>D[5>��ގ/(B�?`-��E���?�?�
i��������0b}C��(�-�WFmW�����"���� ��oSbZ^�"���D���X��h��Z�#p��~����y��j��d\�c,��V�=X?�� ����ME�G���]XE�O=U�-��䖙�;]^��i/��ȁ0�ψ����$I�����>h�f�za��]�Q�]bd�X���z/l�ͳ�b�H7�� )X�7�����2���8� A�Jceg.N�m:���,�m�Y,�uˁ���L����%�Tf�?k%��J�Ǻ��oC��l:�[��@�(�mV!U�Bz,����=x��a g��d�[oB1s7�=d�gf
1!t=�T�Dbx�[�Ol�����a�_X�0� 1��Fao��<F&�T���Sۇ&Y5w�yHI��u+�;QE�A�_���^9|��nR��u��"<�l�>z�l�U��l[FH'ЉH�3�=z��SWďZ�!�2>��fj����P5��<j�P��W���To���H�0����G|02�[�H(�ǂ�#z�o�u�5��*�\��w�c�sE%�ma�u'n���R��	!琭۽�����aDvs>���:��)z��0=6�M�����s�$�\CY�~O!T_^��h�Sl��-�����x��ɰm\%őf�fO����C>�\��g��[�Z�掣<�h=e�H�/����W�>��b.y�z�H?~Y��TN�J���
��4�n�P�Y�^K��|rNT�z�zb���-�/�Ϯ����i��  9fk3���6���k�J�`V�e\�\d�e�������r�ؤ�fH���_Vg�G�`�9�)s��Kݵw8���U$�k9�k���i��Ԑ�J(�f���*�~Ϳ̀��|,.�Fg!/�Ҫ�t�_�����'�`gur7�J�N�"��U˱	S��P�ʊ��:�A��#���{���On��2���]0'�Se�,��?B��j��{A�L��VU��<�"R�N1İ��w�0�on�O��R�3�A'Q6��XD�	T�_�&�b�ؘv�(����A�U�
~%-*�yʕ,-�v�w��r�+�D~6`� [�$9�>��Q#��&Eg��W!6�V׉���u-����]����x���%YO,�u)L�u���ǅ+��m9�.���=q�,�&⫭+�c�ļ8�G�\�1��ָ��u�D�]ދ�jT�о�o��Q'���L:�{2�j�X4]��	�,�[��y{�i0�����M��ړU�.����q�a*�*H���aCL;8�@`!}��}� j�G�u� +T;���U��{Z\^cO)�n��:�ň�I�_ � �Yb뷢o�u,U�Ja�B@���ʺ)6�&[ I_�c��yN*��jhʢP'Ia4��sh��2}7O$9q+C��[��  P�ܤ�;����lYYx@+"����F����+_�3[���ߙKX��;LC皴�FIp���6q#j���꺬�Q�s��"yQ�z�h{;߫N7��T�DN��)]i�:NI��b��e�1w=A=�i��Q-�b�*;w:�-�"�O/�Y/SꟚ-Y>�yݦ����ŖƄ�#0;ܺ}'�"�/jBN؋Gb�u��L�;�P%"T��m*@���[�~(���S�,9�e��$�g�5�S�%)!W(��!3![����hs�Ɇo"p���_:(+s��7�	�∾P�Vf�Ѱ>]��4L!m���Y8x�j���]���)x��р��:/i��(<�ʩ�L?t�v a�/��;*>���V��YO~	�	�����d����_��o����,���C��t�:����Z�8�)�{�@p�sh��Kq�.�/ܯ�]1�����7V�ӵ��	���+��H��2�J�%ٸ�5������`6����m%��F��
$��x��{�é�P"{�'�,2��R�u�P r��ùg=v�Z���9� �,��[Z�T")i��t�-�R��Ós��3E8�a�@m��3���% ���7_�+x�+�+ez��s�s7)ܱ�<b�hG�[�d�N�GhР�� Z�{-�ۆ&��qJ�(��,�q|�$��D����u�F�-�z���b�	�����v�nq�@��d�x-�=��{��,�i������uլr�˨�ʱ��r\��ZPc������;�v����ٱ vϥ}����:���*��F	�����c�F���i���K�x6kP���$Z8ɗ����e�o�5a�f�=�抻��}�lrz���*-�̸�I��X8H'd7�a�����BNV���༭������,7Ѝ��1�k�ϼm{'EN���.������3$Q�c��� i���c����d�i
B�@�X�I�f(=����֧��Sz�^�0�Lޜ]&��A���W�fe�ܷ���$��eY�[�f��Ǣ�	Q��+��iK`����$�1�=�:9Ȓm��{��7,��/��f����H�ڌbh��7Cb�J|��[V�Ymr��śBt�+�l,g��~;�S~v }'�W"����׉�꿊��0�{��l���"����[��������S
JID;;�{x����(�>% RJS��Y��KO���?��t�A$n.�;��O�����i��n�Lc5$��T�\�p�3�{�D�Q�J5#�K�S<hH�Ю���ԥ��!Bc�Ɩ�;K�߈��G4�����*���x�2�T�X �><5���\�I$�D��~aI��n��9��qfX�V�3�]qMG~$��-�ܔ��
r�|�P̣q�Ik�:�w~J-Z�d����^؍���/sJ�/�.��2~r/��s0��V�5��e���4�nx��� �t��/ �ԼN�׼W,�ή�o�q��K�4�@���x��4�p��T'��j)K|�	�M�8tA�	y�����fH?����C	X�~�Y��p�ް�rSI̹x5�i�e��%|$�.o�"�N��F���<�Pp�`�H$�}�~*<K�Z���GXޣ��i�ʊ���狒��KL ����P&�)	���Mو�:�F�[�\I���	�K����_���m^P<G����H�nlY�(�?+}t;m)@�4.��TRD?l�n�5� A��r�a�jN@��! ����4W}(�ۥ�("Z��jמsuc�%�; �c�9n�6Rs�B!s�>�	���lz���6��AŒ�l:S�O@t����G�`Q#".Yr���H�����j��r�=���a����n-A����oP����<��[j����9t�He`ZV�!8-
�J\q7bB��-ʮ}��gW4ܴ�Ė��ƣ�������wso���m5���QQQ�z�&1�nK[cz<�������;�^��(6_b�؁x)�Y����R���+R�ї�<��nK"a�w$�SQ�X��3ŏɀ�o�q���>��*uk+�H�6Tm���/y��P��	_1j5�NB2�@8M��v�k뇦=��E-��i�d��u�KY�0g����DV�!��m�X�;�$W,�2�J��f�i�RJK]3�	�Ɲ�g�GC�4ٖ4�LÚ��,(I�Y����B�� �^��m����v���`%<�����%���>)�Y��lP��\F�AuE�}��40����R�k�թ�.�n��&K����;����Q�+=y�[A��j�({d�|_�P��4pv2!z�(�/�*tX9��!m�ߵ �V�M�̗-;`(֖�f�oRn���HwO��.�D�����,��r�Ta���U4hd9��j�O��8 ��������p]X�`}�f��s������<8q㪧ݶ���+2�*���ݫ��!�6��X�X��m�X��U
Ц�$��?�Fo}��� �ka�`�J|��QxF:v��ںw��hx�9��GK���2ş�]���ߢ�����2+��0#�,^ ���r��i���g��t
�茞qI�YEl�bĶ�)���H�{N5q"+�rC���<�]=0��	�p$]��%v5]@d�{y�ï�+�l"bA%��������8�� 48�~�8�>#��<+z�xA*ހ��Q���Ǆ����+D �s"����u�Fo2�Sˣ��ѝ��Yuy1�d�+!$D��pO�9�P�@��}��hNy�`P����q��!������,����K"T�
W4-��͕*c�%���t^��V��q^_�'L�3u���w::�� (=!O��I�<�Iqc.��*�o�4��e�C�k;�|�>z�H��8�%̯������:0"���蓐TY�*6�&���6R���������1%�����4��0S�zX�]/-�f~2-��Lp��M�Eu���!�D�����	�Ӕ�v�J��K�򣜁P�%\��0Rz�-rnG0�.�e+>,����m�����ل�~����Ӧ�2�Z���KdH�9I>���9~+�9hWͅ�ղ"�
�;F��fH��3ʘ�,��cK� �#n�������Ú�]�]��0)��V%e%QT�K�o���7�I$�A�j{��8F��%����Eʒs��W�haᵘ�y��l]}�m_\�������g��ߴ�0zp�Nt���(��5�Y�~�C���F��4�ͧǞ�t�L|�(S��$w�H%��pI�4�7C$�E�jE�&����m���ǹ����T��u@B��F�fJ ��Z�@BlV��p��e�1��$o?Hɬb��x���Dy�<����U_��u�b\M��~E��NZ��_�l��AG~>yʝ��xXz�\���0TU�V�׈�W����~�U T��I��?!�ԥ)_��)�~	��NO�e������(��e��bB��2�ɉ0�"�b4,�����V�N�����Ql�Q��v�MP>��U\R+�E��M��So�DS��<�L�
Gjѽw�|��~�X6~����m|8�"=4�\f�}Ӥ)�.��M�<�� �ww��ra��po��7I�s�.J�4Q�h����xݏ������a���׾��w=�*���1��w��;s�:�g��1�@�!�Z�[X�:Y?7�F{j��c��8Gj�C3t�,�� F��M}tB��l�\6�욧��^ְ��+ӃڹN�t?t�s��ILlZy<Td5�����宋�t�����U�D7>�|�_N�z�d�"f�h�~VR>g�����M%7\_o
��t��
�T4a
z`�e|�G���9��]b1*������0�S��rS�m��΢���p�A�IT�U�L�y���Ow�6/��E�:Y<�%T���M�§~lܬ�O�D�������G5!�,�ffr0������N����Vw� ��`���z=Ћ��5qU?����6�H����K������f#˸�TkkzY��
>2;E��A�@S�u������V�y�$Σ��f��Ƿ>��wb"���VqZ����׏�A�븎� ���k�\�˸��_fx�FT�U�Ǔ��F) ��J�m�b}Q@)��]��$��D��h�@� :����$��a���#�������շ�@� ���J.3Q"�9T�]�R^tv�LȦA�?��B�1h��֡���CM�T-bBKA�k�8Ć�QɵM��� �֞�� u#�J^����:�;B�������:��ȼrI����eU��o�RJUȴ�K��a�4�Ve��"��Ej[A�>^��#<{�(��6�k�I��E����R�6EK{���)@���*��4=q�h�'W��eH�]U�����-8���i�AB����K|<t�X� �s��7�	׶�M��#�>>��Y�;�,�����!H]��Z�p�ͯ�p�boMS�C��$A ��Rm*5��-�:& m�P����[�	��l�)��h�o����?c��\�
�%S��E�jYی����E�nh�& �t�՝(�Aӓ��$�N-/�	*�z1�$e_� ��#��u@{M7��Ů6���u��F�h��vL���8]ZH�돺)2LX��G���,QQ�?��)-<J�����oO̰��Y�s�o,O�W�����c���ǉ���Y�8"6�s��X�P9eN�����2�a{5k(��;A^��b��j��ID���tJ�� ��V����&E�:������J�%�38¯p�"N�P�S�^���XBc[�z�0߶���[�LN�B Bi~e�����q�'�}Ɉ���\�s��,p����1I�q���̗���k�s�՚u@%�[mE��N|#7%�
ێ�-\��D�O��E�����k�G�"�G���vk�_]X��]�0����2����x�7.xbX�B
����~��+Q`�>��a�ii/���~��A j�F�G���':*U��Nz�n -��#����^ ��4��F�e��Hm[�Hb~?����l� ���o�?�>��ض��B��}s�O������SUw�H*��`���p *�
&��N�<-�5;��V'��u�0�ܠ�U'�������}Y���S4�a�e]#>t�Ͽ�7�PD��D�#�K�w���z>'t)�wf����瑽���|=�O9�K�jV�.�\b�R���f�5K3�};;U�6�]�]����u����Y�zZ�P�L��iZ��zh��@����=-$���%`���;�[��Ȝ0�,�}��~YH>�H
<�A�Yq��:����v�D	�4}8���%�8�My�������y����'S��B�C$�Z��\�Up��~`~�ώ��kgp���Ŵ�XG:���;�b�A3K��A-zF���e��0�e������	�߳Ae�=u`��n��b8z����z^*���-ڗ<NÄuށ�P;"���-��y1����V�U�p����{��w�<2���@�I[� �֫��l����4r �Z� ����Y'�VV�!AVY���9+��Ʊ���vM�%�c���+8�Ɛ���$R�i����+��3�+ �~��3���Ǒ��*E>%ՙ�TJ;˿p\ahh��/'% ��ࢥ¿��-���N��e�[i�;@�o`�-���=��Qn��m�j�5�ױ�9x-��y!�>A�y@�p$.L�@�z}s����@�Ν�`�J�{gì枣JH��K~����q��J�	 6����S�*RfBȩ���D%��U��Ƒ��>d�~�EU)����5&7}�3αL�.k��vBt�ġKD�޾��&F���/�I�P,��>S�i%Yؿs���i���	ȱ�/+n����]�lA	C�V�s?���Խ�+N8k؊��4W݊oE-U�s�D��$%�{�^"���Z�v&&�G���(��Pyg/�C��.����c��9�.��MHD�~�C,M!��՞��	뭺>|9�'��ו������@�Uu�_f���9RffВX�0cl[�9�Ӣ�b�
s{!?Yu�*��ɉ[�qa!s):�0�´�]��2)0.�D�n�&2�՞a����P�ٳ~F	I�K����_HK<�ۼkj�����X�v��p8��:'d��G�y�ܯ�ǑL���?c��h�g��}&�U����֬��~�?rzw{��gn�ۏj�S���SLPw|��@$�ճ�*D%>q������W�fޟ�	��GR�Ga�vaq&�"p���f'Oپoo7�x� H�%�����w-�r����u���z���<�A�@\�p�5�F�%������Ώ�T�0��_S�Zꗱ�0�r׉�8�&䷑O`����7S ����x�8S�3��]4��<c��1M�I�����X�����)��^+ົ�gTܺ���O�m݂�j���d�������{��P�e�����,3W�+Xw�a'\��Nla�/���^�	��T@�n>2�![ܻ0��K�K���C��k�W/�s^Ufi>[��a�<U��bv�'�!s�'��=�׌ϼD�ܬ��T����9�U� n�a�ǂzT��9`JPiy g�T�[��}�.�����k(�"�9��ZŨ��ˌ
�.�	���R	O�����S:�Mn)���M�BS��ע��kIT��9�{H��|�k��"�3?�՟>~Җ2i�-��d��(7�����
d�_�<
zO~Ct�к��L�Ah��{E���EANjb̶�q;%�A`�!�9�ȟ��_e<�s���uV㴻�@ T��Gɮ�P6ZI�Ҏ^�˚���U}���f�:��"�e�G�#Z�]ȡ�Y�'�S��U1'�&��펐ZM��Q$���G���q+�H4�+\�	&�>m =5��"*���I{Y9�t�?n���\���:�6򄈲���p�x�J1~~�lhc�G���X�c�ȷ/L���&�����P�w��k��������z�D��Y[�L�:tv�Y���1�͵
�ynms�i�����oN�]	r|@E?��Զ��6:��b#l��#s:c���M�ԕ���Ѳlm���M�Kݍ�l�mi����s/����^A$�uX�!Mnx����<(e�ҵ�Ų�"Kֺ.�PB�r=��3�R����!�܁�ᨶi }�#Y�yGk\�.���3��&�}:ș$F����ku���Y��O���2�2w�&�|�wɤ��'&��Q��:�R��Ƥ8+7&�]��(��� ��4��h�����M{�x�2�x>���{�X�\1�V��/e�>��e5�p�;��]x�捋aщ:o�nkk6O�}NjlR��_�,�E�/{�51��JaA��<�６wB��0��t��5	�_����� ��2L|���M+K�����^�=��\\��քľ}�y�֧$��D��8Q)�ҁ{��e��Zw*5w�E[�2,�w�.�>P]G��K@��� �'
m��U��eC�mCY�t�i�dL�/|��T��#��j1ۣ�!��aָ�$A悤���x�6)0�.��m6�jR c��/~.҇^���ݤ>6��S�9�O�N#���I���-@4�3�iu��Oj���6�g؇�֡w]I�c��J��
8�e6�e\��]���n�=������hJ�j���Y͉Q���w7�?9��#(�^���V��(�K�Ǚ����k�el��K��M��ɭN�%�-���7(�F\��,�g=����ܯ$��X��=��R)|,�<�w)'�H ����Q�t�-r]KU��~)�^]{�qt}����L)�}��s���o�6�U<d�0���""P��F������.�yc:(��)4�?�x���׺���U����Q`.j��Aʥ�p˕�j�<�s�OY��(��x�Qc���u�S�۰��A s��|_���9>uc${�7������Z��nQ�귊�������h�uG��$c���A-h������\y8(���op@z�V����t�?��5�ݙF����v��~�����N2��	"��տ-
�F�.�����e���|b!O�d<݈���M� �<����LE���T���@�6M@m�m[�K����W��hYv�hw�7�)�L��wӅ$�^��5L$�����?��;"��K� ~�w�Vt[���׿~Md��P�8m7��0> ����Z�fR�ag�i��_�U".DJ_;��MVq]��n@4DΌ������"����^��~0��<���~�q��X�y��`�n��Wr�Z��(<�>M��-\^�iƚ�E���+z�f��6����vᾊ&�c$Tf]t5�,Vd��"й�b���8�>�4ɼ� �����$:,RNV�	r�%욨�t*M:�=�6W���(�H��MA����9��AvW��;Dr>�c�Y��;��T��
�-P�L��s'��.� �?�����~IC�7ݠמ�gA��a�����>���R��F�T�VLQY�ܼ_�c�n��&m�渪a�������Bid�r�����gq=�ř$��d�g�f�ޫЕ� |J��A��\�i|Po���/��}����ȳ���sOS�X����pk:�u�$�?������s�p�t��w�]�Cu����-�ѷ�x��I��Sq�K�tc(�ͭ��r��~ӹa��n��q!��7Ԕ�+����鄖�$0Q�n�x@b��=���os���hH'͈Q|��C�!2j5A�^�(�O�;��2�M���Ӝ	�#s��H��+�Jl:�,�#�Lk�k�\�X%:����ڽ'��(4��z���T0x3oYoti3}HP3��t��(��1������oꭜ;|������b�A,�郦P�'��=Y�d6\�Ob6�G�d�Rr��ڦ��)���W$fԒ���P���zz�p�v$$gi���<�����W�K#�y�@��[R��eoM�����~β��h�ý\OĐA	S]��P�d�) �l�A e]�����}��^�HI�!l]��lS��K����0�|�a_��ky�_H�_�T�6+��x �aO��Jj�=�O�*����+�p����ɛeQ�f��e�A�l��>-�����=󍟴MA?`��4ԳN�����B����hQ������T"+���uO�1���eޒ�~W��u:[P��l�Ȓ��C��� }�DV+�7K!C��3�8R�Fp���#�g�1�/ ��</�߻���;+�\b9ǖ��? kɓ?��l�͠��/c�$�S��R�s��g�w��C>�Y#
��I���Jl�=_[��7yO�4��M|q%x�2�-� Y�WC�V7,�*�k�Nrc٠���g��"�Z�9P�VOm[�j�-~8�B����h�4-i��)	���r���\_��]m��k��`���G{&KZ(� `o��!��9�������V����Y��b0�e�yX�xä��!�Z*N[����/�pN�����a��~��զLl��X�H����wR�����?æ����!���`�>͈,�ߪ4�3��"Z���T����q����0���:p݆1$C)�]uU��VZ��t+��}�Ԓ}�U�U�Fx��� �寛 H�GvuTL6 �NX2D}�O����B����̦��09s����\��~pƐ�Vn��N_�P!���
6_L�Y9(����X}�] �(�����w�ۜ$�C@f-l��%��\:��Q��#�$ɷHo���X/��S��x�Z�b*7�� �u�#�}[�<�����DT�*L�;��BD�Cw��׫�s&ȹ����t������:q<��[��M ��U�D5[�
i&��z��Jcz�'r&�A�]~�M��Gϐ��!�,6| #�t]F2�Rh��?~��*
�B�����q�� �w �G�4�V�&]�>R�5x,�����ƛ�=��o-Z^��P�Q{�4�����4�P�OC���0Sx�ٍ,
E2^�
Q��t�z����~<���w���������,c<� ��I�}U��8�*h�!�uˢ�WG�G�-��i�����X���n$[�'�Q�삓V	;4#�0��'�D��؍�+�^!��ԁ�Y6@���������?\o��FF���v��8N��-���84��'3n�AY[l;�v}�̙W�
����&u�K��0�%v��1?��~C��2!����M�����)�`�^3��y��4;��5���Z��t9�1��N��o�x��|�,����yl��3�o��*�����7:b�:���R�ˍO&O��>�w�@��r�6s�S�0#KC�'�8{Q�ENנ
w����`ng���}�	�f�!kp����G����T��@#��6���������"}�8�oH������z�:U���ݟ�`�޶�g*�X0"s�-oYRW�G��նy`ⵏYվ�	[�VD+��\Մf�~|�~H�g��ض�H	��u6�T�O,�>X�h�r&�E�'�o�0�!- �u�(R�����q�[��F"��QX$�
�=c�BI��|����OP���Yx$Q�	�R<�UF�պ��
d����,�Cr��+���l��@��h�wׂ�q�0 p,���N��d��t_�j�Is���Y���s�_�j�;����25����HpLdM䧺�s३��"��LR�!^<��>�Y��J�Ʀ뎎r�����Bm��[��đ�y{"�S�"HsU��a�!0���g��l�.ə$"j��{f�\;7z!]u+�\��NG�k�j|j�C����K9�s��Ai���:[L�{���`f�� L�&p�,1C�۱Y&�npx�c�4��F4�=�B��/<u�K���2��OXz�&Â��������)�VQeSF�7Z�K��B���w����A�@��X|�)B���8oa�#�ŗ���@�c��e�{g|t�U���̖�����ڨ�xդ�����N�@��7w��E�����+�z��frp�5�fo��̢��K�����ġ�xG�ɺ	za$w1�ߖ "���B�Vr��`r��BW֭sry(b*@:eb,�W`
;��2H^�u|n\�c��,<j�xh!`�-i�ԣ�?0���d΄�5\�9"��W{z8&P#VUu����V��0�5��=�)	Ӫ��c�#�Պ/��Z�2�R�y�(v�OoMj'PKF�V�k!��]���>R�5��?��aY�w�wm���ĸ4 ���T�UU��m<���X�3Ow�@��X�HI��^Л���c[�՘к�1f������s"���I�a5Q~C�vU��͓�Ι����"O��t~퍲��a�+��Um��+��*iN�kY��7Q�9�u_��)�{b����@P15�~0<�%`DL��skZӸ�I�1���;�_k�]��wL �u����.W�2!#b���C�����i�P�5r��L5͚�/�?S��ICI�lдM���'[�2��2t�$.9�V�z#6�Lu�ѵX������ln�*���'�:[2?���H�F�k�@烈n��U��a�D�Zv��m��>LJ=�Y
��C�%�V~B�2H~nf��J|�:g�,�F�ڍUv=�D�Z�8��f"%��������3�`�D����'6��C$�E,��*����q�C�˳k��h r����Ԕ$�8*��xNG�..Q	>^��α[�?���%��u%-S���Gt&��������r4+�z��>��L?�Χ|�YpԆ'����B� �@�� p���'�
��汇�'�+�%�bJ&����tDK4��Ȃ����HK��N�)�O�@&D x\�B?�$�o3�,����?�d)�};q*��2ߺf�^��'�f�QpF�� �G�z HG�1Ga����W2E�������e��� �1�ʿS��U�VNL������'����7�ީN���ɍ^ Va�<U����.A�#���p� �}��	�T���9 ��P�g?(�XU�G���H�W�.���\ʈ,�a'��J��Pi�{��)�k佱�Ӿ��8k��Fj޼�W��������u��e��.g/�폑��%%o�I'4��T��U���
��ԏ⟀��8��i`�*Y�p����@��؛7!G��U��]^|�@�8���ԷPD��U]m*2Mw�r�\Rs��-������.�0k�3W\6�?�Y�(*2�_.yH��v.���p��)�MA��Ó�O-\�J�;���w�1��"���p d1����� `�����Q��!ܨ�z�W�y�;S~��.�	4�����
-At��s��fNC�6�'�8��/I'oՉ,�+�[� Xt';|ٰ�_�c��~/+�A�!��/���V]z�ě���75��X|(�@�7=�$"NSE�yMc�!�H�ͧ eF��o������%��Li������Ό���mtEVr��Ȟ��xZ�.��L��2�������C�Xb�G�l��I��>5�f27P����Hu�ױ�L�FaS �͔0�۬>�n����oR���0�|�F��$�Q:��[�d���s_ey#+�����|�P���4��э��Z��M,�b(�'�S�eè��.�a�$F��ڑ��?f�� �	o���d��\/���+Km&V6���xa	��,E�s3g�
���GsT~�0���W��f��	Vß?Bh�w���cvZf����C�S���/���[�U63��^_�im�)Qp<QQП���i�ˮ�do����݊�W]�'�g�p\�D�����f Nn�=����/OD��~e�a�<6"%�g�P��Q���d�Ӥ��+c��]HϩZlI$ऀ��TC�lb�s���r@1�JB�����Iy�,y�=.+B��r�c�ReH���g%��腖b>+�3�?<f���3|g�1�OjQΣ�Z�
N5���(3�� �� ,�ⷈTF�T��Wp��r��Q�����X�L�����A�:U���h~�����u12��IQ��;w� ��>�Zݺ�sy֭�]:Q��� m�e �����_x[ya��1����"_˘x=�"�䋿Z��ڔD�SB���;�B��,������vͶC-��9n��.�+Gw����	���ʦ�Z�{�}y,|i�B�}�v�a��K맃�%� �#Z0���\�cb�ً]������ltnV�U'�@�lИ�4�V��������(Y��}��g'��ѸiV����1�@�l���z5�-9i��q�W��j�B=x�;��\F/W��x�FЋ��x+E�{|���)���#}.�n�$�*�]�ҏ+�@ص7�ǕJu#8; w�6�[����2>���a���%��3��k��%E#�Qb`����Z� �b��v�\�f�%�ѡ2�ϓ6�t.�����`t�o?�]�����AG���>�^�� ��o����T�Xq�e��'��N�L�5�+��<G��ǣ����3I�t�HW(`6Z�m��!Y~c�V�HTK�k��W��%�+�Fczv���We#�f~���,ףo%p�]� ���l�.4�cw���J(D�2��Jt�W�o\����q],��6T��b?�8��A��D��3謧���	�`�� �ю�_��n8��r��*�-Z��4KQ�9%�6��mzO�/ �p'����M�\��Љ�E��9ְ��G�t�Rʀ����G!Wo��1c�	���g]�/�,��G���6A���D�O6��|�F;)"6�Y��Z��يQOCa/��ۉ6�A~�\�����^�ݫo��3y�%���+g8Ww�f)�J�����嵯�U�o�o�\q�9;�xTX�p�8��SFu�Y��F�?���	�k�0��J�Vs�F	'�	И8h�>���`��4���}=%���@C�-���v��q	x��O�g���̪�p����0YP�ù�s�W},`�&<͉����޿AҺT���t�<��k&\h��AUB_CG��7]G��b&�C<�ށe1���I����y�)_B�zy�ź�@�,����,��m��`V��[� !G��g(W�5ڦ1N�D=ɜD������@,/�E��y&��,�<c6ZBuQ����E���Z��,��(����G=k�a�Ș�A�a�2�8UH� (1��Y�.��2q���d���l-�k
�*���:&�r�)���s��:��2���gBＱn�6=�9�%1Jb�/{\�%=��3?��|i��&l(�EZ�hV����EH�qw�K��1�.�S�j�(!o�����S�ȤӔ�5,?�9]�����\G��"V��A.y/)�	���p���+fע���0�o�����)F�s�o+����Vاf��������/ʥ����e̒�G����p/>l�Ş�7һz��Q_�ᏹ̀F3�A��f�A�|����Ϛ��h;9�GYۄT�U<Dd�\�$���n��dDk�(2�Z����3L�/d����NH�qϒH��w*�h$�����e���r@�m��){�u�;���'��pW�����H�aZ<��f�)V���"?O��v1ڌ�C3��]�II�D*3u~��"#�J�@xj =F���G�P���gͭ`�p�SA�������� ����%��|�)3�G4���_;�˹�Ă��>4{�.���s 9b��_�uS/����N�z���g%t=J�զ2r)�����;&�!V�!a�v!\a�]�CW��l�� ��L�]�Z��Ӎ� B(�Y��w��v�<��o�L��K.w*d��C�!�/��y�6��1+i��4)%�^��蔚=V�|�.����}�8louz-�5��vjgĸF��*<�ǚ�T�20^�c'Q��i�r�؀(H/��� bD����-���F3����+�vPN�ւ��pG}�gR��#e�BV��$�d�N�D{.;�l���h���#���L�%N@�\7x�f!4*!*���4S��X�e����垺h��yjm�Q��r-%�n�(���Bf�I6�$w�ؐ�`��J�2��3�e���L\V]�G���Sz�O,��ຠۘv��BS�[m�M��xa3)� g�%k<��(�Q�7p�����R���8�@�A���
2�M(�ν{4��cpw	�M���ǎ2R�%�!=�+IȻ�tLζ<i7^0�:�\����Cd��u)K�M�y�[�筭S뗙!}�a!qM�[v�X�;�m$����^G��6���쥓�yf����<�#SZ�=E����`:*8T9X1a9��8�$�n�Y���`���-I ���҂ZK�=^��u8
R:�N����t����#�.�̩d��%?�r��-���o�5����Ók����t�4gC:'bE� �!-���U�����	��	\T9�:Waxa��^��>e��C��0 �] I�D����C�/\�T���8p,��ݾ�<\��xp.�6�W9'�
C��G�/[�p朎��*�P�_�`K�_lp�6��K�W�d���V;W`L����#�2�ױ+��6��l"�9�*�qޒB`ms�t�e:�`[^>ۀ	�9�^��������<*�MI�t�/�^�C�)����N-5q0o�B���s��J����!%u��nEK�v~,�ԧ�܅�K�f�~�r$&��oR.6�SI/��s_�NO�N��[aF7$Cp���~�jҼ'���r�$���(��q��DK�#J�U�����r�L�_�����0s��Z�'v��c�VRf'���/>����
�qtƲK�Z����%@��B�� �Zf��uy��k2ڿ�.X�T?~��LF#-~�{Lh����s sWi��6���]`��e^"f�B�:e0� �6��+p���q,,�٩����z@?M�[Vt�{H��x��ͻi�w⣘�>:��g���FS��ٹ �=��"$`����ڙ��ŗ��d-T,�b�ɩ���1��J!�zR-��]pK�����Gn�	�c�M-wy5�A2,����P5��!Br+ؾ^��#7���nq�5Ösk�3n�*��r��(j1N���/��j?� {��v�Ѩ����hŮPG�����*�\|0k��/)Ԑz�y�~�vO�џTִ̏Yֳ�ۓdB�4�����Dp@ �׀{'��$��*�8�cF1N����9��P�ak��A�x_��2\�"4�����vN<*iOd��+�Q��dì�).pI��۫�i�(
Qte�D{[6��^�(L�aBo����H��Mѫc'�����{�}�=+W�e�`�x��?��1�Cj�������k�G�h7���RYDӸ�Ŧ�v���>`U&��Y���*��k,9jE��� �Oa�*����#�x�Z�����=�4��<�o.5� �������O��b1���X� ��=S�h�a��H5�ħ6���F(�֊��F.SW���t�z����"�
�( ��kO�G]L0Qsx��
ʂdP�eנJ����N3v�WAwj�w���0�c� e��qs��˓pW�1(c�a��3I/hh��Ba<p[�������DRz�#3����i�×�E��:Ε����\���q/��G;�)�?� ���E1��q�ְ�*?�g���������e�{�Q)�[���@cF]�P\�����;�8J�����=؇����U��ԏ���M��*�X��ธ�YȬY���SX��b�E�}]�0œ��3�*0X*�L����q�%����?��O������&��?�=}��a.�b[�q�Z���ɜԈ������Vr�7G�����r!!X����?�������s��5N��7!8<z�N#��$k���rk�%GO�f�.�q=9�X"�'�x<}ԝ���<
ܨ�:�;�2-�Q���V�	�!� ��$���k=w��\������Oj�0G�d��Fh�:5U��0��T�[����[V]�ƶ'�#�yy�<�Q�t��˾�C:do��r�~���5Z7rJXM�D��k�6Seo��W���~�"!��� d ;Fp��*|*��u�-���\x��B�*9��ɝ�������K=��"�v%�Y�Pd ��,\�[fں3��ZEy�U�u>��'?�N���>�^�p�a����`T
�R.qV��W����T�4�L�_��:���C�8?�0Y�n%?�[1AX�'�P�=��%�1{�ʹ��]4?6`��R���88����-	��۟ˌ w��6E[!1��`?�������]�M���M)����P�.mf�����d����k�р	����x9�r�>�}�5�W���{5T�N1wkEN��	�l��b\9�y��(�z!*�l&>*�?�kN���<%H��n#�M]��%�_P��M�Ylݲ��~yJ�����BV�"�	�'Z�I�W:S�m���5��&/4G�	���^��Q5�j���xm�4���Z�Z0v�骏0�Q�kB�܊�U��[�9�R<�� j���9*3z]
.��/<FC�hq�]�y��ُ-"���	�}�h��>��joA���Q�84,�)3mSq�,�"a�ͼ!�C�@��w4�i��\�B'.d�|��A�ٹ�� ��ku�k�W?��)����L������ �鸣�m(��ܛ#-h�$<������J );Tx��~x߼(�Ｐ�I�v�{��*xP����
M$SwQ�xZĄ�g��f>��m{��p�/��+ˊ\�&wr��{�b��\>�'��2��.�@���#}�?�P瑣̨bXP���gE�1��2߭�8*v����GR׹��(�`��"2_8����D���I�ey<�[���;Ю}#L5@�@"a�2��,?RPS��=}C)�DI̅�ۡs����~��ŉ�����Χu�t������3G�b�� 5	X�����Ų!��9��[jn��&�-|�����`4����Q�&����������ēP�P[��,�o��$R��0&��;�G�1���b�i��
)�O|�C�*�,ƱП����}�׸��~���͝y��Qwp�!ƾHp�����On ��N���b�1��]�OT�t�C��O�b>C���.E~*�'��7��a6��Cң��]��6��]U��������<���q./�7⅕Q�#9'���|Y (=WX+�pq]�B�U���~;�U� 2��z� �]��^2��7&�v�/ؖ��<��0���ҭ{Ucu��g�+�Z(�GI��y35�����O��9k-ɇ�Z���2����OͰ���.X���TRBQw��ަ���-щ�ʴ����2X<�H��%��<�s�����D�x�s�+����'���*���Zo�WL�N���YoG��|����R�Ei.B���u�^eв<�w��g���3�2C�mS��)��撢��l�Y㇆W������)�N��z�}x�˱�~���uR�7	����S?LZM��� 2w��7mD0A���]��ۮ鏇6Uq���<�:�ĉO�7�0���]F���!�����{BҾ��E����%����R��A���J�O5bV�Rp�]��R�rF���F��pD�k^�)��ٳ���_\����P�����`2�NreM*����+���LZ#�H;�M�W���M�w��%�˟�Q���&�e?ea{ly��܎���Y&w<B,���d'����燣)Y�;V{F�,煙���)�]x9)Ne���x0�����������=�į
��V�I��gϚ�fO�n�ٺ��P;���|X���п₥XT�L��O��������TۏK���}y)���~ź�Z��'��'AXǆ�x���EP�F���K�K��p͞�&�bd�X
O}�K����CV��JLrzp���ꑈ�߁�������s�C���T�fV:���N���
���a��l.�:�F�{����b�:\��!�����{W�%�q(:��NT6*�F@����/10�B4b�e���Z'J����8ݏV���' |j����B@�k(���l�%jS�wˡg
J%)��B:�;s�V"&�"��jt#0I���,M��Pn�d9����T����Q2�9�����j��?��^[T�{y�ˤp)c�9e0��0'�ɺ�K,N�y��u+��x�Y�Hs�L",�ewl�.Y�G;�EZ3>)�z@EՋ�:|i��'7���0���D�Gk4}��(OsJ�J��S�<���Ą�_��wҙLn����ۭMݰ�򥧮��J�{"k <Y$Y��Ȧ���`��7�b8V!�{�O��	!чL0��꧑�=��k����y>п\?4B\*���;��Z���o^a�{��:]�*�\?��Џ2{PC��^:��ɀY����V=�c!1�C(;h��mbt�z�礈�[���x�~#śn���)ꗞ�_�1����%h�%��r'-���F�������Cӈ��'��2Nݙ��)'1Og�u��B�k[��;�j��вi�6��'sK���o��u�n���;L(�ֶ��"n�_�4W�c����]���T���_J�m����^?|��#V�%WjR�ȻG;�L&h��ݿ�d�>����gs�D���RS,�T*s��%�H��e��K]tzS7~�O���nz�{*�T�w��3��)ܗJ��l?�Bֹ<i�5�`��?\Zѧ6�b���:[xPʔ�Ʌ�C��wF�����D�ܳ"_Vعr��L$n�GWTI;�N�� es? ��mG���S�~��^��_�PΆK�f�a�+�E���uz��,�E�����PX��5��b�W˴!�~�#�����J� ��T�u ʊ93Ɂ���A�S41�lcèLw��024�{�ׄ��@���h��躳�LOX�#;&;�x�RgS e-f����X����aYr��O�G7�����>����O.�S�L_.�^�����N���]���9p�QyT�M���������	liN��'`Ng<�J�H������W�u��4�t�
����e�2~�j,јOǹ�TXZ�)�Q�Pt���+o�:�!�81oY�輵�y�
mD��:���L�_7 X��n4���)Z��Z��lJ`��:"r6V�@�7:<ۉ����Dm*`.ѽ�h��N������;�yZP~�B���5O#��t����m�  ���,剄����M�w����H:m�?6���I��lvU��Im-������+���9���@�sF��J��F�;H���G�)&h 4��ͫ�yp�V-DjgY5�w�3�����v�L�N�2vͭ*�eþ�=H��S�^Օ���g�Bщ%��ΈG�&�z�mWC4J�5l6��c
�0W�hP	�!�m��ײzX���蔋�)�x�7W��l?3r�Pr?��	�Ա�R�;��K7�F9���+I�m�vx�LNMo|�f�鲌8� �:����X��)�G����/��D�#����r)�(X������1`'J����"7��R�����.�lC8�{!b����� ?{��t�9x%F�.B�������,�h�{�N��^��U��8��V���HG��Ci�_R����@<����S?W�[�b���qd��j!�t��d���������p������� e�Cu��x��+�/�3�aע���\o�cX���9���5�F6rgW��@H"`���W�eK.�˵��"/�i2�~pXΥ���������w���땶NZ>��i�s3t�(5�-8�a+�U̧�*d�?w�1��m����Wx��~XL�����n�j�+���E���	�[�y&�"��x��M_��%�#5������^m���]�����[�m���-3!:z�Fk�o�E�jU���W�7�#�[z����D`\M��w��a��ɱN��u	;a�F.k��"h>����(m��Nd��;�X�y�Ճ�P,|�|�(���醲��L��� w7��d�ׁ�,u�-��{u�3D�\Y�#av�-��&7N�?m`�P���[%��?�WQ�<i�jf�VL|a΁GS��K�o{�t�"������A��-�>�f�eҀ�>ǲA����a>3*w���9Y�,M;�L�_Ւ������p��FY��C��|�=�<�3wN�)g� �8�Ӆ��V[+q��Eךa�/g3BPF��\�et��*)�8�;#	Qm^b+$t��k]4PE�������*�:�X�9i8ó?�B���6���@1ë���[��!}��`+by�!�:/�i 5���I��7j	�t���E�7�����l̤l&��Y2���r���AsRD��<�}�է�nNse�"+���g�a��T1���p�M�y;�����~ �+%�h�<��e�ƒʀ�:Q.([�B�,VC�j�V=�F���N� �R|��]�d��m¡ٝ��֓������&����^��D���ͻ�5 ���A�_:L���ɥ�Ʃ���T�T�7�Xp�> �2�J@�oN����M��W$���q�|1+< U���[�	o�{�z+1�XHel%p�.�@O������o�R G�S4�v؊����L���:7r_��"���/���8����z1/����S���&N�-�t���Zmف��ק)C���P������B2Ι �28�� c"S5`�f���>ʏ$�JxW2�v��!H��s�<��+�e�gz�x���p�
�ߋ\�5�s�4%�z�λ[p�E��Q\�=��7jLY�kk����1Uj�}�~�a|�ф���h�j��Q�y��<L"4Й��Jx1�b��D�ÏS����x��ߺ�O��K��S[�d�ui�aWh��q�c^���U�J6��x�7q��4����"7���J���M�33���F��4�p�G ��>%<FB7��S=X3��E�|�sy�s���h�=z��<0� �t�0�V��j3͑�jŞ�n��5PѤ��FS>�x��ݚ��;'��`�������Zj�c��g�P�Q#\��v9�T��N+��vsf�I��aj����O=�8���by�^�4-0u��T`� �e#Gq#w�zڄ����J�TX��je8LY��%Z{��@L�f�:���Ԍ{)��`B��T�O������U*�W|�{�
�x^��2�:=�=K���Qύ�?R2�3����n0;vX�)���x��dJqՍ����=�p�ָ�4�oAu�hŷ�5PSJ>7�fS %���$/ŵ��sR�e� ,�5Ĭ��nzp�$��ٖ�rZ���(�u������O�_�~��mR(Y7��H�;R��q�k��-�[̘5�t6����g%b=8������08)�ɥ~Sf��%��{�7ퟬ۞���:��a�.�p�K��pFbڡ��H-�%a�^����(���੩����[���}�!�l�q!��#�C\��� 2�f-�����C��+U)*k+�Ef�o� }zY��)Az�eӆ�s�V!W���i���F���t$��>������
2\�y&�-G�}9�"Lƞ�VS��/m#˜w3q��YhY�d̬�=?+����O�����^B�_3N��fU��V�HYѷ��m;��Cv���uv�l}�-�)���*8õF� ^l�l���$E�����H�_�����<������ӣ䎶��In����#���]Q�d6X�5����2v:2
���ޑtk�V�n]�5ؽ�Qg&{��$?�8�b���l�����kI�X�j�G{*��.���;n�{�=W���$O��0?���9�ӄq���n[WO������].���]AW`9�ܪp5���1�TY��,p�q���K�������(S�֏���ǭ`\dDP}+�8�ie��*x�&B|��瑸J���If_?c������K��ZM�����e��n1������h*=�H���3��M����hչ´�#ݽ�a�R�Ag�/�5x�=��Ȯ�x�J�hT�T�M�I�D��U����f�۵V�hOV95	r�M�(�T������?���]	��<Kqsb�v�vèX����@8�2���V#.-�^x��1��?tM�L���;T�i7��T��_����8#�2�����AWa�	�Vf�3^ l�v\�N"/���yX�����X=sn���X����a��X$Z�[b|�պ��6���)g.��q�\�o�"���W
�t��_��Z���n�����w�����7��3ʺ_�?X�㜼pPB�\�7����'L�J��hԲ�i�$��&ONu�ȅ�LWO��頾HʚX�oK��tB��D�ĳ���~̼|��	�(L��1
������6�kǗ��{�K�RB���f��^�$�w`_�WU;:�=KBpJG���b_^9\����NU�`f����g�ɁY�T���kO��Ve�"��0r���[v���N�_8�N���ئIj+]N'�6� ��L��Z�F����sA�Oa�W�
Q�h2�>��R ��\(�<)Q�4��鎅w�M�|�̫ ?��+�i��Y�1{��0l�f+TT�̴sXg�F-�7H0��X���F�e��0�m�]���W�h3����7��Qx������

B���W�b�;L?'�@��Z����R�[��~���p	��`U��Q��둾����c�bK{F(�֋#b{��nH5y&Y�ᴩ:��Ҧ��[���<*rp��4�=#>�;&����_u��܈lX����b�����t�`&D�.~T8Ar�VH���g ���QD��n�{�I#�FXiC�O�9k�p~.����<|췹�b# �e�m!|�:;\Pm�/�?S���դ8�z������J�9����w%B���J��T�>�$��՗ˮ纼��3x�ѡ��XJ�|j2[I�b�t����|�OW���sWM�����D�c��}d.�4dɓ�q���y���E�1t��&�n���g6 h2��ސ�L�ز$��]9���%�zn��!y�qҜu��	��vffh���ĉ�wD�7��̿qj��@��z�_�z�r DT�)��BE<b����߃�t�d�贃�@(�
.]K��zV�}v���DR:�I�PG����T��l&L��?bc�����������jh�=����9բ���hp��)6v�g¿��z��uSx���Ŵ=:���!���c�}��E�b7�Q� �GӖ�e��$z�a��34N�H��z��°h,,@��`�%#�����޸~�ql�"��#��S�Du���H��r�9�Т���ު���6�׶�u7�a@K�����#b\\G�p�#n>��I�RU�K�"�:�9o%~C���e���a��Iۛ���b�_�h��D�9JC�Q�=L\4�<���@��cT]J�Ak4�޹xW���/|�6w��.j`�o�`�_^�< �G�R����fy�=:�i�����C��+MF����i�/�ɤ�v{��g��)
z6pJ47�e�R������b~��$�I�YZ6�E��6!��#��DK1+>�ͩ:��eb�4&N>�'�v���M"��BT�0����P6L�J33�m1����/	FY,�K0R�n9œ�a�&�6�<��N`(8xv��X�JSv2�Lz�i�54J�ʙ���d�6�IL՟��dhʕ]v�^���
H�4�r7܏]�y/JdǇ ��]=��H���/�$�q9��&@��Z�SB�dX�:��L�k/�-���8���M��}��@Ն�l���.�4�fi���b�6y�7YN�9����:뚱�+���vڅ��5{�t���a�Х��I����_��Xr��%���v�C=]х��ԙ�3L�H"d�/��t��1��H~��x�����P���B4��'K��q���9�m���g�u�](J?�F�U����Sv�����E;��D֙�O���U�v|rV/�(e3����n�5�D�P�B�쏛��dI�q��]dRM�Fl�C��Ip�������X4��R1WoX|��;)��/v������_�]W����0��B���C��&��B����L��k�K��z	L�=f���N{,ۣޟb
���y�4N��u��s{V	}���h ��4:��c3����b�u-����Mpt���n�!�{������6n�N  ��/#�� к�u�ǋ�c�}�<E��ʴ_2_x���:p�������yA���T�u����i]ƒ��-zJ*9���o>�O����\��N��>��:힑�	��A����ӗ�Ĩ�zl�]:B�:o�J����^E���C��*2h�����E���N\�߷��l�t:���[
���I���p���f�&>c���I�~����?��Y uՖ����H��Z��֥�ݓoI*�dJɑ,��c�*3Y���:,���Y���Ƚ���ۙ�=<_-|�c�{�����u�/pQU$�΀cq����%bk�"�~��'�)H�'=�m�izft��-;Ȗ����\$⩟"�g?U���Qg��i�*|�BNȽ��wШ�?������HAe�C��=l���[+�M�2�q�x��A�� IG!t���a�`���q��#�1�+Uļ�:�Y�6�Ҿ��`Eu�$����"7&=�Gpn*�]?2�Y���zp\��%�J�20����t1S"�s,�*Aէ��<��G]M��AB�@�k�$mI<L�j��M�u�1{���+7\�2�9R4i�Jh���T�ߌ�M��"�jc��Y[�7s�<�r8�o��w��'���W)}=ӽ?�ӎ��?	��<`8�^[~h*�Gm�E�D#�:��0�*'tR�:SY#ֽq�Z^���_½4ٳdh��q�s�� 0 ����' ��E�N��=�$�3V�e܍��%cfz�#�J����>Lǣ*�l���=M�#o�%�������ZP���<�f<��"� ,�i�o�u[5@��{m�9p�.���RV{�~)ؠ�	lIeu$�B?0FJ����ط��Y���+��ø凲��4�o�M�D7(E���5��w�.稍��9)n�"��I������PKXq�e��� K�=w}\^�jo<���#.s���I(0r4����U1��kq@�d�����nC�M�g6Y�����G
���r�q��qԃq,(	�6�8������F��/��!q�FS�x��e�#n�O){�d�5�M�Ui��͛O�$��ԗ��Ҕ"/�`N}N�Nz�0Zu�둬���C1FL�^~F�I�ך�d8HZݪ��{�;�w��'�Pg�JH՟�>_��N����FK�I?I����]��>K�I��+j8T���Wy��ܣ�̓��y:�S�=/IL�� t�2x���e��f��W����h��9Ɉ�%���59���X	\�s�̵�K�4�u�TaN�ކ�ʻ����g]h,mH2���>k��i�EF=��=0%�T/mIL�gu��j@��X2�{@�fl>��LX�gx�����|F����~<�#٤���(�ձ}�H����[�L���߃�]P8"<9x�JugE.��s5X ��\D�����2���ZڵG>���m� bZf�r�~=t#bI���� �qQ`=M��}��/�2� ��˚���U��ƥ��CsJ(��۸���"�W+���y�ߦG,P�~�1���e�zU��ۿYVϯA#l����5q���2������i��ZXH ���(EO�����n-/��< ��K���yR�Q�M���Z��^�v����JA)��@|��s	
3�p�r�V�(ʓOo޴Pn�Mk<��
�-	����v�s�`���� b�3�/Z3uF6��VT�@mo^Ypt�H@7t�'O�l�f�������F|
*��o�D3cH�I�
u֢bՀ�n?����E�Y��[��,،a)r{:�P�N[�ɈR�o1�5k�l���g�~�wO2�3%�����~K�Z��V~��i����I4��א ��b�s��P^�I������FMZV#���E7_� ��r��XD�˰!5�X�������������)ݕnZ�
�Y|������R�u@FYm�2�y�Q߲<�A�0�S%�a���G�C��O�c.��r�E���y^9���l �.P�n��1a���݁𪒺����Oɔ�'`�T+9�Y��Z���]&=*
����y �u�"�����G]�}��ىz�흏�,cn�$�?u�Y٢����Z�^������f�*���B�q��&�j����eO ���nbw.FB�n�/�� �Z�;Ϝ�3��2��w�c�9ݏh� $�u?BZ5C����)-�{Ĕk���|(m����6B4(�O��3��`c���43�;�� F��Ɋ�BO�<�LU)��-p��Ä���Oc줠�l�-q�ic��ץ�:0)Ë �rp����AP�Բ@��W�}yA�F㡃8}�`���y��A?n[Hܛ�C5u]��z�α�J�>�F�����:��7�d��"J���c�Sؐ�B�k�{>�/L���/�"�A
}⣧	9��
�F��O�2|8��I���[��][R�R�i <��Y5f����UW�3����W|�Gm�m\���=�z��S�~�w�e��{��s�I�H�& �ǣSq#��L�u>�Dg��lYh�mP&����_�n�7�ip�ݟ�h�em�櫵�K�_�e��-Če�w�~�+�۽�|�1F�_���pfU��E����>�axS��7��*k��k�A�?'i'j�T�u�~��Ȧ�d�MqG���%;H�s� �3�2H}���l_Ӳe{��c2y�o�aGz;1.�kF�z�~�|��D)k�D��S尾'I':�i����#MH_�ξ�С}?���Z���4��}�"�\`q�h���� �����\ȣ��M�����Fx��w �2�4�[ٌ��MA;���!��!�r�J'��o2���_L�ʝ6H����C6wC��8�Ny��Zvch1t���q���	b	���>V�F1R�O����{��:�븓�!C3��Lm(ՊR �b��=Ũ�8[Ğ�����6&D)0a:Dg�������3�,�����5V�1��x�0��X�T�r��;r�Gl[(�u!�~�k�^&������X�W]L�ֿ�k]���}��,����S��wI�\ ���&c�K?y�q�Ú����Y�̥��D��P�n��7��ҩ�y�x�"�2.I��>˸��>>�FT��h��������<���15�mJ�A��tn�ɋ��E+�02t�hB�,����l-� �4Y^�eCǓ^��h��M�D��q1�i��|XӸkd�"�H��ss����~�\6��S
���cʆ�7���$�j��Ú�Wܢ���Ȱ�ý?�5��9�����M,��w� w�Eg9���.�Q��� {���d>A�2��o���Lಯ�,�ұB��թ�P+9@h�M�`���!쮧�Hq�ܐD-�K�7`������چI�;���o��$�?i��]��=$�]Q
Ɨ&E"�;Ҳ�W�������`���*�v����8PP�5�D�e����*��Hk�����ŭ��yL;�����?�E�|*��A�+C�"H�Sʄ� &��NI�;�;>n��.IR}����2
�˱l���R��Dл�d�N}�g����nŋ@!��=)�Y��0�M�t�Ε�X��M�:*�f΅$>�o�,�r&~��lY{����8��>gZϋ�7�x�G�Jbϯx3]-����)��}W
G(	�&��#x�Ą�L�99����t}�7U�䷏�2t������(�����~�͵��?���%�?ݩrk>m�7����C'�w�SJ�':r�o��:�lxc��z�>���&��rzL�E��&�+o�Y�@���?E���>-ìu�����n�����tBn��)ڀྰ���xE�N��_���O�5i�| 0$��a'��g@�����ߚ���Ǿ���_��q�Qէ6'p�ar(�_���Z��M;�p�I��^�37#V�5�*�3�Xa\���̹�]`��+�(Pgr��0� 8�S��3d�Zw�܊,}��ئ�5�%6�j��	t�~��ю~�ߝ�u��p.R�'�i歗(d/EX��F��Ĳ�,��,���]EڇڹMB��O�;�6�5)����m��`��tZ�C���6��ԑt�W��w�%����@֍B%����K0UOj����9�m�c�?*l�{��w@�G��?]H���L$&���[������:�[�-u��0˛��ACuރ�o@'u��h�����T�lI�<��c���|��(���p�eaI[rYarL@����#V�7>���ͩ��<��Yِ����]s�k�![��m�W���DD�{>	�] QL/�h�6?�/a��B���
C�*�\ʸ�F��@����@h#&� 8G���έU�pym� $	<v�:B\�ֽ��tf(�K�"~.�<5*���w���n��tv#����/JT8*�7��g�x>���ش��iڋ{��X���=��c��w5� $�CvM�8-����~�Th���W�@����y�Hcwu���N�Xr��� �l�u4�Ш���k�n��P��x�o�W<���2��8��U�� vj���!}� ���j���f��]�E2�}i���#���ߞ-��B"HD�n��t���w�����LSxi���m����F�t����7����o?�����W,"bRZ���ML�X\⋦ �����w�*�J-��8�o��r5I0��l�s����߾����C�v�Bw~Y�l�`"}��qbKW@<�/;��`�a�g��8��Lc��B���l��h���������>�P�E)�����r��"�@�'�R=U7�ޅ�nųq�.�w�س��`�,Ԉ(�� ��*2�E��4򭨟���n<v�c�>~f-�ι�Oj��KÐ��Hs�)}#��̬$Uc�Pz�B�����К�����wQAF������ln��4w�C��0n^\�8��[�	��,#\�Ƚ��&���3*�Z�)�y��,��5�890
����*��3�Q�F��bL��P�4ʂ�H1n���
'���s�	!kJ{�NNV�V�+��P� ���l5�ӭw�
.�J���k�9;V%��J��\�O]C���`Һ0F�c��_YR��&\��?��s�œ�*P0�@�É�0CEḨٖ�G
_���'��T�V�?���(yrL��+u[Tv7�R3;e��ֽ[�'�T�9P�0��[��2����j�;l��5��ì]��K�����a��Й���w���EP	�2쩃d�ؕ�=�^/9���w�Fy�9{�r)�>+��p���o���8f`�H��t�}VN�������ݤtMd@[y�L��
 ��̠�(�j�a�*�b����ԇ3@���*bR�����"v*��;�Z�p���`���ǃ职n����BǇ�_\5~G<J9,��'�~���C`L��%�f$Jz@�'��ܟ��v7a�k苢/Qk�h��;��]��38?#O1�/��o�=.�m�:O�%���^ͩ���W�a�!O�ð�R�So�b��;F�0
��#~$�N6Ci*N�6�l�!_��JzN�ө���h$4,�k�����卼!T�N��^��g�F��ntrRO��h�j�:����*��2���n�P|��_�(�������%���9q��p^EvvFt�G
U��9�>�
�_Q����ƥ����-a�@%�n���H�/v������-���(+�d���dt�D�%-������$ގ-�3%��s-xBǥ��F���@����۳���c1��-����$�mtc/��3o]�_{0זb��̺����aB�je�i��_@y-��QF��ЛV�6z=�Ԉ��� Qg�|��0��K�������X���qÈ)��	��f�����r�V�z2���\]�֜�lz��&|�h#��n73�|�e�
�Qq3k�c��������d2ܰV'��0����6&� g:rfq�F����݉��A����Ơ0 j��ǒ��%�h��j�z����������p��t0i��li��@K��y��>�Jq�5�b�L��㘏�Ԟ
��S�IY�Nn�K,x_���o}%)��w����`0Z���=��N�Ǡ*�JY���B�
�w�Ɂ��֪��l���#�QK��ܪ�7�X�7���:��*�%�@� 7a�B_�� 7}�9������>3��n��s�@h�w���B	:��"�Ȕ6�k��2f�c�1�ʚ����K5���^l>H��jZ/O���Ě�����1�$��m(��ށ���0f1xi����y~"�gd��DI�4f�Ke�.������,�+~�O��\�f�J�
�/�o D>�O{{��}eV!��RK����#���*��8�� @�wɇ����Y*2�$Q��s�A����WmŞ��Tm��b�)�6��K��.��\	�~{��'�� ��u6��X4���N�ov�6a��ptq�`'Ȁb���WU�%F5�"��$�o�����1�5�Im��Oӕ���+���K���.���ߗTp?_��qC$��M�m�>�\�4r�!�?���:*T�<\��6u�����t��#��7�=���i�!��`V��6#��6t�g��s[��Ht��t6�(�<���hk/�K�-��,�d5e�UQ�Y��4�R�	N�f2*�Ő1�F�P�,V���A�u�)������ĭx8؊�$u:
������=�Or#����p�x�`]^|�����ry��T�E�$�*�O�����J�Ѿ�I("lyLa=��?t7�4	uY��Nw��r���\����s5"�-�+�������5���}��Jق�ԕB���vK����K@,��á�Q�Z���ڐXG=�z44=�rq�a|���D����9�&��P笯���,�`��Ӹ!��f����J����1�	������{ef ��a C/%���ڪ8��<��7�]�8��_p�$P���5��%h�9_�5����kJ��gN�v��x� ~�T38lX�ԃ�G)u4�dw^���_��F%\���9��,G��fxwU���CX%�46t���QB�:	*�����\�rY	U��|�Ϟ�u'���+Oc��YE̓2�o��3~��}��cݦ���wMb�+G�#�vOl���R���Ȼ��@g�
�g����͠ۀ��kk>1W� =�g^ȿ�^zʡ~�{�#�{���-��x��9�z�f-������$�4�I$;��>���|�M6[��o�y[7*���פ
�vr��X�>dy�������X&u�PF��&gw����!`���^��h�v��V��ϻ��N`ZV���X�<����Rh�ԧ}P���_�u�,u�±��5�����z���'/.�R��uj�q��Is{� �"p�g�[���D�Q��J����LKή��8jw��J'euu���Q+�=�kp=���y�6�Q�����^���b=� @�󊱊�'#�A��3����Hߨ��Ѭ��]�O{����Ѥ�/�R3�� ���$6�����C�E��#9�
ߨ�S���0��b�V|͇,o�l��=%�Bb���[�6:�b%,#���#	dpqQ�8���J�+d�CA	���͸Қ_�4��!\.���ɦ(�Ln��3]\���;��៿���iJ�
�e���ί|F'�����H�EK�����0%؎�Ŏ�����NMT��p�f/�"��Of�Z�[�ݦ;�s�0S;C��Ym�?`��n��q?�L_"%C8 ��{�������)�֘钽�������]FbT;^�3Z3�$���A�+�˨��ХH�)��K��R�����02~�A�Y��T��Q����p�&��T���G��\�*��+Je@��L�׼	"�����~#�pPk��	� M=\�F�B��ԉ�W�=K5�ț�Έҙ�J/�ecƍ�̣vb�6@&l�b��7^�W����J3ǰ��.ԓ�����DC��hg,6y�����F0!)�$�?{IJ��ч����U"�N�;���I^� �S�xv�-��N�m�O�bL�� ��j��S�D&�DB����.�^��,��.m�xL��h���b�;�>����B���nA��TDfPշ�o���*OT��`n��#7B�®_%�.$u!��/ ƧN�-��7�Ù��%\[�p�X��?���;��>�R��{�$OTQN� �R���Q8��А<\P�e���o��:ֶ�}�;̇����S�g'��V}��0��+J��{�n�/nS�ݶ
EpD��)�O��O���8f6���mtɾ��'���g�чd`P�J=����K�7xVTsٹ�BZ��lq`*����8#���Ȥ�yD{/x�يP��x���ľ|����5�q���E��˼dN�!~���%sN��s����x
�pZ���eb�#�����$5���W+bˋv�%��l��Тe�<�e�xK7���ǫ[}����V� ���A?U1J��Ng�ߪ"��53��E�J�P�:)���x9��_ō�*�����e�s���3=�MjN=��Q��TL%��nn�a"� �n��
���s��(n�]J���	�KV1�,�'���")n����c��gW�5��ft(���$�v�0�a}Z2�D�X2�%��s�=0�i%����?��%}j�8�L��ޒ�,M��a�n2L=U��B1���B�u���9 k~tH�$�W�f��P<h�7��g���� ��D� �q��\��b�~Q��QY� ݫ7��_�g̠ĉu}�Lö���s2�P2��78��66�=- �%�x�XLAG�W�E��Cv���;F��gaPN��4_�Q!�8���S��ﳞeX�����B�L����S��"5y�Rl�.LURX�D�q�k�����RQ�L�C���ﶦ�vsNw�T�0b��2ܠ����<]��ś#���$��8�d{�����U��&���F/� &��}U���k�F��D?�Z��׆��(��X�~\��=]ԐYQ��v�Lbo#E*�|��#�g�' �֬����Z�]Z	#�g���U� 0F���ʻJ����S��0�����᜛v�D:(6V~��[2̈́����'?���X[Xlw������#3�)S�w��/�����=o2HB���;�����u���3�aa�)�x=���諎�S�o�/�,&��f뎻r%R���Ip�v{�X��#����9h�r%��ann�6��0f���Z;���`���wk��5;�M���7�w��/�fjxRv�!�X]%	;��A�J����k�}f�7|��[_�%I9@���v�-D��ѧ�B��.�����p�G|q�r����= ݱد�F��q���)<�f�<���D�G|�6j���$J�j<Q���B���8 � �<�&�k&�B��<�_���)�%A~j���$�3 @���\�]��ka(֔(�f?��-�\�{���	o1��Q�1�ed���w�Zˆ�@���C8�,�A��^�(r����.ɱrtS���7s;8�?�̩�Uo�X(�fQ�FSĹ�պ��VA�8.�K�X��Yoo��A�+45͟�g�}-�=�ic�6�^`���O���8�xK���J�P"��8i$N���@^��>�K�Sc�6ɒi��x4��7I:������<��詻���[�}3<<V{RU���<N��oQS�%˟LC<�����~�g�1]ty��Z'mS)��C��ԫF9�HN�^8��2"��oc%2N�0��
��.Iǹ0r��E�R��C�#s���t���72M��E���G�$Z�a�����#�Z>m�a]P�Q:X�(\���W�R'��#��̊�6�������NHz��G�ܕO&��%� �^c9����;G'�s��&y�N�W��� 
�*eŋK���|�5��a?T>�><f��,@9XpN�筫Z�9Njn�ւ���ĭ�F���䋆�A1�L{�Ag�|`�;r�YLd�����S���x���4�{�Q��zd( �z�c�f`l��q�]8��1�۝N�� �6��-��q���#KM\�����9nuhzƛ7��{���x�Z{p6�� x���Me��>�������n��	|zxo_�3���?2,r&�zn���$�~�so�'r8)�;����'u�W�9�� �##�o�'�Q�\	�d ��h��7C�j�,Q�C�(߿+�� ��X���YO��g:5Lh���}��5���,�!�h��D����e�Rhyrtu��o [�-gwt����a�oT�Bv�.(.Ł!B7޲�]x�Sˆ�z�A���b�e��EmP�
�D��􅓠�(�^�\M{�
_�q	r��\K���ܑ�[&�Q���<��,�s�g�h�����)a�ّA48�����2��ԯ}�}з*xr��o5;�h:4=.��f�ZO	�C ���c0���9�b�"�?L87�П3�c��L�54a�xI���1��*�J�ǡ�i�.5q�Z�b�{0����Yz���X�W������g�<�w���)�h�y�`�fnZ*ږ������V���w4�줞WUi���,_)׺��Hz֙����ԭ.i:/G�?9���ȳ����L��e�7��\�7�!޺^fJ?�e��idZ�C����m�ʹ=�Հ�L8�f��S�����:7��2�M&xb>�jE�G���j;$XAe�Q�������8KQ�*w�"A�8�6!�|���wT�m*<����V.��)��^�se�(d��e(�xS�ׇ�k��>U��8z:BI�238��k�S8�q45J}����S7l=��A+v�mzh��U�C�6�e� qn�b� z����yt�B�&�4��0&�\��]6� �)x� ��L�c����	c!�Q�>�B�5��������&�����O���yY��OLx#�r?��7���Ӓ�!ɯ�8� �Mg�T�j���Y��٢��r�'��� �Ѧ(�|Usp�>�ps���"�Ro��d��|`�0����h�΍�L@��g,�RÒ$������SVpE� ��i\&D��A���Vr�輖�2Y�3Zlk�l� q���%m�~��9)�ݱE�W�]���)��y��?�b�{���A&2��̥� �n��GrN�����m�ft��J����$\+p�t�;�H�r�06H����-�â��'ۂ��{A�����d ��%���\*����VA��T����)������9D�J�9�΋�JAn�H�p��㘰y�^�{�T*w�Wc��͢���矖3�;P��C��!��*�e�E�uu��E��q��P�ZGz�s�$���=�.-�Å�b��� .f <�FÆҢښ=�E�g���T�e�|���؂#�8՘�D��WR����$�?Sϳ��n���]^-eB~T�l�s}e�
ڜ˻���FO)�1;��4zIQ�!��5=�i�z�UE���fű�K_�͑J��`l��6�]T��v�>� �k:���ڢL����EU[�"��B6�:�|2%|!�,���ҥO��?V�!Փ�K�v���B�S4�qo��@�9�!��3%1��YȄr��u���٤��|'U)v��@.���es���Gw��:c�[�}�<�7���G鄪�m�3���R�/�%��a��V�r/y�S���\�p	@������B��w��ӧE����Tl��^l����պH	�'J�����`m��<=��o�� !#��4C5�V���a�#�Ǩϫ�~��˞R�8D���r�j�rt�0�٣���"�?��}�۠+��ޟ��q�1p}bH3�����z|$�A6�:�5D�\mS��^]�xQm>�%u'J�/�m��lK����^�_��g�L�!�Lq��9λ�0Nb\[�[���*CS�� L"�+�S)r
|L�j�}��o�%z3ۑ˓Tތ�V4M�]bκ��6��-��I� � ".˨��6����̳���(ԺwmBUF�ؕ��N�L���864Ƀ_aS��te��V�U�2�{J��52�tJ��xܥ�0�,kcƂ]6��^��+H�'A�Eȇ�
�G�>|0ղ�gN34ő�r�4�j�Yڙ��<��J˙�h~�P�����lw���q��E�a��F=���7F=�m�\M����q����qSW��e������w��!��~)�Q�K`��  �������3/��{9�FY�ࢼX֡��F�N���h��Ø�[�j�(Ԃ�t[^|a�R�;qGB�e�u|R�i�v��~�>�Ϳ�CRn��c�&©qv{R2D�oI��a~zs����Cd.�*� ��4u�M�"��&��s���d�ˊyU3��0c��c>!���Q�W5�L?g y{�R#�r�V�t|�v�}�i#�U��o�h��f[_��OQ7Of>%V�n��2yQ�푺����t{�U_	nܒ����b����&��K�i��ʶ��a���p�яrb�7��nfZ!�"o�g#y���G�l������\U5z���?��5&`-䛄T�ط�S<+�n׮����kL'��`��WjeL�Nm����jQY�7	Ćv8YѢ�`ǑE �g7�+J�p��{�4S�NVH��?���Moxf���÷�d�Ix�}1������gTV*ɖ}Q�:�VU]����}r���ث��V�@ ��|m\��[J:c%���w��5�Q���Z�����a������홚���%�y�Ϥ��F��*=6�z��{��S�oؓp
�~��|��n��}��}<��� �p�}I�[��E� _@��h����*!�q�ʒ7r͙yұ3:��*�h&�}&� �FĨ�k˨XN��HS�␉N�$5��F�i;���m"��Na?��\�W�h���7(/^S�P�Ъm!��<1�s,l�J�,��y��4�ĶOʊ���x��z��R��f�3Ya�y�F�U����ϰ��nw��Z�����&}�2u�a�j���1�/�k-5�c�R��H�{�^�Bj��>������Y����7�<E�D�{ԭa��`��ю���^��]r�;Pa����K��?�U���<vػ��;��z,s�͎۸�+�V��i2���Y��d7Ͽ������]f��ޓ���{L�$^)��������x��(�˝4r�����ρ5�|l� ��I����E��yh�d$�5�Q�Ȓ�(G�v|�g؆&�t�E��+ҡ|����Gm�H�}�!}%�\��w6��)϶-�)�m;� ��=Ƃ����-k����7$/�G躞�ƥ��F�4�m�GP�._���R���^^��XF�%�᪠J����`��ՉY5F�� L�]�J��;Q��e�d倨�lF��z�=#G1Y�\�J_Űg�&װ�!�L��*�Λ4^S��	�m"r(c���"�5Z��_F�����Tٯ�5ͫMk���:�� A�PJ>4#d�(|�XZ���G�#�D{[WxL+��[9�g������c,4���x��~/������G옽t�A�7�����$���F���2
6m7���\��5@aA~h�oL|A,o��&�p��Wb�d�s9�{u������+?�`�_��p�0��ԺzHt*������ �Q�^yo��j))|�Dkk� �f*w&4�ҍ5��=.q� -�9
����	���y�dy�k^�6Ď�[��9�Q�Z'`����5�/P�����Z+��>�'����ұ����@�<�|������b��	Icb�㨌��|�>�'��5g#�р^H����&�NXb�>�k�i�����	ko�Z`��r)7~�
0��	����F��אy}�aXEz��[Iʕ�?��M�[����Gf�n$�h�8��=����u2Z�5>B�b޶�oR�V��2��2��TF�D���^�Տ|&����(l�<,וl�)�@����1=���,�m�Hj�s����Q�׫��^��k�|�Y�J)�֛�YsR_\3h��ey��6��Q��y}���"#
�Zi���j��tD���!|�fθ�?\H��P��P�n��ɍc�{��t\��Z~f��MO0����g�}mVߑ�hz>J@�Y�o��>�����U���`��A1;��o�w�A��E�|�VkQ���Uĭ�s�qi���W������6��v��S9��ϯQ�Le��6���M99O�6�Ź�$�d�P���m!�1Hw�z̛�tJ��h9g�଻G��u�N~<�ս����hB#��7�l�;I'ӆ:�N"+��y!�\u-�MQ�n�����<b#���b*�>U��̹�$=wD`v�ӫ��d}���у�eh�0��lQť�]��/��@��)�@�S ���&	Z�6���e�����'j�/-4K(xʑ����S�bin�q�2>�E*����,��Q^<h��]�m����C�a�*`�k�R��(>�߬V,SRvP��Ʃ4%�@~�Qa�a�g�|�t�>�Å���̻X�y�j�H3S��j˥�M6��k�H�F�;�4�����i�WVT�5R���ל�z�*�;ƀ�	�<Y�v�7��jCO��C^u[9SU�����0�4E!�^�¹V`��)����`�w}+����&���,�Rw�*�U���V���.�)��9��q�Иn�V:x)����6P�i�r�+xG���!Lnyl7��A�bE�oKl �67�;�Z�Ё`˲��f/�~}1��AG �i���na7�6�q
�#�¢{E��UQUg��2���W��P��{��h3�^[�!��-��8G�./>n��ⶐ�a�oˮ����g���]h!X���w��h 5�_V�N��a�l�eTRṀ[��2���u{)����=!B7ǡx�M�Fu��K���^{'$lX܃�<�S�o5ӹw�U��z������ja����W�7�v972�c:+_Y������n;(���y�W����p���ڦD��J������9BhCL����׿��0m��I��̇��a�r��+��[��>��q�4�lEA���"��7����a�?|W{ʵi���@c�d�W���|�s�,w��}�k[\䑅7%�e�>�'>г>hZ�VЊ=+E��-;��/�-�Bj�>��຀b��K��9��:�z��e=�]V�u�ܟnG��@�X]�I��ڻ�Gk 2l���(���wr�Z�V��x+!��ɭ6��W�	1wW��	2��9f�7$��o�I�w�rRuy@N �20?vyh�Z��n���ǾB⚦l�
�D7 ����	4�'*���,��g���aDNޓC-nׯE�����̖_���n+n|�"�Y�Y�C �����S.s_�g�y4�2t�f�
6�xo^�����m�:�王V�~��VC����Y�D^7^��p�T�k>�`B��B'�p�����c�F-h�#q�V�F������9h�V��IW�Bj����m#��N����ngr�<�FÉ����A�!t45�4�L�(�X\U��Ku	��(V�̃��uEO���i�y���^eo��t$
n��Y-B�,������#2��ʇ�3��PIt�o����CI@W�Z�6���XB�(�MG�s�ǝ2#[�%G�8]�˹�Y-�.�>< �=�� rH�@���o1�.�O�cIh:;���v%�hn�2&�j�q��^�p 
��"��ڬ�ҠA����vRG���x��Pё�L� P���&!_�~6)E=�I�����y1��m$@�怨�r
��f�H'�Pe3�#�og(�9ݝqo��]W�42�+�9]�	=�!��xzɽ%�*U���F�"�:��ՓlTY�f��n��Ҝv�)���N�	s����|��H�yY���wVk�wٗ�� ��~/�:j9ѡ7�,k��������������r �1�����k�`�����ҧ(ep��(VN������}ǆ;�q:�>�Ev���=�Pa�����A����j�s�}�v�^aH>�h�&��_U(c���䗾E�r�^_��f^�Sz2�1�Y�ރ܂Oы��O4�S�=��@I&W��Y����r���� =ĺ��w�˰�G���&U��4����J'|�ۢ�U�������[Bٲ:�|������iEf�wr���J��/j��&�ay�QJ��a�?`Q;�Z����#��!>��.��خ�f�lI�7Qf��vF����O�Э�87֏w���a�j%�S�&h3C�?
�Hz�'� �'5HK�o�l�r�ȧ"��=�j�'x�R!\��}`B��[��˕vq�قO,�'&�0�*o��_��+���n��0@y��W�<|�qD�����xK���{�GnȦ�Ղv{{5�i3Ru�*h`A]����Ft`�e/>�� �.=�+���C���Ȍ���^��ne: 5N�RL([o�����tpb&�=��'i?7�Z�ZZDm8^K��"D���"�*� �!^��B�ח�v�;T+c��6a@Z�{��(LG���K�QG�o�.)�		[����=�Y���������
 E֭R�	����x8�� NZ�����2<��.L6��ᎉ5 ����ZB�?�Z���P/�������Kւ]�w��k�a�}��pqYH%���jZ23[T=�@�o&�����\�~�u��S%��9NP���=�.!�ʺmX��<����ڭ+5�r�X҇n���J�f~��Ĕ�Y��2��rs��zq�_&R῵��eXkx1���͇k�Y���4��p2Ŗ>e��Q������0/�'��Z?=b$�~��Gѱ�x�+�:b���`&�m���F =�.a��܊�΢�	�+��2bT�²��lJ��}���	N@���j�|�i���������Չ���<���+j�ʴ��DX�{��Li{pR�E�3O���d�7���+o}�=㒔��}��2��FxT��]��d���t_f�6AK	�R���5�;o(g]�m
gvqÞ�ě�:1�PA]�A�q��$�ږ�K͢�K���'+�1� ,��C�6CQy�WX�R�m���i�9��B7χ͎��o3/&D�`3�.)�gC̎�H�+z�Vc�oy/�bFyu����bX�H�����"^�O�qR���־Cr~�������ڏ_teDwؒ�"����4��hG�HF��ޢ�=CT?c^�/x)�1���?X�B7{Rs���XL�H\J��A89T��Ь0�8cPl2�8�FP���[��c���K#L��ް�9A3�mqv�����Ϲ�J�����/��Ҵ������i��g�;���l�RBҭ%[L1����4(�|��?��W!ud,��'
�|��S7x�m)�ۀ��;���˾A	���xO�U���!��F�C�؂-Z����U'Cp����,"��a�x�<�����A:�����X3�F-����8���<��cs�xc�J�S\���?�.2Z,၁�E]dX�T`kg
J��M����i�^Z&>��I�iכ�mW����c'�[��9����ĸ'����s[�P�Ճ!;��\�xA�M%����o�KϚ�/�	�U9�;:fi`�����|�->h	G"t{�Zg+����"�`8��t�QBL��5#۽�,�i�d8������ܲD�I.�Is�	V�����o^	�9���D+��֮�m6g�N�5Q�� oRf���d�}l�Ҫd�Zy<�rk�i}����t��]���m5���3����sa��[�+dtf5.Sտj�!5q������)��q�"�6j��ʺ�K}�:Yp"�3�F-S�ˏ��.�S]�!���^��>I�:�3fǼ�&��=�\�Yu	��	����ؾB
9r�+n/��2�؛����"�^4"�Z�;�>��1[�5���n��`���s0�js-��^W�<��@�8A����`:[?�g���_m��B�1�*d'�,I���^� �;i�p%~?Ϙ	ۿ������A�P�a��؀����jx�j�on�m�g�i�Q7�_�J�PN6Yy�2��K�V38Qɔ\:��Y�*zUk[�]>2��v.��b���}��p�<��o���KŞM�f5��`�9��;9%v�2,���xݴ�P>�k�(Pr��O�����ޝ	���˯p��)d���3���}�+�>d���y�s���z��e�� f6I��u��eR��z�PZ~&�{��4˘yqR�`P3�xcU]~��pc�R���(�g�Mŷ�4�U�6R�G��6IA�i�q�2��
fV�e��)��Wo8H#���}��✇ңk��τ±�K�p�{���S��^��Ba7�Dr���5�iH�RA�Hr=�Mzu��y��#kO��4m�q��� .I���-l!�3X�3h�#�$�����^��A�vu*�JYC�F/�CF��l�7��P-)D�4 �!��%����
�`À���^�v`��*�ٯ⎨��4�ä�q��`c��ɖ#���4���������-v�>�Iĳ�� ��υm�ȉ|��獞�(Բ��'���2������Z�/���3����D��������w��8�xr4��գ�D,����L�X=��Xӷ��U��;�`!����v|�?�q�P�-�ڑD/���&9��+0�Ev��2�r���}8�cf��a���R�-$�쒙�D�D������V�nmPf�x��Ĕ�m�>���-խ��F� ]�x-�I��.fܲ���R��k7u���g�v;;Hb;i��V���!�,c3�����;$Ԍ�L�@�l�%T�T�w�2�ٸд�h)/�6_�~TH@���V�R:�䇆>ic��Uތ��������  d�����&��!lPQvF`a� ;��T��s����������8n���d�,߹�+nD&�K�]�ީ�n@٫n��2���uZ0E�Är5���hY1�6��$[�.���C�Yd�?�-4 �d^�,�0��w��n�P*.�}��������fnr�������[���>r��Ѵ}?��d����3,�pHI���0?&��qx�N1� ����=��CY!�3��O�����l�Xt!�8ȳ��	�8��lH���|.��j�<������,�p N�O��-�I����˫��ی�;VHL�@�߉�b�'��5f�?A�R���o�*�jy���.V�֨-��D򒽸����>;�m/���aH��s��m��+t�~���p�ٰ��o�s�����r�8Q��<��e��EWG~�8Iń��4��m{`�a�y�����j���Ls��Z�o.�ܢ�J��o	r�h�y��o��z�-.���Mx9�QC���n��!�>�;CQ����E�?'�����ĉ��ȸ��G�y�!�d�
D� �4El�$���@��y��k_�
x���v/��@=7���*3�xZ�����*ƕ��A�ζ�Ñi��ϵb�Lz:H�ݨ)(�Lo�v�4u3�~�+J����p�>ם���&� �>\rk���5�Å�b[2�ipp�v�\zl�D�=��S�	6��B��[(��&*��j�~�_b��Ӗ��(�,l�2y���o@�ךǞ��\q��^;5RE��w܄�}��*?q�B��¹yTƃ }��(`)HG��қ��z�:�/�+�X�\�V 5"�=T���k�翳���q�@K��3L��Cc�!6��NX� %�F#*
�]am���3o�˰���Xj}C1�Q��Gȹ�nc^^auy��Y�e&,��D��:��0���o16�4����5y��*�\Zݚ�㷔hy���ϱ{ٟA���{s�r�����s�H�#wZa����}�͜��^P>d�wi��^�N��Ĝ�9լ�*oT%��4,d�n�.���eg�{O�d�dK:�t�k� ��Nd6d���H2��j%�.6v�`-�)����M2`�H�v2��f� ��!��lT#7�і �M8^�_g� ��(Jϵ3&ng�+f��������?�ԟ5�6�<��{���i�'�uU '��-f��8g�K.7�Y��f�	A�PG`�:'E�o�<l�jfkD�n	:�%tM
��4S��4�j�Q����]��u�ޞ4�?��f�A��!����K�tu
���9�V�g�@^�� >b���e��ں����|�%�y5q_���8����qy���H�׺��{ O��P�r��;Ӡ��wFЙ,�T�p���t���u=r�E^"Q�~˒kG9�U�����T~WI�$�i��
K���5�����0L�����t�+ppK���#�T:������ '=mVy6T9���H�@f��3�I�*G�'x�7�f��R1Ӫ�3�̸�i��X�b���̶���!��bˢ�Yt�:k�B|k����_�wO4&2��ar�����[�w��o���n
�-S�|�����}�K�8�0���!�D�*�N�4��b�2@�KK?r�3k��s�5�C��A���TM%�sϮjT4���;G�Ә�bLW���nkey��X��w,K����h15�I~�1�&��v�J�D�� .�iǜx@��/��}d\:uF@A}u����./�|������o,
��m�cr�^i�yyx�C )a�un�o$�z���y*����E߿�B�f�3�C]� gX�T^}����e���U�[P�0��V�cȚJ�1:0�*�Ųm aM;~��u%@:8���� :�\xݙPo�w�]*�ƼRpHn�k$D��@�0X��f�C)�	DX ���0]V������;M%��P��q~������9�Z望�w�sl �$fG�wl'�5�c�fߌTǸ"(�����my����7��)��<=�93��'�H��
����D[|�x��t�E�����7*��{�Ձ�˰��9�ΠC%�z��v�ԜTeS���m|Â���/�=W��.��O�yQ>���)��_}�+1�FHx��!.mU`�'|i7�c=?fQp��->�<�w=�M��1^2/V`�z8mi�N1�21�w�]i9PP-��̒�������q�I9署Ӕ9��k�MV+�Z�e`Yf_�M%w_���aHW��Zq���Y�ʗ4F�|<=��Qf2t}�>sv�:��4-�0���b;��"WL�[�y"��*��D���<���_�ԏ"V�E��גL�C��Jg����8F���'��Y%z.8���(e��(̤�~b�&<�S��Qz6�z�p]��H52���u�,��R?������	��}_9�bN��̿*P����DQ���I,�����oj4y9������r�7�%��aL��[���SI�ms;=�C���ŝkVq�!�c�~l�l8���� 3�{������A�8(��t�\�6˅�� �޲��X���q,����{���x�}&��5k��5Rk�6%�+A�X!%�ŵT�q���	�Wm�Lɟs��5���Wǹ�։�=�4��������5�h���0OJc�g�������)�6"�����e��7��2��d���ٚa�v�gڮ���]�M~��iy�4�^��Pd�=��$2
����\`�\��ןt�ߺ����ԗ��<'��J�N��[�@|s5����r��,�"S�O��S��th��nBB�{a������t i���5��L���CD<�}�Rƻyw���C�+����(����#x����gY�7̸*u7�g9fı��i��;�MY����̠AM��6����^-���[b��U�yUۋީ������0���T�w�U;�eQv��ାf����A[Na�^C�϶A�w<\�5�:����80�VZ
��~��-�<J�c��"�H%�W����C�Ͽ�­�aaw���r7����'���k�ª��2?������7��z��Sv��/y\��6����1et��#����c�B��;+m\�g~�4���5���r��N�hSsL����&.ͷs d����{y�������w��|�ٔ�i�J��W==W�#m�>,�s�m�$�w��1	�z���<�O���G/d�}2Ji�����d�Ub�0X�P/��H^YK^�ނ��B/���g>䏹�Ch9�g�z����X'U���R����Ͱ��.,����8?$����1����Fқ.���!(��3�]�)�+�4�/����zz�ZD�b�ֲ:���c���ν{��1p�Bc<�-N&;]���07��q�mXu��}Ͱ�d�O�;�S��Ӝy�%��
�Ys��B�te��"��܉�(�}����%S0�g�Ȕ�s���˙H&J�F� ���A]l�a���,ov��+e�MR�6�g$�PG��HM�Բz���:z�{�Qun��m(��FQs��VY=�sh�}�j=��"�a�m��{���z��С��.�	�򀷪�4j��<V�@��HD��r���u��$�#W�dmgs�4�=Q�3^ ?{�2��s�s����#���76Q���`!o���	G�2�|��������c�I���E�����N!@����(��aYv��UFS�Ŏ�%�Q��WxSwR�-�c�J�0������V��w˶�vY6F3x��PļZD�3̠���U�FN���B�N��úE0�%AwY_��dY�fg\���i�忏4J��@��q�����W��$R��_��2�t�	�22Ȋ������׽�̊&�1�İCV����RL��Pp1�y���5w�����e�!y92P���U�,�0�ebü�p�Rp"����G=�%)r��	MI>��	�a>)�0���;߭��ȵd\St7@�8�<��蕝��
\�)�P<yD��ywd$�~��=�c��d��������w��-f��K�V���
)�5'���K� �5�t#x�+�.��O6�-$���Q����-@m�*s�>j���u� %~q��=�ݹ\��x�$��h-�˳�����F���&ֺg������b��׫{rfw��b���z��x�a�S)iŞ�� \�@H�Aw-��]D�|��x}�0,M̭ؓ|�҆�������N:�C��nm����dOM��� ��y{q.�|��}���ۺ����q����+ܪn��9�
z�0
V�.�W9��w����Tt�&���$�b�CE��YխAbH�D�c��D���%
�������L��bD�P�bZ\;��������,���PO��L��@��A?�^=����d��PZ8��by�
5\�l�'��ۓ�`Km;L�ө�#x|��ظ�]HfE㰁(K��3Y+���c(��b��"��C��%&�I2t���76���N{���/���B�1���X���:?�7��Z?D�E�}��z�@| �<�k[#���jϙ&k�k�k�k����ɔ��ݺ�JUO��jz��	!3N�hvT���:@��"�I�Q�cz�"f� SdWO����2踦5,C�x�[C��^�C3)���lZ6i���Uֆ���^s�z�-?���YT�Rs�'\�A��4��1uۛ?Ҫ;����g��g|��P��_݊���^�C�+J����R@]�U<���L�y��湋�dI�~����8�]N5r-��3����c>0��,����r.���I�L���=��ژ��'4�b/6����E ������ېYƠ*�v%�/�FURt Q��s%��8d})B�u����=�QY��)�	�*���mv�R�|zt�Pƅ�Ʃ�Ep����|bw���K�Eq2Uh M.\�m7��Dc|e����kR	����Xc[���+[�N�~�vv?/�'���VX������|Ÿ�P��W��U���R#�#2��?k/�K�҇��<�5ݦĆ�����ɥ��A��ۦ�I����<�,x ,�i� IHAN�~����H����u�����Qرa��͵����c��t�5[�I��=��1��DV�R�R�!P!�K<�z%���\30L�?m���
�Alӧ;w�y3�R�v����╴���Dd4��4H�O7�(>E#�h���.٤���T���v��Հ:���?gx��Q�O��%]._�@f
�[��1���=�9�W]��ض#Z�������U(��,�w'��
c'��Y=����1�9�R����hD�M擺$3�q�r>Œ��4�z�}�>Yx3�d<m�O�ш�>su�6��|W>:�>�EBN���J��q�Kk��!����3P-�c2O�-����e�/+f����ր�	c����?o�;V�t�Z@�QӐY�D��� p��!�z䣳�G��J�"�a4���s;����31���E��i�Yu�J����M��PL�90�;[L�Z�;��g�I W��g'�ϴk��ս��7"Bv�ņ�b�i6\��}�0&��&�m�Ӻie�W�ff���@!���%��#fa����&�eE�]kR�rM��1Lxz���YIG��cIJ9�1ٱJl���b�A�డ*����/M��:�E��g_K5ԢLqkۄCM�Ӗ',$3(XT���v_pgع�}�ZM�U��Ǎ�$�����߅�����{�$d�|*���=5?K ���Ps�� ��b��4�%��a�z�o�e��"�y����~�IÍ'ߑ,�_��W��K�,���TL�T+�ty���	�_e�Mg("���e(�'�YU��8G�o�'�l�5�3 ��%m���J.3�Bo��N�_��kZ�L�6q��İYd��Nt+��ɟ���H�ffb�YI9Q�����1��>_��޴�╻�a�G6r4훸���Bl[��݅3�C�����H��n1���~�"1ϝ���g^��#�k�1��_��Td7*뢃�S�ݣ�'fx�-�����)	l���s��C���u���E�*�
��E��������cO��v�z�>K��y�mV��r�İ,q�MM�;��k�Zh'������������ �����-�����xy�r�gG�/m,�,�)��w�ʳ	�Z~vu��VJ�b9��_o2���(��}����8EE��!f�;�F�`��DE�~�� H�.�q,p�3qrZ-� ��`䆟�% �����x���P��L�����̧�,
�	�������nZ���	َ��LR�F�Q3(t(}�7����N��[N�Ѯ�%�s��|	��ٻ]�xZO�ZsWg�����V�� ,��;̹\�c	�,(o�dc�F�4$q��]�n��ѧ�C��LqA����	���6�{�.�Y?�:�.sX?8T6�W�F"��ai�mu���ia�,N�!->ۥv<��cˏ�����U�̄��7Z�zAed�o'�y}?	����rs7΅z�L��~��R����f/f�s��an3{?)w���@8��g��3ɗ@u͹(?�Z#X�����'޷��^��� i`�u��;�Y�+�!<�r��ɺm�俋�^��C>\| t<5.޴���~a��aMk�;��4O�3(_�t�8Еu�.�0!]��\n�k�j�Z�WY��^�r�x�5:�u����
���o4�:��p��JfN�ߌ� �E'V����#}rT�η!�8A��C�2�����F{ɼ�8�a��{p���T�E\!�EC�Hu{�y�A�ȷI`}�L�1���2� ܒ��o+B�P�~��8O5(-��fr]��B&y�Ae�9VV�����<��s3���2����:.����m��G+�������g�:�ߣ|��"�",{��I�{Կ���w�6��Gު��3�W�m�O�g��i����`��tw�t����C��
).Q�g��X�����U��#�]�Ku�`�ߖ�6�yE��L�'6�::{ι��W��2o�� $>ъU$��n�ckR�7���t�T��5d�EZ��C�����A�J�c+�z�baN6 ��T���ƌk1	�g��k���^�p�h1�uC_k&�(J�iej�cܳ�����i⌘����X���%��f�n��0�+#�&�a�̄ȝ�MR�WkOzg�e������}�0�t.[�(7l����)���í�g;d�3
�Q��D�?��; 
�0�B�����+v�x����C����S�nMf>��x�^���
�Fw?�lh�m�@�? ��H��y4�U��`�BV_���7vJ��L!i5Iy�T�I�")`��Qȗl����m�ʛ��ް>�\��90�b�;�6l�؜��I^RW���x*dR6���YՔ
�{�%T1J._�|!��L���{G��^�F�8�.1���l��_����?�C��R�V�]]�K@J�
������4Y�����a�ܛ�H�蓾� l}���z���(�Q�jE5^j�#�H5�$�W(��MG��N�i� �l[�}@��vl�0��9H�%��m�Й,�k�5�C����t7��BAwa|��0I�9���a�^�h��!��N:*��/�Q"��0�d��<���k���^s��Cs_= ��xirq�dꕿ���1��C$˂���f�ի��r1�������{����B�y�Jᦆ�b�-���o&V=����5}�,	ﻠ>/�������2�Q*� �{%��<=���A�w�&��]i�ՑT�F?&����]��f$���*�v�i�3ͨ���4<GV��sB���I?AG���H��_.�#�8�8�|T2g#��xr�Ji<{�o(��(�4"e5�c/G�]�bu=0�љ����U?����Ɂ��SX#8C���:q�2��<�����M��8@�P*ňY�ƽf�����H~߭�vY
1s�3��tӀ�yqS�������R��W�c����b�iP�;���q���Y�gn��� g�ˈ��4_��D���t��jU$}����5�zZ�R;���,f��M���\��V�AeĦ"�Z��:����~zj�P��e�s�A��]���J�
ђZ�P�֊:i܉����p�G;r��Ӧ��`W;���Ar���h)\��\�dk_��ٿ嶨�n�s�(Z_�c�[)�d�X���at��z�W����Q�a����
e�vR���' b����P�򯮐��?�P��fk���"���Mc���wd?L�V��wu�(DE�L���)�pK5�(b����<�+�Q��,����m�����ֵ���X�~�t��[�x.Z��uf��Cnb�:�h����L��3��Q�`�b�h��#��t�?w�ر�혅X#g�rƪ��!�����+�v�M-�4��`�%����۸�J#����a�6�>l�[�P
��\��~¡�5z@(�q�p�<�~8�\���bn4ء"
�f�V#��5�s1k�!�>�iyڧ�^�_ۘ�� pj���^�z��Ц;��N�Ԝ�����&+O�:�
�`ˇe���Vp����d�{��6BdI�T��- **������%*QS��ԫ��%���M�"2J����_�����f������+]��cč~�?r��I�mD
e-�b�*�Х_Dڱ,��<]������
�,%�q��0ܴ�&=}�?�+���4���GOB�Y�Aa�z��+�D���^�sO3c�h叆�J�q��+225�yP���=��SS��WށX�R��� ��΋u�K���H48��D���:UE��55�x��9��Mܛ̍�X(v��~M!�%�Yq��:��b5��3d��]����7b.��o?�p��2@�����,�p7�s�<�X��0]�a��b� ���H޷h�!��"�X�vyX�ku�?d������E�7�A�'���_��Y����náS�ʮ9�2K�[*��_ccPť�8�}T���ЃШY���W�n�n4��(\`ty�q֣�1�3,T�.X蘫~�ȱ�s?MN~���pK�}����H�kD�ԛ�20�&=o�P���iw��	�2��	h�[kF��˨�| �	����-��x�`�}:���3��'��*&l�Z��f�Ê�'��n�rT���N�ʾ϶�O��PI�ZnZ�$7���]�^8xh��t���3MJ����j��;�+�Y1"��0��Ԯ=�L���]������G�}�"� 1����~����j���\��uȃ�=��۷Ww���_nK���!�G�g�B}�\��vR�)o~b�V��#9� ��AW��@��
TU�Ǣ��æu�1`�U�H��å����*A�O��=���f�Z�������x�������$�j��lV��-�JD	{�(w! Q����x՜eh�l5���,i���~�֞i��6yϞ]egu	��5��Q��w�X�Έ��<��	Z	�@ Y�k���aC�>j� �vX]��t��8�׭����7�ĕ����si�N��EXZP6�R���O�*S�9|�uy��z�/d|U�tqi����d5Ai�'�H�7������?�m��l0A-E4?IJ_�B�y�<����ç�eMBм
vjkF��T�$F5.�O��Y�=�9B2i͌�.��8W� ��}	p/�0�Rt��{bT��Y5�X@�h��񪿬Í%xڿ͢B�Ϫ�UP�To�A\����"�h��6��)_���wz��/I��8�}x��`�7J���=l>�t5�����7lՒ�io~����Ql,K{��M��~����)6nJy���b$�����N�M;�=�\��X���s"�m��\��@��QFE__��pZF�����" �<\x�=u�9u}�W/���v��hE�6ԇK�J��d�z����4�Z�G�(N@��=:��>��FY/��q�}n�<4��z�z&ˢ�70�U�E�����r�5���"�o$ǏvP��\�pu��~@�W�?������&���?>9�y��Ԧ�q�� �uم��wl�0��G��!X��Ȼ55
Yi���0�i��qD�H��Xƴy�qs�{�V�P#U�!�Z\̇����_��&m�&v91�<�����~ii�6�o��������\"<櫾͇���R|�oՒj�k��y��(�A���@����}�QBҰ���&�d�9�9gɘOkr�kN���dH�݀�1����Ć��j�bV��a{�>Őkg��98w�¦3)}
u�\>�+���P2�c��R0p����s�1�q���kt15�Q��i:�˱�'3,i��S�qgZsnz�g��M8�zI;E?7��Lْ�Ql��8���~���(�2y��ҰH�����<(��ޫtM���$n�)�7����œ�{���ߠY��K� �>���1��!�E:��T��'ܧ�u@8C�gL|�lQ�j�k:u�a�^T���%�G6ǜ.A����j	��GO�2g��%����݄�7����A6�a����.L�����Z��6��j,� ��DzmĿ��|�eꕥ^̸!�홮���3�N�� �̠$��7LH��vm�}�	V�a��2�T������*�{0��W�|��'�?�)����5�=�h#ce>g12$�Ed۸|�.���yH�i�% �货[լ֤>g]��N�W�夜������n�/�p*�\:�c��ƕ�hќJ���E6���=قH+�/����eD�S���q�q�¹�m�_&�����A������%���[)�T��a�i�t�+��Z0��?�r����n:Z�Ƶ���O�@}�3���Aa�KO�,�[+l�D�ƭo�m5LT�G�Ӆʦk�~�����e�2�N�� ��}y�4��PO�$>�V��^�_upٞP ��°C%���~'�d�����E����S?0��4�@M�D�N;�i(���3��	$��`���JMjK��:]؁T��NÝ�_H=�4Ha.����%]�5�A7�5��툑9�?�X�Z������79O��4%1� ar��9�?�%[�}xuV�P�Q��r^`�dˉ�h�w��#<�3����C��x���̪�]�]��-�m�J�����v�Fs�8�*̦s����E�VЅ����q���4$/��6��@��K��݊y��ݲvr����h��~5="1o]�x�Ʌ�����:�O1���/VXk4��v�n��}�_�
0%'�V��r�83��8N���%� i����v]���/m�׀�#tȗ��t���L�!׉td��U[X�Ղ�L��� �"M	i��O�?*'C4�*h�r��팮�fN��u
__ﯰ��h����4׮��`�o�o&�wW�˽���W��_���MX��m��T�d|���ͧ�h/0�)�R�8�j6������v���Oά~g��P�R�*I�_X��]MJ��1$���8E=D�OX���5�xIi3@n"[�&�UJ���Kd<j�gn�h�W[{2��M|�v�;/mZ�}�D���9���8 ��8� ] �"�T���e+��r�)�h_j[f����A�ů!�hFO��
�+�V��YM�s%7c�uN~����"Qh�l�s'E�u��p錵�¬38۝�T|?c���K֧YA������G������w88���Ru�����c-Tw�Pg���mU�K��Z��hon0�}����E���t�o��֗VN�`XZGT��%T��f΀���q��`X&�[-�Bf��c�O�P+���?��,��I�J4Uŧ�zh<k�܋�Er�%q�P�Q�� �'��H��)��B�>���/ʠP��_2�+?��>����5t��1"���'?d�K�����k�=���o���݇2e���;���IgL��V��
*L��-��jL6	ma�8E@fFC��PsT�խ�,(��R� ����������� ��qa��3�h�M9b���y>�C��P8��?0+��"���B���&g�����K�1C_md�:{�/9��3�a���"������,g���Lx|�!�.��*�ą��i�x3&��ҝ0�����<��R�\b/�6���}u�Q �ι0���;�q��Ko�mm�=��%%F���A1��'�8�Ϩ���q8����h[j��9�+ӾӃ������o��`ê��~T�H�Z���n�Zן��s�`�uBWZ6[Z�{�H_8���������3��u����Ps����Y�eW��i�N��UbOR�V�vf�f�Y�vV�V�Li�̏&�?v�����/�_��u�i6":.�bm���7`�n�><A�_�ƍF`mF+��	�M8�
�ϙ2�Ҳ@7?�����R�9O���FX�M�9�DОw���ݑo��\kT	�{���Z�֔��'�iXɞ����wΐO))���U�3>�\GL(�>�ג�Ԋ8@ւ��fv��B��t��w�4�q��u� ��@�`굮Y������9�*A�YO�x=:�u�6��H�އ���pt�v,@u���e�Κ��o�l�Q�%zn�ie!{����}U~:pB�k�gD�=�X`��L�3�x�F-�3\}t����tWA����A}e�~{"<k>
��)�8��[�� ���[֧��g�@�/T��Q��� 

��U��-�5�*��l������dϜ!O97P2E>��č!.���}5F�W���8#n�_����?<�O�Ŗʿ��N;C�2�����楃��;	8�)������~ۺ�������	5`��-���?+�gA���͏�2���~.��k\�H����b	z������(qvQ�Oܯ`ʳ�s
���1I�mP���AM�l"+��D���LXX ٝ}�I�X(H2D��R{���3���	�a<��0 ����S��0B�PY$�AXMN�Y����onZ���*V��������k���+��+���6B�{߭,@�A���o�et��gL�C�qoU��2�E��h�����&��}PGޞ���}����.g�%U#������m�n&��.�t�'5:R�t��A��7(th���;��]��{��r��%�όl}�!��	8�~m�Q�X��[C=B��?UPt���,l�w�*�����A���5�le5��5�S���1"dE��e�Hn7���lP\���i$�r`��Ǣw�85*�h˞`Ï��*�<B*%KZ��
��H�d�R-�����n�7�I�b�R��!�u>�IS|�ض��n�>p�}�/D���fO|���T'o0f�*�Ú �/1�'n+w\U���Z;��?lH��D-�|���� u �_�Ѯ�e��������$�SKV�NR��K�x�]Г9�6��«0?�,�+m~�� ���-�eF��J��پ#��[�]�����u�����2��O�n�@+�O�1ʜ��m2M����WQ�'$��2�}�c�����	~ʉ��^!��1��Q)��Ȉ�MX�Jj�dl}��*"Y�͂����>�����M�{>-sP&��!��Oh���<�4�0��wx\:�.�|��ĸ7��4�RCyC��K��|��%��)�h_������K��b�j tN�J@��#��ճw`зѥa�zNH�y���Դ]��5�����J:�L��1k�<ǰ7Z缰Rӝ�N�z��!����'��;%Mb�v."i�[$Hh������vv2z,[�Q��߼PZ�C�࿌�U�D�¼v"~�p��p�1.�z��۸ը��x��;�w%M��@�ȗ!'x\�OgB������D��.F�O 7X�)�t��k0�g���Jt�C�QnX����a;z�-(�sI+=��V��n�l��hUg���i�b��V/�B�g�u�}d��"j���Թ�c�n��B%���54��O�F��[��e�iRఉ�H��<X����j"�U���cM�J�e�Ef��&�!O���q!;>C��N��T�5�Q���������G����n��rͅ�\g7�5��r�������D!�L�<���aث�>�b_�Ec7a-����N���t������ ��,.N�Ogߪ���Z\�39S�������	��W:��k��6Қ�����Nnx/wF_�fM/Ft�&(闞�R*~vm��Fe��H�F;L*-�%���^TK�)�5��z��E�5��S+���m����l�~�0~��r�2���^�ݵ\ELv����#��&��}��B�B��1H���p⪒*����͆�zT#���w9̮�C���� ���E��������xѾx:�i^�d��Z�a��̍ZP��,S�S)�Q�������ME�U���w�e�����7A���<2�M
5𠏪6���ݫri]��F$���-0&��8��	�6��������Duxrc���.`���0����y�	pz�V'��7��`�y��y��P�.	3�:8)������,��L��
mhM9�����6#�g����3�����B�,�2�D ���Q2�&�:F>3��oK�Fn���/Pf)�q�<dXg6��2:`��1Ů�~�JK<w@�����T�r�j!��$���v�v5o��ʢm�N��w��|B�ɭ}X$Y��;�+~���:?��Vg2�G�OPLB�Ė�g�R4 $��Up�3�(z^���tKRx$t=)
X�rۓ��-�O���*�F��qqnk�����*�4�x��n�i���}�M�d�M�����1��`���g��9q$k#���]-�Q��g�d[񭸖eZI:p��@E�}7�t!���Yˤ���TXu�(Ѥ-?��cq��|�f�/��o�K�F�r�3K��<V���_K9{�y�� ���������2�_c4�H��zx�H ��Z�ʋ�k&�.�X������>:0��F�z0m-4&;�\�PRO���$�JǾ-��RU|�A�>�834~#/��;�S�_�(�uY�08P�U�Gko���Jc���a�≷��>��-�/7x�X�6���ͩ���P������Wc��I��d��
.��� �R����q�ΰ�lUd����E�Z:M������3Zu`KŤ�]E���P"_U�e��X���h�T�C���Y	��+�|�6袼|Ec	��U���5V�P��rg�����B
	���:m�*kwD��=P��;��e9��^a����yzE�)��UqƦ���q>�,�R��\�Q������3��y�:�n�`����ҋW�`�PvI�F=�R����{5H/K�z�:�O`�����v�]r��+F�Zj�-���nP����MF��;-?"Q�S<�^y3`<���j���XM��Nb�*�ak~�#K�O��;	�K��=x���29-֡}�.#:7��/X��hp�$וw�߷{�_���Ƴ|)3v�@�j��g���6<�x{�w��k�:��PPw��f�}��~�C�����^�i ���(�9$�	����x�j�3x��7P��E��o2y��f����N�������G�]��kYm9�d�&� e�Ț���Ї���K0q�,[T���6���2�]�9���
�vm��;:i�t��3+]�)��x ��PrH<}�������e#�e!��O�*U푼n̝����vf	�6IB�H��;n�	�7��d��[�toZ�Ȃ�ܒ���|V��u�q,��!C���]_�;��L����"'���(��y��3��Z4�ˆ��Љ��w u��ú�j찰Yd=�	5�f��� d;��%U�
/���!�r�җ"��؋-� 7,�p��<��f{�퐰\��<�&k�m&2�kw�q����2�E��������éL�x��]���,Ib�][٤�h�4��h|t�ŭ�7��Q�6X
��"I�3|�i|����TV�hd�ZY��X"J��g��!��X���A~�.�u7�RKu]OH��E�;-�;��9$G�z��1�?Hu� K�"%n;�5%�����|F�#�A�iԛ��Փ_�Z/V�~������K�c�No���5p#��2�ၨ�2L�{�[`��>��[�j�$�@�#I���ݹ\�.ڃ�A�t4B�y}��i����:^G
]�Gٰ��7��X�y�u���4����ܙSӑ ~����RA�l TmJ��k�Z^��:6�RD���N_X�L"@���b�D�寂5?�W.g�;��b�{�L���:P��Z���pm�D���*DK�<�I�&�d��ؿ���cj��^�`xU��uIu�׌3��d�wF�H��
Z�A.��#~���*�p�^�'���z�z��A� ؈`4W.���`?����8��Z^/�s�p���+�ӊ�K�P�u�z�h0JFl��t2���w�%1ږ�Z^���'�d�'L~��½��� �_��0]�YA�|�w�J���#H�N�����z�
���f=��_�ċD7�	*��R�ŋ�]P�:x�D澗��Iԩ����xf,��FFY5�]TV�}��vKt*���cW�㕋��z�#�m����R*u�L�%���do�)"-����ͲKI>}�8��Zviᨏ������@����i)Y�݂*}w�A�ڤwno�tq�y�n�xqCf�6�T�j5<���LMU����p����'i6�d�������]�����2ʐ�2�+�d�H��*[ikCA�q��0�AqU�����F���=��:��O�>5�P�ze���Z+�f.!�Ky������۳Q�!f,	'��pR��v��e�x^��[)3ДF����aq�D
�^J���a�-��e�.�\vT�d�.�t+��_�sh�dv�2tr�`�
����OuR�����0��s���W4�Qz� \P�n����U�!g�T�r�L�S �o�ƙ���^\qJE�j����u���l>��c�/kE9��+���G����K��7)��붉�J@�1�r��D|?_�z�ݵ�L�O;�f���P��y ���Z���
���fu�r�ˈ�z�
��w�31;�dl!�R�t�|�mM���W�`�t���	`��_�ۇ�ƿ��O�U��M§�f0���*Q�J@�AZ� ���	�<���#Xm�A0��R�hF��o�}�YU�iu8��Ǌ��ؘ�JÙ��51p��q�O*����`�Pmi(�ki}�R�\(�Si�Gu��u��i�@�9�M��<՛�eQT�	��9a��*e+�Ǖ�{azn��P�C��go���/lz�vz�[�5#�3:�v#1x\��*�_mLd�&W�P|H�J�[��!Z~C�P�������<�e���'��t�(<��E))����g�=B�Y��>)s�
�"���� |:6�^v������J����-Vlf¯�6~;���g/ʝכ���R��%��qBsȩΈ��Mҗ�:>�!��A�Xz'k��͂�vz񃇠�:s��AF�ŐF�9�1}vDn�?�w��>�hk�p-�� �=�8��Q�U>�^���<�%]zBC��.^��F.X�xe��ߎ^�"HtU�Q-ii&����j��H "r�W�Q��(��in�ѵ��.F�u�F4�����4�m��Y�,%�&Y��M3�U������͌|Z��B�ǟ��P.�흍�{"�p��5-]���\�dy5^4$�Щ�B���fxgL���Xz�k�B^6�.>'Zbm����������#��3���P)��&�+��D��������ӕ�kdw��������U�"��`�I�wv�e��r%Oy�4ۥQ`}�	B�l|Ck�yke(l��Gl����Q�D�l�tu�а���o��N.��\Y���S�� @r�lD��r�\�-��C�	��Ə�w�2�Ȼɮ�J�Y�4`��*�����1V� �UMQʧ�)pk��h����1�K�o�����A�6%h����r3t��[�S��F���?I�熂�Z�`��zؾ���E�>��#ޭE�Gk.���\�d+�'v�<j�=��'4�����Zu�M����#�6�j�'���_�| ��ߑ�o-fRB�5`���n���Cbo�SN����{����FE۝�vK`:�ce��W�~�Qޙ��k<Am��5S��O���@2��s�l�^Ց��i���VMQ��y:��A˽5H��O^Di��
A�Fs
U����E����=�$o|�����	`��mV6��1��O�/7��F�g�>nmi��&K)��܎�cCN��t�S�>W�Ѳ��;n�y.���6^њ��X�,L\��_���� ?�����l=>�./�|����q�q�� ���Pe��9P�ŉ�Fਫ�������	�;�����y�A�)Y Ȁϸ�"��C���$�࡜�$�E�E��aD�PU���^ow��
���H���K>L�����\gh�,|d��$����-+���X}�������ƽ3G����^W1'����l���xծ��E�� onR�%�OM��� �0c�A� �	<��[�z�E͏�����E�Q���~E
I^ƛ�9*TS�Ú�5ci��߲L#do_t�����$��)��6:��6�}c���,���ږ�L�yV�	?ݘ�u�E�fr-����S=��5!d�Jܡ��w� @Q�#�����/���|_��g V�b�"k�f�_}z��˽�?N�����}�5��eVk�ܲ/*3��+���)�B4;�p���UH��)�->�o�6`/ĉ���hY�W�t�.G͏�����KsF�˂�SvY� V���v�嗭���7f	�������!0�8n���´)�*T�f.4{�dLQF4f�qlj2`�72`���Y�{�����zN���YP���YVM����^�ߑ0�.6�E�gk�������TV��&�c�0��"���[�1�е��z�fP���փ�ΰXޖ��T�W�!��8�x.���\�4�+9�9��0W�č�a�E���W�M��"}Y�o:B����^�fx^���j>i�Y�oǏ��m��l�1�P.��Be+I�>kYL�:�q���W�=+V�H�a��cBrTW��g���v8��F�����׆G�%=��=�����s�b��D;�A�.a��o�e��d=A������ye�H�	K�9lD���8 EޏT��
ȋw��4>xy����+ð�լ=�q �oV�s͡���Rv������׸��B�-<������/⠛T=�2 �e����Ѻ6���藐s@���m�_��7�ځB���R�1�T8Ƞ�`�<bC�O�2a��W�_��8��u�`abu���$��:��Qs�l�D����6�V�3,d�z��������-%�����,�^bWn"�h��5l��p� ��gH����o1�?@�q���f�2�<���3�#������x
)�b���\-��	�k�� i=1�=�\0�$̔�3�~� )ql�DE��)]��x�,�D�=~�F�D�	W�q:���U��`{�vC|�H��w��!{����ͮcK0�1D�,MB@.Hx�VT�3ru�u2�N��=V��r6�_|SڏA�!¨�1����
Y�"���!V��ϧ Y�`��qL0_	Gs#����W�pט-5z���7��69FЂ
9���s�C�O[��D��?�T�v��V�ԯ��#��ړ�ؽ���$s�R�]Jf��]���x����Z<�����b�򭚆].�5�t�Y?�"����qd�,+Yr���BA*c��)��X}{��o�hU->l"��왪:3��< ���\X,ԉ��şzE?(��Uz�C17���^Z+Փ�AZSe ��ؚ�q27���b=WCl�[�K>�6�.�$Vt@�z]�}pes���29�v�5���n�^A���D�z� a&^!l�k��X�^ہU�2:ּL�B���'�%�'��R�����L[����Q���	h����oY�և���xQ�)�\M�;v��r^�Wg^�lZ��\d���	bv��Ԏ_�;�����5���N���Ѣ��o�w�����(�A/�@܌MB:0И��4d�C C��!-	�0���4��{~n�P8hhL�o~LCcޞ���#���Mha7�9�$���)T|����)�
�p(�t�p�_�3��k���䩾W��j�d'[�?�!^��w����Zu�¾�jɣf	�N��ް���'��CK�K4"���p6�
���%4?9T�{5_�A�/n�i%VB� [�?��jΌ�D��!M��a�F�1�/2����T����og�����_�����j���?�%'}ū�t��S�6Z,z	��]�o��3X\n�ͽ�7���;�Q�)��E��/���b��Y�Dp��6(�q�׎^�+I�i�o����#�iwI8t͆Ԣ|Ua�7��@.=�Ŵ����h:
��]S4��e�{đo߀��|4�\�v���hV*��K+�/c���T��
�d9r@�i���C+0)D`��c���6)����5I�c`�w��<��)�����f�{|ѡ"�$ڷ6�ۯ�S����.u����� xYT[����4�F�Pf��})�s#��Tj�@�^q�~�B:p�i�Mz쨰u�C�`�Y�|�lQg�Hx��6&y�2�̽e�b[���+�$s�	fҲ@ARZ�"�z��x�>1Qf�-�s*l�k��qzz��c�FjT�C��~5��zR�\a����ה0
X��z�'�q�YX�b��^'8�H���\�bڭ��wI�|�fL{�o���RA�y�d�@�	�����Dt�p�d-�ä��lX-9�>�H&������ȏ���l���\Tի�QU=VL-�]ٌ��%O8��̵�ֈ��E��E����E��|@(���� ��l��r��#Tz�9ܚcC��<�,-Z��z�"�;j�C�Y+���^ k�����̽�W�/E��	�Y�Dn�� "��B�p^RTgr@h����i�ng �|�1.�S:��k����I����H������D��4��_(I5�e��ݳ	�=��ӿ�C��H�rIڞ8tf����%*g�#�`�p���%����
�R�Qe���ׅص���΀d��Hkå݅�4� ���<i��{x����iX�C`w'ᑀ����~K��+~��b�=
�{ɫ����k���U�ڡ�#`|���	��yd������7)�[�!�H��T5.W�9�w�|������&�j��؀�Q���<��d�g����� vI���K���u���	[������T&�#���5�W���<$-Dj�9�n�ㅲ���K6�/��wP�����}�����zfH*i���(����JBlI�{,{�wX^��R�z�CZ���|��+B;�5n�����*@�P@QJ�Ҕ�I�kh�.��	PlM�x�	Vw'����.���DpҠ/�Fك�E�����z�1^�Јq��4-��jcǶp�sJ�y��5P�m��0��I�Z�3�rn��'+�F�_�qQm�b�Mjߺ�GH>7:�� ٴCO�a��=��t�UdO�f;P��T���`�����W��-�&�����Ι��9�~R]:< =N�[���C`��'@Һ溜��<d�t��>������]F��9Q��r��$�g�t��H]��H�X�+����7��On�6�����[鐴��4&� UCVK%�+7�Ÿ<�����kW8��jO�0�]F�;E�Vӧ�0�w�^k�F"���P�N��'+e��6rʇ�4X�<mGa�� �rn)ci4�XP�_��{0�^G��d���"�(�ve�4��)4�D\ޗ��p��U�|*+��dh:�&��C��
W�v���}f���b����g*���*�����w�8�����b�4���n�Tke}�y�Arå��(�di�U6wA�gW �U�t⡂��d���~O���Y���b(�1L�Z?S�>�V��sr�<�"%�3Ʊ�Lc<z�.z+�y0�|��yԌN��vbJݒ��Z|S�R G��U�dT^jsaݝ75�z�K5ƃ�q8�P.O� �/�
����3Dd@�$
b���0��F�p���\ƈ��y\�IRf=����ˋ�P1Y�ɕ�k*[g�S@�~O����M�$:�~����`w:�Is�D�t;$�ȯ�o��-�"'��l�8$��f�ӛ|e�����M=s�����Bu�@�Ȋ�h�k\��J�Av�F+��J^Xn��埄�ꉌ\�����+Gz<�Z����xP}�bK������
m/�� a!r�Z& ���2&�ԍ�Z��|XYg@��=�86�@��dSԊKFBf��6G_��LJ�'�l��E�D*�B�+��Va���2v����K�a��	W�Ǟ_#�w߈QS�P���;��΁�v��޸8�Ɔw���RU��@�<r}e����CRJN��v�!���Q0�i�3'���2��<~�s�	�뢙����AA�
����fk�՘�Ԏ�7��5����3���_~^�Py%�rdP�%��Q4phhR�?[j`�x�Ƭ���@��XV���b��4��5y���]Yf^W/��?�1�2>��o���K��O�B��fm߬�(��B%fq����AR���y��9B�e�.����=53a���e�U���D��䔅h
[��5�4�-Ժ��4D����$G�8=�����h����r���4�G�#`*;�f��7�x&B�'$1�jD�/�4-�V���PC����F�NQژQ�l��ĥ����a�LSSd�F��zQ9��!�w=j��G$�F�v�h��!����ڴ�X7,t¬*m���#���5@3?1�<��`	\!1O�J
,�V��[�~LE�'����E���AKȢ:8��<��kj�T�?`���mUp�d���k�� |K/ܱ4��W�N�����2�4�em�ĸ����0	C½W~�y�Nb|��E��\�B�& u�#1��J�Gt!D��p��xV�Y�R;����}/�b\��K37��kUDػ��k�ͫ|���ޢ۸C�⫠U֙�p[z���{�e����Q�j����,REU�-[��b�MϜ����Jx�6��yz6%��%bgn <Wb�2����`�4N�<[�`ֿo?%V�7�`04j���BU��ꭝ}ˬoS������L`�k�݉^ʸ��Z�o3�cR~.�vAd��t����i3m.�G�+8nV�5J]g"TI?��=��W��������Յ�q�9o͙<�xO�c(���,<��`W�;O�Os��1���ж��!�¸]�h�E8i�j�p�L�����EC�4;!-i����'8	�ޓ�$='��G��w�x��Nw��"�$v/��Ȗۿ(i�R�T����ڞ�����x�]O��~�7�E�msJ��\��T�����ܟ����J�Q\B������(>�<B��tH�C�ok�kb�y	g�K u�=ξCX�'������I�9��0��Q	*��MT8p�ȕ�zw ܡ1�᎝���$�߯x,&�d�O>{� "�����0�q
��NF8�Y����ƅ�������l���[A�9�GA�1���}"�Ә�{~��/��B���I�L;�3<�d8��a��e�f4���M2����M�j�x7�P�H����bL%�a�!T��q-/�3�!\�V%��	Z��0�u��g��.W#��C�,1F�]�r{Z��w��>�oOJ�-W׊1��[-ѳ;1�=�o��J���E���k��� f����`7f�Lh�Z�"����G�i�l,p7A�2�F�vv;kI���x2?�Э�{�݂�R>�J�E��O�l��h�o�#�p�'�$���_B8�;�,�[T���ȓ�-$��X�@T+��8��%���vw�J� ���-�fl��+�5��H�; �	0x���@?��5Iв�E�O�|�l))U��`T��	��#{r�8S��i��r�&�$�ƨr���ۤ���ס������݋h;��|xe��M�d3y�Y^x���]G�F�,��#�Gg�kՒ.c�ߴ��~��?9�+��hx��m���/�rl��\�.v1~-�#�o��$)��S�C ����*1�-�df}��/FF����n�/���KcrENb��"@��W��z��jЌ���QwZ$�0�Q���e'����ת�Hq���f|n%��l���\���I�ǪK����	���48Zr��)������1���� $�to>��Q�^ɉQ��Kb�����C!-�Q�<p ?r��l�:�l!Y�fY$�:��t_�
t��r�����\��V;�Iי=��A�������n��6`g��m3pl�O6F9t���2p�
T��Z���K�F�G+Y��]��v�Ma��К*�0_��1���V; �m-����{Ď���}�b��(d�F�b�p��l�����<��-�dn%�ثN�<� _k��W����2�+3�DW�4�[�u��c7���˷�n!0P�(��ZTfXa��3@ga�Ay1'5�$&:l����i#;��GSit5�� (�9s"d �a��x�~
�9Ћ�
�W�۾%�avN�P�ty��#c�k���p�(a�sX�~ 	k �4�����':)5+�W�R�s `�Ԛ7���F�z����q���ҵ���y	�]$�L�R;)x���!�ꔓB�$��|'� b�	�>&�D �&6a0������?V�`�0�*z�q,"R9ΔL��ӵ؏�,#+�:�Dd����+��a��-d�@�E4��T��h��,�S��OZM��Q���n��JcCD�����<)��U��W���c�e�e�'�����7�,�le�
�D�3~]�,���;ᓡ��淉�UCz�빀�A��Ss�2�����@�̦l�u!#����'�N\���t�uE�F7)~�Z䯁S�4�\a�6G$ӄ�<0��X�z�ҚfgX��a�ۺ����'�d6�G�ߪ�vkD��aN��2v%�����%ĵ�g�2��U�\�B}�p$�V7g8�������:���{oЗ>��xnXq�n���݂�m�d�m�M�H�GQ��Rw�U�ֹso�^�3�ΒP��n��ơÃ���s̒á���/Q��%|�P1�v`���hʹ-�Ѻ��f�lJ��6�<�g�_��<��s�\�łNqU�L0 ���^�Ŭ�<o���w}�<"Z���q�J��7��G���b@�
X�U����ڽ`�4�����I3�$��ؤ�,>.��`Jp:l��A��o��.����4�h�6���$�s�d�@MY�T'x�6��-LŔ54:M��%<���oy�Ag�v�f�|�!�"X��^q'欫���&�a�/�I	S�µ4�#�&�$���'������%�iր쉰��<tr5%P~ ����
ۤ��=u�jWѳ4��5�sד�}-Qk ��:�X�(o5�3���̺"��v��/��z��]�*쇆a�Z�>	���G�{H1)���q���I��ԣ��m���j��2/U�pY���-�~qQ�
8O�;��>3�$�םC�2��	�(�vi7bz!��7�We�^��/_� C���]Jk�0.�����'�L���@����u\���1����=!�>���C����"�9�i���כ&l3<�=����8�ZT���>��5L��w�qC]�
\O��1��Q쐧��u~�(��^E컐��@C�騯���?���;a�'k���<�Dy���i9X��w[�� �%s��f%)�^܅�ۏ-�$���"�R?�^_6�+�V�7|<�s���uR��H���u��n��*�>�n�:(ߨ���īldQ���!R@~>ˏ� s5���L��n|~�V�?��X?�x��������d�ϼ�)�!v��*j�w>�Sb�n�X��	���d|C��q2��*�Ofɚ�#�y��F`�w��~��bpw<)���p�r[`h��i�q襅Q�m��$����,���)�0E�ی(����IU��cx+B��4��ơ	��db����@���.}T>C��.�:�)#! �j�� 9�o2=��鏙u�L}�����F�ڲ�N��AN}���.���ί� =).IZ,�g��K
�o#� c�z֎��7������̒8��H���X������@k�T�܃#e��%>�|!�QLϰ��l.�p��IS)ACґ���������F�&�PL�m+��-�isc��(��N~�����n�"�!p�BA#b:n9���i�1 6����t&�e�V$�����#�<<�,�d81m%��6u<�〭�wH�2
�=��Ɩ�2w(֜O��E��l�(ͻxK����8�L�/�u�&�c��7ǋ��"	ۦ>��=:0�#K��I{~������
B���b��/��vG�q�|=��Z$C��M٪���u��wsI9��v���DJ�A�V��]�����AE�n
��$��O��z���"���c?g��W,t����;�V�Be��j3d�s������1={D`v]d��i�T�B�mq��~ "O!iV�F%5�=�"���ׁ�Bw��C$����e ��U��a��c��`�4i���^"+�B�A��0U�z)ݵ���2q�O��O�ֈ!]��
 �K_�N�wg	��]~}�n�QDa��p�5��	�!��N�䩐_hϫi��?�5H��
�%�Z�oT��z���<s����J���2�JDܙ)]���Hg�@E�lH)�U1�1����0�Y��s�Y�Jbر����L�+��E��
�陾њЧ 틪G3��9�T���G��a-�Z�>��9��"�j�y��2�׊�����
qlE��$|lw�BH�D��������n���c �T8���\b�n��w��%e�������ȿ���lc�?S��V�r=o]���X��Fi����*h�T)�9[��Y9�6"��>�8���"�%��W�jb�;a�ӭ�ܴ�W�"��+���6�����k�DF�Dz �>w+�%\��κؘ��-����d~�%=�n`���b�F��T���h���b���s�F6BW]�l���bO���F���Hb"fT�͆��`��h��(R����5N�P�Pb�/b���v5G�Զ�̾N�=ݹf!����̪@�۬V3�(�]�A��N������7�xR�GAB`a8�N���������~k!��e�#�C�Z ����r�60��������ز}܁R�C��dMZ;�Y��Tb0E}�P�S�Ǡ�k�mCmM�.���y3�h��큚T��L؞�ͅ2n8xH�ڏԏ`feS�m"\�svC�Äi�EI���O+@il���ҋ���w�*<	^���x�#H��O_�>f��m�+}=�RV�b�`{�X_���\�g�}a��߷֏D��6 �9"��	�&Þ��E}�p�T��\gM�^͜\��Y��g5�j�m��~��q��*�+��m|�D8*U�4Ig�
F�B=� �\�U��!�8�{̵��s�<�����W�����Z����Y �g��Ώ$E&�=B|�t��`��.\�Fu��uf�@t{���f>ۃ��Oz�J�m����!k���oW����'>�Tj��w��t�K��1���_��?t��/$����-�W0?-xO�,A��b(��<���&�Y��3�x�i)P��N��ֈ|߄�U�
�*?d�g�k1�-��A���`+��O�8cŽ�]6ey�|�+��/b !�=�,	E�ڨưk�� �,����u��O�����������ۉ��Y�	�<�9�uZFB���BA,Ye����W�.���E�.�[KP�|[��޷���8>��Z��恩�{
?�_(�%�#Mc������k�(F�2��*u1h�7R����97���azE�׏����J�]�jB�rBCS�p��=b���D{�\��z�4�Zȕ���p���m	[�+KG�sr�������B�C�x�\���;!�̫~CGF�\�n�62�I�s�]T��? �6Z�#M�WtG7AV�b�,�vxo� w%��/~m��u���C�_����w��3�����O5$9+�ߴ������s�=�$60ōy�T1����+�b� ������Q)J�h�����]��pN�a��m����a.FȎ��'+7�&`��J����b�?�.o���#t�h�`����#��������y�i��\�,�
\
&��Xu�� *��64������Ǒ������O� :�-����yk+ă�(:br!ϲe��Z�T�[�>���%����Z<����'�ɇC�thf� 
&���R9I�b�a�@R�+ND���blɛ�ri(�h��6���P~GG}���5��u���E�����iPP��u��	?��Ӭ5�/N�C9����m�I/�Nʊnc�>M3	�beôZ-����(Ƀ���.�Mi��6�H"��e�
��8��f�TQ��m+5:9mD��!p�B� �+�j�gH�b�u0���� Oj%ϼ����ғvx>[�	"p��v�q�1ZkP�X[u>���hp;��il^U 	�r�Es�n�=1Zy�F�B)�.�Ff�J��T���������� �X1|���c�������D�u��wM��(�X	���&�G�
�����_]^�?�2&p��mÂ�S:�3P��SY��b��i����(��`�{��5���=�w��5+�����4|*���7u�)�?U�I ����Ci�+?�S��B�����N��̓�T�� c��]��n��5��ΥQ�ү��oSل��YF�GcW$��[���=֤���[ا�)�:tb�(@Q�v����`+�o�S�/l���'׳"Z;�/�}�&��⎼G/2^�� �N��{-g�����`�J�i+f���>x���z�m�6�KVS�~Lu�O@Z��^V��م��E4Yy����M���kU��m4S��h_��5�_��!~�v�Y�=ew>��������SHu���yG���؛��#A�Ax���cE�o�:����9�x�V��c5x2�Mjs�[�����;%;ں[6c�oa���e��(�z�A�ҏdպ��/p���ʷ� +�ճ�g�a�DgtѾ��h�����l`M����n"�ԁlw��3={�[�l2g�z���w�����5�kZ1���9� �2�b=��G�K'��m"Vz�<���	�e׵vPG���tQ���i���&w�����Բ�g7bQ qC5�Ӏx5q��*���Bח<�/���N���4�?����/���z�\�J�%�k[����	�������C��(�h$���G��y�dS��k!kF��K�"�XI��B1����l��� �Т找թ%���0��?P�ze���V�w�è��+qw����O�ɽck��-�**-�.�a�l�ec�9Bº��3̚����Kx���Je��/��Hϗ�H[�Ȅ��R�#������?b��M�����g�D�<����K���ʅ���6O�k��0��p������G�"V	��R�j��26���6�)�O��l��,*6W��hN��H��"�M#4r'��s��ަ6?)	5�W��3���w�-g;�ۉpg���I����_8@9�T7��pF�����/8�V��MM4�J�M�&(�d�ǃf|[�#w�+A�����N��?G 5�Č��⢾�BYu����[t&��#X&n E�T�A�	��>@�-e�1��6h;G�%{A S5 ���h\x(��c+d2�f`0X���������TŹa	qn�3Y�ѕ�:r�Z�n�ϐ*��fgτ#z������B#��(��t�(v!A�
�ߐ���²�^�M�{�?#�G]�tn�#fH-����t�6k.���P�w�i&Q�qף.$�|�q&̡_o[#ۣ�J�C��$�k�(2��ˈ�-2� ĭ�v���q��ִ&}c[�	�@b�	@a�B�]9���pO�؜�L(�S�g��{_�XNI݇��H�1Ӥ��E�W���E����ۈ�I0b4���D�T���� ���� &��l�"x��A)�ͤ&c
�8q ��s�}��e)���J���9���(+��SEf���?&�N��#=>�1��� ;Ȁ/�}q׻�:.c{c�Z�zU�k��1�\K^tT|c*O&#�6�5]¹#����]ԡ�`)�Fz�>��JM�1�7*|q=�Qo
}�Q��J��MͫV&`	��ani­]�|LI���D�\V�Г3�����%�-�9N�Лu�r�W���cF���uŀ����P%�UF�Y
�̵���g���!2��a���k��	σ8�®Fd�+f<���6"D�E�j��g7�y�Y�I�jG�֤-7S���3�	�ثȭ�������͓}c�i�ީׇ,�Z
��ފ�8�ی�q/V����*7��� ���?��K��d�@���l2��t�?�H�6'Ҹ��5Ҡ
SW$Yc,��?�ڤ��W���~��ߕ�/�o��O��q�Dh��v��&-�a�[#w/��(ڤl�=�����Z�6��:�g�ن~�`�T"�C�&A3��suW��E�f۟��.�>^y+�e�?��e�,���A���I���98ߏ�W���חv�D���d?G5��IqR�S�.`f��8����zy�݃�rf���u�����*��O�sC��#Q�3�D�uGUcuÒ�� ����ȓ�.\�
![)���KU��.�w�xPp����� E����|#�����éb�9$�Hy?����L�����nS�yo� @��B�x��3�Ic�N0�TDxH�1K�s>cT�}�L�C��:qlQ�ir����3\�v��3�I�V$3aH������f*d�za]���U�����	j��^ߡdr&����C����Z3x���";��L�Е��(��Eֹ7#�]{8'��;Y��'t"����W�c,D��+��S�D$��փ����]Rxċv%���C˹�	���$����C��ɝ��o��V��z	r��'KjF�0��ma���"q,V{?��J�Aep"�j�@}G�% ���fy�g�`���7ۦ�16��,#�y�K�Q:{�T���<n9��7�U��:���]9D«
N��~��[���q7g�]�;�3W����P���E*.��G�:���������P��/�Wt�~އ�>�I�bnZԳ�M�Y����@���|�-�= J&@C�>���|��2�s�����@F�Rf};�rgy6���|kj���t�}P�L�V��H㍫58�<^���0�b�}�]L�z�/K��у��4���Z�O�5V�+��߀v�u*��M�Na��E�+�#�RQ��ؕ�jd�.)�!�981�r!wK���~L�&S6tk�T��X�����qD�T� WYDF,h�Vk�O�'/�D�o���l^�j��/#rUq4c�����@���F3!�4����vزB艘��/{��o�Oulˏ6n���֌�>A�ek�p�T)��S�@�b����b�$�T*F|�J���%SG���l;ʤ �]�h��O�X��聎�d����&�v\%Zښ���"����m-�5�h��ȅX��B�֯t�Mr=�~Ȭ�4��<F%b3�I8�E��'q8�Ov�)�i?_��'����p��D��h��UM�1t�  ����j�N �k~��%�Eh�����O�{Vs��乘i+��#M�a�t:�cdյ�_57^3jN�D0De�T��В��u�H�����\e3M��.
��Ln�r�{Lۤ��CUj��´(>�k� 9��?�r1v�
	-��������u&A��9E�:�i�_�wB���Q\p�d2W��'�sW`�+�&�%*~��,M�I�[�Ԗ�y�5����0��S�Ҵq>�	H;�e,���&���F����~h�,#��ѣ-E�"N�n�@��G���f�6���xEr0d�2r#�� C��WI؞���cn�50��ml��$݅t�b\�k���h�"ޤbC���*f�x�c��p]������|�� Z��)��+*J���蘖FQ"�0;Xic]/A����������'�S�,#r*��5���b�@��A�����Ey��#97I�RJ�*Ƨx,x@��&<��Qf���!��* �C0��j�	žPt�0Xn��'� ��5����,�lF�T����k�е*���v�����������7�D.��ŋKc�E�ъ�}�=h��Y_Nl�����F����@�Z9M5ef7D3��;��Y���ad�L�D�}n��^�'�=����%��j"�� �p�K~
&�qT�١:��,}ℯ��(dMꐾAU�AjY>����i�M݋mG{J� ��	�G��$3ږ���R3zU���D�	�?�a#M�9FmO��ý<$^�8:�y�π�&z�-���2�S����f�Z��t�:�lv��o�NP����=W.�v�9���w:%8���R'c��Õ�P�,M�뤜���	�퉯�e1#�Ϫtq��`4��=�����n�Ȋ�[�����,z�GD�^!�4�ד����`�o@�-rd�4�/AQX/˳�VDё[�K�	C�2��3N�����B/��/���Z�o���e��:3�=n$�f����ZE�@ٍ�S?����1����b�V�$G�(�N��p�N�&جƃ��u����Q���L����4�7`D/ʹBA�p{J�k'/L��?_P��S���pz�d�z^sȃF���T���K��2���;����O���K� �j�*�h%�tD��^�8�n���%�9���'9��N���R�Z_��-ᖼ�����5�/�4�3��Ԭoh��M������n!�K�y��}���G�����yXvLaS�����Z�۲t?p5f��@ƫ?���4�2�L#I�:lq�yo�g�{`1�
�u�6�L�[p�Q�Fe�N�R��k7򌠼1�4f.:���q�����;S�I�i��;c	��X�T�{�y�遯5��{�������2�o���;�c�o�G���S�-���ۖ#vgh4sU�����X�7�{{Īf�`1���SoB�����Z� Z�����?�@���N22�bK1��>��˳�������nm�/HW��b���ن��vN7��6���Q��,�ۙS]�N)�UOo	�-_�-Z��y���%�>�%n,F��V�ʅl�0N��G�1Z���4�
��Ԕ �B�ͨ�6�$�n4mCD��1s�Z�u�]����I"��PXν�5y�<	�')pM�j����7>�i
��*�fû��agM.x?pY�r���|��1X�X0`�b����pq���Z��6/�ҁ�X�/�i�Rs0A!�V�R[/��Ɩ=��5� Mms�j0���JE/�G�.]��a��W�j6��ZDߕr��y
ʽ�	p20�6�wI���hg�\j�@w[���m��H�b���$׬���j�N@������-n��5��5��љx�s��Q�0��|��\����)�`�g�1�[����1�=�)	3��X�l}���ehۊZ��r���K�%��LV���g�#�^"?n�,H�)3|���hGd��|���۫ς+J��Ά#J$�m�=���W_?T���0*��C4�������
re�g^��*C�r���#�W�5��~�����@D��b�C�T�jׅ�M�+S�h��;ojf��A����t��%��������[�R�ًu��lb72��\v>�@Ѧ�N�x�ܞ���2K_h�T�࣑7A�A�"{Ӈ �3[�j�βj���3I��no!F���d�E�?&�
uꬿ�x�=���a1>�iQ:㑄��^�:�Y�7�y�(}�LnoUYJ!�'�U��X�����/��z�noE�!�II"�d�ˡ�"�` �Ϣ��l0��
M�)��F�_8��̋eE�'l�>��G{��23z9�|�"�I�|����| q��Z18�{7�n�δ/6aQ4�\�؛����x�gn�����i���b�7�"��>�di��o&s�%�)@�Є?�6 -��#&Oj�A�GJ�=<'}��Rç�U�aIm�V���]��������<t��0��*��bh�E8�{��a�jg�!ن=+ټ;�/�'Qհ��7���T��I��E|Jw�5�髳/��J�;��	�ꇒ�XEj�P��90f��l+o"l>�<<I<�U�u�h�Ч�ͬ��AF��t���)P]+6:��G�pAq�S���b9of��,BD�p
r�oS7I͛[�?�fG�D�C�#�Yg��[oMk=�z2c�*-ǹ�o�5k��9�`F���Z�>�5�BD��
��뚤�~R�~�Pfsgs��đ���\���?>N:~ ��D����qѸx3���U��jz���#<����4Nż��R~Z	<�`k�/��_C� �����(�Ud��pv0Y-몱$^�m*�AC�<��n��kz}�O�� 	�s�'��g�'b:1~����`���l�)���I|�qϾ��|q�eֽP�O1QjaG���h�0�$���[-��^�0c���ƻ�S{�t3Q�̜Xm�������Y_ÎM���W�z�9v�H,�y?�љ�����c�ԯ�jP'�X[v��[�|�a��i',-�`�����7��L�����$�HB�>�
b�Y��z�"��x��mI�j��fh+~��e�#}"j����5���kp�. E�*�����;��6u�<��V��݄.@�����>]�؏J��+�:��q���?�kM����(<��A� �&��M���!���1vo�-� z	��o3���dQ�A�"i����8^%jo����"�pUm�Yy�p6-I�`�F�� v̕�ʩ/Bwrf-��;'r��7/8ʚ���&oYI?=.�B��)�
TE;����/P�aR�2�O ����\>9���ID0R�G���*�2�Y�ũ̬� d'��y��J����s�����_���l�σ�U��N����TN��2�i�==�������3��,��饋]�HJ���/���NU������&q�8������HL>5��1y��/�ց�W���*��]����:��/?���<DP48�� ӻː��e���f����)�!Y�
ʽ��W�uaH�>����q�S��2�f2��A�%�F_����L��F2`�A��j>B�g�oD�l�ծWpDD�:w�=�{`U���F������e2ބD|��G�!�%������}jn���G�IߖD�2Şh�x�$F{���È\1~��Y'�Ovf�N�� ��>2-$�<̃��/�����\9�B�`ٗTvjZ�ӿ3��+���NOs�y��;���^�
�n�%��������N���C��G�M~߷�f���O��p�L�]c �.�*[P`,�)�b֜�@��wCR�^)�����a:86�8������p��'��Q�r�c�@X��@f�0�D����:P��9 �r$�q"~��_�0�e,@ ��7�\�vM�j�\8{
 �Z��剢��M%����~��v(�l��֜w#�=����&[��ߢ�������p�ů1Eay�&tv�Y_uM��7iO��$̮�<�$�⾧��f�����# ^�����Р���0����1Y���?dQ�����\ l�:\�H!?��A|%�FL��v�銻pL 185�ޟ�dv���������Ε����SKӀm6����=Ρk��D�M$tܞ����cN
�
��s�%��Z���en��2�r�؏�g��n��|b
Ӓ}����n�a�A�y$*�.�7P֪b�y^��a�@��l6L,�X9p�=��y�R���T��Kl&PP�Rf$��s8b�;R�����bS1�/)�R����ީ�����3�XOds�_���M��S3�O�	!5�$��/8���N{��o��&m����#����ɢ ���N��O�a=rS~�C�{�.Z��dK &��m�r��d6����g�Q���qxfrސZ��[�@t��N� G�����m�@1�lc�"�CWͤ	�K�Y�챾�*���m���@�{ �u����5��sl�UXz�z!���0>��7�a|\�-��� ���c�-D�3]���+37T��1���v�>si3`������E�}�TT�1��>�jɝJ�^�:U�)��Q�.�8X��ǒ��lp��.�(��T�lz�e+xN.Tၝ3�٬�^1�aqk��&C��Uw���h>RG`;����p;j�HD@U�š�Ɔ��.)�����J)Q(y�ۘ���8Sأ^Oa�4��e���4Vs��̚���	�
o�����t�^|ٌ���쯏�E�z��S��g���w(��L{��N �p1H�\W$��Q�����B�'�m��WحFdEY��c��U�s ���5��'�	��'�_Z")�#�o�ӿ?�W���-�`�-{���Y���~?@i��N���ݾ=R�G�W��U��hi���/b:���)�^�t�ٍ�®mD*�����r{h��ku*"	l�u��6k�H!�fg��U�;��N[��K��N0v�F�@�2 !��$�(�8���w�'�Z|��F���ED��3,� ��v����-��pÁ�	EK�._F�R�[���M���;�*ZaO|�J��g�&ʉ������pb���I@h��)k�@�����]�2.���8�Rd����6��Ȅ����?�1��9g�F���B[�떕{�EbiHd���[�,�����5"��	+��&!�����{b�7�,��va�W��8K��)͕��~`z�!�|RR�F�h\�2�]P��)f�`��)�Uo�Y>T�GPs�P�.m����A,�/`8Ѹ��;�V�D �u��?[����LkXWJ��7ß��Ɋ���h�96��7�wA�P%�����PƦ���]Ճ*b�d2��P��N���ܷ�u~1�d^��rی0� %�щ._�a����]1poErN�- ��V��	f��|'$���Vm��QL������������,b�'����?L�9tK��y�>d�3���&;��;���c#r&1�!*Ͽ�>�y��m?��g�iK� Q���	B��aUY¸�O�v�>��}���qZ��g��MxH����f"~�bHWE���-�Bǃo�_����(-�鍝,3�C(h�	�����&�J��G��ل^���+��U>����'0�T�6k蓞Z�.E<���<}�#�>�x"������q�LS�.1�v!n�K��Xq6��LSWBUo�}X��vP������ŢѰfN��t롋�e�/�q�i*$9���4�L�ь��gt����CQ�$�����"�Ev�H#��łF.L���Q����U3+u"�ڹU�ұE�y���J�qw����>��t�H^I���jJ<����+�~-.k=1.C(�	vz���Hě��-"md�����J������R�C:ut�}�J/�O�USq��uݞc�6��E�`�=�>V�۟�=��93�L����V�>ȵ�{$�0�)!WA��y�R��H�^dZ�!��
�C��:�vգ�����_1�O������:��J�c��Dc�r��u�N��e��jF�t�5i���	��j���(�����~lc���Ӯp	��+FI��-�&:���E��72���VYxE, ��¼� `Uw�$�[,��R~�"�@���-�N�pz��6'���`?c��X�Pr��?����&X�M��E�>_xع�=@��[�[��w�>�Z�}@��y��2jUB��,����V_��,���`g�Sw@ne�_�2��Qw�ۦ�|�zC˘�X!��w�$�J�v~w�I�
+���wa�3�� Q�h����/_�p���P�50UB\��J����c��*D� #���`�\��@t�qO��ǀF(�����x��bx6c�n_3��@tr:��}�o�ab9D�"50���Z�^�H8'�D��ϻ5R	.���?��_�TсS��1�n����C�A\V<�A��3������7������rSTii����_�o7+�z�3�F��fZ��0_��^D��'�~`I,&~D� q,��y�eV�~	��f��[y_KL�� ��MY"���1L�O){�v��J�3�ؚ��T�"�,�HS�w��}&j��΁r����*�[��щc�#ƛ]��9y�����3R|�Ĳ0��s���ӄ'n�d��S�x1<��>�؇�w�@L9�/��1����-i��f�����xuT�������[5�4�ʊ����iMtE�Ƨ
:�.2��@�X%/�栐�Z�>�Tu�FPC�r���N g\�����GǙ8^��bV�;�g�������_W6��u�qu(�� D��C�e�:v&�\I���|o��MJn9L"2e(k)~�ʏ����q&�)$>��zP2�(|-�ZM����2x(x��1��H���r�М�~Ė�2�����dZ�ox���a��rX�K����V���o��ϙ����v\�PC$�D��Щv��֓�q��ekf*��F���`�%�7�%�)���@X�kiZ{�f�ۜwWRϏ������k�k|����v��xSWK�eYH��bP� �X�*2h�3=�Fʉ)]��*��VW_ڵ�&�,X��	2���(��#�UCe�K�c[+��` ]��a ��]�J�IOܳ�eGϿ �����Z��	��ӆ�W���#V6WГG�=h�/��T��]���A~���?�q������/Fۓo���j�'��Fc�$�,�г15�Y���0��R�`�� R �U�}u�,@�: ��f��J��YLM��ot[N����^o�9sf����A��H��i�*".ʹ��U�߹\0��:����D��{� [)���5lx�o��:���6�k�5�e��=8K��l�2��WLW{6��M��0���RI�*��m-.p~%��3p(1M�p{�I�o��������iǌ��Z������	�������2��s�{�)N �)�����3����u����{`��XcxK���ʃc��$S^�Ctp��(*�[@�=��|������d�Lm�ȗ\�� U�?�4>Ϲ�@��a���D@ѯ��D��K�xI��i�D��l-`������U����}%��$�ִ;�T'I��m�Q{�ZL/N
r��@�s��z�aF�N��a���Ge9��ksc��+�$b���aI�wo��Ҹ�?w��I[0iΦfr�9�^��u�n�wl��SX`��{!�8II"���׾�P7��b�ć��U�_u�v�<�� ߰W�]:x	����kΛJ~�� �R]<-Es]j�Umj�Z������"R�/�'ˬ)�Z�,iN���`�c�m��`b�_s��B�܀'� ���/$����\��Ae2�Q��q���@����I}��"���TF�4�^�Ԫ������ �i���Q��?�~�^U�Y�n�t?hE� O2�i��VX�y�l}�</ҁ5���cS/%pɲg)�Y-U%�G\�\ �T�FOCR�-���c_ȧ���h Q��s�F�4Z~�u d/��i��4���G����[5���m�#�ц�l5� e�'���hw|T\\%ҧ�+���'^�+C�y�#t�-�ڄ�!q�N��
Xm�U��<f3N�G���:���]0fGd�k_���WƜH�P`�L�Dĩ��Y'����B{���1��>�%��Wq��l3-�t"����!�/��r�7�3�He��Q+S�or8'���U��ʔ�V��H���j5?~-V c�]�ˡ���ڼ�E����^����<�H��Nl[� o�K�O5m��T`QH���E��ؠ;�����۞���X`��뒿V0��y��HSW�L,�
>n�c�^ꞷF��/¶������w�-a�/$��!{ujV����i+u���*(��w*��p�Ly�Q/Cb��KX�=h�b�hU�,��-p���0�g�Ǽ�vnYx	���J�*?�"U�E@_:RIdjHn-�m����rB�J�$���j���yeF7���`��o�5�K�ܗ1ςa���Rt�9�"�5�g�N;uPH��fQ'�8�#i�}Ϫ�p��Qv3�Ko�v�Ru�� �G�U#Z�ޱ^N>����C�2	�ЌԢ�}oTۆ���st���0��4\ݐ+���b��!jn���{�S��#3|!�0��2�~0�Rh1J�]h+h�`����|la;<O�g���UR���$2IՆ.ו��&7K���5����c.�{��W&���*����f���)���xʙ̙�1�F������o��CR���5��ed;q���7�~���w@��PJ�����@��G!�Q�
�zN�޳l��r#.�E�����%�Y���֚K�/Sf�j;��*#`�_�]��5G'�_i�0��`F�����FK�%k�h*�3��~8��o�G��рw3�PX#�	�4�Wn��@7����O�@FV"�*8�P��_����� �:\������(����D8N��H�sϻ4(�t-�ݽ��qU>��7�O��(�g_Vģg�~���%�T��)�z��<�%y�K�B�q�L8�E�F��N	og�vl~�7�]�-mX���T�9��2�<2c��؄�_���9��ᒝq��ɦ6!�T�$���	�ˏ񞸁<�X�g��#*e�P|��e��D�v���\�Jb6k���
>�o��l�5gD"�\�gN��d�vZ��ʘ��'�4��WG��)��4V���Z!_�=�Zd�1`�q��Q����8@;~Ya�m�g~�,����NU����"�bh�*T^o~����P�̃X��E�yr���QLh�9A�}l���A���4 ���g�C����j�Rǵt]0���"���*��R0OƔ�u Xdf����7\M���~� غ���\�^�R��kZ�5� &�VJӡ*���8�yV��~��O�V���4�s0M;��}��Hm�zŇ�*ɗ%�{�Ѫ����{sɅ����� �ػA��>�� P�[�i��p'��H�9��=�����`������/�y�	����2ޢ�:�����Do�l�p�o���w߷�G-���=�-��䶙C�%e��j�F�d@��]��)j�����V�(63EW�>��\ضSY��9�
f>��V�=�'��k����R:��\a'� �2�@v7�&�ʍ)���ʲ1��}�	-����t�N��\�=�yh�e�A��L�/�ؙ4��.18U�6��Jf��Γ�oO���\�3�6R<+ɱ+	(�j��iO��Y@A� L�U��
 ��Hz.�i�������[6$�^��1�Zeu��V~�M����-w1BI]���� �LB�6�?��[g2�e�2����8#'Z^?(u*$�SO8�ǙtX��Y�phh�������C�P�
�x0�4�4!E�R���\�F��QZY�欋b���%�_�N�g��%]猲�k�pu�QA�!/���p�0D	'�m�]@6�8��8����h����t���O\���:�H3�NfB�0i�vAcoa�zՔr�ɧ�6Gɩ#�d�n��pc��}�|z6��v+�Ώ���q;*�Hm����F�A՗e7������A���t�Kv�
��M&�C9IQ 7�pnԛ��t{@l�
�qq��%eC�W�8�����n3C6/��2�c)=<oU�{��ޓ�'m��oywu5)l	��[i믓/ŕ�@�s�3V�:|e�5ל�33�.��^��u:=���G_�~x1��0)ζ�ٴ���[+���a�C������qYG����^�*HM���Sɼl��9S;)�i��9��]c��&+u[�j��7��O����p�n-.�ME� �������7A0���u�_�!YȬW�_�C`��_�&�<m�.��5M����SUg�q�D�7������=b2J?�˾4�}A�3��:�\W��5F�\�sۭ�N��@����\%e	�!�W�z�����i;����{��G'7�=8WR��3"�����-}el�k2h�@���*�;��em֠{���JG@H鑜c,�'+K�;;�z�J��"�m�\P��ʺ���c�|o�U��teI���3�{�m1/�u4ׇr8r�BBc����J:��u�w$������,^(D��Z���2}*f)��zN�E^��ށUb��,��b���pu�e�n���o�m�^�a{���?quO'�>�~���>���(ڦÃK�(6I$����>��^���蘯���O��Ky�z�����\.ա)j�t�Ĺ�4�V�6��I�ƥ�D��5%�T@0x��F�����Y���a���������&�>P�
rL�����������&���-kA����I-����4�5����Ѳ�C��c��a~$�k{m�6��$=cX��#X ��N慯
�t�kP�����ѿ(*�����R��x*���> I"���/���AʓF ������o��Ϫ9����ѡ����_�̳aO�J�#Mְ���VX��:X����m�&�~�s��y>��c� ��K��G�7�c+�٨(��R�.,p��W��*��R�w�Չu�'I;����J��@�X��z/R����m
ϙb0�h_� ���"	6��ⶌ�c�r��z�jn۱�l3�_�!d��C�ۿ�x��2�\�{#��HKU ������`ذ�벯�>�<�2#�@�GR�r�f���jl�o���f�In���b����������̢
��~���e��k5:w�D�i�w���P�Q �>sDg�Hi��ANҊe�l]���@bdF$�s��8*?ڰ}�4�k�r�	Z���7� ҫ����3و�7�M|�L�5�F6���<(Ah��D�~��?@�!�z�
�b��� ����
N%�z���tE����'l;Oq:H_�]��OJ~J*BB�.(�6^�*��R�+�-N7�6=q:�d�H�\}NL�L��^���G	���Ի�d<?.���l�N���6�I
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6tffw3MM���7E�;R;��Zэ���2Qn�懙��D�����*�8��P��cO� �8��s�礎V�t鋜���]�oG�|�w,�#��w��rH=�ϵݣQ�X��՗��N"<��q�B]�=2\f����2���ϖ����	�^�h�o+r�/i�`wP��/(�U������Q�g�O8f�Υ0�U����b��Hf!y)�2\���]y3ЛFy�Z�
�$"�X!Γ�8�O�,s��ڷ��\�E��rkӊ�:<H�����8�n1��[�>�4A쬘@�#=�0@�T�ԉ3�\��M�"��M�}+��G߅��MT)�r������(<��r�m]�.�3�@7�.+(@}���JJIU��q������4�H*՝�|h�Oۥ3��CMjh��_�1=�)� ������h�#��:�kK4��V�JV�!d/x��D<���f�Y(�d��*7����b/�D��i�o��V�i�����u�o��~ꐖ�u�ٗ��m	2��;�,r'�����V����.���,��<v�����7A6ݟ8�Q��ro�s�;� ΝO��<�W�z���+OVJ��EA{El����H|�8ڇ���,��F@���w����	I,�ČM��ur��*������������	y*���>��4�$��{�K�v	�Ƽf�#�@1+
��
Ŵ���"��)#e10,?�4�#�� S�]{\A�r���W/��L�@ߕ����IH��coAm�n��mt%��v��/uc��ߍ;I��P�O�u<o�ߣ���e�R��T�k�`o |�����h���sB���UtE��՟l�<��D� V�������u��f�s��8��~��\��7�H8��ݍ��ǡv�����h���-f��5�������ۭ<��/��8��w@�H�?�b����.12����;g���d+�7U@-x�`��ОK�95�V��'n&S�SU��c�ٜf�/�GPQ�b�Q�(��']lv�0�I)��dΪؘu�_4�".e�g��Z�����"�i����[���"I947:��G��� d&x�S�6Y�)���� ��kZ����<��|S2`���K��mj[`��c��ǡ`yw��ҍ5*?����J����gj����?juŜMy:������n�in=�Z�:�9?yziJ��:�HyV)j��,g�zi^N O)��Ďz��F{�-���Pɍ��u�+��,���ml��g�{��:��7�jg92Y%����wTc��qt�U�%��i��9fF�9񁱇���u��4Z�J�=ޣKCf}�K����t�U^؁"���������Il�}��eK[�
.��RS��x`���wV�q%P�n��Cy�u��8�^1�/��4��"X�������u��Ѫ5g��c����=?W0��E C�H���(L�$�M��^��˫���Ǵ̼RҪ�hNV	*�R�G�����"?K|��QGֵ��%b>k���/���L��d��w��ݣ���r�d�E�����w�V���6n����g�!���3l8�ދ�nBֳcp���v�6+���j���/�T�~V�j~��t�B��k���P� ySi3�ݙ\Bܪu�u��f@��-IҟȞst=��Tc��� 
��\1a0^^������eA�wI��O�(A�"�j��E���r?� ���Q[�r��eo�I�%z�F�iR ��JaD����K���5�����wM�k��U^}�f�b�=���A�D�������l����N���5<G�|3s����f���kI��7VH6��F�Xa,�
��׳�BsT{J*df4pP����m���&������e�-i��,b!�D���E$�4BǶ#�Y����>r��;_Co�B^���.Ů{9���W�bK\A&`������l큫#ɭM�7��V)��7R�7H��$T*_�?�>�L�:Ԕt1�i׼�s��I�7�	sOq��W��!�+�O+9��l�#�����Z����آS<�F��2 ��P�,4D؞Z�6)�(�7�
n�6�E��r�N��$�f&G�ͧ׺RG�\A��U���%�K�x$��N��uH&���q3��kr}��܁&��M*�#>��ܬ��t�؝)��� !��" ~��g����k�<\�c�,'5�M&�2�K5J�Z"a��-��&�z*m�!���Ո����fs!�,a���`�ϱTҮ�V��<c��߁B�6.$8�)@Fg�~��Aci�M_�;�y]U9T\y�u��KQ�_�4���qĒ�_�M���|&�A9�̤;��֚�K�JKJ���~�ߟ����{σ0Ĳ��'}��k��	�Mj#�N\Ym֦X���}�ȵ�t7H��[�G[)�ʰ�4L�*9�<�@�eL�Jr�k�"�Z0ƃk�m?B�q�%(�F�圊�_��>���9�����,��kbs��{�6 q�.�ʁ�n�x�Z��!�����I�ǪNߪ�����u4#�Y��dL�d@*����5l��&�,:ؒu�Sl�����-���������#Mi�{S��ܹy�����WF�:�Tk�+3�����#*Y��0ֶ��"_�8�z��K�ǚ�7U��he�,`�����F����uZ�"{�s�Dq,��m'��::�rW��m�ޔy҅1e��x��°*�~]�@-�� �F$6#Lͱ6jZ�&��Ғ������=����z!�Ñ��@�YpXe�N�7�K�=�݁}{?��ni�v�&������p�.B�4З�$�qf����`0�Aa~�P^K��>�qڜA��E��0�)Kl\�d9:�;�?)q�X�f]����m������:�"?���pˢ~��)n�l�1�֒!�$��mcY aH~{�b`�x��)��(�":hf7��4���*�jp+��C�Y�YN]"錙���g/]��Yz�{�)%�F��hX�t���T���]��5�}&+�������{�|�ӭB���i��X��Y���U~'_�l^�`�n3�X����m��6P� mEݛw�Y��Ȧu����_-I��*׭��GT�m_ �{8�F��\��S�}a]s&&h'
U_��0�*5@��ߤ�
�f��h?��b�a �`��&�ٿkn���PE�{��j5��O��t��ml�9d�Q}�$�9��%KfdL�gj�nM�2+�\Y/6�*� N?~���=��\r0�һSX/����Bv��"Xo��.�}y�<pa�麃uš�_��D��Mm�:0t8�|����8I�]���� A/5�#h�֭{�7�u��4zD�����e�aA"��}:�����ִ��S��3	�uP�Ձu���n,���%�퀾�y
��K�Z�`+��((k�L�;ڗ����aYCk�s�"2��@#���[�*Fb���fܶu���\��90�@\5hy'=F�ٺ��L\�#癅�lR�7�Ձt�h��ϼ엫����J�����aB�<V�w����$l����C�� H/g�BZ�O� �e%G{ݢ��d]V�A�EL�y�d:�į�[��g�(-E��#��l�����%;z��w{���s�T��`�{XyE�t_���X�+�����4T͇��8e�9(��v!�C�HC��㧟��
����"
���X
B��\�M8���~Q#�U����{ �jjߟ5?]�ù9�8[_^���ӿ[��9M����2�Q^������s�̔ݴ$�Ot��L��#��hg�����_x��8z���i�s�'��� p�k�Xp�7]�ltq���G)��V���_�~�͸=dC]���V.MPt�!�9���{S� L�aJ�
��\��8��b�����ER_��FM����|�z��;�恢Qp��N�R��e���P��k�_��y��h�c�A�[n^;X�_��^�#���1'��h��g��CS��}$��j��3}���'����C�����܃c�-P������hp~2ZN9��\��mc��3�^�a����h`H����P9�8ܜ�E��X��ɹ�ħV���xL�(��4����m͟):��ِ�R��m�����P/?�G$��
�@b���v��ݨ} ���k c�m���F=���uEW@�B<��T2In��R�5L�l��N�0҂��k��p��a�M�K���[(�AM#�H�b�u�&K�i���+c������?�1���u��L��y��`m_�+&��o�s���`�R'�%D��ֳ&8��e|*�*�|�t��!�	�U�@�84�Ǐ�,é�IPw�FI�Lc>{�֓Y4rLsb�Yr�H����q�/��a���GްE��|����ƘU
ix�#��9u���� �
?B�df�p���l>�����_���$ן(���� �X�����G�{Y���b�Mw�#�C�ߝ�Y�XY�|�W~�J҈��Ă�����9
�1��%�a�OD|ihVM> d��E`â�4���6F��P�d����S�[�����b~�7�-�JN�8���/	M �9��Ȓ�-s�	�����A,^(�T3	ݞ��[<ަd�0T*��W��&.K��}M���?|���K�	��Eu�My�`d�s8	xo��S���$�]�h��'X���)[!�>���3
/+x�� L��5���ݡ�v�8.r�z�m{NiN�B��6n�|�ռ��P�n���F��)E� *ql4�:���IYBo��$����0X��r쿕Y���|bj_� Iq˚��.��?�alSi.�ˠ	�E6�V��O��Fc&���y�̮����H`a��a�q�6�BX��tO���=j�w ʭw��w[���oM�7,F�+��p��V�a�[3�Z���f�q����=��&u��jd������8��t������ړ%���j��(8����.jS��3�pT6۴Q��2��������<y�h"��i��@Kv�4��Ȉ��qK��ePOϘ���D�:;qTZx��`��!���JR�|�K��B���5��E0��OӋ�I՝���2��)0f�c�I[���� (�d߄���e��UG�=�3��Xuw?\i�NU5�.b(7��א�+LR2oz���.�/Vh�� G���^YQ��h�a��4D����XS������ z�L�O>��0:�/�:��k��*=�{��3Y\�1X����ϋѺ�ۂ�Y	��~w�|�>�v�1��.a�H���{��z9�R�l�$���x[S�>x��7�����������M��7,kܛAZ(Oɀ�Di'��R��Ѿ2ݲoc{�Z���w`=�nG��|��իh��/��~"���� �F�.�;���Y�e*z)~�Ԥg��~q�W�"J��5sL�d����a�����/��i Ģx�B�p(����u|�ޘJ�M$B3V`��T��K����B0�� n�N�	T�\��|�OY���ɓ�����ɾ(��ǳC�x�bnzd�B͝�>P�&��<L(�4;
��ad��>@6�-��y�e���e�[;��N;m���:��p&#����RJ�G�f�{:�`�v��;(�TI��� ���4� ?�S�����x���������5���+�'k��T
�M�PP&K��p��*�c%���V�7my��a�u�,EMʋf��a�f*�loCǹ3}�fE.\��%��g��.N�s�=b���i+V����}`@�p�紽l3W�߫L���Ǎ�kD�p]���I��L���'�����`�!U�:���<s��J+@ϡPpkY�����Mo�EfJ&��EJM�]��wD��kmx�����˄�q�-�Zx#��'�la����	�9��esڅ��IOzWE��io��1'�(O5}�H�4[�=�u�$�m��%,���k
  �������t������ �R�.����gn
�Lxk�����B�AS��%g�cy�F �!j淥�&�+,�Ƅs�L�(��Ӽ��b�؎���e�ǿ�n�B��R��TZW`|
��K�k=��h�[8YC�P�'8���&t.n����Ѥ�hϬ���_��Ѓ'H�Yu�Z�跻&�8�aff��@�;Gad�z��1�2Y�Y̙�6�|j��_��5P�
_�=�z�Ù�'yC亡$�R N����P��kN�!���> �&��}�kV�47���ė�5��
�
J�������{�5�-���)�@r�ap���!��9t� �H8��c�0y��Ă�H��2]���h'a������ ,��� �����l���꿜���r�_����Q�|�A�T�XχǦCgo3H$�`8%�P�GZ5\4���d/���`\;E��n����HW�l�C Lw�?�Bj��_��ɛ͊���.! ͢���o�@���s�#�~{�e��(-�A��;�"�*c�f!�T�����,m��. d�6�U:�~�������z˧���7b��M�����K`��!e�n8���\��O-�j&��]O{�Z ��_�V�	J����5�6���� Suc�#���[�:a��Ra�DT��\�{�Q�tx�u$�7o����>�o����\@�y�Ƌ�:��hm�����$�̎Ѳv?8��o
�c^z�>������%G��v5��w��h6��.kTm�]6�ښ�}rEӄ	L;6��zTLu �U_��+�*���<Wv�N�JO����|������2�2I��I�j
��bs��!Q�d.f�?��a�P�d����οa����Y���n�@C�D+y�G�`:�[���wi�?�_�� gYh+�xi:0%�5�I���%�\z(�N3�!<�r8L�?D֠޻��q�����6�~.<���v�ގ�g���Y��3�`m���13�7�Po��t�:O���c2�i�n��}��*���80�;|C̖S��0ܵ�L�SY��;OHazJX$U� &��r�F�ub�w*�?�)�� chZe�o���_���.�$�[�o�]0?˽�O�IӢ�������A�\Df���W!�� �g.|�pm��2{F�Ω\�����k�������!���i��YХ�>4ÐД��`��v뷎7K�Ձ>4� �������j���Kȣ�;g�h��%*��-�3u��Bh���%?pI�<M�5��AY'%�~��ڒJ�e�_��NKXd��N�a>|��<-��ӹ�d:�?�;�'�	��F�3�"�L��[�(����!�O�A���+ё�g;�&Tr))�ĺ�3��@���4e>��P*t"@�
�SH�-^
�oķ�g��QWv'~A�Ƞ���ђ�zs�������/U� �x��W�JsLB�L�tk�yIs��W���3�@��c��I^�����<�s��Ir�������D��\��D�X�Q_�|�\�h'\�t6B���cQ�b�����֑�}�~�L�0��g��s���	4{ߌW}�c���CfH#��<$����E�DF�mQOjǥ�B�����j#�]�
uv�ù���'�s�5��+%?�RbĬ��T�� ������ǫ�d)�����븽nE����5B�~˘o�Q�;
}6���Y�x�p#~;D��^�?�M�kD�k�Br��jI(d&��@�%ON{�wWHY^�Ӈ:�氐ߪ���4O䦅��Z	�`_D����J�zl��Ҵ"�ek�/v�E}t��bv��+>����1_��D��&��?�)J��kҗ����j	�p_��dc��V��lշ����w�K&��ch-������%���~!����؊�Nھ�F���ۢI��?�x�ټ�v�
e���� �$�@�E&�	�uQ/Y@�k� �bW�Z�C�-pxrO%c$H�#��âT���Y�ҟe��������0TQ��u���ٰ�`����Β���bʱd3��-��n�p��P^�E��wŌA
kRɄ���~-jk�va����;�^�8�j�ͅ���&��2�S�q���u��1[���L��1���/�|_^(���9�T���b#�^���5��o��8P�3��c�!�8}hI�8L`6 �GV7u��)�N�vu�;8x,�͆���*�X�K"�}��&�15z��*�sQw���%QF��7j�l���5� �-<��z�'j\L�7E&D��S�p�%�����q�._���>��xZ@���Tŝ�J� �CO�p:A��@+s�l��mp�4Ag"3d��Nj�̐o�]J!{҉�߷<���o{��99Ϋ>:�l�<��o��I�+p�-�OI�I����df$Y�	�?�Y��b�zv��lF|�����P�,�Ҝq� l�l��ȍ7)Y/����?7o�aq|i]�3g�ԝ�l0��H]�axzY�Ib/;�8a��q��	C���0iĒYتe�ڀ�̯(:ꢂ�U�LH����%$~��H�B���=2|&Eܦ�t=[	N��uC��H]����<t�Kɹ�Q�9����o���M���*�
J��!���Y�f��ly��U�z�_���z�bx��ڂ����Qe[� Xbj�# [����E7>Lz!�s���譭��J}>g��wɢa����J�b��HbҞ��j;��7���:�4�0V�v3.U���Z�����]Z��I}3Gy_���d��I~o_�l4(�l���h�'��n��nf����(�;W;uuMg��ZnMʿ	o����*K7��E�;��a~��;�?4���!	�����qu2�����H�y��V��Q� J$��LA��v��0�������h��3&+������"W�k]e=H���i��^nb���sx���Dw�Y'%�m__/�ctd�N��L�5U�tLt��zIFfc@�zp�#m-F�Sn����T�����|�3�d.��_��a�w&"k���2�q9Rȯ�L��1�h
7E���{�UMa�i��Io�dj+r�dy ����m��wХF���ܺ�@u'
'h��oD`l�-��\
(�������1��A<�P(�V	��u���P�bG3cಇ1Õ�*�����l.�7J��A{+���A����G!<Ԝ�ɔa6Lʶ
��K;NrCZ�b�`>v��������o{�h���O�ᐗ����Kj�=���a#�^�[�6Û|:'M�F�s�xT�Ipz;q�e�̣1���}@�����9�wx8��5��f]��,;?���ex�6fg��N�fRC������W �d)'!���OK>Rӏ��d����۪75�tC�˥)+FRf�`��^�F����"}�e�����y�!�a3@2ve���Y,�B"e�-Ϫ����&��L$v<��$�(���9_�p��Ն������2�g�>5}���ΈA���0��7ܔ������Ko���f��58��Nȴ����49��P3 ���#"�r��2Ί��� 1`
�/�7<3>W�1�W�N�݊%_���m?v9odN��f7ſ��v����sB�
�)�K���i���o�`�i��[�kh�2}�VSx��5C "r�)qc�'�MJ��H�5K{��X��<^2�M���DAY� ֭�v����`�r��qs`�n��!y���z�r�ac��a��2��bg��ms��w�\�����63��� �§���8�s㘦�U��ǖmN1z��]%0�T]Q�c�x����P��'6�p,��gb#���'�=�\�nI^Qfxr���2��p�^`zP��t�ߙ������z�1��C2�������cKg�Ip{�ZC�॒�M�&d	z+^��^L@�����-[bc��yg���=����c�5��Z�ʱ���>Y�3Ac�^ϞW��z� ���/dU��������g���:$^j>�ic'E2ŋ�\���t(��`]�����;̙�D!3�B�c�0��HY�MDL�ȭF�r��m�u��7�ڑ4ߧ���n�g%-.������3˥�T��;�ջu�dw�wt�����Q�ç<���n��@�[�yS� �%��ha��;��Wř�/Ҩ���M�z�M=)'�G��r��d\A¸!:�����D+� ?y%�$-�b�����:.⫔��B6��@j���� �'��w���|m�\�M�/v�{E�c�\?�؇�?_����'
�Z9K�Q+�L�9���֓h���]I⏈P:���<���P�%q�:�W`w�v��k �O����l���v���2���� Fݐ��I���a���u!V_�҅[Lw羝��m][�oO���Q[�D�M&��_�jO�d7�9:��,+ô�f�K�؜L�����G����Aю�]���.hlY�z���]�Yp懮�p�x�k��S?�^F�0R �4���\Uk��fq�f n���Mn�mp=�Ug&\���`��ko��Y���x�z��+�Q��5�_���܆?t�.���ɀ�UG���Հ[���w|����V�)�ۯ5N辶�"
����y��B��-��%n�Xё�m!��G�*�j�S'���](�>��&͒��/_�C�ZʟR�˲�۸{F�^]�&F�J6ç˽��|�9����&}�������ůJ�AW������H����T��u�R�rG�A\���+���h�1z�hM �G�4��,�/A�P�Ɓ�{�J�L�3�4�'\�@7��z>�r�pŲ��4�/��9�T(�Y]i�)%��W%��N �<�nQ��S1�=y� O�y�+�O����銡ϳ,�9=�7+�n�o�k���:7?���<Cݥ>`IK��Ì�t�$�<�;�׻n�(��VH��/g�K{�h���f�_�ԗ�i������������w��w�%pvXߌ���NN���A.ł���gLT[��G���;�QN"�Q�s9����;� �� 6X�}�E��=�ny�Ӭ��&\ �"/����C���ɡ��KõJ�KZ.�P�2��wH��p���!4XM�V�V�<$/�4UZ���T�?�K �]��q������]8-�:`FA쇟q�l��]	��Op3�>��mtfWיI�,��GD[RեϤӞ{���,��\�uǝ�Ӂ�˻�J������M�w1�2�:8� ��W�h"�Z���q(zl� �Yx�s��' m��\����O�E�1B`�O=���k'<�K� ��A��5�-��.��=.Z��;�y��Pڻ����1b�"+l���4�s�0O�\��3����1��~f���r���J0>fW��Pe�<q�E��x�ys:�k�G'��N;HU_P���R�j(�]�,s27�%,��3��.��
 8T��jH��*P��j;�����|\h���G��q�ƔD��U�A��I� ��~c���D��g�h�,��!�A 4�kY�#T:O�CI&�� �[`[��:����>)]�`;I�4���+�eJR\�2��WJ����\�ꭐ����w�_�jG��e-�|#��U�v������j�
�ҵ?1��o~B��g�M�8���o�E�7dA��t�K�f|�JJ�)g6Х�F�ba��OI��y��|�[�?�f�+$�̙����|:9��k ���K3�{7�C, s5��_i���h��W�M�>_�ÉŖد�̫��T��% �%eЋ]��[	�Pﾴ9��j���Ou���\��7��)�,�s�u�7���<tv�T�M��AR���v��tpk��X��x�G`��K�0TE� �Ŝ�g�6��K��M-�\Ymq��� j��L�*�8�UL:"���g}��A	���T���p�������a�́�\�:R/��I���a��iN)
k˦)�>f4r%�^���Z������Q��#�]�'�/+��?�V�k�W������h&�dc���p�j
�>خ���<�6J�>�q���Y�Qn%���][��ys��āO��?䤰�8aX��a��^^P����o&�U�H9��F>,8�3��m�3�V2��*��U7�Ē.��m�|0�1�#��;Jn�g�w-&�.��˸qGN�V��ָ��!��2�!{|ܛv�����w���,|d��:��#��z�3f���! ��>Nm���x�0�WmF߹�	��Pg��	���m�F��W����6�� �m��|�K�����/}�FN[d d͸�X��8��� �AP	*���1�,�����+�q���	e��ςvꩼ6�	өȖ��5 ��?F;m7U�4����E���@ȡ���6û"���K�Y �����2���纐�~oߝr��:�V]��_��T5��i	�}z��:�`2�#����hR������_�.댛�H�PպB`��U-�,�#�SW�TC�����I!7MX t��k��(�,��Ha�z$gY�k��VT�L)]���'����L}죏ܦ��	q*ef(\�ݚ�[#�홢E]�h=S,��ϓ\��yJ�q��Uq^���p��ڻ��j:�jV�����a*5׍�!⹮��g�WF�� l<��j�a dUm��P� �F4��Uh'츧�k"oGdͬ�{�7�O<�:7��,�Ͷ�����	C�U�#$��ږ���T5s=��ii!n�Q�И�Gݸ}��Y��w��uqά���Y�L�c>��ꙭK}J�"i>��_��+�Q����Cpj��s1�T�Fh�ǹf�C��k 0�PUf!�a�S|�S�d�
g�
�(��Di��k�� A�e�l�'�	5R���G�L/}KE,���~�����EB�Z��ۖ�C)��o6K����~,��?�OÜ�Y��y�تh\����R��O\����x��1�I��k)W5 X�^k7�3�`"��RI�b��m�[�A��xX�9����B�|T��,f�t�
����v^������sƙ`��	L�NUU����TsٯEKG=E�ćvN�bp{�ׄ��w����ye"
��3p�E�䆆+5�_Fǐ#�+�Ќ�[�������9Յ�	)>�1H�i>��@D	�����b���1�N�er�F� ���	4@x�t /���O�Z ��R�s����
W��|,��[��<���*ۃ��a�X��*P��SZЄ�)T�vSX�i��r�U����ʁ7�����3�7B�}ͽ./N�/M2��T�,$q�BD߯�c]�g��@�lAeP��9@)���I��]Z<e:����&���|�\�ߐv���(�I�'�u�C�9����M�E_E[�g���r��4���fj^�U;Q�N���牒�Ǘ�.����Sc���<4C}=�5�)[O1����X������t� ���������O$� @4�$����Vwu�c�����Uӎԙ��|�x�ZB@�u6'�^�MWM��[��Ŧ�1��1H]�q4�÷狷��ɰ�E�ֈ��4��Ƣ�ȿ6k�v� �YAS�����ћs����t�ҵX��I�z����
������>�D�S��_ H���燞��'��>�ynG
<��+<�đ(6��T'��J�
6n>�A���ޤzݑ�ڶ���kXr���U��r�n�Gt������|K����ȧwS�5IOãH�2�Ԕ!�1���-3�~k��x��W��)¾Jq��x#�� 7�ߟ_s�L����I���c%�G������[%v=͗�#a+oK�lsb��v'�?y8_:��WQY�?�Pa��Cs&qpM����]��'qLzK�����%&��F�B��-X6U^��=b��l�F��	�S�:�������(����W��r��I尵(�o|+%�x�p�K��0��wv�s ���#�Fz�eS+�	��F�Q����)AUѥ��x҃��˔^=�-B�C�.�JP�Uy%�"�ذ����]�ͪPјN�����:f��cy�(�"�?�5�(�i:�ؕ��ѣI �`1��Z��#�-t���&h���<�v�k�g�׬���kߑ�m*��vD�k�tb��0��Q�˨���]e�u��$��_�.a��~лi~2�,a���Gh[��c��n4?b��.��2�t��T�N�Z8�LN�d�z����|/i�,l��M*.�k�D�G6����3��w�ت���R��"RjQ���7�n�dcWe��2��D�bD���d��%j�VT���فG�0AO��U��.�7��Z
�Vd� a�q��6Q�eN/L���3�P�np��	�]��Z��M+�hW����<�ڑ)�@�׃PF�w,/Ŀ"���@��& $!��j-�ٕ�D���i����3�`�i�����$�]�Z��;�MI;�Sf]��LnI%�&] �X���`�	|w3�������nPk(��
���|�^J�J1� r�)�	'���f���[k	D.n�![���2>�#�k�����?Z�¹����ug��-��i���x��X۽N������������)�r���^��_�/��c�6��Ԣ�z%M�z�0��D��յ�8G<�{�U4�I��АɌ)7'7g�[3.�r$�̼F�_VQ�Edf��X�3�K$C%K�4�`#^�6D�)�v�}��R�9W��
i����(&	��("���N�Y1l��XR~��	�sMfZ�M d�EP\4b(�/�5ȸ���.�L����W��r����捷P��(1��&��Z1�F���S�>A�g�N\t?�E♦O��i�����У�g���&��ٯ~���pۮ�!�<��iz�Q�!��r�#X�K��{��J�_3$���;�]�5*��\cw��� q�J� '��(y�]a�t%�E�au������n�/��V���v��6 =�����P��N]��T��%�=�T���w~k��t?;2�"Ը!�P��%Mo����w�8���hi��*Q{�!Z?�]GtS���u�f�������/�|�����b�M�3T�_\�����3*����j'+����0���a��#ݑ�i����Z��+��Ja�(3��Ϳ�8ȏP��z1,�"ύ����q�u�VhaR��d��N���ɞ6��L1��xXX��-���I��bw�X�!��5�	o��rW���9��^?��#�EI-�^�$�~��d�����m�u����𬐦���"��4b��d��tb54���H{-cc鉽9�pA`Ɨ�i�EAk՘~7<3	^�N3�".�����I2��>��ǲ��V��-�8Ak���v�x����#����M��@��tU����$~�� b�O���n�?�I��O�-ø�(�R��p���]��:���sL�*R��is�#�����@��<���b:w[x`�ǐĦz[�/���M��ߘ�2�MW�~�=|�vo��kǈ�?��f�Em��l6�h"T�h&4�T�^�=K�Ϩ���c?��T��#��a���[d�@ ��l�U�;��М�7Ib�c�ݩ������"
�B��M9�z��'�^��8�Ybc�l�0R���¦ID4�)P#�%����{����JG��U�M��𷙋��C��؋��R>�#A�q�kwJBT=���>\�vVJ����'�Y�����6Y&�5�(GK{�5w��-�&A��78�P�Yg�z�-Q�ǅR�d�h���A|)m[h��8`�F��T���_��N��Y�6��q���������o���0Ҷ��Ģ�.�Dj�H�����"���5[5���8��vC�����l�}� ��%�Nޠ�;:�5�d�{7p��Z+0w?h�f㜸up&��þ��3�K���EB1� ��og�;C&E�Y�ݙK���wh-X&1�~���ҕ���ʆ9U���LpS,�NH�U��� ]�_!����ƈ�ǿ�&�4�V����-:_�)qE@(�,��;ѥK�RU�fgD��Dfcᜫ}Y���U�mbIQ���yz��s����M.�s�*$eu�x:+2�#����Y"q�	Z�����]� ��#?+SVqn��@��nƮd�p7km7t=�r\_�Y~4����8�H�,ݽA�GFo�l��Q��Bw���a�����	��z���_�j�[&5��6	�~E��2�Rs37�T��q	�gU�&~ ��x$R��dQ1E���@��5�n�a��σ��E�\�6aF�-�'j�)70y���D
g4��;هh	n���t	�o����(��(�M�*�� Lr<˿����:�ޏ�g���5*p_�A�%�k��P�=K2n����.���_�K7y�. �sC?��F���^wqܥ�D��$�&�
���%j�D�i�S4��7��e�秝uu��ٛ?�h��
B�����ά���l�h7�U�[:�ٿޥ��RZE7�?fS���k���TH~�LI��'Ki܃�먕+H��ǭ	'cX���d��wà�q����zj�����0�	�o�.k��S����Ͳ��Zk�VL7�"�7? 0O�o��mJ�=4�an|E�A�:��!Sa�mt�B�X/�Z����Yҩz�7����!5��[W�ڭ�{��;W��ܶ�9P�8D̞ykZ���  ���`oA������)������n��V�vV�%p�� oQ�M`�����0de��� ����Jh/�7ޖ�M��dil� �3;F��@ߪ�v {�wg�L, nW�`�e�cH�e���N�J�g���E���d�}#�#'��QVgI�������S΃Y-��Mˢ�j�Nw�@��QD+�ĩ��S�!�+{ӈ�ǩ�!rS�-��^v�1��0ëo�'��?{�R�Q�I��@!�Ͻm��"c>�_�DK�1�#7v�aᴯo�X�i�F6C܎Do�t�$�����z)�|Ħ4U=ǼJ�?�:�;���
Ƕu��j�/���u�@P!p�U�l�&,{���N|b}�`�`���Ov�3w���L&����#�xHB� wuA@��ڠ�G�y�gZې���#f��nu�t���ZV�S��S;W���;��=O�1-�haO��K�����E�i�bI���7���gEa�-���2�s�]���&�LvDm&)<rY�`��"��s�X�}p�:c�lxR=l��8p	�:	��p��-�> 9��*Hz5 ;h����1P[�`���IO_�����,��]PZ3�Sq7VAn%�ĉ�s�b"�4l0�bPL�z�]�q����4|���l �D?"Q8���Unt��FJQZ�ԡ$�@_ \�|A9�T[��n���Cc�p���T�wz�N͉������u�K�p �d��T��ѝ�M���
�̒��9�r��"^���;�iS7�<���'3z\�=�ia�g1zh�vODAQ=��o�*��h	h�-���v"�8�l�U���!�[�y�n&Z�-�����AoT���_6辴���d[��u�E!�7�M�*�g�֧��IlS��c���0<d|�*�C&�"���/|'�τe�]��852���2K���&K�!���Y��d�ϣ ��-V�� �O�/,��ͭ��s�� i8��@���܃�=p���R��P%ý�UB���O�Y��'���НWR����kDǘ��_=������(�����2�O!�8bQ�J-�`vAӒ;˵C��=�,�	p>~���:�R:�=SL�~����º��zC�1�f]�P� ��W+oLp'>��A _��H+'�l��c�Nkd0��:�߬�I85I��@u�$iG�Ļy���xD֑�l�S��W�}B¿Q�aco9�Kq���fs�}�D�T%
��5 ��O��6��(3�˴�-A��������'C�G�eq��!V�m_�Iw�WN�F'һ����Dm^ԋr��0u*��
i1B���Ovh�Fg�A|D���U�"�"-W �m��� ����Z0
��yz7�<�,z}���Y�'���ށ,lw�~QØ��	�ɦկ{?��]+͐<8��,�������堢Ẏ\J-Y�P��J����� ��-_�$G$XO�ч>�����l5�HB�7)���	.��`�D�ؔƅ������~
���= 5�����q�qUK��}< A�4���~�bY�:#���l�-ϪkԼG��ܧ�ԀWSB���*5�K�ֻ +?�XD���T�i.��G��?������Q+�3���>�.���t~��vtٍ�q���GV�׊�����}��l�.����\(�®�׍���C ���������v*�dk�ζ��rgiq�ە�
cӟ^�aގ��A�jP�Ϣ�ػ�cŊ�o���L�ڎO��G���'��`=#�q~���/�0�q�t乶��TItTUެ�h +��f ��.ˎ�Ę��5;[-�J�3�^n�ٱsV�S�+`�ROq�]~j_��a��O���B]��x���l�Ęd6O�ʧ(*�i_�Fn[�$g����#��Ѿ�9S�0�l|���ޕL��"�L����l�\�ݲѺ�7�,�p�F�$�N4�P�[G��(�ү�� ?a���7��@�[b��-�����A]����z��F��/��ff5k(H e `y�ǣ|w�e$f�oK-\������*�V�N�=���ղJ�q�cYf4	���}�2 ��GŎ˒1����Է.��%>�XQ/`����f�ILo��=_�w����}���,�]�����`6
�7�g�Ψ�y~G3���[K�E�J�[�D7E�v�[�^|��&���f���$K�#�츠Xr�������D����_�s��[����_��P(a7��m�/����@xʫ�S���	��iuZ(�:�c�
��xb|���㹠rE�L7t�v@m�&���J#� �~�/[�'j,��]�Yo�+�#%����֢��.*�i{��ߣ���d�Y*�J���nDW�AL��� 	�T�q� ��7!(j5�����1!A0�g���NV�A�BQ��BESrN������)mk��9�W�v���������l0w1Br_(��`)��H��)Vv]�p�,V/~�����C�F������˗ŋ���ҒIje�ڰ��::�v��>����(j�^��^w�c��/'�V��.é�4�"7ڝ��z�z  Q_�R�p^���-<��>�}���M��Mo�-�	���u@`9��Y��H��Za�/�@fL�ɳ� ���Eؖ�`�����6#��6x�z<ah�v�w����"g?����v��f�k�u�b�n^=����Է~P{��RK쵊����`5����L2�[��#��%H� ���C��v�����7�+;[�s.�ZZIs��}C��s���C���װ4=����� s��0�pE�����*TF�)5<�KQ��\!ا̄���g�xǷL󍱫��@�������c8��x�5�)����J����I�ѧ"2���Zsj톣,t��p�
l�jc-�|q9h7�!��q�j�wCM����m�x)�61鵔�TF��:�d�
)���:z���0�Ě�/!I����M}2����U�,�)�������tş�P��K2zR���[?]�M�0��+,�c�PM�}{���S=D��\7�����b(�E�X�m=27Vwu���t[�ʷ�ꄄ^��>z���Q���E>�x�Q��|7�	�p�i۽-y5��5h(��������6�/ZQKV�0��A/TBj|ٸ^��i�(*!8.\x�
�ms��ZD��w�wҠh�ptN�]K����I؏4��rH�dp�(� \�	�3z�jV���a_]�������j>�䓉%~�g���'�PMqw�jyz�FK�	����D.4{T�� �S���I�����m��T ���G�G��OϖHk��
AtX{xQ2X�;8ʙ�k����w@������c�d��0�F)��tK��et�s��3����F�wբ�8>2�>�ݝ�}�K.@k5L��l��`h�9h�$��R$����#���W1��M�?㴍���k� �zwz�B7*�룱-�p�q�1!yX��
���^�k���&	���_a�^��-j�/@2���G�W����E,!�}Į3�+�ֵW���ˍF�T��E��IwlP|'<���dU>��֠m!��ゖ���o�%Z��h���F��)�Մ�ղ	���絶b�䱛w�NN�(W�%���k��>�#�QU�TLcy
�
C�<Ʋ0�ĳh�<Pn0������q�ܿ�d&uO`kϔ����3��r������x�?7ݤL���H�0�n	�4�E��T]W��@m�
��f� ����C(��NҦ�sepp�&�rfJQ�D�fb&�h�S�X�c:�,��o3_��0*y߅t�e��p2�T$1��+fI�x�t�mX.�!��6CGD��o�W�Fs���(�G~&|R�>}[�f�����>����ES0Mw���*L�
M�ϕ�{�1�A[��,5�/�D�Zp��'%^j�4�ƍ�����b�V���0���+�#s�����'<���b��͖�����@twRtz귑9��t�eC��e�l���o�a*_�����Q�r���LfG��#��K���T��j���-��¶͵I����ԆއiEA
/tp�lp�w�Ӄ׊�%��C|eO��o���u�%��|0PQߠܿ�q�^!��8%�i��!l�NL���Œ@_0�=��*���Q�����+U�+�H��@�3�0=�V���6��o-�k}X��i.�IN�������l��%s+�[}G���Sq)#wq�Rv7�q�<ɴ��vC��=��$���1��l�V�Y|U\/���xcˈ'�V�E��7�!F�qU&�auW���|��K$�U���N�&�]j-G'�y�j�U;7n�<x��O�č�:�ȸ�\V �uo��;�_����[q�wIN� 3 �Tj�Ryچ��z�}�`O�Q�z�b]8�LD|J>q�F�*���3�ߧ��/�d̉Σ�"?�mnS02�e�Y�%��Gq~��>��V5��"������ڻϔOT��(]_'�ì�㺛�j�sj�V2�Z��JG�e�x�;?�W���K��t|N����'Jm��/�ۻC��a:�v��
L��i��j��C{�@«����+�q�A�3{d�I�Re�~W�A4����1B�O0Sr�N?Z[oC���i��vY��5*n��;-o�i����6X�>�wb58q��=;��yy(vu���KW���O*�	���8_�q[R�)�!�˰����}��>N'&�+�|:�F{5�u�V59χaW�?n� ��VY�Ă�[�R(Ƞ�U��t���zf��G�e4zF��Wy��^d��U�Ó�~ץ��U;��Y|�SlY�OT]@q�Cֿ��-̤�v����ťu��Ɗg{�eTmZ�<�[+�*ȍ�#�l�H1�H�������%uJ��;�eW�H���Ί����@j�K���Nq���b�������
x���.���mׄ6d[[Øv��L!]{��#îGJW�u@��1��4&�T>G��{l��H�f	<$�Mj�"�y��K�"�6�'͈C1�ˑ�l��ț�'~Ã����e�>�}h�'"%��m�x���k�y������Z㉿ti��w��':�۸e�7B+�m>�rL���@P�U]�镺ۄ.W�aq��\0�J���Zk-Y@"��J:N]���h��2ԢS'Ugu�&^`ɶ����6x��!�QVB?��
���aX�VO�n�K\iD�g���F�l�	��e�B���E(�OT�}���y�G!���~i�bǭ��
��n���4���ID�m}]I0�B@�9R
��O�U`����>Q\#=���g���	}���\����"�&���P�'����;�WRZ>�z�;��Z�7m�4 �!G߬�ߴ��Ai�p��d�%�X�Q���-pθ�x���lx�"ж���w� n9Yga�"�o�F;x��a���xQ1E���UZ#��췅Ѩ�D����5:�QQ����-%}Y�F	g���.{�S��C�L`�F�q�����A7��PI�Q'!p��C5�p����;��[��%K���K�#{�v�y��=`u�/!��Y�>��,�ɮ�'�>���ă�<��ٱ����?��0��o!��. �M����HO��0������B�P�M��EpѢ��'*�������X����A��4@�!ɀyNbvZ3�@�1��c�ǲ�N��E��-{��N�M!��R3��:�����o}�3ۃ�z�Ơ ���}�h��<3'Pr+M3�G�ջ#G]4����Ѿ���e9��Q��,9^ӇŦ�jp��-���۹sm^:L��Lb`%�p��{�$�	�&�U6���|�����d���*�׏��C��:�cB_v�-��1g�^CV,CZ[��B ���<_d�~�!��B�j����`���:[�Y0����3��!G��?�=�4�oʓ���ɰ���z�bx���܌��;ͳ���UT6�[�Ғ��.d�5��u`D�������H��;.�i� ��C�ck6��.B7:9O	��p� �+�Xc����W�$x琞:hsR���G"�?����W�$�[�Q�,�[S���~6�#ӭ*�l�"���54�P!�{��;~RKsn�"'�=
�ݱD�l�ܦ,p���_}hokͽ�OrD��w��aO�e�5S ɹ1�tN����[<�L[Ealѭ����s�x@���2a�z�nP 9tt��H����?��ĳ$��k��o�K���=���!³+�m��itp5ĢNLR���l��+��З��-�WE�2-W?i�L�%��4Q�~�knk¹�-�5ԩ�.���K�y�O�ٻ���Eӥ������_��ž�b��������6.I���� Y��E�A�����'P�Vf����s�=�G�,C("P�5��^4Ɏ�i=��D��T��ŝ��ƍ �P�|?�Uh9]�:� �����HU3�Ï��D�Q���.5������;�,�Q�(�t;��
<-t`�ʝf������*�m�i������?�t�� d��g�����d�zYBc��Q�}aɥ�&���8�2*�	�<o�ulR�����w���n����=w�~P�סa�lã[n8*�,#�[���ͯ	��I�H�e@�b<cR�y]�� ^qo�0y_(eQ�8��!R@r���K��p���3�Ł��X��7��c��0�_�o
�L�\G>�x�_ٞ�3����9y"��\�W�"���UĜL��)�S�IC=eě�;��wc��OC15x
�D
¶3�L�3�ϧ �5y����W�m��.:4��,X���̛��]��X�4+�#��zi�����%Vr0��0.@X#r���7>����E�'F�{�J~p�S��Wl5����vvM�c�`���/r�q&{KH��s�DBR��~��/����z����
�<�9�ZK�1<�oK�J�7	:����^����^���O���hәL0%��AI�Ch�Ǭ>��:Py0�1�`�O����rs����gdk��b�5���rH���g|�hh$��Ų�Y�_<�8qoQ����az�w�?>�ѽy�xX�O ��j�����2��&[q��:�%����x�^E�w@]���	��r8����y��O� K�W���5�:�b�F����y'���(�Z���Z�>6Y>��%�s��5	l�`�a�w#?+ߛ�����l��U�4��W��=,��cIaU���� .�6��D����\9�)��p�%W�'�kIO�q���U���@���:m�7�I��f���X�������Q;&;���Q}�Y��ٵ+��һ$1�h!bɻY�>��yu�ՂJ��x����A�D%��"����MUs��F���b]�̦l�ר+��l�bV��	��x��? /a��W:b�NL5 �у�ӷ\4��*%N�d�%�n6���SH�xXծ��e��l��VH3�(����g�39�}�T�/�`e�@�a�9m|9�\�K��{W>2��̈�R����� ��>Ա�����P���ayW��l��<7������Bu�C8����a��$yP12p~5nf4��e�����<C Lw0�a�9.�%�sű�~"d�����D�y�t����D$H��g�ʤ�3��ޠ���׶���p�!�ǧ�ػ�������v���y
�	�0a�͙���>��F.�a=»�d}�͜R�t��{	B���	6��ɿ�.�rK�޲�T�H����2�{q�ƞd��!|蔫�������A�G.�>I�
W��� �y!we�.�kǉRz�/.??B�S���ٹO-X$c���ȫ����*���;�gb��@Sz�l��y��������{e]�`
NF2��"\N�|�{�vZ]!<���D�ljnPVP$`$�c&~�`�ȸ �VK��C��g�^&s,+�ag��'�P�������Z(U\�G�ںŬ^@�����xr���Uǀe�S���1kh��7��`/��R؞8z�hrb���~x�_���Y�,�J<`���)xU��~o��߱�@���n�m��*#�E7\�.�����H��a5�Z�xe	�wX�8�D��)9��.s�y�m����'/O&�C�v�
>����͑��~D��@�$jJ���б �T�6)W#��P��0�$s4��%A�$5D�~���V���g��K�q<�O1S�^�*��_+���ͪ���MHEC����>�z�Dll�Jgi�ތ�23@����'�VI��/�ޗop�\�+x��t����%�H�`+����q2f{
�S��M>�����<�`~�5���.8�I��FJ��'�uhKRz��Y��E`n�r�B�S� ��*S�S�E���T��g���B���/J�F��X�l&�v�S�2]B���\�IV��=��όm����?�i��^�����������)w�L^'3�I)��f�f�K�?��Y��%1N�<o�}�n��5�����3��io��W��BϫP����G�Ɖuj��L�,V뎼�{�:.j�F�ع�y��R�W�%c3.�q�TɆ����S}�
׷4e�O���d� �U��e?i�j��q���!�os�K��=И�=W��e��FH9�!e�Z������,����MA�T	!�8�60�����72I����.]	��l~\��K,�/=�fY�+	n�Ba�����Q���t�u}0k���&��j�;R��7��M�C�ux��V�y1:�<^c�-�FFO�ؼ���v����k��1@)�����?R� akC���y��l�JS�%�k���\!�G�3�z�Y���3�$����c|BO]
S��t�N�>��G�'m��I��I�ѿ�=˜P+=��؋"�۸ٷ���/K�lF�������.݁�*3�?_�w���83�_�>���1	��N�2��%�A����W�ܕ��5�P2����(�,�{ ��_��Y	���)�FD�m�Z�"�a�6P�c�
>-B9��V�@�@�fy����@��� ⳱o�ŋ&��Z;�S�
n�N��+��P#0@�$��G��ÂA;!RRT]��A�խ�Pa��O��fU�wB?�� WsN��<��϶�b��	�K�~L4@��"�|�D]ߏ�ÑA�Dt���ۣD���/�%���<�Xs*x�����%�qq-������Ɇ�V'�CT6O�w�-�Y��}hc���D��S#s���R�p�Y�9�4b`:��O��9����d��kĹ�&<��Q��^ۻ� �1�r!�5�k��R���A�E)C'bW�g�ϨU�tR6��PVt�Ge5~&罼@����}�Z�+t��IF �k٠L�0`YZ4yH\ZT�":���ը�<�hǝ�.�-acD�b];[��w����ǩx��Χ-U�R�������q�hh���|M����*�}�rl�Ҿ5∏wf�T�|H�e�@&��h�s�*�M������e58%�%C��gwvEC6lw�^�/�־CJF?N���i��}��l"ѓ���w�~0�����+���I}���Q��.\6?�#�oH���/��`|���W/%Ƞ<��u�#�z�9Nד������ ��UW2�@�X�^zPZ�t�-����Ny�Ad�i�%��fM	��3�1�Dז��ծn�Z
���id���%����@{��͇��+�A���Q|��l��Xψ���ր�`���]��X�G�ŽL��ށ�ǁ��`5��$RA���);�7��)��;
R�i&��x�T9�G�߃pѹ�;�����p(܃���TA��ByD�'$�
0W'�`g�[��T�{Kz����J���ӳG	��L3��{)��v_t`�����T<��n&K��s���82��T} �?�oA�M��#��bUi��8<����⥍����68���+ƿ�X|Y����'�Olh�aAE�����dVz��zm�5�w]���o2'o?��_۫�:4(3�!�~���o�1'U�䳪�7�ĹS�j�T�1l˦J>Ӳ�:�ɫ���	2��=SÉ���yϿ�Gh��]{�W �;\ J���aZ@�Jex$��un?$��"
xg�R�5�W�;s[w���ޟVƃ|�l����Αכ��J�bde�l�_b��� �R:�@|��q�+��{��ln�ajݥ'�&1��dU�q]g~L�Z�X"�+�n���9���������L@6l{�qd
@[����⨇�����~�C�G�=S�������-ZK���z<6�j۝W�9��1��u0��X򔸑ܜ�y��$l���+,����V�Jn���eZ�}pWc��i��c������t5ب��j�k��P�,�?�.*i�h�dE���M��p�+�G3�X�r%���f�D?�ʧ�R��P����uِ� �V�&:�rԒԉ
�ԃ����(9��Ga�>bq�
�c�}d�ث(@b�y����5ְ��I:��k'=����_�l��5�t}�_�'O�X P��p6jI�N
���q�객|\�C�1��^]T/��ؗp�״Q{@�":/f�v[�4���. ^DR*��&Puff�E���rjp��4V���4E��%��tT�,��Mڦ�XK�����Cw�)���-	�R����W���/�~Ab����7���A�X�}��~���E�n��Q�Xn/]�1����.���uU�:L���k����4�għ��;�oJ��{
_��^�T�ks�{ɭ���"˳��#T �� ��7��B���i����Ɣ��2��cQl�M�s,�dª
����U�6sM���4������Lq��c��T(f>.�B��Py�����ԉ޸$��z�����܏j�"�����ϫ�g���u,��T��i���Lܤ�&Ui��[C��~#钎L)}�,�9�_�)�3��)��1(��B������bc�<�c����5��^p��_�(����g��W�g�U���%�M�Σ�M|8�g�w��y?���R�ؠ���F�]l��@N��)1�WTu��80�9pt���Ua�Ӌd�4�$�/�z4�����hh�AR�<�쾻�GE�
խ�XO�|�P"���u��U�d�1a�d�4��7��S���d�������W�7|4��ko�V��y��fB�����G��ش�5鲛P�G1��W~<�3�w�`hy�`��\j��4f�o/��P�S���2ߞ��qɬU]n�F�0�q�3�>dn9�$�lյ���D;|7'��/m��R�Y]Y���]��.��y�O8p� �M�{]��PC����@���բ�X��'��}��5+o�*��-�6ϸ`a���Q�Mj�ߞj+�ɳh��u��� �ꥱ3ud�)=��I���k ���GS!fM�a������c x� Ȫ�LSZ%Un��g���{�X���zA�B(�8"@c��ە?H��ʵ`%}��0�$�.acD߱U��1�v�8���$��B�(7��p���\8���.U�끦�#��XG;�w�*e�WYz`8��ݲ�a͂ޛ�6}@�X�R��h���k@�ƈWU���h��xr��%.�8v3���z#n:d���rf�����@[�Je�p�Wh0*2w��kI�����>G�Yy��Q����=�(�
_^�.K����ֈ� IH���6	j��k�ߵ�h>��(�]�Y�v9[B̚�ҋ�!���I�D#�t�(<b
�����}���A�C%�Y �PL��Vez�^H���)���$7ue���{�b����"���P�]���m�uj������={���:����b�w0o�N�~F����ܜb�rH�w��j�ĖӸY�1�0�������(P�8��*K�zc�{{;d��d6��&)�b3h��>��I|����HL\������3�|����Q=�a鵱������f��1�_r*3��ud�����`���l=�ibU�o�
V�\`DP���:TNj`����~��\{����	��1���e�hZ,e����f��l�Z6@I��vpxV�Q��.Z��t{.�X�UZx{UFD��ae�0��%e��by��8AE�� e
z��3ӆW�U�aK.)Lo�>M��WE��b��V����@�[K�͍r� @�3��"�C_x��"�l&|7��c�z�'��9�J'ӋK�?usw�"��;�S�l <�7���*0��z׭-����^��}���9�@J��mt^ �H���ZQ6�L78N�e�l��88]�lGY��-OY%�^S`�:�� �0�W��3J�:|P��f�C�zNv5+���a��^0�ߪ��iN���@xV�K#Ϛ��%W��W?C~ϛU�!��R,��	��33�`�k���g�4F�Gc�*��/���#������E��R5��tXM��M�ݗ�@��"ZX1�>HՃ���T���e��p��>�fl:�L�F;��ʛ/w��j��� �7A��&Ľ�ޓFK���I�n�CU%[~?>�n�	�����GQ:��S�A��dS�h�	�<�"zƾ�����8n8����8�<.�ǘ�9�\���#��.5�����]��\�0�H>����d��9@�Gp)��2}9�{�$�}�%�>PIu5;����o^�5���ɳc)�M��O�3�[Xq�*��1���g��ສ[��6�X�����ۢ3�VQ�z�"��Q��g�ؔ��}�f�P�ݙ
7�XBF�K*������_�鿀RęK171�Ļ��kJ�+��f($B��+������Ⱦ�*Tg�� h1���y`S�[�dtte;,�j5��u�����TL�)�
�9lL�'���1������!�D�9��I�E���M^��o �����j

{4��Wɴ�F��w:��5
�PF´<j�h�/m��B���x�����]�4�M���|$J��A�1j&1F#��Z
^3�rw�$)�I���	�}�<�Dx17���,2~�� ��B�I�����a �d��iP�c{�Gs����[���I5x�OɅ��'��;���T��3ꈽP�9{g�xO;�]����Y�Q��280= �,���a9]M�b@�3��V��}�#�+��o)�Y&���l��=0�;]ϋJ�!XQ�ڠ����1����X�s�H�궁��^���³ؼ&^�k�:!����]��V߮��vH�w��~�M�%"�d�Ӡ�Q�u��5�j'�`7��^�+��SYT��:z������X��1��↡���	�j/�r�\���I����C�{����=o��=k5L�,b�2x��yS��FQv1ӱm�WV�B$�]1���]q����Y��B��>�����P�l�L�M��m�x�qct���C�^EIEXQ������5r��}a�R�*5Ŕ���A���ӥ� �)�47�NkO���H���Қ��곖֣i�����j��8�zKlZH���O�}�мw��	��W�ȅ��o�p�Y���u@���I��	�� [kh���#.�A�Z�C�)|Kv���E8ڸ�s�wG%�=���q��zV[�q��kL�'�F��-^��~|��<�����5)bGm̏D��\	̣���b� 
�&X߱�%��_Q��n۴�#v��8��G�I�qZ�bCLj�U�{���U�v��3��6mͬ���[�d\[r�J�!���>5�g�$��\��t� �ΐ[�	��븟�k-K�<��}�%��1�l��3h�1/�����b��X7:>eW:��C���_���W���`(?��񲣛�?�uQ4���|s@���P�� �B�%��@���V9�l���	� M�� �u�@��?��>�c�'j�$D��7����ǋ��h<	�bHv��7����&��-�%���p�<:�]�_E�O�<�=�aY������N�j��ց���(�
�wL���@a��[ʙ��-d��ZG�1Tm�	�8V~.�_�^D���lP�SL-*mg8g��x��<eS�HN
�f1��@�Y6����J灰��^zL���"OO�9l�������A)��-�շ3;�e]vf"�+����8��㺇f;�y3���J7
Eam��cY�g/�o��)��.�UK��'}�x7�U��h� e�������Nt=$�?�Tp��i��;���U��ʄO:��Q�q(�������auҔH`�S�0L�$ě�c�u�9A��VM�A7��^8N �$s����G=4����,�bu*-�L+�ݡ&�ꁉ��p�ؗK���PY��<��W~ޣ��L��Hz�~�W��;����t�nH����\��|�gE����=��l���FL��E8�@�teJg�e�E���Oyb��i�!���Q�$Bn�a����M/T2�xZm��R����t~��y��E�P:;��&��k���de]r���K%'V��i<3NSe��h�4���l�N�5.��y�e�H�4�2�Y�ɵ��4�Tx�,��6�H+�[��"y���N+8ͷlh��J�@��!�=��y`<��n��7����ҋ!�㴩R��1	I��KŬh�֚�>B��|s�E�- ��g��O8֠�?��E���t0U0$�c��a�Y��9�[���
��B ���i8�#�����t��.n���3����/����
ol���4Du�/ k? <z#�B+�b���M���9�+	p 
$V�v��(���0/��6S�F�_�~�7���"��U	l/�c�a�&l���z�UY����pmdA�>�z�\r�B&��e;���G�X�����r~��_%�(e��L�/�g�0r��~����eR�7�=��
6I�0���T�;��d��H�{���t}b]0���SԳ���xA���]�>���ׅ�,��ض���k�?U�`@p��Vް��������ݑ6����Z�e~��N�ċ�h����m���A�o�|�Ɖ�`�������e�t�o��I΢!q��3 2�#=�����4�T����OC��f}��� �)o�bO���`��DJ�N�Vf~5Da:Y>�#�j��Pd�!�&�ȴ1�R�
�o#�O#yp�8�B�`��m��X��əw�vq&M�pH�p���VkTNʰ���n��wȔX�$ޠڥ���l�ӅkLLNS!b�k���7�D>�Mf��Zi���(c?�Y1q��v8���x������-mRN����il���)z�20M�'D��iż���8����y�=���m�0� ��||�i�Cu�=��]M�ƈ�{�
��훜	��u~�g��jݟ{.����+K��w�|IS�_ˈ���o����M�� -���8�Z��Z�$-�o!5�녺���$˝kB�j)\S?FU^]b)e��=���K���-�Nk{�թ�|�oid*����5�L/\_�.Nx�l�e|"7�E�Zt���m:4�Ԃ�h�^�h��!-�t���P���(p4��3S�a�-�;1�3r,�Q�W����` �jfUC�]�dnm��ܣ}2�&�-f���D	�|��+�d�R�
���y����g
���Kf�n��V7,2d��&ߦ[���J��z�*8��=�K�:5�V���b�����֤~�9�� ���+��w���w��x���������O���tx��+�IaH�����_�9��N�H��M���拶�s&Ϭ�H�!�ۺlAz���A;���Me*�1NP�3FB���z�i�=Oɰ���r�79'����dy~)mf�+��<v��K׬��I�ɩ@�/�L-�	��dr�~dhw�� $���ک	�I�FO�jπ�i�~�ጇخ��y��BO�n�p�g��ܮ|�K��[(��q1{9��Lk#�H7�1C�{�"
��F*�n���[ϔAS79���?��Ī���BSc�XHʉa/pI�=�H���i����WU(nA���	�Vp�o��՛�f��Ѐ�6���~W����,�{�h+��,u1Z�f1����|�� �˸	�=`��R��X�4�C��E���|	|���,�yJSLa��'En�j�Wx���l��;�G6�
̶�N��KNӮa~� [H����~V�.C9�efG=��4��g��04�6��=���f`�0����e]�;��H���E�I[解��P� I:t#�ި�^�Y�I�u�¥	�$Pt�ƍ$��\��]��R�CB�zK�}�'�ω�*#���)�D�Hx,}���%�JO��$!`�sO?Er�]̹��pY�m�yW���q���Ϊ���3�R�&�z�XK��_B��Q�w,n^x~�	Q���W5F:+_`�E�6dY�i`�b�RTp��Tɓ�Ҁhwc~����~�S�v�5�W�Ql�ތ%J�ǹI搪���&m�����0ϊD"���k�����6>����7y�2+����5��U! �w��s f9�ǎ�_�H��;�߭b!��q����b!ܡ���0��a�˨K�P9����3Ǔ�aS��iC�꧗�Gcp|��L�����qx�h�!s��	�\��yX��z	��Ǌ)�&/�m�
b�+���\4ӴR,u_+��hnG����~��k��|5zRK�=Z��4��i���`���e�����{
��e�"�t2k3'�h�Ko��� �C���Kg�j����	C���耩fgp���_�qץ��	�E������4�����E���:3��%on g�Bt�X�UO�9GZ�dyްh�ݞ7b��F�D���7t_��9���e�t����b�ʎ���RL�Ɵ�1�����"��&Z�r��'o�V���M����e��<�瑱��] �Z�H�
x�n��`M�4�[�YF,�e�op��2e��3��^%0F�;�"�I��>�I�;�����^]��d�{�G/&X�R���Q.�FUAZ�ĉ'Y������;)���EIV9����XE� Q���>F
���F��Э�}ɀ vo=�o��$�@� H�)��v�Y��IX�W��b�	Wtƪ����.[T$~�f����*& ���	�s�a ��
��es��gahu<�T%z��Ȫ��S�6o�߉毁�'�ü���:�Q�5t�@�	�倐*�!4.��y����K~i�w�8yAv`R4���7����N&X��uZ�Hh��^1��O�/�f�*P,+�i�}�Ǒ$ 	��O[��OQ�n�ԍ&܈t��!i;�Ol%_r����ߊ�B�K��t����I�p$!=�u2pY��î�AV°ً��S[���0\/=L�e�MW�P�ޚn�%�����u���>Rɓ�c��H�)*3��qGM�ܥ�D��z���JFN��k�dA<����֠===a׊;�����Vյ,��r��*�O��}�m�����������;��!�VR���<�3���3y�Zf��J��]W�	r��o�_�4Z�=A�@Ʈ�Kg���#.�h�#�I*�
@�4%�.��@2|���@�}e8��k����7?NJ��nY6���4��8��2���\p�)�NQӉ'?'f�U�N�V^�a?�tus�Y܉�1b�9��~x��,� �����v`M��+�sFm�m;�����+�rb�o|�Z�,�-b�{��]÷#r��?�!�4���\�mр��Ӓ�%dȜ�wU�E6kzԁ&�]_OR�������AD��U2AQ��_�-h|����V�_ZԎgejb��������kR'��S�£��KF��s4�{�<��Z����z<�8i�9q�����X����*�\�+���N*�ԛ2e���"©k)���3�x:�t��ob�.	sH3F�	��x�m_e�9V��BG���>{־�s��x]F�");�2�i���V�.����ӻߔ��sG���g�Ny��Gd�G�2�e�yJc�(�c^����`��bJ���β㜀5zL�`T��/ܭ�d�0/���~�0"��1!�p�Aew?NeG����&N��|��E��i�s�}w��y�C1��#F,Ӫ�{;����L�:�u��v����k�}�ؽ����J��ڱb^e����;2�JClC���be���x����O���QA�����K F��R7n�\5�*!��,B�9D(�R)�լ���G��bɖU��_�(g���� �WI�1��6�O��N�l<jc����hA1��Y
�Ur�?aWJ��r��l�U<��
S��
��W���)o�U��>��n�l\�Q^V	>�����Q�@Yq��]��t��))`���@N�x��e2��60�pɾ��HJ��O��R�4�T�[��3�q��\��8��������2Jwm;]U�K�xg	��aFb��~M#K��a�!�ZY�A%������ �������%	RɰP�J�*���d(�:CD��í��czE0���[aG���O�"_YX�;���ͫ�W*�F�ZswZ�y�Fs�w��=�����כ�A��!�b��v� F,�LN`���h
��,ͮ1Yol` ;����]�*%�#iڴ���AO�	�A{KQ��?i�ǚ����*QvB�T+I�U��_P�åmH�V����k�,قB	�!x��-,�tj�AD:�մ�� ����o����X�À_�߲x5�ɽ
�l���\����9�@�K݊��#F��u��QT��Ѐ��=�?��h9���@_�z�g�;��{d�8&]o�'a�#�E��V�
����`��tbǂW �"G:��0�9\��������uTa]Pv�s>�,ذ��	�w��\��������,�v����b8���8@1}{�$��꤈{\��:Cǥ�����Q�,�.��%����Y�c!䋪>pq5&��/�h/�9*ʫJ.Z�󛡨���P\��O�Ds-����ڜ��+b&��Gl�����B�o�G���_Jk�=m�t-ۥ�%]�i{G"ū;��(�[I1_�pPL_����>�xE�rsD��rgN��1ϰ�o�8n!fGb�^C�BG_Me�G�齧l��w^�/��\ލp!�Lu-�|�l��o�O���{g,A,5+��" �ʤ����П��V_�TΥ�>5ߡ�w=��!��f�����"=\��#�>�Ҍ}5ڇJ^�Ȣ>U=��P��,����W�3���*쵯��7)"����
|6���Z�4VpWj޿�COUrX�`/Jǘ
�ңXd{���!<��3Y2� 6��vs>���&�b�����No�i��Di�o� f)U|Uܲ4$Ї��]w�EՈ���1|C={�&��}o���$GC�pW���܂�|�|V�6��^��{M8�ɩ���պ�U/>��� [{����g�G��|�x�K%��bE��Z�ϙ���{uh=�DdA�Dx�qp�<\D�<�?�"�̊�t/�1$��P�f��9d���xf8,����&,�(��C;g_�B�StZ81��(�|�v3t��B������h�7B!�aD/�0T��X�ù W�nv�R��^�Ȍ�!>�N멭����vs'����Y��O�Z��L����i��bLxx5��0O+��=�$[�yQ�:g뉖q#Ʀ��/����ɽ*���#G`텯%�3L]���ܕ��q�C�~\�\	�e�䃟�]�Usԣ��=�����*�<)�24rZ��`D�!��u�ؾ8����l�X�i�X�35���cz%
oa�`�wZ��g��c&ʈ$̽����9����a�t@mO�?���>Y��5-ȿ�Fqf}�J�I�?�����_R^ �4��-K<(ޅ����BOQ��D!8[�� �d�kB�b���U�@Ǎ$�cçL׭��C��bE�ԬL�kZ�cP������P����q#�qɇ��H��B~˫V�%�7���3�E;w؊r�34[#�T���S���HӨ���F5�b���T�41��/��)�`�lH��'��l,[���˝�	N�'i"�.+-e�M�����w���keΓ���K���o�I������+#�#��xEew/�y���3U �G�� �n\	�%�9�0�'S���9|t�11�/���h�`[�ݜk��
��b4��\5�H���z�%�A��� �q�~,�-*GO;�eo^Q�Zw)Im5gl�SY��7:�܃��^P��,=�w��^{�{�e�~�3k'G��s�,5��I�BgXt��~�t}H��l��8ȍ�l]�S8Ů�����?_��[�(���[�D��UO �O�a�����?����9��i���x�uQ�<�T�Fc�(yf�b��;�	�#�T�(�e�w��D[B���S�������	颖�%�YNQ{���&�����1�i�!ӫdi,��0�cl�4��ﳽmU�`֚��`ݥ�E�wA�ϐ�k~<7 �ɛm���3��k�,�q_�.E�l�pN�!zc좰�@���R�����&�-4C���߇_R3��`�!̫������W��j\e����8 ��Y;톢�B``���p悮Rzg $�p�6�2��2ϱ��W����I��ex�o�YL\�����r�v���>�|����*��	���X<�;�~���-��<��s;���H�?�z_�u���.�E��0�?�=��#U�X���1�T~�o��	;�����C�ak;O���b�5���l�}�qT�@Ku�����8:��������!�ࢂg�]k�|ĭ�����r{J:o5u�w���
���q[��|��~��5�Ol��c�%\�q�a�O�N�J�]�;��Q:�����v	��Y�(����ٵ�@����v�z 
e�� ߵ��@�e��O��d.@ۜ���>j�|	rC	,W*`��F���T�xR�貂���O�#����U=�p��g��I.����jA��>حZ���[���ȫ\���ң�j��Ha衃jǡRF����9���x�l��3<.s��cw�q� ��KC���I�!cw<u�:�*���͛<�2o����P��&F�&�p����ՈSjG[G��������>K�Z����w[m䠟mn�5l���h�P�ȭZ�XC,��;�Yj����{�j�~`��Δ&[k7)���Oܔ�u�!��#&f80c5��T�'�2���fpf�����A�]����=�Ln�%_�j3��z��9��~r|:Zib0vB�n(���ǧU�MT2�&=t�V�K�ӕ6�w�i�.���[�[� |Y���C�����ܴK����E�g�/.�@ʕ";܆����-6�*9�\�ͤ��T����t���K8��5
kʤb�c@�~�sP����>o�[6et�1ܗ�s���3q-*�|3�]�Y�@d0H��Z�I��Y[@{�}�%��\5?S��l�)��.���>[��pE؄�5v[�к3��Ln�_��%q$��j��˸��ۉ%s��j��.V�}[mڱ-�, �B.�g�r*� �U���u$h�O�	�I��"�(~�w����Ҿ>,�En���X�DY�&�wہ�HRa'��ч�e�}u�U�1��r�-0���M&�j2i+�| u}:��3q�a�\�Ē3��/]}%4��T����Qcq��d�'��Ѷ��]E@}�4r����`:�D�k�R�p�ґ��ŕ?��"f�f�Α��[>��Fj��;*�A�;˥��2_��kU%r��#� ��'���	�����ncK)Tx�4�)��0�)�s�d�96��X0o����I�)S~M��x@Ǒ�U�	e�z���s2���;�p��jۂܿy�U7~Ș@��;�~�tՂ��E���{��h��z�3A�f�����rW�C��`�#���K�_ېԡ^e ̓�z��j��^�ko�|���N)i�-wp
���g��c�[2��9��EOS��]�)��b{ �pZc\ �8?�m���m6T�f�U������|��*ݡ��
V���ݛ�zX�����F,�28É:2Y���s򊸧�j���W����t��T���d����,�p��bi�����+ 9+�����FA��&?D�k/��h��0��}�*>�,�7?���r(�>r: �Y1����E�ժ���ɽl���{��x̿�7�K��b�s�k؎��:Ǖ
�}�2A�J7���K�ER=�`B�hh�mc;B"\,M/��yXk��g�ڼ&���z�jV�!�um�|y<�����UJ��*�S&�3��U���=�!_��$�j�4�@�	(Z$�y�<>���E��fi�`2d��
�<n��VSf���e�Ρ�hN��`+�2���O�h2���Qq~�#�B䐑� �D5θc���WB��gkNЕ�fg�O�fO9ߤ�g������1�IG<�D}���k8�4�TQI��7)�T��^�v�5��CWx�,w|w�q�u��#R�N�>'��؛��V���(Q|�Y�0�SæZF��%�JH��	<yT̻��u�B�7sf�5��En;���:l���t��"�<X����r�'q�~����J3��U��A��Ol��ܘA��Ȑ�e�z�)[��rj��i���'g-+{O�jft�Pą�09�D(�?\nr�;���ɮ�h*�� E�&��Y �[
��}��]�L3]�1�{�o#��?�#'d��"9�����I�g�_�t�Kif;,�)`���$,yN�rmsWI�뾪��D鈗#��]��*���8�/QaB1
��(J�19y)�^����s�n��(���i/��9����D�@����$��.���$��}�H:��7�m�',N���K�c�#|�~`� ��SC$!֎$��{x>v�G R��U�B���Uw�k���#w(��:�Z�sʉ�0�C������]a�̜�;����Hc��0��n��Ʈ��F�<1��S�n��~�Fwg1�<�'��¸�P�k?��yq .3hP�=<�
J��d�3��zi�.�.�c,�;�|�H��3�!���q0�����jΑ
�����0�|��_KLK��"aN`������[���DY՞jL�4� s�@{.KI�u��!XY� !fF�,�"��#:^���D�z*�Z���9�k����5�gFޭ ��灢v����G��QD�h�~�}�m���P���B����e�)~�?��!��՛6A�ɟtX�S������t��E<�h�]ò8��Y�=�b/y�m�M��q��g�%�+�T�G������AH]���)K�b#��S{�S��+�����5bݕi��+�"�+{���N�X��#��)�Iv�/�k!��q`@\`/l�tt
c&�-����џ&+�L0%���p���ܠO�hϼP=,��{ӻB�'cd�,�M���C���Д#0l�*rz|�ߨ�V����R��A� 1N����h�F{���)V�?��Ǝ�P2ˤ��!�-���E�,s>���E4�Td? �	���>�¿�8}���<T�Qj���i)�'�g�kS'�b�}R�SLEĖ���6:یXɾ����`�2�Uu�Z=��a�a@WG���Vfte�ՠށ<����A��;w��kcV��4==�C��O=l��1�ph@�ֆQ���%\�u.�<�p�чyWȸc�:���m�y7�5q�8e�~P��{�^;�k���Tz��%n�%�p
f2Z���`6�;�WG��7�6��Z��ٕR�P�ԧh�����B�J�������F��Gr0�Β�cޫ.�*Q�t������T�gy�ڔ��kä��Ɍ�Z]������=b+�.y��k�;�'޹I��G�G@�c�yh����fb�SZ$��������v����e���Wmp��jk)�������T�d ��(s��r�A��k���Y���(3A��5�s�)=<���} 1.�W�V���gc���.�������A��Vong~?A�F��~���Ok���A�35Z�u��ڊ;���׺��+���C�2�Z�,�b@�o�I��?�	KQ\N{��R|9�����fw�J� ^G��ډtެ��#�۽k�KqK�.5�S���	a�ڜR9�3i��f�H�� 	����W~�Z�M��T� ��̽=͗��[ɵsCiO)Du��a��)���DcF����>�M7�Eu����6�O�j�T����:�y��tU�9��rJHvRrZ�L����A}c�Y��ඃ ����W[�)��b�-��
��r��N�z����gv��F��B�c0Lj�Ne�Ur�E�,���%�աȌ��U��Ҏ4����=��]�5u�x&�W�������{gmW�Ey]B5Gfu�6rV.����z4kjHӥ����|�3�P;��/N�)6��'�-:V�����[�o1��#��u����ж����/�c�LD���x���/���%����JX�񏴓�j'k�
�!`bi�Kf���e�[�V��eu�C�Z��׻F9Г �B�`:��(��т�ǥ3�{�?v�S��F�jz�!d=�G�u�)��OT=��SJ��w�U&|�ԣ�~�6�n&ѻ�90�������H�
*��v��0�h���f�P���� F�7�Ó�����F��.Run�{��2(�Ni����P�.��;�˅�=	�j,	Bj ����am?91��h���r0��`�>m>�,$�����7ݞ�.�����ͧ�MU�> ¡��q���ƶ�<k�V�x��^�l�Cx<KW=������N���A�/�*�RZ~�����0���rc�^oM����i�12?���SzאJܴn�9#�#���``O���g>R L��1�/.�}e�N?��tp�|ʈ�۫�>ZF̭�

Zx�P��9�����M.�,�ã�?C<��/9 	B��E�/5�[oD�jBv׭Fpr�B:J���NE�R4��ʏ�f�24r�v�v<0�껰a	�������7��6.���,�)^�H�q.��X��;J"Z܄���b�Ըt$�sL>����L@�om�t'+�n�Nr��0� i!Qz�����f���t	A�6���τ"®��&�kЛ��W�k^�����Ml��)�ǂsP"�Q�NȫƛПц�,���ww%ݻF�b�����\���2!�>�{p��?���T��0��cbS���hUOH]y[�Yq��2�x�#�h�>5�����Z��K�]l�(|6~�@U[���2�uʂ��� �B(��q�	ט���[��z�{�W�o}�v���X5~�71��X1Z$kW�ݔD��bM���<������'��)�].˥vc{$F_�I�?���bA%w;~�����as �A�Gk荸|���
[(qTP�ur
�7=�}���P0>��U��fQ�7���I��M<�I����rZ���*�.M�<�<���IO�4�k�&���6t@��0�fhT7�#i/�7�o���}-Q��c/�$����G�ɢ�ɤ�Q�o݇/a45E�Nd��2:S��GRo)�PM9G�?�4U��n"������: �wd����A���7�����4�MM���)2�u�5�u�UC��B)��O�9�"�*�g�4���֙>^�gw;��L�v�ٔ�9��>p������੖x^��������͏Z�ݗ}l%3�̢�/of�B�}|H(+��1+���(���q�]�����T���Ɓ�/��Ģuȿ�3��2�5N3�:�D��k�uq��*�^����Г2���hÛ&���i���p���Rp��=_3m BP��%������z����-=�v�r�G��qs*�6���(y���d�����̖I���	�5��UU9bHD�h�N�-N�\�y�DM��'zؽ�+��|�S8	}��8���N*)�G�	�a�E��$���e���c�wx2�A���n�JT���H�[a��)��u��	��.���˶��C<w���9J��Z�<(�чfV�����G��Z�Q!2�})�0#��Ʀ�V�|g���*�p�~@�L����H���;�ƐA�$�aˆt�QsN��]�~�J�^�.�`O�7�L�Q��h���.�W�n��_l W�B�?�A��멋mJ�{���PV��/?Bߛ�%(�D� -�
�@笥���ג��q���@�k;X�C�g7m����^4����*�V~�8xw�v=�S�##�J������u9U0�J,4�S�*����O�|MȬ��1iu	T��i��� ��Je? �#5�ܻ����U4�������<{�}��:��u�*��(c�_ui0�F�K�8�c�?:NI~��6�S���Gu�ṒE���_xǗ~��q�5��h����ƥ������wqi��	i	ri�
)v��T9"_�]8^��E�����K�� sd���R�5��G����0�2tl�}�N�Zd%��n�O�,rU�����^L�����qJ���+t�#���b���F�)/��
;��. ��"�6k/\��G��T߆�-J�F_�����tSD�c����s4�zs�`���u&�_��F&�ȇ�0����LrǑ.:����	>_\ɑ��b��xS�!�>�L�y�Z�a F��9��3VwD���(y{8Ke����vW�nx���>7+���O�Z���G�	�\�}�:��˧$m�{׸��o��S�	��+�E���.ޯ�����U#��B��_*�Zꀟ���2/�7���P^/�&���.B��a��@�'�����hA�J�כ��P�$�&���VHi���ێZG���	�Z^=��-Ý��&8�c�8����L�,�=/���(�U ���a�|���ѥ�����5�r�E�B��ɠ�xw�έ�޼�ŕ%�7���$M����t���~����_�퀬Q`�	��2�ͼk&��l(,��-r7�LEB7�I�`Ր���3Ҿ�]KO$I�3���O8��IωȫEP�--Ww�KB�A����u�c�$��O��a����4��� ��C���������}�h���l��g��d4��,-!�j�\xĮ{�̼)��x|y���%���ݙ�p�]k�Mk>T��Nc����!`Y�sgA�.i�����k(�*��T�]�g�Nu�*��!�D�͡b���L�B35.IR�t��M�S�IYz՜���i�,�31@�:J�����t��j���	�Sh��E���
/����^0@��o�W�?�u���9��t�d���aeZP��� +����N4�$��R���3�+���B�9,z���@^��xJ?:�S
�6BW�Pn� #�]z�|�U�|�ղf ;�;��f�Y�S��r�L9�!,.�`3]T���`�K�\��o����;dC$��^âE�l�f��1���S�B�E�~pq���_t�����9;=�St���"q�J����������!�\_��z�'���d����hE�'��,ˣ�ѥ��kz��gd	��çp�= �.,���0��|�7��*4qn�D�C�dрj1Qt!g�$�'\e���d;�1�u��p[�����J�=�Y-����c#�0�NX��%1��S���������Û���V^H�fL�P�z�M~�Ķ4遴	����h(օ6cr�����\Ϣ:Y�n�q��8Aʮ���j�����
��^�@~��^�����ip*�}��53'E<�P�Wm
�S�.ц"B��L��Tf����E��c��Љ�@q=�/��=�W��f��.3�
r�C#z��~�w_:L����^���z&G��N��`PJ^� �zw�m�,<�,���f�5�uY���3¸��%>�!g`��5f�2"A>S����{��+�ʣ����S6(�'�h޻��|c���mY��������rL'4���J�Q&���~<�q��oܘ�h���%���6�{]o	.]@>��3^�\���J� o�;#;�+�oLVT������!�����N�G�YEj�{���٬��޿M��4�l^k�S�`{�+�2�����Q%���Ol$-)\�#:�.�� Fh�b���?�M�\f��jš�>�&H�Ʀ��>���De<�[�@{�:�D��	= ̗c�:uv
�T�E�_�&h`�U��=�)���p�[���}+��m	��MD��"��AZa��̰���Z�|U-9�u���<_+��<�Ǫ��>��� �4n�߮[7	� C�r��qs¿��m�EQ�h�T�����O|Hk�^(c�Ĥ<���(�Tvb�@y��sM+�c�T�yq���7��oMdm&h�,f���KF���w�E���?�����s[�(6�r�2ϴ+�,9��S41ONДF8AA��AF,ƣ���	9������@�q�C����*��c��N����`w���$�t�Z�$ڱ-V`:�--�&�q��L��G<?BMż��f�p��.� �ZЙ�ݐj�΋��F�1ʍ�Al�?g~��`��k�{�چ#3�����,�G+�Q�(`ZdHYE�ahW)6R����~y����UfH�NA]�*r�h_�4I�,�w+�]�"0~�_vް>�ێ�:ej~�_���Y<Z�I���@:����0���Ъ�֤^��kD�`O��8e����\Q��N��ꑚ$�>��Fu0͒�3/�,���X;O_6	U��M�۲��}*�_=�H:	C����bc�.̼D�8�@�if���	Y�l�Y���wym�N����gP��h������]y���9'�Ўo��-F�ＵH��;c��'',�Q��;���s>�����U�\�v|����R?e&:�F����L/dE�K=+m�z!�j��MJ�8��N�� �����z�:�}�˸ZQ�Y	R�'��J�n�HIq�B����W('�kCR�@?�`6@��׸�gZ�l�K��V��TCrX��M��漳����"�<�2@y�gdX#�0���x�p�.F���G�>��=�S��m��cg�a�LVKє�ߧ�����4z��9& z|r%���^�7��*�����Z|ZiţD���8�C��,󸟀Q	�;Q�U�)<*u�~f��YYK	�F���d�����#ZB�#��R�񲕛�&��B�hY�Z���N���b�H�c�i�E	"��9�t|�Þ��{��24Px�o�c�*�eב��ޔ�~���7���7���e��0Ǜ��4�X{ ��^���/��砖-���IK����]��Qs�׽����~�7ڽF}N'�μ�JM7J�5���ד(�\��f�������BV��'j�h�Q���tմ$��y&~R���x�I�E���u�9�W#�T^1
>�0u9! 5(8aP$]�YN���qC�mى�����a��&1k�ݞ]��H^8ⴃ���0}k=@U?���%�OnYlg��!/je���N�DI��T��]�ٲvٰ&�$y���EN��#��^L>U^z���I���{�?��;50�l�k#�����s9�kU�$�>(aGmD/�7�x������f*�?u4_^�J��]b+�]g�/��t�Ғ23TՈ�����ۧ'�B�p	0�H巫%-�te�ڄ]�v���Pq�"��G��c�Pү��s���I6��� ���W�;���S�},a�Ύ�mP���>)�`.^�}[s�+"���(�lZ�uʠ͚����~�P����? D>�L%�س�
f��(YJ%��#}�C�u{�����-���z l$�?S�.�~�!gwX񚅦
��$
T�����"��{���a��|���Oyt X���,ӲWL�`��
�#�t8q8��nГl?P��)Ε���0��<��<,&�^y�1��|r���x��P���{ND�}�y��D3�vP��e�vW;86K�7��"�,wUsL��I�=��[)�ۢ��@�xP�������I:��<x�К%_�!�)��&{��8=�%;R�5�y��1	�����Y�{����TY���Õ3:%^dE>N��߈~p6����sݤ'��``+w	U���쟑/�	a����������ԸA*��w�0�oޘo���}�I��zQ�9Q	i�-:-����@!��x��$�S�H���� ��:�K���?��a�w�ë�� �l���w���e�+��9�$E]?����6�����u˂u�t��u3�1��|�^�����^�v:7-(d���tƖ2�c rCȫ�2y _��
'�e��l�����'2!��_��(Icd@��b��<���Q���o�(�w(���4`"m%��s=�m�c(��{~�z7���Q�z��̛	��H�2 4?;���u�ldGoo��Rڱ�B��a�Y��\�o�Y7�B�H�ٲyh[�9PK��;$�+4c��r��Y��#5�RZI�bB /ϣ����g��"�ߢ�F}#�����c��`��h�YE��T��$x_k+v�Nk��x+�&�6���K`L3�]��h�s�A��������KZb�R4�x���M�����f��Rt�_bϘ3�H�!X��\�"�I0[ջM	xU-��h��k�ey�$�k�Nh)ڴ�o���cm���\G&��Lۛn<�h�����ۖQu��	�;��|4d*�ud3�~�;=Sl*~F��ź����S��s}�����1��� �t�SG�q�wx4$��da��6�>���D���۫��"�	�c�>
��̛v��v�@��{�g^bMԫA3g;�3�!s
3�ͧ"�Y�Tx��S���Tb̺�r��t�pg��R���/϶��k��6�>i�Y��]�FwL^ ��d�/��	�!ʀ#ʇ��?���a�y7��LQ/U24�7ɇ�uK�"J'K��e�Rc�{�}���j�$S921n��F����(�'����� 8�F�̥7�(� �>_�(��8>�3v�DMU���Q��;t�4i2�?,������в/�E^��֚+u�8�_�{�&��(}�w	�&�޽��ĂY<����H�'7����_H�^��)��i��Z4Ƶ0A��� A���	'~�a��\�EZ��ͭ
���ȿ�p<��!��(R�i�ϭp*�ڛ�>-wEҾ���:C��`L�ۥ���{��h�긂F��q�\nE4�޲�_�&A��</��%1�69@P�z����K����݌X��_��c�`z�\��*����}L��"a��t��a����X-����U�S��|[�����/K�u���N��.(+� ���2�B�q �QU�� �Ȉ��Pr�0�v�g��ۙcf�V]�m������),U����?{OsE���qX�� ����kE/��P�u�\]P �E����,u6����E�G-���w��5v�j�4�Y=O��to�
�|ǡ�Ζ�u/+8*+Sd��x��6:��\9mo�ݚE��RD6�AWer��=A���G}��d�Ut��./ZMg�@N�19��U#G�̅o�;o����[�%nq��sBi=���a?�vc��wi�L]�%��<VrX�?l�}6�/���r4T
���|�?�a����W/��4�������'�i��^�y
�cq����B�Ii/Q.��q*]��W��/�3wj�O��͸�֏����%��-�v��_�<6�Ay��e�̞�,Jz2X����O[�D��ź�ɼ�Ͻ���p���S=��o��'>����V��
?̰
y$����:Z�Q�Op�@�i5EI鑏�
�ҏV؂��-��~qJ�h�Ԭ���R&~�T:���|��Ui��CP�E��b}{F����T�\�!J˫5x"��_�0<y����`�����;V|l:�͚��*�ǉD��<�Z5��-4<Z�
�`зB���CnDQ@�}��`��z� �8��9�<X�>�5��.x���9w�m��7�w�1iQ�i�k��D��\��=$}�0{�����ñ���җ��Ljԏ�b�؇����.�ԉ��m���:��Ȳ��Z�h�L�$�2Zp��L��k�K���
�%6�=�e�oz���w�jC��ץޅ�VEe���+	̅-wKgK���Nd���S��)n�µ��y��n����zx�9��?�=ݾKz	��=��sڑ�۱VgT˂z����"��wq%։��b�H�[R?1W�A�A��TF���.eրA9�.�����;�Z�F�5w��n��7�����ɔ�HW�'�%l6$0�DܥG�>�8���Ki�����)�����Hqb���h � 7U�����H��ۥJ��5�n�����P��"��yK7b��:-(��YS�b����4Ɇ��a��g`P3�9��:��սz���c���7�2Y�jr'h5ȥ��R���*�O�glGXG��p�Rw��7[%Q���!���DQ�g�8�z.��!������9����VH\���b�f<�L 8%�ziy@��R�;o�RS������ � ��cE�똾Ƹf�~���I���n{9�nN>����4�K���/� ZD�a.���g:�ζͭ����k8`#����E�z�9A��x�z^mXb>F�9B��E�����'Ž��E��j2������s�P�PV#��c��|�C��R����t�"�c`�
7�>(r���닄^�O.��xf��4k�Y�V��^?/�0�ݕ��._E��Y��!��l�;�~�V(�NW6�BM�y.���u�������:>;�h*"TS�E;9��Z�ʘ���nS�'�5�ѭ�P�u�5�˷�؁�M%;NƔ+�l�k�8��r�8	�(ef���kecB ��m1�%O�F��s�CI��^܅�O�<��	��L=Ų�s�#q���)�e�D*�)��;L��T�n��M�~>D(xÐG���E]���.&�{N
��p��w�����s�L��N���f� �� �+ #��X�U�����?5��Ks�Ҡ�xH=�N���7G�7>
�s�q	z�%�z��J)�����p��p[c�ە�r$�;,Fjč`��ʈ�}�2Kj��z���z|"��Xn)��J�ظ�Bנ�'9�>ݖɺ����L����Y7"K&�F+G5q�%>YB�_���YJ��DB&l��w�/ǢGȚ�CiC�E�>a���?6#��� �b_d��9Y�F�2�,�a�����%�f���i�KSJSRn���F���	ˇ+�����9HI��M����!.-�-���Vj�me�e+�@{��S��p6Ÿ�9���K޹�Og��''���Wr���N��*:[^?^�XT~ :����������Q����5�5[����#5$ݫ�m�	�����i�#9.A�\?�6$�����v��/�u ��wy�5�LC�zт�7��]�׎�K�a��+�������%��	w՚u���P~��b�ѷ3."��? �"C��?�u�#V�%L9$�ZP��y�w�)���.��|,牋(4A	�g���B�Uy�a���zxB��ב�q��P�F}h�M2)âݣ���!��lYI
B�_1��`�qD�����r�H{Rs�I�-�g'a�\q{� �TNڶ�&a�5�>�==F�a�o��PB/:@ت��$��0r眬0iKIotϋYP���!���\jC]�!�1�b�p���_$q�Z�9lp_ܴGğwȊPi���T�T�:-*�g&�m|��6co루���o!�P	��o������R�Z��JTЃ�Ke��z\��CU^���Ct�jvR����w}n�b�_&���z�
��Cp����1d�cc�!T�����4e|��=�L89۵�85�l��w%�s��f_u �|L�k�S�6(�O[f?M���}u��όܼ
����wS����uta6�5�Dr����}�Jk؎�b��'uf�A�j(�k}��a�9FR�߮�Ȭ��ED��
m�h���@�]f���&�8�A�@P�(SMi�?�q��c_��l����]���� ���� ��V1�N$��	��̞[��^=��I^�sn+Ê�[ն��v��4��Π���2=�j�[�����}*�Ho
C �i�����)$F4�WHsD.(�j�8Di=�,v1��M+�m���'�$ޖx=.px��)����'<���F��!��:�֏��:��z�� ���`R+u���!�;�W���S�U�Q8����S9��:H�y�de�kD/����uj�>���K�_�Jj�=p�D�%����B�!�ʘ�a_h�A"�n����Dm)����NݢY��\����P�Ь�;٤=�-^�޻Nˆ�%{���^�].�6��tр��cn�����NT�}?��:�qj�#Ѐ�a��G���&D�4��[h	���탃
��[dxҳwq�d� 9�4]l5c�p������ퟓ��UI��ʝ���o��p���<k�M��2Fb<�9�#%愖?�O�,Fd ���Z��˔�6ܽm��uƱXxi�^��,̄��K�����'�x���Bɦ_����4��YwhM&� 2嚷��
d��bN��x�۪������;���1��
!�Ǔ;N�x�d���K���J���%�KU�J�6�um�{��xV���*��	)��b7�q�A�ݓ��#�}�����s�R������p��<B8ʦr�b��	^��3� �9�Qt�G�i]m$yh�&-he�V4��>�,NGsgq�������w~����o��/}��� ��y[#^�J�Ί܉�PV�٪z��9��/�fSj�mD�o�q3(L�BV��&�����6�f�/�2!1 ����c#1_G� +/�{��3�Fc��J�ݝm�)k����S�ARZ=4���g��`�J콴:�����w��!�ᣫd����fa�%�wxhi�G����yxv`�B�9+PD�O!ZY���pgn8C5��	xE�Ԩeͫ~����Q�B��f�m��>4��ad;c��׭1ݩ��0����â%��0o<`�	GA:���?�zS�*����kyN�h���_��VT���W�]�g��K<2�~�ݱ�*�?�I	�^B׉����>L��j��'a��]�{t}�0�����v�uL�`��,PU�̶+8g�d�`E�ܿW��nv�����(�������3A��+YD����9$%�Vd�.�i=fD�i��I�����	�c��~ ��S_Oz��l��¨�����ƾ��F��S����ߕE\����oz��N�7T��	���į�d�P&B9��bO��Ӱނ���/y�]5;���m�4�ښ�w�|r�y��)}��,Y��y�*�}No-�y '?<�X��$��pib�\m(tT!���K����(�S�Rrߺ�@�.X�s-�E����P	�-9���.F�c��+��u�,}�{�c"�*M�pƟRx��30�WbI9�	��t�Y	��V��P
�7�:�>�RD�"�M�����7���xr~�6a�� ���@*|A�D�lgn�^����+�DC�\�T��"��3c�>�J���;�%�[��w�h��R��h����PS�$K�gC}"�|{L��'hA���Z�����$H�d&�2۱�n#(;I�T���Νi2ꛏ�7�h�� � ��� �4i`�7�@+x,��(ZԻ��=�N���~92��K'ը��BF� �PN��TEd}R��X�ΰ�ϡ�$�k�zu��0�Fw�eN�*�E��Fj��E�'����2��� j=��7���6�` 7�e5=��������R�'��"��1��3�Q�m��
O;��;ba���]z�j�L�u���W������{�.뒼�â�t��K���Ҩ.�P濄���Y�C��8Gؤ>8ś��y��u��j&��Z@aO����p�	����L3�٢A�S^5)s�t�[fr���?��`fH5d��ڱ3��h���=E%h��fmL��\-�I2)^��7��_�rø�m�C��ʪ�TK�&���#|�vڇ���`fwL�[d��#���I�?7&�A-��p�h�������S�Y���lxh�bM�!�Q��#���_T�EO��&���Ʉ⨹A7R��K�<�fx��f���+�T|˱|�ܡc�P�mN؈��;~(�.��1����i+0V֘U��O`S�14� e��s�Xl�O�u���0�U5��`-Ԯ?b_Y����y�<����ߚ˱��tAx�0x?55��ͮ���&e�L<}�KZ���SއC1���.�hY���e�Z�@e[��R��z������IAO�e�rWn�-T>hyU-�0~���
[e�����RF����3��	\��)T��K�L� �_���@��g�]ɕ��1����g0�s�����-u�X0���e����O�;\ݜE$�A��&����>����Τ���}�0&�׉��e����lp�5��B����L�'3(��
N;�*sqDݽUE'W����4��W��s���p?��/&G�V8��n�m�e��A��Br�Þ�B��:��5��@��p����
���j��f^d4���\j��Q�	�Iϟ�@B��4�i�cO�Z0���F��01���D0�w���NA��4���:�(|� ����2b�=��tVը�BbX�Ok� �$�ÕA�8Сxki�أ��Y��aƪ��ͺ+w�W�ő]+_�2#P] ���R�y:��(���;�mI���/���~T��)�ȶ�#�v�>�xj'2`h��ƑE��m � =�q@_4�t8�F�i��	���MeU���X7&RՇ��H�y�<Z	u�,��k#�/<�%�{�pm|a��H[<A	JENF�A{Y��4U�@�fa����5�~a/������̐h���w�gM�=):d���%T�}7B���%��"(��:�&)F
�/�Ј`����F5|Z�K�cD�2I}ק�Y?a̕��KV E�p��_'��e_��XQ�v����o�i��Yc�D'����`%� �}fQ����n�'��?����g,CyQ����@�}��a���\,�*�ҡ)s|�1垲dz��{H�G��+@0��<cS�� �'K��J�19�=�"�`0[s���K>���0�B!$�ɦ�NNn���fےH����>�5y�G�� ?%�G<�a���h�n�	M�9�kCpcV��x�ܑ_��)��p����f�P]knEB�^#�,�1�r�	\8�E���p6�����^+�����j�w��_�Eԯh��?z~�S(����2�q#��HzAn��i&�P��:D6=lM�<O�V�&�t�S>�+�a`��>|���d�_y�6�Ȋ,2N�0��'Ζ����ZC�E�-��m���ën$XZ��	L�����@����Y���H.ONt�E�U+�0����L�Q��	��׾[�#te�l��7��y U5&� �s������_*Teu@���8:u�Wفeٽ2e�D�̏k�]
���-q�5�7�X@^<�Y�Z�e��ԙ�C:T�m���Y�6'���VZz����N�s��=&���ܐ��s��*>�˕�:_=�r;�~AW��`L̹
o��'�cq���&f�f	��U��d{K�����s�t@�� � �Uu��e��(��*��=�_����gm��fH��{о�x�BKɭ�&EmM<BwHF��˽7�K��M/��;9_��:5`vZ�A�vH�����]��Z�0�W�&Z�n)>��Q
fJ)�t�l��6l���E�~r�B'�&�g��it������/��!.sL��2
;&A L�	��<�z�I~�0�R�b<��;�+a�)��V�҆��Z;���J�Nk�6���׃��!\i	úӼ���1�/:��[:�J����T��3>��\p����=�6�B�/ڲ�βtR���O$P�P����m�)���Ҋ�u�-2�0+�>A?T .[�Hs{�$���C��#VR搌<]_�?��]t���U��,r�R�&�Q��5x)8r�0�W�~F�CD�Aڋ�L-rK�NKd�k����7w/��w.�M9���w�59Zya�*�����-�����/0���^g�/�;��*!�E0�ܴ�B�Ո��e*��f�/�Ȼ��Ԗ�v�LP�&�?�	��*�{��Z�N�`�*��͋�qkJ�$s<#����vm����\I���fMv
i��t�->XU���e>BTl��p�R4aFi���#���\���1^=���`�ڬ=�^��������2�,�+s��x_T�)�ʬ��%���smGϕ�ȓ`�1	Rh�p��Vͦ?W$J�}	�Z�aH),V��h�����ʙ�T��8����qx��a���c�&��g�z���&����2A7�3~�n$M��p�Δ6cy�&K�d��G��'�M��Jp��G�R���i܅n��k��������В� �-�_Ɂg���5� ȕow�M,}>��N�v���y��c����P4l�x�mflz�^N����
�!���#�<O�z�	$;(UD(2\������L]걼�i���7��j��k���J�[q/��'�s+/�h�%|�E/S2��eXD152n[W�и&5t�W���&]*�Jo���v���Fމ�����8��Jŉ�Juy�Ɉ(�v��Ԯ�؜��6���?����������wq���Л`FS�CS���(�5JT�4G<dE���@h�!�F���%[�ɉ3�	cq�a�U�Q�\�ߋ�o���~@�nH�����%M?��]�?���.��@y�:���/�=M�zJ-�t��81 �Z�� �����oJ܍>�nY��؜����V/R,�8�G{��p�6�-f��Y�zK��S~:���.X�N\��Zve�2�<8*F83��V�����ц;�o�k�1$-��TEҡ�;�����@�U$��e{��F�Ǉ㕿����ۅE�j����2�g�w/������w�hXqZ�y����K�C��7F�����(}e9������?�2�-UF?8�:�����$�g}Y)�ri�B�GO�cf~2<d�Ml���OS�J7��e�0ggO�(����q�X$��cqpɦ���͢!�����@? �J����@
ִ�sYOZ�����h�y6������	�v�LV>�ﮮ�p���S��Sn-���V��H�
E�!7�����π6ԮM�Ș4z���(�H]X?&o�\e� �����ϑ�V �]�|GIX�e��(�|=u���.M���1�1X"�u�'���V�P�L;�<�VX�k�
Ǚ�6�4��k�ͱ��+r�s>��%��#'����l�q�S�Q��,¸�H�*'�ɉ�2|��Q�b�8��W�̔�k�ְq=5�^�� �睫Op}��&�M����K�ʜ��/�����%;��^�נ��W�p?�a�I�:��I�,T[f�(���\��l�pL�p�����u�tH��`C�ƣ���+0�m��&|��ۈw �P,����8�w�&��r��'�+��ec���9��i�)7�]����hh�5�ɻ��Ȍt�3 ���7�i���t� ���-�N���Ic�H���Q����H��C�� � 4�5�]��duB��"�:�R�
��;,lX��U��X0TY��e(���C�?��A�&��,�l�4�s� jlr��6Ku[KPL��Hmp�Xf�P�vZ�/��T��d�l��8^
���t}P�Z�u�Ť��D���b=v^�]g���ZVb�0~JfCy�w��h�eh�5�~�Cɍ�'rQ0�P��I��><j���x���*^b��(���5��U���6�qf�w����^sl�#�U6x��V.�
�u��Z���8dI����,h��b�f���bo\bp�1��<���� �4�jHK����#����p�ʘ�MU���cb���R$4tK���r�kK F��u:�:ħ�x���Y�N�}�Ɲ(�{D�x���ԣ�9��v�<4bc���jF>�@t��{���H1h"��o�x���]��G0�0�����.��������O�Ꭰ?l��t:4�è�0��ʺO�������\b]"�Z�����naMP$hL�+�6�'��g_2۴��N�UoH�x�hIJO{�6�<x��{��I�����8+�� +�|��K����5�x~�<�4�m����Qc�K������D��~�!SC%t_]�`?/7[Շ-zK�-,�?�p:�&�n]`5k�:�v���jY���݈:.����S/�s� BU#rl�{�b�ʮ�o��I'� �;/\z����(��I�RkK^ޏ[?Y���t,�sd��ˉ�����!P)z1?fORh�a�ׯ�O���;X�r��:��#Q�+Ywc�pb��l� ��B 6,�M���E� �q��5L��ώ ��4\�����D��~��#���Κ=O ��5q-�� ��@q߇�QQ|�]hX�w����m�I۱�v!XoM����ː�-�u�E���S����z���k}g8g)e�^ǈ�ޱ���]PT��y�?�f�mg|��b���P�_�"�8��.y&��Cԡ�t)��1�\�B�I��aM��ğFE�`.����B�n��_��ΰ5�	·�Z7>/>4�A?qC�Y���?���p.t�:U`�f&�g��g��E�5���=�LJO\��lء�Ґ��,ø��]J*���>3�k�P��+�^ |��Y��=���R؎A�Z�$e�b�h�����>�����GE�;l���uָ�#���q�x�:�U��j��Ԙ
qO9�s�[�+��a>�`�>[��U]�Z���^�|�w)�8�/~�ݸd�qNd���S��~:.%�`FMM��~���'�-8%fQ�Nȉ���*�G)��K�A��RE��kJr'��?�$�*�i���4M�j�;��܃L7\�ȭ��T�tI<�"�����v[o�������.�e^�_R�=I g�n��Sp4��1�)U�ݬ���G�9��:���8��1���f;�b/l��\}�5a����Z̪�V�I�yT��8���+�����3�:=ПT��PU����(��N����{vTиC^Ts�&Â������p�糽jG��ؗP��)�0I��W�c�K08۔�����y0����{�p�U�Ժ\��zY�]����~����]��m�A_�)����[�U�\����}���!Mg�����q0/m_!��T!L`���,,��}._������hy~B?�ɣk�AQ������w8�U����Qȍv��F��N����2�P~c��S�v�h|`^�訫�e��ɻ�^�F|JTp��S�i|M�۝d��Ȥ~�,�����q�'�%8G�b����%q3"�8lYo�si'c�:M�k�����Z���R#�Ix�.3A�k-��Z]HE���!N��Wq���� )�D��~!>�ʱͣ)x!��!5�rT>���~x��ɖ8#�����ĝI�]�B�7��uT�$����̷��D8������?������K��<ٲ2�o8ߪ",xj�"����D�!G�OǸZ��
S<f�k0Q����Hx��>s�0�g.�Q�]��mI1�K+�3+5��߉���s �O��B���!��v�m6yP�a�u�֛Ų����1�p�w��$5ϨkN�]��H���gH�z%J�H���A�e��-�{ߙb:������K��Մ0�ҕ/���-�l���+�?`��"�9�j���� ��ߖ-K�
����;9I��y@��<�8�_#$����b��V��Pӌ�	�A��	�>�Ƹ��Yq��,�(���`���4M�VQ@�8f�1��
`�B�orW��U/�E�4�0���)h���X�R�t޽��r����U����3�(���7�VY4�@�Y9�ľL	���$�%���}���{�<xb|�+����մ��_�kJq#��V4f,i��O�w�"���G� �Y�4�W�Y���ܽ�E�Mw�cj`|�U�T�y<�XN�q�_[_�íϵ]�a���5��F������RO����� �*[-L�2Zь���	_�aS���L��Pۺo�&%e�Ü��Ϸq�Nd����d�B���L�8bf�0׾����➑�AA+f��۰/�����%��w����8���_���\T͊ʥ^n��D���VZh(z�sz�x7fM�}L
�,J��h��$O2��/��*���>���/�2��%Kż$�b���C(�R � Z�
��Tw'\5��/���S��mx-N_-��;�{�Ϟ��R~� A���g���o��ʵ��G����Du]�"ż*�#
?M��?���J�Qut-�)ô|6Q�~�p���7N�`'G�bnS1��7>�6j���f�i����tCe����=�(��B��anN|�������bNR�֩I)��e'��_��ȃ�=[��Iۖ���ؒH�V���zQn&Mg��;PS����M���m�Q2���yc���~��{���*�S��+�l�2;]fE&n��ύ�	0h����1��U�\ȧ)dq:!�B_0�&�����+���4�"3�bJ��RO���s8���6�q�0'I�l[2���Ieob�hǡ��WE���Zt��E�'�O4)K�Z?�N{��T�p@$QO[k�R-�d�}$@,p���4Rb>�i�G���)�V6�J:�Lch�[w/�͙��M%�9
����oaXdY[��������%]8��E��N:��[U�\��u�!C-Չl;?N�W�1���y������,ul+z<̪�5H�R�y Ur|�"fa���@GT�������%�J��m��!-=Jk>g��ڑ�4����R��b9]����N#�/F�n�]ؓ�i������C�`KG1��`1�z�z�k�n�3�sΰ��aaԪ1���,�酓�g"��b�$[A��N��\*%K�{����"���������2e/������j���Wd{�
g���t�C�&nUM�����n(ͷT�?ߊ--,δ�E�v��4��N��x$'���~u�Yq��Q�5|��70�����D!)�B��_�w��s^>�)q��7�Joo�n9�[a̧O՟�V��jaj-��42� ��96/i2�h�|�9g����#{�b�/L����!���f��' �	4δ��]�Cw|T�HCG�ޤ�2��J���3`��E�z�N�B�}IS��n��"��ZO9�s5���C=K=�Y��P)��vLCۃ��5w!Y�%��nF����`� ��3����G�U2�2v� �~�O�<Z�D�+�I�R[��_
�fqٶ)0Se�hw�]b�`��a|p�G�ڽ^�v��Rʡʞ�8��l4�����p�l��t�|�rϵ�8��3� �M�ƽ$R�2�ek�<�U��!�ZS�ngՏ)����>P��~Z�@S6��u��[K���J�UR�ϛ'��n�ސ"��|���o�����m1y\�9*�s�Ȫ���U�V�G��T]��K��^z����1�^�N���	`�gOﳩ_�睄φ�����b�89��4&�碶OPg ��a?gE���s��6+D�����7�w�-&fP ʨTYb(�u�w�IPT��T�(�Z�L�X}�1��e.�&$k�2J��$�=�Y��kؽ�k{�UX�|�G�����z�]���y�ǁT�_���\��ڎ�t�[h>��bި��MXrx��?�<�4�����B�^H3��c���Y�]��{ �&8"j엕�)|WF���W����Hneuk��>���g�KJ�v��V�Ag�ȩ$�Dk�kd��0k�~��"ε���ܓqm�CX
q5J^O�NgXzj=7�43-�v�p{��F&���{�<����.��l�H��"����b\#�kk�D�T�ĕ7�Ր<����`���G�`�g(�����X�˗&�L�{��H�|�^�DO4Pa�qGO��;PA�I�.�4���X����ȱ��"�M��ؘ4�}�w�[�w�6�澎��Q���ԅ�7:`;ZW��(yr�@��^}��uaJ����ď���Ђ��~�M�nDT��A�����dH���/E\˥<�:�/p���z�^@����.��VST{�/֭v��ap�,�.�R�\�[-� �|ǜ�Kv䘚��D]��r����H8#���M�0�R��X�K�oHȑ!)$���si]Y~���ѴE�DP��U0���b4�縠�m��?�ٞ�~�����~�Co��'7�]��K�y�x�"���)%^sj�3-ꃇa�{���\�׵�(*�m5 �Q�9�Xh�B`�$���"�qp�ڽ�����З4��&��<=UM��Y	��<b��P#jIdD�@�{N�b&��P$��L#B���5�i���	�R�h��
iI��i����`#c|��Ms��.ߋ`�M·�#�k�X��X��V�ǻ�\���I��C�DF����%0�]J$}�йJKy�Z*������Lz8�:��;�)��-:m�6��@8�9�E�Ǌ��~�~�_�lV�~I��l4KNkҡ�>;8QSdτ�W�'�f.|c��60���"X1GSt�+�w��{����멞�œ�,Η$hN"]Pv����ۄ+�����Q0�>�2��
v�i�_�ʖ��_-+���B��4����Nەy�R�?�9�"wο\�I&��mh�>3���"���������� ��8ܙ�� a����ũV&�m \�w�r(�Z��6�(<tZ*|]��\rۗS���h*�!�[�\�4��#\M9�l%�_��B?	�鳵�,{C�16n}��*��	u��aG&`G�;�����zؕl1'+o(+ʄ��������_3�OqB��*待;L��X��r��E(���6����f���BL��񁧁E�v��iŗ��W/�sa�$a
*7s���ȷeŤ� FFT5�]�l��֘>����St�l?�]z�6`Y4)@�Q2�l��UR0�C�B,����'�D�Re�<����b`��N5�l�\_Փp1}�Ѻ-�$�,���r�E��Xns��-d�Dl~j��>(�I����Q"���c6�Ba=�)$�!���)��E
#���O8��� �$2�SK_��+Ro�6��&��M?.��� �P����MX0TcA&j�"s�(��u����;�d~nY�7�GA�'�k�I�x�'���N,޽�d��AUK؁z�#xQ�)}U��,v���$�.߯ܬ�m�R���~��=%����^���T�U-:ޟJ-����|�5�L��JF����܂��i��JD����X ;�("j��v܂��c|��tћuL�n�?0p�>Uc��
��0L"w��$��E��LZA�������9>�ID%Ӓ�
�«#�:�9[M�&�pg��(;<iM-�2�U�����LT��D(^`=�{���Bf���m�6�U�p㴓DG4%1ZC��q~b�<�hJ�!a,�xOo.��� v�CJ����*��!�ThJ�EٶK6T��R6�A��3N�?XH���J�JU ���fyx�'��ٔ�lEX����!
Z��koO�b84�Nx�l�'$j�[����3;\8��QR�����I[d�4�l��S+���߀�ܭ��C@̡B)�0�G�ȉ��BX8\�591�y��9���H��[%�J��	i4kReB�t��Rf �� �(Rjr�!�w;)��W�Ф�0���z6ň�|�U�[�� v��rҋ"�
X�� ��u�س%�1 ��I	�B���ı�S�q�����	�81)kn�� �i��Y\��R6��|2��nyc����j�ǖ�g�h�m{7��>�ne��nV'L������Of�	 ��m<W	:�R�;g��R�4f1���!�K��paBP��ƫ��)��g,�Z����}�E`�:�7޴� ��"I�:���?�4���Q��2feY�=MCS��u>ʡ�7��6ӀV)���[��=!�7�¬��ze2��(<�j�u��!�ݤ�5��:�z �+��6���v&�I�"�c��VFT?c�ܱ�)�Ґ2yՉ>��Go�ۑO�A[i$�Rg��f��9����ߑH|�����<}����L Aw�.���G����?�5;�O�ù��P-Y_20�����;�4TC�4L�f]�#�8�,�Ĉ{�C}�=��iZLŅ�B���j�&��zS%��ޤ�h]��������S�h>zl@ZJrW�߶��0.2P �?�9[��.�8��X����?�}l7�T�,�5��L�Ӭ!�>�I���:B?V$�\7��:�Ǭ?R�p�b��L����0���HS|֎l�ccH�¢F�id���u�fZ���c^v'z���ߨ�f�*#����ݻ"�zt�+Tz�:�R 앴q��ECD6�������s��d�8j�ͷ�qK��A�n�h�H\��S[3,��4P�p��s�i�����1r\]�y��'�jH�I7�j��E���j4���yu���ɉX�j"J�DͶ(~�^ݭGBu��
�>g|Y	�@����C�\�2�UP+g̓4�O�0"����n��n�J{})���oHV>L�p���a�6�$��xw'���FSI�r���iqNFZ'.�8�2k|[��^���+� �@L-V@���'�r:O�k�J��_������?�1=ϭ���-��Ulo�ۼO~�΃)4�b�1��g�w�2k�\�#ǁ�4���_y�N缾��Ӥq�Lo1]�`�cc�<ۉ���~D�D� H�ct{����
�_�1iò����[�Zr]B�͇�\��^2f�@�©wi�{^�`���'����wg��#'��ԗ	�Õ3R�mV��7*�EEJ2?����v���J��1���tC��J.3{�^�Я��k �pS���+���yo lݟ��f*����I�P�k�4�+��@Ab�vh���I�H�Y�QW�&��{���t�h傴���O�:�n���~j��8׫>��F6�~.�8?5��Z��Ca�B���~�*uw�Xha�@tr���~� e���ܤ<�R�5H ��Ч��J,�T�vR���[���>���Ӱ������#�k��5:��o�L_�k6��CҰ����c���
p���Q6�|n�lo���{"�;���5��4g̸3��WS�"/�ߧD3PëR�(W�8�\��U,�"o`g�nM+H����V+��Źb�|������h��L�g'H~�h��^�?�0�~����o`� <*���`�*qe���+�N�E�Y�wn��'9&�y�6�s��ն1�ac��=�R�:,��;:����j9��}}K�WݛwkTQ���>��-"S�_ Ra0u)��șKMU����&h��cڮvK�_�L�� V��2�z+ݺ��IU�4�jU�a��LA8�`����#ޫ7�	�즟��o�&t��Ǽ�#H� �@rN�j]�^ß�l>%G�l''�xL��>��]���l���f�_2�%�U�|�痥
��kYs��XV��=N~/U��O�X��Zs�f}	���D.9���WF7�ʐ=�8?��]��,q�~���Su<��*c�'�����	��N!�``���j�{�;w&��IR�������;gY��
y.�/��*/�z��4�%���*�s:x�x4�Q����|ΈX�(��@���L.�e>���++�&�Z��*�5�]D��g�R�>��l����M�<���2��yI�p"�ߦ�'2�O_@�� �"&�m)���ɪt��(�eI���8�������-5�&X��f�%�����n����h�`���w>�� Β/\"z��������
?�^v	���#ɍ�W�~(���ak0��0ݙ�V,L���dz�~h��,�)*��t�������̈́폃�����c��cb�BN)Z���)����Ԁ�v�ܲ�"����gb��$4_=oYW��MK���e�2/C�Z;8����ivc��ʃ�޻�o�5��c����$Z��]4���h;����W������.'螸��"�`=DD򁼖����t��h�2�}��FLEH
�Y���B��@�#0Ǝ�p��u#� �kD(6�bA�6V�yCd��~K��2 ���ٶ��4�k|���v鴶*"N1.�K�M��jN0�W/u��Y�ر~��r� ���?}v:�u�����������sB�VN���T�٬?�_7�����Ls��Ӱ�8�֎�Ϡ@�'�@��E��q��hO�.u���v!*�\X��PcB�{9-����5׋�����ϼRɂy��!�-|	#� �'�y�r�v :������QATT
�_f�M܍o�L���΍6D�c\� R���hN��W�2%ᴯ*���)�,����2��|q�1j���K�l��jY���6uTa ]�U�q��8�	_�ܱT���X�}��.�ʊ���M���lӓ��4��k?ʳv��0(Y�s���KGy�� �����3k��:��QL���ދ�ה���:��/���O.A����_��ތY��	�x� -y�y½���)Ё`w7-�kt�� ��A8���fP'4 �cAq{��A��Z-�1�F{(��wZmo���ol���B��h��#xg%O�Q�M�{��B���S�nM�4�[�L�����*���z�*=��hA�GӵUxI2�[uN~E��y�0d���~�����'�Rg�'n�]�@o�?/v��e�2&4�����y⮄�iR�Ok(�������E�p����Ox��y�(·�Hj�+�X�����Lyy�����횕*�����m��[n�l-��Xz%V'�&ky�6���$r�6�{,��ȃڋ����a�9�{�0�����g��#�V�y;��ӗd~Q^�u�(�����̕��haF�}����.X;eb*h���
�ǷV�{�.����s{ �?&�%t|.�,Tq&�p����2	{��s|���gO�?��Z	d�KXp�˘^����n#aC�с�>�ݬj5���4��PV+ޞ�H�H����M���j������� ���Q��!]��ɉ�Ԁکfⱋ���֩;��җ�J�Wl�����lH%���t\@{s���7(��֚<AZ�t[���|~��0[1d����up����o�����Ҕl�nS��r�-$7��{]k���_�d��=VI�^yIHv�<$�o�4c����xr���ׄ�"��˙F�:����!6Y~kT�M�p'�<�� ��¦�D$/��h'v� ���.]#�h�o蜟�����X�2��#˝���	�m*o�`S>��_���o�/���	c�#�D[�k��ʴ�$��E�����ҧ��'�T���l�r�e�|�����K5Sg�ѭ!�֖���\�J�	�3;����2�6���!]ZX:%|�k-U�wá�N��m�G�65��G���?kH��X�ѭ����w�?T2�� ��@����r��ˣ������,�ؐQ�!zr�-ֵ�+�|�����B*S�#'�A�����N����&��`�MŒ@v1�2پWv�T�f��#^�ҍ��^a�x�o&Q��ah��u���Y��_��'�������ݭY��KX��;�0�{����Q��Jy+�11&Bϛ%�&�~}e�`�MK�!jv:}'������CUDP](*�����(�i�4�\�@�6	&�~��~R�N���
d7�����)�KB�y3o�_U�1�)@�%�Oa�X��1��a�Ů�a�=��РxY�a�N��~���T�������p���
v�M�n������������y5;�I �>e�F������U�������"Oڴ>���8�˹��A����<^����)���L���Xj��ޙ�	 �淔
���7ͽ��0)ċ
N�mYg��&��@b�dg�2��_�)�X0�`]�$q;Kj2!Z���	���;s�?�O��F��rXث����O}J��X�#g����"�·N��\wuǼ�"���W��'�AQR�x_�|g`P��e�� ����;(��14<]���8�Sv�Ծ%h�o��z�4/T\������|�u�'ŝ��JE�X���9����b��*G�DMe#3��E�/%��"eP%��G�N�(L�ХJ\��wX-_R� ��fɣ7��j��$��Y����(��r�~$�T*=tH!yH����x5���>�#o��t��
�`fE����'n!NE̤h#{E(�o�&ﶤw��M�����r۟�G���'�#�V�xHn����/-�������D���~�F�:��g!�۽�ś�����2ji=H�u6�S�~�Q�&���0D�tX�|W]��!�f���uAR��ר��)J��B:�{���KB���A���V�e�]�Tϛ6�g�7�KIֳy�3'Lض�������#o�����w��X]i�Z����#�R"����%��8*�L�7���8���'�yu�5_
�k���W��:T(�آ�X��loZ ̟ԙV�`���ͥ��������0;4\���/����JZ�=���O!�[�8��[S>�
�I��m�ɂ��<��NZ���Q��ڳu�hb������\��~�o��ݽ�j8��b���������F�k��L�ET��*�"R]�Bj�7U���:I����w_[������#�(�@@�UT����tmv��P��p����Ჹ9kmo_�^��Q��8L���Vc�k;4��\IS���3-�h���Ir;�c��q�
1E�!@r{�N�5�n���,Ɉ�1�)+�24B��$&^Ύk��V��R���m7FXG���1�������p$��k� �@�'�'jE�FB�������G�E]?����i.���r�G\�Q>�O4��&
Fi��t� �κ�*� G���G3�abй�e~�8^��ʖ�������x|c�|��B�p4��f4��ڹ��%�I��@�FAa��UAg�U��ľ3ʓ��]�.���v7��7�q$�Y<��6�%��:���x���;S�N~
�#�mn�&w��mJ��Z�c�S3y�D�	�K��'�UA �!F ��M,G���*r��E/���__��6��"c����}�F��M$�+9��ݸI�T���qw����\��s��S�.$?P3&ߕ���T�r8��ބ.@����+��m�z/�]r����g�j�:�u�;C�7wTQ�\��Oh< ,�p��K��1�6�F>U[�漀Rٳ���� 6C1�	��[�����L&�f*؆j�hm{��`��z�
��>�r�N�Q3����F���Rƙ�+�jY����)O3��0rv���:��g�n�r�s�u�'De�_��O*�(�͔;E��gӰ�K��otvH��c�#{>Ln��!$`z�J����^ygA����.��o=�u3s~�g� 3#��I��^��cWYB�<52�,��h|����9V �	J�_�F"z'���b����i�೟[Է)ׇ\�	�f�)��a/84��� 3���+u�6�R�Jy����R����As������g�d����6�r��U?	����1kSKD�1��.�G�J������4����R	�@{,c8C����F��q�5��/�7�ں
�ۙy���F�n�߷g����
p ��<$�3Z��I�=I:�v�����~:���A$z������II�g1��~��j���_���;?;��y�I�8�!Y��`�����zfc��es���N<�^�/a��[V�`,8B>]�f �7�=ʌ�Ry��9�L,l^�X���"���{7�J�@}�^H��3�CbnY�@guY_��CeHu����53��jQ�#��n5�_��1q�;�1�:%i�{���Rx��LU�Wx���uo솖7Z�>ɞόp�#� F�R��r��~��v�z��}M��������M<y���<Η�M��ډB�8��-Ӎ+�B{�u��ߴ����za�kpӨ�0�u����i�+��R��ԩ����\�.�M���h~�D#Hkm�i��G_��U)�����Fƛ�%�g�k����qE&l���|�zҬ�%E,�F����۽��`%�f]�$�Y�iH���`1���F&$��{^��<��P�	�{��"�[e7h���^���U��TPH�2ߍ���bp�+��I!���~���m���G_�S�Y<[��{��Fc ����s�x�L��b�����'
?� �Y��K�|������ay5�5N�ҿ��/Q�]Y�����ԡ�ቪ�$���z�����]�|�a����Z���/@�� Ƚ�*�Y�4����'�z]��i��xMo��~������5��/EF�"�L�6����ǜ�͛�ٙD�[��ur)�q���m�Љc���J5ɢ�I��ڡ�3��j��H��C-����iǌ쩁t�w	��g�f��:�D�����W�"m�Dh8�w��0�9S7�O���O��~K�qO�<@9��e��m������È��,��`���96V�L 4�[Q�X�S�^�t�����&�T��ZMB��-��L@�[��fu	�={����'��=.%�P�/�h���Եh8rA�[�6!D��[|�����!�.x�N�|8�w���TO:��
>�{�i�䔦:�/���׈��&��)@�K���G�fˆՍܩ��.��5��`����F� Z��F|�@�-��O|J��oyY��>�	z̫��[���9I�-@��WNˠ��=����욯S��нR�ܠ�i��MR��HE��e05+�\��u����B����+�ڙ��
��#���3k����Y���e�)_���-��)"��j����Q]2���O���4 �ܴ��A���=?y������'���=g�e?�@�bM�V�?7�e��a��7�um���1򒤦����r�]GX���#��Gw��<��m��q�/P�h���ST]5��W��mpgDd8R��ގp��ļ喇>��p^х�g�5_������j׮g�7�Ey4��\�p��:�j�Z��I0�=R��h<9z4Ք$��Z�v#V�?4�~~߇g���D`|6�I���`W4B���زB����J�:�˞Pz�05 Ml�#�:�ha6�$��΋iZ��R	���W?�o��8�,W�[�e"[t��=�=�c\��!h�˚m�̝�(�O�2L�GF���z�@�3/r�J���Z�a�7i���۝�s��5K�UY���N@y�۫��-��)q�_���*����I����I�R�4a���P�.=[�$ �M��פ�NƳ�!�]Mo+�ϙ�Lq���V�8��B,��N(�o���1SM�t��X�u�+*ߟ��RVY~�w�&��ӎ�
S�kePl��0�\y(BQ���l�s)c��^���-opb�&Yl$!���ݎ^��������)db+^���,k c��'B�jyb��d�
F�m6ty�3��o!��~�/�(5��-)�9��yv}m�����˶v<f&0k����c���e�5�,�� k l�A[�PI�&le��>�4�%:�����5=.�}���:��fW���Վ�
p�����3 y
`P���������)���cbwFm�T�)۱<�$B� 6�AYOx5g�4�����2�ޮG4�C1���!zڰR��Hre9�4�Q����NBt�0�m���H㐲��kf�Vî$8�����,��"0�<���9�g\}-�����h�ܩK�(��r+�q�kh����u���~�g�3�� �1�OFS�sh,��*�2!k������`Z7IQ�%�"� �g�(��Z�\�A�(��i�9�����*�Ib6e���b�Y���ɓ�p̴e��?���'#O@���	�ҫ���;w����V|�6��hM�Rk[����\B�=�S�U�G�K�h���5- �p�%JFs��aZ��J��cg�ʿ��+r���ኦ�]����`We@]��*f�q���)�B�/�5�S�u�#� �5GD�I2 ��`-����!�Ⱥ�E�A��n�����o�3LD�a�=,��?&������|�Ų\�xs1�T�=W��w�a���9������L�z����v7+�ծ!��u�zS���IuM��Hg��IS���/�:TH$��������j��Č��!�R�Y� ĩvus(��yQ���(H<j[�`nF:VX@�
��q�w�Ɩy#N����J�5$��a��˪m�����g?���(Ua�J"&�h�"��.b�Gz+�ĵ��G �eDk�@h��L�DG?,y&�l���&�ʪ;��n����J�R`#I_"r���,�w��^L謜F��#���NP�>'�|B�c|v��'jC�g�������a48V�(+�լ�U��m=W��Y0�>�
���0ՇxJٓ
�@�۫��X�ϐ��4AN�q�7����T�m���@���[L#����n\]�0t�t�P*�V������HF �AHh��~\��������T����'U��g�D���wW�%Ud��1q��:+�^J�ъG �|��5��r����n������>�)_�Ѧ���y��K/�Fa.����42��H`7���ª�E$@p����Q[�_�P��b���׃wyZ%oxo�t�9��3 }򶩾�I%/%�~�	_��ǩ�t��%���?��5�\x��O#��+�2�p�]�95�v�iC�2��y�������ܦuQ%�{T�$�Lv��i��$bQ���h|(6�1^6�x��#"I�$wtM4;n�A�(�
��t@v`��,��&��~��{�ۑm�N��תP�G��5t� G_����ܭ��򡘀@'�����vw_���]�1CT�� �cĽ2$mP�)�eP�*��h]3:���lW��Ԙ=��1�c4�OJߢr���-c��޲VAV��A�0j����o���n�nܦ�;k�Nw�܃���������32q�~B�M��qY��N������F��u��g�� �:���~���h�C2C��]`���i>�EMȐ��oC�-9�We���3yީ�{u��a��T6��J����F�j��
q[����o����׫=���x�ч���-�5�}���#M.�WR��U��%��~�Oϐ$����3��(ʾ�rFW��ac������9���&�u?���;^��������zY��E�.(�\�)
�Q���+�ʑ��T�޸.�Pڶ��d�cù�圹\@�2ŮY���q�N��2LY�ﰌ���A�Th�R2% �ד����K���U��w�	DR��]�D��Y:A��?<N\����#y��'�ԕ��.��~�gw�l�]���h����a�����tr+�z�	��L�E&��/ �/�1�B_��9	����XǼ�V��s� P�-�����%���]b���=K��+�K��%�GvI�R��n`��
2���W1^ah��@�qa$x��$��S���m$-r����+��!t��UJ݊q��~ƾ�_�_i%S��hP'q��7�D�Z�.�7��2İ��&Ӊ��:1 �B����[4�n0����<�;��y�������46̜��>�s�z3�&>H���a�@�2*E�x�Vdl�x��!�C�
(�o�2����	A�>6L�������s�y��Ȧ3���i�"Dw}��"�wM`��M�l2D��'��cG��H]����R�?ƙ�L�'!K"��e���ۜ��0zJ�,n*�J� a0��!V�T�W�%p\9!�C Oƍ�����/�^F��7������]�hH�L��a=�P轸�4c$
'6����l�P��7��e��+���~�[A�.�x5�O�S��4k��̭H�v�� ��hRl��x�C�Ez���4F"<$��T<Ƃ�7������HR l�����������~wg�䘪�PV7���a�5�M8ٝ���l��1����`�YWʾF��ܻtO�v	;���Ǫ)��N��ϱ
�?-|��$^��#>�ڝqǰID� 6)�k���̗�_76�ڷ&�~,��"���t�Q�m�/B��֎C�+�Z��:��o9�^ 	��6k��J�E�rnzg��(���y�:���l���ju�X�(�n���k����U��W���w5W���~�LRa��>4�aͦR�j$�;��eL������WR�Dl0����£�j��t&`��懂�r�k�2A����c�ؕ�1�۶u����I�Q��͛�������=�)�����#�:���4�X�b��/���"|��ǹ]����	C�O�Һ S��uaボ,���^�
�px(����愆t$�1D�.we�&����~�c�Y��m�
�΍�<ys��iHk-M^$�C����/�Y�h�/�4�{�\��$iY.ֶl�J��>e� ����e����X����pg��%���Sj�tf�C��I�����po��c���ba�%�)��(ӌ����~ �%}��fbr�4��;ℑwǫF�N,�a�7�mX��%c͞hT�^zo�sjI&��hR}cG��*�a�r�E��>�\_��ˁ?�^ސor�NY�|�I����j��ᅀ�w���8yJ���u��j�L�͌F_t'�٘��
c��:`ݦ�\�;./�@ ��/��մu�Xul��5ˉ��l/\]v�fH��C��K�����%�:�̚M߯�6�	��'0�{��x`{��`�0*���P�ʥ �3r�hTmƬK;/mPnzȇ��_��g�<��K�n���z�ƞm��L�{]	EF�t}�%�-E�������ؒ�̥��Q�qv�眒3`�T2�K:sB����V�ǻ\#6V(�t�&:P�1} h#z�O�l-4D���#��mOΩ!f�3�!��'*�#����$���O����k����M,i>�����+-�ɡ�Z�>J��3�	� �c��W_o�t���_k �Վ�aJ.��XfE+u��.��V�����ߒ�3�O,,��9x�:�.����7Ќ��#Аa��'����VRL�p�NH�H�(��ҙq���)�`c�5 �y?�2?T0��\�w3����_u�����4�_k��h����C��MV��k�љ��	�oY���ay���ef��L�qX�W0�*��q	f�q��-����yM���{c4��9u�z2���G0�_E�2\�8��JV��`G�&L���YE��+57��[�帨��}� ��ޣ��?T��@E�=�d���*	R�?���K�~�����J�Fu��B�]�D��Zz�գ���lKdO��L>�q�B���D�v`����.~X�Y?�M�Bagf��(�܊����d*���6��	����	�R�2s����G�.lV[P��|��-�@��c���P
 5e������1���p�
}����ځd�2�e/�fOʡI��8��|R��vB�K|J-X�ӗe�fwX��g4�|t�fZ��j.K�֗uu���4�S�@ػ��ٽ0e|��G$���Nw;��h��k��Щ�r�0P�7��<,X"����=T������'���!�x>$_U¿��1���iɂs���B'&�>g�5��ec��Q끮�Y��.?��o"NI��������Y�ѯp|c����Š�-��L6���>�E�����5�3����=y=P�s^���P���S`p|�� '��pMǐ�2���TP9�D=PY��R:�Ъ���LM�ˢX3��&����/��wHX��0(k���]�L�jj�P}Jc��&���D���ǣ��'�2> �U�(�K��W��E��	��I}Af)�H��~p����,km�TM������ɫ�L�s,�@�\�T *�'e
~݉�+�h�`kK�G*m>�Q+rW3�̎��ￎ��xw����ue��4H)v��T8s��4�ν�1ךW.\��]hqe%[r���í����+p�a��e^ ����g��Jϳ�6,�	!���|��v�&܀`Λ)L:#?��m-ӆ����<ʜ^s���/��x>�wd�(��|�2*�hSZ	A��ZT	ʚ�gi�{���߮je��8�f�̥�ݗ�����<��X�.��fTjE����F-���8�-Ⓨ�� ��T��חZ4�ꝠĪa$�v�\�6��|���,UQ-�9�~g�+��)O9�$���2�6'�Eє��,��E�8���i6�T������GA��g���T���$�L���
�p��g������Q�{ݟW��9���Q-�wSy�(W�?؝W@�b�M}��;n�M")�G$P����3f�3�'b�C{
3QLq�w	^����}���M_�{N�[�%����.��^޼6��~����� ,�aV��1����gb�W�� .v]/\�v��/� �"x�`���L58��!���],
��r�\=����{3B���
�8�}�p�k�J�[���������!4k=	�lJ6	G�`w	A�%��r����#��:ڥ��R���
?{Џ&K���TL%�lm.�9���)��T�V_��L��Cb�(�P!��Km��/���K��Z�lB�8�E�˃�h��^Ѷ���ΐͷ�/�o�>���9������>�T�g���DP=}r.���p%T��vd�K�u����_��k���/{�@#I6c�L�?ЧT��7�4C�cҋ�|�x|]��Su棯uT�6r.�$��묧5:Ò62}m�@=)|�?�?5J�Ġ�X�Hވ	Ĺ%Ѣ#(���lP�꫉e��Q�ev���>����6�ȅ�c����Q�"�U��[ߞB�*�S�_����Y��uݓ�F�fH��Sl !p3��$��ߩ�]S� '����/2X��@a�4��{�+M$�����Q���^]?����d��@&�F������W� �uL\�)t}+9����$�E=�,+��o�~-�-=qz�A����@�p�ٿ���R���B�!bA�d󞕼Y`T��.i��+	�]@73 �yCl6 *����z:���E"	.Z�6����> �F���r:ݧ��ڧ;U�L69N�֩�'���$8�"��C�}-ʜk�J�H�Fd�X_�b�K��)!h�s���k�-�~ac�0�>XB��rk��~}.7�
 Ƿ��l��l��8j�������ߚT�7o1YO/bac���yfF[/�ps��hA[�i6Wc�Y�y��`�y�ːܨ[�g��0�R1Y
>������Ԇy�8G��"lg��6FS*0!̹+T����֭&|���-#���iX��`"q
ݣ>%�����Y�;��&�����d�	���T��\���u)������yK�%�N�`�l!T����{���u��L��\S�2I{���z3i��U������7��P%�]��������2�.���XVo'�~-ވ��ݲ,A�����z�$�}�4��Fs����p���� �o��Q�RKtb�{�q.���a3E|]��$41��0�T���u�s����Te���%8�l���ڙ�H�楂{�~*#��M~�$�g�}2k�CM%a�c�����!e3�H��+�yS��#ZBvQ�+nƟ��̜�9�i��2ԭ3�QH�,�_]�P4P-0<^������K��^����5CU��+���L"zf̧^ІH�񍬱�����6�Px�0�E���9k*�����|� }I���o;R8�"'2��`�����%:Ԋ�N�7Io�e���{P�l�w_H�]/��E|Y5��E�)C���@��%��}�V�t �����4ї~�Qp�'F~z��U��w3�u�n�(��w��~[����<���O�����r��g�@`k�I���_�
,����G)��F��l��c������-!���q��O��2�C���:��`�h�KQ��	�8/$�8�ahے�dI��M�b�t���3�V,/���l����!�-U��'R�mP��򾂮s�[)�J�We����9��+���(���o����IG��Wc4eu)b T�t��e�â}E��70ku��Eh�˙���,8u����Y�gK�X��J�.��}4_x|����,���`� }�\�~����B/����8�|�DC�Й�e0�i�G}���ʉMnj�\��8���c�-N���U�k�YE-HC�~bT�GO�ű��_�-��Tq.*_}�~�we���6���<������!m.�Z�΂�"�<(-�4%;�K%M�x?J|�Ǐ�EBY�����!�$��)g�:M���CQx����{��[SFC;[�il�g�J�f}�c���w��j��S�&�����ғ����%�P�x���q��]�11C�p��6��������kWr*G�!�,�^}x��L*���k%2����ގ<�y��du�{�+w5�{g�6���=�'��l9�c><��a�itf��"�Z׋H^��Z|�F����>�,�#����+/q(��I����%󿁲1 ���[Z�h;<��s��\�͈�J�&�"��U2��X�x�C�w�ޱk+�xK��nP/l��RGܔ׷M�5�� b�c�x3�Y�J6x�P�*^�n��~�M隣����f��Ki"���ͷ�.u�d8c��.�qˡ��P6�������bk[t�G�B!�8��ǌ�]�^�%ڤ��zu��T��b����@�Ol.B� ���g��6U~!*���.�	�L>�h��Cv���ƞbp�l	t�aϼ�!�������Z��5�F����;��q���Wy/���{�Zv�(e�5A��9J0�n����T޼��T�����:��]���Zr�bѤG��m��RkFj����[u�X���Si@�4I	�\h��0=�;�R�9�b��'�0]W��L��8�N�q��קV�����L���/���G���G'M�*4��IA�}� ����QyR�_�swPb�s�J�����J��{7� !�3��ڵ�o�ڭ��+����אhӧ>�@���f���&"|��)dN�+�bQ�veXv�T������� ��݅��l����󜛝e��� �4�p=_�~�\q�[��ߪU
�"W�I��)�ۍ*���t��a+��\A|g�D����/����!{C�����chx%܏�5J�@{- ��B�\�Ăh�'.@�q��gJ;-f������P-Ό��$�Ms�>����&�x<n������_&�/��@l~�Ͽ+a�	sUP���i<3 ���iH۞%�Z�d��nN�ԫ��H�p�ʚ�|�Y���J<y��`>捳���]���	m*����;��mo��:r��rz<��H�-�Y�7N�dgQ������ז�w����L|�7�4Ū�~�	�K��"�6�0j
�����2N;��C�U��I�7������N$1���t�ȋ�B��;��e�Q@��Z�U��fP�ɹ��>Lq�*Y0!�_�/U��n�8н�'SP+Ʋ�W��V�j��z��g��	G|��m���K�t�^�|F�O��!�#_�d�q��I���-㈠���Z�u�Qѳ����S��G�	<~�g��ͭ���Kˊ�i"��!�y�g]��ӥ���?�`8qG|�Y����O	�%Qp���2�H���(�V��}3|;I1a�@!�h����� ��s=:�=���&W���-d;��iS�2u9#����u�-�K��˯b���������{B-�-1��� Y5�,��E=;�K�ǠM���Y����s|o�����U%th����hX�n��񥝥ᙻ[y��~��l�I�-`�d4z,� Y"���3�����J��0>�>
|;^Ɋ��L�}
�8l�Jj&j?�j�Y��ǌߓ�!�&#E��!2@���o=��]L;���tnT���(�ֲ��r&o�h�+��+-:��,j^�wQ�%%��r���{�h��j�UW{�vnj��0Sf�%U~�UzY)Y�j!�@�-��~���מ
/���Tт�H�^v�o�H;��#-Ճ5��(i`���r��(�+�6שb�Sؔ�T�5�=e�C]o|-����hz�$��9����n��ʧ��nHC�bRy�A���HK���G�Lg۴��TY�@��s	�lY�*M5�	��w^�ᾞ(Q��ܢ4v�f��������
h)iq���$F�O�2�X�xCh�e��2`�@�5�K�4r�t�in��{v9)�ӯа,4\*�Z��T:M�01���
�i�\񓵺����c��.��P��]�I@4�$.��s�]w����͡�H+/8���N��q��WU徭D^/n:[�Sή!k���[�M� �ݨ�f*h*�ւ��b�P�5�D�nՠ����eS@��<�u1�Ȋ	1&O �af{rf^3��@'A�Wm{G�8Y�:��0>^퍬��s�f.��~�Ck��dx/��8�W���p�
~O�a���W<�k��f�R{� +J�;�>4{���,u*X�4��Mk��ul���##��#y��=.��K�? ����;�F�Iy1�������v��>%�<�J�ŮG�7�T����%-����~n�Z� �Z^�c؈��!ܚ��dUv^�4(���Bb�&̆8t�X��`�0�@�.��^*�Jhc%lu)�\�!���F�4�%]{8���k�k'[�m	�=I����	򎟵/}�"%�f4b�-{2�/�-~��Y6�X�2�4�7���ޛ&�C%��ik#/���Ǩ�jC61X�R\^m���l�'�_�G�{+���4���Ƨ=��ow��a��ٰg��{�P��>X�85��9���7��ܻa���~U=&X;�G��l)l�)���W�4�9�Lm�[�J��I�\ls�z����f�s���:������Ѓ�-e��c�E�?ݠ��*F�nb����iֽH�:kJ�l_�ΗRF�����}/%��yQ�7��N-��CO+�X:١�Z�Ɨ�NV��(�s���RΑ����,4@�	�@�k�ᏁO)��Ĉ`�����&�ȓ � �+������ [c�6�蜉Q�'֝]���ځ�Ċ0=�����ec�<�
���yPs����W���yE�A�dMΠ��`8�� }��ǰD�.�d�n-���Z�;��ᒔ��v�K'?�-��ch�jBϑ���e|K�^�M�c���tBs,�~S+;dPF�#�1�hG����K�N&��s���J�ys:��G:��I�x�@n� ȒY	O�-�B�U��5��n�м����A'x!d��`èk�W@2^%��h�v��l��r̃i�f��@��P|��aڔ�C�>�r�	NB^h��DM��ݡ�?u'D6(~2A��7�����H�6�^Z�X�
oy�6�L�> ��]*�Q]ꯊ%��"��f	!���G|��ёC%!Ʌ��$`��q��+�������3-0v����������?�L��c �l:�eN�jf�l��T�^����<��3�U�����o�P�	�_N���K�/aJiۀ���.�C�V�vƷ$=l�=�!k��TV��aCƈ7�������Se�'y
֋�������ݵ�f���C�ݪ��[?��>��[ǵ9*��N~h�X0��ҧ�go���=f��]x"�x%\t��,N��a E����~<3%��n�O��ݕ��dݧ��Q2ߚ�E�锇����i��Xz6A ��B֨�@���v�IO#��Z^��J��;��5�4xZY�u$�v�b���>��-�	���:�@�gc�to������$V6�GM��Z�Sc��p���J������i����="�����S���9[�d����o-'�)��&5{3�M'���k ω��^���Z#�4��ᓅ%����}el�._��tK�f�9K��������.���w_}u~�����g�^��B��R��郟O׮�e��o���㎚���A�'v?C�L��N��V�h!�������X�L{��k0����i�� �ۢ	P�#h����9���@C�=��b��~�}b�Ё��6�#�}�,l<����#�t�B1M��s�(�qL�E���]U%n
���wq�xNp�&��p��*Vl�CvA�&g��2�Wµ��lh#�kK�V����9�n���� �����Ȇ�%dJ�UD�����.�࿜ˡ��"�j�:t�-��� T�GSE�Fz�%�Bs��^��%1jË���SJ������Y7ѷw*}:��5����F%wb�Es߿�9p�HbJj�t����հ��|���s����i�����Y��UR9�S�Tj��Ecug��.P�|�3˳�s�c�
��-�&9�
��0VP� :"��,�ݼu�Dc�X��Zϩ؂e}r]v�РG�����$�[�N}�QQB���(�WחYm6z~�ޝ���č|�?@=�#+��e棈Z�7�D�ȉ#4Q���=L�VL`��ڜ8VPT���3q�	�B����9(n�z�B9o��O7a��Co����)�	i��4��kp�׹7�ܦy<v�d&��?6����������^�'���ƛΏ۵�i
���춻˚y)�:��P�c���3;��t�u��y��#9R�f�W|�"�:`Ҕd'�u�0���5�j���	��=�.Ӛ��ϧ�ۡ���"�O_�&�`��d�Km�fl�pJ��
 �#�4��}�Ay��h>Ӈ�!�I�'ήmE�����ڪ�j�V@'�5Az��I���Nx��2D�� [Q�4�I�����NR}�R*�(]]�����aد�T@/�=v6N�f �J��k]=|�����[;.+����"쮢:Y8���/ǹa���
���֧�k��0�	*,����K��$E���&�Z%�n�7�@v����ҩcOG(�Lx
E|J~$=������P�FB������kV�Q`�>S�ǁ�����t5CjGF�ܑaI�t�����YV�TF�0Gj3G�Ŕ[����X�em�I����i<n�e���J/�ނ�����8�j�w7���hl�_t8�1����hXJ0[�l���*>�-��00Vƚ�8�By��y�CA��hD2h�:1��c���\�5i�=5�ъ�ߚՁ]S��I�Z�=b�
jx�<�"���D֪d���)="+���瘉1����&�]��fK^±2cR�Łȸ��W?^7/!�h8o�}%�yLf}i6~�Y\�m��i�� Q3B�&��I��B����>C��B $
�<�1���v$��Ue�A0�Y5'G!U��فn�����{	��@��o>Lh�%+ːO�Տ��<}�G� �]%�7��X�7����ؙ.X��+@͘���k�-Y�1�כM|~љ�1���p4���:�Z<��c4d[w���Gت��M0U�����Mm�l�t�X>�����ݬ��A!��c<��sY���(�]�ژ�}��1�);�CZ�hC�_H���,�������� ��0�'1\wjR�a�y[X���d�����Rs����������Ws�J�/�j��~�]f��;� E2���<���2i��*����~m��,����'����k6��d4mkq��Ϋe\}��r���^�~�c�a�1c����P+�S��nS[N��r�a��)q_P��t���_����d�!��6`��?9TXu#��^~qR�c��)�D,1���B��|���>r�5�bol�5�`�)��w���Q�0�̓=�/��u2�txuI�x��޾b��E�#N���'A&o�[/�m
ӯ\	S�������[b,��@�D�*c0l��m�ED~�v(?���[���gn��)u;'�N-�LQF"�D-f;�%�]Q�'-S�`GDv��~@!��*5�o�2�Q�����{2TBi�wX����T
�,��"��:C�}� q��\�͒�ت���5�Qy�hU*X���S���*�%߱$�ŴUI͟B./��\��7 +�o�®�y��nu� �Έ�Dd#%��<H�*���c3%�H�6B��J-E �ùqʽ����#e#�q�B�K׳�Ņ%����5��ݗ�H��j���Ї$�.q�ua��@�7�Y�f.naz2�x1�)����>Z-��h�Z�.�*�X��I�w�;A��Xu��q�=Yї�N5mz��7In|�4���ҪD��*vh{S��L����dOU4�)�"cj����v�A�`�iCV����Ƚ--�����K��*7�/����D�'B�(�ikkl��	��3�	O\��]v]�s��������C���x�~�$Q>������/_l�\��H�9����W,�M�K�l���O�%���Q
�.�|��t���7���L! v[{���ZC>� ��{m�w��<�<�Y�7\��� B�Tӣ-��oD��_F<�[�\D����4�"�1�=��ᑸ��r��ҝt�r�������]윌zW����q�}��K�`��Sq�`f����y���(�Y��*D���YF%��K�[������� <~UD�xP����Թ�"s�����7,Rpە�"�r������+�"c�Q����T���cő29`�n07��3�'�w��bW�-��Ӣ��ڐ�I�`)L��u7R�K���ӫ�*j@��~�_ C�PH�^No��E~�H�ڔ]{�s�	S]p}xyT*Bu��*�9�ު{f-��>K�?��򯄆�~�S��U��m�Cԫ��(腔�..���Ţ߳{�T{O��_9��ŹǓ���Sƶ������d<����s�$'q%Bw�)G�Q��qg�*��Z��+�� B��H̻���S�����̐�[h���m��m^y��c�;gNF�T;iMn�g��6�Z�� !q�K��)��Qu�
 ��?���
��\�խ�7�1R$�2�8Jի����M�A�֊f�^9�^��Z�1�4�9/����(YF?O���g�^t�k����~����@�]����>!m���q�x�K�Ւ�ˋ�Cf:�����h��m�'�Ⱥ�r�=tj��#$��&�%�=Q��� �դ�hN0\�%˅�C�b2X�z9���g�4y�/pW��cejF�L�P-J�� �ε"\�u�"��':��^��D�58��33̍�e��J9��D6���x�Y���nCK/>�7Q==�pV\����
�����l���W9��[�P�����j�\��G�ѐ[�^��\��m3�3+G��\y/���NI�ٶƼڎ�*��!��~M�)���,��}��f�]s T���h�U̾Ay�@�8j6�í�0}6R�Ņ���0s|��^���e���:�]J��|~Â��������1��v��C�t헤qdU��4#Fi*��Vq�����q�QZV5�逃�$���a�G��}8����.�N3�Φ��C��"�k����c�ݰ$<�U�_�ƽSHg�	P���a̵�A�����g���ui�Ԝ��m�7��a�R��M|�H�� ��F�̜��P����s@Bf��U�XAnYS8�������y��:��3��:Chsa�e��{Az��P�#`IN!l�����.� ��&l��V���*7�hA���d������]sy�s";"~���9*�,�0��d�
��Ax�O@OLeha��AQ?e�gE���9A��Y��+��v�>�y$�'P7Ei�2���;������#2+�;}�`�lH�+ZI0�
�ҙ��*�_�>[P\PGzb~���,��}ӹ��0)q<����˙Ή0;B��;\	g�{�t^C\�(0�Y�\.��Zi�&��/����׺��&�ԿN�Q�wCS>�]��u´����?_Ȏ����A?@�m
�z}&�{?�x�=�46�0^C|�5K��v�N�$<��`�m`-^�@Q�����bͤ4n���aٔñ���t����
�����^#�<�b�	���0�<\����Zo�O����JzY�KҸLpYt�)�$���	2r�"��y��k��O�(bvN�F�M���3D���t���U(�� �rK�5Ul��L[��\׈H��Ț	3PQ�[�6�N����!@ޛ�l�>���ۛaćG��Q��	(%�/�cR?�7p�7�?��@�W��%���]�@' �@$�m{V��6ю��:�,�3�����;q=�c@��ǈ�1��l���9W4����������`z�����bQ�v���5�Nx��?1@IT2hyQ�=�i��j�n3��i��V�pk{p�l�E�?����e!Gg��W �ѧ��a�tR��+V����)�<�S�ZߖF�.bއ�87������,$��"}+�ܥCĦ�S"�:RcU7��C=4Tm�����l.�T}�G;�y�����w4yKӶ�0JAn��)~9���ѡ�įM�s�S���y��λ��Ĺ���{j�˴;��J�����X5_�-��s}m;%G:�������Z�D`�:��]"���Is���Tdv�O��ϧ/�������3Ӄ�S�L8�=yx����3pg�ktsY��e�	w`/,F�����rla�KVl�@{w����x>����YK}a�w�@*:�h�$z��Jh�*Ƨ3&�L�&kz�K�ET5�+��Unʶ�Wީ��������~ٔ��Ta�o�@'b?�!������J�����p�&�?�I�Oh��`��Z
S��^��E�z9��Mk���ʍ
��2J�V�!H�e.�����cz��(��3���	4o��ɘ>%R�e�]�G�y~��R?���Jɾgt
����	���Y�a���j�T��8���A����"�����:�oF@�����Y��a����E�]��=� `5>Wq��dzh޵�A'�����*3ѡ��h���tZ�#��P�qB�eŃ(���.����Ю� ��>�)����Sn�Y 7�U�Y�k,n*}สe��g��U1$#w��B��/(q��"��5ƽ���/w�Q�.���6�_L�6(�����q�ٮ����A��{��-*ۊ������0ʽ����\h��'>s����
p1&�O� �zi�����q���.�Cެ�v���'ĺÊ	���y��i����ΐՆ���ͪ�Q=�&�P��`J����a����Q�DS�̩5�3?��m��d
�7�R\�����J��;�0�n�5��*��AԀi#��{�-�UmFۮ��W~��p�7�v��uCp&X�сqTK����Վ��7���0TZ(+�2�2����-�}4i��9���1d2j����x�N�U�R`ވR���:��W����)��BH~��T�7;BI�5P��6�d ��4�fl"���Q^c����S��:R\I��ԅ���]6M�Ί��X^��G�.�C���o�j�����õ�W$��C�`I�`i&�;������@�]B9 �8M��S'���1�fwg�'�\>C���A�n�S1u3s��+�Vz̓��e�Q{�3� b�
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zWxa9U67ZC0+Fi9yE04gxZTs8+o8VyiLA6C89V7yOfmd2ncC1abDBmtyx7Hw/rJ7gCfasl0GLskq
2m7hqXMNms6pbfL1imXVdIQsuLQscma/ohgIg9uLlw0NlvxinQhOcy+2jru+a4LKGECDM8dc5VrG
LD3V/xVv+aPakdWykgvZP0vOH6rG65h4uFfSZVE11fzbUzoPZWiOP7jiH63y427gyllOMeZMjv/3
j/ajJOCWcqGfrqt5S05C9pnrtv8nvS5NE+8OPgV70hMHz/TqMEWcR4w4jG+y8HBRGMPN4RArlwBg
uWKsI7dQR2k/tyNCDLEUcBCFiaMgPsj+aD1JcQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8544)
`protect data_block
AcBp71ehkRaL17u0aCiPGFVkv8RHGy8XAJAaJgMTWZoDdDQm7GxVqD2njcXbBWGcFIU9Mnw58Kui
bNBO0Y+8fcu7OaalUXDNoeBkGKPOL0l2zQUaWEJYM/jpavBkl/7wZ8/TgT5ye2lQsnqmuMWgw15g
PhAKHR9HMcrSd8Exb3Ba3iu/89K1dSniYy4LIRuk4JUWZV627HUrdCQTXyZrrT1GCE7BBCvqMqi7
g/aKLGC73BpIn734rSxNNQgHlluhU2eZ5hNP2JVutkwd2gOuVCuwBO1tW/sA0+CB5KBnrynVWZ6B
hdCTy4iR0IaWUXgOuW++olX/RyhfZi6pCELPOQlrOnSfoAvhc7EFLxABU/NMmhHe8c8wfZHt1A27
gBRuiv6NkkFYEV8du/LK+6ggJpdg0JCE06ALkvbBWPMjE4X2IbZUVUt9NZxFMWCp3VNm7ctfY7Dy
dlKKNrntiEN1DF7YlwdKy6u9YEHuiZN87nqjkRO97qx7uVP2xJBreyoj6AxU2toYT7rTJCrTqZg7
dD4lRus78UFTvWGeA9jsA07JSHlEJ+QmtBu5bBxx/euzV6iDFYavHaU35JswFlMLvgR87bh0OLa3
cBI480NxRyqboyyczlNXzBUuPNs5JXigiav4sKO/fj2ZVvVCHRWPwo+XJFfCPNS7FMixjRTmeHcV
ortzdz9qtDki2XmgS8XhaT0InXSnCdFReyqi5G8Yq5fto0++0Z1poAcz2RCBgJd+XGeb/ErXWti2
i4U3PQiPIt+K+gp8hTKbp0uh4Mw2D+mQ7tKI7JyuZkdw2WZO7Q5dfqKOhNtwbe6NBTek3uQBdMsy
TT/OtfHL1Ljxyf8303NlUf6oSo+i4tdxYLLpK6BwIzo/BQ3k4shRSo/XOdekQDpg+riDJwI+EBwv
ymuzyatUGYfSb+HDrtbTlWBuso42DxGHYamPd2GS6JIyqeqRdUvyD3q3NN4bq01GwXSBCpxLe6cN
B55JA6bfPh05IT6iuWA9JcQza9tNyWJr83HlylnsuUOD5GV3+1hIeGaCnX541d05qewhCrBKQSO7
i60NFPapbVUXUgYPgttUTng/xqbqNSXMBRggVubIohbuj8LEryVnJT56boLHZnKxKmZc6tOLlt6j
MuuCu9XEwnbR6muL0H7g1N5Wq5NFZ0IZ8xBfjllwUkQ68m9/BF7ytM8MN75wGBnOU/fjZ9v6NwpI
5fD881ObUnhmKFWZwmYcpxzHvJfjPJfl4h170CDMDnThqunFLDF/GdyoBpT5+7TCwCnE7TB61uGi
fmrru+ht0lkKeh0GcPCQW6CjXpiBogZGg2rzYgsVtYJfksnEkqrZHT4FKhbbVjTv0uGk/zsVGN6E
NPN0kd9IjjMo7ZVrktcwxk6yMqHvC4qK8bCgXBiSzUXT0cHAvyM1qq8agzPT6u/ugz5ij3VU/HpY
VQb+oGwaM/vZjHNu423JPNjc8HHKg4yrftAPTXmUZtWT0wpcwQPLXVSbn3GXFBvZKRkJChg9rJVo
osk60MeuJLBxYGsEH0CBAKph5rVtV0oSs6EA9xHBTFVAW9BKa/loG+EhQY2YU2OVig9nAMIWJzLV
V60a5mWcwADQG473bE2JFyPvCi4EORfaW7RcsQ3is2nRu+O/tC9apB/AY3VLV5U9jP6gDepV7VUV
myS81zkU4ncmX7zHkpQQd1qbVMkavJpKgxsmG1kIcjppMR7rpI8EZFz9J8inFRrCHi1b8ITkIbxE
rThT23g3+1ESR1maqP3foDFSF4cWq+XcBRDk0mF6Z8HX92YXFFb629hZHk5QvrBLjj5esWH8gSwI
6PgPl9cUi2Br6Ll7T5ObldA0rWPdMukelrqQzeofzvzJciYE6eOAba36NEFj4i2CeIq/3Oh4I/le
l4m108h4UawPTqgK0Xw2OJVIQdzhALR/9vyomm3SiQYPh02ibhISaTqytCI31Cj/rA8U9WK4D46x
f7iRxbG1m9Iq8XchKqWAWRCcQsbIkpESu77vNjF505IV+iG6YxkHUH4FFt80SsHRcT+VF5Au4XnW
s2aPHFXC2K11ULhAXsHagxHWKJ05jrjLxvqgRzFJpsb28Ih6PDFXjCAWz2s1sIKeKoiEwakhTQ6n
D8K7Uy6SxQK1M5CdEzl2uNAC0Ma8cMUh3x3XmS7koczHhiMYST6UjOCD+U24GrQcf35WMdFPRh89
48dXfrYkeNIe8HMtz+5X8wqeg4b2xeIHWyBSX/XnG+dx6jowCoUnJXXuoMaMS6F8E+XdMd9imS28
pXL6ZgSgb3fJAWicmHkzHgPU5gtybv/6EEuAQullUFw2AVORyrSBP4AEARVyoZ2sJuf6CNn4jPYw
Etz64WrmszlFseZciPWF69el2MJTi9NC3qRuqgqXPeUnsR25T1yDX9SH+7N8Ty01Hfwyb+qD6osV
dPk2sThRVrC9E9t6BO+M9vPO/iQLOD+SQvYiNZ3jMBY5VdZcnpDbKU6d91+EPEzt7+BYnhpxF81f
HVHWBrpGvuIb8UOfQbM9IFVxVfEd2oq+YBctOFaPX/ZAHSJGgXSJZ8cfMG0HQgSFpfIciLHY4zSR
4faO0kUh7BYPSpth9zikjU4AmjOKnW0s7D+Wmyn0cNGSdXxYE/ilRnCTo/imK8lV3UWdcuPjSpFt
hBN35BMFmososRT3dd6lHYlsYm2NeKdFeigErS0W3Se5GUQnF3iXxyJm33ztW4y7dS95ZWhQlcRz
LYpTXHxphlcam7yA6FM0nymh1fzMMFk4bNNvcdHqUpUzfY6cLth1KgxLusMzy+3LIK17AH9gl2C6
dYVR/2Gapv6fXoCA2wu7FtWMRyYy3Bm3l3BNc1ezqEsbHdphWVRa9rF5ep5pzg57SBk6uZeJg1iS
COVLibbQa4lADWGIlXa9ao8gZdrMgTw7Ag1U6ak6/1WkfUFJJS5eDh/f1OYDI21KuuRqXmlvACuE
NvxoCSQD14Kee+fO7fNcZvC5h3EorX9e4IGooH+ei41KFXXtXuYRwOb4PhGFROAErxKZ1M5kU7CJ
BLP4fa5dm6jIdS2u1OtiFJjRJ0681+/6yTg1tmka08/DIZv2ivCKiKW4NKE6FZ55aY+xyVUXXhrr
q1bkq30D8MFIVKv50WCCVH7YqRiHMMRiL0FYqGBHvvG4x9S2fZ+ACq8ymb3KrWUDCOR89CW1PSF8
IC3isBpnXrlgVTqYFtGdEOdvxykLw5kzFhGrUdXuecqgBuUj/bdw4/At8g7KwxeyuxvW+JB6sUl8
x4itJcTlJ5EUdCg6SDdVTwk0Y19xdipURaJpiz0ppodNMI9rGpx7Sa7T0y41dkKrSbiuMLTSo+ul
9bhdJkBsuAiVKClQn4jN14j+ssdEZ6ikTZqh1+cqgMSGJPgCjtexN14cvfeY3yVSUtIUIx+ms1cY
LIuiBRKu4U+Ye+3eRO8T4fHru0eZPtmKZoXPVB8UyR4uK7qQtNQXZ6+Np5j5SDoE0l395mroqjCY
f9FtvNuYqkJYWQpAdNLWEK4J6OG6mScdUmBkoG9+6JLQTnQ24hnw17b84FZ3TbnJYV8z8NHj/KPh
1aLIpaouuQyPVForn/upGSvO7T8PfCAN/Go77qYFtUFw0qVatjUYXDLfrLTrhXCxeoospvzW+Vle
pOO8GG9Ym5YaonYuY6SoLbyir+tFUxKnf/wJd35ZYxuwpZrMs9qakqM1S2adROgqBhmSl2dXj/0+
7tcIMWPNxBe30NNmK+WcjXSWzNM8y/GrQ4TiYZCCrSxjgSUYb4P5myVmMH39RPnWd9lxpKE91r6M
Wd7P8pBFd0gNebJdgUTvVomu3RuHfG40hkZhS4gYdxcaTzqy9GdoSWn6xnlqKI7YtGVSgnTq3TQL
GtyzN6oYjVJVG0oiBJu8owszdn1c9hBGnCeQkhD4I2xF2BHtqLmgcvrURHQnrHcwJhCrR8/os819
TxxOvf1B+LwcrcCq35M98rKw5C3AxDN81OtKgfOvhcTzuib2pdOm/cg0K0sGwYKx5TdPdxrfK/BE
0SmPqllgMS6Di4VeXwSxLhetJ0S27/SEpBTYE0drMELP4KPu7pEtvYASCL/gaklAHQOUUoJezCjB
8B7J41VA1uO5HUk6hczCNzCr+UOQuCVD6NI9YglgYlk0ViIbF2kHyGcQp4mf1zx5OYqGNnhPzkpC
Zj0HpDjvzlfkRN8mT7XM+xmIerfAnWyUSmH9H8z/WMQdHINvGk5Fl4ZUAMGtSZjeA8meDyU6iakx
HopFQMFoIMg4xkSN56Z0nEN0UV2IkKF3wL8AeihlFDjD7IwzyoUoQEUdG5cHQxIHDPOIaBYquyoU
+q+fHbYbGg0X0CUEdl6CDyJ7uGy3/2ZlVbdzxNaEYQnzV62Rne10+aOQB4rmkYonCqhGK9lwVFl1
NqXMyuIgcJ9Wl3guEUXVBNjyr2b7A+qBm7WHPApBNMsmD7XNCHk8PARsN4B9LziXfrfxWkvu+Lfm
8Kd4otA0+ZthrU7we+QBFRchtpW6yQIqJ1A+qZE0d88ff7iQec5ACajpmEGed0rsw1wlWhaCB7Ej
TzkEKVc66EyIJKghKzKS7dxU3kzsk76JQEsIoiwyC7VdKLLGAXpaPyohDMvja7KdB4h/+eeWdo2U
Y1ImDD971lC2i2xynVPR8n4YIKGGtuKCGS2em3V7Pht/mHP7MLtgWOky0EJhz3pvtqpuIu2XqUAs
RDhkT7RBvjzQkfKHbDtYoBotF3Gy8S4tdYh1EeGWJI6g1sOAa/FUksL57qpM5rYqeTSEoaIMA4c3
Fjk50FpUC95qX3/IBYouBF8muXrA0JqsNdaFUcsOJgY9QAnDroG1JnPs7+a9Fj5xVTfSfZ0nuAYs
/QIeDJHO155PYETNTVuFWHxUp1w45nSX9QVKWdbZFVx5GZc1jssnDNZ6Vy/rL0N9XFlHXHtgYIij
RIbUl9a9CzV/xy8HCK+GrAFf4GpdJUVGNg0Vflep9y9rFFFElFJyCtSsbKs3c+q2lx5FyY8+TPwO
GfKXAZCzoJ+nO5aRHx/ZxZ+PVNzRynfcXY+Azv2CU+3JZaF3YiIucYCf+jK23CnomDrs70sUuPH4
ww0+E63RyHrdj1Qt68PCLuoZ7mOuwgar1ufupTi3onAgW2QWN7w5SETbG2W6dqVFXCSMl5yEnb1X
bLOeJw3twu4zy1WJl3IM9ugo0xy0DlsE+9/MnQzkfnYV9MKo1CfIM8eIeW05LZrwFVAwApJI0fKo
0d9I0D6vX1WyDuc5US46QlUPB1Fwbx7GR4zfHSk0zvwkfEDB2ZTCfmbR54mfYGT3tu4B9DXV95UH
NtyE6woYFBXrTR+71iqhu7MA9MpanApxY6kF2kC9IgZy2p1hO6T+/c4SpernL6fDg+K17S/l4IIE
BzeQDJmVB7R8t5aPLtgZKnceKeZBo3hd5CZljsA7KzNiC1evhdLI03wKZs4x01FYZQM0YW47vsBn
KGMnLWiLQUZlNe5AQU00pkRk41l7hOaU2NxXB+GxSyRmkFgbHoyPVITYekC4x47LR7FMb+fmnie6
kTa5c4WY89iX4qA/q2uJU2tznBrKjHG6IuF+pvPukJrkRlGqFghyRKtXC79WP36zNSGKRdf3gop1
sBXNWicuoEwgRw+5aTv2lHurylgqbhlHm/C1RTKcP8cBoAoZk4Rms1tdbTaaO/arLAZf9mgCj2fV
7acxUfpwxN6RFHDS4D69ZLjOIys9kimNXlx0fXRxLlSSivfsqyY9/V8blLgeJt2qwp1SQlVZmgdY
ZQqKiLsbntfofgaP8ECuPZuSuS8MHu5hGyCzlyxmSCGVliDfLOAbMvYvSmO7oBLDhu1PjyZfZDks
F5CGIbqcRuwy9JxVKwsNg7vrsZMEHBLTj+9bKa9xSzvUsvr6iiGMtP8LCnl57A2UpNSRRgj1bKC/
Zl8jd/Wq8cLQuB3D0KViasRIDGJlXUZBi8IhOwL0X2vUdyybsGDqFn0j9mFlKMa1nwuaAWN0OZXR
z7FrdH8Xzx1EjIl+aXATnf0gVkz6VLv9cdaZMw4+QPUNdV2H9zyVBaN4MpB2qbEi1e1vqpIRfDzr
+wTboiNqWUERaAy/yCWA4jBBvg/n0Tn/KxT4Tni9BNk/7LBDOQC/zyhuKS5h0Zqzp6rE7XlQXxuL
2nrw1p2Zp1JoVEofgBdQ9XtsiLU5gA/j89OyGQfsao7AerQAk5wLbWflHkWej56TYytQgX8Et2HD
IIEUkHdcsYpllpq5QMnFosbo8RYfiBPql6fDFtPYUSeDTQFDUaBUQQIZRVdUfDTLQz8qikoUG4pg
D/A1OXPXXxwe3mq3BdyQK2+Eoh95xAqExjtne4qfgg79LyCt5DhTk8JOO9j+ssoX7dEkHlKkOH6j
6FlbvTw/BbbhKOVngzDVCfdt510N3d5UKY7DjFK0sjkPD1LgwCuuicsH4ART2wVZt45Y5I0TcOEA
YF1dJ2WpKAzmBBDfTT01Vjtg7vfEzXOlN5kZ3B9/NPteHV8lms11t3hRO11C4HwyjK7Nc+tHdUCL
+IUlvikdqQ9x80iMpzSIbC7jyIXHEHS/bNqUzerzUJoVa8dvvM44WuBd7Wii/izVGxBTVO+PBf5T
rQMWXGkSyg5CBNtTvoI1It0VroU6VJE0GRwRz5I8319zB+vPl/JcsspRY8IWot9YEYxRjfW3BX3M
e15UiPEb5k91qYReaN7Ekd/r2nnwY8eiWehEP3mfm8mlDRLHe10zLQtKGnVBcS5z3px+ThzYOztD
JKhYnO1nHoHDuRjhOLo7deQmO3AOoZpezv1FH3drNoPrJ4JxsXXFIOWHgzZiVb0wLb6tMWTbaorM
S464PltFGqtt2pC1WEoRc99LpXyzjCwFqsrf7iKGwz5P6opBooBGcZOJpVxi6bKhpqKZWniaRHDo
7OtCiXias268sw6kZLzOGYkDZdlQblEAZTeFhFEgGxC/zzmI4/k50aeXm0wDdCG1Yl0zKUkT7mlu
N3da2ScY05liRvgs68HT5KJEJPzE+vXLRUHsMo+VDtIytnqWqTx6KMxJxyLdYfBSNNB2UZmVPrRf
eW/NdXc8GXT6YC9elDaJBUyoUNkvCJg0MPtJgKliL6LXlSrSwvejHkr8EimqC00DZfBYyPhNKfw7
wnuqXAtb2PWbnro4bAWvnFaWfCGyxhgoN22EO1SQiDQjdq5XJdHn77feVmklaU6eRgizTe89K2/A
U3Vd4ViYoSMXq9yGxQP9wBoQN/+wHzt9whL0RCixol7B5NfYN9ledJDBjrWCcfLSz4Oxmg1cTnEc
UubMF7Q6ZFXkeeZg5daRipJunH3dVdM7u990lxkByQ7rAOxvAKRAIcOuWaF24ozBngbM9yoi7zrU
90EXyDi67IWxlHgeFsmcxY2wYNYZCFPUE6MzFwnyjnOuwp6xrA0IoMPQm3eLdFyaNjqH27+pY1OL
tElV7XkAodJG0w+LH0IO282JN3YwLYaGqafqf2dgdusFZrEr/xDiTZDiull2wq5YCh02ckpxK9o0
ghiVkgEgMGhnWdcS4bW9lbb9jIqIQxuPVIQPYIFdbtZI4NQtL2dEEB6aLmVZunbMt7pcztfnnpSe
wnthWpXHF34oEZXq7iPN0pJq4sSizZ5D6vbehA0llA9tzK6DRkq9Xqz5nKp/aIrWxtC+3Uy9EE/L
i/EcvAWfzAnC7ki1yjs8HtLhTnTJ/8lGnoq244nrc/r/tvStDqKHGxP8cVXCTsuJXf9WHoNZr/9C
+LqSeg8ei7r1LF3L8NVDTPYCcP4N8E/d/eWrQEfBLLBgig70HUW+CV5LDQRVp7P2VAswBj5u4Spm
aq0P5Ifd2iqEqaKvNra9eJ5iBUddMtKoVLl2kDgoEZDc8A6uhDnU7GScWXOB+xEMz7FaTFiB9Gdt
xDuLkZnBrINtzp2LdJ7vmqrvwc7sNAGPz31I/xzeRTwxaf8BlzHD5Rpk3Ve3Z0lHVVqwEHiAyyUN
WMkwM6m5iOPWQFB9QSYh0OhDcPPgbarfB3nIwzDHcvhYKrMOuGZzy31FhkDuudqtZHKR93l8NJx0
L8xxOwfk+ze64nJrYN2eRinE4iNAJ6riugifg3JPQVsuVwPatOlfxaGgCtlUUz0bIvxpPciuJulu
AhyCrQ/6/TWfU7cnNLtsaZmYYs8VSl2UdppBPrP4Asm2ANVbjc6uLb5L+i97LaMVs0AQQhwWnVcM
BrpkV5aA9Hq7Hhfyv1qnE/d+IhhFzc+8FCConKY2Cbl7ml2WRRTI4VqSi0kE57jy2uIlNopkv/xm
C+Y6JG7vGKUoz1/KdiEYBC0ky5y2oIjBJlaLY9zKcvEX3rEJ1xdJuBB2tAtZXlekun5ew1vRuqAC
DzUkR+Kx9PTiTZjXVSL94cNsrBB2EsrIN3WHen6FCzpdyd+eu+gQj4Bz4mDQXd25meqjS91XVsZ7
mJ9uhZqrvJBSKXteLh6y0mBbTVTZFjQrWKzq8gQEHbiyETVDTmdmC8HOkI6kbtt7NSHVb152eRlR
gIOXX79vbzy6NIcBQ2BElA8kY3Zo/EQPRxsiwvenBNnASfjcf2z/uer64oqsr7ktN3aqIU2GO2cT
Ju6mAZi8IYH1pFAmMqzpVaxIteUzFoTDAEaWsxccZE+JtoQ+7msTg1GDK1sBGYb6/o7BRSdoz+29
Id5qZuHnc7LQkUsW+2stTdMAJhAOhVFnfOkIXBJpNe3gk66abXFIQ10T+RbuJG1QNd8L4SKs5/Y1
AhwE8dFTJb5VzE5h3cItZfDoWZONe86Jd0wEm+STIBwrciX5hFeLlzgmNU8B5Elzkc6xO9XH78hx
hGOoXnWC1fJmyHY/dJ1kVq9EoQvfkMbFDo+bQVF2WcL2OBQBlcoTIf6fhrOEVsjzwjeDoKxPt83+
ByW7lzToFTdIQUTagvdzLrLZ3XV8X9mZ8BZx8dEPw7BfSfAozesUOnQY7j6IHWNKMuW+BPbdHH7M
yoWs5dn7A0upm13Bne8DWSkT0q0URxkjUEIM2poEUAUjCWio3VopN6MEeMupHaZXz5k2uy4Cu8iL
FhRNsXa25yQnXuBxz1K7f0rPTYUeBo30QZs9dWlYK7S0utuaY0OCirpWBPQzLoC3083Yd/gYNxgM
o1qcB+zOSmrOWK1iUSmPyi/Pnr1FZrNEexPMZLJPS2gpAYZDSETL9ETW1PglvbzMubAoXxDZiGs1
LVr5Z6McW1vBdvlnSKUK0b8e61MUySc8GQ2vppLb1B2yh1NUhPRbbBRCrDlEOW3l+6XUZeRF8hWg
V6m1JisOCtqWYKk5/hyGk+D9QR2/n4lFsfSHFeVvsCk/TWbRwTADML+CxLH43ZEvVxFhJZpvRgt3
/4JNms7/zSZCUTl6ao5Y8x6kpeozQc2BTayLrxZjJy5TJDyGG5FW0nBu6ZMOkrFQWruG3/X/oxt6
+xNct2vlWcZlxAxxg/tR9zdAR+IY2wjjAgCO4kJaxv6jPtUfLk9AoSVhyqS1LRUltsQrKJThmKOD
yyF2AJVtrNPBqtpPdcCo5GpMkrjGrybfxDcvHKrki2psk/BEMMGlDnAo9aacm3G6JUgi2nWU9/HE
98oCY7QLVSPv9ikZqIniYXB6V/K20d20PWLEfoJ0bR4Bc1Kd2lFOqTTMnuX1JmdYl9DrxGLOtCcG
uMEhGrHZ0NiwlmXFbQzJNoyvsecSB2hRyaG7TOQ2nu5iB/1D2JKmy+1JSFKQy8n11I7YjLSLAbDJ
KYBNvtyAF1R6pR4VdYBSoGecxGwl9uvzV1pH8T7WYacLcp0HThE1U+YsaXNigOObRkBJ5x1AagdG
a01WLlfytjIYn8rw5yvOZa+vKw4PF8oA56Pv/jsLJbWtqL9UwLgl42wMkMcLVcCNRC8QHbNKuomw
UsZXkLVV01dltvQyVzpPo5+hWRLCsBARFVZsXDXB5h6u+ITDvAc+gL9/EAsPpjchooz3MzQT4OiV
VPVGsfKjr7sUMKnCDQmHxb1idlN1jUitjWj+0mLrIjcseeYQ+tLQJwcorJLQrJMuv4Z3lzw/Vsju
NoBvi+D+I55DjUvthmgg7j4gR2OhXGUvtBWyPiSAE6EPmdfPSnIvWUCE1gXd/xECHy408fx7JyUa
vN3OxDIGNRy7B24aLhMZszdpoS85SZ3hsaeVTJd1NHH0FPGFHgFv477E7UyjAuHVcyP2hmAz0NIm
iBz8RBbFl/QpQtkC0TXQ9SdfdaExQuFbWZa3jiT7mazP4rSkWmkTpI9KhilsSehviykeo28FE68B
7geZNN8qgSmkjRieREXN3yMr2T7QaxExUhdZpKv/YlF5FMh6X3pAuZn0+4/HsQOVchtY/h+IrQZN
b2nEcXhEM9oINS4HYdS/FUkvC1xCgD8Gq9742gaBqdahNK0Cubji6620g3d8NRukwttbTeNeRDGw
GUw+0e2KeAHmvi6YGVNLXw1s7Cq77dmxEIVkncrqmjPvpvND7Rco9beg0lfqmn1NrUJlnOGC4o2M
+tygM1BJmcySdPigHDYVZBqafJLyAuYxvdfpau7PqnXHyR1n8pDKJ6Aciy6dPXUt4W81lFUXo97x
rBczwXepfuALFHC7ZanACTN5Z8mEe56PJHlI5u1VCWGg+FhVzugSeUckJ5257sIqpyXFzzy/4IpL
+M6o9FlzedZE+CT83aGFxQqCtnWlM2R6sbQPLVzy/U12/sKNp0Ybf6V10r0sLUfSYcZoXJV4D4Sy
OAr+T1d9UpfOL85YkqQmBJEZDpDji3BLsZeSxaWXYxsvs0zQf1TCBR/2qay+GaL1UIkB6go/Qykh
saMCWaDh6Z97oXbxCY3bFK24s4sx+ntNeQ3t4RiihUPu+Y21Tl6FUniNXV2cyRm1IdqHblOZ/UxA
k1hWsbbRNV0JSGH5+YUTymBmkT3WrUsEf/ps2V6iguJO2ib1kgog3LIWaMji/9xfa0w804h031PL
1k33kpvr6ckOvMBPVhMTakgL26ra0NQ8wUDllKOEW9zh+51LlGOB0nbUvy1LMxewbFkd8gcPFsHl
VjiWSegZ4/MaNbCtxJjt/gtx+AGCPc9Uc9QInP5mDoDsU40fSO3XK8kT7L+1dOodB6Qq3rCTnVyn
VrLyzi3BOnrjvK0H7TkEh7Oknqb8HUM8mJFyeIEpFs6YxVn0wxx2u/0XPgh5+WDJE6D90jQFhgiL
dbHq3BNmUHRcznlcBlnmX5s/E3EgH0O01TNf4SR144F9YqWUsPcQM7RDx2yC4wsRvUclpnoIuqog
nK/xpO0elT5Jc5IkTP2uobrvjyIwk5bPOeLDsUVf/Yui2G/peJcNx+xukh0I4dPIvvQ39CFx+fhZ
jrLSBh65nT1j+U7WXgjzMPUTrvHtWWgTPHjOpuqfT33arxsK/vQkN3SisalLqilAeoFv
`protect end_protected

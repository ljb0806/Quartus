-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nrLrSL8ikpS5lmSLjN0uuo+nn+Cc1od3YJ6SXa1uCA7bhFcJP5b+4XC4xHbehnbhzZZ8THD3Vwu3
Ow2pl8/uIh7vRIr6nK7T5UtxXwy1Wz0PzLSD4Qci5R0alJOyiSMYKbTTuHfL4Cn8AjmV9QkDgb4M
2ZH8F7ayROnEoAMR2mFzlT/jcN4yimwr22W6W4qubj5xtV3wStBYH4h/Bd8Wq9Mx/1CyeSXjElKS
RIcQO9bnMV0iT21JH4ff1EOQklq4lGwjurdzLDITnkNwxGoc6IcPp0ywhVWt4vv3eoHu2/2phsqb
xLTmd5jqerLFVJOYd/uDmwyYgZtcWbf/GRPMcQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
emglKQC1qHqOA02CRyxjU41n+B37NXn293bt6EnrLbbQsKSa2dH2RMoopbBEiiPIUhQsVlqLD/0x
ijz7vHMNSQMBzYZpZ22RzV/ByJ52r6bdfJ6W50cc85l9+QdO+bbg0H3OjeKKZNWWjGm4+C9kKeSl
pdTw0eL3otxiNXPx871ApfauJ8qegAKeGCNPRLH5fwwdgVzeVk8js9cGwuHOmSDHGXt0fkPTx6vS
OuHiBUCDprPfEYnfK787gWO5Oa4+WcpzTWEEZKmQKkwWMriNt+1ubWUg8PGrKfCKe7ouUR8V+8jl
CpzJ13kl1jpHcMWirINcF+TuaRWCGxj+6ZujPGT52O9A2icOKVO3vZ1rgBbfgioMnwPx7BNExD9N
Up1oKtitRE1Xgt4tNoAOaf6ANV59y5Wn7CFC8kHgFQB2053k+f0raOu+AzPJFW5JHO7ytDIHVtfv
1fQ5EvoEBz7f1uk7+s7xxClEkx/28eddYPQfP88G1P3c3PZqeEG3/eNqyjrcdhqd5+pHF6r6CMVP
ZD2yNqDcO/5GJj+mIx+trO3tVXYROjKW9EIPEiMVZOlcDK2Lw9BBBwOpC22sYZbyoXuBmNrOTxOh
4R42bidDF8CS75fwV0fhaHQ0S1NF1Iu6Ko4p1pf32F0la2IqoJqgu5MkePShrUrH7odWhY0QEtOi
8WmaBjJI/9SQQyRmkkUcefvcuH+94XUHgvFV52KmwYbYdHi5jSqT0g+Gymez2qT6Nt+MejuS5XhM
LR3i+YJizOV6U3Nr67Rr43Z+CiM4o77D1SMjKxK242WF/nDoBn0GlpIhcVYyeUwKBzNHraqSeY+K
YRz5FgV0CagIgl4jSA8OATcRgu7qQTysv4Dt3ZZHTmABPHLd8328vfiD19wCBxedz8+P2iGY4yJ6
OLDFfA5hQI/qGeqwfs3gEdCoo5ySr0J3yKfE7keiP8Rwv0HZvHXylbm8CBdV075bj8ddG3iPnj5g
+mRkqR6YFt6IhiOE2sEU5PIp8sYwerHA3PDb/uVJUEjvbHvGNyj4G2xRjA2+gKE2Cv+K5myjyxNX
HHoUmRIcpqrvS5LGG+5kZHQAcumN0dcHOF1tdIqIYaSaWivSLWsTvsqAwCiv4Bctqug+qkcNdAmF
DvSjpIkAE5zLuVLX/7iKDh9boz2nUMikF5Pt6R6+nXQwyaTtt2xdy4h/8qHZxthfKR71lRG0yG61
eCJtZRGBRMhbKcpdIHaApgv+eoHFi/qeVGo6K53y1E9fkLZyBl0aECklIrpChyOBH7grx9qpkGBf
22W7DMSue1MA8cDzrQvp3uhd2dknvjf+FzlVcvfheUlBxAnBKyXToK9+xf59uyq/2SCH83XFqPt0
y+5T4i7fztcl4QS5mA64Bph4mxbfqlckm8fQ5MMHIHt5JxkQNwrIvKY90bf6qcfkeNBIfB1pMHhr
6BtdAaTdPkBDzjBiTZeqXsPgEF4Z/Wp6EI6XugkMw/e5NPiC7q+/cD9/B7IlIDThZIW3nL+CtHlU
YLtpuJNqk3gzODd+H8xEU6FtRetzn5K0UxjQg5qz1EMX1XBzane/gycFaJbSUUJBLs0UkAyrnq0a
rv7YO6a40XDCF18zpwQjmD5hI+BtrieqK7HOrh1HmjLGKtBezpX4MbY/Eid0xQMuDGV1VspVmSxF
VqmlEmq6F8diwwmykZ0rZODB/hU7ro1nDqE2Yz33so/t+M881aC4aIroQcncEbdLCIM5HzL6K50S
LpfH7NNpKjhu8Ca7EWN7ThdRawcntA2JspR/xIxAdnUg3KI46KhRrYITT/1+FOegqPMfyGKYDqTM
iA6319HcG/fwW5BU3yoJx1NNKM1bFUQyynxhgvxacrdS1fzQU4NLOktOqFsvL7gSBmOpchK2qiDf
bzYKsQhcXUBJ6V5D+JYZoyvF+QKuOTp2kBpEa8+PRslf7xoAe4FLglwcwR2AD5kp9HADiy+YRUkv
rdoM9IAvbhnbxbhv82ijGQdkBJ4xh3bNKaOCort5/kMvnFfgkuV1JXgRd24i+xIl5ZPzjXHQM5Q3
gL+cdIMAvLbm+nJUbyPvz98pDoUvIg4iy6teTZ06zWRjN7rxExwPlHBceX5DpKmU8ZFJsU4cvJbI
ARA0+SS63N57ilKurbuqSSrkbUVtLLS+9ictYiBuxVE7dgCmI0hEHg90/DNxk3f+VAos0Ed6RGw1
EJQQ3ppUR5zYeqK8f5WihRg2bV34QHn5ZEAvDJuA/sMvRtocv3cjDm0u46e9JQMc7HRSVeJTHq90
pACUkzZld+k8kOaIBAIjrxb3BNJPhNXB9L+kpttFzDW+AYIwlQcyeYw39fnvkQPY0/O0R2mo5+HZ
I0WXxwzBiSeXfJTvi6rn708uRfBBRz7z/EwRG7tWLTOzqBbnrm5HK4QGXzBi/TS/Y8qK9rVgzHLP
zTM2xGzs1zwHqymM3eCGYyxlWZVS6P60vK7HPSpycLRt/NTeFeKizcKLyWrN1+RCMTqeApzy/mmg
WwPE/8O6dUw3fK6iWUkVchVD/z7xYbU4hBV6/SZbkPN4fbG36hVftk4uDljtLpJhv8GZ/BlZFNPA
Oz6vMZulnJFj7TRSX5VJ8/3FSuQkxymvTQ/YZS/MxvhJ5kTCySqRTRPZgMW8ItJsYV9Wl08Vvs3y
GUx/W04ks8hJ5v62mAec0trKxsBdIkE5B9DB7UwdO2irV6wUXXcy0Ii1yzBDAUxlIq/i6ZS6K/WB
cAGVKWvptq4TvY+HVd2ytwuGcNykhT3Me/XJeF/Ho47jtJc2oxLh5xLGb+7tMx0fS13Nltg9Z7mh
sMba5KT8iCmT7rY7yRGcXPYv7SpycW8mxhJn7sQa5HvDNpV+q2YByOMPjDQnrNhyJeu/7OJA5ezI
ZUB/YdiKmwYRVG2DeQwAV1t9LuMR7nTVo0vxKvmK8FHhUeV6XRM/IMdH2GueL1FEfyFymuVS3FBB
moX/K38KoweAxWQTAUD47qVse62AHwUt8J9iWiPu3RSspNazyTulm6D48XPcptKYlxC4ZYq6owLm
iG2wYzUVicUaB1mx0xJk9ifunu5EwHhA/fHr0V6sidPd4VKDoFI1uq4sEOWMW4V+sYqLMqCeocec
5lTiTkJwEOsQkFB8ufdlC5C2e+4QcJSwxG1yVlV/DRoqmI77cvWKJzChZlHh5AMlQy+Mk57VvEFc
iSos9DUq8cdN7btUP/6Rok0zaSJPa3JZ4ptdRj9vuZUfbZ2nBg6OhLbdPsluYAw3S4F0o+ugQ/VP
Xm4Un7zYI4CjgkjUwSTgKNM8kfoD5tCmgIgt0o5ynAO1/d8d52za4SvRxmYz9pSem5dE4W2IBlDQ
6UNUoNyvXJx2kh7eo844HASQ1O8WoDyM67KpBOzQ4ujDt7q6qIcRyrhflz/GhNiLWXZHluT4xY9Z
ldt9YDv6NfN6XYVj7TbC1nCGlV1VwwZM2+yGtuC7GnUPGYsW3+0tdLe70cTb0YQwtSDDtGpYzmIy
pqbA0P5y02YZnq4u0JrYZDJI4G/4WlGwEdaMABNMDn/pXswVMyPw7/cxWCIIvZ/Tempnt0R7lyOS
L3VnHvq/YEJWsEe+zqnt3nRehgDszoekiQGXTFQd9eAVX9dBMAV4QOzWxmShDp+g/txe67CHCiSs
hd/L+YP4uFVUS0L6htINeYzG5vz8P+Zd26hu67QjH4J2/YD1mx4czrcP3qZF9Swa2NmEXSAJqslt
Ln3R/mEbsdHH6dZfa5QDWwF6GFJDbc5jJ5W0E1llSjU573EnQb4E36u6aRoKtvDig16wO2YNCiIQ
qU4xusdcfVcOl0UneWBEAhe2N60w8zYpi78BYyO23nq7bzcSeXnPVSfVTHr6/HSvtcbmghsi2oaw
OhE1G1Dv2aECDXLHO83cm46y5e/LUm8JQbRr6mTOQ7e9vJDw2i4FpEkIXtQQZ8/z3evWwx/9F9pe
9s17gLCVfcwi2cwka1DIFxbKCn0AVSPq2YaWbCsEBecq13Q0vvJU9rpqDEiYlZAdNlc3DCljHinC
J/pK9sgRtn6T6v7+iBowItxZArmMvgkQoh5TphisEDzhbn+Yo31gzzh+qOFomAjZTyYKG9oftXCU
MeTNZL8D/J+ENanZviwXIPCB65d2+NT3az5fLK05RHSiv2N602D/96MjfezTgtcsxICq7AIzvPfw
vN2TXwmkXVevkjD75MUoHBoWeH6+yhfLTOCftlE/e0N/gEVsViyNpnEP9ikTUAh6NSy4VDL0JjNT
Rw0KiT0mOZuJ4y/8p8Q5rR4Yfh0Gz5yY6MQ27Qm7mFwlo4HrkOU+a/VCL240l5gULqBGEtRoVGKc
O5Um21+aWAeBtnirbE0hS1mTqELmIcZSUNv9Np8sDtCxoncAUr9Xv1S5AaHmlP9WR+6zlJp3I36e
7XOoZoe3PAJ+nl+yLxHxDCavNtgPn4iVSEHYNBOK+7upyqCdhqcBmetDLywyGZLm/UjujX27RsnE
6LmYngN/En8z9GvrBiR/h0kfdzaRWwqs5ZW+5EU1asQcpojA7YgMTDT2J4En7fza9KZDLmWJ2r7L
0dnUgp1nkP5NEH+X1kHzlPAX8NbudVqm2KlU3CdXcVKaybLXn/Zz95FJQl2DQqHm0CKy5GE8SKmY
c0XVsVDj8MV2H7rbBzPWXIUS/BDm1BtJ/xeoIh8Yjr60SThExWs13ywONbYiMu2hiNFWARdJcZoW
MGuJu+N4ZNKY3QPr6zZb0OuRRmjYu4Hz/ZUmx1es/GtquAww0dFKkMASGYIbccCPEsv9JPI7qCJx
DoI5LFLont3stlBFFCVIkk1IrrGzHYUlT/8l1Qn9XaRKJIiOLRSIVzVkND/u343TdakSNPZJcHKA
O1UeLwV3H1ArcSIpdBdrD+AKwB3+1pjUKDufOZ9HGWuJNENucJVt4JMxber1TKxSNJPiMsf8K7Z+
vOaBdDvo3SqADuVUH2zpTzePjdvLFNH5ckrK9L9C84dal2qK4DwsMx7um6GE2VPE3kpPsJNiylkS
UHyPla1/fiTnZehwExdOMoXCxOy9D92PhnFS4rW15vqW8i1LklAnJDKitUC3TgvKEfxbPQhq8lmb
inn46o4UgzYLgGLFGdiCCyETXiPOcRsY0l9JrbbrLA2V7x0XMMW6vMM8GAO6cPe4NuUzW+KTouUZ
Z5GgOCrE2iwaQ115X3A+vpsDLyQ8YuB6akyVFSn132wdl5x8QUuXeoj1F7ASpMtcyfGc55FS/Kx1
jpTXwwne9AqcMGlBKcZOJZiQwGve65aIoHgUqB8AvSiDQx3IOElQBeDvv9IB9n/brJHI3rhI5njU
7hgdDs9/qZHSaAVRziJKjpVFyBu4x9LrhsE7SyVY/LhSPexiFddnBHibNicxmxZspKy7KQjM4L0c
vZU4Li3gRLEwFg10l0gOPLfnd4hzL4FedfHEztXVsRaSJuFZGX6rdFmVCpYvWWfZtbVF4OsDpMSm
TCCyHtCEB20pCRqOLqRBws/jE7KB9qigDUiRSsyjKE0WFTTiUay5tSblvqA4wRIgjeckL4sf/Z49
85n1Qn4+LYVHViv/QQ4l54RAitw4BxZnLdGr3+Sn4VWAn0318XxqDWm79AhQfm24XKegLMdHIcu3
RGxpjG8S9YRjsH9hpQT8mHMw4uX4Nd/5rcpZHM3nnllKQZDgNH/JnmPp4ro0ggYxyet6Ig6mFbJu
TUHXMW//+Ghm4qFH6WfosV6PpWknyPhHEl7xl3NREeTt/o9LIXIHsckIelffBSGbMqOld47+VGVM
n+6YRkVm1aFQO0lbDQdWEvJS92IAOYm1aEoNVkN55x5dbf2pNyS1kDCD7i1Q4Yqc5LQD0YUH+gDQ
RukBH/AG/pvhN+T3vu0wCD/w6BsuyxxIk3Tx2aLyU617J6J9CZ+r5y3T6aTsnwne4o+gLGIjq5re
iOL86hMZ65OseIiRZO1PTFZmrq28jyUXkbsy8f/yDeOly4FMXayD+JMGRluY2PlPB2CdlnLog9OX
tBlBpMgo4FBiYsCDAvankMv8exV7OTujdAJElBNjUaVoVp1ReWK4FvVdcxPJVMejr9vRDfoZ3C9x
scczLF1YuhtEgYS/hILsgE0Lmb46U2AjtuLkLwjLe/Rrdwv9FekCeQSdLB96G8P42PJNsT7vf4t0
jJYfwk4NCc8P2wGsvl2H2qpKLjzEuuVgVsmkMbHgZxarpCtKh7ljGIxLwTouPXWoidZRtUmyjMLs
5dBnR8HlmwKU3k3AEacBahQqvqz4UW/qb7kAvmI1iVc3hD1J55xReLFOb4FHhxDt791G2TRh+ovg
o9w1gUKrNqxH65HUTw0rxnD3Ab8hN6VWL3y7TqCrjZVZy9X4nl7VwShSdyRYnGaBNJWPyjQPb6sM
a/FK13AZqSGpAOmThfsGAQXLu4KBCFz6rQ8n1J6Y0/txIfMWOFnThjKKw5rs51mLr18mKEpzNTs8
0RLDwMpeAMb+lsZeOFo5NIvzazrEZKBfH/Pd76OqBB9ym6DrPj1jUbrFnO0Pw0iCz9l1UmlQsrLi
2KzyVmEaMWM0CkrjwFF3kqI4Gm3nAKHya9kTTFfz85siRoRRqLyZhAXGM7szyaXKeENiRgJO+6GF
BPqyffyryfRDjjDtmkTqylBBpHj35RRWvu3lFD354bqrIRdh+5HKNWWGRTFNWozNgTG3bb5Vs53y
A2rfOOTG/QqWNPCItqDPgiDafv+5fWACNyQkX5+NXTzXuqRnhyyzcFkl2KSYR1Acu8MNwq7BEo1X
2ZEoIT9BvF+DmHVoTvneGKrvBV8g82rXK2D9CINlr2pLhPbmKGWfw18nqQpBPrTFCVjjtD+2EhQ4
xQLyJedABauat6sGuoiiID5KTQcp5BnPZNKzLdZx5wxYtqAhIR1CVe0lSvS/+MH2KY4XlkVt/5Eu
/tIvWw5Pu7Zdz4prDFOSf3QrYrcHnT0p9EMTz4PRjjBV5x01i/zC6udgjr8uJ7M4N7TKscPSHAX1
i9GuDZ/IM23EMYi3Nd5nYvVely8dXrG5+dRALLH8tWQoJ399g0NtOzImF4jt+XbtBnoIDZh2Bdch
t0UlInMWRYOP4FWHyzH2C2jNCVO5RizppaZHKkBESpOwOmvw29wviJFXvyBRaldvYVdz2uhZcZ1u
noThopbzw4MXIFKfy/9VANH2iA3sf8e4NA0B5iJg4GCS1pJr48s6u4RXKnDdcjqUQZoARSsH4qT/
nlXtqveUxZIOPEGWAYNtvddLF4StDqwfXh5UE0nYv6kBmgWb9OPQ3OQtOl9KkgIFeBm/i8LMYkGZ
KcHGU7QXtGH5H+Qz+8mvYZPW6xysC1IV0TyKpmEZMeMDNuSaDBCTqqixSdJUi7LiJ8Oi5BoKPhyi
bRjqwM/Mr7ohBCFN2d0t7dZrcIBvnqL17jFSAwnMIbcgMHKQerYC5C8WcxUxGA8NowOhgf1m9S/1
a+RIzhiiQh7DjeDu0b1Ol1cXZ99z2ZQm+RgQKPfSOTljbQ9yrulcUe4qNyJz9WgGGjKomLDhz8Nt
fppYf2VR+p48J2luSq0l23dYowrDcbETGzI5qh3JUqJsb4rPH2X8QM+pRZNq/JH18xu6nQMMYeKk
IOxTBNeWzqHKJQR5Z+0eZTw/Bzkj7Wy5DAoHEzEe2ybv2K1v2lVQ2gmSCVS0fJfG8CSl+9Zf7vvk
/Xr8i9mlVBadh68I6ca6b4YDE5BcdXOjBvnOarfQ15HjXPVfNcuvzSOMMpJXTcTWlxcLUtteRyy+
R4QsjgIHlvubbVi2WTF9B3DjR+pmfWBQFPF1dE0rdwV0b6VvASbQsslVywjqGqfgeXCisSUFbSyI
yMOacHAI+A5fJCraKO3+qX35WKyAKCG7EvQ292h5R1yoR6yhRLLicpsbJ8yBs6Q1J5Wl2C/QhEnw
lQmm1Y8QAaaFd3L3wCsEFwipFHPmW+I1woyoERK7Wwjg5uvustMNz9D1gxvwUXdrscaoelDjfL6P
8Y6iloykajMNfQT7HW6o39W/gi+db9H95fTHxAUixIIB0QNTmpM3eN7Ws4JFVzxwCocbYS0d7pYb
c2dVIz8Bbymcnhz9pgI5mWcKnG9ddansbB+uugR0qUKpfz0QUJWULtXsAKmIUfJ777rIVk3n8vKM
H91sIWqNSYL+0z23mevqZZsAnZ77tWs3gwUoZPykVXQUcm4L+gXj0OE+Qt/h3YfZhTyW7pHqXXnR
JGeHKrcZ9RG9/xHg5tUCM7DIEBOH77uL/N+RQaT79ZAGoMudurU2b9rR/J54z/AK2lNYQqOtvTLL
8VZpQBE+R+dxAJ6BuYQNGk5dNOsCtFgxEGmPILocFXHYUvl4xmSNekd6l/X0PvmK6fKCNgQyI9RC
3L0JP5mXQ+tJyrI4EgPO4DipGHG64eg23Olz3m0YM96c0Xcdo9MxuBZo3JGe/phVcZ0ffBFGrnER
22BdWRXq+Sezqc8F5Htbr4DjxaIk4CjoBA/qQTrmkItXTscnoBhlNkmdlnQq+DatzUWmSZpwcz3t
K3MHpms10IH/kFlIkRkrepBeKMNkB4+4rmKdhXEah75Vdlu1ytEs8OgEZ8MwLtXbd/1kAp26KJ5K
NWX6bogg7ekye2KpPW18ulJYL0y1hOlCicooeGi96BdJl3hqSafLSFdpO0XXcVumbudibn59LgWh
PnNh18B2xKBAcV/yfZUhqxAeIO+hYg4Md/X9RhkKhiramIhkkwiihiPH1Jjx2H8NrvKTreK/Au0/
TUdUL4p+zvQkqJzmaZmHIYWva+IcNAVLN8BSBYwpqlHXtyOH2fmMA3S0yvwtYv6mizXNRkn+gIjw
LHP+Z9br/FegMnvCNGuAqU5fzHWDtaoknThZLA3xjZ/3ug3xt6ANz6KF75w2lWdQcYRP3AuQdZMg
sKZPL5uewJzMja/J1GPxT/MM36BCw5dxYR5COW5mHfminwUQ4B7B/ZRZFFJti2xCJchePnCeuL5J
UB+05X7F9D0Jf0TnfykE39NKVIWEIodKs5t35mzn3aSHFtatFCiUCuk1rdHmyQ6X3kz58scmdqf4
TyJYUb21uaalYFoaika9jZB9xt/CEVh2hs8eaVEyErfhlKfrsk4IAI4I3KheA98pgaV8RjZXFj2a
np0iG4Rq8b8FdMbV3z6ESmAFL/iBPP6/IRfvLxwdAa1ixz86xTjKwI0qsbKEK4mep6gBL85dW5S1
3NT/Q6xxbZIfFrZxkrueLt8qraYnEXgsrDlI5+Xsj28bZw+Gy79r4Au/w3/H1QNPSu5NXYlDHgUz
KWAaBHAh0PNkYCJ7+j6lt7Se2nwMIsMEiAHx3e6EzOldfp1dKbqF0U+yreMv9B6dO+Gk6mW6heOE
4aoJiknMerZtkkMHtEMY1DUPQ8F28/ehj/ecBePwCgZmB7mF2SUCSMLDD+cCc+u3GaN1LDwhDICP
ancir4iPUWDKUbRRiW5Om0Vv8YCm8v5tj0CDDMuQgWWjNMsoXtlkUsX4ylxtDtqopgS/3bi8Yo44
NzQgBKSFebrivRm5oZ+sVKBxZPWuUxpmdSarbPwpnh3R8g63iXieCsUD4A40rNdE2GyR7pqZy5rj
wmzMsB0knm/L+3izVsxPGghOfth0o5QGdLqSZsqQuExvpScpNq2C6M43PzVYFGH5daLC4pXcxXGR
F836pTKPpqBVu/UMdAaY9bmNgN6qrRzhJ72MgbshLT6TktaPAEnoJm2tUl8DVwtwVKa8Q0xbBXmc
CNM4faX6S20PtabfZbIXk4+juwl4THqHq3adRsIzO6bPSCuIv/Ac56EzcSySvqdj2W6H5C1djoDF
aJf/gOx98eD1jogIfT28Qyd4oEnOGJizcggK4y7Q4S5y5DquXIjYDE1BwwLQKogzRZZ7hkEdp/Gi
9M7IYlmYZ7SQD+CPjM6Gf/ltSWvXySN0YdMcgzQmBo+noORkdPaTjcw99lJ69uHbVASFjbALGFwL
dTgxvEqyPhdZ6O90AW147Hn6qpfjLl834/eUdBGCnOiuQblRg9nNz/4Ng9oQj2kfBnH+qiLGxaF9
ZQdN3dex/y99aBvLbjWRDrXAtUnamWExl3DTf48pcQy9L+OWV+ZZ4ysCiAw5+wCLflKHGjPoIOih
LkC1ur7X9DTAPs6OsPqZJmGlCdt0wwXEGvOpSu2pPWNjJmgzSArbykD3OZ/CEYpbC58GtWFxBh4f
9yF+4mRkOE0Q8AFwayXTGvPAuDeTMwxIGJ2mI5J99ql1TU+5jFW+SPrrj/EK0iVRek5BQShOnQo4
orEVKUcDdTWc/rhX0SqHRiI=
`protect end_protected

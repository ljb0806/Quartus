��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��?:Q�s�Z��@��6�W�����@u����Өn��z�'��Ǖ��"�ݗ^v&�N�����X���g�gހO"ۋ�X��Ϲ�㳏x��0�	����d�H)rpK���(��pg�5�Gf��i���+��>��{q�,�K�6s�46/�>���p���7�Tۻj_���ʒp��I�(�sQ���o��Q�&���Rd�k�DTꮸ��t��N\# Z|��Ӻ�ȈQ�QC���
���1_��Rۏ���j������kWB+�Ɨ@�^o�*���O�Um�V�4wS�����`�/�˂G���̊d��m^�bP07�s�grx�s*�2=&EZ�m�{��W4�!9[,o�x܂Ua�`�.���?�@C�����ӳ������jG���$R�L�I�Ե�Z��
��6��a�8F�͜ �CR\�:Fú�Y�	O�D���(:��X卿�H\��G��5Ǻ�u�%{~��h4�����۱��]pܮ���f��V�"�_�8�o�
����*��j,��K��F.Fj�s�1�?�,��$"_M6�&9�2�@/�ra�<O'0���E��:�$I���M�������@S��ָQ�L�Pe����o�����D�r��x}�y��'[j�J"P�ɸ���"�xꊧv�Q��3|9���A9���4>�ש�ʂ|��|�����04wR�
�#�	j�J�
�j�Q��U���L[���珵�a��1�c [�{ڣP��V:�\�B𬬝�MN��SkC��ߖ�;h�p,�<�,T����Zxi�5V�M>���߂P�*�x�H�!ݤ�a�Հ�ai93�Mo>�qӧ�x�FC2�MWSE�h�}v����TQ�}0�}�ٷS��Ɍ�KH�{����n;0�
�Q�e6$�Xm�~#��<)��-A�j�%(<굗�����OV�K��֠ �?�>1$���EI^t�)m�\�nk���/m��|;ZC�-WB�y��El��DI�$�Qɣΰk{0��#�G��FJT�\˓r�}�+�G
��(�{ը�`��X�x�����A|���N	�L���(��ߧ��c�7�ە
d��W�y��H�A9_5�+S��7��{���ԋ�w��j2���GH�.�hl�����sxʖf����D�$�s�!T�pd:�Y�\�"�0-�|	�A�֩ sxtÕ����I�)�-�|.JqI�X#�"�-���XV�����o<4ͨ�����-j7����Ƞ��$˩����p�gf�䵪-�\m��k�yu�#���k�t ����$�n��Ů'`<���@�G�h	'i�(ߵ`�k]�xȡ(БD�0���0Lo����.�������`Q��+{S �J��Hy|(�4�m�����T��jd�u䴌����]�r�"���T/�'~N��A{K��ӯ5�ROu��)j��n�0T�RM���̾�>�s�2�O��be!�[�0����eޅ%�԰�2O����
�d�s���oƊh}��f�'r�@�Z�e�io��ԭ�O�U!�t��?Aeػ�y%@�����R01���j�@��m���qܹ�ʲ�hWwxc"d�
04{4���V��v���+Q�2��-��r���
�5 ����-�?U6����o�MŔ��8�9&W����)z7����b!�dt'^��(�_^ʒ![�wj�1�����<w�Q�k�Pxr�S`��軖hz>44X��39��LF��Ł��<�:$|������@>d;׊l�G��TN���q�AU
u��M3�r������Ѹ��o�t�)mHr�[�s@��B��=@n���Ԅ��$ǰ6Sm�(�ig��B9�x�!��5y�a�%'��3�W��Oq�{��s�V2�ҡ�%��5I��^O������I��Y�n�!s����C��A���@�$���8�\W6B��s�����lZ�sJF���F��h�S&�amS�h�����I��d��}�:E���`���ae7�#Sf\�д���8^⎿J�ȳ8����Ӽ\+�7y�t���R�zK��^���`�� Y<ZY��-uJ�<��,;\2H �~��"9Џ`�:��`��T
�������; �G�7���r���=C#:��]Ԯvj����63a�@��O�*P���۝���19N�C½Jw��1R�V/�P!*%՗JG΋v�?	O�x�� �e��Zp����]���l�r��<�h�%>�iK�%I�ӿ�mE�=���Jz����%}s}o�U�F����V�0���X�)�ϥ
���@!��<;�e�M<�p�V;2dǏ����[� ���V�hX��I��#%�d[!@�W�ܖ�"�"�i��_:�XCe��\��s/'�B͎x ��*��A�lb}�m6�����e�ߵ�H�o�A�i$)vQ���P�;�`���`�$̪�&�d�M��99B?�y�������ki�@�5�_�������%�h�|�SkZ>W���Oͼ�*�*�V��O��w�?(�B��7
�o��P��׫�=��M�{$h��r��y���Tɜ'�c�Wql���	`��7����M� ��~if{&I�a~%[	��2�4	���`V�[���VJ]��h�d�]xĨ�'�X��z$�f���:G�Gac���T���c%���``T(� �B8��r?J��,�����rP�`"��A�1rwNy#��ac��v�.�[��3�z/����3����_�+������@��s"7V��zc,��'F�-�=oB�h�DS��@6�όك��7�YH��Щ��@�?��k,�+�B��cы4��B���@�S8�JO����/k�2�����:��1rB�>啱~d�/��o��0�C0J�K���;ȣ�Eͯ%8���opҩ!�:��Ј*#f��!| VGrDIw9��y}��/��-����n�.��L땛܈3�3��UC����@�b�I�(�p! �E����f����� `>D��c���9���ͅ�<��r����>��ݱ����r�j:��H�A�V���Ɗ#��8C)2@Os�
ښ�N��[�K�}s�?�r��:Ep�wq.G��=�?�G� �ڶ�K��y=#���;��ܛyf�t��H��2�����Ȣ��������.yo��7�P)�e�[���4��g<vى��OU�-��:d����u]~�ev�y6�̈́[�.)������i��J�
�&��H��.��&�R�1H0�_�^s9�f���T��M�
eB�:5���돟����\7��8����W�
��?�o���x1#��Cu�kG�_��(3�6��*�Y��X�;u�2��H�R�^7�p;��h3ʿB����`�R�W�X�����Љ�p���.oPQ�	ku�Z�% w/Ƴ��	�D�:�D�^-?T�/ܚ�b�J�L�k�E�On��%rqj3� ]M(��� �.��\�d��E٬�����k�U���C�����m�PH�I15�@���o�e��4��H�훐�7j�����uT]�GL}�?�DOC���J����jW��S"Ͼ0J����40�"x'�pa��U+�	�ʮ#���X�R���"F�=4��O[2��=)���ڃ~9�`����!��fү�qF�&��զ�����B]����/!��^C�MqW�7�,�
{��=9�߆ xA����{B��)��-#����x4m���ū��e�N0����]Gq�ʤ�J���@�p���D��m��0���������c��트���G��HZ�1�;��[��6�vm+�f�5�6�o��99�[�p�f$eI�9����~ �h\��+!kM�5�f��x�����(�ry8�<̍NC{�w4�/��Ǔo�K
ruj���(Jԙ�W�H9�b'���rP��Ui�����������&{��\��t�Ý�y��~�,X���cV��+?O�`� ^bm�A�zܩ9~u�a$�k��"�Y���v��>-��������6>B����&��R���0��cyu1���b�w3 f+����_��\eS�_�w�a��s���~����4��L8�mΑ8�zP���ݴ�tP]���<1�a�\-��tܰ��?;��Q3Ȩ0�����1%�}/[o�� ���k�Ȭ|J�5z����N�.-�t��&�9��]�������3�{�����Boԑ�Gd�+4 ��fU������ �x9�o��!�A�<�f]h��T�q�_O_�g! AF�J�\��D�u����Pt�4� ���:�Z2b}<��S$���m�m��H�L��$���+b�zI5	C�2	s�e���iҝ�+ R�����L	�pg�Q�uz���)��?*!��Tc�3���"��
������}�KS�e�.�ƅb�!%U'Hޥ֧[���E��l#��a����	h�B6�#k6*�e<�?L匷��#֬.�z� ����/+R==u���!���1s�:�+�fU��z�L�ƾQ�ᒙ�2�P&����j�����E��"�=Ϫ^����Z�(_�ބ}d۲�Ƕ�:"�Q���YVvF��A <��T38hK�C�!6����i�����r��x��r5��Ȥ�ߐ>����(����N��)
l�Z<��Yr"���0p�606�%�`�kE�wI���y'+�B�:_8�~_.�>���4-�a/eЉX�(_�a�^|/�m���`<_�gx��{"{�B��2���P	|��k������t�{�4��_r��ϳ��l���_a�J��%��j⬧�RKs��4�#�m/8A�pݖc�/Lj��LA���
*)ۄ��m4Z�����`�e�����j+$�:}T���/g�89S�'�{��Jy������+j�k}hI�$n>g�S���-%ʳvD�6	�q��C+��~�c�(��Q�j�&
�")���}�rIx�:�|�0�����I�2��;PB�_^L(�m<����x�A�_���>4�W�eH:}�jUC��.���dZ�Yw֘�ؙ/�-��G�_>���
o
id���z@���!�a�(`ԑr�ȱ�fmb ��Bqkq�%l���H��Q�c�^z�E+���9���"z��R�d޺~�̶�-.�2��r���ҙ��:�˝I�?/�k*��yN����_�4!=���-��T�o�\��!��,��P�:��=�0�~�7c��Oa���.�^)�\.�@� �2~G���Pj��TtW�F�I&g�gA��yQf�&5�z:�NM�a�����d���=N�P&�>g�M>���%��,�|Q�l��_$9�^�6eP3>��H�����7�h�Q	��'�0Sȍ�H�\�"|�F��:j�$��s�	�==Ga��:�U�M��Z�X>C]���U�ը>_.�e�Nzގ�A�jGpm��L����e��7#�1��i��x�VH�:a�}w[��l����_B3�L�4�R����BDv���̥����f�p�p:P��m���֘&��ỉ��8'b%�h�]ѣ"o����dc}��$_���
;�!���e9�o`����-�p5�!�Sq��IY�1rJ#�wc�"�.E�zt�!�X��m���l�V۸�ѥ%���q����J��B���]�~���i�����2>dٻw3�G ����/����u��ŴV�����q�~���:�=������I0V�R�����`�_�`���#��h�x��;�mw2�č�cRSw ^�KF����ً�|�JNY�%�qxFrDk��
}����";2)S)����d0QG��f1�r\d�T���ΪR P��P��!yQ6�����ǲ&;�:rh�5��7r([�saD�~�#�i�cD�ަ�kd�[�K]fއ,vDw�'�t�;��J'�I�z�t$C-a��� ���`7�O-����0�@N�>�H�l�q:�9�����Cߣ�%�Ǽ��d�<�.�\ˏ ��r���{�o��z5@MK6>���"���#n���@���o�ܛ1�:ΜȸGr�I �l�M�U�X��k{�2�)�U@�N4�V��)F����%�sb�J�1Tʷ�b�e;I7��U��|�|��v�n��o�Q$�ŋ#x��k�4�*���K��TBhWs��S�<�^J_6r'xI��c�'ё/���j�SfB9jo������A��V�D"zȄo���A-�j~T^���=l��3��W9P"*ua��0�l�0��XA2����T0��2���~��
v�^��l���e4=*�?�J-�xJ*1_@��# �$���DM�V���\R��0X�7I�7W_�O'������½�8*��\��~cJQ9z���<����2�g�D~���O,$ײU�|T��֫*w
��Jq[��|������{H��S\(�m�m!/�z��xl?���#��"�Hf6_��7&^� ��Ś��`��c�׆����S�X�O!ڥ�c��gH��yy��b4z����Z,UoEu 5_�����&p&��+��9�.�&ItiB�s-�DM��d���#�����&��9��K���)m+x�"�w#�M>�H:\��@�c�Xy.1��lAzg�>�����4�'jЍ��e���x��(m�A�0�A�\��rLV(n��C�=C��x��"��PM�~`۷���5�F�I����:�(���y�$��W���P/u�
�O-�)���X�5�Q�Y��1����^����rq�bf���E�h�/Xo���a/r�r��3
@��L�fm4C��5P��)��ݚj1�{�*a͵�h)�C�h�z�l�;� y�n׼3�Õ%���`�ii��qZ)\��N�OW�@��<-����Jm0��ZS�3n,�Z
so���&[���c��r]�D9#׷J`d���c�,ф�ʘ��hPaO��CQ�,�=����`P.s����m��!R�sRM��u�ߧ5�aPW)-��fQ�#��=��O#��R3�ԗ��>c��(�����[d�Wڇ΁h�v�QgL���#��U�[����Zf��/�m��_^ ��W@Z�y(��V��E��z���IS���K����Q�y�p�U������?��ƛ���r�
@�n���z��r��Ͳ�L
�ZRZK��	ݧ�k��-c �F�C�<j��PdCU��<�>���k����AV����ih�]1F���)�Gy�>��8�0�`�
��w�w�5�8�Z:(�p�S�_��;�7��/C��_t�q���h׷J����/p��oU˶PЊ�쵴`˷iyG0�;��ա<�,A��;���f���y�m<�v��5��F�"�W-b�q��M�Dj����Ʈ8�Xi���e�W��%�Kת�t�������Qp�t�7[��gl���;Yh��8��qWZ�{�n���F�Y��c�)���I����"��a ��x�گ1�LЌtH��Po�p'Ϯ��+�P��8�Ѽc!��u�My�%��zOkR�2���By,�0TJ��\V��^I�hJ}rU��q��Jx���(��.�y�Oy�L7A��z�lϚIZq�!��0�K��cK"��s����4N���3��6Y�;�WM�\�X�$�('�J��*ר�9��|� ]��E\mI>�i���+I����_����ݗ۲��4�l�Pcw�$�f�e�]Ǌ��\E���u���!�b
��~��E�8�M�p��Bd9�
c|�I��I���~�ػ:�acыR��M�M�kf�9^d�n�iBۛ�Ӎ!�O����\N �K�\���P��6�;�_�������k�@2;����y"��xdy)�0����i�D?l%՛�Y��,ɹ.y:<"��C�[��$���_0�q@;�����P,bg�b��Ρ���;k�1��]�ͅE�,�(���� !
8"� ����Y������4
{Wx�q�*�Kԧ���M�����
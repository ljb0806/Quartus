��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB��1��F1܆�p�~�2�"�����S�'γ,/�'�3l�A�Ŧ�{�}�7Ie��T���h��v���2ä��>�"[	p�*]F���Y.5�H�bcm	���>�>��pu�X͡�Ώ(&��Hr��@/W��jje$��o$�k*X;Q��Z��� ��YIƥ� n�96�{�?~��^Q+�ȫ�|�E*)��j#�/I���.C�I��B�n����Sjd����R�x)D��Z���;x��^��0�;F���8J� �p@<�l�4�t���R��h�}��` ��G�m��rwp|��0^G���W�v����p�w�9Z�'��p{���c��~f���"c��r][�z9�8�aH^e�9��K��Y�0\!oڧ�7�1!/��|3*�m��%�oX��Sږ�=�n�ʜ�mޭkT<����J���zj���0`s��$�O7.ܔi#`;�IǢ����䋲FCm���]!�y���tϥ�n����y�k4%�a4-���#���7�o�����֛���K#6�@ch��ɽrgR�+I�HU�	���uc�]�W��j��5֌mƝl>��%�U?� ��[���'m�s�a���d1�^]C��&{8	����c�Gp�h~�uO�����.	6a�^�Jϭ���9� �.�`?����j����⹾�^@�tq�z#2���?$����@X$
7�3�a{�0P��e�J��D׉�]GO
Qc�� U9᎒��|�)��=K�ʣᜣ��g(/��w-�RB�Z/e��:=�/WҌV�Ձk:Cҳ�%w<`x#HׯWO/�������~�x�J��T5�lˁ?p��	�ȁ1@SI�����5��c��|�K���\�8��ʴ/|��R���	aL�Н��2��j#��F�ԑLJ��ar>�`ġ �:׍�i�Z���WL���pKIڥ���[�R𶫾��s��h�6*��\�����W+q�E>���pNo�g7#v�	��;�\��~V�bS98�L.�ꨑ������n�J�Af����6j��'�$��(�L��3{��s���{o�7��j���ѳz�����t��7_�6��;��O6S�z^��9�U�H[�[`j���{K�Kz��Mi`���O0�w��@�Q�^�Z�]��r�a�Ƙ����Ŝ�Fh��N��'lċ�������n��6��Q	1��ә�4�+���!a���a�ޓҭ���g_�h�6��S�4�E�oϖc��m��'d�>��?"�Ӷs:�:��G�&�2��u�13�����e�������?�f1Ic����-��ӹB1P&\�l���G~<d-7��i8E��,����i��Z�M�g=�ͫ��$uN��k�3�˧��m�\0C������e�}�#�90�:K�A�mC�\텡�?�іG)�����!����ި$�n�m���58��S����>��	�FŸ�KU�ՄFX`IێHf�ў��9zߕ�n05�<����n����E��.��.3�R�ܧΏ��@a�ܬE8*Ƈ͸b��H+L�N����z]��w�h��a&�����$�q��T����tO����۟��Q���Vǃv0�k�E8�g�M�F*P"�e[紞�h�$�&p>��1��Z�!l�y��B�ly�������$-���0爯��F�S��8������YB�r�k4�����Q�-�I�����&��*��b��.2��_E��Ѱ�n�}gP����Ɓ>~?@��xk��(l���t��z��tM����03楨���;�F�;�4;zG��I�A' ��!t�l�au�{���<鬟�W�s�|h��˱�����O��"��c���y�[�:9d�+��׮�I�qV�Q;�NR��Z��6%QjT�d�-�Y���iR�PY�M�)�o�?��/����c�� �e�j6.�o4��N���1o�	��.�M�ܳ����XT	�'��4Pr���
"���L?�W���n^�۴	�b.��\�Ѯ?"��'�e#vc7(�\^��s8�f��Jx��G
'8�O�g���2*�Ũt�(B�|����(x�'|Ҡ{+q���,��J�.���B04�V��k�!����ЯĉZ�������3�F/��"%�F|f͐��E
\߶C����Z��5�'��]S����2q�)*����;Pa���h1���.����D\��%q�P�|�
2Ovyjx>w��+4u��`]��R�6�x�Je�q?&.\D�4u&�ˮ�`�7G�	x� 5������G�8�.p�c���	@��3ݪD��N�����L����9�ǦXnw�ޖ���o�.K�
Ŕt��;�?Y�F���� q4�+�QCW�r�	{9�O_P�AFj��Bݳ����{V�d������Z�ĀD��B{��wr�0q��;}�"�<3����\��|�nn5�u�b /�bZ	�A��~���+\�$���ϡ"��{��)��u�N{���0l�� ���:w�əO|f��̉�۶P)0��'?>E��$�ØR�񱽹��n����I��qRՓ������o)[��^�H��ټ5�x�<`�:�~N2?Y�{�[$�6'�l='��<)����'�DNb���WHz���v���gy���ˋ��pL�(����[���B*��l�-�ΒI�1���81b���/��O[膏\� @��/U���6h>��@M���'�ޝ��ȞJ]-r�z߿����ܱ7-�8�a�EPO�2[��dOg��%��R�^�<ި�I�.k/j!Ⱥ��c���E������A��+������c�ӝкQ�s���@M0�Ųψ��2p#1��QwC�_}{���Q��L����iJ}�G:�8�2T�Z��/6��}���f�'Vz�-�H�����=VY��B�]:�3�:�������ѹ�d��SíOθ�a8=<�P����������u;tF�],��[�M_���G�}B^(��5�'��SZ����_��{�?�e Y%�F�l�TW�Te��û+���a]�B���	��J�SS��xՈ��P��F�ʗ�Z���O,*�C0�	W�O绮�_�Җ��D��
Qk]���
v�W	:�w\���p�CE��(Os/�=�L��4��<����G�*��v���n��X�.��n����:��1�g�'\��=�pv��%D>�(���Pc"z7lw�����7	�|J�:Հ{l���e�7�_}+*�&ߚ�.�\�� �T��IA"Ҝ�,x��gO�c��Adbq�s�_3,^�!�����8��
�����{���؃�D�j  |�n#�Q��Ɋ�؋sބ{�(�q�]Ъ�k�$�����ԥ�hV��8�	��AO)�!j��*E���^�S�9���/lgbw��/��u��o>�r�����*�<1�O�G��8��!1��^g��Rf���bs�Me��Ȣ�bŪ@��X���b�����R���6���c��w�sR?\�v�,��p!
��t���ޛ���&<�$fu�f�W���ҷ�v���k�<� X�%
(}��)ހ�C�
�*��M���5�;��6��g� 67���E�vOCU�*��w\ �L@�!�xA��2_2�S]Y��߱=7�>��M0D��P�}��{��jq�v���o���QPi(=�$�!e�o�>MӘ\Eǣ�3�Ӣ�\#�
8��x��&C�� j���r+���������j�C@�͈��ޙ5S�Ayː�`�r�'��:g�8��
W��m�;����l����4.#���0�	��]�q2�m�(To�n�x��V5�K6��ǃ=�1�Woɠ{7G�?C��������t%�Q`��d�������Y��s8Cp%��-fZ�CR����P�T|��|a5���au ���t�/'�Zw�Iw���@x<�Xzb�Ü�q@���;:I��>�.�A'/�ʈ͛M, ���`�$���u1���Q�0��@�QI]�O3�}�:e��8��Ư�����1��z
7t��,���?��	�F�iM!�lf٩Y�~�<{D�"7�������oT�]_�_zu�3Jr�hb�~������r�?GAzT��\�D�_A���j)!'��:��"��^�b�C`S�;C�x�n�#�Yh��㋎F6	"��6�D4���w���F�Һ�b��s�#/&fƫ%ab�G9�z�����8��������i,��yVT�з��M�b*;Cs��Ja�@���ZZB���B?:8h�r����������&HU~����Hb>՛�jc��@�(�좡�@����} T(z!9lqt��m�2�	���:]3���m򘟸��Ȑ����DY��l�~�{>w���]B���1Y�����W.R��Pv��� ��)ծ�(��̔�i>L䔁�"ݩbQw�E�o
&�(� ��2����ռ ����N��l���b��bI���I��Dّ���S����&܏��d�����"~ioZf4�G����Z�$w��I��ԼiV�P�1g#�D]R��H8�{'�?�ym�n�t��q7Q�xN���� !����:�;��>��U;���gX��Uގ��/5v���e�j.(jU��%E*@%��r^��`I��B�,蝮/�`l�3�y#f܂z�����u�����1��yI��=�X���~W��{��xw�G6��|��i)��Îѯ���	���Jqmz> ��*g}�3�47oWW[��M5^�FNQ ��Y�4�'�:->ݩ���X��;"����X�����O�ό6-�P�D�[(ɔ;}8�݀�|��<R�xi+r e��݂&{��G���C�$LW��f��}vJt�wDN�u�7��+Y�� Ȼ���w��q;0L���5���yђ!8ΉW{1ðvܩ/���:�)9!/߉�E,��2x��U~���O&Fةx�Wx������"��*�F¾�ͲH��R]���*�a�h:C�|��X��͵�����So��FJ:P	idM*�ȅ���ѺUⰁ����b\i`����K/N���4���zF�
6�d)ǫ��.���/�Gu��� 9Y�y���=����@����=Y��i/�ҿP�������*Ҋ�%��t Ll\�Ψ��<
UqKz8_�6J��b*OX�?7G|7h����H����J*Ɉ}A�}�>�*�T"�W������*"����r0h�z���ԬJ�?�]��@�}ol�%�޾@�~�ȩ�RgLRg�ZT���9H�"�}���3�Y�"���̧e��6'q�C�&V)�Bu�XdHY�����}�&�	NQ��16�Z�z6gq�`Z[�WAKWJ�t���1�;�A�讵��E����`P�Ȱ�n��[}�ۗ�U=�9Q��%_�7��~�(�鏻�Y�����ٽ$���>d����
22��/C��O��]L����D]W�N���z!H�R���Q����C�X)K˭����K�W��xG��I' 腻��c3�D�����0 �x&e�h�o+�^0J�h�iO�5���-&�Y�Rx���R��`�WN=Z�������Д㓕�E��x^��V$�8����m���?"��01r�ˈ�T~���j�e�o����2�1�4X�{�Բ���%��ɐ-����"6Aih9Sm�~�����Â���p������>���R�S�-���C/5W�N��5y��t���	��ʰ��Hٗ�Q����/�4ri�P�z�|�+)QQ1B�+�}�fĈ�m�X�g�v��0����>Fa/�u�w�<
fZ��I�F��!���,z՛<eZ�<�G5%��J����YӚ|��N�ԫV L��0�ap[F/�^��SN-|2�t��_�W�����#.��(����!���[a%ő�qIA��Y(�����+!�H	�k�l��h�6�7KJ�L���>Z!���+��Q�Nb�v�q��M�A�1\� ���I��J���~z\�_���U�1��#m�Ki����N���S(��b�1-ƚ/�1�Oꄤ(��7�;e�{�4�iM�+��ͤ`�y� dp_j��2�%W8J�ٲF�:��J���6'\��̐�!t�z_��[�eY$m
?O�����&y�[L��Zt�&����ߦ�w�c��E��*]�We5��7�{oavG��2�ٟ�W�.�x]��9ڋW����f�:�T�Z�*3(R�����8�O*�O�:�c\��.���w�,n�ߤ����G��I�xE�A��+Z2��	v�Xz��6�r�
D�BF��|U�4%p����7y�m;+w���ņ�G���yj ������H�h3N!��S??�XBzk��e�_�G�Ap�����b8�Ʈ{~?�y��\mSP��4((�4�\)�ㆰ����4%�D�N 2qir������㷂������; ��UW"�ze�wF�G�Ƚjg�@���^����.�6��q��'�H&��K����j��|Gq��ʬM�XK�%#rB(s/�Fe5�K�Ϙ�P�5[�p�b`�I~�\�5h��mh��$��7���(������U�7�|���h?���Ս�yp�9s����ɋ�D�ƾ#�(�g�����X|@�K��*���f�xߊ���G�[%܌z/�XK�EUG�w�^��37!I�62<���A�ö�p{��V�,��L��t�����mh��{)�A��E�{TK�b���;���uV�\C��Ɏ�s�l5�Ϥ
���ڂ$u�ٴ�^g��2�
���kw�K;�=�R�����k\V�tH��R����
�ΰs�X�Ĉr��em6�ʲl�?Seʔ���m���[�d�N3�~��d6̐W>�~[  ��{�i���U�K�eA��3���m7���8��a�U|	KՓ�Vn��0�� Mu#�+h����'~��d�v2�e�W��7��d�`�F����>S� f1	�e�qן�m�g�lU���I!�Ȏ��� ��4B_Vg ��)�'�<iD�u/��b��ķ��_��Y�/v� �"R������S1�a�a��v0U�9�5UM~����v��<�m����y��z�a�5�Ui�X�]�^E�	MG�giB�Jq��́݊�����5�mL�0b�Es�
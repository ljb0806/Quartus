��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�"G�k�sz���%��U������ƭooY����_�`�#�|ԨvP-�7{�t���|��^�����ˑ`XD�[n�FP4��� �t�x�k� y�>>}�zX��UW@2nP�D�{߫�V|A�32��X��v���MV?�r��r,�-�^�|�߃|r��d5#q�)����$]����5����2�W�/s�s�_�=W��J�����Oַ������������W��`�����6$�H'2�(�sq�W�ǫ?/��)!���C��Yc�����z��Ja���l���(My��v^60��Gq˝f�����V{�X��2kQ�C��v�n�U�l�֋C�#ߑq~�jb�﹤]�4�ɍ
�bj���́��D`V��n�4�Q;SD����u?)� j08�2�7r���aD��B+3BY�lh��~Bd'�O+z���U�õAm�c���c4	g��P���4��(���b���BEٰ�FA�ntrID۶�î�����e�7����w%�z�;(].y��=ͬG� ��^���{���B92���:�1R8�8�N��i�l�ĤNи�ݻ0+�iƿY�V�hp������G܁�|k.��3�Y��p�|޼*��a���V��S��^�\-ˏ��8A\�}A��h"�7K􊦻܏�k0`u��M��G�ҳ� Q��I ����y�a��ۉ�{��M�4��x4aJ��~ ;=")�k���]��_09Lf��`�w܎����5�^S�Nnj���e���������"!9��}>}�=[T�ugN^%¿�6;ѐ��&%�QwO����.\��W��)����A�"Х�L�N�(@ح�/�����P��2��CԖ�=�� �y i.����{�h�|u�@){�C�9ѭ t4��i�ֿ�P��Kv��T�]#�6�(��{z��G�nHVS[
���"W^�\
�hM����l����7��ڲ��Ŏ-u'x��3��o�{�?��ҡ)o�ڤ}�c�U[ڣ�_��kE������n�e.�}B���U~�HQQ~4v�D�έ�b�U
�	xA���Q�� �ShgMM�S��MS�%+@	��K��7�Y�����@i�nR�?�`:���{��7ci�1p$�~U��&J ^.��t��v��5T"�os�z��/����P��i��~:;�a�Yy�5��C>2Ł{���:����u˲��j%�gj���6���0�Ԁ���y�!� S������)�����uv��!�zv�Dc��E����Hwf�M��\�+���y7?��':�oK��Z�S��FW�s��a�6�����%
��!���M�EY�Vg�0�\���X�\{�`�k0]���be��Ae�s�X�GJA"���O��4�7=�Ƴ�"	ڞc��s�{_'u���ޘQ����	���-����Z�I-Ǳ@|�5m�঒s�x"T~�;8j�ƛ�3فeL�!2V[侫��6/�m��W�7�d�W���//7��.(����%�'��Ck��Y��b�x��wb�H����1�wE0����]�zW��R�)�[)��I���Wo��Aݸ,���I?:!�b@�}�s&�m(�������4m.�Fg��g����nV�P�fT�s�"አjϗd�	��kj���4�����C��w�a���C���qb��o��*���W��k���$�ҾĊ�����blD=�-w��5�����*%WUG#���W�(k��m����'77��D�P�,o�x�D\�Y1���8���q]��ş��{_G��25�F��0x�#���̧S�U�ݨU&�+Y&K,Rx
������\���`u�����ʺ֪k7��VD>qR�Uʉ`t7��`=�ee�����g2��]��.�����{\?�1��ka^�����)�5Ѹ��*����F�^��AM �{m�w6��ɪ�,r$��ẳ2���n&�W <��Q!� �ي�k��a�_�J�lgjN�`��{!a���g���g���c������A���k��2�Z\(�]����x���%
�T:N\� #���|�WA���~�J��0MX�R/�CrS�u��xgČ?�k{��J��G��N���~����̘��a������Ƙ+
�U���L��SZ �`�1��t3᎞+�iFM[â��W16&}`I�9��5����~�\0�#����r7�ά���s,��鸞Ku���iY+��XN�E��������5s3�k�J�]���Z�����B����x�@~��$�?p��5P�(��R�cON|���M�d�5y籎'�s�i��"��ۭT4��h�UM7��"��b�-#y��άe<I�4� 7.����˹xVq!aRv��%��PF~z"s�w&`����ڼ�X^�a�A�Ӕ�)\XT��]��?�J�?r&�t?z�c��1�G�:������X��Ѝ�/�[��j�{�>�� �֫Q4�p�~v�7�r�;'x9R/_�@��7�,�R��a����u��YlI3`��l�����%�7aE�
ad�J{W� ��]ީ?�f�q�1�9ZR6.��ؗ@�[]}�am֎�6��{�}��"Q���7�i��?�.�:Bd�N�M�$�.�FO�zS_�ӱF�Z�*#��۟@�w]�g̰~=L=20f��6`�Tۋfw��|2�t�B���Km����L��o�o
g�e�߹~"�g_Y�!���H�ݩվ�Pe�5ׂ��<sL0c����.��^̘E%�v�~ov�OFo`߈�j��\���Dr^��ޙɬ{����_���g���aHS��&	�)�&���W�!�~����XPߔL̷��U��b���q���+�<2���^�W�Ug���4n��#��Do���L������p��uh�i<��`�H�q�
���0�񿤔��&|c��PLCZ�Sl��O�Z�e��޸X����kE��0�/��D��f@|���M��!(�k2O�x �.M���aK�7��Ya[Rd �TYr�ß��P̝�go����o�E�O��4�da�#��� &Z�О�g|��
^6!���)ř��F[֙]���_�	��sh۠XI�K�(>pS��Gՙ����!q�:Q��ZC�����n�����H�@������Q��� ����ZEݐ�t�;Vy-|�[��$��Xk���щq�,�s�0nW�|��%5��L3������ؗ5���ߋ���ٱ�U��>(�˕�����¢�	�a�OV�?�Q�������m��p3Q����5\+ls�I-b$P�۔q��:�Y�W� � ojl�Q�E�~݋�����w^�<�4$n#_hQ���)�Y�.�J�W&�����峝�e�.*����>�W�(�d%���u�խDk�s�Xq]\����8(���{̟u.]��lM*�1��2C"q����g����4:�G�}�!}��Ke2}�����)dm��pQ�ז�����[VѲ��=%�'&�=����sH��yΝ'w�S�02��	⹠#��т���L\S��L�M���O�]�,�F�U���_��և7�p��+��(��^ʗ�!P$6xI��-��j�*�v��;���B�2��-5_�Sk��X��Bv6<Ͱ�C�7��9y,�����fHu��$k���8L�7-;��B��Bh�A�WC��ɝ>��}����XRZ�*Rի���{�v]yJ]����_&�D0��ӊ���h�rg���F�K�����ؑ�n�X`o��(BP�c����;~B�X���7�G3V�ل��������J:��q�����*�'����P�%���?�+F�a�\��g�k?	�@帣ʫH��H
�g�Q$oOz"�lV��X���}�<�ZQV�Б���='�P�%���w��V���;����ء�N�N���������쳸��!ht�L(� U=a�S��I���k��Q���ғ��ME���k/��d�	շyy�e�+�m��A���;��N>�\���}+)���"/��O��?���7[D�oB��K��@/v��$�}�p2ƷeV��b��`�ݻ���&c���u��;t;p	�vZ�.���0�myo��El�C�@����ߤ+���
&S��yˢ�S{�[g�?�,��E��i���p�!Ddzv�/z����2��p'*�0��n��,~.%1F�)/~Pi
�q����)%񋔨D#�\F��[�&t�ehV�u���"">L�����:9�JP�"٨�7+H��z�rl���D���QW'�{V�S;&~h�� F���B 
ڡ1<��n. ܏.E/�	��[5�mZ�����3�|���Ln�,sA����\#��>��׷�R�H�+GW~}~I�p�G�I���:��H�$���}(��ҙֶ��Ѳ =>��A7w@k�2:Pd��<@m�6Fk�����}���s�E;F��d`v}m��K��|O޻_}��/Y�>b�Ɩiw��Gւ�6�+��j� �P��t�"��x����R*�o5��=kV���}��z �7)}�@=É�S�ĥH�M��T�D�:|Nf/
 @��q�-����t�C;�p��*��nk&�3:���E�� ���j�':J��J����7�OL��}�E3�2�[/}@5�5��sa�^���uw�F�=���+K]��T�tv��<6�g��k����[��@U����P�F�Ӽ������"P�;X��4<����L�����r�; Q���&s
�*�O^K�����
��GY��o{+	���9*KZ�+�,���.��C�+h�h/�"����!eRO���;��Oit�� ���
0@(&tn�@wi\GSL�/�1��]hWԴ����»I�i����ڔd�~�ƹ%x
`EL���ش��J]��S��$�m���1�9����Df���ܷ`0vT
}�u7K
6��"fj'm�Y&�e3цų�-�-��S���Y�ݔ�����|��<�\�._Ф̸�p�S�g�?ѡ�(dIN�=�^^b� �OH���!���P��]�+�Z`���Q��gN���S��ı�2aG�f�Vk�h�n��Ĝ�׏.Y2)�:�F��P5�q8���s�*BM��A�x��]�`�^��B)�h�(o��7�݂f4�(n)Lγ ���_7!��R�±v���������(�a{� �K�q���!��{�%�lm-6��F����
tLAJ�90cu�Nr�mŃ��m�i��D�=�Q�V�9�7����m�T�ؠF��=�E����u���9���mI���&���-��w'�c�c����p�z?����_��k�}���r���,�
���߄�}JA�I����_����l���=���OB�PM�!(���QSٚ<�v��^ʭ��[�&&t���%k�g�np)|�]Po
�T�+e.���\�:����|9����ܙ^���!�c.�+��輷���и�z�3�wU]딭LPԥ�����������j��ё��%�.f@�	�V��`u=��"�4_��X�U�1�o�L�4�`�6����=��BOV�1�M2/�2Uv�QE�^�@/.¬)N �ь��bWF��Tm�kg���fٱKU�[I��r�M��v��N,��6�箔e����[*a�D��Zv]�TK���� �ˠ9������/>���������+4wc\��k�|��7q�%����</�a�>�\��׭�ˑA��1�=��f��h��H�5����@��9��)���o��d9���g���Q}��*"���V��U��W�'�E�cQYP5�a/toʣ3�=8��wB��R���i?�N���jN�����=�c�3��f�?�!�������
�d��9�tU]��-�I$�������������{������1z�9dZ�{�M1�\�Q(�|p�# !6d���������;?�������.Z-������m�Ӟ6_�NG%�[q7Ns�
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VBXcsPvZjKbPHMxB4itdizkA39gbfajIY60Vq8ZzTi5ixj1SGKOOF1IMy84GA8IV+GGugcwCKGup
hnZZeNY4N7fGzNfYuOF1emd1mRxRFCC+bRUvtZs0nvol84M9odaNBS050JnDU1knn7YSssk/qxNe
/ncguzmDRk9Gvl0sBmgXYToBK23N4tjrQVV7z2CPsiPuBvaIb1EGwbgLewrF9aI4W7W6kMasYJw5
w3/K9ZXkPApVVzmJGQPS1Nb2aCjZBdyoRvMD+5pkwBE0EpVvrYIT7G0Gb64NKMMtwfepxY7Vgx5Y
rF54ejZbOVwvJ62PyIAcb7hYcCHYpGQTE1v/VA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
do/6844GdHuNToFvaXOrTKpfkeOkZtjPd1S34essmIvn5il/VgDPTKsohwvRdhVVdKo1OSt6HEOm
7TCxzKJO6mRQUmU6Z6ANWQevt/GuC1OhZNjCHru8gmYYz5fRJMI7uSpdBrk8xKZjJdmPWqavqlOO
xUHaepeGGhRC1Th+vyL+bPQ+SYsDKz0Rr+fSmqL3grnbQMmd1ID/E5lBscbKoiltTf/sRe69b+uB
uXyKeEoiIDFOqbQ+4Xt5HEF3dNDgvem5HsZs22Vka2+JvA9WuFWtXZRxkKTwX0dbLT8gSEvg6l8t
7wY8J6XkmRkgb1ED1/StF5oWh7MX9GOPh0/nHRvPck7tEWGjNEDlEZEFhv76uC8GqxPR7qCHJ4FD
mQUaYuZV8sIaezeyO1brcxmmOiuAT39t96EymmYw0WTMorF/y5RrlleBsi0Pg25Q9lPm48+kH2mB
IPO32oWDhc3AJpd/WVK4TcBFF8l8CQMgqPbFkxA4lqdNdfCxqr0duqap6iVmgFtL2LLb+iUbo54o
PzvB7tTv2GL32tncMlrRGdfgjjyQCscN5eAzsTUUZhyPlOxbW8ar7w1zTp1V+MtBm7SQe+xmh5ML
Qob16W048fKLvEe4SLK++7liQ5dQM3L83fDnK5G7dtQVPygTb+QeX5Krl6F5XAxJKY29UpWEcpCJ
tWckcBFxusd+qWhAQprOqIAmu8AV5/x940lTBTrByhjsHP23zVv3b3+2sHTX2Ybv36XaxDKgAx0G
uQPHLn9S586BnU6XO24XOG+7sLck+fF64CAcg5FFLokGLSVKtv4bEWAI/05cCJTjSJ92lcuYoopj
fqsuqciJOfasEN5m7Mu8aCLgU+4f6deatbSX5eudfhzI7dlWGRpQzgm69BNGG3n8sBGbucN7vcmF
H22noSsgiWPxoIbo6on66rh2ct/fL6eiupTaqjyeu84t+KOrQyEHoXLX+O6eOyLQWoH1TfFSzKzn
kZjbB7YfOXHCBf8snKk4w7oWOs/8MppZ7Gf3LL6yp6aGUY1tlS35U35/sRV350eSNeIO9jjc0Xbg
Pq+SDhbw9MD4NYmJRB6jm3cW+piSqJ11S2uhU5o/LIPYLXg4tuxgUXQm982fgytOqR8EpSBoO77N
mqma2Wh1kboyCczNj6A1zWHmnhPKbhC07kva0go7X1y77ATnlNVaNv6vBnOl9S6UWKYOc/Pz8k39
XMxc7E+aeo/uZWW6E46rV3IfirbfWndtGOZuL/+EmHVF974cl4GQoxaYNqMnqKKhMCwbNcSWBKlf
BneLOH1uxqkY4xYYz2I94Mhopio4yBpq+q8JTqFM9I0i2adzLIxD/byWu50nAZCvtiqtJ0JRY8Uo
XYgq7afIrAn/NvFyi9es+tTr//NlupUf2wPHKz7TE5+uhkvNRxLIrlpM5Vdf5tN+rDM+gzi2v95Y
gXjt+0yr3p3cznPcgT5Vs4nnVtSMyVXZ8O/JAonwc7hds68OLjM8cv+2NDuu9sZHlBJgOmt6uoEM
Qan7Rmmp7o+3HbWwMBwY82Ae8cpRJPyZYZzz87ivmOZfbm7+zGeLYl5mI3gRhop3SZjmMwt4I1iF
G45EN7Me+p8b16l31Show8CHhbaUdJHLm6SYFK9MJgGZYMwH4liBkOCXWcAzuwG/AhzZfI4rZdHZ
ltNAWimOW92T2K0jCbdb8/y3Fhf+2vxI2vjwJhozhfZrs3X5anks/H3hwOia9BaLIdLpf1uKkAr2
VXlFnhQYCjBi/iwLpRZ1/1GSY0iDiLvecnxGlcNF1dZsGoMrwjiCvoY11m64snNKehCg8BogHPRJ
5MYjL6bjfi71VspyFjd7ax3Gf7xA7jKrgV9L2wEFKwP7xXl2ajwS+9KNLDhEdxz47zQsjkwPl/ug
zeeudvEUX3DOqVnj63m1/owVOggyKH1TO9dd8zc3v1NgpIt7F9BbOl23whwsLqCllg6K/hwb3lGy
ZO5I1LEfqhlCIaSN6d95rcAerIe1QDouT64TV+miLdPH0uqnYqdwqYguUDAxQnfiK0fyM5Q+UFUp
PvPSjjTgAZ6vzgyHY8dwaXdnWJaUbZPd7p/Afy0vSn9iMIYdrTmY7udx0vU998r1Ez95zEClgtAE
aowcT68lCledU9xMwzilwwOsVxMHgIBBU3f5EJzzbrvG+W29LbN78gWEHcBshqPZJtJJ8t2+7OE+
Xef9bYze/qLsK1w3RCP6cnER9xV3l1aCrmZNJuvwCImO+0NC55UQw6Swqi5E5ewNJQXI4xZCGqme
SZxM+SY0tLN7YdpDlJN0gAVMA/Epop7Gypb9RafxtKSqAEDuAXt/uEkP6ajLrNMV8u3G9TvQDklQ
+XREQrnAX8U2MObXTf0BJyVQaOY8oEFOJj9abPAhIYzb2Rvz1OMbIucZPwV13t/G1XMWcJn5I+1C
ssqKbE17Sem348k1krixj/RaM8jzojQ/GWXJ4v4bfg+EGMTCJxbnOC70MeREw0Q2s/M8YZ4DK7ud
7b5kHW/mDT1yy6MAo7m4S5n4G1z8syjMYiukcqxbMP6dtPkA0UCsvG6hHjVgZ0G5kqsE7efaG85i
g8LOhlIAMGJF6hbP9I5Q2YcoD2e7J6L7kbgnHaBFgYUeKsPmTee3+sW3iUfGune2dx2/+Bee/4qJ
rWWloWmHyo6UhNlEj4D59pj/NqAyu9R5j6TRXhmNUg5vPw8sHTrPLdGgQ+353t/g33JSsHBFsCdo
R4v7XSM8QOp+odOKgPl8775PCV093h+1WiBs9LtZ/GiWrGxSmtWvez4xITd9Hpvm3YXbju9fZj7W
xtdo6Be0nyRrSJRfeC8hVbNlTSt+sYI8alTr7h0eXEXpdWME7RXVH4Wf/itj1QT+0wdZvNQErqRO
aE1ikrlUGd73zLOtrZXu0/8D9qRPoxoGMnP8HW41RSeixNxTaOfbGbyUAW8mEkoATXirR4iBrZwq
fmXKuBwBlWQsLyXjtElz2IW3K/ZLU8DLZ5RNXny7CCIdVY1LBo80Yj43zsNnYBow7aCcpi4qYjvv
aW/EPdCRc1NnNcUir6glHTWDe/uwE4H6dRk3ZgYqkTP7tA+xH1OqgVQ6bW7n1obp0NCtMqsTrhd9
8BOGcnOST0q3PGDG0Xik/4OtS+227ZFzIUydpmRfApQw+xEiDaXQm8KpUDPXFcuF+mzCRm/Fr6ZD
dUnb0xzzRcY5b9a9gCGQLCUk7BsFgRarDGbX0XokzHAMOGEkioJhfpcZNHnZcYj4uXTKo55QdsG2
jbCEt7FUOE54WyP+/ALsdZyvzVpmgAdxSYQG5KL+kD02vZxySwMzzrQ/bfDPKaHbPUZb28uQX9lp
4CXLUGy6S2f75n0rxbroH26mE2w/D6Et2Cddu7Rl/IjqEfIzVoiSRsRgIP693XMjr24KRdWbLTlg
bjmGzNB/7B215VBHUjhSpfMQRreGInwHA++nA2AlDtMLw9hHW17qkUPPVh+KPvUVw0R7773bsr0I
+fWQFf6+TQ5aZp4JOkDKUBmPQJgRlzKqNn8EfSpWrP2Lao0CmQ2lh6ZEynbBD0unTuR+5xnRHkkT
JZlHkEWGt7Xf9wmOdzzTL+gDdzAAoyS2cziTaGwnEKl4BgJ4mshBUU662f0VQPzeKRqUKOLbdIvb
4TKLO8blnwimyLj29MR9h/VbfFWedYIMBFyxawAu5jNN9Cg7/t0ey1ic4EQ7mHzBy7v1xRhB1q2e
uCg4TuvTEnVCyh0Lve6nmFU7UBwMO1PKePxUPwpeFIDZd7qso+9BbFUVlx8/JZwjTxozQ506uBOe
4SXZ+Z6MSaDP9g17E3dDrrgZOpPIUYoEwzoScwXDA6bOHSNeYolS3n8LJMjEdU5gZtSFcQKEpNG2
GboNjaVK4Iy5/B6MvtTCTroknj7yfNygXDtRrEB+mnYgeG+UJ+q0vlxFOi0xCaBKqLEE3YYQ0SuA
L7cIpoUw1dlC92CFq2pxCsay+C7KzctELjJ0dMT3HIXoA1blRO2V7GK7J/sSW/4PwBcY1dG9Wq4V
BZGffh0xdxKtQzreZgzIKSoP6ApO7pN5+iNHPZVlzJT+1ale0uaiLX+cG9IYNJ8rLzmh7SyMgHuO
Kr8dSAS26bzqU2UUlUEqoYKXct4QV/rgwZU600jXCJdf30zbnyi5PhuW43dBDWo37qPFEwv5CdRF
2uU7gYN2kEfQ4aU4g3gkR5he04I4cPDwbThIr/xaev3exAYuxMqdC55iXEBUxh54o4Woh9mtrmZ4
ydh4fpe7l7qIfwAaE4aFnELBaC0qLXHnBQvf8YtHaYcYuc+OULs1llT2QQFy/+7SYDDlXlJEO+ab
m8SDXx2f4bBJS6Kd0+59WHBB0KSgcEECtokksVU0AmXiFN5zn1JFIrZLK+yfxOxJPXCRSdhNtILJ
a/8F3HKPFHMIPwz43KoakDrUHvTJa1zu33QuvzXCxo45KEQ9zPOzZL8KOXkhjEkzh2z3yENLYh6g
MR+F9OavGJor41ZixeUyxF3x9nKRee35LlfEIs65or1dpiaJkpMPr2jMxFcDHtOviPdc1NTznfF9
ktGcTm7jyieBhBzgxDUYX54DpaYFjmaPInNeKToC///aTQ8foIubz0dPkJ66RgmOIu0NSOFXmqYQ
gp5UAeeN3qdhjJ7vx9cLE4CGjcWAw9QboqpxWN5NMekyxvC8gjbWcxbcuJdaKzB+ReEW9gCbuvwo
OFYuEhERKU6CPYlj6oCE59YAJpyoS7f/xoYd858+LqkupbIUoT+Y79sVuVI4oX2hQ5jlejq8eWSg
rY+E+xRlkXC+UE7A9bb1rK0t8fJ2IX41wpK52E3pb4rHoSmxJ/N2RZ5KnqIxXJrQxbgUls37buj7
eEvO2tsD+7XjGttfSqdpOUa7rRBlg4dNjZWSbSfC14KgY6DsZKrBMIqm9USbXFQ6G68u3t6bhs1P
Elu+dHk9Ei/EooINhnQ16v/UjljB6wHi1OEzSePW2Ph9AgAaKuAaLvsINHOTLyTJ9Rnsbrml3lDm
GxINzhdyBA7VnhSwsUGXfRyxlEhLvl6Ra3My8RBXGdJlg0YGd/eXNo6kojsLwZEW4/4dYASQ7Iiz
itCVqEamMl85czvYBCXRuQnZf18K0RQ+F8xCEmeAMkCOREzRqry2YM7xB/EgEku1mktHuQ33tpMy
itRziuq+KCYlD8fZM7HqDToJbi+8wLNnYFapUjQmbYR3nDrRjvVUF9Oia5AX2Qb6DiQlmxCqcMAI
9Hafc9Uu4G6MDDDGJZBSz0aXqd8A5j4OcbQ5wda7EWPYRZvyPW/OntAkx0P3oTLnO6E8xn7q2o8v
AYeMMgRiV3eAnDK3wd39uZL0iHLY7ExrUnrrE0NjpcsaBkzGpg2Pnqjp9oqiq3FF5P/6aUywIZ14
DnL79EhUxooj1u8vy2kyD+b4PHN0W8CkNrCyazEi6lIGsEGmjar3dd8RnDqISgiuLyVfVeniKxmq
6S/y04RQZ2ZOjygSRPzqxAhspapPOeWxZ8XKCWbStNJVilvfhCeDTwiDW+OdKJ2LGv77NGcPf4cJ
KblRP1hCHFCA/nVkldreKb8/hvvS2VOS5cDdG7oVm8hj51ujWPao6hLz6QAwxRR3fELGIifvmUc3
qFNId/7RoIW17hBCY6BE6bioScJpKAqjJcML4EfA03Rgra4O1SAyzmMzvBHrTunz3y+2PLk/h5CB
OBGrxcSD4d/S8aM96b66hguCITx8TLrpzS8oyGoFnr9KI73HnVA8YlMfD0o5UnK/fJDEXxygflTt
ydKhuo01pZUQtUcSYttl2EulrdEjQxKlwEQ7w41TA0ypplwVLJEZ0luJlWiYvcNxe+hxQbMz68OA
DYjNwmlPBCHE473dtBL4JqCLGaR+Xf0GeDjIhttgLyUei+rjkqfy0CR68tJP1GyHvIZzuSp20lOH
MNd26cmHY+4dQQnkoe7USzXv1gx9Pm9e1AqrxQU7SMUXDs5PVuM6wrmt+O7p5Zmyemtc7AF6LW3Y
qNswX3o00SysNYNlu23IKx7enHEcdMe/ujKV0WcUsbCoka0quG+9snSzF/eOBS+tQ+xcN9xXtrTs
RoV4SluLqjun/dbvMkFqLcm+KFTWlkN1fTUXrOM0S+13zGsBxRVG/0Q8mkm5w+geYyVtwU9UZjKc
xIe4ekQQ2slkoIdDtf4fr3DZOjLzqfU8Zz341w/x+02w6pksj8dqF9pH6z/AVXfthLBSL2M5ILZO
S9K8axnn00dMxYIjz5is6aEhTtAtVR8+GTjEqUABKZ44Zw2CIoC+KBBo2ve/QLVEan0wZBsLlW6k
2gV8tGucVj9XkDLv2yPGRXo+V4+T9IbaqDd8TALby4Aar88BS3vPg1bKe1ZEw8eA3z6PEXAxSCHA
ukAQljGXU8gj+MwGH0giCddLKV6hVweRmulv286gC+CpQ8fE7kdrIOiGPaUjTHLRYtAg1TzeinWd
5smT3NbcvWbvuCrMcBHnliBquzTjCgGIwK2U6c5rtwUgXiygS96MbVvGfg2hi4xqmo+XFsSwtX6A
BA3MZ7EX/3fPQLypFSjHr906eU+mUS8+t+dODwI9jKxzcJXtKOHnXn5VTlXaHQoV2ua1LS4gAhHe
XWc9FyYs9w2NuSDx+eO1/InKSra7sLWT6HMXdi6cTP8xfthmKh+EuaQ6d8+4YdxogAGnuUwujtHz
nTu8f6myaaQz83fYGxQnSgwNKlqpSw5Kx/7IIbHg3vOkVpPH9mdGUnQFVsL5K2NJZEhS5fdohvX5
QBoyjX8tYDomB3StVW9cVNDO//S+clb5HsDqQbiBhTL+HdbWsERtVwxqmreXqKyf9JkU0TLPsGJp
9gKJasQ70KG8nIBD+qqtad841QXdRPtELC+rFbBq7a6cLq6WQxcCtVUtHvtZUfhhpfdpyV52Hg23
X58LowfvvdaL2BZt1BaKwHlErWW6/cGFdjB57lwePQoUqriYbAsSLtv89/dzgR58O/DDYbMGfFoV
lDns0gHiY6eweIeSUE02RqgxUQNxBikoM56NfMRje+eF+E1lBwviPx8zDCwsCzXP+ZveC8ytNRHP
ZgRkPP3+w7jE7mLXwyDE8UWNty4jd+tdGCvCL9ZjSYJeFgzxjD9ElQ6yNf2ig7vdJkx74890wIWf
5q91+tk1A6DRUz6Yy7/UB1dqwy/kzh7ekakvaGRx/ytkeI1gvTwCmo4hMF+DE2LerlLICjqSspQF
DKJOLykwp7b6xH0pEZ90V2jG9g+jvcdBwh9l2u3KhgS7pk9p6wRgHfg3ApzSsILicUTrV97GGv8c
YRpROhNHatQXby4Xm9ubROSHVE3PTy7Vdjv5v4YTT4Gdz/8oBsXy3NSYa44EP0dRuouaUhhTRXze
BxtybO+NdWFd0cKdfEoC4G9xvPv84FYLtVx3drDr7ihuBGNHw70y2fhSB0LVkHXupjD1Ad/2goev
MnLGS1E7aWf9d4mnTy9vr69W9wx/l+A2gI/gRR2W6MJs8HSrSyC+7ZwByw14C0K88XtSkHT4eBXD
gGQ+BywIP09WyKFegVc4we+l8zd6OyTwvT8qywIepPjJsjNr1WYXwhQGXbOhuzNfdtdgXEkRMG4U
oIztlATRLhckdKHSuWxWMVq9QJdVDD6SFHoa1FiBam2kK4U8H+Hdykq0jap4aZobf1dWGNpMu4Qk
YFTAmuLGQQtnaLLjx6OZ99S3DlTKZdclvLdBzj7I+lf071qQ+8l0+I0LUZvTBDWptekposKyZdIq
Od4iG3A7/TFV/M4OZDdgGtO5c+BUvFCc9Pvv8Kwp00OvErKE5b8hys2+zQZ/aYvtzA1Smi2ZtZUu
s5eRFQyAJ49nVmR1z1XdCkDcNLwVcZQReo0AJket0Czy6c3+Nkwf4yY2Wc+WvbR6/MPs3DQJXSEK
Nu49MUNisyeHy6aQwf29TwkY+cHX96Z9DU2kxnzRDGYdkvuL/iMEr5cfilPVnvBWdKxJ8b/mU3ui
Y5Tk/51d7EXfebRGB851afnPngQ0iCPX3yrv4NU2iuKWvgXmULYzNSgUmBuco3JaK/xu8boWs4xe
Pup4t25anZ2djOabXiVpoEce4hUF5TFwf3vaySmJQwirYNP2vd+koW+d+3py/G17nCdAlRq+iXl5
1xQHfiPRpOVGWz3y3UBYc6QhlkQ1PqDXXxavNITKIBTUZSXOH6bP11BmwlAZ+ATIbW5mar0YSwwY
wf6EsOfKHEZOxboCtHjL8ZjLJdc8h8FDUTZm0N3tGdd/Hqx4OWHZSydmiWJmSz7LtQ6HGVR1CCSJ
RmjGTEUBxB2xtEAufJRe7AnTewLl9CTzIVRl8TO3ItqJuCQpfQ7JG3XOQepxnO87tlKljnjd8riY
mfK4irXtQ9LDW8jgIqxdiwjR6Llz5L6S327mLummofr63AAYrK5Z0n3KLNngfHyacCM7qH3ZPZXi
ya1tyFzcPAICP0f3cbaVGlWHWfP6GkXhWH3/XWkeBDLJVmq74iPFj3rdC98ilkuIgkGgDORIRiye
5d/Jyia2vkJOLUrePOUkNBMAmyAST2+C/d3kfUkF+RUyyupe/wvjNWNfZsIma5twNZYwuZEdrkwq
l4BnfVKwTSDNiKIqVnevZzcIBcfZLA+Q4ux2eZaToe7K3iCxLtharcr/fUJS31aXI3ggFxKugIum
dBr/WWjqRYCw0jPs8YpK7USML9ihAluPvlvZMDK7DH+ZnkkmsKWLFgkQVWcwEIrNIXYjCkhcd6Q9
DDSapIi2YJwWoyMs6q/ipr9eCNtzVTqxc59BKy6W+pahmyi8PS5SNdGXk03ACbQam85g7W1pIkW5
QDhUV0V2zNtLt0ZHm72HE+jGU+CruP2Uku5SPGbf7b6UbK+O3mKW1F8cL9+8KW+2DRkNjoDx+68H
VvSFzkaCYL+KD8khsqKl1o/6yMmjZOcna9Ko/f7HDUcPeMM1ekGraCSGmKoxTVnzhMLuIiVWR3Ay
teZHnIL86H6XVKSIhErSRCW+N26oD76cQwN6aq5df5/Cq8mEm0Wa+fz4HcgWcZg+l0EL8Af9agoM
k/5DMNxuyrLdRJeUJJcmzQKoLilC5cPagABrGCrpHdbVqNR7zXHFbV+3+AWre+Cv+rTGOan7rqg6
zhxKErMRe7ul2LdgbITS7id9GUzaoby3x5J9bwrxx1meRfIsKGY+9kDlq2yEwFv4FeRzWjbym7r4
RgvOON4CZH+zHsq8fDduED2OHTMdowU2SLNGB2XIDvF9TlCIfCA3jQXf74d++ANp6RFQN+4fBnVk
abh8/jR8I/WvI2yEds0UfUEHVRWfLbEdI0Qhb55EcjyQRlCOm88Wdd6cBgM9+j3b0wtlydEydbDl
jUD4A2luTMYhhNhYCGH/Iv/hQ4CUiKrJvViCNc1O3hnjoMPBPPvYGD9CkzfQoBO7uvSTBNZcfvEC
edFP37Z8OMQfsdIdi2Owm6zXgOgpjDa18yPn64XkK0gJfAUZ1xcSF3fZTj+HsAVU4aET0NOqMiS+
grRjAWbIacdxv0GjUXJ84fRRhVJhlUHGiusExWAWxvcQo2TxmZZ/Ik5PYn+s7hR0r1vhJQs78ovR
6uzMct2sCmLvNdCEKGShhrtAD3l0DEuPML3ID7oz2zmtoNir4DDXxJlYJqvRM2xtoxbWcitH11va
2Nf/tJKHsD2FVSbJ/k5HckHD35xoJFOjiezVl1OzIJ0qJ4/OV1eUOqFXJ7W2soXJbW/Nzlglx494
8QuLleHAd2/mFAMvRECT+EmYJwyQTcqRfLF0nJhF8IO7bTebqgfOsMNfP/gEtLzRTYRsmSBCC0zy
Uc6YA1RCdWNZvg11uQtB6dM0ZpWfRRIlV4TndQyL7dmfdPdqVLgvCbSCT1GPaIbqomrAML4bULlM
2jI1+mbA5Uk56GL8Limqzp8XZnAoD7RkKO9Kkmo/cjYEqyc2YkMgiTzsI7oiLM07mJeMbfwuegAE
d87yBtdmRt85ESuz4SjTN/LJQCZokYHdM7J1U62cS74BQbr/NQ/xUMI4Qzgs6VcZLICYX4WvqG3n
3nI2cEDM1AkbDLhP+r5TpqAyBeAH5P3+3hSZ8XF1UqYa5Oh7ZNWwkYzsl+Qdm0ilTk1JKHThVRiN
Ke+OstPTV1WIWiXSpMs9hhifkpi2mJsDpQeB8Gmq+ZTcxPZsVoketxp9Pe1wtxmtr/A+E1uFztoh
1SmLWRreHUmB+yp/i5rqk8V/FzAwjmd/esK3LuLciMPUX7QklNllMP4oKLZV6SFRamlpJnA2nW7N
tLIkXNz5ApyrhX7mbsK8FDdzzte4BkFZNKFGPve9CNHBxSWf943IRKk55NlaJFL0Lc53Bg24xQmU
8P2/AcBWDudFI/UdAU8vIMv1qhUkOTSJaQTnrtday7Xf1dYek3jsaDMGagcg1br9apXZtT9GyGhS
t+HgRkkUyee9sT4Exhwzhkg1Q7kvikkwmXvjWswHk+ftCOPP2IWE0romBSyIYGPKakAMSdCy3Eyb
j7KzVINzk3icJQQfk5HArLsrUwHER/9+FE9Q/5YSDVmNNzmP5GjmhjkYOEcvl5ZEYEa38rcY/u/y
IqDnqycTn5TavnuWKHp06503ccxRlmJ8W47gNvct73NDJ4B3Dj4Sgqus/aTLxLlEsUY7zC3TAgz2
u7yUlNTs3CNGoEM9mRzjPfVdA8lqHzAOF+g4f4ewfW0hnraxw4v/XsElvf3QIlzPiQ7UBqKV8nXh
phupuK9S2xJ8/kiVBbmGKqho62eWbqREHcWF1rSJ+qdu9XTsLG0NIo1bfzbh/SXVxLuASAXKUUAt
Wyb+XSln8WSsGw3sBjOLGIU1lRl5CAbvW+kabJIKCqX/BuSR/024GiO3PT5V9LEfW1lxp7Pst7vA
/bAqTHBP9ehW90NIBHCKXSHA6fD+7tsVuyGTSPu9auHOE96JatGx4YWss/MfzjRJPcC8oxjIC9aq
agEqRpuAYL83KfkHYZqotnrhapdEqCd4s7n1nje+BMigcR/yMi0+Zsr6viwJSJt2fnFGuy1XlwPc
zCEIj0mg+mduV+GIb7ZpnCGdu/cnss0ntRXzObYHFP65hX0ckesVw0frJuw4kl9rjgQSCZ/QKYgK
vlzZX05pVmamPF73ZLCEYtVmMAW6tmeTm4wep55/7ShBEUOGdATkRrPXMQ+YeRWpNjPucpB8Pr3q
Q6/Z8DAriYrrovIWA/afnahWGcKfnLBXQYxQ7lf8fEZ6PL8x9HGXKtR6bbLK/7hpJfMvi4a//C9Z
nBIMDKxE7jh022leXgs9jPOJgxpVbJiQjquFG9ZgcYb2C7jEbxeziMJYietRcheluFBhIBI0oc3D
6J23AnhIN71h+P93WiYaNcWCsz4fJV8To5oduQ4rzoSGW1WCtOPI/po2YVM4I7bfRrMnnjwpmFAu
hLM97SgR/NxHWMpvf7LkhGgF5hezjBGbVhRSfssubK6wzCIj1YTmdaCFBzp5CACUw8p9Z7UOWA9h
alMFrpIpV9PANhnEKEELWvMuomPAtOa8tCjq9x9+eDK653eUHMRzTaZIeipQ8daqgiK+ToNCpQ/8
Ynsv8tVj890b4xYKb7rjdTUPrfD9nsGBhsd8GVOs+0KW7OCf48opHggio25NE+aDj1U4m5lldftL
/NCnYDlFhf9aSRiFWPMCIvueGCayM+PljW3+rPwqaOjxEXYNVtdo1VHHzEpBhvVvfLrSvy6Owa9z
74eqtv59A3fK9N/3ptwAoHa9EZODtdZdLAPUmfEHVBTdj+aMwu9BGTpBjqMpcMSZ58GnFFmlPppB
K/zBv33OlxDEBwwK2Q==
`protect end_protected

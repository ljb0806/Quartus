��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y']��=�Y��w�*����6��L���]^�f�y.LR�m�˭�+T�%��ׄ�Sp����iF�Ѥ~�G��Td-(�>���E�u|���]�x���l�C&��I+��ֿ��Bp���x� �����WxvpІ�	XAi*z)|uu&w��nC��7��t�ĚQ_�6�83����ҷ�9a�y��A�d';ɰ�?��G�į�����ǟ�@�[�dn�g�^��}�zjW	1-5��C���B�^�c-����mhyt���eG�����+~R��X�����s?Q�*\�R�쌠��裖y���C�ɹ_�舘=O�$K�KQ�i�:7��M��-�w�A:�)ѹͺ5O���,�TH��qI�H������j�i�N/=��h/�͏��ˈ�] ��OSp��WnJ2M=�^�L:s��!iMh��6/AR��<��d�H��H��97F3�7?X�z�h`>�9�"��NAU�?� �	�.���"%�������ݽ�!����*�r���&V��;���
?0m=2�8��N���erGX�z����22 �d�H@S`!^�A�[�xr�����J�㊲˚xW��`�Vv+�x-�ǡr7!jQ���=�M&UE\<.��+������<��}��!D�j�t�*ܠZ��Ӌ����l~RT��A�tH��?q�$��m9f�����O�T�̀����XQ��[��X�(���#�����x/+�-ɲ>�x�fe0"w�؜�9J��� �NN�j9t�rg�ѭ�e��-�	2B�Y�`���E�0�L�-�(0����"���-6�T�9o�e�f�n��\�s�a�db\(�����H�rp���\퀛	��%K�&�^^0]�3LT2�r\&���G���/*��Bb>���)�ż����Ys|Zb���/`����Ĭ�L���o��{�;��J��x���:R�Be}��jP4�ȾOk;S
��3�8����j%
a*h���`g��e�㢄f,�bD	�<��@3�)���Fq��7����aY�G�f������E�;����>Y)��ע���&.������؞>9�Y�P��� ��O�Cz��g��I}�U���"^����ԗ?"��������*W�Y����jg�©��)s��l�Oj�1�$?��h�������yc�R��}a�Q�߳���佦��g>S�@j �n���0B�����jghmE��;�e����B��\�Ԃ����6��W����=���"]ؒ�;xO������Ow��J�G�#)�k��qÐU��B\����'���a�T��8D�rS6�J�;�V��_�S�0wV�9WF�\����~ �S
7� \ɭ_N,��P�Ɛn��=�9sЯʳ]՛��Mn[}��&ٛ��/��&ɓ��ơN�{���ttX�_��n��
�ޔrNQ����X��E�L��9]�R��W^�$ˮ���o\(�VV��3>%Q\��lX̄��Z�@�#>���܋�ĳ.�l덜{�?�}i��!qя/n�lK���E
)Dк�K�6ݱ(nj�q!�D�Â��|��T��)�+�V���$�۶'0�ݽ�#M�Q�n0nBQ6�������I�t&��� :���L%�=q���˘&5�����!//Q��ٌ�J%0%l�fWp�N$/���ɞ6x�uA B����T�zv
��R�H�^cPF��H"k�@�Wx�^���#��T-��a̪0�pQsg��W{\�2Ѡ�^�`)fʨ�ʌ%w�f�4���!!0�"Ħ])UO�we5�����~tz��h�}��>-�����(����׍d�b>�I6�~/�@Խ=��B��J�	��d�� ��_�ף����Ъ���K	�C���$�p1ɠ�;���*f�-z6���5"ů�(�w��cB_bX����82GV�'��U���)gQ��)��m�k{7n�Ғ�<A%N.��"�<�|��G^!M~	'�� �;�ks�b������ �9?M_}��_n3�a�'�3END�) 5�$Hծ2m��U  )��Vx�X��)7y�y6�'G0*�n�5�S%�t�*U�+n�.�S�O�c��0�
mYW���#2�y�� @I��n��j޳����+0�'۔�c�+�0ִŖK�O�i���!�Nh97@:J^���Pa��єH�M\�7`��*l1-H|���v�˿N����EcB��4�r�t���������Л��m��1�K�_����n��%��PK%6�l���W�ȟ�-���l�\�I�i���[-�#QV�d�����D���y�8�{P�*�U���0��:r�����$aw�tHa�t��	��A�%Z��������#Xvf����vCH��I^��NȒūSK��Q̴Yv\���͡� m�y
�����'!�	"n�XP��I�m��=Ie:��I�䅻�ۜ�@���'�F)��	e۲�i�����J��C�F-F��V" ��ǹaEX��S'��C�D���x��I�jmME�����j�ݗ�)&#��9]3��f(���
�l��Gحu���e E�=J��ߘ*_�7Ex�����An�L��D���$��;J.��kù��cN��:��>4�g	X��G����� ��&�=��S#M(
ʼ�>��߀s�Hޟ派��~�.֊7�`�i`:���ލ5�ē�tPx{�^d�62�����S	:/f+��5�x�j�:�A8�-�v 7~��cq�$,)�|�m��b�$j		giy�V�+S�V�?�g{�����侓l�a��~J]��@��"�<7����� ��!\��8��gH9'�x6_�́ �o��x��/#���A�	X�n�&����	N��B�ʘ%�ţF��ɢ�����y.��hp����#!��x?�`���;���}g��@��LBu��o@e����*���!yy0�;e��`�;�R\�_�~{Y
0���B�^��������l ��4>��k�Y;2���9�K��,�j�Q��W��wD�6�8�����$����ꎟ7ҡ����� ��
ǡP��5я5��s�Dc�i*�$�ܷ�]ibe��<vP�պ�Rk���$�0g ʈM�)H2�׻����N����*��]�8�g���f=-���X���$���y�՜(Х~���s77�}��A�5؍�o+�Jk�X���u�ܼ�jL[iVK��@)`+uΖ��x�'�����jM�|���X��0:'�I�AX>5DZ#��T�^�`=�nc�ݤς�y-M��^��1н;�z"�5��	"�-[^z�H-��mY/��ja]�\��������/�S�N�VШ��	��x��^j4$!�U�V���F]�2Uv�����ܔb�f��3�RQ�[�S��5E�yR?��ߴi�Ӈ�ͬ$T�ĳ�cC��^�f��wA��VRe�1U=���@�"����d,~�{\Q�%/�)4��ʟ������G��J��8]���-���Az�YЍ)J�oļ��M�(1�8l��$�m�H���>$�^���Q�7��,6!����["��=�t�Y�	[�ᵚ�&Q:b��Ej4�9V�x Ѐ�,zx�S�2a�>�;v���$��I��XJk7	��;�Y�ce����0j:�|�a"1#~�P����͌YN����������������=\�+ˎ2DCL�ml���
�M�M���̓�%�4%�$� ��G��/^hAhL)��Q���o��90x��T�I�^�n.�{�l_m,B�iٌ �(G��
"���j�+�-��.����`_�?J?.A�P+�k�k#���:HC����$�.�ܬ?i����4��Qtl"B�KIc4f�?T<v洟�
�Ub_�FoQ���U�!z��@J����kb\�
|q1 �("�7�ˬ�[c���`�(����fv����~�m��{?1�V8Z���OT� �$�&a��~|�bp]��.�Jj7�4�.c>018@iq�k^S�z�!��x�� Br�*X����s��AC�Ԃ���MQ�,��njĊ�5��W2�7T�|��d��	�H8&���~�#@Մt8��l�����q��XhWy9,1������2)n���e��F�2䴼]N=�R>�)��=�L�\��n��g�O�1g��$���Eag��i�����-�4U��們@��d7�Jݬ���m�Ut�8IN��(K���Nl�<�LF����ȉ�Q�Q.ah�.(-��C�����ߚ����
s4ORQk�L�p����=?.3J/M�1�T�d�hF[��ᗊ���>�A�x&iKTe�N��&+�׎qSjF���n�G�kL�퀤q�P��mB��������晖��^t����ڞ��d`n&+��J�W}U/�Iy���3<��5m(~�S�����CaXFO���x�"�٬gC���BpA�!W[��#�]�<#U�&?L�tF�س!c�~���A1翇���I!�,� d"�n���l��n��"ɲ�`>����C��'pjjk2J��/��'Y��� AY�:�V4�T�@��,,a �S�i���x`����m;�<��M�� WĞ�E� ����5�$QL��S=Ƽ�M��o腱b��РK��Mm���m^�i�)�P6�M��ଯ�(��S�r��;Z�c�1H(aAv��xԩ�|�����������x\�Dx�H����}�� �Pmg��V'-]�7g��c��n��@�Ƕ��Ud��bS@g+�S���4���Ӄ5du��P[T(K��A�0�OZ%Iј�P�������J�e�Kǁ��{!��5jX������#���7y*�j !R�Ug��g�onG�l����~LU�:]���0�ZUh>`ӛ��5�����Q�f�{�L��]?Jo'�	�l�?�L�Q�.+��A��lc�ɡ��	��˓�,/�];�i��Q�pY��u?���:�qB6z��@��RBt�ı~3Z�:�Z�]1�&�3lqW�a�V#�����'���"�|>�r�W�KO���%���SA�-HϘ��f�_c\�h�n��`�P�Pq����:��p��Y�Z4rN^������S%�L��*���$�w��a�8�ʓ�	}Z���7��|v|�R��-���N�+�Ņ��	!����q3?�T�5��ç�o`�32�Ζ�ޢ����9�����9���F�i3�bZ�"=�ϛ@I��mc��~DH��F� �2Y�-F�ϲ�k4�ُ������Ȳ��RX����V�[`�-��݈�X����~���6�%O8�d���ƭ<'�~�T?� �a`L��� ~��dK �࿍94�|�Hhz�8����-�hYN��/�|��{f�d^�(�ԏ4��%����q�Wͺ��aՂe�W9ȍ���#�-�0n6G�����%���	�JW����,��b�O0�)��Jׂud���;?�CQ�����}7�VO��8l����u��s�%q�b��Ws����'#
9�P�i�
�W��>X@.wQ؃Al��]�L'F��6
�̩lo��7L�<`%��B�]�;�L�u����m8`��A�qx����b:�-jڎgC�����
�3�05��J�c�����T�g�R�Ѣ,�Hok<ۚ����+�c(�j��u��b��(�E(���tf�h?	[�H��+vj��;�,A�a;,��1�^1��{�a�V�3Sk�К��wŪ����l�~�u�OA����V|~h�.�l㞊~�l�K�H�E߿t�N�v�X����#1Q�A�7o��w�,��Sd-jQ|U���[C5SZG�����n�ໂ��6:W��`�������Z������V��7�j��b�&O�:7������b��_�j_�i�?y]IP��O� .F�wP�b��;�.[`\�X0�C��x�0���i�ԓI�.�Ma�'�p%�\�C56��t���3輂5��A�@�7s���RЋ��E�s�]VTy6vе��A�����]C\����M{eo蒩Df��b��A �N6�*rc<h�@�>U�i4�ܢ��C��ߪ�QiCi*�:hj蟌3�/��,h��QH��,<?�&%حQq�A�����^&�M�؟��y��_ 4�vz�2M�%�H���."Mx�>#�%� ��P�쫡c�,Og�ȞR;f�?��B�1�:nm����~j&ڡ�����ػ�.]5��
}��C�1�����^V�Vj�����yb��uƺ���*�����"��kš�����?8��9�V9;hV&�����פ�񔂉��:��ҙ��0�c�H��*P��V_%6�Y5�ג��S�y�����s�o|��s�`�r�E����C�!$窺`e(0j��ʚ��A��*��8_ ʩ��{)����i�9�����dp��+��>����!� H�%M�H{~�b��D�+�@���T��j ��ЎcH��G����Uq�ȄX�v����' h>�'.�"�P�E�!��W٤�a�� �-���f	#��:R�Q|#��������4�s|�m-��b��-�
M��	$C�c4��HX�
ز���D��qˡ��MfRۛΝ)�q�"6��!=ŝ�~NP�Ǧc[ȃ_�%L��t��m���Ob<��6D�1v�uWK	�*$�!��E ^��޳5y�ys�4����-[r�I85�@�P�y��b�j[Ⱦ�˱)��)G���{�A��}B�����5^�k���a�w��iC;h�y �C�i�$_�jE
��S~�"ml�W+�&��^����B-���Qf��V��$��^��� t� �l�����nG⠡�.�+�X ����`�S��~>��r��X��u_%�TW��S��=YVe�t-��j���2Ō9tu��Tj��]���5ң��p���eB��n��M��B����=z�^�T�j]H��p甩�`^7�A���b��WW��'	�;�J��� �&(�L##z�d��$4�=_R;����P뙜��������]�����W��l
/�����W\&�eׂ�cʬ��N���.Ƣ����B�`�>56�dܤ��E^�[�d}ޛd�)��I��M
UjcH���9�)0H"��T?���|����<S7�ڬ�Ɇ��~�&gxd�k�%�Eu���6_t�2�w�:��F����҈�8C��xv��_�v�E��5/�&�����Cϱ�����nm"���6\���Q�����3=+Yk�+c������=׋	\�Uj�%R.ho� ��@�����������Q+�~�6s�S��$��D�`<WA���ԙ��{�	C#J#�����Ɖ�q�*uӖ�fE�,��&�/�*���5;��f2j��Jd��֙N[���7Al��V&����88��~��D�a�Q�%9.B�M����N�u�J`�S��"����|XK���s��N����;x:�Ex�~R�M��9��:p>�/�?�=�#q��.�ݠ�C����l6X܊w�}�D,�+�B}�)�
91�I�W�܍Ky��J?n^� ��̷�qwCqo�����������*~��2�,�j�����8{%�̽UB�adə��WB�� �-D�!�m���k)�xam��2׸$~T�ތ
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y-=^��l�y�KR[�q�$���`L0�y�T��2)Ǜ�q�s����n����P�T���#�W{��2�y���]��\(vg�G���a���P{rx�^�\�*�L	�ᾌ��.�.-�LwCrW��.�xs�,-��j����	_���k�d{�WqV��	��l�305���B�Q���)�q;_�_VTK��/�`6}?��j!�ZsG�X�	�$�Y�g��&��q"��@AZ�����k(�*�e��t��;kh������'�Ͻ��u�PN�d�S�v-P2��t͟�#P�G~YH�
lo��ۀ��>�bu�\}E�Z�P��5r�%��Do��/��3���``�cK8�M�qO�0�_'�r�X������γ�3�~0Xx�I��(�����(�f�����L��ki��DGg�B���պ��`l��r��e�i���;Σ�y}��M��c���6|�JT��tU�����9
S����ϛA���u��C�Z����x���� @��_�󅍻�y�t�����0\��k;{���'��:n�A ����+<h������X8���X)Tg&��-f�_2�a� �x�¹�����!��ש�~�`���-vF^�!h�~K�Kmo�ZE[�0O
�e�>�p���p�����v<e�_v��^OJ,����Bg�������6Ԡ�*&W�X1����F�Q�R]Q{�?���}�Ѧ=��d`o�{UВ�wN�~�nZ�+09SM������dd3.��K\T�S�^=DL�<�I�|��H������T��N�{r.j�b�C��V?�HgL��tCA��L���;�]!඗��#���V̐̋��w��I~��"��/���PW�U�Q4J�� 9�����k�Ɗ� ��f��"�?!�my��)�|��]�G1���5��i{�O����U&�l�4+�{s�?�=q"ȕ�(�O`�Pc0=W��?�b�����iw���KU�2B/]����S|a�}Ø�9Q���7e~S"v�Y�+�kY�Sx���J,\H��b^H�@8���o��J�t�o���k�l�2+�p�\�=�Pp�K�VÌ��!�@	NY���U yEf_�@�<�N`��qbz;>�J��X�M���z,0�[)��u�S�N���&l	be�q�p
d6M�g�7 Aq��HO1�ޓs�f#X+�}	�὘��Vj�w奄l����'!�у��+�����'P�୒mb^rC��@�1�bh~����F�!Q\�3�,�A-3���غj����4n`�X���*	47�ֈ�� !3?M��1�\�����Q�h��~{L�va�3f>O�`�'���r�9�	L���`iW���d��V�?������CXV�?yD�>n���d�"��p��'}�Oؔ����S��Nc4�ۣ����b�v�<�EjI8�}�j>��:�ђ�e(\�0n�|�I�\� +�O��z:`:N�� �����g��Wi`������}�E�0s���;��M<dz��X>�ef ���:��<?��}t��M/m�-��|���UUH.ʎu1����/A����p���sz�.���fl|bl�אZ�&2V2�� �� `����4X����V�D)�����:*}�3��̭M������h���R1|��'h�ݹ�|�7>�ΰߖ��I���7��Ce;�P��f�\�UU̢&�@�UQ��1��6�y3��X�o�_����Ww�Q�u ɀ�L�=�4���l<�Wz8�D����T���R��2g*�nAd�rG�;u�I��&��5���B���	W��R�&����	�/�v���b)�7�&yؠk1ùy��x��Ɠ����t� ���	�K{�2��ą08����
�etI� ~Ȋ�OP!�d<,{h��E��3���Sn륽�b��L�K�9���O+��	5~��[��a�'��^�poZ,��T�n��ץ�P[���ZAՒ1 ���]
��SW��g6�4d�/�F3��a��ɢ44����υ�ԙ�e\�-	,뮬"��"�\�X��f���M8B�Kn��w��__:Gی��[�R�0���Ҝ3Nb5D��9|��Q�>�ͪ���l���V	=�X�S����ze��3��@|/��t���1�ya�9��ibhaıK�4[����L�yۚ�z�,g�/�C���x~+��j���!L[
C�[��E���r�N���U�n���0:"����j)`��-*����h?'ש�Ʌ����h��ޤ}����;�)K	ea꺦& �Rd�y:�`U�2��DΕ�n�/�&v��yH[R:�i�7�r�=`9Zq����g6�io�.D�c�@����3�E���ݥ��lp�ް��y��T֦r<���TC����D�(�"�n|%}�+�>xnt���{�#���q��`��n>uW+6�I��V�rU���D��1�#�[�eā+/�A�)�c5t��4غ��n<��R8���^ڋ �������F�����$��l�װ��W�߁���b	�r�]2 =�,L�p�,Xu �o��s*~
P�jE�dDm��Z
�G����6����7��<A�ϵ7G�y
��HA��=�l��ƴ�|�W����������1%�
�3C� ��W�gJ;���\7�~*�Qԓ ���b��_'%#�H�_y�ګ���ع�E�&s׸�y~��*�%1�R>��-�%db[����Q�,�?nz�j�a�`���J�`9*��?��E&_�_!�K��v���~�U���z2$�e��$�8Y,���0���8���s�jw^p�0D�,L�g��FGٞ��2�[묆w,�_�v�~nV}�G^�D4� �E#Xo�ӈ�����|6�;a���s�� ��<eR�o2'��DY" Q�NF$��##�� ����5~3�Z9�Y�")|�,�R�\僨9���뼐^�m�E����$w#�	P힣-��v{M�Kʞa�#zUÆ���5�-H�$)�Hi��N��+�Maw-���<��l�L�i�-�����j0��1"?��E���V�v�h�LU�A��w� C`�v� $�W�D��7�[�%�$�cCT�3�C>�����؈)r�	=���~�Bb�&�8��\��&:�g����GĶaV����e��A��L��?8!�����#�&)�X����~�:_fmm�ܴa T�V4�ť��S��J���ZL>��G+,�N@/����!j�QF5� �����w��,�$�׀�7���f�D	��f9����������:_���ۋ��Ҵ	52z/߿�-��g(���&���3��W,�]'s�,Rf��m�����K`�1hÍ51����#�R�7 ��ldKz��`_�����PZ]�m(���G�}���s$w|t>�#��Ѩ�^��>s�mț�_J�x6q7[��y')
Y2GeW8t��po��p����H���-��9>'�"e����H0���@7L��
�\��f��9���/�~�
��f����*}�%\i^� ��,1躍�W2���g�ʧ��� 8� ��Lʆ6Y����Q�t܌{�z�l�U�s�����w��Ա���iDT�@��g+V~1��A`�n5��FXieg�w�rxZ�C�¥�H�V�n�M
1�=����;�e���!�]*�Jf|��������q������h����0Ა�,��+� ���/`k�
�nR�	��d��Lw'V��I�a�1��0f�(2(�<&�+�\�H���;��6�)�8ñ�\�WC	�T7�.���@����t2��.��>��W��a������9�e�x�%��[��<�:9�"�`���׭��-����(3�la�I�3؍�xM��E><<W�������!³q ���rW4��J} �����q�N��N����Svjt��-H�_�W�����*�{���L�$dz����F�2N�Ū.�|x�l�/���gA=b��&�&�wY�z�O��ύ"�K�qw�R<j��)��Ma�­wbm�H��5��Ͳqo�9���>&F#��Uɗ�H�dQ�����{t��|�+T},��o4v�)�H8C�� vzLƊfs'@�_��40���H��[���!�x�
m��/dR G�V	��qO���AH�:�Yj�?Ձ������!���U���;�/�d��i�U�7���u]o)��C�p/�����܂q���1(�v�A��g���|�d����Z��c�2��{,&k^�����Kk��<����h�������*�O��V�f;6��4�X�e�����J�)j'��tV��[�>,#����S�E�d'K��䲵b����d�hL<vC����+�Mٕl��wx�ó��^���xz9��8N<�Y�- �k�v��n�l�Y��ஃ�w���`�Ջ�b��߰E��IC��� ׵�0zHHw�:�o�O�.-u'��m��s@5�}�n��xˮ��/2��:�)�0�#�ϣ�^�
}�n��6˧�p��~?�Ngևk����6Yp���7���}�3�BU�n�hd:��Q�^Rr�7��O��;�9���0��b+
¸�I�$���g��E��H<�N.���Z�V��3��H�*�D�$4RVX��5���8{.��Ƥ�}%$�R���.d���~b-�*��?�c�>��{�vwP#xʊX�r�
�S@���`~Z�y02 ��㨳6wtlf���A�ٯn�������b�x��yB$vY�M���������H��8��Fd�y`?��jZ*�i�a8&�R\7���	�P����Հ�y��XB@�}�oq��j�"uu-���Dr16�,M$�j�0��g��)�ga\��P�}��@>Q�� �_�S��G^�/*�;Hd'M�|���u�?��S��A�X���IN��Nѝ�fޗK��)�.��[��s׬����v�����N�d����8��Ξ��jJ!,-��f�},�5�Z6�ޘ�Tʘx��R�0M��/�ذ�'"�M�\3�A��'����T���q�~�w���[�=z�A�[�Q x2��~M޳!���Q����NI��^a=N����p��Pb0�c�!s=j��Eʒ�f�)�a B��VL��;U�"��^�G�q���N��F;�6�݅R���e$_�r���W��9��L��b� ���x��g0kz0�yR<��<��sU#����r�a%�ߩ1>�T�>j�yU�������@B�/u#����$~��
�����~�߻%���-��T�����v:�C�d���L1�����4Ҝ�Ff�"6W�\�)yO��^Q��e��vtA@�ˋ����m�ʥvb͈�S��2��h+p��%������R/����U��1
Yxc[�&M!��\�b�C���8�KC`����r�n1�e�8.'x�9	[��Hr��X�湗�h$rhx�F�8+����1'��V+5H	�}�n0g�G�a±'cr��x�gw�7�����!*���8_;;����)�LhV�l��~op��H�C�~�|L��S������?��O]����ne��}i"F��	����¸D�L��[��@��,Q��f���!}�$YG&��7�K,��t�W�2-��D��������rDv���D�Oe��ㅃ�`�Ǹz��?
q���AYҾ|(����=:}���c�4�l�3����C��m��Q������s���&"�XTy�Z��Lѽ�� b
�v7d�2�e2;X��/�XK?&vG-�-a��b;��Ki��Hf�����v�o��#��C�ڔ����vL��B�������>I���L$!�Th�yܡx�������n�p�<�B���3��.=-f��Ŷ��I��D���E�>Q��M;��6�+���gS�ir&+�҈+�	���oRr�2+��u$S�{�=O�����.��5^¯,��zt��qY��
f�xd���F��u�؜����2�ras��:��WQO��Z7k�Y�a�� ��}�����1��Y��sF��_C���y��+&��
f��� 	H���[g�I,peev��4�B� �,ԃ7o/�wBF���Ы��E��ۅI���6��z�go4����뒸OQ���S9��x".4��VO����r��w�j�H]8�h�^?���j�l2U�a�Q���$���ݥ
�j�j>��ceZ�u
��Q�]�qA�{˿9Ԟ��2�s���m#%M��(��եVb�w��#�,j1\[#<9���,iT�®p���%>���5���m#�p�c]�DX��!��f>��#<<6���J|���h�����=3�4\f� �A����R��Q͉
L����-���FJ9����iw����{%��� �D(����8���/���4k{u7����-*tp7+\ȿ��� ���ok~C辋����$Q�7������v2�1�?Ɨ}Q6{8����Ll7VF���ӻ��Z����'��v7n��)�e:�B`�#�5 i��S&w�ה�"���=��|x4�6�S0(0����4�6	���\�<z�Fw�
U+v9KwV���?0��;�Lv�,Cm-����}��z�����F������pچNf:���Jm(,f&��׫���*ٹ��%�B~�$9�5��!ʜ����nv��y���Ŷ��R��U��-�C��Dڅ�)����!Pb���uX s^	Ϙl�7ag�!�3W��:�\��&�O��"h�	D#���+�ʅ����>;���%�b�>�)y&�i�%�1"r]��q]��p�+��������qWo�$ �jKH;œ# �
�Znf�v�Ӽ��s�Y
�d�N'�zr��1*�v�y�is�Ë�����2�G������\����S�D�5b�nt��I�h@��jZb�LOޤ���{�EhA��N����oE��,�pw�j��|W�2���V�JFk|�0�&]��B�5��n�=�iZV�0ϝOQY,�`?6*Po�㳊/H���ZXd�I���S���"�ZtG�r�*p�;����'Qj��GA$�"��8�	Ua��I�m\~��p4:c@x��08�サ/l��h����d�<֖��u�"�0���{�\���g��T�
4'Gd35w>:ĂN9�1n[�!SB�k�� R?g��MD��v% Q�`׼]E	����%vT��O��� &#�%p�(�E��)�Kp���ʹ���a�z�p`��	PAx@�ͳ��V�y��rS� �I����Y--\T�%��'�iZ�\�M,RL�z���Nۆ�ع����$
�`��.3�)�QY�QwE���v�*���h��Z-�/�!4(�"EhI���<2~��U��R�����b��I�ؖ�����{�-i;q�߭p�X<}� �l��o"�D@���/��sL�~�_>�e���Wy%XK)�_��T�#�`fW���ƣ��(7��im����ɔ�Q��7CJ����>�>��Y�h��o-�xq�49�J{R�u�����Z2�ކ�UwZq��sZ��+`&Cz%N��0E�Nͨ���]O��pTVľ�@�#���%�4xX%{���r�`h�����
D������-|K&&��m��H^(FlG�ty�H %��g;蜠[��H�f⪷l �u���\����n|�+_H��������F���l��۵ݐ�\��5$f�|/:�4�"~1��e�`���zkb�OGK����$nHj ���<���O��Zkb���ٜ^��f�V�N��5�޺��}�����?�o�_no���~c�pU$-�gM��]pĈ�Ŏ_r�D�V�{����^��?U>���yңcqfYc�t�mPs�-2N�Px{A��<��CZ����1�&����J�V�~��=/5�u�R����mؾ\]��w.	��  ��"k�-5����f�
E.�t�&�]�����+ʶx��*Ä�H�t�> �	��2�OBB�u�v;�d`���hݧʧ��.�W1�R��'����¶�5v�m�~�	y;����0��)�"�Ɵ�="?�n���y�ʒ�@�?�y�����$:�G��n��&���K�1a�:>-K��I�Vy���B~B���j��-�Er�R
C�H}mQ�L*��_=�����7�GJ�s�D�"�IZ:&æOS�Q*\(�d
H�X�TE��+N��1/�}��2A����7a�j��\6��h(d��*��E ��K;�,�+�n:�W�W�n�ci3�}
B����<���zܔP!���oE�|��� �����
p���2.t�5%�>؀�B���3>ި�@��ߑԚX+����7�
>R�X�~��~i	�O+��զW?�����<D??�7Om+#��^.��:�8��:H�l2�;i�_dUL�=l����}�e[�x�9E\#�S��A	$!
1�"�E������;�=�y�5'���2���΄&i-t�y�<'��G���n/�[{�+��ݓ�+[�e����y�"^ ������a\�w��������V� �6��#�̞T����{��Z����Ԗ�J� 4�4ݝ��E��l��0��0����m;�-U�aZ���+���E��"�pڶ���� !7-�l0�	�tg�	���ގ&��='�V�QO
�fn����d]�'�g@T����ŵpl%��Dk��
�#1j)��t/L5ء�����{�O�.Q#FD.�P��G'��8��ɐ�_@�織���@��
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
123DNDKuCD6HkUpfrzLbpa/zgGKn2bpDCmIIHwxe9ewJwRp0Djq2OFnLrwboVs0v9zsY3QTSPiYW
smzlPUFKfw7uFYwlMoHuYcjRgL8I9CEel+qdXOuLE7/Nw/GzNVQR60SXT/Jx81nQVTqwDFN+EE4S
Q0EmJxjzCnyowGklnG0Z+bkYnLuU+WU97W6x8iD6cSK74AlUM9tzgBcJGbYrAgHnyqIqqXRGJhvV
QvU54TJXz1wyqOJMLj7sP9lqSGmyuXIZCmKJmHxRUBQttIzdyKrYM8c/PlVhNAX1DzNU7JtJHvca
4EZVNAEkaLk0riBm5x34JJ3p0UArd363XetVNQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9472)
`protect data_block
QPmyM9i9xxr0jQK56XFsMJ9LTWW6zAgvAnDf1qf9diN2aplfdGyZjy0v5DL4lScP/pWCNj/QqXt6
MIH3k72886bufROtPhDnD2+3H8774uKsJ8Wg3C5T/gA88CuXJhoDNQ/xDFo9cbbPbguYlZWTaJPP
CxJQfIqxhs2I1AllG+CLR5l9XuuGQ02Y4s75zBDDQU+vt2mj0GFJZwOWd7zLByCImvAhiuCEX3kD
xC+nmUuxQneVNyTZ21P/bEq5Reu9fFhjp2JPsn67xosPYkZg+rDWC4Gxrm4loECmlm4c2zQWbKoB
VYODtRfwiv13n8IyxdCu/bmWeKiKUzDnTeIrZuBIw1+tMcauyxMP2nAk2uIqP3QgeVo5ZKsv6o6Z
fiYJtNELcIOU94XHZA9z6aFEY2P5X4vsS5OfU+Kpc3V2T8jooLTZ8yinGfg/IUTmLtdNwwrF7PPO
oScKp7ij97ZHo8T07H0RUsXJNgFvrj4MpVxEhoFS5DtAIdMMDzz4wbr4Z5GaPOg7YTQOWi3bNkNh
CV2jipkX0I3OPWjuLmFFH4Kek+iJtYNbTbgXl4L7QzyHmjD8oHuAmPni5mWQ/O+R3CpKFMpDKGJ1
Qjc2F5spIU+gPVktWQVl9d2BRBrkIDbaUlDA06gnGuj+5kd+HFl/+oZHgw/8S6Gz4GstCpQnd67i
5gyPTlV1PAjEwBIB/7a81xHlt/T93VdFHoC0Yno53lF9vL2D3cVJY7KeHKM3hDECeA5wAFBo88zV
u6wpv9PRaMxk30a1RWxavs2MHYUixAfU3b0mODvGwooEXPAqg6ksyi0kEjYOQ/SQfTcoyiDk5edc
0rJloBMLYjkvQ11XEr/KOucekXOqQLF45/fgyKvj7pLjH48uxVeMhtp0Zq6Sn3uN7suFNlz+nAcw
pVsKXdrHWBlQFASLmW+SJMTn4L1B70/Oq9IXCeg3jsxN1IE90XLwOwXm6603ymxyFVUPdxDm+M0T
KHJhKOrmbo3wp5x4fdLJwjte+/gBYhZt2s6QbchjOoBMiJ1cBPBjg8/1HKipsShTJvX5qI2ecUad
aqUogOPkJndM63+VEW0rXdP6WyMnuO6npiyb2JN79OJwMe+aUBF8kdhsgaLhhuoBc/Bz+6aqH8bJ
WD4/wvcTvZKs2iYZkS0gFErJCT/p/641VS+5fPyYC80iIDmweKfi/nyWHXAXBOCo220SF0oYSozl
VhhrmuOi49US1hCDlbmfG3yegObLo58RoTbvUttqDgywVulRF/dd69n0i2XAEcGPWl6OxYWWfoiH
wx9xYOn4QIevRoJc5RsSrRFcDjDEJZU3dkEC1OyKOVcm3FAFg8RfIGdtJWoqVyLw0y9MbZJAAaxW
HG6hL/QQBsCH0WxE71FwHFI+o/1qYcpQX7VF4oeja+1uR/LW3ZrnWAn79vSkt8J01TniY1yD2AgB
7+r0KcdIHZRS6uf3MCF2mpxVMtrKWA9bB8nN21KSVyKaWp0bNMmh7aE0u1R4EK5QpbefVO0i0q+Y
hCnO+EDitLdTFBxQ5E8MW4kFJC+w9a+LiGibt1UlZKe9ld+E2jHEC9Zyr/CMZgHdY/5j55ALaCqM
T3QVj6vneQH7JD9DXA9MLQS3nBC8OfMrGmk27OJqzTpEpeXzZPKtCoVizflJflrmRuOHy92XVLBB
DdbtjhkUTLf6AHo1PLQgmXilZueuI3zbf1fClzirpfJo/vQuUI0+QPbVvKnNs6D8i4kqZgMRxPJa
CvKhmjnEaP25816xIGjMKGlWtdDQnNqh/vd2sCoMZpIITNI1SO2Yu1T0lM+23k43k/gqwcfLE3Gd
7nsru2YRK7kbfItGdRUZU9XAB2HagzxtwErOU9Yf79es9wXXrLE75jnLOmXLKihYwVSJKNq7+iKA
/+cGbURideBX2lNKYbeaIiQPOxxf1/MLQkqnajIZrAKQ6S8cIkmR8B8sCiU6LP4MZyZGC3gUUm9G
d8tEU5ABu8mqBZaFgbRYQqEqA6FrYrMmRfKqnuLxGSl3CoHS6X1y4amvbczX+umGBhmckVnoldkX
4a2hPtKXagmFjqdbb/GcIWFV6UZqdM4VQGuBBif93y/zjyW/zCUfnfvPNuaHnho7RG4SYcXFoYXW
oNI6QGndFZeKkbcV5Lm29m+N2LrsdFZfgoqR/3KQwhcNigUl0WuHBZtmg//EtHYDTiDYCiPeH4Yl
+kTVGznl4tqJWRjNPGr8gnsNvsbaXrGTCHFvoPvHjfJJ+PITujNicnBXVi034/2cbCVnZDd4cngD
6BMBE/f1XqP8mkLZ5ziZBP/lxKGQ3bjFjLrkt8kA6ipEZkTopqZwNc8zbMFBPTVELyY7XIfs7aqn
vPihdwu4IXCqy6tM+yFdYJnXDlAckXLh9F1ijuzEnVU9skjwFv+NZ2voicFp5WafXfrYSFuYlESI
zfP1dwmw2zUUE2bQh6YKWBv/7RmrGHNNrJTPBCdi9jqhdvqrjMhKLV+MOxmMxcppYQ/vLQTd7aMO
wyxDa+sojT3N0fv3+xk2LvyG2pyce88XpII71s6NEvmf4NgOchiGfa+lhsOQXszP1WA3VV990rRN
1cY9N+f6Ld5i/l7wLznauNH2zObE22P6WxHW0eRu7NSblh4cdEvZPvNHxjD563Xj8ckCp4txEk4p
kbAupM50JTf8otKpi89XyYWYD0ZZjhrnYzZC9VHOwSiYi6ZO74a0CD9i5K1DXM3bi8hWX24L0Q6X
yuVXLquJDw2k9COb/YZhmpCmQbOIzXurqV9ONNK5d8S+1FWIE00IaD8sKlQuZaF/jBBz6RErOXdN
8R5uGLYSL7QmIIxs/BR0rkBByj63fE0adkfxYXoV6efLopHSgCE6vCqDxstMGxkI1mcht1nyrYdy
tOxZ0+824eys54dYOeLI+Dl78OoXAXCqpNpDzXgsOp624x/bFHFOifIUOEfY+WI9mfO9w8HfcJLf
Aw5ZdadoM59VP2tm4+g8Et01tqTE0tHpCHV6bWD8u0lJzTdwSAXuI2JkyQImLMogLq9Ntj9/ZkSE
5j2GfmtTRDYGn1qMIBg9nhHZdaEZsoJtg/oSCAhYQ7sGw9OggFEoIx+PEomM0M5yzvKaaOnQH4hO
6zCQg8u02mbyn9SVunI82BdKm59YN/8SPrNqFsksPbhnBZv/AqNClPTqmuTluOYDdPKQJ5aIri5A
fN1xbpxqNrkvxkJGMYeL8TobrLZ/quy/VGdShxwaMlnVbgwYmLgfeQimmpGyeEbIX/lKg06y5KO7
GTZt29iAnwc/Bd7XBqXLUApmZtRhfircaBfza9f06zU0cUza9cXJoOWD3D9asLBwJ/vjcGtrp32x
gbqaeQV/PHe5Q2D7/z8yuDiZquHy+hHklXv3zCs45v/OLPeA4bJ9xQZjzbnEVAxkwpvfFqQFYj15
RPUXT8h8QbeO0x5jnkhlSp4rPF2J6gObx297LqXYU7qnii55Y7JU5pMIhrCj3IwVPjEg0ByymqLx
3uUr5KYmgdEGbFQYuZ3otHqQgDwW5Ln0Jtxmg2pnEE/qvfwYh7gVb3SA3WL5jmbSDWsc2Hk8+NRm
BR4PE/wYt0ff1YzSqfV2DQYW+0K+UU/QofAvd4uKTjTcyJpWwWJf/D+rQafwenY38GjmK9qv3P6w
oGzDzBMqDw7Wfy9MiUV9s5qv9ZDVTp7ZoEBm+oF2UARthjUneWPm9OKR4HtAHRP+xbrKDFiQ9O8e
y94Up4AgOgnsGaX2Og9VYlCGvLRBQujXRmN6hOcQ7iacbtj8QNDlII7wEh11RP7zl3w+SA0H4Vv6
jtXEdlKsaFNl/CYKDHnYDKzHZZLp4gUWTPFstopqaIvm1EK0FDXTUJ6T+5q9xUNMpgxNBq6tkaqQ
aNqcEkzF6Q6Ie2r6zObaV5PAhPfoTbecOi2r250tK8EwVTjHabqxx6QBJL3dMVUPvrHM/Npf1lF3
lLn0lW9XEYadcfAJyxEs6a11mf6OOQYm4yO9a3tr2yU1qViuSyFwjExJbbAAx5x2AM2/O5X8sW4v
LAqE0ptXX6GgVjRpk2G2ZAaQc3W+QUk+mCNq1adjSAYPowC0NDthXb15WvoNMoaFC0PvI2UgxPzC
Zbp/PrHwJXh24SWLGgrPA3Aj8DuzDqHEpLr4EdJ9xgJtOVm/IOYcTvQbM47601EwiL/BZa8F+S1f
LR+x/B1e7AstTnAe8PlVyGIUqdMfGB0Xy7VhnDqtuqhJCND3CRC9lSwv7yg7n6xDH6SCCYsPlbjR
H83ONb6QksP6g0eBnBMHsdYqkco9ARD/3z560yPmXXPiJYPaNmhx7vp5WMsFG19dzJQ2Ba6HJJ4T
Rb/N+nivqWAsy0IUhsQfs//9hGhYrmmJFR1u7UsnEfFGufTqm4+J/V4jBJJrwHwpEw6kZ2S2ZeNw
KhZVkjYFiMbDeVev/t9LUe0wGLCYnzXBen27FlynzFUmk+qnlKyIsZXb2MrKtmXaYgB48nKCh/ay
MWJwaj00vqYaBlrzk4nbCcIf05w0QvzU4tbnAZ7Eup7eHLIXAjLg+Y3xpnTUNdCy4J5wmYHLlJg7
RhZuWcs3Z3hZvZYFjAC/DEQ69dd2OQ2T98zOFAqLBAwEzlLFye94iyUJRzgaOKbJQQ17FUlYQZUB
1iIMG5f9GPwAE+D4CvOTSulW64PxgoBs2HW0OpMEDTRfjB0SYdZbdFeOE1D8MXMD8/ffI8gpzmht
p1kuIVCLHwq1enuQNE2MOlgyEcx/eeplrX+JoGNNBDnBqI8k4+fWFIUwOsKAMILePSK7t0D9dhYl
cip6+7tQyq/x2hAr7wbVaXF61l3xAoxlAh+N/HfepGS9HXTiudL4ozyMioU//hoYnxRLf/GizQ/1
CzyBfI4HGvN2eV8EDdAjUF12mioB0A1XDwQLZOp/QeYMtWy4oUcEONZRNi8IgpYOoorzVBK9PqOc
WXnDr9tLHadSflLAGt0ZEq5Enx6Wgl4jrTyuIToiPFRasJkisUDMPAgM06nlVPMv+OlG88Xbu/n5
nGzqNcpIrwKe/HGmPzMA4C5ZhC7X0b81bCa/1PMAzPE3bWqVWfAhbgOu4dO4QwcxiiwS7rmKsxUj
3ilS1aGggmyFmlSWcoP+Zo0I07Buibe0X0P4OtJtEuyoYBsmYtEQbPPY899L/NnEH2UbC3mFS9B7
hFilglB6ZeyThl/IK5BvGniRkw+15vMibIkrtYoyT4qATMm9k2Xt4YYQ2C92TIJUUnXo3WfrArmW
odI3wpUOKcPve+SDl3eMGCnw5zzzWTjrk+vZ6V6QAIsPEliHRN3SZ3Bkppcwz8xS/JUXUsKWTBOC
vcPcDkW1mx8DxVCNBQ6j0Khf4KMnjg9GIasCMq9R/Pg7pFFEItTMlC71ATH9mG5up0mQm10HIs/y
EI08e5BMs9h57dqOOCgNlVa+7IME28mdO+AlnJzl1+iWsoUCGtS4sVjquO7vh1dwngmTl1MkUIln
gSEEi+A8qIxzaFEvajEbbiUnimy/wek8/zEhdcXvR/BiV2uTWrMwgrcywifvAj5Eotr8hpd9Hqbx
YDYJng5U1IqJM+ycrYTsKNQtIRWH9mg+jX4/Il93768cNWCvg1X0SkUmKWyoqwxWnTFDMP5l1iPB
fBTBCrb/JcGl2cbRy/MBv8M8aAOpGpOSbab1xHbXuUSDuApnEJacFFC3zyfO6aIxgzSPcpcX2reb
NCiMQoNwMvHXvDP6PkK9b1M5YXfiAXOT/MjU4cFRTMYypaGwxsmvh+I2HZu3iDuFDZbjMZG/VuhC
dnE47ct/LnV+NDuSMTNaJio4lZXuOjXcxb0s13vKRxlIaFerHqVinrz6V9CBHBgXNaUHZqqVctsP
Qh+sKXq6faDwWeoL67BS3kT2ZV1iDNJOgAiEOiZk548NNUs8tVOopQamhmHrlMQ3Y8WklGeNiUp5
8Uhgv0p7VVUewtyYsx/xPB4xJL0Xp6jIZ/LWYruk64ztaUI3KrIyQTsDLoh/EvtxiT/oTQFyDhc0
5YxoGAVntWlVrb5IxQXhWZsMpfln0igzP4ErlY38UNrdNpzQKVCNkaYPnA5GEAsmErL/Oa1eI4N3
spz+AZJW/OyTzbFPujFVWS5d+QixlucnLlYDsGWrNOIDgvvjQEAPS2t+f5xbI7fgIfVohnogOqXS
4GjpBhCc2E+NaDPlnrlJ3nNs1beQYNZkf8LJL2+A80l3e+mFRIen0LBIW5y8IJWwdycN18ur1ZSv
lEykGKYNrKv8Q3v9eVHkA8osL4G6MiChhvi7ah5E+af4gu+VbvEwFf4ZPO9Yd8WDiXnGTGpELAjK
LagNQCepiw7kKw3IjXBhfDOJqWjho++C/3MRV7y5CMK4vSqJ1u3hFSvoDCpFF6bVJiTi6oag33Tg
r58nu2FBAeN0daI7rdcNBNvhbQ9eaGOa4VYyGZ02Ctu5G8b7Ge4x0+qTI1XiOi0DYz2snBy2U6+/
0k2fPSXmKLYxjJPuovZDAy4w5C8AoNbyDYcEHMN7zKSZJUUFeTSh8GDI7s3XafwqSDHdaajIiwFY
ezyleYY0/dLTHuL+JNEWraVwNMhg+JMoRBZW6W9TRp7b4TqMDdsBfUwdyV64GZhRpd7RiBclOt0v
WewiwaqfNoWdEQVTF6sGJrzXHXSCaBtP4PpZqvuE2FWE/6zUZqDH38Opbq34EbyFXZWsy+Kosn1Q
wuRkJhs5Sc5cDoOEIQgyxVNmBP0tCBsh7uWVkNLmjk/vSxzwchKt5B23SkCcB1xklXiE/RNyucd8
oP0/z2vUhTaXG7SvZAqUz7uPHXk79bPR2tNC83aw1O0W7zBkh9c5AmrTnd3zGmAOnew/dEIdTaxp
DttUwmDiV0zHumhfBGm9BtjXzBkrlg5o2DC5T55IxbGVFM0Hs68ImSISJ9AiJ8etlim4uc4qJmCI
pYOw+IBkvYv+WhBRjpQdofpswqLMC7W9UP2JEw1hPDtMbjdXo1qpHj8SvziCqT79JORpAXdpOR0W
3dZgNcoLcrMx8zVFRPhzh5UTNPozFWD3OMW6E8hcw2MQ1vzBiEQZ6/wX89DHNlYxj7h8KT0OU39w
2wFjVNy2eB0Y4GiiXvjN+hByoBN7ikKWjnktwAzU8F5bgtPoLvWfzQCPTVhC+iQ3alGgE7cv1MXT
8Td1YHbbu7CILdSlwCwtapARO49Vdo1CbKUS+VJc9Pg7crw/hGyz33bg8es+pSIecQqKkGDTeURj
CfuJIqMyU56rLbfc2+pwmtpoVwohgogigspgbmUjiAyyq5YwfVPx+bkeGlpaVq8vuQI9/KcYk+9a
LJX+X4HtG8MPajeq/ENk8/8U2VoffoRjappIALM/xdCv16loWGV/NDomaWjM4pTtlAWZLqpm/7P8
mW+QY3G6QfpA2ubLv9Y1tMGR0xfNO84e7Kd95joGDaEXS3yoif8VjEzG9TW+eqOCtlYconlnlYx/
jKM9k1/Nzx7R9WiySYyjV0TrTkwPy1K9HGGddwyFvk/ycVOPCOliiIVzoVQx+9r7EKql3dEg0VDa
Tav4TGU7Pz3vhdD6IY51/EKOLXfcG5nf0q+rNEUIZZZLsQAbr53/PHBeP0VP3vsd9VFu4bg/231+
02K9Ye3aJmT5ilWpaJxpkMatJhTX8fRjZkeUrf5cT1su4ytzOXZXADZBHC9TlUV33Ut5wooIExii
HD2EhOzLv4dPrDAUMTHoobqOqeM3hF51akQSq/DsxHhHlciBtkCKLlTTPAIWTMc0AZ+caiE/dL2I
OcoRm9my376xktHxju0zEXqiWOkF+fqg1v181pjUn6MIHZJft2BSJFaK4Qepd1jrkHRR8tU7adZM
hqwk0ka207AAMvA9EccijjEKO+k5Ts//cpiB222/pC754m4eyIVJaWNHzkH+oEoTOX2sBeooEaKf
LQHrqOiLuPm0zLR5m2n1gV3BZX1e3QOF4aXDReAz+hgUqqIXVud54gTQfyE1VlgtC2I2fKK0KBVr
a07A5Fzl0dTJn1+WIHBPOblj9ijxHpBuRh0RUJHNF6JzNe7vU+d6/wm4FbX1PU3w7ij1813d/6PF
QbGj6JLY0oqMN7XI4hHTUuQ7uaCRjaOtn3JIAQP0/avXbzEAEPnLEzMGB8wEaAq3VY1WaYA4OXmn
ERonvYMG5dFk9iBlvvhHlsa8agayqmIGamQ4+v03EQy+de82PkgICLipqjWBlcMDYY6/UlHJ6Tsi
88xvxOOK5ptNZIwbP8jlrfnf7xUU/p1cmiaX7runESPJts47N/sQk0ck5aVtaU6E+h9A8ogZ5LZb
BC+c71IAUkC9MEmj9zAdegnHWWeJk3Wz7E9BEgp6DXgl6tq7rDqp9EO5D8yKK3fjAVhdCyaoCT4o
W4xMjTeRjlAYbfh/SkqJbRk31hLqedPti9b73T06DZfGrq6XgFhS6YAk59yiT18JZ7ZuQei9Bn69
S3kYQbEaJUdOt2lmsf56frLAfQxa7kS0thL7hilTzyEugkKOOCSgzd/PSXBzRFLJCqJz982tk/+W
RU4wg0jUroXMoKda5m843rhPxqQCNgdCThTkxlIcWG1xXyTlEt0SNzE0ZRGDMxLYDvSSzNDy4gYw
RE0mJKhJP6ZtshsdKnoR4Sg0ht1Gb34menAf+5ZmQCDUsJJ97M9XrGGnEss3Wwcsg95h3gBjTbaX
5+XwX7d6jVD06fREPmW9u+DDuKRbCqn/3ngSqj+EC8NjGMrvjUlNpd8ea+wUrH680XRhnD5lh8Eh
e3OB7/Us+ym+u4dA9bwsZMBitVug1TAoTlsTugh0W6AGGEDXBH3/6I1RATGXYAZo2Nd8+TR0vYNA
BmDDwvcPI8sdSYmHSVZn7nHXMYGoWeyWgxZh/Mq8vD9WkJL96CaZ4zHu5mjnNnua/JWgvWmcB+Y7
lPTtysQNTUk3TJiI2xOFwH09eSGpAjFz4y8fcoU9TkCLqImYtfElhhqrhcTc+Eoc2o2EMU4gsd7Q
1FEAqImbmTBYz11P829NisFaSfVQhiZLi1Eg2DbEB+z3ogECUQ5e91j3qXMxuFQoIHEqixaDKPXV
qGOUYRXtKpuxR8m7LxE/VxWqae713HExGtiday3Gq6QiU5t2mvBEs3NfH3PS+RNwciLpUB4Luc8k
owobyaM6Wt069X5TxY++FeEdLjONKR9d6p9gpIHx0pE+HJrI+2Kf6pXUKq94mHrw1UZWRjoxqRnT
4Jn31mcmIMHu2ob6hpy1EfEwx3EO7omOvMp1fas/fyS1Vz7PY5c+3vn00hHot+AfDzheYC+l1BCO
5iO+hmoHHklQbeVzpJl6u6gpdDw/xUJ+eoX5Nh6NjwHym8k6twwFrbmwcDdc6ItRMzJQeH7j+euE
p48aT3lD0U+rmvTPHaEPTIueGBIFkZzxxFdyIxoyWyIWpZ2QbWSWU5klXlhV26p37Wj7akOvGy26
GIJmng+MVBNt5RFvqJb7gdNK5OSnY1N6cTON0nUA5gSD45Wn8LNqw5nfOoRizvVeKKzG6VOY1sQc
rbh3u/wMjVKQnvZ84U0NmTPrwBFeviU76FbTXOjjWVdWPr2e+ZbOdng/jvmecfHT9k1LMzXlp+pJ
0KOu8dkhWnx0akzGOWktuZwhX5L1npJr+OACRMUCAgVOnf374h6DXaSi1s/arTsjTz4ho+TCSC+Y
RpHtMjlWkiiUMZWOh5o9xIwFQ2rCDskkYv6GFmrY+GpJ4wsbtKCvNJG5g2seeWUA1xBr/gaNqC0T
9uSf9on8Hh164Hi22ahl+zYm3NmVYCeEAOiR4tAeEhijVliEKX5277mito6G+JH+SiCuLlVQaX23
RoguydtCVfsBcwL2ursi9SWCgo/Pr8ceflqao/Tdd2e7HB0IeZ7Nkdsi5NuOdaa86TBo+ui9oIAr
xtcluoOuvkazD8MF4p4hlaa1LVEKRAvFnW658waeZvGYKark5kvSDmoVV1JI13/Hk6CnP101QOuf
kE0R7REbFsGb9SLcumnFh8cfBlhB041Y9VTpUhq6eEA4wv2Eq6UNzoWao1UwDMoO+tQ/7PnueAL6
nuvzx4GbvT+UJy0gcy8QUBdeCjLESMQRDWBYn9rf+ZS54Ee86DsHoOVCBVlJfAcUzGhU4qBgEUbj
Bs5ko+u7oWz7E4e68MZrGDeVBhn5pTzEKraPf4BnqFZRuA0Q5zoC0MxpNVExafIgkkSynSvUGwpH
XxX5qy3CQy5hdu5zS7CPInV688NLza4M1FqT14d3fItYZST9ah5+HV8TRemTEX0nxVrKslgu5Od3
EH2SEYIAiGW5w9M9TUNzFp98cpAYQbzejC660JJ5GbfclbaiulZIOpYsZnbHvGRWkgV0p7UmSb18
adD6j8ccT3JaVYf6dA6V0EBAul0wZ+OKeLY6xxPyXWCpkZ4a0NrTU5edSs1dMZjI+fBzRn/KkYtm
GHoTD7x+6pMwmtHQMnmCTJMqkMa4DU2IowUK02X8o9NUdjCylbgFThcwxoraQrRDmw5YZDL/xnDL
uFH4kmmJ55Uoys2Lw86Uhmsao1DCMttC6moTu/beFSs3sffNOoEo65+85k4JohQaubZ9XE6YUl9E
NReZTc7xVHf/93QTJFKpkEmv7rbvju2V/+HrAhh2MbYe2tpRmYZSmVEOCpywRu7VKNaJtHu+Z1lZ
SbZeTbhRS3VdeEJsYDY4CPa7eA1n7Dri3kUY5i/KMYECq55ut9yeKOi65s8NzENK4tyPvqflsjSU
+3GsRRX3B9gIBTc2GwU2dLk6cMdgHa9Q0R8+32IRWe6HhVhhEm/9VkHNZc9qZ3h4gIlaaERvLKrO
8NRD5VT+FF5kz01RUqImKqjvurvcg/lq08gOhMzF2GN4a3LsPvVnvThdp91pwuEERw8vECs+5ecZ
jesTHgyGYnShdhAWKXL9+WyXKwZQBpmCLMn6NN7zVS1DZF8oaL5/lIKlvGtyabfIVUcM9OOM1SxA
9qxbTn4zjkv02YftDNWLPFx6oft/G1ys/B5dLuf3sK3gOeLPglVyCuguPVFkBzaLbp01+tWgMf3y
c0uyzezeVOW5aSp8TvfrwxFEUyvy7XEVOI6wzNiCORRFedHHCIS327piNVYry2MWNNeraCKBYhAR
ReUqZ9k17xieJ0U1Uc9Jta7kuW7DddxrebM52y9H3jzyW09JWee36SVpST70nzQDNC9+bdENq77g
+KlAgb1ZLS2BvByhQ9FPdMCdsfFWkZ3rOrHzMK+OfdAlt23PQrife7fEGVtiVNErfCXSKOVaSNnu
APVljetzJcQig8eYFsIWJ/t4jpGaeYda+9h3mxVx/u2KI2ol+zAXwPyQc4UDK197mPe1Juc9btzd
xSxn8qRz9teMLXAHoiSMvQ6QrT+kyZLuS1Oc3SGzdFCpBroclfOFfhpYn9MxAINfrFukpHXt6fO+
kOYjFYStQsZOtJ0dsD4USiBFZ9/1bntaJXMN/LyzZBiuJzpi0seLIxHoyqS3rcd3YMJUzlyTjNUi
Tde39xLoI/1YgxJS08OO73RqbVdZtI2G9EE8koZnfmm9MYvQeLUBeCljQXprZd8/KWjUvMc6rFm7
hhvTq3UBaPxdmXMR67tb9XYnmEv8YHhpsv+LCXRVbCC3GvMCqW+K/ExbIZeR14prRMxk9jTzmWqh
cat1vd5nNfDDYGnmfCuJ4Cqn6Zsuq1GBNNX1P92+3ALMxIEV/75tNOWE85qrnFj1SqCSgDmEZD45
kObNNshJSuspJXwBVboIjXaylAysSL7MlC+TJMlaz+r1oiFSFci9y6XvV+/2E0/eltjQFRrDAWjm
A+Y8q0ZLvXlCm7HR+QPnwJ4zVNTgQr0vrsFAYuFA6dY1EUcTwOOIjKJm/3ghQ0Z2cqJtr1fKl8lv
MXBC6uHCSaQJlBTHeQmGht6UobOiH63zPaOFJoRD6Fl3unNECZOzgZ0r+2Ciup2/t5SVOMkK6KfP
MahfhYFvham21YiAMQSv2LWW2Cx+knb/j4ogFH5pAgCe8YcAZv8brqFvHS3H5vyoQ87qUe2wMDa/
ZmmEaPK3JPYQl+nKqSJfMHOE9kLjQp7DIf7U8EWYV6WBBLvR86FQsXFOWyaFkFQL2aFJ6ApPGggP
2M/qxdkkeBi7Nru2UC9CEYSPtwTM/cPXrBhwgFDgL9tEoG7cBlHu3c+ZjsgIurMgEJi54NX4vkZf
+zawfpsN4Ebt141LmQWRJrEogUwiTlAo4S2jajCzd/kTRcElglB08Q8in/4A2QLA+73eyoCRxP5v
E4Z3UiovAwUr2TcSz0w8D/ZyPd0rlGBqQG734b9K/nwkTLKRdsFStE5VOFmUsCYmNJqwJWqXSy+z
NK6l5D02rWkukV4qnVLv0TwuHLQwBMkBbtF6P+huojUQVvSXIvhgLsIg3TWUSnUc22RjDJ0Jkp0i
VYAPjVNSRMLOlTWxNUAq8vrEDd9NdPN5O1ZWlZXnoZpGT0LvRu2XmsZ6PDpxZgjYGwedOKcx9+l3
6TiW98RNRyptakb57Je/M0fhCllCxWqMBD1GNgCRtRi7FmwzjDNx7ObNwgS9GsgDLj9Dksr8ELH7
Fx0K7fMkKTaGjGaQQ1c79AYZL/J4qO/YHW/9YquJGwW8MdWdD7LLCVC4GhC5ppmojnnq9OVj1Gih
pj9oRMTcKwKA6Q==
`protect end_protected

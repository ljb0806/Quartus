��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB��n͖����:����E�w�mLH�Qҭ�b����.b4��ǄC����~�83W>��n7��̌Ḗ�*$��c��hl!�CO�����wPq���cs�|�"�;����+���)U��&��?�;��*�\0�Tȡ�""j�0�7����͋�k�p�g�l���ї�s\���p�� �f�{�>�MfAF�C�/���i`��}p՛䑶4:�\�,>P{7��/��)�J���&�P�(���I�o�����ٙ��ί%��чj���j�H�CZ]�C�qҬc��Б��@���Pj�5A.�x̱r|��I�^�67"�+��c��Ȫ/��5���_�Fr����`���� +jB:0�5��l�Q���l�r������gtf�6�Eՠ�Zid�+�O��~��g:^-D��	�/2-$i[�c��v|A�)�*�V!��?��ʱ/Ey����@�s��r��M�9}Ǥ�b�_D�pɅo�(k����t.6 1�*(;��i����j��^�ezG��*���k����a۾���e���������#g�8���j<֏�:��ȠWn[]�Ů�e$��>�(e��]K[Z��j��4X�oLY�s����b���
@3���q�q�����fVj�=���b&T\�N��=e*#��R����
r7�r$�*�x����ƾud��"��q˽�U�Ob���}��Dճ�
�������C�|J�^y/��鐴��DA�WaP��}7� � ���i峾�!&����˖�+?*�7+��hw&T��.{�oeS
1�[�ec��%$#�fd)$a����Kn����kFgQ�W� '$?yi��#�� l�nl,��>-85"�L)�hy�xa\yØL_n+���Y�O1�9y��9�{��˦=���>��j����l`:7����Ks���֔�r����豂ݑ�m�	��b�+olh`�"`���$WjKD�aas��ʥ�
��8��BG/�cY�c?���]ӛ�V6�G�l�-�C��m"n\k�!fE�P�>�Xym���ҹ�iL��/�G ���Q?�b ���m��yb�b���7���Uf�!�6$�ښ��|���5�h�ꤙ����T[�S�	ow��k��p�j�o�TU�m�`C�қ�^��M��<�� #�y���u@�%�7�l���fkH�~�/�/��6���p�/�7"j`e&m�E����[9h-B��bXNИ1#e%8&l�V1<�|9?��k���j()��.�Q{w$�c��$����ˬp�u� �3-!j����j�G�xbs}*%i��0������	hs6�1N2=���������(���U��;�Sac-�s�!OX%�}E�9�-&N׍��k700Ics�Yjմ�=�9�6���l����a,b��0�N0g���}�K��h�m�,*l�'������	�A³���pIg�e��P�����++V�b���y��Z� ���B�v�w��d ښ�IVnV�p���4 �%�t;���Z���CJ�����=�|�bǕ}:�*��-S�ҽY�ɏK�7jP���.G�aQ�lv):�T����=r�%���P���¦Y.�_��^`��0�PgZƲԒ~D��6�̦��l4Y��ϕ+V�Z���W�aŠ�1yA�P�9i�
Y#�o���=���N�I�oj�Qe�FdPL�O��ami�g�)2V�A����5��O�aJ���с��(�
��ț�Y��S�-ʿ�:���eK�1�H���H���ֿȱ��R}���ܔ�{ ��a-$X�>���iHH���>�Fʄ��%�����٣c�YTwchTr
�j�%b�`��w�CƗ�i����Z6.�e��?@e"w�K^˛y�9�~��$e���6mgp׽�����2FqpqJ/���M��FkQ�a�5Fg���	{�pe�`!�}���C���Hz]~��,W�$4rjeH�YX͖��`f0�#,����B��g�GkW�V~\tYq)��s-#���$�o�ɤ�;��L,���;�I�}2���<U���0�I�9�(6���qqqu1-8�.���P�F��X�e?N�8G�h|�����Ū����䷑�H:}j�����{ǃySٻ�s{0jv���hؐ����ºǳn�f�6�b��P��� ��G����n��l8�`%$3K����/�v?.@q�Kd��p�M�PaI�h�??�2��9@���7�/Ѣh���(hh5v�'�1���g����\��%S��"���a�mO_rdY��K�8��w:���ɯ�.s�<�E��VȊ�y8zq�$aH���4��_v� ��)o"�Dh�ZN����k��\:#ŭ�Wc�&ѝMm�����h��OF�^�	���1�,��Me�-���0,�P0;H�@сr
x(+��.�e�����,E˭�hN�ӄ1g2��C��Dz�)�cA>:d��1L�u=�5[/vU[#��k'��;��ﭘ���28�8��x�mIp����̘��_�L�r����̯Q�ְ%�zvac�]RCAƷGi�2?�x4E(d~;pw�+z�X�D(��l�oڋ����[���>�d^�QO�u�u�~��Q{���U����Ǆg�-�3Ӝ��yu9l�R,~�R������:����
��)�<$?�7�Pb�P(Ք�=ol�����[mf/|(ĥ�38�G�'����E�������>��G%�(]m��c�]��k9QS��Q�͌a�N�������P'�Rg�A?Z@W;
�����q�y���XҤ{����n���=�Q��q߂���X�ݺ��OD!չ�Z�>�o��)�1͗�3���&�#`�8�D�r��2����'��K�_��,eq#���T�γm�}��S)���A{�b+ҡ5 #��ݎ���=X�ϐ���&�Kj���Ɠh�6�
�9蜻������H��f��GO�ۖ�+��:o�S#��RO��&nP��d��܃�C��������F����4��m��Y�K� ���/��K�9	
Odo��`��O��o(T8E�&�s��*"�hQwUp�WJ7�Rh��_�Pi$$
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sQNPBhZRH1Gpp05/zlNWnIhDOsYGNty4pRyXS40Brm4PKCpK0xGf9qW4Z0AvWJ2rC+Z4Qi5IT3m8
4HtwoD6t10NGXh3ZYhn10ogfzogdQmFettzoHcpwYhk7iG2iUtgFxdaS6r8iq4wCvrKS/2oLw7yn
Z6CtK2G1A1lkuQYnud75aX7aToiEQqyywLzWNM5diFavKDDFIiZr/lelWrzaDMvzc1AdyQanLiZv
YOgE57JLJfPBUVSHZq2LgH2YE4GkRH2+c1OkHIzc1zT+RVerr7bGCDY5d9dS0+U4cD/drebZ5a3E
448L6+XWAl5dDJFYpfV50DtLfE5LrMPvTzGCyA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47136)
`protect data_block
yoK6+9/JNVIjjia03WH07Mty1VCiENEigKe+91xgdk2S2tU1lsfj5ZOs8G5JZugZ7KyXIVOq+F2j
+9OjySVKxOqlLvGmSUM/j65/StgJMYF9uJY4SOkHi0wE5d+0X+TO0GatJqINhCDi+tyYKbzI5rem
F+Uh36B+PESV7VL5/JTvDT5xroXrdRYDCMx7RhfY1aidGCZ9U4KnObyZe1b5CaAbdEn7A0NdDZSM
7sPszRFxXTGlwKavn5CgEDZUqPPPfBRQAf343rI2x5sgntgbrIXE5jWNOY5K6wy7Oh32EF4hrVzk
MBjcEn0FBy/mrK5ku+Aj0FFVLwTBdna65y4WxrOpJqcIuxHbRrkvrYE4UwW06bh3ymHg3OzXlvci
Ni1ikTaG+pjlgolG49M77mCVJteU3wMNPBIh/I4x7HBIMAiHU51tTUDF107g7C5y3741qkRkbLSR
toY2BahqMJG94EnpwfbpQ+wRx0GMWy0bbt15tEoodJFybPkCc/pR3R74Sy2jekTEN9Fdx2Zv1H9U
K8piMpM8wyERcZrjVDSRoW2GwG7GPQzyRkZIcxy5qkzxiph77QR8mBXgtM2pWliNm10qdyOztx46
9d8etpfrgSnqe4ARzRaGmfW1wYFTzACReArhge0GD66TYSqsCo5Ynts5Ix9ElqOOBmmTkM/CBO2e
6hXEsRRIiymWY/vgS7DvJx3WkD+2vajfvsYoTiDiQnwVb/tUZE2MdSP9fRwVcdohBBiYkQnEN45J
fXDr+7ZWMo5e2ZO1pdUejUKngOpsTB7wvP+Tfkr5dY4WrX5d6AuwAiGTOpHP/PSXcSmXomdBAqq7
Xgiabv60lM/46n1dUtctOK6vMB4Yipe1JTT+jMEUFRK52oig4cEUpzZ1WihlkeqWwXL1LstGFOMf
0+zUJ/1UVeoW9BU1Wp0TsVcJDc2tVmKGskHt0B/9JLkgTnqvOpGNLoFTrnRQuDjtgp343UdJPRNj
OjsAdzeNkolrs/g3U/NukK1J/HzOBFZVOo7s4J+XWvdaxQtsiwWqgOkwvaWHTu7TuF6jDQAcn/0F
/5pYU6p2RqEztEegSztnvcuykkmadbEVXSatLxXf1S+S+2NiB7XTTX/C60xmmHMhmmkG1ZAocs+r
MpEV17UU7jPORo9GWwcQqC+rVMhBuWEMN1F3DPSAR9KuSQulXppPd1dVzbTjK9PmagWYUPo88Rvi
EBwa5+8o48kkKS1Fb30vnKM+GJFYi19szm0XdKPR7F/NJxliA08/h22GItQ0JcZVEwicCfun1zDw
cbpZjuGKdR/CncasOGPcYEcuQ4QuSwlP81ZLTTdSBMzYytbP+1vu7hmuzkvWo21PypKn7Ot7Ua6t
HAG8MB3m4sDMVjVhVmKJrvE+NLGxmFlyYsPW5kOSZE3xrkeBAhwmtKa4jSnGpsPVS4tAdR8nysba
5mUiJn9oJv7BVQOCh3xST++ReC7Dd2FbvaBp+sz3VG3dxn9ReikE+xvNsuim341VYOGCz6DfUzPe
jYcSk06+6jsVuIIEJvTiRqc7uWOUclUBr2kGSkqTTLKKr70xqbnP+KJT0kvznDd91HnxSsyKwpTC
BuF7oQ5pb1SA8wDto41+JtKeTsrmS/bPTNhGZwxFXHUQUVubEfRQO37iaA/HaBnDdWZpUSiBcht3
4gjoNPxj/mkvy7mnHhg0HrWhtErKwv3/j57Mr0TfZQrun66m8A45Dv1iTlfc5E41FlLGl8OTAc5P
QpTqO+jTURTNcalpogfYHTe6HnkgwdeYW+sqTL+MD+V0YUqFCS5VZAPlqox9PXB6wqfHKCKm+wu+
VeT27+kDTCFWn+ef0chXjggkg5VKFKQBni/Rp6RcsT4BEFxeUrn2u5ZoFh+FCYBx4yEO0S8lg447
uI75uDT1ecD1Fs/fOGn+e9osMbMll68hnrjFSJQjIC4oCINA/ybIkQlw93zicOXtr51aMHRvGZXM
xEYc2Z+JrxbjmMO/rkOi5vNs9eeyGH286Gj26nq8fIpYJaQI+gZcdpmqe6m5MiIL7k14IIzOzKUY
y5aTI52cQmDePZ+taoq3CxW0NTMoqXacJ0xB50o11hslJWEi0wpbgfwXyeMKcOdMsCHT3oisuoh4
G485yUw/9C9aIatpI0/GG6t0nW69/EE1eTgBiArJheswMZ0R7R0lssdX95x6FIOr6WW5w8FkveV7
O/XEIqAcpPm2s+64CtfrcL1YRyL4vIJq4XU1uwgSJtGwXXZDhgj+d+o079HZmc5RSHjTVo22naqH
sAgj7k+jHzv4kZXapehVnBmFtD7y1jaCOtl3SI9iXfrapTf4ESczdrMCJDYohw5ppXB/EhyZGyAc
BJqmo5EjIpClCUqJ2p86fLdEeJdX90rPFiH3LaEeA7Ux2D+bJzUK295Dx3M1a591lFxCPKuXx5SH
UxMQoAkkZtt5MWDPk8xJCiL99bJ3WLaguOZq2sEh0Qu/J6e87e9puFUM+3p7/1V9/amFzlEdAjsm
MaPOWT5tY877Ic/c4CTkFABT/QCfE0YfGrSmbVQBzd8WC9aP3bECQkKBnK4zDE81FJDLmO+FyWSq
x2QODmZYNwTVfwIIL3EFOn14TLQX0mLQVng8Q30ONOIYrsMwTYAGKgBm4sNAcKowqpcqpzgjlNuw
e8NPQrMOHudS70X4VF73Yj+NFzI8zrIsRnz7h35PEXk6dCC59ZhwHrk6QTg0il8AN8XrADamfC8m
G7+bVpeMjlSvZqT5oUgwnEXiC8KVAS8lMfbl5Ygo93MQg3+2SwPS/7+YW3tNL8sXR9yClpFyAx4j
VehmghEE2lOUT1NCjR1TxwNAnsd/Kj+90Uh8xSMCpafpk0LlVTTtkppUPMSE16ImWLWTXNI7iGnF
AXJJIAGGJEbQKZ5DD/yBkgVKiVHxa07R5A4tkczbBDQdm7ziQMc8J5+4IXo1n7Mk1O0DW9HBziYL
/ow+G68AHp8xdv3GunHyIOcoHp/YbaX9jJlsLrRpUgur0jJ3PxE6ZO856TYjJ4wkhcY9VjwIwNeE
AIT2GKCg0mgepGym8o8FuQyUtKSYj5f0B9Lnl731HQiqEGv9zbxfthoQ+ge/Y/lhzFNtpgAjKID+
wAAz1vcWo1J82M2yCWoyz0y3rnqnoUTL9qZZztUV7G/mZE3wq/cvPcc5iMyY1CfeEXI2FEUHTMeo
B2qb5kXy8ygjfUty88vOv9z0hTLD3vjJ+VAZFavP+2mdW6HFIdb7w1g7y3pNkwo+OPYNNuRvYO1m
R90LsCLbI1qEyOtD/Gp60WfXS6dAUlOZML724fTcSmp2o/NpTnOwryTOwNb/F3WiSfYHYbjqwV+o
FzN+ad4z7pjE+tqkLPrdSIT4CI2ACGsqJxhXf1PEgaTrOvPWIi6+KthLoUJzHC2il6vzfVfhMmFw
4ptXnNu7QjRJGRSZZSyOkpXZc9vN5qHK1O151TLJRoicFJiUGMO9qmbO+Qqye9R9BJPrEd6OD2aR
Y+H8SiwzKRUhCXk4/STP16s+6cC92iq6RNwKsR5VKTzJKe8cQdye8Fvpa4It/+dwrfOv7/lOCwnP
JKyR7TxT8wPR6/IJ0azrH5D+ZKxNbhkj34eAmlcXf65Z/JJ0Xs9BGqb4Xelld/HPaeCUrxAWHdsI
oNmNVlV/g6U13+22tc2D1fFUbhOJbSIxva/hDCkEfC5D7PCsAHJIgZMY+Id+xDwTwq8B83oHJEeA
lA42+UqLiZ8ZS4dUm0NYxUqlQMOvMSlezd4IZehJGOiUo/o1C4lqVvy2OiNa8e2zVqIuzKzL7drv
gmYgADeuSgXSh5bufKXLCIPKO1mtbd5xf4UZDSTbYjE3WrRdJ1HwREMu3pSTBigzNltuAZJ/pQG3
MlMA+KbV53G/BNfOufKzYwV5e8g7o+a5y/aEBKiJc7HsCohbLFeWL7mLrebnffHL4vRk+/JYeq9c
47Sh9WuHsW6ConFK2kerXxjksu3o6woapF1Ou4r97WiEFW+8Vr+3WND+5vyUIZfDIvjXcZN3aQp7
+GQf2c5JkFI/oA8yGz2EkRdCiupDoi0ZRKzWC9t4O3ORCIExLRZGquxv18FZNtXHUuB/UKYqSu1Y
Rhp+1R0JhX9WOH4o3I3HQGV0J/J1ShE7HXSc/cHXgp8JNHSrM0SHU7sY6IZKiprYBguho8QaHv07
zhhEW+xX/2+RRtnWmFutSBJtc9A8N4GTSqFJAvlU0EY/Jw4v0IpzzPlbc8LP3uISAyV9TWiajkXP
K7SCIYwIs72sAs9dLUedutxPozRlrHVa0BZMAye5sgDReMlh4XPG6oavHN56+qtvJ6qS7cOLbVf6
HaX93DDKbxPVf/kA4S16nBr1mB+Tjx8Dx/RbnmiLapEk6M/QMdrVWRzT5rQB6CYrboyo6opwOSfV
C4h9suCCHeYTc8PYZzMLy5WQdTWuuRRcGtynfBXtfzi/XwUZ9Tr0NgBbX3rHQPJqttbt737fLt5a
yxorHiC0N+Uoojgpf1mb5ULqRjgFdVNT838wReN4mVpXmMRtLIpGozl2BgBoosPvVtSNlq4+DGGB
wtGv5kV+R70hPeme9UjCwbUpk1iW5lW+XC7vpFvHw4jnmPkCeKW9YU+6aLpg0DsGNq6+pc2rcZm+
EoFiYq5hA0Qjxf/WsSqUwRNMuP8l6IMOMZ8AdZRlBnR7kCrw74THm9YYnUtpyTD0LryicZgvS/cT
YBD1JzohxXS6yD15z6aT4uGrFsne+Dx4rqb5+k2pYkxImNcVl1XFQ7X6dyUizJ5ydBAWGJdMgscJ
FfwHvj55ZpnubLGqIsbS8E+tS7zlbwSxpJy0kmPODJR+oMr/iSA2PnR7bM7fuLakGWDmqn4y3pwt
2z1hFZbqFV9iZdwLtpV0c280Hbex52GWHUMxDZcLBtAnYDITYGgk75bFRs3H7M5Tk/mGsL7Ad/Zf
B8G4zZTLjHQPeAFwQkmygPjMPRQoVE/TwAQB5CfHGU2KdIVMSUq14xKHfOOBEERvPP21MdZK7iB8
TB68LhJkLmhKRXkJ+UcCqo8YIUVgBnHUXwXfyArXWSYmB1fLPCmu+kTZxmwKti7kChTRH+kLQMbt
+OXm+mwnmZ+LupETlDIyESKrgy85tVb4hQg+RLyhsVdmunIMqNHo3Dkf0FqSUdNur7FQy1FlLnau
ik3Jv+wFHsxIyzenj4162m1tpfxGzjza7/BTS/LDIfDPfiO+CpWS3iJcw64k+udQY5jnB9QjDJ4X
Aw16tl5NUjebo4YsjNlq3/pCDuKDfO12VTRkoZJY1ZQOLyYXY9k3dQo3dOUiJx91Mvim65MVkce9
gnh7XSl5ISkkHMI8DHEDiu0aD0b1FOVTIIH+vyKSTuwsh8+03+1QyB17nzGhyvB8sAmvAjHhMJSb
FZNGvcPCWIexWWDyU3yzZqaQYHvHMuGDD2nvynDCxaTjI2Z7ArsTNJmM5iwDWFe+S4Y6PJVGfLxk
C0rv15SAUv3Tlpmd+fz4i+J4gO7FbJyG7X9AHNrqYIvc/J3YH0mWSPnuras7WlvQ8LCI/dhL0OuY
OAqgDyirJDqDL1jKbwWCtaR/8bTPXLgdiCBiNhICLb6G3bWKTiIArv2RPr+sKBgXrTICwUvsmavr
fdCLDl3Fio+T5OmPkjEVvDJ8k0+UmBWkGdCrBBErlEKPCZ/wNsyvikGvuFrKQIbgg9ZAwNDOblKO
3yA1TuKnM0dNsIgeTrd4PYygxdTYZavLUQ3iMz47AzzI7Ks6kkEtpJ6yHDDMCLudtS6tAaHzvZHG
C1ApKgzz4n1hYWRiUdmPEkHQA3EUAXxqXqU9kZVuc4gWPu5bbrCMquH5+yUzq6Nor7SnU1EgHekh
a8GlpSJWUDoY/6dgViDj4IxBnMXSsv25vK3qqEWlqZ3ZEvS60daKwx2ov8LduwJaXFgh6epuW25e
Oq1YZfeO6Hq6jfTORd8buLH9Sgwp33J9sGQDDVG9NM6udGI3FfGipTDNKbjnMcQBVpZJltIdh9f2
44iZKYIgVtEm9L0u4K/+jFll7o7tU5yVA5PwUh9beqHZfqiRZ+Ya/sCB+kPvWTQfDR5/kgdxJ7fB
VrWnCFp+kSKk/LuMBRrPR8E9F6SIO8y80W78hZOjXy7l1s0JYoAXYny20DfbgdsOGdyxgynCCtJH
pR8POmJoYVbRKtXSbWVwVTgX7/BpoisnnKN0ZEyLW5JkQHZRFSKvT2rTGkcfoa9A/ZqvHPnhYlcU
dTozd5EJMl8Y90iu31obR7WGh6zoWgvtcoD1GsbdVX6Am+hihV5CNjAH+Cmvv0oiTdNfgDVW+oF/
hHEHDzBxKwEz5MMyZH1XtFGpDhu9kNk6Q/gbVYKJ4/j3nM1Tm0e+lZuAasXVx3yKG1ths8CjiPs4
5fMrFXFLVLnCv0B/3shruGpwdRYmleXOqILy/h8uqKVBQYq4lEE40zwnba4hNrasf1n0611GX7pm
JFVGFjP59T+2OEedS5myPzKHe0rzKd6UDEn89Pf7Pr76wuHYLa/UQXZQXWrtkw7yw3WgJSx6mptx
z9oxaZi0VlGsVu5jQ2/CiSZZaT6Cky0y4Stl5IeSLbFU4kPJgpxrslpi4uDQT47FwLec4iC7S97D
krphPINIVRZAkVxktE40vy5/yJqNt8yXZ1+TVg8Cp7/OOhkR1LzYY3W89fhEvlPoQxliECfSXXKz
KmHvlducqHcwh5YCjE0+aclo4VBl3+DM/PYhOslB426vbp+Qdj3yd2+qumY/rba2Qw/HRIfOpsUJ
Umle6+2937tyOX5X1O/uBD4vLi6M5m/1uvJMRB2yBAkx/xrld0cEYdcAZ3+RbrMgmM+20Gb7mygr
dNipcNrJ+favoT61jXrYGmw1Jr9T84rJLeN5v5DAfuBo3ccy4jYwWEItu/nj05xI0nQorqTW9iap
h5t4g4YkCVPxivtqaqVv+uNAzZfNk6TLTIZBnOam4YKCgtSGVT5+SA+R14eYvu+UurEZI/8EeVdk
1+A/YO/H2fLaVQVDnYjWNc0qI21JuKm1jhegr7hUtkz5uMhjAwrreWncS8Z1y5/wfvxI+ZeKclSB
upI8yQKEU5DcTBcgUXuv0ZK8ou/voQ69OXUfVdawkKf8wAfTAVh6cDjqeWEP7d6v2yytUQOSAUzL
O458ENmAtVft1dKoGqG5YCnOqKXk3j181bl6bNwZZeo2FXBquQpBEedk9lIBXCZq4+XLE6D+TuJd
4ciUmj9OkDcpuDHp5JCp+ZR6EzCCVtBFEa1IFg4qHUp8u/ZeYIQ8t4UjutFrNfa7ht+jhueVnZky
wCpj8i8gf2X7XW5OB0h8zQtsSzGDi03mkdz/iPk/4jTX0cNho6+nEjIaVqBq7ajSf1c3luN+/Zlq
l48L4SKbzgpMEQO+wK+wlQjEgpBDTu03Q4JYrHcB+aS4pe/F1HfpztVIzENENf1vb/YLobTblgJ/
BwKiIll7TUF3C3T1elE5v0wxz0wtYUyiyKWy8MT4/1sWaSL9jAWfvDlG9VIw2eb23AtV9z7QJFt+
H0FZOH/vl0I94QzXKvcAy6y6BMbQPcLsoDSAvkqqevUYovzSo4/nz1pywLpUPW5le/oGqVlLbKrt
CeBEMJKklrOq+9bpc0MgkxIu504u8+2mKYEcd5zkUC5AeoFur5WI3cll8N09FggF4RMetQ+8CE0R
BNkYs13lELzwLRJU7Gr852Y1NbxoYH8DWmlAv8i8OmVES88iBu9jFLjIO4+jxxRXYVaHoc2f5+pS
fSXhKbZapTaEOKdPL/gM4DxKYW89MrO0mftKo/V0a/u6w5pa5Dx1YQ1W9lj1RwGgW+logpo/LpW0
Wnv15FlxH0KO4lzMRZQjEou6Ug90BcKQdfoy0hg4lwi17oeFYVWM5CHmXfRKK+L0bdv0FPxYCgjD
EVtaHo8aLLE8rrb1ggTXostfjvFwzG70Qorbew3IyiEjCZxSCxGIb9abfu0hgGAbei/Xr24Yz6bd
PqReo3az9YRDABqiFKvTCMB5IniEaT75foJCasigQ/PpC65winlAG24S3mH1QEMxVoLQuJTUaRu2
bUaMNmKWJPKMSKDyWpA0w4Z5iAaZDmtPfKLv6BqkulBduVz7j+wz6j3uw8DuwUMGo1AUETwt1ybZ
GdN4mWpRM2rr81yUXb+6RG6q8uGrJ32yubGywkkNG6IPkwQksyPWuOeHC4XuMzU/POGL2WiLKv2d
rUgh7pLmf3zNjgNEDZBqdLQcZfqUV3jj+xE56YmSTh8eYi7Eq7+wyzf6UJJLE8DSWe9tENiAo4N0
RJUzJMfwzjHH4FLrKTJ57P7cehhLOQgySnSCOVWfkk8Aw0HX4uNQmGW/BC1qPTThSxC7OwXtfT5v
iF8ZdCtBCtExV4DYisTzev0136i+b3LAxwvcda7agaYRqpiIgPVh4J0Aymn/YQ5ptMKAQnkZUOxY
MCA1QySFH9KRwKr65UBnnBe3rARs3jwf42yQk0n9VaAeU2p3Ijp0kPMzqnzD14Np1ofBzWSlc85l
TN9RaAEHSVbd/rDYflKNnMqn4/u3xq9Uj1QlcWzBmHHTKApesm9+WqOOJG8D9NzjD0mym9f0cNLq
FfEaH60z/E5Yjxhbrf1+jBkQYJYQHUnS9vqSrNQ7opvtritteQLpkNJpvvsAaqyz+YfoEcMFRZWN
5wUIXsf8syI6zw4I8SRbBPGXU+XvADTAjfIF4WXxFmssgGASZRsccNj4+LztYTX/EdWYUCmXu0jz
srD5f9FCjsalA5QujKaWUL43r6hbz8OnlyUjKCtMvQXb/+s3F5JkHLweOhdXTSI8BTNDIEAJuhQ5
Ob8hIfG2niRwkit4balwHL6CZAIg+wyfsPa8jgE5/Zpau/O/R6daopGmrTChFsROGlLAtvNLgcAX
NncvYalXPNAfSWTWbWxRPPsC/B/VdnXRDh87bZVHX0wnp/hnL3wrPAzEpVMc6KWDR+OgpSCZ6ML8
osjTUslJ8VzdsBSsf6C2MPlSzGtvPGfYQTKZzId9szaoS3k7IaHK39c/eF7eEdcJsn3iyvmv/lC8
/tH+Cew9WifGoriUBUgC704geeEdq+SYAOgYjhpAytIOWPNsuLeplX+LJtIaIJMchZxsKS25l4+W
QFZ/Ya/c06CWc+jbGkCBnxZ7/O5WVlmfNu+ur55IhG4QVTsXC3ofhmRI6tz3NiO9akxaS1PBKtTX
olQAm+h0BGs8Y+S5c9pWiRwr3A4XSMX1WUgnlFKVu4z6uOKtQK1c5ggemBhHQQTJdaZbpzZOQqZA
FNEqeXi9Kia1rxQkDaONuf97cZr197+AXN6qpwBGEKQWSv2KnZ0KeptNKxBvTAFSqKyRlNSfx4UM
1vmoEkiMn+uDbYWJZx7E2JHKA3wpukgFaUi6GqAAdzU+liCLkmU7OTFjavDtzR83bqFy3ONO43ix
Y7F6D34RnQmZTFavxe6wAuPr1PZY60hPmFouh8ZZjHjiVvwXSH7r0bLWncqHZapD2L7SmhFxy0zl
PLU7BGTh6bBv5OnGT1uIAOtiK4rjmPE1JxDxNxdXFD09RJovjxn9rfksQ3ESmW/nzvOGeNvaohIk
/uAcvEw7kHExe43mc+88037dkVCWyQOAveMbOqXLPsxn+dyqXF7hZBfL2Y0pDrnuPYu2Kf1GmVpl
mJHE0WygKiI9lT5ABjj/wiNDTKrOJxQI5iGPkGISNC7yKgDa3luEGf9o7LbVZduuf2skQQAO8Kcf
2pI2cQXRi0gfiwKVPtDAcP+3jhtVF2jYBA+6MhkV6EwiJGVKCYZDRmCBt92WuwMso4NCFc7HQBj+
aeS53S8cRw4t/o50BVNCuBGjsixeDUPGOKkoyvzy3B+4wUgaS4QeJg+tLOwUWPJHb8wPwB+7aJ9A
6nOC3TvQllp+2TcXDTdZ4bHxaWXySS/ad/k6UcNM0njij7dttl0OFY08WU1Y542cMz8Yt1ASoitZ
QKNLt++cf4EtNzqL0urxFe6nStiJq9WBDjyr5Y9KHehW3F7nut9ytfKBf27FoJRVug2eqAUSlzB+
KpCIA1vXYoSm5Lw/ecohPuucWX3FQtu2KMW/hCQdF190aDwAUdLjq46BbQ0cFdIAwusdbTgshUk3
RXeVvnHVjXiMTNuJgqotjwJczqxaBrMH1K+gqgDhTppPnV6TpaMXeFbgKax/dTBZxbvePQ6nY8oN
qWdy7QuC6Pjzy3vSviLnExwpbCQPmpp83uKo0GPHzSMWf4Ke6Cgd+fJs99w56yk1qmY4znak7s/f
vtwORBtOFn+AzfFCCY9lleVEaaPP5lUavNAhVQIn2QJE7BQ6bTAKnr8blsruy4Dz79CP0WUxMu47
8rqOHzWI8HXrA30ZSpJ5Qz1iRv8EGTSwTQ63QGPxRBRa25MC7yk/5Kwc7X2Mf4rNV1Haa2i7X0J9
j3YesZepjWA9RRc3SIOy9fA/G1UsfTlQzm1o4qsq82dE3JE8PeQixJqfQPFsRuaYEXPjykF9/iNZ
GktHT3garTbM3GcZGp2KKyGbVPOTtBfgDplZ3Tx/Vv9EJjwFTmW3Ao2O4/LSexjZb+DFcA3R2oCA
NpCqmopdaOvi9w9tqNcmnOtGz5pko4U1FDdYKZH0o/Rt0q0fHITasYOzzDLFQWxNO1kjofYOIksr
YKI9+JnnZquyVDEp85E9NnzSpa9BS9nEg551oNN0pejdhgs6QwDc6j6NWoeC7dixWWGQgE9JsRpf
0P9G1mw/CAWxLyNWM9heBGgEL5hOGfQFyew0k7eYJ+Zso9K1Uyac2jsO/xWUnQj3gJ/Cxgt8dmpr
zgFYQDuun2Euy7VxgC/31Awc0Uwl9jqK+Wx253j32/oD1QSeppGp1CXaKDK+qF9nV4QVeTZlzl90
s/Mkc4cjBJGZWzNdqsaMBdupgzgcgDeDCgNoTOrB6tiRFYT4QcVLEG7B0ojALZl2M/RXJAdiMsUh
Jx+QaTkgCu/fHdJLOhfFymWRvF4qHX1at9Gq5Buwk4DFRiG5BvJ0GB4uWshM6N6t0BuT6oLay/An
arldEO4S+j+nXcngbwjXfpOsig/uLxftfP+xuRZmynbgcPcYc+hS+tQmXnBQ/8e63hPsWhVse0iv
BABzyvyq4UQqZ1tTo99dbc43+3ArFUl31Wq2lLj3HmvmgoKxeEIBcEundtaQAruzAZO5p6hn4EvY
NRzYFQxK1bEEZyi3g1AE/qaGzreHDU5JUWeHQbDLAYVaaOehPYq1FC670nqxd9S7nkOfn89TFXqL
rTjVVGVnU/wW+bqLB28pMZ8n9b6oabznmy6rGl+wKUMB/jTh52AtIZm3RwXOhZZ5TZW7kx4YT7VP
q0JCovDQMzHxq+YZfunpZVpeFDGlUvO+f+F+SpkhwhN0az54o4kWOyv+YrgAgpVuEBL0SH4a/gs9
pDREs6AgKGGXIMBBxcAz8L7pyGyIyUydInw+e4Y316aA76Jw4MK2KuAeVu6tuyjRHgVlTf9R4geq
lnoRK3Ayn70XbW9af3tbXapOtZj4CnEDqRFFUidLaDDEimO+jrpBdfvD13x2ml0sFrIjhS1PJyvf
rDX3Ignhsw45XbdXeucMlivGqo8krMGxKJ1R3ACJb4tNoV5Jwco+5SwYM+YBa3cny/jL0tRoOYBX
jBO9bWOo4vgbXhZUFAUbmQxNwyCg3f6+D/ncS549orlntdcKoWLaQRVRpX7QHJ/0J66iASTsSkpm
hnLC7Uc5cnjlajXwvgDnjuPQlU5B3E5mC7sAorVV4hoSRukH2ccAEYLPI8Yj0PHYa6Lk/7Viv8Uo
GexSL6wdRMfn83qgXn4N95UvDxzywT57Mbnm0cfQAafPWQy2TK+EykKXIx4+r0bxS4rEY4E+f+tB
An82uw49oVhjfBt3lM3RU3d9d8J+qy0775HMVQTJDbskLIczBmiL23SJxkQic8GXNlwad25akM3N
9ihHua8Vx4WlMfcNXvCjjWzE/xiR2L/3bOtMjRZ/dCcHqC3FG7wXpgX72HJo4TKIzkX7JXhWWhMz
5JIeqPgTYyU1RSgBHMdMEA26IyUdIWTAAvVlY0GFG4fyERwlgdLR7r9WFQ9zTC9aw8Hi9NgbOCDC
FS/68KRUaDASew6HJsV/gSOkSu10zQr/BVbF7rYO18rYm5f8ysCAnC/fEFtvq4x0vU0nmBTHwzIF
c2N0/U9tIpQxaBBlQy5G0QcvrGnIW9bgxdcQnpgea5SNrkxCdknWqGSaUK1cWrYuU3LIZr/vRhv1
qbilaWtVHl37qN5iDT5S5k2YP0niMayP1gjdQyeQPYcc4y69qURZTsjnjedCQHEGUr+esDJ7tuXY
WNWNkTTr5ifQv/iJR/Tw4QwemjSAiVg0BpSbpZRB6gcb8x21HAeSgawtbNzZSiKzgWKryhhBJCpW
5Dj0yGdmN/1RAZC5MVlgNO4Bd/LJdu2N13vS2w3xer6WYOewP2UKlryjqbjU8UtuqGTdmzEVhd8Q
GefT8J+dt197h3dqv+C2Ig39tOyu2oHZqdG8SPo2EGlFfDCb1aH5cEs+JOR2owOTeyjr3R1njO9H
zKhEZ6SMkpsYpeDf0W9/1j84uR7XaiwSBna2j4PrF96AglXSdKLl6r0bFlXVnKC5Htf9/SqThMQi
OwdvRHo2bHRQUlg1Me4r6vt7iV2O1zNgWoHPkv+norsNhewTJwiLVHT+8blt+8EdxAwDzoB+JkIF
chLZ/nEfJPmF/BcXWJeGy5TeUxrAjU13RgguOyIwuxTK2D03wcyrKtygChezyyveJa+dJieaFDZl
+oMH1H+od9Rmmsps07N0Sg2g/NrslMj8BjBeBqCy5BVr2QxZ65br10H4oxqOJ6UilBRUIBE2mTR0
sN5WEnnt8DHF7pDuccPn6MgBQkjT8oyt0VRwnlxkDpLTcI7fCbGbv1Kcb5hUeMxo3GCnlxALBGKC
PR72yWej4kt7Ef0dRxnRw6ld2sBVSBtJ0+ebB+g5QfIVRxEhKOZ0BewHYMjjwViXteVqFHp3kSyg
7tD8TMFlWYqewDGvtuZrJeYz00S/dvUO7veO2SFgimHUvD0Gzt19fbLj/k0SVL5CVJwDeSTyoAYK
Ip1QeMCZjlXXKmSZsMjedjbzNr7nu36L83D0I5tS+oUtrmF1bvMq6iAUgiXsxhArg3P7gAOc0ooU
yUCN0Qi7ys+auop7qrw+1jlj0F5TOHWMfOp2WJLvydZQrqPHmCa3PD0AfUr7IjrD4zen231ZzI6G
Ehds88Ur5cVt4Jq1n5e+VF9kTxRVaKTfJFU/tm609RThMYUODhRk5cm3c5uAwuX2Rx0/poKIZz01
kIcUnWmCqOlO3Zm0WmGtyDftLMJULi/4xAgWQOpWaLoFovJCDOxhhUCLOlzoXwoyXItdNR88P+Ko
1Pz2OAQBt8Xvd/ByS3vWBurHQUqklk3NcWjm68sPa6osEh3OMDnT9sPyspNw+lv8Xu99etYS3Tjx
Jt6OP5A+iKfWSVfb2x/cvF/X3iDS9Y05rastlVl5pfyFL6G8dAUXn/f8ddJMWHx+UdHXdl2TjwXb
/PasGYQjRTq6UvmoFaMgol4UopVnBKqmsgUvh82juqGu7YYNysj4Dce4hjBpxbrXqYvNZJ0lj6ZW
t5/d9ff+jJ1m2SnRqEH59/9y1Ww7iMNqCVUzzzMaTZVp8ZeE9wxI3SqtarBYrqjLIRaBJJVg0qZz
KN090x9X2EOwQ24DZjakfYqg3hCsowGLu2NE8hTyWPqPyTxR70G1bZSb3mlHadrZHeGwm3KV3shE
qi3/OzAhSAMLC4OU+MWeXruRxNVLaLO+N5XN1BhgntC8o0E0WxDaAFCSgnCa99oUN6ZFiqPN5cOl
NHMvrI94hUFei8jUd+5ltjd054HRXYu4yEPUufMndcaJOeVc6cTlNSr+jyz+ER7XfkYfDc+PEkt9
IPPPiA/9Y2N2Qz1Ql8XvhZXRplRXVaR2R2LjKaZcwzQ2DeWH48TShPyAa/BjoAaPSRW97l25FvUv
0nGwN82gN2LvsJW2pbdFjUyXy+2QnQVrjV3p7B1/fN3Af6w0+ZllNBFkgv6DuH11R/46yp8qh6s+
dkuBcz3kAq8yJnw89qzRHWWL/YKBncmMLCbV6TK53eO8WS7wjfnMsiXjfWNn3VVqv2OzihUz/nof
yQvp1UWNO49KENgt7wkvdJpHYiymvnMd6QDlJxLqA9dvcX70S061h4sxEGGsArm9WhKj9jIbiTYQ
/3ezkel6q411WFN9gyAE4cZtod8q2qyoPV49fGaTavjDVSdsDXgktTE9jwD2W5Yd/C50i8BAIetB
wShQl/FP7yhYdnvId9Yn3vMAmbDBbvHGD8qnvh57aozXpPlH6voWu0/5+Oo2arRB4mNobdlia7eL
kO13Jsfm9Mc7I+Tt77NC5BeD9sS3RcKmFrVir7ynsj4j5OQQD3BhVdgWakq8NCjFtr2l3GtaZ9YR
hKJ5kSITvxwK03tezKewb7zTJjgRNpJMgGhIFLSWhO3XBnan7f69UNpq73sovjGH1JpMVUoo5oPK
KKVPB8IaVnnif94Be2cimiYJtI4wvmSJ/3T8T0KYrzyCH+LWK7qSARqGhVKb2dL7vakEMJgtynCx
fAZpEEvLpU/Kz+4XPk5RBR8D25g5d2Us4R7/QIsKpesUw8HXMJpQ+ilYLpPXx2ecz24wMblJAEEM
FhGv5jk2Yi/l8ruZhTdPIqjJR5vEitBzN3sJ03ja+hjoos8Fq4+XejjOK1cBuYhJtQB//axu4G5B
jeCOuAjZQk0froAJOwNIBUmT1ZKWyL1kLd4B2j+qxx+/IyDh/Rq0w15OI9nhlqoXllxf8FGexosh
PrBX7B1QBdhgFAnTQitFKgmuwTOjfL0/mFFu5bsoznhYzgTVat7MlweyxHGD8RH4D2N1sb8kuaHM
AUrBy23p5xkbpS9K+O7ZUxRK0PSBgk5+z/yyYv/bSEVRMXMiWXRsh3xcYeDEOr9aXuwLTDK1XHP8
9UERWUzSYYWLjs0HUMmfHktbjVCNndUIKVnv9D2vJbISynAavDbyotPZx2xsiicU244Uu4G6AjMk
HYyG4BNfw4puG3+LRNxRkgyFSKhDp0KqnUJFEZZUmM6NyrsrtJlzIwX4vSq4iVIvibrFVYmecQN5
LsZ8gwdowY4F7qtSBGorlCW0zWRzajvOJPzZFpbpjrQTs9TG5VHrKZD7LNWF+PSe9padYbDP6LO7
pMs9z9OFrTcSfIlbTPyrnkHzsp5gOONymdklJf2fdV1pOxW4k+SI9/49Y8q24NrVAfukloa7Thvo
1Wzicc/7a9eZJctKu1SvknN3cHZp5SWuKtQUUUbga8JtjpxE080oXL70a4F1YFdmcEXJ8OM8eB2D
QDisFO4FlbEyRjfT53ITpZyuwxnjbj1TW0xHCy/rcuiEWpV4PLVzGC83aK2JHseeHkx58Z9ex7tg
dNJl0tKausExxO9kqfspEqjoGp5bgMNv2YM02Oco5U5Pcf+nVgQ1swvcTyP+vseRxYvaWSts2pyJ
YtoXG2z5X9/TZkKh+mA4DC3wE6wBRPsiJbguxPsrdHSYyavPd4mzPj5vDU7L4MnaSb/LjMBp0riN
dp6NhFl65UZFplZImPxpQc9A91f6BfNrxCgzF8oK3V7K/8vOiW2GpEK2CT5XpWovP1egLYJ04V9Q
IeGtRbQT9Ks/RQmGKExstIpucfz2eGSyyNHCIi7Qr9IjfgZWcKSk2VkvRz/h5xDAgiV2auvAlbPj
/wmNFfo+sMqZBFHRXAL1kv+GxojrrJ94rbmCFAX1skbG+plBwOkSn+yl6+l3sv8gb/qLe4otpNli
ImqlCoH3ng6qX2YipsCj/80noE8XSaPqdnhT/MORJShSED0qYegKIUFui0bO/zSgQaUCNrsZFmEs
Wt0oBwcYRnFZrX/iupWcwxKFE4vyyApCTAXxbOyuhm5Q1QwNCf7lqs9THMMxvZnUM17wRmZQ8RsI
sZKjxmmx+vbzCk8KJfrltPboGOlntMqNQMK0/VKnDkjI0+5Rzu+mTYK4egat4312M3DSn5epPLTZ
0zw2m09Cpq1Y/s7c/4WoS6ecjbHHK78U6Jll+uVSz9NBttg31ELXtJNOICHTcb+Uck9FD4La6K+d
k/xKOZuzKX92TwVneIPi3FhB8LDJTYa3aQVaZEUf0zc4tL+5MNMpXQk6e9Hj24hVHoqXHZd+Cogd
cZZH0Yy+3hbdHQldySq1/5r9NCUYeDNkEL2XwjqoOdY7YM4WKeiWSEE9gGsmV+Im4jiDzi+EbH3+
G92Bn4BWLp2yVqxZtkmCf3fdJOZlCern8SxPZxj1rGDDtHRj7ADe/V0BxQ7NU5A7FTrl5gAKwSXj
5YQpE2vJrPEydhm+rUyPtmlE6eaAMf7b+CHmWe1i+P8PN2mv2GW6jYG/gEV7t4NZE5r852r2egDB
LWt1zZe2mmGSMuWOl87FASHFn7D2rS1K+18J5CepYN0aSdaroBMiNSVAormehR6eaikba2mj2IV6
UpdJzrmnsy8BnqI11TWMs+xlRo56GVgx2vPOtiF1KJsh2aNZanL44fponBn6IJHdTlWzrNqPTWeN
68DBMLpUmmOGlluYlshCom7tYKFF54Aw8cpG0o6eK8edJYZZffyjgTl4TpZcIQZdnWHVsiwNVp0i
RQf/PMQcY0R6Sw9xRA5oXc3CRCTPdK5EtNV/MqzjB7U6sxhZJh73hhb46p3EfWFiFhclJ1ros1Xm
ZwJn0XKiea8qwVqH+Kf/8e+whpnO5xTyWtzxqXlFvZNq/VSj8EMp9SHyRhZbTQ15v7DxvotqRYd5
VDamwAEEpCnQnH8C5tsaQssD0B5DlRmrtCvKUDW4R/I1w/OwnzSHsOumpDe3LhyiBsYEDWiUdJ6V
MaFxjiXzVQ6YFj64ad7hFzKzJTdiPdiiIklfrD1Dwch8NFDZcfxTa/QEGoEfs3gOfxTcBR9Aw/AP
Jueb5+GWpYrVt3w6taCySk2JLtE0/p2Q5gXIFqFQZa9jqc3pXuoXqNWbgzQEXyvC4ndqy1FZN7t7
qgHXnrG3RDjaUiw1p+4AQZ1l7JVDsI4hInjIHVCIBrFMm+RGONAzBJH5C+m8ku5AfgC9BI8X6ZLF
ckWpyuRGb8+aCj2aBze4mx4rj4vxmY5dslxkG74anI95nr2H8LM8DJDQmOuyL85/fn7LZbKGa3up
tCbGSqb0A/1gSeus5dYaBy5TvbDL+wERak0hxOhWfHgn83jVYjgDjbFm8gaBMD71ho1UMhmibypv
Q+fAobvImDcY7sY2z+kJT5YqTNQl2vzV4imJb3huNyYrny2r3kHhMbLeehJ48ONcSY8U1Dn2TMBw
hTAJjGx5lA4GlZzJKCq3fQThaKT6nCuVU20xjDRojFiFi7fzW/bWIXddugRXd8HeqD50uZ7VCMT/
UsZazKB+NB/YkiN86oAVgn9+Ra5uy2G0QBz75N4eMCi3Yuh/eR3QHBZc52su6yaYPnV4ut5i2N/l
pGSRFWknS/TAmwYnzl2nJ/fb83LVCfs8PRGSdsp+Qpk44gqPfcBkChIGawxFMkTFw8QODQY5MCoE
UHJXAanW6lFKza60gXRDCyeiUDEzrpWQx/Hq7qORbib3NQ1Kv9OFjk1DBhqlUMSdB3fmtx6BMnmh
1vTKyFqBEcx08YNfXAX6yNVidyGaNX/lvYqcTNUqRjXRBuMToCibWNAeAGs89m9ynj0hIV/MJGH8
8xrNET9kL9RaaV2kRDFIzUEvytu/xSCw33sc7+LPzPrTSR4Vk3PhDgTwvpxeWbELrBqAMrG6K4Fb
bOKy90DQmKsKvi/JB0AYIGUOSPL7GrNeMm5AMH7jnY2p+2lh1+Q4nu6L7vJPCSTASeSUm5a49lQy
/DT4zJ75EOSYVr0KrnC2jt8Mykez5QLa6yj24Mq/1vdvbyD6jDoRs7tm21UbkfRqughyUD625gjU
3RWRNjuQtbmSLttUZ/kk0djg7lwCGWEMaVsIpsDkYgZzCv4p95Ufys+ci/DPcn/jq8iZ7KXaOCg0
TGuKrPZLmVY9QPGedcZEKUh5Qsfkf5DuLRFScl19fFlm6HkW52Ha6rmZgsGJahiOHxpHNEvj2iGw
sIv9ENmt57z4BmgsLCBt49h1Nst/fYNZWW2Aos0tvrfeQ238jwdSa1Ggr/wSd/gexqaByfyWnPCp
LRHxhtGRgZKjS4+UZHKxUjOZyBwRdmA3exqtNMM1kZ/Zsbcb1De6P32tvrlYiMPZvY47BRZvM73V
dK0LlO9mepZ79cUG02gH9xZlnZC04Q1k+ilLGBLCd92YERwRSBSX+UGMvGX+r7i+zQ3/XRNfedut
ESVOYFqby5kYRoaIwg6VWOqGqCLzVm+QA36N6DX1d/ikgWywHHNkyehpKlXn9jbXKJGMp8PKTOKh
I4eVxmA1Xt1rmS0Iez9M09tv4sMj+AS+cL1B2Qax1y82MiYqmapbRoEqbhhCACJKgxjdCMouGTqk
sEzV3jsgvBHAq/EGmbj2WOrOLgsWcmBYY4/+zAggbs9FxvBjbVG8nzP2URz/YTq3FTv6E3dUqwhD
M7dxxQLAgKasFWT+pvWI6T22LabPtKm3EtwP8tArt8Aj+ObsDWaDYeIr0LLkY5uzmR5SpTItjbKL
rj6uUmhA8AdOJVNotaw2ajmA/84yE2SuF6/LO1qswE8g3tpylOdXPWA/cYiR+ACHKXlK6S7KA2ow
ez5IMwy9aFfqDiYhb7IPzoC1xvsZkgynxnKzy1BjIdhpezIf2hu/6inbRlWCA6SX4FGH8W9I9K84
gWqvyl22oYdIyFfmCv6COB9AnwC5ucVwVF57aoa3HTXdVjTmQ0kG3LoL8r1CB3IFPtrAb//N8O3u
oXlATndT7+zPxc815f+nuK9e0xI1TzlzqNXKNiz2YXblWF2AXaK4U6jeiK7nnWNqLdHUVAm74MaG
f1sS+9SB3dj3Cls39w6fxC/VebvXCPAmPfomVp9d5CyqOeP/ooUocaP3oRwmPxwzNZRkTRbcipF2
ObE1nDov5zYANO2HFw+LvggHCecAgpC2/YUHJHa4v5S+2sUzHCfJCbhPXNpLB/A2apko+z6gp6FV
bPUY9IYcisXMcQgFSBfdc0FeEsrCCm0JZzQSUieCtvEqDrwgr4D9W9FsHblAZJTIN/fmNKo8q2pl
zdxHQ2Vli7pUSuYjTMqI59uU/v5m+yoKOKcMh4JfZoGK/nCt1qwTN/3PHmZH8mEExwcihrZ10vQk
uMsP/VoByQC3dJeERuZRrppTwnBMUsZoTA/D6yNkDBicJgLB9HLwQ+83tveNKX7Rc+D+hR4PNcec
XeXrD/KIjYsPW89O4sn8TTQocatANKoPUUIWWXJw8B7PjrXyNpRbIAcmoEkZ5ONpu497W12mp7y1
ZD4KOG3TNG6oYv4AXRnSjXmh8qiUFoZ7TPGhcFXtYXU41s3K84OXEjCqI8WCXMWa2iwl7NpbzUTw
ediqveAwoo1EYxZvq49F1oOl0p6Dt5mkgxpkn9BnvneYdNa4WPTJwRdAGiPRATnOOqvVMsqAm8FL
LGodpsGyzUPE1juDscHzHkBdbDQ0Ffrz4pt3CGOULChNxxFn9xCCwDx2E1BSk5/uiVljGXOZgPZ1
IfF5aCm4H/Uq/8vaxLyGo8VUEPp+KePAywixy3D9XX6pe6qbGDdvxcqjZzK00abv4NBSM4+Aqoc3
yxrbq5++RFtQdoApr6ZQh1+3rM2vUR02A/sOA0tprNCDf7lWXwdpEAGCUwRDU7KlK+6ZIoktXV4A
GKfKC/ZWWLikb0d3OPkmxe4/lopbdmnjDEhrNdjWv5nSliRstJtmJIPcdixKZ2bEpN7n1qtLQVbV
8AWr7CSNPRrdi4arS1afmFoPsHbkDQzh+uFiup1MJlHZHAbjFdojuNDrF1FWQH9/SGuBTPSjVkyJ
Nm/v92zYG/Iuwaufmzahdx9eaxaVQvkhvZ/SmCStCeRsr/7Bb+6stPxLHQAx/qYuhnmPkb7Zd/3z
l09nUxMLNLNhn8DbjiFz71h+VSpMpaD4XgCiFopUEkOEOxvSxnr6af+sfeFhX0QSENYu7brrKDES
McoCBtZJH4erf4SADpkdKbbddcHAsMh/ll3BxQPRUhnZH6CUML07mHBG9c93+5vKtmVocWnT+vPY
Dt0Nc7be28Z7Ww3m4u82VP4YT+yFYYjhOgLBNOXaHvIVdLAVo5fotU8Hn2CLeajOd3684Psanqmy
Jh7YLGDfN7EG1IzGm/UWE3fbvsjE9cXKuUuKQXB6OsBY0rLmeYliaxQ1L6Hdm2WFuGhBsvBHu6qk
8Uoggqdnip2MDR1P238/eDayA2PAuGL3QyaCViRdgsXjlvRtSy8q+nVCtmWcU9vceeP3T9ycf/kM
cJOYOozTKEBwApU3xVqV6yVEUkghwU5pjwoxnU5nkkL/Z/EQP2DBpB7aQ/8m9ULcw3ehIuKw+/uL
9+UTnMt1iPTDHpcmAFTinD3WTzq2fG9ZkkGzKOTYsBWBqMCr7qaJQqRNMGZ4U6g/aQA9cxp6ZD0T
mnMEIGVICIHoFDeWd1svWl+A5j/Akq0RYJBF8w5lqBw8scKNyHCiGUjNiYo348X4ThowZZqrSwz6
uAVmPd59OlEF6hqYWFtXAdmOU4PLky+THThjvEjx1yznQCtaRTZAnN7vnPAAXUS/+Ig1FkwsnZuD
dicv49pz764yD977lIYzOfu6GVEOoqPGoLIVf804gpjOJESLuYKmwe4Ncd/A1OAFZsF4yh2qX7wB
ZkpkDfUYnBKdllPX/+XSVpIZ6GmW6zm49MCqWBJ1eI+mpxA77LGCxBMUha1K5wCsYJaczX+lZow7
cIgfAtb3AEhNZNM1W0VW50ewoAaF6EtU+6litZHdI0Hh6OYTEdfPX1GpYQOxBj28I+e7Pu7Anw3B
9kNmGIYlyKPw7XTjPNw3cXFaWtEqvcVEVlRXd2bqhVfc3ktMSA2HZPcVD5zb+HASQwVwUtjlQkwr
kP9dImD8qqyq+jldCuDlP2vaMz7XTlpZylY7dMtKEwWkUHUotmaVdzqmr7ZXlplCM7xOhaIWgCQ+
+BBXzgWgDOKX8VTNSNitEW90APlzpCjYNDJjS99GjbH2Y8Zf7ibeV0gXyDzVcs1ymhgIRheMZktF
RZBdpMg0X6N+sE8TcUeUJrK/ComCIZaiHR4w/FSshqEBPdsXTi5XlHjSGnmfshJaHi67WtuzThPP
FGtilYJsednOvDxoKbkP39cRjsJkAZnUEtQWCtnDQS7W9GzKbH7HYBE5NCpB+cQDlCaoNMYLjskq
4LpMCKe56YDrUHfoyqHdO+/cL3Ix04KXFZUjYSWT6ghLDGEDChm8HQbd2pJJ1oqvjd/MethGz3gq
zO3Eamctx5E4+D11kk2RfUzBJaYBo+aKyG+S9NEDKVX+G/rq3gUqDgUA6piJEphUO5zvjkcJDhGX
tpv3ao0uHvyOVaanwlt1KNk1st7gsi7Qx7FFjqZ9ARIAEJF7YM7j2+bfS+wbmamBgHf00+APrJ+T
xxDl6toTabPZ8YYndwd8ZcmSMJKfJy1iLdt/U/07qoXawgzL1wY+C/8kkYOXAFJ1oWjZB9zNkMtq
0AYtvMqubJxm6rSCuED1vIwBTdzG/u42ekTOnBx43idPpWMUxVqfJTrKT8bajRf4+AuWCkSjDHOj
oURuhwcJ1AuchqP1oIXupZj7St6nQGwF86/LW5K3z4r6ZKM3VOFM/WvGXifs9uFGxr6/hQ9eqyFY
laQrOFWDXFQypMCjxKRQHj0kHkAuWXAfz1Xlwx2bOgJkAyqPlidIGliMv4HDsQJlNfrdVRlTbIeZ
MeMRhOpVHKZCgC9Lzvm/DV6IbIazeNM32cgyeOtf9cWrZgidjvTNz3GdCsl5FJiynATOZJG+Dq80
2aYQXRd//HZBmFD0E9t0g12yGUub4yQW73NukHr3ybn7Jpg+gi+1+Pmw4/280Oxl/nI+kXZGzPcC
wRDeFcMXI53Nji6hzXFf3CE5CNvkZkWrLqSoUT5QHgTR0mmnuEGGnnLLbC7AJ4zqKdLX6y9dXvDv
NFqsggeBhU0a6hZOMFyzyGgQ5GvGsn8vH7diZ/xiKpi22UEi2idB1yHtg0GAfAE4h0lIr2dCmH6N
KTgjKtY3IlR3KX/OfRgYTiGrTrKd19TDGx0im3CbVBeJlCnyOrj1/SU9seuPlaiGk+zJEgLLqo4N
CR9SrjjF6/3+W85TpLspVWspl6dJ6JlUoukQzLdoXLShNOYLb88xoG+JQ0rcWd2S7S14MgijBvbZ
4f6RfyFv6Jropkzh3bHXpq25GWe53dEzV8Ow0sPb3WFap5Fm3VoXXEbR2RVxKNPsP5xLGNjrTBOg
lzh00reMiojgxzory8NDL2Y+XoXg5yl6HG0x35Yp+fDWUDX5HEu8N6FJowuXg2REtq6EJbj6BBmm
TivLeenp0DRpY8bsKP5W+2jDwgASQY9GzW56sjpmuWYJegy+VVdim3WWt5cMBVf2U2MO2IvxVEbG
hypjuolQuiRRedGTxBeId2kqT/tK9J/XPn2cmXvmc0esOx7f5WO7LNgoJfT/TMpEku3pbyzuXzmc
a0qKO+MqoVC0Xz7bof1GFT53OHWKAhtQ0RJOUo+Es2X8s9rVipNYSKzxYKrur0glgvKkvE3H7OJT
aM/WEm8QONbJAWvm6QLO3XoO0lwEYVhKfmYuqJpGa+2qed4ogt4ny3v47HkI9lzYOQ0yb9t7+fRV
DXycUT9Z1QRXzeqnMAiKUSSCc0valTZzM7Ea2aVEYozx4D6oQI+nIN5Gv77ddigWxkTXJk5uyCIp
jgXga2O1nneoJxvV/6VUNSQWvEK8IkV1TQSElDVx4NY12uTQor2c0CmlE6PK1+rZav+Vnt0nbDFq
43ttJ8pnMzYPNOzNxFn9lBniyk4KX1jZcyVcQPgkl81AksC+c/ck5mxiSnkMA3cKj0phgK5LT6jD
IkCViSVWx9FbUxgosBDAGOL5WXdse3OT8CwrEUprD2lwk7kknui2tIuf48xqr7GwKg2JCtmdwGJF
QLpUQ1QMFdB7iMK0UV9T7V1l5gTEkfYXDqfDrtKPX63RX5Mq+Rb2BdlIVBr4VxCtCnWrmaZX8uLb
zsvmRW0FmwhUh9ICds/E+qAal7IvBXEypuMPuJ9C65VBWxsj+nNmAS4ILXO/O5qDrzegJJUVcVwb
4fZgfU7jQPrv2GasVPzoSEI+YvAtAtsZK4/q4LaQz6d/pwMZg/YvZjHBEeI3avdL8i4AoJh6+y0p
sO0SaxQxjqI+xxcPKJW0Pu1lRrAX52Pudpj1Ep09Fs1HQj/V3DkD8DB5FrWO1DtYT3Qg26UsXB+l
zmUvEsvjDYBEuNetbHKnwVgWe+Bg4lmqsKrrTb+IbLSTFQdl09xOAMrnQ2X6dksDz3b5R6INGfXW
fg2CnVYxQo6Y+1RpJxiWVHNnG7p1+D+a/ehnojVXrCkssrF0VxvvWQPnyfDzBaWEf2RejnZ4L9xn
KD1tguQtHRfBz6yRxR8Z0gVF45IH3Y9PAfEeF8jC6tFHCGPLFd0oM/CVl1z1gGYp/aIIcvmCSn+8
gD3NgKMzFWoq8yhjl8XaXJZYVs36UHMU574mXSuYKRIr6QweKBLDcS/0u+W3AyE/2aYmbneDeXIh
fzuPR65f3D3pdZaGZuCWQSgHdvb1cpDZu6/VfAWcJ6fI3ecH5DoI1yeDSiH9+DW103CfDk5QDie8
WpsIAn4UfuDUw9uo3hXt8J+aa9FIz1CCQXxydvW/dNeGqVfFh0l9YQ9gkDQYDopqg67BoQITAn90
dbc5tTcC5tNXqE/gG2xqqaN9sL0ZvKLln/Z4mZvbA2JeiPHXjXQ49zUftxnZA2ZIfLNb6Dp0LMDV
s4d+oHarXj/aTSQ/xgN+hsks5QH0P+g9yOJRQSdjVqDZviBtJ+e0PYCv1+xZgEuAPhBRwOOEXWjF
XmYHvwVeSkVmJg7sX7dS7lzd3ForTOrm9tUAb5V2Tdx321xO3uKbqRrUrbqENk9SWDbcX/135zsN
MrlMcxEcCBeFFKgIRNJt50J2jjSv22N2lAYvhw8iuYaoFJlys5xJf+zIdlq/qL6v7noDuF2XzhfV
Tu5q/TghnJF4JgbU545PQ8C1aeH2BUmsCWVJAFls5kdb12yeAqCKDM5oVXwFwUr4zjdBsRLVYoOd
dnAkzpz9a+vZCHs8xCsTcCMg49o0nmm21G3nkfGZXxYWDExyiZw2zjBpmwVYvT8tlKsAQFtCh4/9
qoe8dWFF90v2oB32GkrAKdYny9MMFGFnnn60ZSa+waBBR62mYBAKH+qBmLat6Top8eyifLg3y5At
gaRiNdllYzFIEoW8XxoClFIiLHrZtRTox0ZI7hHVJ2ix5xletsNBYoxLV7jFxMPUwDcPUgBmXGo3
Cz8EQ9fZz8PCJN43aDhe1DpAnZe1pqw1JN295ALO0uYm++cPR4Xzs5LV8uKhrZGULp27WOv7nQ2w
YBpx1BlQadSx/0IHaENiyNpz65ABkJISZmLn+gKtjKTSTpnRk48rFHFHwz+tlZoA/qwaczPM4RQS
WAztxObDH1eMQg80Ao5KezFnY5FLlAxlVZ34akU2etiOeRpMW3DCChENrl9TC+4dzgBY6xtML+y2
wJ3jIaz9CLlONFq9S+LkDi3OgXcaoF8AsCC28nO+HHehVq2iJVsYC9LYfdZr1P46cxoZVlNSg1gZ
nAJXSArS708BLZ4xnL5/hS9BouURcwigxv73CLLPEiiunkrPiODJ5xVdA4eL+VsJ+G19Fh9o2cCP
m6oIannaz/Aw3r044U8CrtfMNnJlBFcmC22dWHUPTbguBdFbNNxS53xx6b/d/WZlnbqV002apb/m
u1PVfwBBKaCagyJ0UyOgrkNU3CjlzOtRHs8CbfDjDiEJZiteRd3ktbYh+bzdCYkpZ9Z9yz7B7Xaj
YLyp2+cEO93707+BcFtRLEGJtDthJnQQMGZyY4yGlu/u0vTDBy6eLlmxmCFeAcNHyQmVRwZMFYli
BixKLoI3iQ8BFvTif61H96hVhqvvLOIgogGN3NC60EjriPvRZiJ7Tlppeh+JDxioX0/4glrJUJsa
c0jtQwro27NderXcNPJta0wcFnHENwDMt7FVidAnwVOkuLak6vbx1fAjjwmBokWJrnd1ex4cKHH4
1TqriZtdeKu1XHnioR3lNXYEmBOypFztnwceoLU3Za/OHKTfi9mjawDzSfGFlZMdZLKP1dxhUK1i
gyerniAH7+nNlPrNsdPJIGh+kdntzzOU8W2Vb1V6bH4GFa3nq8EiyP3qHikDi/+y/TeOE02NeXR9
04bXvSuWKkA5u1+ls/0+yp3bnmiruqsQ9smnb9FrP4ssEG/8XXkc3+edm8RLNr6+Yu1ZMdkJvs5Z
NXZcMUK4s6M3N3v1ht+xT9nQQ5NHMmtSDlmXgxjc2qynRk6KkGyE2FIkYy3PXwkiSjH6bkHHduS6
MTfc9Nk+gBE+slJPx32RXiZIMNm7MA535Q/5EavLhrpRhYxo0NnLv/9YVZHV0XFtmK/azUtz+Epe
GKEfIuvJr0GfYszyLWxkKXp7HA5Wgdlti5Qv8IlEauJjXX3tiCEq+22TDgSWhGFW/amOzIuf0sda
XYkL8Erh68v8rSSBB50Zq2X6xOHuTZgYCQfxnXZmOUcJ2RQFaqr9vfqdGcUgkgQlWsbFHssC3hFw
CqDnKKRcllR5+G/mKc60z9WWiRsufKGPWRyNA5mhCgn7B5W9ZmzB0Vclr2cU4eLeJ7TDWnHkE7Ic
zN3ecA/DoTa2PFqJu9nV6y+lxKxYClVpgDvJe2YPXksIhztv/dU70hGZGL73srP/z//tJBpcMtdG
AxIgD2l2dNHpfhxpNrIhcfXv793FXVhSOzVCvEkRE7dhrOrmbtToGS5PHCMHzjsHbTDx4/43/wL9
T1PSgmK9rsec8TZuLj2GRxc2weUgNUdFZRPePdtcIRshk3E8TCnD/g8Pio4uXyoG/Gjo1OriBuNk
qFpN/g34GmKhpRSlCgBU8EaxJk8xQZlSTi541DBUEoBgSFHQUcchPwzK3v7Mb3hon8HWzNgfWd54
liEiG7hOdRW/ESCWN2SnZTynq/cvcd1Xl3d+ByoaLR6Q0/R2I2ccfTqQmfPzjJ2r98ydiB/tpmdq
HyFBcY5U1yf9s+byn+5irsQIxBSLfziCkobs9ir9BiF5rujMExciKLJjLvV0iWbu4xdDhdPPz7U4
kAsZ6f4NG5HFkgWkNb4kHfM9nSyRrHQC8en5ht+BR88UpeL3MeEjwvRLqEKh7ILmKmo2Zu/Xrcil
H2bT1BTIRjfT7fdJRR5WIZY7fUFGH2RR1G71UeCw7u1ti/q9HQsA0X11nHazDFv0bDgRIK694Bj2
tQSGYdhtpos07h6IjeOihTSAGaWLivrpwzhO2xHRjB4izsMLITVlHXqIhaasNKkGUFpR53kMVcPB
9ETBbOFoixRHhFL0a2l5Yc3ULf1Q1B3x0HIXeVunlYtnR3t4AHRHKX2Q+D3cwRMeGE0r/szF9RFr
4SnVIsl37jUFyNa1WsuohNGZLWVkssR4xG6Xl8wD/R/lRvuNZZCfyXSBKAptPjYR1ugIIIAdaGNZ
XOWlRMcU4pnwEPqhn+FZzw/DHarmUwfdwxvgQqNPr+38y8p5ThcZqTZQBgg1upMPjxlDmhe+ASev
5EGOofP2PSnEeFXV3KwzX9pjROBw3WD6LN8KAAcTnnreEaCyYyb1sNEQzpMl4Ig59IZuXjzVeGpx
pT6Mx1kKTU4NIPWaJwNgrMcbefAC0pOkX/ySMuzQovvxKIvWqNn/lIiJkDUax+IisEw9gGXS6vUq
UNrfcCT9IxApXwjnWJG+gW/n2ylTThUPGscNCX5widEiKlt/wVkt0ESdMFazfLt7AnRgCO6esRlt
8EVR+3vetUC8V72NRCybkgYYeX4bcApl0PFUGoqYm3+tpEzrmYnIoBhhggDXKFbMacS/allS6mHl
6LK/l4AnuXYiT5OOG2j6WQ/NmImThO9id6GnR1IzIL8bTcjjxFJRojExH16ewbMSRjP9syHnTVZG
bZpuTVTOhwAjQiYUo7//+CIGBniS6laHdmZEmIJFWmgYahJ2FcBfjHlQU4e00QUO4wOKgEFCZ+Tp
d7940YXKsJ557vEAGh7UEcT3qkXi7G2BWaxEMqmkeqldUG/1njoSkM11j3WPvlVwbnA0Q5C/VHy0
CyPd41i6+6WeMVe29lrsui3loBm6wg1O2v0uhbfrJetyuAnVNiZdQa4BaBv4RLoGeW+Ad3/Cn8o7
sju93/SDTZZ94WQRcJxeLI3uVmYPoyq3er4ROWoHcGF4+jR2RdDI50RCXmkHUH0nWD5DHaagOh8d
CIxrdIrOHeei9aobAJtQLciariQrh+INycamPCgL7SYYJAEJKtucsgtAS+DF35AACMpp4GZhsrb8
cjwc0vZqYlJ6JGEQDJprUdATeLncAHqqq/avg10f6mzW5uu7en/mYB4hGNWHvK6G0utupLHtxctF
rPudYOtR2upMXXc+YJraWeNzQV2hltJ+5kZ5lQV4c2yNnJNxH36E8SkXt2T+LQJF8eNIl4cvJj7g
RBUDU/7QordQzOoKzE3eBMmSwO9q/A6FnWXLI+Kb9Wdo4acW3oYSyMMWc2GFYOw3iu2mfh888kel
CTZzpLcuDn4GCfTQlPRYgaD2Cjj+l/2AtJbmEN0BO5Zx5QZSZlB6P/tAXq4fbyNsqBcpUW3abJXm
Cnhjj1agb9xYaGuBsdFV/apfnGCdRgOmWGi5PuSYt2L19wIAZs3EseUbben7vg98w9XSFnnAQPzP
xmL5tLWYPc2V5JbyjL6LIwJSQD7ey/CQSGvU62t/zPsVYpW0yq3gsb2/ZrBXoK1W7EY6u3ueakRm
6X0slbKU6OIZLmmS0IJXK3bj+QOHkFtTxqcAaqXXKN3d8hHsDPT10bwt2KMAoTdiAoNbnlSIvbpd
SoCo4F+9vXYkE/tbSDhC4vlqF+9/R0UoeF+bl5nTXVLV5JPsBaAijnYfijXfMEwld7jci9NTcQFl
cTisKQsIEnVIn2Ou4K2bn7Ha1KxpiLzLPTqxVChjHfswGYQ26MiW4mVHqj9XyyhPpy6Yt2oRYSoJ
GQ6ji6IiUQVWDZ6Fe5UF5Ztn4fjSGJTR23Bl5ibZgkDdNVRyOqidUSWqxnVZa1jpn4QENheI4GtR
3ZtMar/DyZkh2NjKm2Y2LDlbNmgh/3cGzTBzRffnDxuw+2pL8xHRm++pWWItCaUJu4KmGc/fQadA
iwWQg78qBP49CjW3Q2NgGRIu9WxpvnszGgsLZAoqx2QaFQ2KeA6/DdpuXPoK5m7LqtbLeL3n9VuL
EdhsSh/yHxfBbk9/Wf5RsxarP7497KMl8hy86g85RvDVAWMYd7K+QwhUb32l5ePuyRlS3JRIyiQY
BL8csk9cVqLXDnRXjsUOMu3ypjyLj+d67g7/Nn0y8g3vcWJKhUFVOiWWnRHUzPsDbriMGQc2x7q6
rwhNRhrqa5R6GjxzSiMyXCBbSD5Nm1HwWi9XxR2NJgB0rdcGWO2cETA+dQakRMBA0+HVWy7aiHX3
2kaVnqwv96YloVVOJR+ubFD27jw4rJiDhK/jLmwC5E0ieldg0ybpXanqlzC3uBW/MnmMNhjaDBMo
F1WXU5nS++2mnk4a2nWDXqxS2K9kWp8Fu9M9W1pLhTBzKTOWYzL33VQWQrXxnvp8170/9ac8IEur
UbHdnidgBsuCUrL9ROSWBpitXtJIRKG/aGalGrIp8iQl1Q/4SkZ5eRhDLbr51OfyZ4cqUGwhDlp0
YIiv5fsisZgQ7GEWjcKLopbe2EdYxd4Rk1IlIsKjPrj+1o8BQRRTeUgxeHShmLGeREQmEfEpNsEq
XVvYvD+5RjotLCmo3kYTpCYcqGVyyK6FUrLKCUdCvVywE2rMTMjqr3jNQkqIjTTu6MPUKHCLjUof
bH2gQSzvoUOSvpQrC8EjXJyCaz9mYsuu1E+GikroPaE5SMTlE4xZtwYuDHrEgduY/UvYmIVcseeY
sfx41RbRrN5/L59hwkmXkCYjJwN9mGat0UKr5UvZRs14Atwqa7IsHK56crGMPXmxZN2OFY6txEA9
uymGpDeGybvV7jEUO671WWFRBQH4tzhU7QOrEzDEgMYBFAU8ScJz58QIdoMSRooztxKQtbz6lb1J
bKMyDvtoZ1nGlS1iy4VAcYmSEh1WbUFCMaAAbl5u0O4ZZ81/Cyv/QOg3alFr+4RCkSSX9ua2jhNd
oU9crT0DDkzsGWsUKPtCxbZO1HCYManRQ8x45k0tzjb0+jPXYnS+3IIMUQVAvzmkYDsqaohTS4dD
jtFk5pg+dT+6106Vl7VS+KSVchWEccEQwrdqZDeOI/AV/iGeK8SkymkWY/1nqxx1yOeN6kmkWuqL
rsQok5Y3NzEKmKOjrKgQYGPSqpHjX4rMa4PhJgiMBthauC9MW8sjkG9Wi3QbUFO25/yz8y6Oax+O
vGFbbipCijjG/41bdHFmh+Kr9s2aTbg7KmKFCcSSswmmrOu93P77stQGh/R+RZwICAevqg3C+S8a
50nXep7+ldggEG0L2LOlNbXG6LXFxLz95nvX2NQ0U903hak26pfSv97m4cVZzH2/d9GGnKX+290M
/yf0ePwz3USr4LX0iQRrbUayWPdS5xjS/lkXdMdY9rXSkF4srS1Fqfx2xxIqrH1ek+XLkPHhcd+Q
yh4/f1xzmDEEhdi6h+7W2Umof/lRe1N/f2vZPoIu9w65/Tft0O+qIcLpcHPRW38AWPaHQx7hupTM
34gtIy4slQ1b8vyPrKQxIKP3Qo/Fovj60kSCW4cI6vMWhMH/4yuQSjZfya/pkNw9HYsSXM/CBwfb
4ntHDILEitB4SHcNtlD0dkBHzE0fvhhSsvu8EXfqxH7cvT66TuCvyD1w4J827tDQGBpWo9/xLXVp
TeDAsFHxY+DKA5j4n9crMzSplctDTi0rlCbnh33LtUryYAc8qF6gGFQEOLfx8DEFFru2ibmju+MY
TFQG/DF/Mgi1rG367K5QJEPaSuQj9P/qtl9nZChgm8FCqeVKvNyQye7b7fjU3LZ5qnklcl2MzM5s
540jO2jyNfNgZoa2SAurgPVv/VH5AY23l9VsdGoHUqqeU+KcAxlyROjfWNfghpppNg0PkMiE20/K
UhA37fI0+nNTGLNJsE289qEKhsgmriWoucwYIFN9QituXGx6cVEER6OzY9vLktxr178PeorAcxN3
DtdHFOSndJ0vunfmzJFmF5OeZYuyzo/bCcZpACJJMq4JtFkxo2Kft/qVsEJfRNr2P4DTcSM+jgSp
YQbhvsIVC4ACprWQ/eh7IMqL4NGwNsu4asd0/rXu1yDW6g9j+VM67rfYiInR+Lgot6hkc+fhocjc
/TKTW31B3go6qUU0u/Ajzf7xP/G6Xmw6U/G0uRGnIIx+G3XQE7LRIQ/eDw10Es4XIfqoHFayc4G6
dF13wBwGy4SWOGffd3FC9LdgVW+GBc0b/cp7sMKOtsPpP4Ste8k9TmlXlaR5US4BE0g7jQtp8kis
NTBZJOTrdDBjhuhjS3NAFiv/qpCR+sK4r7aYNu/CdmaDqtDgkYDXgqY1qF4dUqW8Wd2iywsJP2/7
+Hr59snOPgNlQjbuXTS0mFajKHmuMMmMPcJtN1LgTxVHOYXeI1TLqaiQMV8hKJpHxqbxZpzHDC25
794RlvnUWKvTvoUNGTssanqSeXqbUoIQrIm7NOVCT7Q/+CbbgW7iChQofzvYeWVkisqug8Io2/OY
K3W50tfbQKYVUdsfPKQLWHGQf41NzGn7jdJV/0YTEN0y4pbNHl2oMck6miuflRfZVcWxzNB1BYzi
r8neuT0uZCWqmbd7zxtGYMeNdXnlnQ7XCsJAdq4xEjy5K38rPYzzxJtJXrCkvy/LsI/bBGgN+ATr
tvVT33fJZXNkhraaW6vqwxZ4R6x8e1l8GAFFD2kTuyAx7s8rj/BJlFMam7p37dAaJCXfPs54fNCR
35FfOF/rN1Xz6kxQbHoi2+x6e/qLtM5CyDPOtpbJ5+LChY2XnzGESKXybwOuB+5oNy3EQkMEtUqM
n7LPJDnDhoRXSOxDvR9IF6wxsy0ibuXnmERATgSAcmibmT2pHfIRU6ZykVHDHJJ6S8XUgQkn3vzS
tTEs++azSvVxwIsYRGsDM/k4FztIsuU0wCu8GMHpLk8AtIk25aOyhKl5FOh26O5x4XBYmx/YhvqU
0j8U6X5U9C+kk1eNiXrY0tVC1RWHrqTd2MCnvF0RJbTSafIlbgUVIMwaZYvMt7/Tm2HzO1xQL0DZ
ys+YcZSnacr6lqbzJN55sOoLWEYnQy5z4VYaO74wrga4Yl3XSMzdKr3zNXQZQUpkEuDwv/rz8Ouo
MHuJPVbgFpFXdJ0RZW5bS6F/Np1cgJVin2AyXJdXeI6VgVd9nUcDuKJn8mw43YA4JHd617i4NuwJ
n+QOqp3v0jC38nHuMSWOrs0nJtp92a9ANO23k4jnAtxzWudzr+UhHkUc9hEAxKm2jPk59hjDoiWc
SDbeCiPvANX6sx6SBXpXheUEw3gxtlLV1MTLv75egt27DMhYdnmjiqd1iYGCDzZlMRCWis3a9QEN
9YCR/K5b4UaK3a2mZZPJRp5goAg9coekkmlJorFq+1R2UKmgoNYxBaJb3Oj5dEyi3s8YjnxeSaP2
khEOwJOS0tuB1Ow50b1dE6Nr/JcW8DZXd+K3gMeqzOY9WLyUj5YtfTgfqP4cQqAk5u5SiXUqnzYx
xXkjF4ryC8jwFzSTbM7es877gkRnOJ2R5wZJOBy6fjNpxnl5gazAlG0oLrqyp3EPlB1uocKCYx8Y
f4HrK8iQexCkZF5t8HDDS/CDx7lvCZHsviLxpej57LhmFpJ97lThVVy/EahYarKEOQCaPEwIEsTL
pHOJ4F/796LE8DJrMhPg3CwNNVf6zSSHVBRbUHTc7wAE9GPTuYm0+KWF27fa2/2wgjkBvzsBllMf
uUc0S/0vM4eWwjvupViGZqRIixVuubEdqMzYUu3dfzVdMhE6jSUbPpMPSKvgbRw8zD5w5R16Q2e5
td960d5SJixviuWnFMdTVmai3WLct5/uFmGImZ+Z18pXZCNApLxHpA3ixtHdlMeNaHzkQaAiiQeG
JmPkNwD+CSgId3u7U+w1c3vMMsERMz+o+CxtJtuoZbJP12X5+X1jviUc+TJX0Tjp2/CjAIjqx3ju
4oKbtvtP1NbZUCsm6xxCnpz049hK1G3OgyUCNrijEOlF5P7k66QO7Xs12n+kOEPRVX2hHPL/YDgh
oCWf/LnG14M5a9jAEaqg3R+PAXnU0piL89ms1c6Hg3bbCM2S4mXIU6ivTwLAA2NTdgXOqG/ytyZu
tw6BjXGCKqX7jrzWL2kC//pffn3HXwYM5GuRHGGbN6HZt8xiVPoRphg9b/wsgmoKdlbiixlcKhV3
gCbpzGW9P/0cCEycXKxLOj2hTJ+amVVnROazLV6AIOhRT19dOgv5JQ8OmvhfxbYuctfc7RKzHtk+
KhiU1egFHu/gOG3NP2MOlacXgjCalbZhQUSBMFNXidlYziQW0+OQQe+xgHCeG5QolxbCjJp8wwjp
WCtgu5HIc89JQJ9bnVLhncZUAC5hxWroQZsWSPyZoX3jN/+GyZhkp4B0HpXaxFDtLp1amX1e31i8
GU2UsDOv8b9nwiwu9/T1/+enf6M8dd37Sf+6j+5t4xIODCcO7Wiqn+2Na8STCkSE662kxsF24pZn
aub6uEeTs3AcGXRiV1OSUYJiu/DfGMoeL6cqmS5t/KilMwRN+yJipZV9IJF/8b0ti3E14hIVtny9
TCYF0etnNCFPt+VAsHywAQmkY7cGvvpeKd1fLOabZp7k8nVNfiXgwJLklsdn9xWb+6Up1DLwHIZB
y1M7tiHKuBLygAuE088+gKOrnj5ZeUc3iX3Soo/8TC+J87uJy/tI1Zq+vzMBiLBI8HCbMs47dbp6
MlR5lbz2nU8ndiULcQRXzwE6gtX9wntk5kdkOtkwkxyylURq+4dhIIuR2AxTHtS+6mmSmlYNEF4G
ZssrOPZlfiIAA3sgm+Hpec5yl3K8HbVljc2UhL7rBmpsN8jR7nyjU8974Qdlq+4hxWCTl4Wk/sZ+
ESGFq60j3siKM8vXbjBTRc6/TRQiWYZzGX3GlRR34B3mj/l04oS6VydOFoGRyzfrWLxfKpWjZKEy
5IKkwFwBEs3ErvgKwgWGz+Rzdy5qcPbQdxtZGo5zUWiCIu3jv5OQ6Epgrx1GLs50QLAFM5IlyL3Z
JkS5azBhbQaVhFmi6Sv9vP1ntI3OwUkYfc6Yuzjx7916PFkMN+0zub6Frqq2HbN88vRy1eHc0t9f
ts8NI1Vn4WLH+tSU81Wy74/n0+uxSA+ju6u7P4JCdNIlsdeXUvEPoH0+tDKunYDTpC/9aPXn4lXp
gKv7fEd2XjW1/Fr1ZjlA3ptAsd7Ye/yyafvNkxpLTV1RncWLgfpSAN/Lkv8QIY6q9woolDrasjHq
oFCZepBSukrwOC5CAAC4gz+81I97TVDD13NSABcT4INW5S5H6/9ASWdpH6bEsHYSNuJAcsWKQ/zD
0VAkb6Yml2jGpjqal3e6RGVksD5NfP6L22aBhNJ1r//eq6j/v8ybyrb5rNDAd5tOLPAJ44Hha5xq
Wf+Fanf9iC3MuKbd6ma20o9K8Xq4RGn5Pvz9F+S6GHjvf5f2pRqUEQkP+Vx1z9WbpxTTzPtTGLgX
ZEkeOv263irWufeTjOotJtD8R29b3ARRTmHl9srS7aftKSvY/CQ0xEuxfROVIw3+fC31HK1msLhp
whxmN0xhL1cP8VB0DxIAskApK/t67t9ktvUG934RaHfUDySujY62W3Bw1aWDDXmHSJObSKA+6ycW
tiIiddwPeXRqC/GkvJn9x8bdxKA4lLIGh52Bl/XV2qOnc64IKA3E7eCIP3ipn+ekrsBa2pZ0ntCv
RQ5oi01pRYIlJMEOi5+YtUf505gGiOF0DkZWXcEUsmz6FHJzfiDqN5cpneEcUBXAHel+6ET8XwSE
G1KxkHFuN6x8dswP6y0w7qLFdM8Sxq+rBINluis3KPYaXKsojjrdOPOR3z7j1Vhh81wTbL3b4kUT
D4YZqusifk/8AFeThOQ1v2gYYG7V6ne32CPQZJOTpUtupYfjEYlqEkBdJ0tWiN7DsSEIiDSBNnG8
8NI3MiYEMmsKUSeq6SJ1v3GqUQbU2gjE8b4Cs/z6IXY1H21G0kVOBUchpE81O5MZQQjIs8a/DAXX
woDUlpjNljnQTaOuojaGis77LQLg6WUyGfmFIZAW3ZSm+betgKgKTaVVx3XBo5/B/JV/k/vKuMLc
7Tuf3bJF+9PuC6Am9Z+smrcD67pR0NjLv2vbgaodI3M8n+TMaH++IF2WBVlesoYeuM34KbuSLXLC
4PGeQPBh6fBY86ktx9N0t+qIF0wT91rjN5dMtWORiHVHl5DnydxbZCARXj7CIBxp3Piclax1PMpJ
koRJ/plBFTYDKkCQquFKoGpp6LfAc4lpebTHrXxYfbfKCu0ZJb/kRwlfshBKPQRay6Tk7HqErWd/
41Qv8aBvcZv1k5Si55pAhaJDj5WN031kKUK0iAuEUDPhpk523a+e2N+rFLBcS/FwY9mYBKG++L23
mHdWir+Q7b550F2QVxJF03n82WzdFsYMuTkgEjrV+TgYPg5niDUQxFDDsJC+3wgwxOhY2YbyVbrx
pVUfJmd/p5eQ6MCZPHbp06n9KCzKI9vmVelGF9ze0eGMDHuqoTtVglfb7p+PzJSvkzEt2dRUs0am
Yd19WlPYzG/7S2cz6ucNg7Bja6XgdMaPn3DwE8co5XtqWVHVmEqbcA3lQTsQffjxUzqspouZIBQ4
KweS7ezvm5DxpW4Ke5qO5ZsGeEIqQ5LAopw1ejLIRokKnvQkEHJOK578mxmZ0xIsfNqcyntW06JX
VxMauGjPIPCMDggHPsw/0NM9NWDeu/1DahTnB9hBNsXJd7q5nWudjUBh/yqTCSKvGnGy9CCNLYqD
aUo93YWKL6WcUYds/v/5rz8Tm499ugM34kGKqeBGYgxB8U5Vq7y8BZzOOgnFzczahWtvwKeVdEtq
sgv8OYcmx2UTNnt4ktZyY7oI90+XhWvUScEZYOuDH1JKxCTTD9OCXFHwtu6yhv6DnqXjthR0M6Q5
G8KiCZXgoUQfSw2JQxbvZxmEkPSuSKswILTHsO9ypLvmd7DaO0bLJ8IA7K0ImPPT9QhB4+bwG2as
9mBiDZJqDuIAuICPj0XGW5po7YUVMukN1de8VVH46J+BRZJxAg9qV3KRoQVEqB5QXaJ1qAWOCvsw
NfLWD79FWYTY9RZcrAVNVr/k0kvJEoBifRSZAz4DTwCiLGGiaOUS25rJ4NiMpr+HESOAMGz6OjZk
V03wtXGjnwjVuV/i7SFkBn35h0RYia1YjcnRlHG14fwbpyxf470guaw+/+ZsRZX0+eo8XUMjwMwP
856EQnT7duY0ez1RcNa9FicSyumVS1Fn1qes9NpvJumwIPoc4BAz+laDypNs29sh16dICJ8NM6a1
RYGkXa64/2sr0S/ePgeaCj5VsDdHxDIFlAg8SfMSbBxaqyuIIt4rnRULqBgesPXnpiN777UPGCqT
LG4uAi+SkBgnsFzRwH/y+leqZ0GKw+6jWPRTfJA5LE+NbroIHs9FKpY5Un2snDXdT/QmsZ8FO9dv
EROuJHS2yTGYt8dVj/r0PTl5cJBvoBUSP9LBFovHHNDbxuQpdRjdUemrpLjM3Rb2HsYh5FRYmjtW
PdWgUNZkjqmdSbvehO6jlFahb1/Gmqnsn8j2GfhyVtpi/eySvmg4L1hDTq4LcX9w7cjit0Gftwmf
skXsg5Kc6Wu+8T6Lfm01+CnstFNTj9s3ZmBkkeCJLbHlsqG9WnQtsjp6yk/F4EyEHdvbpitfvvXF
Dt10oEPK+/5lYM+U4+s/aFZH4jp6tKf3+CHQ8f6vpuIRcuV+0vRXTw706MWJC0n1Pya75svDu54j
xy+WZOkA/ol5qG/Tf9+9IQI1GM/8s6qp4qi8ndqdMiju94ZeSG+aEJ1P2xXPq/R7oc+GufYDckpM
7osIYotnb45pwpTh1n5/8/aeuhJ668o1UKsHgs8js//dZRhoCfPG6HAdkv4zc5ays9TR7evQHgsW
Q0zZfejdVRPi69B5Lmh1cWEk0pwan/ErehQQiJeBfN4HhyqYzSeL4pvwrM940hUNmXbWg5uaCnU1
xhHpW9b/rHExc85g7P3wJEFo3cFQ/XX8zAvz/cw6GcmtFQsfHoXVOuNIc3RI9FE2qiNo21H445bm
Uh76sBoO5HM/TOCEa8FBWFofnvee+uIKxp2/zYnzKSIvZPpl1kZf++iLAveTB3aKo9UijeGvsyZo
2pMikK4xC5PVlNFLI8FA7OIvtx2zyCgLHkWyIP5UnPHEXv1DK1glI+RoMXQni8ve/RgwZGDDocTx
cyYibtJl/fnntPeCW/Sv8ZklGuDo6mYFuDKzg6WqVZVBx30qqjP7mEgKj1D0TSfywFc3THQOV4H3
gx7dS5+ZnnBxU+JeOgzVVmVPK17Xkq98yrT+NEBVSg0tcmOf4leNcyYQkl52k9e4tungSSwkA8Hn
X3CB7IOehXkjXe3tbClt7JqFC6FALBK0lmRCfP+/eHWhAsojLd25s3mTdQeLysanu4h5Ur6VcSkx
R9i/sQFkrGg5cKFRUicTfBsP8+T6ueSPJleKEnFWRW19+avE3UUSs1xQiqHmcNyledKaa1YLp6J6
aw/kAnNB4KOtSoWiR7/eJXQzLBDyPaNQxf1U+MPJandZdE1KoCIT1djJllipXh1iR897y78voPQU
aJFxgRRkAB1jrdCw5sembf0JbDhtqhzomyD/aqx1mRRXN7prePq2qy3FmCrJ/McGiH5hxdgZApiZ
RKc2BQhYGwEXkXJwktseWmyJkK1Xlmm87Ccgoiegic6qvXwAFY9fkKcXZtipAAOumbixHlOpOHMK
/yj783eXdZ7Iq3J4paipZopgZoYkjeg8fiubnqupHhZBT+iK9oyettZsQbrKbChqesCIUZOTH4q2
AkbThildP39zHtJEof5X6ahn+bQQyZFkVSfEfAXycyMz9nvSzpgA02zz3+Xt70aqMsyBc7sEaRqP
mrP7ObAV5hCOx/Mq8YwZeXO20N/6oHn9o+QQGTBWVn9HwGURl1yMvJnXkeuzJFaAqdxo/NdZqVHM
QZNz4FW4Aem1HdPOGRlcerM0wzY5tkCzXZQe0JGpDYAV8xPvogNJ97K/9GlqcoqRXJo4ZWyYM+R9
4Kk+R1jXggJTZTg6igkaveXx4oR6JjVWT4cSc6OMiy7yl0hZ1578Wk8GlAUehcenFlkOY+joCjV4
ZIPtkJZMSONrag2IQKLsURmfb/MWyEhdqOUEzsT/am//Wix8QTVoJltuU+SJ5oW0W8XycRfLyISQ
2rHkxBThLliCM2m4o8nsdcpxq8hyDfW9fSQW5w22seYr7fnMfR78a3DU2qiJtb2iKmeOOi9w1C5z
xPFRJwxgZHYZOIyczrF/JIK/Wz53nYgqQMj55XvWKLulrDKERYbnfp1NX0eOOo3qPO7pvz+C5TdO
DzwgHegYfXLx/0fmItn1z0lK9YLAwi0sQniLKNmPoPzgCHP58wihbprOhKfSTDV7CZ5VLuEX1TRK
0D2jjqCJi9q3HCYc2Vn6skiMFof9Waka9bPhnhU9IK7S/w0xMFZ/ccZDQPflqt7x5fihRDtB/XR5
/tQbItIZCvUkZlDWEeA5KnJrQc+Krnq+IkDT9pYnjrRXWqLZB4VUN0rnWIvXdzR40/160Kiuf8Br
jQhCScW+a/y98+COK6IUiZmUAoTDKId4Rlkn+iXWrjaKH3ySqBK5jC7Y0xTCdUa4yRPcHkgF6OlH
XGefklq36/ER2KTrf6Sdjg/cEwAPFYUAiRaA26CCZU3m1z1dWRzxExlZiNr3I2RGCDa3WzumhfFz
/eTPDXDsx8aBghz1Fg+VOPt0jqXrhASkMzwgcgnLgTUVIZZjEdz4zQobuNcoFIXlowLq1rVk0JpV
UFp3kCUtd+qawpU5hjZXcoLAW2fiUuZfwfDMfX3gAF9bfSjhPWhxiTgxmYkWMPoesNjexzuJUmZv
zkO2MJcGj2rBUcALqEgKdXXlRlEHPD2HihL5hSIzjVuDIs4/zM5/ObmOXOcWTlVdfd/KiTJShuw4
5liGSVWAzpfAk/7jY+y9up0pQz0DvOMgCqWdnBlDEwzjLrQYCbheWBzcRN4wKo3/mBxQraOUKo2s
lRXDrL2XV3kJKBcE7v+k7LcfVE2Z/hdTGKNib/+91nEY428tDv8aaWxt49++N3hgNDVrNZ0ufbW3
gFlJLsuOWZwO9wwBgdO4gLqCXCTKBdpOKzExM9yhQD1XkDSJFr53MNJiGAx9YIM0TtGiRVTp0w+d
rSNI4Kwkkj/1ppxbQwdOmypMANBdDCcFNkYggZqnmj9Yl1R6+H8Z1vzHEkTT8vyTe/6CHHslpVqP
KhpwaZ/Ec2KNfi2eWqrP7KD8JbmrfbyIRMRpLU4O5JsrtCHOGlZugTgKt2JazG9RWODsRPae+Ws3
PExYL9rlKRF3nPI+kV1Y117kYkRjKDAxhRK29yXLnRoEey9NApXu8nHBR7FmRtM0bhFnJCQegFFC
vzBBUcXPvflsU8IgfJv0IQV94TosGUjqkRrN5EWawx9dFnXTHGtqaMwnG0CMZNn8uN5e4dDv/N7+
s5oj9GtJrNEeuGP81jteL64a+cFjc3mdINL1euabQKYENWInFZri5img8DY7IJHVvuooseQm4bfZ
AuWKrkDPDpBff+Su+8+C0xlpKhukUz1d4JnOuGzs493kUWmkyLQpzdkp2AoG6mo4ohqhexUSTMC0
D4rewytH6BHffd9m86/qPMz+eqsfyH2dNWJbcf3j7qVIZUp1ANkKotIycf6/8YRiStwqr37tqLsS
J3xC6ckjVBr17rq687UWQyRVVzJtwDmp+7s//u0pOyUjz0VlvGfBBo3uGhRCmZvyCTo5uh60Hisq
Iu9K8L5phmopbcm3AbDk9j+c0tJYG1dgjdgaxhbnCcHHZ8RIGnJ1KM6XjVaurS3e4qRC1wMt1w2k
qhItknZhGZ1R2VzOnQgWdVXi1A7p0Mow+2cFeLs1dP8+ijtQ5kZmOeecUzvPdYqPZbAgi+bbpq9L
aho2CRR92fT30qufCtMWEedR9pR+ULt9AhFO8fKv1gnhUh1CN3XMzkJf2ZkPW7egbEFDfeyFDE33
DEUuXoG60L3Cpg50SHvhqH3zoQ0C8eL5iXlKoo3G9dAMCnKn7Kqfzy8yzzIjiN9tz6uBCncaJxPe
FdTUhnijOjIQc/GJPp3W43xj6TcFmner5D4J5JQqtG9Uk6xkLzUbbKiHYCfgM6kkWwHyx2GOwZpu
rS82apKqmPGoznkgiI202OeagNDsfnK8WjBdAyXyYWfUkP4i2RL7oliBVVQ25ZHp96IgF9LnXEIH
dyPcJ7sIxP/w4MPUoEn70JDNyB9qWdulY6MEjz6zHsFeM5KJrXbXj3AhW+Yjs1EejKbEXxPnGHXN
7Vt5rI6EMGEFM0ZOGdqtZuelUfuJFU7BocjtLG4qCwGZ28DxDGT9E2SBEi/zNoxaIIj/q9R/aIPg
Hw0/GMKcHPeT4u7kGUUCcadIouj4bzMF2G/4ITgyhAG3s4uqrJBl2NoUSdO1erBQ+677vAEzmR9C
23HYkiqAZfTWYMpNOU8JDXB/Mu9iVpMrWQhHgikl0pvdM+P/IScpLNwL8IbeYjTx7XkUmSHMbQKE
RDTaWJ+XsWvQvInZ15U52vVjgcBblMhJ4aw9+ElWvvbneiKz8cVaZWlgVL3xjEghRDizydnqQudj
/ABQYbUCtGXUK6FNlZzYV9liX3Tf/JcP0wLIiCYSTcCdLiM+WRk0TLEIquiUeLWjcoq9ltz49WrX
2AeX0g7RNzcoqVFiRCi4vU9/nGN4rdjs+HkHa38S9Vw42HJZieRSP9zid3vz6bnr1O7zIkJVzsfO
fl1OWGZdSaCkBG7WzaSecLRdUsX8uUbZcLvWwTzFVtfgyeWu5M2xX8H2+MjTajrlSXefex2sen/t
craTVtZSj2bcamD9gj8H33l1os8G5eYcDBCQeEi2+sC2xD0lhNtFZswn2R20rcsx1DRYWqcdw9S2
EmRcMdSOr6bYdtPKJWKOfagDOsqCMrGOxmHUSuFwz6rCOh/3SuT1rQZQT7CgNr+Rdgfvhu9Y+5VP
zmTEFWI0Yk6ZYHahgBgJnkN2QmTGZFReRm1E9pSChDYjaqzzIAse1IXI9FSuN+KaL+7o/jUoeroV
+7JThh3WyJGhJzL5JFMTjXZ/tXUBlgQkjiuER7JmzzOgQVXh07N/xCcGwg2tfU031ldb9gcNKp6p
eBt9Or1ph0JcduY8M+WzxMPLCb5RA6vq4s/4IMuR5Cjy2GEwc720Nlx7JHeQ8FJouCpzZX88UeTQ
V+bd8k0HQLrWGPlGStTz2Ll/JnzBzKdXeTXrMpQD3cnZY/WeVRBNQCRDDSJv2csOKRA9M8Q5aegB
phkuylJkbzfAFjk7ReDmz2+2EMwhqbuPKa8qyGAYSXgZJzXV9GTcToBbGkCjjSOZJxL06nvVJElU
Rvq7qqYefYIzFJaEd9+THLHYRKx7vyz0VfPjjPgm8ofyC0vsPkhjvhtIrzOrdfJNPv6peLQ3vtxd
+bsL7PfpJrAi4GJkaSty6LPJEuijkH6SJnlpR32PJNzowdRofz4e3zp0JTnz/ZVj193mbPy6WIy8
FVP8VENw4e044dV6RyeZRfrdycogNburHsCqpDfKmArK7ToLyVZcN+u1zSyAkNoKwXzxukhTQAV+
qvWdeKmVDHalLg/egmkl3ErvOvu3KBwaxXSyyGRbN+eQIW2Ghukg7FfZFZJu/2UsP8aAjt/bS/Pv
YmENbBvTlGWwtLiaevS5M+MO1Ntjvd9oR46dYEKbBfTYxaqVJD1SgZ8H71+obDpE+AH71Q7offfj
mJwO9Ve/IBBXIjsLWkeOjFjvIjXpMb3gWy4s96p2qa+w64En+ifFi9q9qlx+YynoHqK7gpJuVAMV
PisgiLsHsdS0ysZ2/2JV5mh6TfPJ9FBKR41hVVw62MT28aQCmaSZ0oyFPCf6bTDKfyxqvuqAmQm7
rscL9Pj26Kbd6wIEPpGSHJCvhOi8fJY3h8wr9pwjkc8KjmoyZWW8f1fa589V65NOFONBtEfbzjVQ
6gC7a68ytC2UNVnY7hejl1TSqZQK3G00k/RNVbFCd8lhY/0TPxyI6405+DZ4yTZn/hAX2s8wuV8C
LoZG7CzgnKsTqrhnyN9VWG3J+L/Zk1/i7e46SGnNNEcKieC9wWIM93+fDb+fWh40jMZN3msEzl+D
fxcvfbcwKPQOTONUlS4ci4envFhLgxi9FPDg0R0ouDQXUCI8sOZibUOhK0JjlQInEs8PGJwnwjtd
chj0hcrjgq1DDaM5MkCJZgW3tYw4CfSMGAm4/xOaVOfTNfeKMFUzukh243kDxhiWd2sO+Dv9JoMB
1SPQvzyCccoq91CJDge9ZR8XhLwL4Sj+84Qpj8FAM0B9gqBQboxMrzHofAYihGth6QOwbj3IZEIz
6Oce1ZLAHZ6gc3tPKAJo+W1qtl4o2rm4hkZv4WLnjknZvK01Vg75Qy9ORyoIF7wkVU+buy/Dd7ii
N/hdTbEWTXWG+IElCu2UNMA2asXI+eCSMujqMDx62/rPIHsCorNATOGgMJGwgxFOtGtXEQ2npKIC
T4HrCB7rv4GzO9ERwNaaPqUR4Bs2bwFEZb5sVyKcSjfPobeOAV/L4cN0Jy9fp9N1uYGjN4hY6eNU
GIIvHci3ePa8hf99VflWsmPaxnVHcFY24ri4nil4yAM7U3qobjfEwgtsvW1eK8xu95r0YH/1VjMx
nx+/lxq4MgWaYMejLPdvNDdxi+YwEnzXXJEsc2h2dTdher2hSl3120X2Hoy7J4ajVHmCUCgWVOiw
2zjLCyM08tiuzZBZwz0MKX9J2N/izHWHNEhilumKC01rSqHe32N8udD89FxbyoFpGjBfp7VflKuw
tsACWg9RPloLQum+WVmEMDVf7fGLEbsNWylTP25m7lQqVjjpaYVl/g6XfOHL72BzoRiB9Zseyjza
bSsvvqk+DBJi2sZ/civT/Fg+9HOhHfEJxIGUSbVioaHmjc95+Dulo3Hqe+/RVCgGdC0uRlFrTqkV
i9LC+5Bjbe41n7n0AFMwVS+Ko3e1jqJF7tShcQX/3u9UbvTvi1fLpCi3B+BkrS0a48sAtIdp7VlG
yfzVE6n/lXzDTWqzoZceXDChMg8zxdClnPaqbh7SOG7S1B93m6h2jRYOh5e52VYRTzMvBWxn52h6
n6uYtTRll/YHb6T4vaQyYby08M6am+rJqOdYsUmEYCQqxRBXVRnqWJa9ouELVGx9scpCNmgzOJmH
BNDew43MVuwTHmnT4eZA5X+xrzk69PX6J6sYzgw6R8GM63RVpIlcLg7LXZMWX0ZGEp6b4O8a1etI
yF1X+A8j3wHHY6wmp0cLE2/A/A1fH2m9lnWZaj4StF/I4oGoFS5oTMBFQzo6SLaMUQu7et+dVwW+
3Y2StadbCmGy2cEY/em1+0R3bWQuWA4QwLKo3aVq1sqMjJsDRmKp+kSNozW8g58ZOvGxkQTrVZNy
7DY0uUon4PW0aZw+DViDuFXybzDNjyvHCq0w9EBjs10i+Qcs+Kc5KVK+V/K+nFUF2oDILJFjtv4+
fZmqLXI2x//6ucon5Gt4c3RaHv+hbVgTs0MtQ8xijH5qLTrgw1+qiD5VT64DoVaZRwfm96Cf7mcz
awJ7Hl9K+6HSQaA8E+0tCiAZqVZ8IMEn1tPMNrHEBwFHmckkzZU54Y3CjvLaDwgGHJAv1spw3Yo4
qj4lLIh0wFNleMgaSVtAd8M6WUs1qqqCTRi4siQWQTBMHCfnCPYs7s3RFeVV6Vb202Z0ivcxCPGV
J1vVQgFoMxgcr+P/YuoTHqvRkcy49Zwgcsy8fWlz8LiKKW0f1Z22blhTsukzVD3qjbIlBnn+ADp1
QKOrlLwT3i+jRNdQZACOrTqN/x3cVohBRcIgZsPANj033cJF3ASscOxOnz+iVJ2X6j+JDEjjA46M
TFhPDYsX85i8BYM95Udel8T6SAQeFJhf76ZIquD/A7FtN4M3OwiuNoQMdEc2JXqFFltD4lfFAlJJ
AGqfy7Ypmw9NXDA0/J9wQa577Oxex1AzA8/+fQcFna66n1kLIKjURboZMBuU0W/qI/wJJmYtNkuE
XxbQPNdBTPwoAA7vnhFAlkSSXiqEiXeTp8hmvnetv7ueCqM85qs0f/l//4N52JRg3eNZ0VivUbxb
rJv5o9YfjJ69zvEFIEd37l63c5qL2Yt3yCFuSqFvyy1bZuntlLAamXr9EyHc0X/Lb+1PD+lumhaV
wPFvMCtgJeww/MZls8R/cRCtZR7lKLiX04LD9xcMrjS6zRPt1VrUUc8Lw4atp8hxskp+RCdkbk3M
vMs+svvYVU/a4jqm2+UYJO0rfnb7dJK0qpumoEM9hvJZy2o7ModKoHXbq6sm9O6d93DBPHzVm1kC
d/UdREUOgLyruCgWkQZbQEUyRJz1cHs/kFKFp8MyqD6NNHpMxIMhHKXI2+xCRRlzpbxUC9JWx8S7
JGB2/65tJHYq359AjgQS5nBZk9c38Lh8IeFg/prpz1UK4o3zwtWY0/Y1GezF9mwpRrTyifuOETr9
h3xEngtnekULCp/inUAC0NIYLZBeUstaTAtaFQ11VXptjZy8QDhzkeML+sjATuqlyu7jvF7HWE8b
3hT7Qfa4GJ5MJZh3gvrrQ1+0xBZ+Say2mSjdhrBGk2SGjXxyyrbiOImsGkaDxsyXr2mcnA8YPBw+
OTyiBJQITQ2TG7gIfT2iH2biW1LejUMupb4Wl+ZqFlAxfiY0dgzWPoX+GL41tFAgEvX9nhWGaNbX
BtVA56zai1n+4xBIf+czAxxXq3MYSI1qiS/l62g+MjEdtrKSgJy1yYPoSjTC22hDCQF0+sCB9g+A
UiZfYUU4PzrYMAxBXMm2Y8eiUYOYmWi01GU5fgCcUwf1CaFzOk5bZYu7Otm68iUuRfTMGx6S54zh
7v/qXExsGtQvm/mL4DIJxzpEEEULLGPrVoQ0L690ID2mq8Ar2QoAnf0gBK3e/H1vdBFjn3BhSgB/
7hEfkYS3wstVw6jfFx7vGVMewHfSe1Cp5q8Qh00NRIGc4ehH5ThEH+6eKk9fVcOoKY49l4HLYUKi
fXNGQJttZRrJtI/L1vacwC6Y+UJo0AjTjkLBleMDZn2WqDKNABDqOY///eLQSa32tZETVtv2t/vI
CYy+YLEChyM7zzo5SVqLRPEm7nVI5WcV9Xh9kK03OUELbJAVlHY4HXiUWfC8bocDLl96uI8Oa+ya
NxFiFsGUYEvhgH88qKOdT2lupTf4S0Z45FOzoYQvn3cnq05jGgBjwbh8DeBEkGZPBAek7cpSfzVP
IfrXWNySO9FozpQOYJ9DFxLrTK9agB1YeABGcafIj4SZD051Z6YO1OC8CneDAnYMp44L+g+9gfrb
80Sr+eY4K9bkjFQjirHrFH79HKHJCnsvClYTTmPZI51uSvxbfBjrf/zZ9pQ5SPk0qe8TjpSOSGYJ
NUd8TJ+gYPp7ReJZjysEpWjPBHjuWgwQmWDiKzthVqPDcCitFMz8Nhq2IXgxXY6R9MFkx6hqv4li
XU30j3BVsxVxGeu3RIW2GOuQrpBlRZp44pLx05zPp/nIUDRv+/YeGehVwgL/X1rM36ZXhPj/fej5
jmRru8S9IdzLpJ/iHXggHSPgrwc8bpEEQWiChO5yaGGsxtAE6Kl7ccSlGlVcQ9617obTVdtq0Slv
yQU4vneakDlod7D+XU7EN/g7e5hV1Ee0H9BwUdO0yf1mcOrluVzCaXj+fKBYcruoKSJONzDwC7Yk
76sKlPhZFcFEg38Z+e85mJz+J3XPgZw61O7+B1HFjkUeNuqDe8UD8hyrJb4kOxHB7MI1wFOcuwQT
8CegovoJzLS/Erw5Tdlkd63fqUopGDeP7JFt6ML4ee6rATMh63N/H6DsLuGDabWdJ4/fFhanjKNa
ypGIf5dhtrzgE65ympuv9vYS5cbtiypOyo1q4PFPSnVBCFwmSIWeUIL1U4x+k2GNKEULF7DzoV5F
ijuk65apgTwSqGJWP3Km1rTvIHc6K0wz30EAMUNY56hPnEf18EV/2vaI/IiUtyDEoE1qPdIOUABU
j8zfRuY3CbvsleREf4W3qbA2Ln/7EsPfnD3eg7O3EUlukx4hs87OYRvl0OU5snmPU63JSlxL8CWB
yl+lGGCjSKt1GrzsZmnXCrYTK4IJRpvg6nMZ0ONhNnJM9vXpURSo2St2jacvPnr7cVoIyQv1GAGU
hFLxJ1ShBrPuBidF5v2ApzVv+cuxbOnWS0ZvwiC3Did7qch6xw6viTFo28/PMpa5a9StTsZR/oKO
tdwjq4gHDGhxN/EHQdl0h9DRYmRZmrwdOlvyvOl7pnGNQbJLcdFwQV1IntS4L4wY5NQdyi89uh5p
4FvblW7r7Ti3VOHV9+NVQRWaEbulCIrL8wfI7Xf1ihKhkpMnX0NQwl6uJoJmciYDa95FS8DKjIZu
lhBbCHJaWrJAkTQYiBURPdZKIcY5KBg+0akxlDo9GPYtVtRzLhvN+N1KKFqjI0ab34J9yqbJ+QxY
aRlLRY08FEuEgfK4oGLH1Ikib0vA3phDx/UJ3WxcU0hN7gB+KmVSEkIFbQoRPX8myQXJXNcj4Y0u
ZzyYHmkyfqWELqbcr8WC9m6vjS7RhT2qUXvZqR3X3FeMFsmKUULmjNLA6a7i0oMLW2OFAg60xvx7
3nUOwEYLYQIONx+BMOXB+Q41Tf6/wa8hix17NJG7E5cP553Ch9xD+Q7rQ7H0wbYNh92iUd6E2m1K
wB5KRJ32rkaFa90mxiOKyadzroenk1vw5yt4lFeXIcGKbsNc4JaJCVh3KfsgKBC8ThqTb7fWbRJu
h6XtDBD9ujcKLapR12prYVmVe7jvZ1YP6MBGmGD7dSckrQryF/1nKNQVB7Gw9T0zsg/YtU9AlifF
H88AxH96q36N71MqsRwEAsKBb8Ct0qUMhNxWns0nfZtLdFtXpAhgMdbAuzAd+QGiCfte3Hp26SQB
jd/ui2SejbU3OYhBmLW6/WNbCHdV3/SLNMW4CX0asN1xWGjm5WCrE+ZIwrk1Cnag5M+oIIIx62Ug
HpAqSUFEGB8gPilcDDi6i/gM0ahzexyUH7WzehZddlJp13PtXzOq5cSI+cHpZnJthZlUThl5rymx
YslVddPJk0ic/JDTFkXFNNQiv5uc+mIRGAM6koRRBORgo+bmq4dlhjMgNj6dAFIfmy+35N1Ag+2l
5ZDenyRDYk9kAFiMBajKi5VI9mS8fJfnjHHMqH141XFzkUmd4fj5HQjQvlrsi2hFJmLvXBBUuru5
/KhwjMALtiPweLmAERK9OZa8qT4R1WRL4IbzrpderYSRKRTkJbBq6+qo8vkqyJNuectSi2iCXQ9p
EIxoRnfGFnSqCWBM7P1RreAGPq7NV1fKpMvshV1Dr8ESdhZ9vV7lU+ip2CsnIY1oiKNP8x61bUcC
TO7m+5DKIUtfBuYcST/XipsXLrBA/R1+aVjiRK1ilJQiN4f2zvYj55h1BI5E9RDYkyriyhWlnMBC
gNWwSvhiPNx8x75Rv5IS33gtQasCP1DpsjZfE7WnLkpX8trDT96hXiT7M0hUqIfiAUU8SmOU6am7
ulI6005s108gnD32JdeyMeznK4YVUSyrxnPbF5duM/Vy/M5xV4FVmbUjLEqOMe31kV0qYNkhNQ+W
kuFgX5caRuMAkv68LBda1TxUpQR+9bZu3EhbdgP3UDmTZH3rRIe086qSJKfi0uzPg9eACtgtU18N
Zj0+tXUZYv6XiSObbbNep+aAAqHzptMv739yxuoG8KZ3hmZpiUiAYKAvBU8rm/WjdGgN4go+l9mv
FWF3Pll8ENiq25b3Nl5emYDqGbJLDRF7hegAbu3NXjUOu4LEeJ6NBQBcgpysND5i9SzsmcqGGD3Q
1yKjY2uz6xuXQFdf7zq9qcY/XNTcGHJf/YK01d7nwRG/7YaDPCeUgFQM2qi8mRq6zYJ9eHp5GaRN
ueNHRalp+zY1rQLQkC6iexJ/a19qrzYE0te/EJWMxfM3pU05wod3dQRdcSDRg6beyTgvaQeGB7k9
+7waCAQZ3jVP45Bl1eOlYQxdv19pR/oC0aQmfZXluBRW08Tq3bX2jSWucfpTizxD4fJa3Kyp+24f
bOWHPL9Y0nfdlMLYZX3D8sbuNLAvPe0cIJgTD7LsyQxESoMnmXjBpgkBkRDodn0DgYFN8V17/dMB
GNUpnP4Ta2dwSLjiTFQbam0Ohx9X7Gkvm9sUS38mJ/9TU6c+tUG/gg/J4njtDckVXyqUM55z7ifX
Ep9Zzn+JLcJWujAXG2brdOnHb5nzseQ8I/HhvszQs8RA+bsPlXVRHN+gBSV0EpNm6RQzkA//bmQV
tUfpkR03AokT+9lLjbRD1IyOV5T+oJgWRqac7D7NHNYOvnNHDmw06LJSqPzSFnRqjzcUiRQsMRgj
59vYWZBNeeEHOSVBfa0T8lkLkSRry7tRak5QK8UOF5WOVRt9/46gwMwhO+jRpVX47GlkU2s/l5XI
5erruOOo63B2jmX0DtLBg1h9pQfYXTd/tM1410Wa2JNNK4e2yLWrmaVc6mUbCrC+HcI9FAACXl0i
WCvKT6BkVwfPqNHL1PKkrvUXuDwU/8WI/rodXnLRLMxmSwl3UM2pBD1v9pvZZC0VA0xFutmYOXJp
GqYvpCIW5g0Z6uprHE0rP1Cto0xZsOyHah/FZLE91JNT7rb2yiOJ8NkbostGFPsoz640n6nU2VZR
iEgcVoOOZXatgzkXLb+2qkZiL1FyKxVtZSYCrbGJC+hEbotxJQ0DA62SC2Yi1lyfgsbU1IUAc1ZK
TksfsIOuG88ZbDZ8lcQptfwGV1GP8aOUPFYLgWjVt9KcRXRcguBPm5cYBOnPafsYsDWR/y8tWyff
XjEVqBCMwq04YdlEYvHHV8k2KDB6X1MX2vpxyGOLdL2Smr5F62w7KN3caIl56nyHu+gk+Y6wB5Xt
0ua1qXshbwhFVvjLMXYgQIz8vqxN/vvPPifRAbNKLq3zBdFeuVbsUe+OnmyWSiJHpcffYiuuKVKX
/dVOP9p3S7el+Ck5vJKO1xPsq8XKC0JIPBaGoCXfFEsgAnm0563cK2tbClJ82B6qK/PtDVrHIw/L
SNrIgVN6A628PQxzmKPacS4uxhUlQNDAWjosr4Vw/LQ7b7FoG55AlFhjhiP2dDifOQcrzQEIWONm
g+xVer2jTd12E/I18Ez/Wp+jc1qxINP4izvV0c/wnMpYmJDzi6P8hd/5eFj+8NGucQNhLcHHzWDt
djXmj+o+jEZ/MtghE0xQBAP7HJHu+BJ2GhzJt9XAmcBqIu8YWTUy8xya9S3v+voQBBYKdaYALJoM
/QuNw1hSlsmuapjF14K2dWSiFinERafMITb0Gm5fvKTXhaT/cNmFOfZV84OD1HrF/yCtbpaIQems
BQrWOxa16k3+WdlWgfqPxmwGhKfvauph/ITxv3zMP1wbiYYzJGrxlWkj8JlKDERxA00HTGXHc8qZ
VBi7GAZzDtUl75a9e2Hyj4ZtUrYv5k70RdO3st93Fr3s5MYfMGMKXKJw+mcWpOFKqU0LjSqjHWYU
QSfuv1cGio82ZNqM4jIwCOHDsVcI+cA4djWH+43Kc0BnZtNpfeA+ehYn0ANJsTZTMB/d5DBxABoe
KNnZ1c9rr9NPLIVHYWCJtlQNAORQRV55St5WGd8jiIZBY5wJ7eCSWyyEB6m+GvpUmV8cd9Nuhq0w
oKALBcA7E1j950D1abvNTfgk6K7L1MpvCP/w9mBgeWa4UIqkMnVR14ReTGs3zUHV0vDDQcr/cbE1
6RHLmbpdOYf6FUr9MyzMk1lW+abJ+JlBp/xe8HNBsIzSHiVC93QfsQ9rmlXlkHeWqEViFtFZJnfn
egTaImXpPRczqyVGlZb0Z4ri4IIFhb1o1wwsr3ZnDzFHGAGONOD1P1SLroimHDIOPqU/wkdm/kQW
mSAyF/z0FScauwz7uRhQ+nkFDZKw/SG2Aq25Vwr2I6V3oFdC8ld0fpiWYWyauM+liq30q0cc2gTz
3o6wWsTP8kjgHL2TIqaa8ocUY0GwvRlDZ7eavLlRdEK1+ni7J25DzCMi9Y61okoA4HHl5zuRAofl
9qssokSsA1ocsnsItglf5aEm5z1YUGrkyAICT9LkRE7vzNGyKUlydTRxhzuWyB0A3qwkR6eXclH7
KYigVcWEk8WZbYlJxmAq479/rIZqo2Gb5eTaBTwVnWEWaRmJ94WtvcWCWQe45bVy05PiMbC15UxT
ktv7Cosea0BICnq+EM7mqTrlQobHYHqmBZ3EKzJaobzTRzb43cWyqwlK97bRlCM3AgbCNS2Y7+OV
cfMpY81nQCpKIp8qtZnGW7y96BTeLgqJTnmh7RyLy4tQgUtfDNXZowC94/8xHi2apXLNdamGXqrV
MjHlZj+D2hhlK7xTLZXOlDF9AcCSzmhlZ8H+OPJh5mdw7YFg+ha/iT6+FvJL90HCPho+kWA9x8ja
g1P1a4PZRT4keBK+5ng5Tkpv8U76YBKhr3ZCUKKLTRZcJYriO2UEXguhN3WMCdzakNZEE7T3uvH2
x9vM/E0SkebwkTOScV14dOdEShW236/9CyA9KJ0mmkyX+kMaM2i+XwJPY21fVKSWiL/4HkNXl/fF
+cemBR7Wj/AtfZIdj/M0qieskBPE+m6Ylrh3Gf5r7cEgyQx5DmuY3n5MFjxkropxF/BVMvww3PyX
SA62fHw9wiyeQCWzgiMpQjV2Oq5/Go2fBreRWsgXO/fbjP99vCEfk2zz0Li2rUt0F7Et7lcUdIma
+W8GTkimtKTybN3Q7taVO3EosyvASjuZHozpeTxAHYfbS4iUfqfB9YkbboXZT+m3EWwIQlMFRM52
kGu91/4jvAf34KkEiWHanYBJdDreBZe6eMOuiAw0aNnVnbUG3BMLPAxsxoFPzx1kG3aH2mIjzqzb
ThkV9DznfcOs8pLXQFUw744m4IrXKStCv86fFlF8nyABwzxBxRACbMJQwuwFx58SiZWB1xK67m/d
c5MDGBZJ4J7vdH4upIMnEzuVCg87xX3W3WvC2H3869Aj07iT7Eto6Ju/ETrp03fkhH+cQnOE5g4u
QCeSnB6vRhSb1Yld9zDA4Lyw9d5u29obzJT5lRW9HGq7QGP/HagbLLklvTRCLy4+HsN4g/+0aQEO
rup4NAiLZfGLzmfC4fJVPk9h9LD2Ch7vaf45+/S2q5VGIBBqzm8AyDMiesOGxG63e3a1Z2fULia1
zrq+8XNNb/8wYDbgnLgbUXmJ+Usw7ntSholHvir0Plx+PfYATCu5toNGNiQvY67EcSfh0kL5ec31
k3BFsqylOp/ohBwm2BSECNBUlD5ft6Jjgl1fbcb8k3I0gr0xd9eYj+eIVUvi83Dk3dOmSh8tCcoQ
ugv1cL9G/HeD+L01RaNfR5Yib2MZY9SRrFjfvYu8uPcIujl3E+B3aUIC2nodI7DGjFDInqt8nzbK
areqCFidvc9VMwCeY8DB80qyuXrQl8N30HX5LkBIJ+k7yMh8CR4srVKAMD692458ON1Je7equQ7Z
T44SkXkRZGXErBEgglmMTYG1pcQN7cEbY42A7sMcd556tRo6AR7VquoGTxkxKgeGZL+88I4O/sIR
jdYgm0mYQ7/77CEnPUckLcXBxWNj3eLrD1d7nOaAG82/X1cTKVvSTRXTZ/dpGd7DFpSAgi7VolqC
A6nN+NmlC9P0t+XI/2A6P782X+jVRXyAtT1qCneImbUMkvXk7MyIxV7Bt9Gn18pp7ImZ64rbQBLj
AyniEVrIuMNclwvePDQBkS6+8LYMIIk8dB99ZXys6I40ViZfc7FWtbWxOZA+Yicr4gVu978emoaN
MP7J1yqR0byN91Fp02EniCu1EKUdyv9P0JAdyX8NjCN11zSWwtTAOrxXz4a87O3Dv/uZ1Jf6NzTf
8g5l4aVgpQIDsacNXS2maa7/V4ICkUx2gMGSiHRa7Cn+c2/JoXiUjiBk1YjHBGqjKqhH6WkiLPJZ
/S5KCKG3guZa/5Vq5t/ngbJqOwWR79KPtZ+BxyedzMYP0nRy0AsPghMj3FWFCPIUS271/eo5ddET
96gyKtoCeq13ur4HadJuWOPqdBITLTt2WnODZHIoyLzZqBLjMXCYzDu+CBWRXrCcveI4p7wQMCRA
YqQMtQcMqMGHbtdd8JwV/Kz60+3qYujOOmBTFGCpfcL2uVGtK4XUiaCkzN3NvSZjn2aM5WvQqLQw
DVH3y5XCKxQE6Yg+mzl/2TYxR6I5Vy6741AReP3WO1GkttFmze//4oETvsykDZ1koUmBITpZhJ3Y
57yyLYq8VRrHHxystY9mCWFlL45TD+roc/gJVYzB/xKwQgWSo921Sv5b49dlGlDPA/U1h7IBLelo
HHk6f8XBvk0uUSSw+MxHV9/D6xzbckTwq+hlJeroGpCEykofiq6Wlu4K4FseFL4PG/P5RXiTWEQS
uNMNUK1cztngRnlo0MHfvVAp0c1v0ThtFp7QnLPVyOWx4tIvUGmMk6Puvgsd2d4KhN2QL6QHfbmC
IDnsG5WnMulaNZudl5aqXKEOgpNsj//sCDZSyIkxRliMI1o/COvBREBmtoktyvxg7OSbi9sZdM8B
AckkoUkCDfkHV6/9dzMP09nrjSEhf+xjsB+mY1gtEOTInVbQifoXX2spTNyZEVBeMbSE6TyQBQ3G
sQy2cUEGbQV19UCMyb06ioApz8jnkXnzkEqAVAHUTRTbN8W3U+BjmvpdnxIbIX+ykzWE0bH87Gwc
4v8gzL34NXcHVvc9C8F1TCmqjuyoqhzZwNSpcdD27QEQRRNd/QQ3DHKLd/xiMbqNTjtWKddEcAMm
Eq0ChyO+zgTwc1oi+b0WB0DgktVtTZsECX32yA8sGoxWCVfS3UIxwwvzj0077/BAv3UU9Q9i4m1C
ZQXKGe5/xiXwdx6ck+efiigDrL3A/+fbUNr6NHt0FAzdHEqWO97t3s0E5H+otywhPcHAWgJH8rL8
Gkjkpdc2GTGIKmD/KsHYboGPPQv7vk14aGMe4WFWo4kO9Ef+pREo+REluKwvOdbK8EYOsoEm9Ymd
E7H2PzibPwpFjBAtt+W5FpMGXWvropkDSbvAwcMwAv0wTUNmBwat6n9UtYK4jnlwTMB/xXpPkKoV
LBU/7c3vlFtSh1AA9t1Sp7iK0ELbnpDwnK3exD8agRQ+lDNzE+yl2FEt/PA9Wdrg5dkdxYJiB2Ns
26Pt8G+xWuInU+TMjXhZApRA1dF2VoMC8ATqk/NyDGwXbOwUuNrGBRmsyj5eQZHAf7zxvKWClSgi
sr8MxKbaC/oy5HnkybFVai7wEYX0NsyoOCmbd97y06JeahCQfvrg2XdniLc48fiv4Zt4NUNfnR8V
b+90Z9giDkkBE4UOnhccoEemnhq3Z4H5iJnfvpwAR6qBDRixKjjy1/Ijtt2mTAH7rqvOcUJMy9/L
jZFnDgTmoM0OQx3oOPEaUfyXuo1s3fVxm8EY/45aW+T77J3xaIJt0M+WAErHfNK2I/pXx6vWjRVH
1Z9BUT/ZhvvYlxry1Jimma1QmNNf8pqpCkVZrmpPoVn9xaLEVze7nxHqXqtyoPBDdS4Ain4w3ulo
zcFu+CnL4o4rv9IyochjXj4ux6pvIp2W3bf6R6KvD9zAabV7oBARLu2yOcGvCK62WM7SjkkRXAND
+aKOk0mZbFPI0uJatCIxS+dXbwz0sWISF196a1L5BMdJGNKt7AVjwepFwitzxx5u869UknFrmEvI
/0QNoXLTX/2HvmZwtceCH5tRabTUj/uGkX/NRR5U/WI+kkgyeyLbVxtdVGzsD+PzLmqavgIv8sWF
20KTkjN3OWJhJd7y3cR5hRIi2kZ7s926qKr6Sb/19HjXLohWA0X19Lycyu2PmJQVTfJQ9xen3QIo
tHcPXesVdxAD9Z0CXF3yqZP8uEYxKn2FUQ68tnS+S+cAYips1ihAaw0omc/8w6qROweHnc963x+w
hTRtrGu5DW2GAn4FoiLkHbfQl8vuT0N+ps1XVrfjxZQ0tq7CK5GY62z0QIsKpsK+ojCaZBdcK7IK
uhHu2fKF8S6eXhXepBxPfaIKhFD2zU23rvsbwKpcuH6PZAWn43BlQreNU5t41BxdW+CE0LMvP2SX
S/daICQtt8Faas0n2uPfot0wL3s6mi3ZxEEVO+9A6w8Y2F3fGKCkO0mHW3eUGQhLPjmUMYVf2hdr
cW6iTCmqOe1EDTZyzJyYLM4JfPcoHOZ3NxrGz5ev/iD8uDwYXC8OW/hoFrVm7/rMrKqDzveT6tV8
CtTydZ8aGwBdsvUv2cbghyqBndbT92ye14mwNAAEkUlMFIFARCoQlbZcGzU14o7W5DB8I6evlJ3l
80Cl3fI+N+b9VIi50vXcL+CnZXQtcHlQT3zy4R1Mn9gdqoYvh59bGRaxYFy0gQozH/BKyp7wMKKd
cGZbMhuB+vpXoHZVjHqtIm9MRYPkz/jsfbqAPnZn/h0c5pHqUE8swTaKeawiYJ0uDtFwsbsX6MwV
bywhXuFPikt1KaIyz3p/PoGz/ctQqQ8OBdLVLvd9I7SM0jpJ5A9ldz0aqFqE6jz84vw1pwjJBxt7
7F9XoTdfI3ER/N2VCiI0n0SVSYBNTSM04Q6AudZtMTQ4grGB6vHKP+XZlopdFEwSgm/iytfJhCXw
1EiC2L7XWi2j83rwTmTCGBuhPEOpTh+ssx9hX2aduJbh4UTWeJ2sqM3DASqMiZwS8WfmQnkwjFBy
AtcXUGj+Abz59+zlrpRJgy6lENjLsv55mKkGOjkzjSgX8+BLMgEhxeB1j5t7Z+ALJJkkLb/eMcTQ
69WBvqurTZJ22BI8WbNxhjuqM4KQPxFFysZrzq0U9nOZzUzLcFE7dE8Ao6ga/wF6fON8j8yJsRNq
mrcxqgDU4FJ0rBofLTaBKJnnxl87aF1SbzWaF6ZRhzIuZEBgflhVpgbWVtA1f09TEpdHvyCFnjsv
qpZ2+KNQAnwf1H9KnaUq5MISDSei+XUNExrtUaFDkJ7VY5C+/6VPpY3J0tdkIbyGcDfX3il5od3k
xj1e3CSC8g1h0IeY+wglpmkr6ee9/UN7/fDaEPmZ692/Uhh2P2pH0Y5j/gek4uwpjRxF8M56WsQK
COEGvc0HiWcXGgwuqtOMLvHXWSUCe/Ad/pPIU8X7GAGSJACfzD3zB68XOqq0Qa0sGtCFHi5tEB36
DDys50JpNN29/9mKxD75hrkgRnfmpNIE9xCE9GeAn/+zJh+s/W2jwpLLX/bGWiPS4rAWEoSAqm5u
BNtt+r6ay4Aqv0KayXIwrLyONqLe4JG4xdjL4y2r74woI16H6ffnNn5CyT0e+/1rk/8bQcYfoLGh
jaT1u/xxva48Htcl97MYypZnBBhS/ZT0fyw6h/53oJMLMn8TRuJULwC6YR45DuQzWLLwyRCY0Xbk
bN7i2laDeDQJ8I7D60LDmZ57O3Pex1li8mvXBOtlAu2ktJVh7r52TtrNKmNMO4ZqmjYc3qyPmRV8
FvmE5UebZStaiB79mqsD1m8F2vPfXTBI3twOaRUro/qoomULJKF1Xz/UPMDQcSNsew6hEXKMuZAk
Dh+jT3dfxgITnxjq4KocV3iuMqOX7GqJX3/LXBuoYB03nXKatA5lpMvVmrREXoOKTpD4DQ9xfBn3
vuJcnyjJLl3vXhu/a/B/74b857WpImRF5EF9nwk3F+9+5UtjpR48puqFVjqypaIBfTZjj++ymSae
5aZcrEaZQG1yOKZFpic4fta1eEGHPVlrtcx2zK8gBDpXp713aPvCUgkeRmXV1K72rwszcXmF2kNk
9Dr/aPXbBEg5g/dOfv5Us9/uc+dWObgT8rZ91G8deGnFoz/8i5YmQx/8FsuzUjKUVMGKScSl4dzF
PinRR+5dvzDDf0yVPYuywfo1DKBH4M4lXec1lv7EqF3u2dd9B3t+ER3bp46z11rCMpKOiwujvLvQ
0TUFGV3aQ7V0+BCUUdsSvbDBrLbrzd2fRk14QCf+UvPASIIR4zCCw7avuL6x98kbN3RLxLks0WaT
wzWK5nM6DenCuYm2CcIo/+oHDTfe2NIpEoA2x6GOsX+pAUJAdLPo9/QON5+JBkWBO4JhkfAFmUDQ
vcyFGtFvZVHhAz1G1vSpEOcIxvxn9EHKuIKqLQKKpTel5gQd/XP9IwHxHpDQjAbbx/VTkGsH2QVy
t8duQ6C/uisRXc0KsfMCciExkzdsLpOiD9QKIFMekhuuodOQJIvtGQPyjrUCsSviLFLyqRWXtSL/
vLOgm1Q8CJ3YeIiH0zZONz621EtpAECuW/+Z+P00l4ZFu9TkzgDHPQM2/gNPzs0r7WSFP84hokCc
udIBmM6G2MjdoFmHfPkT/J8PkxJUDO4y4Fneol5V/Hde3+0yj0vGFNqH8XAYq4EVzb+h18jcAFQI
NczcLL6zGbk9gxgQ11uNULwSbRuzCEmPd37RYBNBR0cjGbGxoRkRiZGkSmuHykGdFLalg3/6HjYk
RNmR7u7BmmXPqvsBiiiuTP7j4QEeFa7RAHgV+zgMWmU5pSA7rDQUarS8pXZtBi6NcvZCPYEKzcUI
wvUIfeSuRC/w6r1O9ov+qwFbOtImjBQ6FHHvEzOw7+ZX+YzU7wBH1PsG4IsLdGbQJrbNDc8qrQ+F
ux3ftwUbhlY0OspXDJyVSmTZ6l18uXkTm/qfW2V/YIYY2Cj36eUy18+lP8zWYCLJMMW5jhd/igRA
CZG+GZY9ppqKvvYFGEB9aKvcE3sXbWsu7y9MmZKymkLCwD9peHK1Th4VovYdMzNd2KqQoeefXTw7
St7IuskbnpUe2WLadyJnFQA03SLgT6tq9P6aJm1ZaXB7X5SmyjFcTrk/m4u42bajrjDFZKpuOqjg
0pyZLHJjOOlkZisdL7fbDdrqTxSa+ZwlTUUpMlGBNwbq9DugpTuaj9FkuRsvOJJKof7iKO7+EA/F
wg3o0ad4OLbnbM0VSs4aaSKUx0sGDLw8F63AX/4OmZ7UpqIwRYWiENm3bRgGe4r1NRQ0pWQJUk/7
ZfKFp/TolPwgWrwvWuHLAyQzdNy3/S69Az3TjkQSJTwtdhJbx2vC3AHz8KfZocgY4QwRtdOVM0mo
mvdvqkA5ZaCHCpbmTuHp4iUwH5Du2d2JyJt9hY6Ec1WBrYVQJNUTKbNHmYgTfUra3VsS3muX/CH0
OUEr4cLiJIzyMr8FulmQ+Kzx/k0NwfVowa+ugIQ3dFH6G/YObwhRfVC0SOcfl8yRgoIsgnJ5TzfO
5UkPQ8EHAVU7XjEi+SdENJ7bz/TMo9UcmoarKEeGhbegOsQIwIrK5Hw1KefA+ytEUx4GagNfewAE
uMBI86WCitOw4PLj0+OI5uzDSP8XOARi5fqGqs0r4fbKeJfFa/2lNOWCuH4kUzeGmyxKikNzxOop
JOfYuxJ1BhDHJrSd3h4BxJ83bG55w1uAvEEAGNvk9hMQwV++IwrJ3LhOwKA1yydh3vDa2TMuylU2
Hpkwy1O7iyS4JDBvg+lHs2KI6YzO7d0PgShbJNSU7wiug7MiKVnbKu8PywnNEejxjw72sle9QPIE
7FOrWHkmOgauMXs0JUxjNahetXvAbpK1yKJGxjfhqE7ZgMnpdT086Q3OutCcI29NHg+9j85Yt/4i
L6K6B3h98gApbfAr/ZlQkIxhNVGPjijg4IjtFmPG86NQMThiqsq/Y5Y82FVBEoFEU6Pl3pSZxvWN
lwkmHwFcP2UgcFEYUzRerGrQfdXbSp5TVkgYkvCQLkxmMTPnTHOArTK4oC/yZvxKo5BzZUaMQ6EF
1eJt5aiBjKGYdea/xPBn5BPDTXsyq/n+/AFRRklUxXwa27zUk1Sb/E8GE8FpVB5THbj4UiXbWjiW
d25PgcYVZ5suRaGx9gti2ghP+0yn2uqw81C0Xy4evwsIolcy6WvZgRrqP6+nrMirJ7MvaG6kcJNI
c2Pw3/lR/3w0UC0LxZn252IJ6wi3CeozRuHuZHpjYQm+EDHyUb387oTEpLTMpZu2+EOpRn9FxRjY
jDYCOjK3HLO5fFAAMz33BKnk7ZbCqWrgDHXIpFStCiYk98qnr8kghNhBAVI6VCMGD8K5QdSDMRi4
85NTZ69Yv0zpQgoFWo91O+sZrX6G83QJi1InhhVwW7FY7zUmx3OmCehT35nyfl/K0rEOBF1QXOjM
FAj0kGL9tcmktWe93TTHYa1vpqN1Rxpcdh/rrdjozg1BfCusumP/ExDTHQk4RoseYdyiG9jJQB/S
2F3E5zTORvbMDoRVc+ShAru+MyEc+Xtng70cbzuIEf+jdMbilxG3FnrMsWV4OY6EXjj4oUxwNZQo
uiyckG4uZb1tL8x8bZ6qtblO4GNVjJdnfF3xFORACyQVIZC0b9bdgyZg+0S5kAHQlhgUlHIg7FAa
Kb58/Ps1cf0xlapj6FjRvBH7uTKucOhRiIrpc/jYcVEo66z7fwhqkzKc54xHUbuo0HektKfq3ayM
ICSrx5SRxyswTt76kLwzAaV0aJBIrL3CE4LNLcSn3rPM1fHQayPPGtiK4tC3qoh6FfZivRtD18OC
w53sWBnbfn6UPpirH5fp0Ixlhk4J8+W7oiZpJl7QqeAl8Y8Q+I22pNmSDO/xbgOaxJ5vh62CFdQ6
Xar6eeorWitEzZr+ufdFrqwYTb1UVGICgdGAmIbTOOAIyloF35JHm5QPuXP9/RSHgndVbLxP6l+e
o4/leUlkx5OEzZPGYJsRtGbXCh5Qpw7XGmu5g5Ct2KkP+g53F055yOJmKPN/5sfUaSK13ReXyqN6
A0VPR+04zTRnFqtKgZOV3BrL/3Afj/XccrALhYNTHnGlCOdPTQdPC2Gpbpwd/9sDefiZF+oyl/0G
gpdiQogcENO0bWaGQfgE1RphoH3Wb9b/ZJN0s9E0lddspZeIJEaqToFDjhRtTjB0Lhpck/dI00SM
KrIOQ52dhVrLU6fc6/IpyNPjzwfbZNvf+PDBSVCaRqVbSN/i5B8azdaO+arMimoAO1Sm/bD6ExAB
K04VhJrnC/KZpm+Ru53xWklE7xiSZlZFuBvRjCf+WPXCJItQ2f4uQUrk7yK8KIX7QRDhqW/sIx5n
teaDvGVUZJRoJpfI5OmPHNwYZH4dq4dZ0uVZI0txbd8sNiQNW79eaJwI/zZnexy4NYCQ2lKNPRqG
U/fAf7zYnM0AycGbIoeMb/EFTpmMVFt3+lRBhe2szZC2ec7qEdJJwjy9Svqh23+j7SCco56vyFVj
5CepeXFefNDu+fQTMD1LwTp74WdnzzGeOlOPmSflxA0nQaUJN6nBLABjpvJPiLGggKgckFAl6T4t
HUQgx0N+8Qmto+R1p5wB8bm1gTk5UMw9qRHC38Qx5PmRHTkbqM4JqTmcihWeuNyF5B+F3k1ALEIO
Ot0fr91i4rE87PioAYujb5lrQzR+mNawuDe5HYHNEU7QtWe8xlMuNkB+UmxuIIj6SuCxV1Kn5c9T
8nnvpAiQGNcjFu4jcSSKRLiR05kIB44ALK4pusAswMQW9zS1cJvlj3K/P37QDksoDEN0xY0NDuxu
+ger6kDOBiWfUy55v+Cypo1L/77J3LqdFchSQKBiTMuP0Rn5LO/wSr/HNvjXdCizv04yMn4tzH7B
j01kIDkVAITP0FAxbMvFE99rmtJ5uWLrv2xk10OBJ8/xvZVrpKG1jEuyBAjWummGs7fdDvV2a3r3
/YO+G+KUj8VBM87SlgGuvfKvRe8cOvWkgkq2YabyNal2IOTSdZCoPLql6gYTHWFmYusZhRng25Zq
UA0DTKRkpvjwh4CzRK1ZWdul5LfZZ8wPAFIUWrcRgWqaqXAKDI1AvAKOsttoOzK3kQ0cuzFyv0Ti
eZYnD0XWywrvqBYBUOxZ+4CMRXBsWIqweX/aJXn0yv2k0Ge2sLF/YTOSF0l9c6T55ZsWsEYvicXU
heWT+YUawPym0mO1Q2vyPjA3Yg4y9IoUENp3F6vhqJkT9h8jVA+/uChSR3ERS0/TlQ/NCysKVuIz
wPV7ciq9t8IsmCTGSvGp+4hgVKSvbBrsauo0P1wkgu5U2eHdtxCHSV7c442C1FbmcGfyvc5giyaI
Z3r98xpy9kOCu4QJIMkFlZDii9leRLXC46vQ0+C4cOVUAAiG/6+sLDdl5nkUECKp1kBkLY2DggRP
eVrnEK7bT0H7L/0lVSOTc2yXG/mAxS2qjglh0sJhxbn4Hav84rcal2Dft8SbQUrvduUQJQEyhpLj
TrJ8KabSiyelwZod4o+6zPlyc3ZMdNZG6jNop7INmYU5QqqpY9dDGjir9WA1Af+GFxEmquxc8JMd
FppfyCusNHim8ITzTqSVvqoNha64o8rF3w/EZxREPjFDCkzs9bHpllNt+GDBn8qp9TGBujGL+AE7
WScLajwmFU46k7hgG06roXvSdeqV8V1PNSiYuJ7hkwaNU3DpcwAvPlB7/Rifu2mxd0zZy8egbKeF
1ZILXZ7benFtHs8H89J461WpwhDb2cYLplq33LK/yZcc0oZsB5uAWwY1OAnD3qrnQiu1dJwOjyC1
H/wfVxAvm+1HVMjqfA2j7ZaqYprMiR4auskWkNh/osjpSHs+lLjqapHphRJ5ozudzuoKIP4vLTsF
MTZuPxU7+RY/lOsQscprOSTTKnhNislN6lkIXzRI8uV10SiBqq/7iSWx0PfdNPpBuAfwGUwcOm2F
Wv+5Vsh6KTvDZCICM8NW1nQyGKpQzVDNu2hHQ6XD++ZeWPyk4CfjkQz0+oFLc2HM8cC6XU39oHiO
hx/XzS5QYIa+8pWAlZLUk532g12xSUSPzyWxkDTlvqko44BK7zGT74YK7TekGZwFCCMXZeljeihu
C1AJEUYS2JC6rznCXLvMvsa7EmTWuRq2+azNsLm15cR5aQEFajcpMcZeb6LcuNiMo3yEcqidJ04q
dKeovs5OvF+voAMfXD9tCZKUqG2fzOOVM5dIzN3DtzxKCQ9As4k3bCiprsXnjnmKlUNwKLuuq5AM
hCot+d+0WeRFnH2rurg4p2VuDLSKroF3kWro1FMCtZLkhBQZBR8JfWeqVo7OSbye2FHieVZARWEy
cev/8UY61mHu+cnQaPSoaHqgPXawvZ4FKjDx9sHk152+spaBbuUYsoMBPf7eu8DBBS1LNR8kMeXe
TjJA3+sL35LKWhuRskmAo3r6UVS5FqfOsRnbXUi8HGQz+4YGArJAUcEarJjCClhBUm4/yk0P2sLc
/MhXRFA7TIc4mLmJ13VStcyDnyT5RergetPfixU8h/7iw1NeThZd0u1FJZfdrij8sCO0QGgJr3qq
ewLRVP5PFUZFUbG5peAcoeqxIkJS8Rv8fNT3a5jXzNsWED91pqxtj3yXhXIKe8qeZuE8ao792Pwh
d4+Nq42Y6Sq+1ZqqcijKog4QWHFenSlRdYCDklrZVpKzA654sl7ksBoNcTdkhF26KCxNA7MjM7Gm
hpgmWNqcQOSv1bOsjPJOMUIr2f7LBg8r9XfE+TX6730ubr2AHvwX1oIVynFenceJAw/Linoh102L
s1I67SFWB1/a6i3peUSs+8dQ7AiBacREFILbsbKG6cIUPx+/Qc4J84IeVUMU90qOzSChNS4pB59e
c6P02gf/7UsYL1n0TqeDeMyow6GV7DHVUk2JOtX5vKLgCqbZwQcEXchlF1LVVDhQqow8pQeeV7tP
U6QNFf3Ha08FpqPGlBSK+vZIyKEaJRhR5NVoztXuKZH62+YQmNN+PJnKDniMKd1TAuF6rzu/9L1U
YMKU43BQ4sw96DkHnKGmV0Qc/y9DM0maZKkvg6D9uuGz2Bro1T34PFu9TozR+wPHS2OD97yH6o1f
egUMUoOLqcHyk+abeV6uuuLGp9qxi4NzSMzmBiVVdASJBqHJXIiXCmmkK9vB3yZN3IP6TgOeJp3G
nkENziFnKwaC24PUvA0+qYVeaa1M+j3AZNkeQJTuhDN7nn6VCQ7nmt98TkfwAyHZnqjiIbHs+w7o
/OpBquqgZnDU0xETpE1jwKOqRfPww4PfWzhIBt+9v+CKZtbtwRtN/v/wHyd5zDkEC9iuk4YQXzOo
p7I8V/Pt3T1gYzaxnxLOPpkefiFeCgjgAcmzl1pVn0X3cxeFL7Bk9r6/wnw0tjPfYUFMeDqEeR0a
SUbZTYqqMhQ9HutSc2knlNQkTNkOwngJGYne87PoFkgk8N8W/haKOlyBAsNmY1//RHT60fgguCg4
GFuHlbU9PRjQuXXXMrTiacfNsV+ouDvyhLbyY2tHVwad7oWLzmL5DPwSGEgR2EKXDC4R3pdDXRp6
81STk2HYMEGGD9Wi176BN1NWxEp4pRZJd/HNWBcPhfXXcbBobrHThce7kugpMCf/RspnHr6XKm/h
tBBz2JVC/v6iemuQFetrBl+uDq57oJE9MDCTrO2mE2LT/VYV2Qfo6NyENJx8/O9tMsEJTYjxH3YZ
e7aqkKAZvovPyCNFrgH8pPMB/sVQ2MuW+KgZ4GMmn2v5gYK9EEfLc+0kDGC/Gg/bbIMrn1Xx7FPo
0NnkeM8DPtVBqVzjRjh/WNQFj1Lu9Zol5XvmYAOaR7Mkj3t6y2hhoRHR5pqt7R59dRfzXqSORYUw
oAAfCirax9+Iv0VKqtdTjWxr2potwCEM+eZp+9NT+9Z1bIXjfTkfAxIDXAfSga6QfJrwRpVgZhln
4nnSMP6ZVkGrAgs4c1EtWwzOu5EQd0YzMUyQPgOT07Td8FItR3R8rdWiPdhrT8lzjkMhR9yJUlYo
+TCZHHMznbG5lyOXBkrIdx9Sr6tf5LhwpTL86b1RLxC9aQweGv4l+oX62d+yEWtZ78eS0iZgoszE
hwWW3ysO8VSEqVxVWoIkkSiX/0NhXBT0+ppRW0wGqNt8wzulI8W2+qubCiypHhumaoY9EkYJS+qR
dlNJ7/6eRQT6LZXMt9o0gcYY7OgBUvMRDKsVMPQN3qZg5FIu/6hBDls+N5amFKDmF1tc7mo+NztN
UM3kzDXjd00hoMgQ0SeG1S3ElkDfOvr5BTjg/2rcCwY7K02JPsZuVavSkvC42//gwUt5HzbWA7Ok
9rpwzGQS7RGb5IeR2B3oipYVkFXKcoPrqSuf9i4B2ra/G0E8GsKRJ4lrpGhh0UIXTOD3Cg1OAEsN
vMG8ZfnVpQmx7FXTxEaal2Njtdboca6HuRa0I/4apIXBDS2vAFsgjK00V2ck9BMZGCxyOHrXRX0X
I6oXfh29EoBZOT9Huoewp5Cbpu4ipND4K14EVvBbGOspI0hb9q0dBZ5JBvVExVFK/miQvCpAaMMi
FgtCiIZ528mCHG69C0rn1vV6MVpm+3192LUU50giEOqhmTrOaU8WX87ItWmKgHALXUEAEnG0nRzO
804tAA8qPcZ9GReijxKsH01AuHWHt3rC/iv9je9M1M3aITABUpmB5+U6KlQh3Wy7ApcI+Q7EerFX
pkyLz1ZJAKrYHU03HmWOKGLUjAij1VCfNacSTqjuFVDwIDMHZcVBTK+SQhOOeveUcTTLwUmNkCWT
8+iurQiXI5nJKm+7oNchYegd9lecg3M7APSecB83ItuQZ9cLEAS0Nhfzgs7mXNMRqIIezYn9R95o
NATDCX5/2kR7Fwdk34mZ17h7Td/XvDPO7IY35HeM8u53Agi755UFQndoDUfNfIO9ZDAGEm33
`protect end_protected

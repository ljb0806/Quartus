-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dnmmQCADR6QpcJeREwbvZpqReaqOxwjiyewLlazS9ZAs9Vf0ugg/2mH89TAnfo+gjfxh17LA/1Vk
GnpteBpH0FxUn/N2g7GmpCeVuvG79W+6H+eKWb/xL+UHPkq5pDXgldYnS4Ce1CfRkLuW9p8N+oZB
3GBYpDepQZOobWQQU50SmA6bYrXLb8fEAc47lD8WwTB4UB3L+AtIxhm2IHCG5QuzvJqaCrZHV+oX
Rt8CcxWm7rIz8jHw5d+9N3DAFX8Kub6HMwMGsnLDqbkEnj5Sr7w/8/heuqv48A16y4j1jerZVyow
EI0ChXZ9xmzb9R79BFDp8ubHaprBaS9fYd+/UQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9920)
`protect data_block
zKdXhyGIHzrt6NKM7IxjzGgpZtjzMJY9iVVISCjbJO52qIOzjf+aoAJ7bRlFExgN90/tm9/TY5Mg
dPngX8MxvhTL4WKRKXF0lm9vU7l9+8G9rDVkhBTMjwk7gEBVOGbdAidA8Pcg9UBXXESdsppBvYgj
9rakzB9z2T7giaO1OKZRtm/JO4y+8g7qr7hzz6iKQlnNp0sh28R5GCwZy4mYmwMrk55pkSLtLN0N
0br8OSdj7HfkbVBKkYoApGuCEc/52g5UCp+T3pyILx7E0PWAvwtV+QWL1vFgSX3w/XItxBTyxTCO
JywoleGNjJzynQRaQZBKUrRW2aLw6eJHuLkQesv7jNdJp3oQoXkI9Rp73I576JH3TuX3eN1uXrcz
KpiTiOJGNWwhlx0pN6ecPvA5bLNkkdABtEohD/5fHV1IGsxiM9+ZUg3KnrAQF6mJELCIVYl3JtUx
BnIoW6ww5nBEU1n4AZnbKN57Aw0Y56fCCVdniF7OLRjjGHIFFKcfkIEHTe26dOHQt6VXPI5faRjf
9UVi/vLJA9Vt2/o0BeyrVEv+HglWSHvAtoA8O/5uY80wRfpY3XTj23CeTB6GUbMp092k1w/aSua8
VdXQ6CEhvWlh6W5jyB/iHBQi9UUwNAPQuTdkRs3KWVQnO4j0tB0Wim6bBqxazh7m1g256M/cc+Hm
K9gfjxo5luLIHTGFX4TGPuDudS5r3FXL8N1bUSK3ddt1I2m4K/G8bdwIZRkSXq3HCbEHPtu956uA
0vz3NX+1jQtnY3vXvxtPH5TLl4haenDeYtPfzOBfxX5MhmmqHfZKO/MrvNF+2y5mkJscAbXwKIqF
ugKg0YMvs3tMKTvxKkZ9327sLWxTX7w45WtnqH7QvyQVMRwduQg4WRgbFA1Mgo3TziJYoimoNPi4
rfk/k+zmjUAu6Gg2h77dv80mAoViR0DpqmXEQrHxU8YY0Jg6Q+7BbFua+3YHIEwQ8gS21ncZdjvS
+yo+v4wyjH+6zM/z03dCOqf/X9VyorMFIZz10iYoE+gs5PYc13Mv9o+++MR4gwHbMqdERfWf+sTk
yFDd9sAONMptfaJgwI7tsNEF+YoU2msI70amwMqcYpZLFBYBVc6bp4OQ8t/n2XRdDBuzjIAneSPu
fEF1f9DgoRhWHublLJR0cyN5Zu1c1m611iDX0MATPn6BT70NI35YoxmQ09FQQ+7yHa9c4R3P9O94
omWe3/YoImK8GWj/18kXS7kF4pca3mVZDAGBOKut4vSY8v8xI09ddOzGRHnw4LI0xROA+OLwGm0X
+wdU2WE3w60Hs34NcTGaCJuiDvkrDEHafw4FoMF9ZLdouhW1f6DN3/XN1P9dPbk+tg9FgW5zwZm+
p3GfT2hhojXisGRJ3T9kmLP594cQ88mc2tiAhzP16/nPs3TuypYsAokkPcbWudxNkuVnkf0WmaHF
YYyGezD0ov3R15WDESQZ4iSBbQ8mGkLK7mTJy8TEvRskkF3PFwzcMyDU3owX5qiO7yEbdFZpQvBc
zcrDdiYR1EGvqr+QoKflCcdoo/jT6tsTPFUmJ5b7NS15BTtNs8pMC/I6s1wUi6vsxes+yQC62v+q
vepthSK5HpL6TS6KISeBffNjsSONBQMQHGjW0YQnoB3VgdLadMEXgokLcRvkR3X2FUkWyv0DlpuJ
1A8syi33zdHT96L4P8QIYmA0BQ729mmuZ8qTlFMlqgPZAkI2178OZNsrbfjWXU8ANtUn3P90SAi6
QsiYhk/ioRaVEcqoX6CUabYXv8xdiSI5aN/rJWxuASGq5Uri5aCgLbjSOsHIJ4yC3oByzmNz5/0n
opI8RY2clJ88LIERgnGsdY8LSOp3rtZQtYieiQmewirnUVNHQfI49Jyda+7PMgxcVJnnqP6tbZ/V
I3V/HZoJvtX5lJLBZGHdbWXNlom1CXMHH85Uk/KHUN69/0VW12icXdVwAXVrltLHSYth5Sxhoxl6
ZsH79durwWUfggGfnU2oAgfF+RKNehe3JZxJs/vbHos6nCg2Bx9GtoFXQe1hpMtyuwsonKsGQfg4
gGaP8u/XaVtjWXV7Cwg3WBtgDHJ0alpcG+FJmO3vrApAgnTNuADxxZO41DbaZH7AXsuYUvtmL50m
ZFSIiZCsV2wTBFOXLdqhB8d/XnRVCk4TWaO5TBpX7aY9gh7AS7wWKrL1uU5t5aQ3r3DagSgOhr/Y
sX7PdDYwkadJCX2bkQrqdXnD9W/HNl8PDENWVUmTTDRkvjj2zJ3fvIHMH4ZXd1v/wcNjEJ/Q0X0D
sQy4bTKR+55pL8Camsz6DNlQDxHKbDjHrLPsegZK1vLkjRt+vAnPVYVWcImB+D+dIktNSOoq+4xE
BqsK5vEQli6hgsWLW+7F/yfYTPr+oXmllhBFfB/0HFQ/n6KHvdom0nhArZxhJ02OlhW2ObWr2CdA
Z0sT1RU/66bVejS5VXvio7EEaNItPRS3qEICe2EYUWUTV1UfG6Y6xtV2Op8i0Kdxtg3lGyE1Ycd0
OpxdUNne8QaibWF9wmgoYc1skurdBgRSpx5I7jixBUy3NC0cTnqcddpyKxxzYCM7okmuQ7cH5Q/o
0HgzNpcsulLzedqtdASNYmCtpko9DZ/kCBCO1blYPuXbwvlAxkku6mSY0h8ftt0RqoW/Dekxm1hX
J+sFs+YOCH/qOX1s7YuzaFLx6zgb8YLqdqxME94HSWed+BxvkbAZkAE21GAXcvYXg7ktrRlj50Jt
PvOaABrEREWHQuJOf+7qpa3yjBji+QZjQcBkMfxSZIeGS3BdxE29gEjftp+k1NjDasKsplM8TnJp
4tRFghRTg/zD+NDL8ZkkqL0M5OS0+XcNqFo5VZOoTKXXI1XNnBykvweqpmuJ6thTRmNEzNMmPLSb
yEPAgpdlBPmCKqY8kAOPEUa1vLqckQUM4z7XpsPIMmXnYgzvqpNf+DXujfQ1kA6mRGc1QtBM5ORd
eEXw/nNQ4lTwMgYLflTu3QJOqXbGtYzZFP9Q2cjkMEVXD811fYR2UV99qFUqzRuRy7TPHjUGrfQj
zgmoXZSb5bAKBMV9X6yuFZj2SFZGXlM0gzd6y3lYhfk0xiEjmpRtC8ZIEEworSfK0U8Tui9hUFLy
HcWp4EMpI0WAhqWW6lP/8aipVJh8T5obtXO3urEbVwrhpcr//OL1wk1zfhWdJn4s58VrHA6IyLAG
/u70iXMrp1kaObvE6/b2wNVBfUfSD8e6DtOfK36xBbcevZLniTzsMT7YphtogOsll8WbchpfWCHO
EyO35w5KFKgwLi2XNd6MsgfedLLtj656Ep55R86XQUPteVESIuQ9DrUCDkRsFFssDnMZUNBSCsTL
gscDdOMwnhq9WsSzzjNJ9vJmupcfxHhHw2cWyHRVRr1+drUq/P9n+oGLW9bRXqcp6jNFkX4CeVsf
Cl6x4Cl8RGJAAZEAEIDebNgJahzvIiZWb3bMGY9h3nJiVtrS1O1EMniYnFfgiFz9NKY6uI5H3gBS
flOVueL5P+YUbA8cmPrFrz1F4miP/dC4Aoi3xmRTOOSW7u/S63Q015l28KvHovXdienzlIiylSAV
pjKtqQ1JjauMLMb0mPj54EoYh2mdc+7NDWEdqb489LFayVEnCzAUGH8uxQlejY8B/hUcpNGL2TzT
La/WrlDncKBHVA+8sQNvPcwGk4db85yrJE8pc3QoBAutGd9boXOEpASSOz5OSMgsiTYvQ2op3/ep
rsSkOmVZ4pnynmNWbX0TOuH/sj1Vp/NlezYgzPJ4gC3vQ4QGkh0RR9DCKOwb726d8YzkEinB8bC4
322oQluGBSRjvaR2azQLDtH2lpMTke+4OU0IKifQCWizPc+9kfVfXzjq37d9vUWpm5wtO6fkMc3d
GMpbEvVsXvLzxO4cpB4fnU73gOYmp/pIb4La6Ms2teW2gyPvrPjuflWZQn0++BOxGGJZ4kvzzGAV
IzE0oUOWPY4lBdyRmLiQm/9r0zljTJfoGDc2BN+GeejBrpwWT7gjBb81GabSjBkcLAyX9lj34/qq
iGLfMbjfpCcvaCHy8Eoow3F2FxvfsLGw/cn0oiNFmt/8FEK0tkNhRWtZ8y4nreI+C6p9k2taUnac
nkYZnpYrseDbjKlz01vfT2AXjqCLYsk6GTohMbTd4oN1L7i0Xh9SnAfQZ/1yN8r+1xDFxYVhoeoK
qVPKVClU9tL3DTzW8D+GEmqKHusWX3HhM5PiAPPbk37e4aElXY3p6GRJsylfsuy9s9MYV48ISPFx
eIBUWjOLgMOBRJECsp/2bppnbjcmWZ1jTAp5uqcwO05HtEtoNrB/OvInyoEygiJVaceDMfvL7RTN
kwuspnNlbIOXgSygXZQ/on30mNXjRAJHZicf4HZckkLsfftqM+JXJPRN9Zf1tUob7yBNzGHAmb83
HShFRZRq13sI1NrrgCnh1wpQZpTRTMLinh/6PugOSQgjt8Z4kI34iAcMNOl0SPD9FpRCkOdtznp4
G6VNgTTkkAFd3SHv6e3EJv9yqRTVfIt/6QWNaw5aeEtMYxtwDiKmxXdLP8gmDp9dNWx7Q0HJM3a3
DpVYqDsm/Q/31UuXR2eLCGfDyfNkkWXsi0/sunD9Mrdz0wMOH4RnIG1qAS0wfHmJBsBTR9uuIJoq
vuFJO4oxPKWkn7c5pdEu4Yj/eUeHySnQvMQCLUbX579nlhx4RZZQNVRiNbf3PDxyaHCUWjBBdkBj
yucTKwgQ8cqMrQXK8IK2bVS1sGkpMncdTT06wrQNPHDP1jYNTNdeb08h6WVhqgE7f/pM6H4/19SL
qYsRIrQ63TiqAE+nNoZ7Y/6OCPRKXwBIusD7I2gKEw6uWflai+P+IiTaFjSXxPbZa9escEjBZqHM
ke3komudDNil3uDIL4dM18mKdxSNXxgQM8q8BomQRTwYfPgJFLYde69lVGTC5uOz+wK77BF444MY
1Wam1ZKD2eEatfcDlnEhAl+MIMo35iO4v7nJdxXlij54BhzcToDLSPOGv2Ikw/jkiBLjSVQ3Vkau
AiR0KCaXSvhHM5DTxXzp0YuRVBmN+QbZik/gplHOlLBMuoxySLWZJFkXC00Pyh8+1Wp2Y7ubLOe3
IoFTembGtHhof9moPpMTUdMbrFTIonNNhLrNzpsEnkEmUK0Y9OWJyNl0sgvjkYPNo9tD5DDbDyA0
R+qiGMHzzpUBpJLY7A4OMOq/vI9lHMBt6dg6dmrQjY3rFan3NNc239IaahVlkEJoi8iXwOYIA7hn
fWqZzERLkm/Qry+8NUH7/pXKhZ0mcLeIjGMPh3nlaFgHOdII3oXSDuOlvAD5oue9RsZv7U5sQkKY
LUK4JQB0PEanf6bmtgsJekChCxCiz+tYbbqE0gvR8lbHNoka4lJhxg85zHJucPnJB7xjzRnJddOG
5S/cDGYyEbECN2QP384ajfM5qtmxYOUHHDxGv/kdliymffl6J+0aDh/zsz7liu0dNU6s3Auuc9Ve
VfIOgJScm1ZeXsh8mAYnaB5KQgN2di13AcaUBJqVIlZF5CiDDT/D+prtxPiaC0klfUkai2WRWPR8
OZoep+TEeWjMdqHKcofOSc3YwIGAE4dqxbHslPZmoXXxV0WWXXNroGEQFcBXYJF6T0hp1JbksZMV
z0sOxKG02l5AM6BZfXY2pytUKuu6KWat1y8ABKp1mVnLPDlfX//BAGk27mQzV410EEsdCSeZPqIb
k22aZm7Fu2wYCL7Uh5lMXJmdVmr134n7CuBOlDWRYyNHqBrJQOh3RleLt4wlJsPsWS3VzlYw90RR
R5kR6Dse58v0OoLvZXX8Eqh18Wq7Kd14usar35CT/lBjSLyBpGbThQM0Y0Uz28oinsf37wI4+pTJ
zAE0qxJOLhFIoiBax1gWL0qwYg92wmUW8VjSskXTWxZjkg2exDeXaXOSsKfxi7ypeWpq9Fp49RIv
Kqrpn6QnSV4UGsqx5HHEFih0ps0T+IeHUXnzNLn2+LNV2JrQ2JOZJovnKDTa/mYbem7v60twG5OS
oA1euEt9yzM5NFwbx9dD2a6jVymNISsARq2cBNsFs6yys/PdKcPIXIE+espNgDE56qIZIIaCCxi+
zNe9z5RzF2Akpc9B/IcBd7YLqxCGK6vxn4BtPdBx2a7AHyTT7EZE3Ot03JWKYeQYAtk5bSaGcM7C
74qSYbMFdmiNrZ0t63/DAHxbyoMNweF9euoYlWQ8UswfieR2OZACsCvOw/ymSbF+lSGwTD2+qBrG
SNdGnAJr393rqes+QilneOPHUg+FtQvbKCr39SFx82cPY3M4TOtz8z7px9XoTJIP/d3A+I8elQ3q
QVW9AETNKUGyCU9Ue9scGJ5/7b1ttvrvA/cWi8A4n0opXG9TMQD15WDeI+0QoIrqX/aYYjgSVd0K
7AnmZjdN3wcZknson6MPx6SiPc2Pjq3kh+Ql4p51Pvm7sC+i8M22JpdJkVWhkXpC+ogR+CG4fijX
V2XxRwpfqIs9IwGjpREh/CFDYXFn7wZIA2SeMC3IS/QDTmUEbN7P+VJZL4rOOFkaAlz8oOS5lVK1
zNUXmYXO5aDc/9V2F7v09xx2kNyHV3uwDJXASKBWXYmajcG1xi2twVlWnYpnhQT+ElqRuDySv5jJ
UMKT1yYB+gs4bNVcBbNmHU4sYesXJToa9yXqCcX/6IOLODfA117JD97Eeom7DC3qHn8C9ffEWBMU
paObDTl4wMrXCn89XbeBtTXB18X6h1R6hApzdT9hepBvlao8eWGj/SSQABFIyl/DeFhIqy9oTOrM
cyBSANDUjX0HGsRwzq0bQeB00QwQ2nZXXKwESOk/HxyS2pTz8QKBcuezL1VIKCBykVVxdCeLsHLa
PZMaLZrTUgmpOJBFqFJymot2WSTMijMz2E3WbE0ElHhyyMRvJwQLx7cTsOm7wju2qTc9lisvTw8F
rwhlEVmDMSDhiO0sTVXs4xAidD3sfe7fpGODTHHFNZnHRkeB9or0r7OJUtFtUb8fTSOF5uIGCxxs
9vhrr7xRH+FuVGxbG2V5zC7L+PaA6CfPJCX4N29kmq1hG5gbGlku2NJ3aDKNfTi6ww2o0osVp4bF
PPZYCCwKp1VnpYsEkorlIrLlAK7xKRuqa7JUJvzIfMKhDaiG1N9Vyo5lOZlhGY093DTlsUPaIHdy
67S6szfboST8ITVjhM6Wy1wnMNccCQvo4++ZTURJKU6u7ytZo3cf2lvrIxScoW1455WiKH5Na7IE
P74O6axcuOwxb060pGj6LYPgH+nqSRwASB7JeZAn/4W5WRs3Rgm4AnEzNSFqBuZm1g0ogMlNZ6PO
j1/fYBIZ3a9DxA8FfnIzEF3CU8T8SvwLjyRKczfTU72tC50ltboBKRgDagNezFxijuGggx4T90nP
Ze6eZSOVyEoTT+n3SbC/YD5fnogTUsKoACAEQX1mKTn5a6ZGffF32eId/1DPS/cQBkOOiyKi/d/q
3NHXW8i2O/xkmP8MC3WgPCSBw0DlH6j+eP0ZncQA2eAosUPVe3Se+xEZzgERdVUefn+knSDrh83n
IMSt2ODPPS/tKxIEocMY32dbKpLRidaA5lRP9x983V8UNuRs2IcTl31vyjRLGkDSMeMWwPNG/gW4
i94xRX6/OI1HYgBhUFB37YBNEBwhVQ7EnfzQVeaWS/I6zM5t1FpPglV9YmziqNTvaqP+QzUlKSjF
VqpY8eWaoNykp/wO/ElPPyg382X9b8JZJ10PMIcp4UFi7WkPVsXhjAgcALRJnJxW3WJmJ17wZ808
RZw0rZ5n6NPplTw0iCpzCHBSF6HHhWfK5bwMYJrADEw9P4TmBC+j3GXuHQlGT3Qn69vBi8yeoumD
aqIg1CXcGS4cukvGd8EQ3qlga3MbnXBJjTw14iD5HwHtYtl4qGo2fRKKwZTUrMvfyCromTbjUaVc
W5IlzY6wHY9A3gNKpBub3SUC4/L5YG5/PURFN0Y/dY5w36ZrtLu+OSTDkhL/LeoIuxxDHphq6EUR
+uggTV7b6OUeJR9bLmSxbVu/q4tBa+5aKTA0mBDJBwS48oH35XpWFkQBAnhcIlj71zl8IK2iiImq
PbeIGKa20py3WgwACrrJJd8uIh3iKtAXPi2dY/gGy3EiPqP7moaMHVastQD5ltjhcBnGfAapVmJF
ziAPxQOxczszvHGO+i49llYQLfEn6Dv158emvZHsD6SWtz1JwTFito1++X+dnpLanWnkFxXB/uUt
8gwo0Do3Dzl/14KO44mwcWzyf/auXdSFj19Th16izv780VVKDMnav3HtWs6NZYyeFKAy2t9184ew
Hbn2GXH+/CEVlaNe2XU40zxCDlgDJPiC9pe8id4HCAtoemoQU8kUXK+H29zhYtt1Wne28031q/68
ye2aUQDo5mLMm7LPnha5uBGrDvwrVmcX0FcqwOEaqV8a8N7JOyT0GZze9geTVskGCGPitWyX1BEH
n55YN0fSvPXmRDAkWBsxKfth5Ohyk/7PmlZ69yFyRsxXKdZZPVg+e0qP7bV+vkpXAk3lRVAJRxtm
DRzM66pYKj/LSm/tKsDq7i/uGe6gP4v9dnlIVbfQE3wOJYmgDQQBH3D1DJKBGKs4fDJJjZP9FFcq
e/4Cd8Toqe5Rckh8qY5/A6f/B5hZyJTElrfrZmqS5onXxWnAzjuvf1U21anuqAkQfgqLDQQLac23
ht7sMKTX+vGsQRROjyruAgIqG/par34i4WtgPpU950CZ1riX0ftp3qyjQ81eGgZUKZHuTL6P2h0j
EpYVdAzAClOK+vlbFW3XDICAiER1Yvl96XN7UUHP5Wp5pMgzS0OljvAg8YU2jI8bt6yOXZ2ndslv
ggSN5v61PThsihmQUjVS8DS0vuMqq5XAhShdzx2/0LTpN2Hmd5tOXV76kjtZrXz99AJMjNQ0iHYI
8C6MuLvpVqTqOXrhrpomDJQacRHSqILiObSa0uhr8qDvQEO0BMCPe/JKoGRajnVzhvlS7b4YBmDu
d8o/qHfIA9+pUr8cb2nVCjNYjslRv5jRZjj4YbI5AGrjWFRfPBhXn6LKAWIJgCEPQbvTbS2OJfAW
UPgyxPALhiYBWA1wqFeqCTM039od12giF4vWOyA+nhaM4AvFzHgDHX6qRGVCoE2u7c0MATxBIK7+
eloINww0qnGmMQp44LDRt/7Mdi3yjA398sjhmJqwzG/5boDedQpPd3GeBACtEf54a5fTbspA4hsp
fMwxYXyxpZp/kpdmueit1RAi2TgfTHZU8Vmsz4WTm90LJlSiMaQUYn0yPQa7n69rW3hFcDd3HSCq
lrj5DRcdHvDgqSuwtRkFErdyJvnsiWK2icjlm3pvcL+bqMSLupOSSc6oNd3IJRnoufhAZmL6nTqQ
F9Sx1SWWf3zw8UorDx5ivTE3BWY+aI4IHDerAAUrwOcDb9doWcShNjVurETY+xafdrl/Ej1NtKEv
U8MT5zmRaMqhdg5sH0Hl8xVie4epFC6jWf3+cI9ebGiPwv7WTiYzBuPftvqee9bvhqr2PZe/DZTO
2KGJ/sxr3s1awNqTmXkY2aK18dFm+aJwhoLi7WrMeqiMon4WOma9Xlm4JPTE3FLSQXEfY5G1zn/P
IJn1SjfbqQkDt8MeAxXYam9xazWDcCqxl+cYbVObRTvSNMNfxlwwnwLQ6hl60Xx3nhKXUmfIYB3N
vYaOaYwE5BceGbKQAP40TpIJrZWXUTGVUMhJxSclldm9a4Wms8uSSI4z2lI4GmuibGqZCqkOB8T/
PXeKtie9vrNbAm5eoZe/OIH5yqvk1ZXQXI/ufOCXKVTTSTPgUyLwIcgZHWMKQtddOYnVkFfPRLYX
GQPxtbV0BXtbsVmIDdtkq5FstZAiaA36NBal/V+lkdotmhlukUJI/MzIAYUMGl4sXTY9vf5cJscQ
ZolM5fkgq7MI4/ODONAnASUWZyJrI4PkU6DEMbwfYLJRVMyvtQVQ5T8OlUD6PC8907VZgqusX5ch
D7gHhRYYb1K37MTYDlUzP/XsVLlYsimh5sNtqy3VeKN1nHRSK/wceuVV1j+06fr5Q/EU71YolanW
xCSDeYRcrgHjByR5x5W3f5qlAcUtkw1ZuP0d8R/2ZivTvETE2FmaL61/jnusslsFZDqKyo1Tolxa
7xEiHGP4LQ5DCzYAtnCt6fOT+tCl8myCbJoIB4a0PrfMHxqR+MqwE5mBWdFGNc+XkJtW0Ax+eCJE
xh6hvDtxljrkuE4ri5ZS1fr5+3fmptMJ8do62suvDKAoo0lbFtFzTCCMGF54AQpXw1TQGXcI3SBU
BTqoY0x0VDFHztxNqEpsyixL+V8jjlMSWXWhT7TGCkQd9BqyJozV1NN2L0qcI3aT8HSvUgWk9EIi
yN7D66Q0ccXPUy72BtwjJBtAvntnfJTBlq34IKyjLmU3O8C2KnCelfq95CIO3Pc94uiMPl8n0qbq
8eLURhssBTfkR22lNOXr9FCq+tlRBzPfk7R96jRKJy3l3Sxzl/lv+40pJ+qLcYgyNFNGX/uvIYek
BSlkS6kPkQfAWkxyBWzuzGTdwT+Z05LyshwFnCBAwarr0ykh+wEuiPg7FfCuRvpxKR31Jv0Y+++4
ywMc+PV0C8fFJEW221WuONhzRvYGUutfdnHwhs9LVxCAKwXo5wO6HrZs4jxsrAPMN78VL/MrlGOP
rSuzhvWCG4AdRB1D1L6t7Yak3Mj3gk8K/qA/vcSdpT3JP9KlAaVebQWUSKRpgiYbId+5s//DP3UG
B69Vpd5RRo4VgdTxIYFQlcEqt8fVswe0RgZj/buEBS7pjsRYZV7vo0SMdW5aBA88w+3Oq/HQQRhK
PfLZwGvyy8dRJKEU7t6ptjLe03YBV9SIRB0mbyjx/m+FyFMphK8e1+Q1g+ctDxwAO/iyNKPwrWbK
n5Juw7Xg/BsyrpHnsWSPt6n8d0jRzj3P/1EwWEiENj3Lpij82aY8C7NdFP8yFLZzwPShMvA8ZGaR
nHud9w780E9a2B8OyJseL3RGcJiewmq6hv0x6ie2W2MnBEwdVLzl5k8usJcgMt+8asz2cWbJEyQ0
xgrBNf3MBj2xwLyeNDrJb1apXW2wxVHxAiyFwchhXodMtExax/k8U+D71SDSLv23xeRLy2izIFga
TaFxff1TKetC5XZQ+KFk1QLVZoV7PgOB9h6H90vQ2du8kA0SYqObIFTrLTitJmy7vj4WSTecaIcz
+4e11vVtXmI/GD4Zz4Zlf4V+HAsr6p5YFuePHWT1Gw8pvbuTHXMehNS7FMuaK1rfONavErAsQCLY
BcvseJ+xr6PIWOCqZKmsFkXi5uIPdbo0p5/KAzH1BHG2bdn+dtGGOJGkRq9vSR5Gw0yFpzJLVDu3
yueQPCIKzIWKV8k4p8vOB13Kaga6VsUe1VpySHsGQemNcN+XEqr92qZzSTJDR3ayjOl5b0orTwRm
FAEYpQemdY+1sJA7xETrxqCHHjal+SWxB5/rfKCisVcTSiOCWN/Hsed7Wks2G6o5urzqRuJhN9bb
Ow/6LZk2bMXN70KMWhP1Yzk5Exb6XVvBafNEiO+23ySSHHC2eLG0yE0cJCb45zaC88TDMfKaB9dd
X052vRdePBQkWqTqKYqlKcvxO2XA05TsQj4RyV1cH3BvayK2dn47VVi8t9znC6OxMpaP1X3nOBAI
r+qEs3O2oWwSG19YwgO6Un5te5fMf4kSqWnOfpG3g4xeFzajU+gBf78n3MQq9RTpU5icmzSFvTPg
fJKK08XTUJFOx56XmbLQQVikAKZ+9fTXmtGe0PwW/+4Woq3XzH2ZtRHrQ1zyz9uSKdpBsc00HWSm
KZeTL1XnN99jjW/FJ/knIB2NEJi3smBoomavYWYa55bNGQwxNo4BQMDg0vI7Im50ToaQpka9FK5z
d3om/IulEog+fTvc4qkqEDtiNjfVP2W3L+PjSkdhPXInciTqFIdwbtlm51Ho4chzLplxFHeCIR2R
UGCkS8itQwfcAJrTJDInoohgok8FmHARH1LcacVgnv7KQu8PqtvvdJXd/rTdWEv7BuMs2Zz1UWuj
otGj0kJbHhiqsP1v2yzoRKNGcebz7vJdnYmpI5kJ37c4uPrMAS04ZyxhrDnaTsQ3zt77+gR51AfB
mE8kZEoxWLBj0FvsnL4ZOVE9LRr2KhsDdyrnOyzXm4cA1Timr4zSxEH/wX4330f2iSTzcgj2xYT5
nDQ+eUCqTNEtfSq7igrpmE/gEGsdOuS41IgrQS8pqW26t8hBHpgTY5dG36LbheBjQFC5yzSesXD9
11snRCAq3lPsP+ubS+cpaCpLf8UJbLRZ12QhgwE81yfjHtQTIW2myqxrgBgxrtCOkdrBjY1kosuw
tVZHF4H4Kkz+URieLShqiDRXyTTJh2Hf6s243C8zpo206dUKycWH1MvhojWe+QSsjkp4V9cP9w6E
ggIbwB2z7m3V2vM2QMI7aUNX4Qz8Ct8bRrEKM1y4AXViu/opkrus17sEfpB75Y6hXICEDgZXjtZ5
xXskiuVRBjq+Xz3iEF++Q1h4sWhzzenjFMBSmn55btFXRRqHXQdIjzBI4+Y3TzlbcAE6By6iYNYc
2uQiQCJ3a2GafeOYFiftsxQC8tMfcJJ6me1GELsjIbZ8ahBIbsvMH+4S5Az/k7ZINQQ9MfrrkupM
Y99YZjSp3tDodQW3/HlHf+T0aohBLOaWkCvgnxyy6hmrat3qD4F4pppBkbJw1POsMyuUqWVT6eDr
Pp8R2CKX/ZkHm3FZUTWyaIS0JANiJOxnGlgYn/7I0Ll3GuEoJEcPjlLMDRGxMJxh1n8H1KwP903u
etyWFrz7eqjTDfTNjacDjgovgjwaDYxVYMCphkkdFq3QCAqlvydo5aHMDUw2I417hbAuP7YylBiR
71WY4GAUafSo2ZOuAQNHOF7E9WsRIJ85npbf/UHFvMSWhRvlmSJegGBCbufdvaR41EMc5FKysYOb
86dae3IzCCIGn0zPJqWfW5kgdD7KvVL+3Rbh17MC5vz0vB63NoStEYWy71UhIJnNUESdwzgC3Mu8
IaFYOE7DhA3uIdsWGEQqdixA3njKXqVpC7QTkHTlEeJ9P1gAwac6zN5IKeslS5keNmXk9wJGjuzL
rWYomLdFcmb6d1bL3eqIsVfChTSEyQniM22/seeKKmwMjlnbJC5i8EadxxwhZB2HT8sd3cJnmfnl
drAVtrp+HseSw0KQwt5CpBw0Upq9l5QTnN22XshqwLsN4/FWhRm7nCmZwOep6TqOnBRJokdTh2WD
JmU=
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AxH0yEdHzZ8eBhnH1GwImp9W+zuqGXom0E7fL9Y9HJKku9jZMkoceGYFqC4iUVL7nhXkMBmMVDsC
q//ue/ABk3EKv2EBv0UYrtSrOIn75DlcyyZHo0h6fkDbmeBvWIMhPsc7qBL78Ty0SnLUpt51pJhD
3JFpjjTP+WHs/kodmjHL2INkH56ASw0DDYRrMqizY/dPlW7BFYbk27+iRuYPFrq0o0XXzTAhYrUI
NW6agz0a+WkIOPd/HHn79Q+agLupLD30hJ4MYowdtcUrfxjqijOCRr56OjUWmxQDpc632FqY259t
F6O7EW4mbupE9r7AVjWMp3mvdkL3Bbq42jB6mw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
THFgTeiqbNBZ70sdmwjmhhIGdtTK5HGiz/w4XEp9PwQDSQW6uE7s6UP2kDuHFqiAkvDUffGCqnGe
PPBEDVAzzt3KXnqeIBcyX2wCxRQg72S+sarDG1sVBY/jE8gUG/d6M6tDFmuwREI/DrTohpap2dTN
zigcs1Gby4nJROMI7L7Dl/FxJ9ZA2f1LPVh0dEAsW0FwZx2rddRpl3ELqEwfXhBvSQQbUP+b3sEz
zXuFg1N3uUSWNI1L/vgSFICnft7kv0EEgC1ClxRM+dPB68FHRqGR/mYY1BsEC0Mp6IjMrC8suQP4
8gLbgcnb0DHCrOTzQHjiLgEJeJ+XMlsdloNqHn7vAonl8i1gNaR4O+xMhLC1o7Sa9SU79EVZtzN+
ug1cb0GuuI1PCkWGh8Luin7QGuxP9Nd2wsdgN1RVUrTHskrGJI1I42K48ZgB9o4FEDM4/XwJfbdc
jXIKqbg3bWK5E13xcawOoCAKOTUBVntGmnraCNMBd36Qxnn2Zu4GM8Tdhjz9Kub744BPtSJXm4C2
q9bpCpr9Qee/ZPkVTfx9ExTKhW9LWvUYHJ/eh/MFnVgdZB0UmmmUiHNmMKYMVTzwxUDwz4byTKM5
PPFpBWSlR9/cTmrTWQ69TpVC12JpasE8cH9+jQBtB/i6DarcWe1VTofuP2/kmsDg8aRkZ1jMaPgr
f/hzHSVvs+tH8Teb+VfpxiBb39RDZfsNSpXyzdaO2AuXDRGTXhw9c7cHgycyj6ulL3ixL5NkPJ2F
5N2rHaCIx0jrP+QjecGBAhHV2s9oHx31WyOPxjgONXY6/ccT5AwJJVaBQPVAenBLKliud132V+2G
J2YYI+h5b+ev6BNJw24R8VTEPQPbGXYePBJ+wG/YdJ1Nw1xGZxOpzM8oPdoYgvaywOU9D9Q67gal
P3auhY2pd83ylovo+8wcvUHuisuXBO0/qVUGqVrLrt2WtZ/3bUO0GZY9M+Ja7ru1VZL4Xncwehfl
rQjtFku300+oetwtyoAZne9DXhz58FPmK+yeP5yjU8n9bBszC6XQ9pQ68+ukN5tNqZhr/DzKEpIp
gcDINs64Bml2xsakpwqnc8sWjnME9mlysHmVL55rZ8NaDp7gJhCgzXIkJOALBc+xQKhZqYnLkhsa
h2CuxwiZX4mw4yV6IiPaBWDx5l1SmI0egsPcvgE8pddYDL31WqDA69auosXHNOduad85Gw1nDDzK
TqoJyQNBqAkcJIoO4hqlfDRm2Hd76FPVLHCv375K0MGtkCR9M0lK/BlfYjVOUP1PDRJTXjBSGnpe
dqsvDe73WI5robA9TNtvJcLo2jBq9AERNky8fhUU6Nisw3+p6zydhlPJjd1gVGU+252d5JomjMCi
X97x4j/Sc8Exl8nu84iTFHXhV6hrIAw0Z8NoSHMSrg0tov6Ko+SECKCCtLH/9ROxHTmhxcai0Jy8
sd+2IFPYz5BEDTCHbzuPbcfgmGtHOE625f64KaOV75yd1Wj3EbYn6PBwAHdDvcXsoaxbUGW43tiy
SLViX7ldZX+LA5d3+f89SJyKuY6gAKTY/QXAdNC0U5vRtFb03DmV5uEln3gWAZOV4mYQcRGmfhhk
Kv/0YiHJae+ummYFIDNiRVTamzzGkUl2HSINmYfhqaciH+u8Bbt+w5u4iJwvSJZF04NfiHt5snt7
q8scIoiRM85Ho75yyU2JHldHD2Ictg2ZJZs38dcj4f37aOQ2aUm1ogO/xCbutd3fZSthmZfDQGc7
2C27wyRYBkl3rSeJdIcwer4jzCU30ce2wSAHQADMxPm4e6OV0Vq2Pf9oehlym2VOK+p4WORvY+Rl
VD5QyrMTNDZ5Xwvxlg/nZ6dyMt4Ds2PHRDJ0nh4TncflfBgBfustP0yzgx75x3ar+vNIgmVMMU1e
RalA1syzP7GeElLYxYaEzflz44oVrmqnB5XKYIp4uGrp9t731goEBwvy0CCvLJsMeW6tVkHCfcLN
UKoUMTJmGjP+IPRt4mavAVSac2OStTS5JLDjWEU35TRFRGJ/Iv2W6hflYJKtYvtvg1QnhbqLAVDs
MYKEKPe8FrNMse2bJQxeCPJiSQ1dwZowcf395JYOOF9qvK8/PvwNbngfCJV0fmJByw6Ze0M3pJ+2
VNFf9Zu2YdMs5DW+dJxwr0R+IG4ridu54FQrRdTzSF2BSs+fqPLmiHE5jUt2+aACn8PyFw1+gfTk
MjtgVEcP0RDyKevXiCNnxO4mJcH3ZiLoA37AGGO7DqaTRKdyWitrEVHtrkPtZ7vtTCh9ceFwU23L
PBm35i0VCt/GQ/ERmBXr3oj0gQTMdT42UEqG5Fa9sYe5e7NvBxI9LQ1X8cyU0rQ02O/IXhd3XDvU
scjhGomPjfFEQYaUBDhrLg8JTe1sYlWuEkXZb0Z7N3qPNp48aigsot9GOurNORzAZQVC/JhTUulX
e4f/o3Euzl6eT/G/+vaB4GduD851EPALpYEiT2zwBX7pe8gD9OFagIaOcxta11FUMrjk4TI++XBf
ZKpnwhX27+/BY0q2eVcAHbB5/zRNf+1ypjmUl1k4SYcCdZxmLHJU3HqjkFWL9+r5OYCqICpC9rfs
gZ83hUobAtKcX4yszd4jG+rttZq/svHkw471S6bWnePWjNvyZqNhmhFwiBWTePnxn0VfpBgRDAGp
WAgCTdEN2KDNtbuCer1uo8nHxTHGoD5XdrAmjyunCHgPjUiwhpCVTC6Wx9pZ3ByrVd20SxmHgRoV
9QqqghcIvLXNMGzcRyCqvOwGLNOKhNcTDkrhBuZoo7X78egqIUGLZjJIflS7B7bjxx7VWHgfCadW
+M3PQB1XKY3vqejWiKVLXAga8QkcwKdnSldzQBqKOtRdXUKZ62S42iFM9Fm+s7R1KqRPac7X4+H6
cUV4G7ume2ZmNWJDwiveTIsB0ubMGMOdpQlZOHJ9zyT7GUEpDHC0nEUM+iYXIqtPGyxorkN/3r/9
DPyfxpJqGpsFI+nO+Hds3z3YydW+BQGH0dEeF43RWrN59SnwPgGYJIS8tRA9CnSlZdcTWT3yjui4
9hFJvombxj8mZlg+l9kjdWImTZ+P76pU2UJWqJ23dW6ohYe2cik2audXp9SafZpv0pAW6C5SMdHa
5hEMuOmMewI/rXDXRrrZ4J1/tswe3TVXUi1ZZyllouqzm3t9K2W73lE02wVqz3hyruM2h+hxoH1Z
wvY/FJJ+QDGjMJQeAoJjNT3uyBB9KixsPXLxhHZJLuCR6nWRu4AwcESgScuA6zjEz/Rv05Tz3pKv
Z5fXF9aeipsTInmi0capOQk9OCyIoDcMQqv2nCRbkw/fBb9sESJ3pJPy9ILKxMIpmtrjNOlkxeIW
PLWNCQqsGwwKZGyFJGof0BETgwIlHS2Y2CxNhjF+ScKkgKOT+BS8uf3n+e0/n9xlwqnW2SKDtbAH
BxDpdT90zh0GgCyI58+l/pqr3GzyAHxK3IWqSgK5iz4946sZcZERXWmPfBDkRj0vlrSQRY+1vPm/
heGSCMumagkxC/SM+GzGjfUp/7YyEqkEjE+NM/ROHUtgyDREumVce0m9QQ6DgxgIrUM7/yk01sQ8
/SGfH2oFjQKH0pdmjAfesloaEY8p0SlIrLc1/zoDcEzsH4znTaqnCbc1SKuKzPFzke7W6juM7PDz
WP6IS/4rysoqRbo95qOEz1VI7L4+R2KrPddmnjV+lgRi8gPD12JLhfn+/CTuk3Hq18GrSifXRV1i
D4yN+HSc9naerQG2pf971C1Fo9ko7KtjDvZ75HaF5Hi1TvTLre4RJ+ZUHK+fd3XKluk9oUC9lDQR
+bLe1t62HDcLaCny5FeL1B9wIKVAW5QbO6F4QntrwMGh9tfC6q3kQrcPTel/xUGw5QX6x7dAWzuI
0nyIYQiHIBKjErfyShHs9lrX2FkdSGF7zGUUxJMtJV9SCTn/sA6uNi8b1uReFhHAgu/J4rFkXNt9
3eUmGS5HaCQkfTDOqouSYrm1cdSoyQaZKWeuqxUMJekm8FB8XOL2fAIDzBPNwhT2ouQw+eHxfn5A
tU+3hzAG2+bqFkyFPTna5hftOBDgR246Vex8Huz9q89rDKOPn28J59hhoK9Jkzx+cVegapJNCqmP
9kq6k4pcnjCOe4EH6hdK/9qeqfiKRoDoB4rjZc7gwMUVNBCNUWL13hmP+kQpHpgO/slVTnaZrqgK
gBX2z9Aaj3W9wU7mkz8JGSjJKEdlVygZLx7Om4EfWW+MsbK3hfoU3raz+6+BMGHS4WxKtONkaaYJ
yTI5dkpQ5jl5bfZ9vafBe84RiXRzsuw2V/MDlCocIRmlKWwYk1G6xclJu8q27M3b6V4fMMD5f6tn
NjNrptRPFLFBYwJPgFHRX3QBT4T5euQZ4pb3U8NdQDRHjIaOxF8GRUV4FUg+zDNCFmEsJ/znyXfG
1d2XpOcFUmd0yiRWx5zeQBPPOq/j7Sy4eKnsrL0dRHrAv9vluBJr+I+wLBPt4s17PFX4owuMkOFz
HAqbbM2Y9cxeV9EmrQZdR9gKrmPr8p0iNd+kA7L7wjvjR5rNbLmia88AZCw4hqfLjbyJb3Tr2LgH
7ZIlncvJnxln1VDRxZlGOuJhMFFIcBVXHz8GBxSsp+wF5XWIZo7TfjI00kayZM6rABOjsq/8TGrh
PBTxD7aRZbxPNtI1NsJmvD/Wu7O6ehGdrzBvDq1tVt1ZBpJJVopH1VFfngtCUywngnbjBbMvjyAO
hYV7usZB0qSiRvRUfaZJc26sA04uw2eStT8i+CZBlUAB6jLFfj7paE9oS6hS/w2N76iA1JEVYPvQ
97Bka55iirU1DKchy3Df+/bugfNlfRbXzlJvCGOhXDNJsTCTfpGQmc1zLEL7sFgzSFbqGYOw9BeP
yXXUkYXWn1sF8dCFxY8JrkU8moP3jlpBg22wQ2X3R0uKGLEORaGu5JeUYP6Gerb3Zca2UKADbnmr
h/DfZr4wgeDpjjrgRa3wXD3iRFPtqyCELyMBe1w9uY5XfFiIJRRd+H6gI9tzPdkN3bHXGtAZGfuZ
4uod5E8Sj6BrelZeff55Q9ZSs1HJV79d0MU0JaZfMRXjeXdsw8ouUiNoUcEa9wtQiXn144pN5Y9I
5TenTTOKNLO/czY0QTcNQ3nB+/SlsQ8oYMmRv0lA3Ie18SXgzQF5MGSzthSpTxfiB0RxyYYRIA22
lGroK81/U8+t7mA1rBD6fE0VfFQbimgzCd54NJzewUOXavx1hUVfGD03EiRCUUaOmSIwaXQ7nTKf
E1JbV4nn7hKxxNQ7+eusQwoWgopoSiQtEzxyT4JaBmoDpEp+QPXgJuisq65KY8sRpXrp0enddkQr
L/u7b8FH1pIaXDKpEt/Qj2cLzDMx2wWvXuoMvG6M0SOzKjNtGoLEWFewQPGIgJDqgji2nQHFLk1t
Z6NdslymBuceYm9vosGX1UkilJB6e1dafrwDc0YIXRfwmZFMnIHv4tKLe+/d4N07yXEHhG4EMvuJ
Vz2nWFhCWsSvSZBlUY9uNmi4KOpKSbJqFxrN+rNRlVdioISaIaj06fq/3q0UPa/d7Dy7+P1R44SL
+hu9H6UfGdybRDzOshTdB3MXeWVxNUdNHvsgC6Vqp0sRSc0QPgsu5xozxrYdJJPDj9AzcX5/DZ3e
YwJKeOyOQRR6XRDU2Oeu01potxePnx4xFjmNAOTbJcA/jxtrSPr2UmAhCoaXeWMwtM4+qNVOZUo3
lH0bFbHsXpH/R2T9JveHaTOSxzFv5kCFRpnlKp4H8m/HkqJ4JYRrWHPJkJn2tGaLn9pCNUcVLtVQ
vL1c0VSSohM7skS4a4S676WuADfo5BT7QrkPWc5I13MrLWDvEZSiLRyZQs9+pxO2drOfASher1W5
Z0i1MhzKMH1ezQQ+NP4LWnZB0OFPbUUjV0VaynG1VQmUBRWgZv8r7a7QxddlJWGkIcFJWING1lmS
oZTnCUn1SZzGQMjwf6vKxPpX1nZFgstmPGE/E2V8GGFesKfP6bJ/MutKbm9jiMYYwA/nJXXnBZzw
twsfsKuW+dZQi99FmDZOwg//Rx0KS/kq8ZcQQHjEfoAKVa2CwBCpCxU1jPljP5YhBiqHVzGoGKaZ
FH0H3Xrn2JuVZKY9yjd265lokkKIS3cO0/SXlrlt3emRlF50aSBwq5gf7htPW5WPzwTTaIHZdr3N
RE4OmHQE1kNmAhqD8NFBgLlq22K1/RycUt/zhU1L1DKRYZXbShLzWTogXvLDZpc6bQDCXPtubJ0l
pyObBvLbFlw+wA+0PQqEQBMXbGJeUIjK5nGyErIig0kizrdhXGwGIGLsFRuvN0S0fpiGcUxnUXT1
26MX1XAfHDy/eeVlq5KydugKEBknSpUpsyD6MQAvNmixvcff8yAMJm29e4ZZE/ngFBygpsJJAyEX
knphEGzXt3vSJE/H+GH+ceGwACZgIq9ahrmdrWYXo9Zji8BPsFFoMFgeg5Z+QPPWJ+qeYzrKuglV
vKlfVSbpiYjnKsuXlQPci8jzDLxq23ZCpPzk7/WDC9xLYDfbpV4UPjFZabGsT+nv6NEFI1BJ2+aI
kEYJMvrFiZknFFozJIK+xxDNS7BgSaNlZTYmV3VYqwMc5VJKdeUIaUmX31QcgGHFxlUCs1vabUlK
14EGIBKVjzIhRkigwJRBsRmYzJth8VZHQK5so8rt5skBI4ns4/zLhcYTN/ohKBsbCk+C1bbccGvZ
Ul/w7LRpBoEH+XUc3NxWJl/Jx/KAhs5Q8IeHaE3QZGThNT28JPf+Mp2QRoAWRvohVxfvMdrlhfxw
pYety0beNRouMzsdRVPNb9I8o3CIKkYhEkPDm2Jzvt6GpUiKqCmYdHyHJrLQTwodBYMeinL1z0qK
ivTcdE38WfX4Qpw2q6dltAzgufretddDBCJBr8AP5F90dq6ZWDdLGftLSCo3JQf4EQ040+uina1o
38zyymFon/0YC1+UseSfbR24BHvhGhwjuk5vcucYqRXbpO3JvqsSPE4GuQ5IeTf8l75ZTdcZIgPw
fpnlwdlpLX2xvikSbn/rB1AVO53gI6eP9X/WPeH0Km4ziNpN
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
plwyn1+3E6TMc3YE9fTjVwAsbqGzB3QpQ/gQGsyLxILOk8Hqh29zZ+fvumRkMDPRdXxd5stva8LI
smX2i5wLj3VCeXxCquQ0PBuc0GscJrYfknDia/zdpS2OgBqcPnvzxbBKksRshvCFrB41cMkat445
B/NVMP1C/cQz5Y4W6sWhuTt29Ftrl5RLU5c4pZrvVtpDy5F+pBROKrkTDl229VS6z9BUKA/Wci3+
ZQ+6T/WljtJkVV504CqLBUgi0XSPgXpbpIND0xDRMU78tLzAqT0MIHGcPz7rDAu4bjjTIqu7SGbw
RXCU2skLHM4omqrmV5+r2x7P0y0WSuEu7S2c+A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14656)
`protect data_block
78tNUzC5sU6nsev9bBLrBhNLbkjxzBOpMqQchvEIcYQgVMQosfARIFTvCl3fOFKAmOuoRdGmPV1M
tFqC4Rck7mc1uT0urxzivPQmIhkE0LIqJU7KUQ8mtgvBFoCHCw3im20zCFMYaomd4jwC/tS+Xdwi
tZNQxRM/ja7NuWrE2cxH8NZfhwKWbp/I6gjpM3nSDldqGszJJayhHY0fY+/QanIjFY3TORBQ3nR7
rTCqKMsaDpC3D+zweoACSKS4lgpYQ2mQmwxUTIugopbTGzJRuLwuf6yTdOt0gIkxGBTKsDrcO50w
JXZalmXY29OvZcNcxJHQEXyDCcLGyIBRYK/kGw2nsbpmRJnuU8F6IBIm7QklgE+VRv4LJZvlPZsz
OiT4oIwsA6MujRLCS8PLkSgXx5xlGEuJFbMIThCKJQksxElOjKqSPuLEl1aUmEWUDriaYRFaZY41
ElLgSnArXryHONqZEDp76TC9ca/VBM0K08Cjphr9RbERm7CSCP7yrdN6OretQm2PmEz+UY/0zAXy
qfk5wboalQPRdbi5nPJY26EcH+YeFCUcTOI+2zEUD93HowAEaQFnw34PLztGyBfBWJ4TDVCtkhfD
TmKfTQ8Ac04YxdjJkP03CA2mKpB7jHRjXWTh72QCHSlavSpShGgad64mnW69Zyh3oGvyTLHvZaVe
y+cL8G78IBV2UEuHToDO/BpA4OfPitieMDiWm/J/7vI25qFUAdGUAMRWTeRUNm+7bQZR0qsGXbuF
efPfCPLmxy6MDMelFGcZMyezDtsFhIj8gpTpubmBNoEjx57huTDHtuZbnZHF5j2gk77wnh8CRNbv
/Jz8HAAPpYi+fm+Ph2ukTxLWBSVjaWQXagkfvuDaHuOk4zAKgrwk5HkghXRkRcaMNBYHT63JPx4B
B8oCtw6ppf7fpSYeuqXpg9DvkXJcCv/q2HFWWRl+nTOIa2m+n2v/MIsZdw+v0f8P1aoGuVFIovVe
dDVcTSfvSoMcYIpEt0GqYx0ePkBRc0UVn134d+Q8qOx+rFdfgNTnkfBLgvG0HFQzkzQ18voD6F33
g0/nbtFJ0mV+k98+nZMp3TvYOdfzSrL4QycAB2nE2XoXgT+uSypnwI+VbLyMkNsTd0otYHw382ph
7AkuUkd/JwXzNzACT60W30o9llCgkADv4v5nmqlJzsaoiBjyUuH/pCdUE8J77b845u7BK1nKamt+
AMFbcMxjlaJJI5jUderRvwVoLOVXvDd5x4mXiDeQo6JWaBcHgmVohkFPe1VSSDEY9dOccWZghvON
diG/8cz9moedDnwZaxSR2LcHvNT/9yPUHa5bYXQr9EGRaQYW5Ted72gcURoqoTrbC7FJxynaOMrD
POAHB5OteGInBf/ZI7OGVbd/0urGofbgRNMxb5y50COjpZsTtEim+0APOOV67o1wYUNjTJp7LSTJ
RJ0bluy/wjNRO565nWs1MwZ7F0sOsbLKE4oMVBIsL+OpZlijAMNIjyG1Z3NdWMcPL/PfhznlRhPu
cS2niLa9RbNx1Y6AzdWpm4OwlQDWIe7u967Dkh1FIOfFCyvYTJU9TAhZU8bI5sMGlOHadE0zItZd
B+/Bc2jKgLyhVhfHRDhMyXhW5jyy3wgf2Z0rPnKhKM0sOut4XFHp5hu7KQpC3GgnudOqsiAYM4yE
lPv88OW1wCWkl/XoFnJ5gZRwPkavjJVjK3fO/4R4b90t0wRjwnvLZkCUdBa7pXw0P8EL4rEKvJsO
3jpkeXAHcAZCgtyoqpl32VgiiYZ+azKHNGbIifmJIXTHWVIvrUswkdZTkBBet52rYfwvuqTwZTRo
Qb9w7NQ+IOCOVElghtUzBmgJZH2KOibhtoU1OB/1lN4wEGNeHHk7zjl5NDWO5WBAvzu/6UqejE3h
kIuJ3zqd4N8S+IgHNpTnue/V8CE0xphZSlrYDbo7PPNJX6dipCEQ7ywvcstVqSxpBrFrwz0uv/V6
JBmcMdIF14H5Dd063E0hlDqOSnnLEk5JJqI741CG4yRiUcOtoylSlmXMBVky8/G6652IL/jGDdQR
r579pz4/2EF05dFMjypLRqD/LPCRCvJtaYynM+oxmngfOO+4kLEvx/2/cxghLhFX6BjYTCU+QY+F
gQAnJ8EqsJZZAyvrm0LTAz4vWkov6M+UJ9AxgH6+xXeZjAtEb0f+uDhtSxa5jkJ7ByBEiiimz7BX
QBkrw9TByLO/wgeDapOty68w3eU1mU41PCfDcCSt4qOGzFUOiDtSdD5FDLF82yL+n47rmtzr+HOf
v5s0qs9C/kBkxIIRXcg9cDiUIHu9+Mew9F3y6KpnDpbEfaP5ZRLrPfQaAfoxYBRn6n4lLBlmYfIV
KTrdKRjyH9g+ktO5g0PvxhvJ+iRUnQOUozaR8ClmhUWKOA3hyLhptyIvwrzq58aUy6SFN3xHgvXl
tU37QrrcMJrAhLgMCF/SRFjo4m3D/2tYe1CELIQsX/3Nqy0yQWceH9XmFsXc8VD80d5sF2SFMMg9
ot7yBRadHIZhlDRe8lkNt16B+ttxN2fr7jkf255zt25kekLSWWpBc71b1NDUX/ke6ypRCE3uWj87
CUtXBcdP2p91Zb66o1d+KGCdv44nNoBTWR5HYF87rX8+cC+hn9ISvI4US1HUm1+p+Bcc5M957wdS
bLGbg8Q1vkokoUuXgbMpv/pueYXbk3mmOaebu+pobyui8G6a4S+1HO8yX+JJ3B7hLuvuKJDJ319J
oz5J8Rk6cs9oDrT94s93zI3oIMab12E76Bn9jIGvlJEz/RuwzKx5Ed2ZtzjmF+6Al+vmvhn/ggDF
nlt5oCCNoA5DrjvAafRKXmvX1xXL/2lbfTNyu2Sd3ikYvmQBcR1ue7HC3ptvJ1Ibl3VnwBizeIa9
sM9E+RABUCEfy4pW9xj36XSv4j3yag6XWL3Eht7I+usgjnokfg6L6Sw7ml9/2MJpTHhckOPH2y9v
PNSQgaw799RWCqaNd4DiLDfFDES8AX2ZWCCrOhS+OlSeTtu4AupQXbH8J8Vz2fNuTEo/mVVRosH+
StW6lrrip+VJBL0LGlo/6X0PV30JaSu5Ua3Kognrv5ZCO/NBEilm+J1EjkYiH0yqgDHV+m8EbWpH
XsVfjXh2qUL4n/hRNT3Ezke8JWVUBJKCZDfXzM2h1tVsyEDp9F60eFe6/RZzMgQWfWRDE9sFYYWI
7u17C6W7ts7IxE5Atlm9iMlTKcuvCZFX17RATLJS24nsRdf5hqsBwO7+nn9fxIMCwViYX4p3fhE1
FkIrObLMA5Q0mtybX+uYq19Hqhbn5E8cWhxL0WB5K6WnjsnTpO4aYs0AWBP7wEvzhZsdmSqfVJCm
EhUxiXM6/qGK6slVfH3phu9FU9F8OxMvrg9uZk5VFsZVXdbFUSeFAgNE7QdX6Bz33SwhhovuECc8
sPsSHdlo/znKljXRF7bXKyhqgUvnQSzHkxsJEKgZ5nDvpkYMMIZzEJMFwDXlG+N4buKePsY6WOwr
5wxfusRb7prvqy1EcesfmsvKc5RZHaVt3xRS0ALadrMtdzQv0TWkduJpfQsqlpLyQHnhmrkGsShS
qz8FUbq+xNmrCG/eCh4TV2FtaECI26RW8bF2e8QqrLSsiVyRCJHAU7j5vO0ypqf57fG2NoHd417g
Q0/ux3QjdO9Fn4RDreRPe0dhjGjzh0yVQ+1pxdLjCkFubsiMpQ4wd7OX4XReqzucY8xQD+AT4Ah4
JUooh2rvPjLrHd6z+jCS642atvN1Xk32w5JsP3uQdMuOuJ0w97puGEfp44yPe/2i5gGjJYZzXzIV
7N1h5nlMOBn2/YJBC8KlaQFEjtKr71vaGX83GU6c3bHd56janU96Y2N5AjrRLUZ3/zwBzA7osm7l
4tKdISj59fMjQahk32b7/pN1/x+VEakf7CS3trkARitJVIkWzfUgHhk9f2rtEzCnZEICyHGvnqvh
pLuMcutD8NSabQONz8uh6+dfDrmWhXUHyBfgbVAoQGcgTiAYFtmhRI4o87AqWh9l1Io/pEIum1cI
o1SSBOOhqbXqqFS1gY+1PZH0WMZRe1b1ENuqBgFENZwn/ZyWWAesQLw36ujCX4HlBw2JW7yDFC88
XZaEWJ02eMNg5GXh5vaCv2bjtkKRSWsyVh9XpEkCXDJ9LvF6Wvi3piFElJW45T8eokN77OG1LC2C
vZ1x0sOgPdSP1yolMwdq2PQDxvUNQkRizA0Uvvweyqq1fu5W78e4ApqNLvuBJB3SAIegSkefmi6x
n3BNRnYBXxxowo1yI1+bbzw/yussLugTlKlmo7AA4mfTntprL0fnrz9V9SY2aaAhwB9a1VEA/Jj0
hiWxTVCZ3MnN/AJQDJSKrTF+mURcu94NnEdtytT2oYPoxVjvs5OwxKFoI9YUHPBwYvy1zgcY/Bdk
KGM9Ogxpf3uRj/DyFsEwLW21mn+P9J3Ddz7Quw0YhebS9+Q0ZZiuXPwPq67hr3tvML/KA9i7QuCe
2H+uAV+QWNWBsZbnDTwpNfWVSmH+NXLHYHCMECayQS00rGs4yhbS01sUJmwnL4I2jhD389WpLjLv
THO8+s/rStI+iM2hsZjGLtqezKILZyyjGINXdMO/cUgPAJ2ys4+HXJsV01c7/ivsoKB+UE0sjilp
nCPk11OncQIBj0hesxsLCpoJoVg14Lp13tNRt1jnuCXWpORETv7WFRVsFktI6fzcCOvItkwzQg6b
eYsAox7Vr6DpL8YxK+wbamh2VOFrRqWr1LYE4KPeYXFlZtTGLbAvbWQZ5p/OajIwDULH3lZBa9gV
5E/1pMmmNQZm5O8M7ZZvK+mm8x6ozUid1cur33bfL23LNacSc96TUj85P2kRJGdnKXj5KTUpHQvn
nKwbp+w6/gJ8ObejOCNZ2ZAiseD0ausNPzDmOu7PTi4PWi652DOucT49PIVFZL8Hsj9W1wTyHu0Y
iDrhyta2BRNK5n2EVm/WZc59QC9jJopDtoAObzygUVyxQKDJxCcBuRQARZoft0FskK/5BJGdBjOs
m2rLqHCwxttWVlUFuej27KPqgq8E5OHpLn5WXC8xLynYBCnLDzHJrJz8RVK/tnKXf4LHrCHM5+v/
7iPqH0mkk+f+JkaCfD3xTxdPUbxyM3qTj5gnqxfYzWrRQUUgPReYUbQs3scW9Gfz7srt+3d97CxR
L/hmuasix5R3ehU+C2A2RgeUj3J/fPxmQ0CwUHoZS58gGn/ymjjEEf4e96/ik0odoDCDitXdL1BS
8ha7n96d8nzT3W/r3dt7GTyVPUn7LBtNYCQ5OchZULHXFfJFxSVFcyZG2PUv4Mwo5nf1DJA4k8Gs
SnZdc8BYEJOfKmo3cZ846OYjiRJ1y4GiN2VKPUOO4FIjc270s79sqScc02jMTBDyuha6SCT4YKkN
rsMBA3gto+3pJGpoBwWJNNcLK73I60HigiCllzeDHLrmzX3NO/sF2UVQkANESl64P0o2cu9TjtWe
itfBmlgmCcbRAgsdhRAM6g6wSwLuhBNqBFs/UibkbRu5/zwNVyjqxiG64AwDmkxlo+lRlpcnAQMz
cYa48GsGnEis28/yXhGMDQTUxQHLSOGEFqEGwwHcOYauyZJ6di9MZ1B4G8fFwLhljFCuPH+5GtHg
kdd9zvH+AZufJ/qifmhkh0uzNGmuW2oUZzU4c2VGHyy5JlWqsCGiI9PjZbwuU33J8jzILvNY/CDw
dOuLxuQ6pSbjXxge+cjmFhql7AlhDjwON8VZcnXaILInJEvGIFoj/Fbe2YfEaRTGJS+BINNn1XEc
c7ggWepnuKw+63eU84cb7QanrtB62U0XFtY0b7O5CyihBqY8hv9XAecujJZfOjB9iYFi5rabHi4E
a42jUtQkmPyDwMtavRKOPWzM+uADA/BZ4qplFlTEAUKgO3lCssV/QlJ9LznkxySqUVzkwqxH2pFO
GD9koyHALE0F0C3221pviEmOnit5hrGinu5/dA1wueHfYhmfKiT9sOH/6SYKb2N6kvtTsi3ifnAI
8LwK7zkFMHxTCf831YP3ryNcD5yRMxiUb2pzIBNGdNJdvgJmE+JWqZlQpfhcA0Te2WiVFtaLEWAY
Wee04TNybAY2RLMxULaO1yseUMqwmv9/OysM9UURAtjMunnUcBTbDQAK72Oa5kxFgRrUSNKKchVr
q3YM/ahcX9Gt8bwout8Oa0reOBQ4pK81DbaZOoUEjbw0wspl+m7D8HfgeBRiMxM3/hERBtg237EH
VE8sOVN5dqmNViQjvrGh0LJyYy9fwbDmy38SRY2N9hk2nyUkeNyR5dvTtw5nvDW9JesDd50DozxT
GjJ8P0JNq71L+s/zsHGwfkKKLceYTTF8gnSby0qJK2qehm581U94ElT0RVPUVsmOj2+mNdNIzT5B
RLnKCnx66YjiaXbWQNbQXsYkCv8p5fUU+jPvR9YRnKcp1Lwkt2EDEQnFsXXKQYfA76QaHZ506ArF
sWMTpyGgNtGMlXNAdtK9dWEHW0v4p/tDlIMz9lecAnSRJAJK0tM4ykeGGWixZ2ynb1s4BwEPDsN4
+RNYT09htYUiwCmp0vdMxFZAXykJuN7iAXa/UYMd4Ll78W0RDh70eL7zYl+Dqbc/of0tsOJ9CuCc
XhSYc4EHEVDdfgnSGzjCAJiSG3/ruXbV3We6HlOJ2CyVWOK5Mz66n2x0a+gbvEm2agMBpTftSIOp
YYiBPS0gsZvj0TLBCp2myYGCeqRHvRVda3lCNxtVv9HxXOHiS7W9Ow1qFFJ81bIEj3ilw6Req/ik
ko3zNeYKJdGZ4ktgvctiGmrFNXWGDzzxa6Kja6i0PaDdIlxmHDMf//zz8D8xmF81ZGqZ6sV+o32o
bQSylQlSNkUKUJGiN0rpqRZt8RnTFHxFn1eR+36vlI92GfHWswAlRgxzXGPcGi/hbkGWDktNAHke
MkqbVMkNY8pCjePSUDmjDxHsiX9OG799JPb554zuYMSaKRi7AZV5qFiwz4yS2UmiFx6dJxhnlvzi
S4lJdB9L7D4sqBeHfCBDKoPvtWG+rGb2Ka0eOadw4O+9TCyB4IRAQYsAcPzGP07PyVCnbqjjPM4I
GscK3ebad95J+zFBJWug3wVMAlsImKo0dR484/whWpzEcT2pJTSUaRjIeiwTcLnO1sn6oBuA1Fk/
gBkLmi6KXOedQ7AoY6qcfhkx/pvybDSa6vdjgbEO/+3LSVA5VXZ2C3b094Naa6DGzcgYk9wB/wSc
RR+0Dxwt+f9jPnydg+ZPVjKQZMf2dZSMQzO8wLQh9cOT1gQpYToEZsESNfYa5FKMFhn5/RA7pqAC
yXm0ASMXpCMFpTEuuqsmnNNoPHzGvrykxK8q2h2jO0iND08JyvuRZ/s8S005FPJgD+9ltVr/MQfY
fXgTjzKlKgib5sj4YcazxScbPReCujbh8wCeqKU1TlQBAJMx1Ii23GyFgCP1toBoiC5fJJrxmji9
jcowVOpuVU+Tr27IhS2JovrpFnHVxnNsGdSlzjGmRM4ODYB18MX+aJxHeCesLfHc3XK369erq/Gq
KDPb9qTPYV/MYpMC6AXpGXAo+sOosPGNAmK1n+2f2Z0MXFp65YWmUNd5BEpQPomvgE5ZzQlu7otv
Gr9vkK43seMfmUOpLzS5SHtqzYd7Bva2bKXA8E6/1MVN65FmOensZV6GD7/Eg96kGacJGw6izcdM
YymnIqiVbdqTXuxxYPlCBPOrbO4TKlwFf5lKmHgJ/N1jLA9Vw4+NGQIpSWZ0g3n4sxlP2vTFAEVB
XEp94YJbdEn2g6qbGiW/iSiAuBzkT+D9f4P5XCzC8SZBLg7Y3GjqXI33eNO6jgcnyFJL0OVcxkHv
xoDFkat8JW3QXQxx7WoHAaEjjPXcSX9XtPoeDMELr0782KL0pyl+a/fw9L0XBkXv9ZdH/7gO9ZJ9
dtAZkxJRfyJQM8P68J3SlMu4EGdA8m9UIZVQTg6Q98IBRpfahdd+2PREBFC2uZ5kIr7afvS2ZerB
saCZEsVhXAMWb0BKsV+M7qpr9ljuT+irDHUeeJOdvLVpZQVk6tLY4Fi9VV9El/81Opu2MiSM2gc+
DPmKnOPmwg6QqEyPjHjSEsostXZAL3oVC69d02Ii6ghgmwff8+VJKauCHlhwhmxIGjSQJJgCxglt
Oc64B6eKTd3ANtKp35qVuDrSsT3Cs3UUUz7kO9e8V1s3THuVypbkHm0EU1YdtjVbTKcNnOMKuXrs
2auDM/2jgP8ATH5IO9V8gD4JEQKStT1GPty6TRRci7yGlUt4gB3JN7VmgrbbIplAq6JCiJ1kjhdB
tYzh1Ln/66mj2LFQ9LuApdzJ4YVLv9+qlcHbcZm8ujd0v/KbO5S4UfXabtCXQTN4zQnHd1f8Ajih
EC6NBFL6jSmE55+AZ2C25IgbtxR2IkrXmNFO+K2CoGRendDdRCnhUt8whluajEXO0du/nAia26+a
zHLmkJSX88UrvJwbVb68wrFhoi4Sf9NYf3HkissX+3I/ohZbKyIdb2MXshfaX47MsGxJfh/BBMDq
MIRVGUgSbH/9IW7qoQbhLcjarbF/ulrec8kh7wrWdvOeVB1j4ecZ1i6i4gc3/Z99e91mxCJtGlLw
rGfm47xRCBOUD1Wrx9Y1JZHTMxn17r3bHtmyaWFt8PaHVEWjhJmBVM1bv9aUuWC49wb7i2VAe3o6
7+nDRZiQTRBoYHKzO7INFeBOJzGUno6WGa0mhYFSwe9cnuTDvKzGjPLsSnCJO0OgaPOM+U1zZIAq
0xmwNya6mJw801quA3X5zUnRw8mHSih5DIsds3+QHl+va1MY8EGWgEWIpD4OXRJuYOj5kVuztCmP
CuX6HRbbZWcqgdTD0RbFhroSwJiW+tsaLjOT1YanLrPUqIIkocGGrvXwQhydHmvQQH73/AIj3TnY
Oy8qZhrBIhmrS/BFHo67UsGiDYLXW7EQMilkPP79SkNPdKOyB/+RZArc1Q7Y78cNe+VOR2ANbeEi
gMEjK5ZpGAoisUPNmh4HzcPDx0Qekz7hHOoJkI9KVLZtzNDASCRVEpX6KPZyRxPvTXCQ5lch8m7D
XcT/RvivmOK9WlAAoMWLKajbSadlA+tN9yiBnQIUFxnBpqwZ63W/10gucLSI7IhCuSPbsvUrBZAv
oBlKQJpIWxGzPlWp/G8qtWZejW8hG5HmnqXTrjr/xhNtQDZfX6v1A5hz0mY2PAWAuv4qRxnSZL90
xva1PAQLkuZNalgvP8Hn1APvbbradmFfDqDlUNdw8N7Vii5tp04MPIsa6uqtIQAlVgnMlZkacVnl
FfuXR1wV/mEei3MRSHKqiSqQPad0IEQG3f39r/vqM+POmMAW4E+FGXRtvrbTv//3IxVwY0gY6Nww
BmzuBt55GlZCOvgBlibT8Ray0GvtCvX973KkPU2i5o1tdnnqOYMVDzzN7kf2IGqV7Am7J60B9/VN
gzqJPuS50chAKPROEIU4r+RUZys+iPlEG7rZsmLpzn7KvEc0KtQ0fgRBtcHXZK5j7NvqHCiOxrxU
sp4ObKFNdEbQm5VL752fpgCl2TOjKMImBzZvL3aTMUjM1v2aFh98XwvMz3wxeZDcfnc60cGh7d3M
BZ7wmBat462DPwVyyRjgFitWDG7BuIbAQPOl/ztqson9ZsU/c9takq+FgBTUVhzVfllFnWP9IG9W
vQumB6CoymLLz1yVw23Izu5+zOf4SMod/eoIDMQgmeZdtWyYGugD88RMB52IiepV7jLbJSW9rzky
GEbdF77XafemQXWhAYbPq+rNelt+sUm7kdK9UMmPgSeljXplbSfL3zzKQjz6jcWyJyLMwE+pmdGq
Z90UV5ayOK78zCwYCsUcLr3eYU6EdaO1mPNsbdOhFgwxjTlqdiKlculcoq2rLkwKl79RDwsZQyPc
bA4lfr3S4KguHiRAEHbMH+W6Y4zdAbiUfmg4nqmqOfpRqks7Zzm1o7ivu9KBa5JXgHVIm0msQ4dP
WbU2Vfgb0TrZYZ0sbGkXWYkwnes4KW5i/meSwsQPJKuJkw8M5tAysS1zCY/5HDnjLY+0LLcpHtY+
Nbe7was0X0pHAzLrJWW9SCxhW69qHjrmQbBsBpnvAfWnViy/6zcIwIE0xnF/O3g/Spdjy0pAqOHk
gogDJV8ordXDXQQygTUU5qUJwAsZ+Ih9NPSLFLOMsEAlK1DoQoAMfAFmB5qkYxp4OIylLOvDKO2o
tErnMyMoAR+lnqIwgl+mOv0Eq+mQ62J5JTK5v5+tnilBF4DIOt+V4HxKfjlewHMqQMadgMZgSgDB
3ikInX5nCB7izjJ9M1XLeA3ikHefx8a/Yk/BGFi9g/RKN/1X3i5cEPfQqkKbBQx8hC8S4MdQl1o1
iDKenG7yj5PVa2uaR9f8fLXYVaP9o6ScW/g2GFkj8GcUIZ5AtNOMnq06AhdVhcjy7xJB30xuFDr9
uFbve6nu9coGB2ZOumS9mgAA19MQESirBr4LyPFrtQzwW3J4p6KUz5sbxayCrWK+wFGjvIldrFbv
a0Z0GNCk1VVL2Y+RuUGRyQaBb5pGVvPXxx04FlUXMf88h9kLZX+cggGN6XiRpImHohKpQ3LukCD1
huj3meNrvVp4MwWyEe5x8NX8lrnnqMVhHQ7+Dl6ttD4axnv401P6kzYnxBPoo2MIyx75R0pDiD+Z
0jC3EusV2LcS2dC9yroidV0siehLp+mYwYzHn5Pyitmh0piOzbf/YqyO3PvXUPJQZerIeSs3SMq4
/y3bYg1Zyjnn1bnJnrpsmFVdXsy0Brvwff2GN5m6oOtjp8HRm9mfu3xu+uujdgfHmBeLybmMl4Du
l4q1yEB2G0P7vlCFOJ4H3U4tNa0eHWpkaUWi+5nH/jzs2w8hX50AQkFPQQRYSJBXWu0ATpHBzyFt
uLs3jLUeZVnxKUKaoHSExpMEWFz7WOwl6c9S6Jxf77LoWQe9I2ss1w18wGRMfkmAwa4kcFXedEIO
SXwP7M2IEIDtgErMzOQW20hDk+AFrjUAbPUwQLzL3bJq+deMHsdAY9FGkotO3Vpm4mLsbEs7WUlX
JEaUCzrmRgXu7d98fjk52Fp2izrab/xfb/53FWYzHq/fjql9xHsQG2LeBjb6QAILfaIEURpYATdW
Yax9eDU4UAmmWnw8aajBtPt5rLoMPhmNlH90eEz72pQzmuAeXuo5aAtR048Bks/52RHlFQnxBltD
J2HbIV2kMBdH5xcF+PmgdXe8CfLj/DtrPXCydfq2joMVtQ6h1vi6wAW+/sAf1PpgMrJUWjWTLwxe
BG+JA6aNR5HVOM02K0sA/DEDmiWguKDDh4hryS0i7EQebaPmRa4t4mhGfbFgR5geXbM6j3mx9fz6
XaTAymJM54w6iLI8vyLwxO1UC3RSfB3HNrsvlGfrnQoVz9lcb0TNG5oIPZZ1/T8lUwdWJnzGg9U1
QVJL9gigW4P1tdtEXMQfhUR+PrB3m9zB+jrjIZPDuzD1dk+BTvbMdJzjlaoVTiqBkwbVtKMW+z0W
01SDC+BhXBsTC9cQ+8sthePO7yR3Tui2PfyQUb9cOBdt2XjJaBLq76YMZ9q7PUuFtjyf3CzXCDKF
4ArTh13IVLjf1eZ6JMLKo8Cx42AXc6WHlR+lvDVv/zK0PBolGqqdoWXDSKkUXEcJ7mCZSulbVwIK
vK0IT3aNng/1/mEb0uw24+D194hOXYYf3b4ibiPL24FF1GqELY9UGrFKoYiekGL4F29qI02s8iCJ
ukDLmz6Eje4Uvz57ox1QniG6zo1RGuVn4xsl4RW5li/wALfo4pmQAN6H66QxZQrGbh6hqjvJCSDV
T/tWe9h0nhFJOyYf10kqh9ss8AYACzNZ701cuZOpSuZEKCR0NtmMoy642YwMtJ6QtcJz8MV3qndq
H6Az+8wy1eoWJOGyWZnxThx/MIU996vxEtpnEsvQmWOEZaFfnfhL/TgA4swgf8HlNPyVlYEviacA
dXwdr7q28RYY935EFACJV1DiQ5l5qFoR7qHjX1/iqI7UZPQkgKguS3UYM1px3whVzrDhrp6xpL9H
2Kenkr8NALZoQGBeBx5lcWQ++ZGthoqXZvWPsvFFFjcnRO89llhH3K4rg82BynoMI2ZKqwwdjjal
j5HshUrX3CdgV74JYUnn+VsU/3b44bFcu+O2pxmszfPwymITWB0nkJYRacpEH7k7+zmIkd3vhkc0
0gGltwgR4nfYm6RY8aloNQC7nSsJLSYvlU0IQ5s9HGZRe3bEYzn2SbZRuVP5IkXb7TktOlfiberI
ACwiVHNgwW4EJE3Sq1ZC2vrtCFl2XclXQ8JVVmpxbsbgNfRhIFl0M+xHpUIUY9XgivJF4IaOCfXI
6zNRN2Tg1nbvGEpJwdm0dz6Oy9xiw7IzMZ55P1kVR+6zKSDJKnNidovcZ8e+tbFIGgDfTC8UGA4J
nLLno8m3y4I0KLnNOG5mtzC6ivcfONrJuti8rhOf0bg4RHPCbMTVMzhLmYjslZ7FsQzmaOxuiBqN
1tcWlsbgzXgO1JYTYhTcWx1Xv+63FzmoI6rVFV0mTsE3UJCxWeK4cN4gfCdvbEjNjc+h84+TXLj9
VJxdZiZxB2L7LqEoofRJIVguZtJoyqTyJciBi6yUezrfYFEtDjPiR41lhpms8sVOfBh2yDiVZAmf
DnHeC4e1fxa0KXqVi6ExO1s87rDTC9Rz6l86mKmIJAEq6FycxKliXqOgHEVvvuI9VhLkxGViKZfx
yzzw1toEtRI9V4jr8A3wY14EgdGDIG4sp/yMA4gRPSkrPBO7eo6+OevPen4D2byHJKuA48WC20uy
bHky/shTvJhciuHbcdplAjHrOcyH1fq4jdALozYtXQXm8HK+e3yEtBam4modqJ6S9sKvDYyckHQJ
Y0RllqwtV2jpiJKL0lw4ZEO9OjycLMy0ULAxEP/eLj5aH0rOX1wgobcWDEQQ/dvTfPkvYWCPCUEg
WwxAW9vkcqChP3QvpGgfuS3nCwgV5vX31LhNs69lJpslJw34QE7phUPhFDpMkJRcGrDTxFEf7G1I
+EFSYXorjEXqLRomzaEx5XQHFiryfT/LH6b3gcH2wabnhxGoH6EjmRrFvL9u40ODzNLnQixNdABP
7wY/oEvpY/Bzp9OulwuC+ZqfL8e1MUVruhBtVl25pqqCGhlEkegmk7zQ09wwGzu2BrDdSI7+XCbe
XiMs0zzN41FxSiuhUOo/OMPkvIZ89YBPHfqfqLhqQuEqmXm9cGgpu7b1gcfEaSpwesQaKNIiyJbk
+GmSsEeKCRqTPbhcXCoMtPjDtA9+fEo2EzvfFBXm+Zfe+1df9gyUIXNNW5TiLsCViiqRVOHtHByM
zbQc3voECq1uDvVpeC5PgtIVdxPVZEHpF5bkw4vtAIujt+g5o9lDRwZUaPIUAbpdkIzYHeZcnVgF
IbcnKySeffSZ4vrajk88DefYQ2zSjpQN3H6EombThtWZPmO8I4/mdH8Fdcc0zTuDcbsZ770Drshf
kqOOMXKR8GSxqLlBo6hNNGGtr1JC8hYkHOfBdOseb3/bAraPYS5iOOgP0bprEz8WUg/98QsZO9EK
Gdp75XivD+67CsYYkr3XpCK+5p3G5h+cVKHZjBGjGvlfciGHjTcJ3EUhbqTxSega24v+Awsksxkv
4DgN8rorS5weBsckHqzigJhvYDIzAoF3mJvvMbnIDl/Gdlk6IM6q3ObwvEfP75fOJ9/xgErLQIDp
8I3c6r6bgIi0MCljRIS/A8bZgdyyM4rfktiKYzfLrsd6wYI6JURbYz5EaDd7ALtxSZ7vPQ2FAy4T
T+JE7h331zZ80RJsYqDMwGnIDrQUbuwSXC7T6voZlNsJPAzoSUE4LGhKUXRX8YiJMWcVK/sVOZKW
iyh3OGx9eZBLH35TwISHBDH59QUpasoUEMiv2Z30TTBTAwi7Oud3/4JalyahoVWvXQcp1OGVFcB2
p/KD00vfg/WJsefcalZT9CMMhC1ZL2XUXEWFC/T5sgkA84BzAM2ZTv/6UWBZqFiE5Tzi6D8AeksP
5U8eNSZPhepV5O89KLSVx5sPi9x/EIa2s67Z5xAOVkaTszP882xH4iaOV/Jn8LWYBzKNkl36eA7U
63Y0GnZ2i6CxTXn2LCXQSvH7g0v+ro9pX2h5LDm5Ykiu91LVdTzvvGgGGYiU8oPKdZISEnmVQPxy
u8QaLnb0g9e5dCWc3DVrOei1m1rzAP+dntIWLG+EPT3bKfb2dNurkGXbKQoGidnO5hb9EeMrYIZu
geuzYjrTeD3q0rj9UlK8/x5chlTyWDUmi3i5xU3fFZU5IeJFo+6x+OHQJjyt3rSMnFmpiJmwsGqY
kJjoVaKsBz0XJYolZCOMDbPC4tpzIziyaoxpHgNIleNQ9RPf0ZvbqltzmOh+krR9kRocgZNvBYkR
RMKq5xoP09bOoBtu1uX4B0i79RTuMEG/gLqglHNtW0Q2zXYCrDiiEOkLDYPnCkKiykpKJVIRrLo3
dpIaRPeAOkXguRxIbzcQfwDnEAJpI+0rsZGWyMaRkk7QdwubbbiG69HQOWMqC5hg8q4O19mP+34l
v/8Ot2rLh6MzAJZzIEa0lr6g1DNTSEif22eRF/RIup5vDDbJ4dGVh/f5flrQ3oamNuRrFEmAeO6G
+jUU6cU134EBmzfDQ471jnnNHfDUPM+7mAxpaWBwLojytyAf7HwXVn7qdMytLAQAqjIroCpgk18F
M2hfeJ7vc5ol2LLohi+EYFRh/ldfuK7ATfHIS+9Wv+nGukxbckzc/BytTtdWPEXGz0vPKPEHjZyi
K0ora7W+EZscauQ0N7L3rsjYFQf/HfyM2IXyfLLNYnFBTlVAa3Keo4gx7uRKhqtmCP7cKkmqxBp7
PyBfHV4MlnqLjHPYJqKcsw4MEOc7GAhGHgDJKc4Um3AK4FbrutJGt/uXNHV+g819rF4BfNjq81Y4
Arrb6/sskHkJrL9bT4YqCW83VIdgYbyEmtW1t8u50cvjIxgD4SKJoN4UhVs/yc8y3LnnvzNCoHd0
jvXKPcpAwGAgX8wLH2+wkLoml9WNCm0cDV/R2mHJm6HjsnA0UfGyep92ve6ZZinn9gbUSWKYWDV/
ltcaeO0ga3ypu/HdRG3ds2+1DGTRD/XZm1lJRWn6nERs3SMhiNQeZWakDpsKz8En5lU2iHbTeD6u
bvr0a9VnuzoR+LwVgvQv3WAejKY34sy1M75jUZo5jQuMWPucY9BQvuzvY9dg+NkidR+dxZccO3dj
oF+8VdPmzF/hsdF+Kb8DtMaawyUD5P3bIJklRSjVKaCykhUwSUL3E1W0Barfj1Ogqeg4nMSV3pJZ
RjGa72KgIw66dwDpq+0PHB+DQ1X5c8xyvtj8s/HNgTQU+QsaLJYCk2Zo62ch+TaBE5GaU307p1e5
kCCsmZehABQj2RfiAeRgoxuxxsqSMhObkddawXdmaup1YYMyYwrH2pDbafHo0dybbTBpA83Cvu5D
cy8t74reC0mddgbLqDoUDf1XSwoFlcSJRL11q7GLFGck/DpAa55c7CrjYpArnRdFtuy711UYjDNz
+2PPmNzy8fs9zt3fEtCRqj41AeXTjSQM0fBu8xhyt5EI+zGZtfH+FOSzf38S+zkcX97b44ttHSjf
96HvYMw4zme2skdptYPl6SGvZUevzPHMN/bLri5AD0YX/bTn4NERR9fiO4F77oX+WWpzcrJTLgoU
Svr/8BJyRQKwvLqPb809HLlOmSOSSgJRt3ij7fMMr1cGOgzQa64oo8rVswTQ7xGTP927DdiyzvCe
iBk7ensTUTm1twy/PyQP1OF/yzej7gMHimWKqci5ROv79XQYxAbDEwos1bYDxG+A0KZKJcYU2qAo
ocfgo9P/sA/9HYQ+udPC84roFxLIXSVkIZk9pG0rWKD8DPx4nmIDt0B8vhL0xvvDIM5QFts2O5AO
fY6JhUy6tcB1O4VQ1qHlbmEp6fkaCLJFHC4FRYzBCs9GCTZXiM1lGIUQomK3L5+/HhWykAbAm2OG
jDjaXWW1qI/4C9jHMIQTj0dp8eP42bAUv2z71LUXjFwKUyORRc+C58ZXbR5jKPAN/4UCHVXhi8hp
1jvyXXpmOSljNf5n3rFDJSvYyGXIgXO3HvUWljYN3EviKs9zraChAHv5riQ/hhykIMlaY3P1pGcE
9e3SOPMyALiOXJqx2M8yIu2OeN/9MciorPEwkh5Zwz5morkxe3gos6/F7n5N5I914A1u+c90ILw5
BuzljWXDx1KlKq6stJHXCJJOKsH+h4H4xHuJhKUPFIdX+NhJzj4pi553/OL9TKGjKRCTjR3hbcQQ
Sy+oZBLplcCxGfXSGfuZKijyK8PzBm6L6ALKXu0zp3EcxnMUaStkkSWLkHcDCIrxrm0zJacB8cbO
q3710dLo7L8lv8fp/57Yu9Rt04VS6hvrpt1JlTg99BSUaesCc9uLQ6oo4DJnadWYDqRd/yLJ+V1u
i4MKhqTxgXlcu9Cz9McchO1CYFDbCjXxY6tXjrg/U7z/bXDrinSjVFWXUTCrKkvfpkk2dFbhYPH8
LJYrtv4f6rWvTClxlvqc44JZe2sGesWtjdWheanGXRq5/zxxRImgFqlZJ4FRQNTuHVJHnmwImmKK
i0lOPx8Fb1Oz05DpUzrlkMDY4rp7xYCaAmmsNv7DdUkzb7ahrsi5BJ5vhjhjFp6D3N4S3ouF+Nfa
uC/uSD4OTVZEvpxt2PxIUXyg76HsUnhXpZIL+h4cAuZWweAzq5C+qDKEHvG5LQi/QC2bNi9Ul5Sd
vT8S4du9UKKtnkm9+oCzAURqv3SvJT3YFl7l/3t0241xk95XRtC/bjR3O3agL26k8jlsDCl4jvDF
ESOZwIepQ1oKKBitwsO8s55uGolmjqF9W3Y8GzPbmfaHTAykeNAe8yiAIZBE8iBW4TRS3vqb31uQ
lzxiuTob5m3dac7fHu4DkGba7Owoh6YK4V36PJhEnDazvlowVGQjH7oN/F9eD6jMjGl0m128UFZt
tF4f/nGeDzjssvLyb0m3XsqBIjkzBA2yFIF5uuIwFaUBK8Hxb7zbeYMcrc/4/sZO8gAv/ptoSHZh
Q3PWwnBaY7P+CaIERfxXHZ2ZMitcHJ9otp8JEdRxwMgpg4KVktjSa+4JwrITx7Rknj1cQnA/+SZE
VC8ptuI8tPXeJ4pRoTF6fOTCd6TE8VAujEmH8rLbx9IrkqAdu1MmwFMUjeifxR6h2tssdsJ+2Yyo
eoZHHZ9pJz0hUXo1Cg7TrqF8HWUW5Lo5iS5qcd1ewL7iemmzdg1XqXd1LCvZL3ilqXbVUH7k+2oB
quSFzR8XA6WpNnsjGWPkmCBaH4s9mcp2fkBE6jirvey6d4ejsD6XvZT0NrVXO9nmlyDOaJaFbez3
QRiPq1Rq+t4pBBd7KCJQ8FFFqjwQHPWsU/LacypWvzCFUandSXXw7+k2ggS/mhlGCnmRR9QIRlSo
yWCcIDs7vm0I8iEJKAeGTSFRIqtbJ0xSZaWnapPW7T6KgyPqPxNQdoP82moY1ACF8F1B8Izaeuqs
BRpFGSN0HTDQjFfE2pxvwqSCkfu74SAFzR4XVPMl3xixDipUrHVFH9UWpsL21Ua1QFMbPvgghuj0
KKOzl3zfqjaY91+ZhHpslEnRP9rfOo8/hjgjSXx9Wdjc9Z9Ahx2G3PwyNj7GH3gsmMxhS724U6hZ
By1XpzveczQxVdmaWEdgBv9L9yo2lzJGjTRIJ771f48SB4yQ2kmIKAOeKKopZ2gnlGShMZYsizjb
1kjHE/WcizA4v4K3e1GvUtRu/DSLWBM4SI/c2VrY0t/DkZP7bhBTNnYFvyvxI/p0Ddkjck+u9f86
tn9pFes3V7QdyT5grpd4rz829bLC8R9+UV5oJUTf6RjMZ6Mu9ddCDLmiPSQlObGX5hMWvlE78WOh
C2qHKzpUFhqWOwY6ycPWm8IR3WXGMGBKD8yl/FqdqeA1jxIqpU7ktqoZOoDMXCfL09LQ5TxLxM4E
ywrTWX343pPkBOFlMSM/UV0qVQExkmDbCRAQ97cxq5x+b51aiRtWruYb/ekb4uQGGKZOJslVfrAq
xnkK820tYIXDqYwDJF7GZrGSGePwZ93LiPvhSee6B4i5MzqA4+dVCczzf4KgJ/khKx8TUuyDjasD
YiKrOXsYnOxpiGMuNpl8Bup8BBUf/WNB9ASRNYwZpWFvKvCXungCsTlbnfNxJwfBUDY+hkf+Gz2N
FKAi9e+1hKm8dwHKmMXHg1Z4ohUERLygeUwz1C/SwbtiA2Tvn4wo59wfQ8ZxwK9mA+iJFWVkGsHm
dyX4cYW4jDhizVxgte9gXp1oH49kZNTV+o0SNHKLOmDKdngWFBrcKLj/pPDrK7CVZpDLBQx0GJaj
QqS4WBxMK3zlUQF2LwXUTjfsKBO2w+oBroXMTYZE+48/G3OQZjizUBD55Dpztlsv0JYkeJ/fcEHy
R+0VoMPvuDBUWayACg8u35a0470kLRsVcumq+YVbvvrawjUkxCyomZm/YvyKm8Mq6Rq6k4Mym8gq
DmHOs/bIaDc6DNcRMBfgxoa4CTrY0rRphNGlan6NkLyIAB8LohndnBtX0YxcZTtU/yiy5dP6CiB+
Vnwx7LxBXN8FN95cuOmEaoGM7SN43E3JFk1/yHcdKKYsBrYhfM2FtRlNUUvA+4ySmxoil7G6v/OK
pVHuF/IvbSAzozMcTDXl1co7LU2zDhv8LU+1OqT4yVrGFdMfsckU6UJC6KSN3cRduIYVYTgj/JJc
C0VRrXGrgdbSKuUDitohYMHT/WcxUJAUnO9DYdp7KD+R58Q55GONvWhIWdqcF4R9eiOLMZsNFsNt
7zs7PHhO4dM/rOW5oRrEG0mylk6K58tvclLX1sKCMTRMRkUGCRJthOuSEBMa9wBkg2DLZH+Y1Be6
RozxnHHEa5fZuCsilWjY8VixTM4SE+sURQIzOWUPsFsHkBfN9Ujp5b946ohS0NByEZ39v5LjeALr
oMvlVrFrbLw3WKDrulOPoXapHL98BCvhIxQwFoHka+4TJ/UK5CO8B32cFj77v98z/Ujs2kq3+2R0
M1lLo8EOgkpioc90v495VH/2ZepE4HqP2eRnl43fxF2EJA0evvDPffg0EBbc2alHxYWm4WHyM2JO
D0Qke+MmykLWC305Ha4Fd4TTwmgZgJPFMtqYIHS4Or2Zzh+H3HxBQQLjfNUgwOIQWCKy49GhhmhS
MHvjuvUbFYVpFKLYLCuaU6GU3WA2psA+WHH2pzo5dgUbrlDyfSELWLy2XsUXBqu0O168DfxhYB6M
x11BjsmM6V/8Pa4/DWhRzu9mXyJKcljo4bAARJSAmdAeKQzifIbTSK9VOTk+JK+mk8XzWLdpqRZ5
OkShRWqnJYxEU9gaCSNOij6sLgxJ+SNGQsKejT4JKmclKh+qkdVhykawYXAj59nSvmtd+HVgRYBT
ecyTPoxJI1SjShqMSn35sM/sHukrDVxFHjEKWD7tX7L1dgAYbrBh5mOfvStL5Ts3Fz+B6TiGct8z
gCI/Z+konsO+iM4kzygpOeWcVwVW2j00JvU6IwsKCNUH6IqtJW6RJ9XUrQ/QEpznK6OvRNsTcQt/
LKzbbxGoog==
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fEWPiMjD5sBfHjGljL528SUIyV+qGZGbhtojn/vtwhnO/5hCiLb7TqibNFtYIja6HwRYGMrhnkFx
mAllHoFdUO+zoL661i2K+kg2wf9exBDnn7Ef89nmkvTUSyl8dAp5hUd9oYtNf5cUOuing23AgJxV
pZfT60ont3aVO74BA3RS4pnowO4NPNXo4LRY0dj5g4nhAXiZaMbRxqRD5DII4xpEKH0R0V4iIrIY
v6GamsBftO3KurtZL+kJHQmRLhCydjyv1PjrhFREOFEprGDZ3/AeVn4a/+1pGGHtmGfFdOgyPpjN
u8Kz/192LpZ6p2QKF0uv5nlhi03ugNKLnYhXfw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
S3U+dc/npk2aHXzrPgdjXKYDNFOy5qgej70GGnoRmVi7KmZyLCffkYraJ+Vsj09QZeP2/an/tMjA
hjBYWMm0PJwkqWfuWANks1hDuURfUQcAryZSgxhlFhJXMf4wToeZ0i9VfwZ7NDCdF5qbdrVAQeJV
JbcR5xDiy3KW9aKJkD49XW6q1KmhfohddCv/DRA2tqv9MxLyAw6+3jwssjHMCxFH3T+dhvEkNBcp
oLs9isY15yv8WUYnNzTKX9qIqJjU8xnUheZ5h/uic0v6MdugVKSan+zUSz9F6HjAP096lc10D9+8
WOUDIm1VWqiJWT5eKrGAm/5H1rtNgoNj0yZ/9JA/iQY+K1SReHkRlrqahoB/q+9Vd/EctdTxa7Jr
TM+t+lZvmBtb2qcDqvg2PH9JsMWDa+gBetY37qsYqzvhi42SAZAU0IOIe+lyaOQ3CUjxLJWCO71y
HQVfcsHPKHDWSQ8hDWU25jCOp00DJONDkldqxoYYL/bzoncQlQlgoxnRlxTa4mLHHhkTUmiBxWv5
ENRhPAEOLLnLLXOqoUjJpnRQe4ild4x632n5QfE9fZ7RemjNXezEwzVpP+LULNKpk5p0CPstTD7k
0cHEb+p1LQdyEKNxpNoEiXf6adFF4m43kCpUBVcRJGLBTA025kqnszD65YDa59yDqrjOWfdXgNba
Y7ZM9tr3roxrD6VCWMCWLtJK4k8r+zZrWV18vS1L8aentm9EW+IelDK+6+oP6pPbbK3zVi4fdmcd
sF/q22DsIt71xS1BODKg1rttQEOAK8v8o3P8PmWbKuFRgAGYLoHWnsGsZdricFsIdtfrhsO9LUIJ
IauR0kr9CJYwqCfa/UOf9DOAzrMNA0tJEfVtnyRQHmfKYK8SDgFEa0EidCW7R8ippBIEnpnkzMFB
Z5ubUr5dnT55k809H+l8LkNhZzJDlXz40L6goXgAuRxa5GC6NVkUIre4VbB9eK0d8o1Deo/NN/6Y
NXCm4WHM8nhiyR5YpfcFh3JRONZXCf5/HDng/OySbodTurnpbjG9BzAbMoM533H7/HUozawe/hB7
mYlqyJP0PT/QhinHlh/xAyVQD8h/tflfOY4LrXE8S7ov4rig3VenSzAnId0GnjB1DaqbPPB8s23h
JymlQ2jGKt5Buc34IpUnxVY0ko8K862qnoN/dIILSu2MoRKqJsdzHD3X+151yzF1yzzHwGw/hdkV
CBYAn2otaFG5q4v4oOzzSXaeu6timCzl/PbqCdfYqsoyfSnqKWBvMG0Iw5jy/YPbg5VYpPjPfYey
BHKpwIN7NIO3KKxtJhqmG7dqsQJbzDv2Ps0eoqITWKKhBAAk2ngBr4riYbkKZV252iLDUYVtisLR
pPvYsWcTuvK4w+yBIiqr+ydiFuD1t4kOdK+9Wjhk7frewIOREFb2tZuqlTbF5A8Pn4hL1Lihvgy1
o9ZwNg0z2aXPQg5ibNsDHoHIM9uTMmZBKsa17v7J1VrBFLlZh1UWaDGSoo9fOP/e6nyGRehwsRZa
kIjxowYgO+b1IzixCdUEMaJJFh+RnmDF0L+PX3zejHrmpH02Xc9+OGMEB7kNJkNNoMvV67Fj6tP4
GxK2IlwwttVG9MwBwHLNpcU8MqZZ+NA1yLD96vv8WEidMQM6BGtuI8ZnjJz8BIYfG9XRu+/w2Gz2
kO8oCtWQxzxh9Yrfc3kw8cR/Nla96a1I42KqgUjYPZDZPCtHEP90IEaWaKLxDJmjd300uyM2UE8U
i/spTDzfE+IHnLzhHpiLl4kteB3nCaVwsP3Zyyos6ww7itXvSs/FaqyqsAkYuUSJoyBGY/xC46ri
Tu4Wb7yg6CY53eXvaWHEHzK1/U58E7QsOv9WYH6Nfxdrf6+so+cCIVg73aVA18OJuUZSaX7fHVQp
0w4Mmti49IzkDEkVLYHPCOIt16mNJWBQmTu10ppdxTn2lH/UXNucwf2WW99syAOnnDyacDjClhcm
PdD4vjPiEN016Y6YDm0rjYxul19N+q6PmhJaDRenjtxafEQ48/fWNAKOX0ccDIjAkWrf69jE04j9
9wLlqZXi0NNdqqMv0smue7m4fA+mwhWQjnSRLCtW5yFYgGpyX83/2WTLX+uWTfh1RM9cPeurYEVG
RrMAQBao4+seLLhOc5d8WdcL1DB+/KWyvOx8tGgA5pOsXKRgW1xXOGIZBXHq6gV1ltS+FVf0FJ/D
rblmw+wVId/uefgYndhxrHNzhyH/CGwhl0NVx5Wovzl5vadIH84ugPHj2QwM91MDJ8Mrs7n5vdTw
W9gBMLitVacP1IVIf1teDPZIDOjfQcE+UJ/gOkwdLHFRo7kDAkLqlqfsnVfHEDjPD6Re4KyaLlZv
DqvwABn1tn1zEs7zlYrk31SJ12isDwsmU/xfDslwQBn+zga7OqkmKqoQpss60uu8jQJXapIyRA0J
EnYJK6iUAwX5OnwyPTprWrdc94hi3UXXs04/rpE3B4c1LXfGXY+htr7kdJcWyW9WdS/+ZRXMK4po
MS7NM5Stt1Q2S2mQbgpuZnvMOaboqgU0ZoKck4z2o08NIPX59TCFbjdahgPpvxT2o8mS1L6pOqbz
X4tPIp6blZyODV91yKsrQTAJuXQVZdQNIVmhYRaf7Cc2dTmW2Pm8QqNL6906ui29wKRvA5aiCnJ5
Kc+zXouyN7pjkSZC5i2zRwPHqH15MZbbu78I6DoWu4lE51JrfIi9/f4ncojqlXdccz7NodlemkeA
aIaefbwkWyTCsyJd1nMQut+LHSqAnWYQwI5NZ/D6c0aGPUIyk8sYbG4irsgKq9diwrbehc0kzTon
8LY+DvkpES4/og4zKF1/cETFs1YahRufgGrdjYCd1iM8Yk+PSpCuzZPEGY6FaZwA2vvfYAFjspzu
axkK7//6j1/3/MArzrB6Q9DjKlKp5u1IgriuWe4ir+jJumH3FGBwGGdUNDXGmBKReQMRVUrB+Gdk
ofUDq+RVjhQzXmgWTahzjzx9aMd2dDXEk/iybytmuAW3V1rZ4HqcmMp+LTsHWxGo3MIoV1+OHaCA
JEn0oOc2yZHjFJLcBCgYkD622Qni5VCR0CzBWNNThyueHrWMJLkVRjIflYmd6oGxm6WEDdOfoUhg
Efdmp6k5NGO+cxADmY6S2JtdGltJjvwv7KCRl7eX2hBluNVobAKXtQITwPFXNK+f7WyYriX3JMlT
S4bB0zJYr9I6NwVThgIlT3F8cStsW4RoNq2tkkEuBbBPkeVYEkmNy8e2VcMFbvYXEq8X9YwMj2nY
XDuFdwxbzOMZarmA0kWnMu22tKOZ0QVMRV+DPf5csG5VO5feu6to2JX/8qCk1XiLSUFtW7dfji2F
oG+tC3p4KMf7R2b+LMpYMfnTUUsblkiFH5wPNVHziBuEmiEeCb/8Tq8NluwdmEFlJWusQih12v9g
9V98njAUMM6cX737zkCgCfKROLoZOKxTeVWX5clxDLmgGNDPIKLDUuMyTcjVQjeA21MiQO8SM3jZ
A+JyQBxUorL4GdL1UTjI+6KCjH+oomyX1yAFJ+0DtUJhT1ycCeGdTxrCrlrIvEl6ioj9GazhcGZ1
JRn9jQ0jiYXWHd6t2Wf8IBMJKusGIt5StHtdnB2/sFLjBGNq59TGV7y493v64ByiG6ZSmGrDSqwA
ywXlEBknyuyTN6eL/4YHS5NNtSJl217bLrdEghJMVbR9czTvFmSAhznDkNkkLdsVCyf8hw6MQA5s
DdmT7UvL0+C1hp9EURr5UkoJ4AQnVS2is7YZA4Jb1E6/RyAgnbCMBqC8/Cca7ZItivt7SlY0Y679
PcqZQE/uDzSTOLt9qdK8L/Bk3u9sdMw9joFYMlXLdVprWNTh+gvqdNlEIxVdFfqcry4QozD3FHMG
7U5glUr/mzBBCrMVCQffTUiLchMzfVlxDV/XTKOs3IfIXAVOYtHWEWuk7yXH9NXod9jm+G/AsH/V
+hV+IqAIIMcpc5QUparA9pNV8ShuyW+0yeDqJtFghbncVb5AMslBqVvYdmq6PYIwCcoiLirP7Tb0
pXUErvYu1YHkuT2cv84yzlDGuoy7cUCy59Loiwn08O05qcDnOudOz0fEwWzTtAxIhpiQQdqm8jvA
bko6ItwpukrsLmRbfsarOXQ0bc4cjBUXcJnStoaegCDl8Yc4XcIknt20/nC7Oyvj0Bt7pB9ZVxxF
KFjJWOrWJa4rAqqz8pEcY0JlIDfDlgqrEr83k0oUcbIZEbZj1QA4bhH8k+Z4GAR4GsBPumOEDRyD
dXTSulC8vDeh5BvVZpyEYx8eKDNTKrFHWwcnZt70zgKnlsq/mbIwT5WRk17Mhjzg3dbjkDrQyr1K
AH+Bew23v2Pb7C30UydwSCbRyfnFu1WFrsIGDulznSy2QslOQCfT65dYadPWqCCiVCnseFudEgwU
dO8s6VjE9y73H44fWoN8/9Z5L6P/RpnD46c/dat4Um0MA0jzpOXjP3PRVQN5RBOTUifJtiguKfus
JaZ1s1T74Oq9wc4YJ6hqsgCsjJgpt0n2dfcfl01lnDAEGDUabvaq7csrfkJx2NgWW8pOL52wvV8r
nc5TySdnkLAAjMEUlpX4IbCzOJjGPgSm2NcfZiRQq5ReiwP7VU1Q2LMMC/TKMlv50h1qiyw9LSJs
8APlrr4TeC9Kw5HhvrWjXf0eFj8vJB4iRNy9NpBkUL/IQ+Vc6E21/52MBhKnMAuYBpFTkmxTeyns
rnbMk+xifLCDnHzeGWNgsDdZpyahOwAuBclmC5XFXIgRk7zloyMSuOiIUUWmhk3RzA83MF3DtSm/
IAdf8xchg8ziZWB5UxlS9ZkpVdQiz0iVqtZfIYAMMwEZXW6yTlTScNZQqe+L7RP1d0ygpmMhu7jT
oSpei2+qsJyGtPIR/upxcpV+njLb5K0svL0Ck5DIW2HZGRbzo4DhNus3YuWcKnLoyihuw2q5FzzW
zI00hS42E05dbeBnEMA53vijKCfuIFIFn0s5XZHPmACLIPrMbnXg77A80MQrLbgd8+yq/xJbLrDI
CRtCaAZZ5+J1ZBi94Vpf+j/7ehAy/0kY3quMCKW/yqqMUSCPxwMderi+ouE+LIEMGvP3w+tn6Z64
3umeAaf/IxwS6egtdnZak9jB2xsRv7IeGIlS2fdjPzipHbwgAx3swfjMSucf6JN1FQGvhGBPGZfj
xVhupzg+vwXdE1ftAFfKl0OIVOkyCR+xm99ZnhWSP6v4b/vNlVdRb6NpZs6aX61ocI/6p78LFcAz
3PIftXDtDrUDhWbkzDzWXNY++ljCN2rDyyv8AtPEZ8Ibqs8vVjbPUn0i35I6sLSNqn8KDvsmD6l9
omhQ5dXJypInV6PE68xmDFniCajvAiGwkDb0q22KHMGYw3ibA+8opUd1PJenRvpuZKdwHv5Lyic7
XuQpmJ3mj8sJ4cHnP/E8DyZrLEbqT7TGg9anWMjsgBAs1/5zxYJ35bQhd9xlNK6X2QR0lgCc9p+T
+r0rHy3Fg9GTXmHf1iYdWcA9/ZH8flHR1emxqUMctKbBZb+pbMVlnhCNVEy5uyCDoYZKi4XFwoef
FL3cRdXvwSggzk+S9L/6mUcvzsihsJdzhFo1t6E9P/DqlR32j2tAdRDLFsI/OojGtWTKS+yNMspe
32tu1gtK66pggblyd5Q1fsnibKl5VfQ1BkbEllYEb2DVimEBwAmiLgi/TgTjtoIkesd1sb+uFave
SI3K8id3JxAWxdo8/V6m3A7I6cM2MhdlcxmaLjXJ5p50aFScE43+ZcSiuen3ftaMKhroJOomEf6+
xIqU8lq4Qsw6NuQ89o+aq57jbnta4NG+uHns1PtWpPoq3V25lAuWu4RxdREw4q4l5j6wDfshyvwr
Xzh8J7d6HYaSzBSPxd1YWkxSfXm2GhrvdlwjUvKAu4FhLI9HmhH1Eam0ppWJ5+tJcOBQbd6PIkxV
qEhPB8YC08iyL4xm3bZmkhu+iah2MVtinlrDkZru7ALa7ccy7rky4mm75SmMYKbTjHEYz1QrhGPt
cgtOObeAH/f6R+Wb9ldulzk+y6mPgMLqAgX2yaIYsLSHY9BFmx9M3t2Zlxq+OHjJxML0m9pqSR3j
SnZKwjkWGXdx2zPu8Xah5hHpvUaKxs5JUiRXF6oyyS/MnwFEz+E622fJILYwrl+AQyDQM2BITFm2
ZVBtlZtJd5vFpdgi40+DEe4fQZIqtQEoF54P4l848XAJEHfBG9EeRnw72g5QxQa/i8ImOP1r4ieX
DzQdS/drHnSzsZQSIYLRwBbhp+2r5Lb62pnd7b+DNSbXI/y/kdKZwS5xUToh0A2EmpPqy2sGdqwZ
P1u9MZ4XMlWYRbA18t6iMLr3u/eIP8Ra0zOrcOYhDMLxHymfNOCyE3an2VWfME6FSp9xvWeyj51R
dG5o2O4jpk/pSgz8jkOjCUZXKpMJzWvefVjc+OGF9BdviG4eiXW25tU8Tgsn5z4AgdiB7V2xBhDk
qwbE2f2YIFas5Qd5D+bJUbfXoECfLejbR/Hn61AQBdWAx9e2c46tnqWghkOVvplkKnkBZ/XY0yey
K9eqe24tsQXZIWc4+4hbgT9AIQduhmM55gEb3y/KwuAX9P0b13PL2RdFBlfU3mFc8LQ9X1Y9ekBV
Wzo17eigY3PP9qtW5wnmuoQDvrzNVIyQnr/aJ4/IdGAsoYKQyzrHxehHxt8O7pFXk0jjEe3EmTs1
KUi4Dj8scMm/w0FxgnOiZ118Y6//OBW4d4WiwWw8oHYFTnzwfb/EV9B7wslRo64f305J0WNpsq17
edDGaKnK1u4Xoat36e9lFQSsSpS6CA6WiZy8b/ZrFCpFMDFmkfpbBdM+eVyjjUG04Z1RC9UB8tQX
HO7X9N7Agtg/antonmdKjEX8jov/JZOTWiIwO0NR4KH69BTw+hXm5WgOSi6/HFHx8RkXzYHPb/Za
uccEDMeaXJ7/05l9Lvxe8/5F74yc6eFPW62BjKFff3Jn/r8c7lZN0Y1+s/NL01jq4304ghjEQXHN
wCIBWI/DzSFrk+LHJFkHCB6e+F9tc9lDUTw7KE5QR4m/NEDF3gQDu+CUj/2xub1pkHL91iw27pJU
DIRU7rsD9C/GeoGmNCDc5QjsmNEH2FDGFhuS0eyEQcQZQp4XDXioHCJmWpOLzGUsfRjKO8SEK+RV
7+Cz4GVqzC/Zod/Ta3AZ0fZSCp6HvvXyG0aQgrgVgdieYOEWzpJN06TLj9hGp1/tujc1OphbVajv
rE8pyteuCxnIPvXLrk6P2f60ldACtt//5SK75z4QcseLceawW6+uTcy7g+SzIawbu7885nXgAAKM
fvQK8QOsPI23NswsV9LpmmoGnbqJNACBwRMOyH9AwdeEUhpHOz7dkBoWlgS09OIx0ZQOdgP3MddQ
a2VhnTT9blscsM9cX6yERSTk3VDPVsEUlMa7vST6XA8VQQfJx1yj+9x38au2baL93zIUxSbbYKQH
KAGdSgsMoxXFzhFLmH4frFlbeihtKCIjEo+MXX2O/Z66c8NR0m9X8VcgKXXKD8Ly/IxqUkzIXGcu
wn5uszz841ewQfYoJNfXB7yGoXthrguv8Hg5+3TokjAau93Y+QtWV5J98qL5mC9ZvLCYhrE353mb
cqlcY+lG1b5Njiuf420OH1voCj/+NUeKeL6ivFGgTxHadQRiKraZRroH0C3CMSPxyGb7BUv7GbQn
2swMROLUndGnZWS/9MzPea+sUYE3QbnRSOyCcbuo4J97agwpI/DQN1vLvhtQmfcenyaei5uJIADd
ex7D4f73+brKNfa+rmOY1c5YxCAvQFxOx8k0sVAyl22fTvKH4vtyUiOvQZXfct7ohZwzGKrp4rzB
PAsRFNk8rXsboQ54/2dbLxSLmtk53vd3muY8M+UmnDdnYz+bymkKKdTq4NCxEGo/yu0nS/9tN75a
ZWDOoMM7GC81EfoJnyFg66jFi7ogtfxbC/nEYsY8h1/Yvjl40GSRDzqZbouopQS2RSRg6/LG3Kgz
eEoGqXywVBK3jSm97SyCSyDvFmcett9ZGzMrOCx5Q7wze5JrEkWB3O45PrtSOOrUwKLjnw//H6T4
qUy5jZQISZN8AGynmCJmFYU9PilOntcoaZyLmjM4JAlLmoJSds0gaz6/kxUxGWJtWIBPwQ95Vd2c
INcqawzlsUQARj8m3ZVt8/YyMlVWTmkjfAPGPZO92wZjTlsU8vSBc9V5aJ/yv/lWXhe5HtAmAbpQ
nm4dcLgwCvsDeRj5FxEbdxq+hJ6auLkqXvPznnC4reQUPYEUSTomjeCOIc7cLmokVh6zOKiGIj/U
0eEK77fyZPpIOfjWh4Lh7jKl493UTCv0HAJyvuwdmVLyRemDr36l0/9nnI+qmi0PdgrC99VuAHs2
Q7vDB+gGi7rOQ8AiB7vc4qzybArUt3Pn4NZIWYwUtjVfd24K4wto46ca7ObcsM2f7Cn8NnxZelW6
9kLJtAOnzGOxuQE7y8A9pzysSeoDimWic8BioLdKwDoAxQWG8u4lOprX3QQqoxD75euBdMRiDCJQ
PgyJ1anOwbn0ROmGpPFuMZkTn2uY4oiRTbPjgc7ztHbBsgPoVsD4HOXVeK7UQ11oB4h4PreCQlpX
YxXNldqJfE0ccvdupA8WZo4tjgFQkmafB/KZxDI5/YO1VK11S7rXnousuRkC90NyuKI7XUGy27Zj
6jdZWbv60V/asHXFtVHz4kgsb8LNykgwgUzELc96Ijh/cA9W/UuylKWWaMsRRr3hQ7Lgz39QM1wl
BY+NcKKuoyx+uiq4VsddNeoFHw35fX3mL7ZZsD244mbTvFWEnQT6vz7wpd2prdYBy+A0R3rFSbjx
jhw0q3rsl9zMHxF9my2ctrwdErncKlxFCbu8t9nipReFAlOqJdONp2YBe2lk/JUaZ5C54edCt5v8
pHIj0k+UMkMfdCI+2/ahgtf+y/qGRjKRuR6skpgju1szlaYntUjPWUnqqq386PIdJSkI7RFIPQTC
KzJKz0cWripZX8hZ9ASISmMSHA4ByXB3CG7WK9lBAQ/BlfEylufQfhrDDVrU+S1myk2WJXg/mcAr
vxMMNp7ouwbZFhN3BA2yBZswqqTVT3TkvwGfP8+5kIWxf+yjlisPIIaw+wrDBtgbkM4k6738zyp8
AncBUVynNF/edqLY7KtIo1X9mwC18ocvYYn2XcaHWrjzcmHfHSAu5L9cdC5hcNJdKsXwNP2f3gKK
mT4pu56VDizC9dTga/TvJyhGbSl4eDe3T+a9FrGcpA27naHZCuHvz3+azcmhrEwI03lgb16vHqZx
bdBHQ+PrXHBzRFQLzL5HLa4u6DKTZuVjVDy+u4TOP2MOSnCpHM9kKIcZbjiVXwv3jDW2zgMv0HHL
J4G/275Jb8Y6/o8BIo7ifJuDj3jlHoHUmxKsErp83Oqp1gTHydCYQG+rOe+f2OlBDlM4/FArKR+R
g30RKMx9k9lMszFMCMCgsvSL6yQpsMv2B+b0in/32JJflMODB3USjU0Z38pxamIG49Y1yD+uoRmA
9DJuxua63L6WrOUBuU9c2dB38yi0rtD6wrmzvulg5te1R1nas4d/GGUloakN6TiFUAAxG5oQKBs7
s88Mz7x5XkWZAof9nwpIuBbniortKW1Azr2G0VXACtd98i8fwOMWNnksFX0UpJwrXV91NMNOFcBw
38Ui+hLBSx3Q0MWxbSXhkQlO4XMlYVVXl7Yj53e7u+a54+9wNLEgu6HFSZJ5OuwuBtb9FlahHo7J
vKAZ3JANvdFUczUS+JQHbR11r2VRWA4XJ680utcwM71bk/FLWDf9xzZD0bNBy7OVQux3YroRUCij
85ij25odIkRvU8pJiQLtpFtFqOQSLsP+vUv30+RrhY1fo+DhSpEUObif+cJOTPKy6blQNvhtNOBh
AGsRq7pFcQE6jX2tUu6O3gTWTbqcWEkTPMq2xHLgVv1MqlBaL/oTxX0uHwrPDg0LNhU67n00qo0h
Yn4De37kVw2EWgZlyCcw5mr7qerUe4tC7g/pXxhBYHKo7QhHdK3Up+9pjvYAbeq+tyXIPSyoMr4N
buGGCfaLok5lwedUV1BwRsxqsjK+gQQ+sUvQ7KqUru84Ap85YP/japkYTmh6RUU7mcitKCNtoj4P
axNRAh5nbr0GgnH12KLln0HTFVWAvrp+kKKWupWbQuOPnbrmc7ghWDg2eC8D2sNwJmiP1BZJBsw5
nWvkq1m8lQeJIyZEdZG8qqsEeF44dsBZpZ/CbwPI2u//8Z6xU6T7qH805GWT7aZrCXwYEWcw1lcw
T8B+chFtlEWCnAd+9W1+ZTW49sDG6NfyrlyZrfbNFJX82BiaFFXPrqw86kxXdaA5OLA/iVJBQsgW
aXNODoQqyMP27T1j9Q8iKyQ8vvqZM38fXz7egiXxiUw+AG5pcBzu/5Ccg2UnQhMR2f7bQPCkIFBa
c0vBfi0WL2V/Z8PPAPwWcws5JPwYK+M3dogRIHGkjKwzexwhbjvJE22O6jyclCv8to8FmtmFrpP0
j2J4L8sf97DOscVe1xL/qhE+XqFLCXnGCE7TYfwULV0Q4RxqC4GitQsDKPQ11hHiSu8Gv0vOuBNY
JHIPAIvqR2+6dqOdy8VMidYpfYmiTgghiWtmphV9NatHnf0nHk/OfYsDa18f5VJ8y3H1OU2q2BkO
qL2zrT0c+VDSLAod0jHFnzp7goolSrxRk5LR3hhKapxt31IMzm4L+dmPUrBTYyE/+egyQgzjiXqt
QDHxa0/NhFxh3WcvHiC3RfypM/BEpuxGQn/QduSCSuSNsLUadYCudsYSznTZ34EVxNywA1hyPCGY
uRmVomIT3zQ2NSBH9Ve0oumFa+nJPnGgfNejLQeojFYGu+q55CZgkH6lKHtKq8bk1GhG3w+QA8UA
5TzFInuWMWJBMa1Bc6HWLCkkAJW0eI5Qyi5Zy284V+gGKw66dYA/AyHHI9DqyD+UCTsohNxW6AzI
j6SpclpkoSveSbvWWWUIJRGX/hc5ZQy6rw+IZCg2Fz85L3Q2dF+J0KLpxJOT4xqzX8G8z9rVif/U
kVlQ/LSVLcYiouR0DrjomoTCScOhXbrBmUzJ6GrDHn83JpnuymgpdepgOa7IJqity58Dmjtq1ivp
kejraVJOUvsFstSFhsCdseM1wZTEKa7WRNGo/hnR09aYqDiYADaQx5+EYhHlUV9agj+jmrVofq8q
tfE4sqhtqZE3ILDsZWILVussVPEr0rFPrg9cP6SrJ6BQZR82XFhS8uR5AVHGSQaC5IGQHZG+tCDC
anlp21YrfpFs7nnvxGqoN1+4tk9RuSnzpeDWeCNPNB5B/7Rqrqyb7zco4p28o/TN6cpcvxsGs/ut
rxhENkfxaXYwUQVeKlov4LVxx/lBupe9Rd+FsUAe8BXz2eKtWbYJ4SJaIO7ehg/7N0ofBpbZ1Jwp
SqNyMOZKbeBt8jGDNkOjwL+ThaMMGclCgfyc+m1M3cMAz0LnG/5Pv9YyAJhEdqs1srLMq03nPTWq
zypmwiavQ2kyqI2w91KLMwVmxNJLhxzgnO9s0yrd/gmTyscm+2hb1KYwTkmJ0RqTSCrw7VnsUjS2
CFDjDKnDX1TDrUT6R1oVlTF2afzQBe5XVYrXlWGQl5TktRfb4Q+zUqe8fniJMxW/8P8FwxK0KcYs
wn3Q3uzEMcMcFECfWyesMqpFpof7PUms2BJ4xyAuX1mXq3XNjlEPTDIjl8I+T+MvVN6bSio1pQTL
RbNcbafkIN0xsbWRC3Qtsiriap4vdo083nYYSo6N3m8Fxe1S6keR/yLvtF8hh0K70G7P/3dAXGHv
ATMkHGFeClttva0sKzeKy1tcM6G/73gr8AdBP2/LXG/tImVKzr639mGvpXvvBuVSsvMUIt3wZXf0
1LOpOr58wGW8mf1UYHoZLgscyHk75R5UoY3kdJJVHT5dggN+UfAP4yY4rKUlBe15/QrsyoPvC7yW
cg73HN5l31y5aEvCTZsCdpgyHYiLtFPIJztBn29lRtSNhyU7cV505aFycuaQMo/jX355ZCxm83ea
5Yk3xjApwsqVHdDyBjCqPD2Wkv1iIFSv2TiK3CO1hmbaQW+zlLOGf7tpQeEL1nL0+rWRO88Mt5JL
zJFO53O/Zp7U0eNgq2/z4FpKLWSmey6vF4Dd92TkZ0smr54reXAvBwybwuA4odQR5zkMjh6ztATA
t+p2IUSt+KYZvlrWuWr++x1CdHSrXiJvNDhgHxlA2y79E6i7EY0zQ+z/MFZsJz6ITmUK5Wb4KyOg
E2y4+v06UgiKZ8TuX03+5J2wYwvWF5QzpoOy7UXjr0SIw1eNmmC9sNfxMvMZereOH42mQCTOteXU
HbT+6N6t3NgambItI1Ak75cxGLPHS1620fu0zYjVRwqzImjErI4E3EAQTTofKhsh+7gggjWWE5iH
zTEwpmYb41A+UPr4QL5XQEP8PFjymRsrhpUfsUq/BD2COvvDc7LddC8Sw+9JilA6CMIli31lmrKF
Ui6tLZGWHwhfks748IoBb/coQ8tCP05/kLh+J4gmTajKY/tYt210AA451+5DIUPszQEDfh8vh9g0
IfldcqlkaZj39F6olFIFaUieZ8a1i54mXktcBUW79bSJ366TQofD5l1W153nL8z3Mu5TTxjJm3zw
xrfHgWhRUa7megjMBHeRLtSiTMB2xIUwHazQ5RucN2yEPqZ/l938KmrJsa2O3PthfX/Au0Nbp9uQ
JSN2Z+MOQ5QfOgeYwLilmGxD1sT6YIKJFM1e19PcaccTqOtNYTar0SJg/W14ffCVpIyiMM4lRldf
x3Wbe/cu50TutjW0Q/rx+l9NsqOxCQJhHG3aCFSZzxrEikK/AteZhEOG2RcaVr1WMA3hJHaDH672
r/RlHKKC5txWXhgSmqrIV5YoAe2uGPOdVJ/BJNuc4odHzz7HB5DOmqXzoFtLJEkFrzzvJs3KWxSl
VOJjcG6JnLdRjK3Yv28SQ8AezFOflLy5fmjaMRAIs42fIe9nT2V6hXWxyZBYypJvbOhXHBsyy8V1
Hn8Xcyz5+uArPPZF0W/lsfsbqvMaquq0BUhWa64tDdshhDWta7D5oKCSXSm/ScG0w8IlWkHyh66P
nC4gBN8wcDi17xBmfe8pTBabjfclZ2f+B7IzuP7sOCvizGhPZttPXtsRXcadvO2HIySe3EaUPVWQ
UlsRlOMdSYkjnE8Yy68EzcO+PuT69vh/OkrWe8TftYKWRzFh49zw8hDldd0S0vItZk45gdA4O+HL
ysiOzxXrwop3w4Bna5pSgboR89H63MItIl1WLRedqsj4E7qXe9p3knzWc2GLbZatwyahBsFxtUuI
VYoDePYQl1bwbodbUJ3NIRL5ZE2jIkOemua7UfdtWoNaJInadZlA2sjWWkU11fLv206G0IGMH+VE
pflloe7otilkONY4bTcFE9amWBQHBslXfb6EPUDQSJfiSe31l5sB09m5Tn3TgdST3pm1/i2lOyGU
UtJmYr+31eSN51rijODLB4wSL17E8gav4PKeRInqXB/CyGLF0VmVtZjIRhh0Y2AYMhJ9uF0hVlgI
9CL/2dicXd42NFRhIJ+SD3HqMAt+NQ9QH0uRbRmHrTNIfDcAHV6rqHVQcGea+OwyZZQkNag2rDON
De5LZ9YF9RObfkeug/uJoLqiv3Gs56gCBombWbuQ5Kezs0DqwsgNzJW2loj5gwxxUZd9dVYi47jJ
AXN8lomeCrQ0XqcTtZUsbE/XU97Q7v81TAzK2tkLT32iXpWzVIxyVuJhgNXtqkCABvVJLEphBC5/
6bqrSUOosN6yKT2o1kDWeGPmf6Bc6/M24dMckL1Gg5c44jkmoa12IL2aqZ8OqQ8QqwcndA1FOR+R
IPXrG5tzpWytrKNdbY1yDokzp4z4BBrdaXEOP6+mdgtMvPVTD0eXh5ObWPVzMq5R5ISi+gTCrt+I
3g85wXmoTzlksDJxSr5c3CXTTjTgmvzNgRgTyNuh2ggI3uu28tcfyYQ8kJdN9akKyT9hNagZHdzl
ztPwG6B9DL/WS+eSZIrIALb/OC/S0nbyOEOf15k1c2GsJ9hYKdUln7JCchfq59E4hB5DjPvsNE2R
hvVF14kNZva0i37hZ4JSdEs4xCnnDZffXRCczdlK4lgnQYUZrfI+22HtW8FfUpctmYEJu4RN4rY2
0UMe9Q1E
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CmfYEHNItvLy4TKvzFWgvxDy6AiUtQifYjIjZAFSN+cb1WYNuAsBTchKK3PgeuFu1cYW8Phh1HBY
f8QENrofS8ENbhr7YxJ4geHF+1Fha5IxSM7qnwC3SLfXoSvsmsYORW3zungS9IUY7fjPzBPqNpQr
b7i8moAyjfrMhqawBUdpRg+Q0NJnehgZrP47kd3cWCEnznalmfSJDbGrbIckc9iHTw3zeCbM9s09
a6RLkGcSuyBtsAwXVfXzXkXFExXoNge1a/OUz9QQT9wzpAUhRqByjG1mISAqfoVH741YHGuy9mQU
JovfL9BmMAaKddRQrn1Q8/cWmSxNMYKFOMLMyg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6256)
`protect data_block
4BrK0bpuBS97mtYjH9Gvc1sNgYXCO4w49+ZkafDDoAy6Uaz+hE2/i2vx6dmzO1fXBQ7WQgdBLhkq
WyaSbGf1FTGrGkeoGcIYqN8waLhSECo2ZkPb+KgJH+QJwIheqxBLmJgGNnymlziXCnxnS6Uguor1
2CVdwdjyw7mVgykCHUSZCVyUghmlG/dlhXTpckhR6SRuE0N2j0vcyu8+MkJbt6gMsD8H25qxTDL1
jV+A5+HJvZamMu6BFdWzLaBsVjNOe1ykvETl6FbUjOu3vSJ4GvKxdm6Q5xTmJL0DQzTRDBQg9omA
sY8fJoyk2C6ShVLPhGWsucAqF4gHYRMWfK/OncvzVOXxSXQdN78JTErIdYZH8q6dGx8m/XEDkPbr
bvIQyuL0CCiauhj1s+052tCc/GbPLd/sZ7yTJLHXFlAbn+Ah1PV2wfKW6r9lhxksF0BDwszo65gd
VO+1Iu4MnXxQnMwh7BMdTlhoneUXHTqAVLPCzS1f+LxMSBhtmyMo1FFkij58aKLoUUxRWG66ACoS
qI4FxXYN9bMbSnOtrdUHdeINhaLgTKIwWALEko2jWmdWe4CBeVYgt/qK2bEf0ImoJJCYPHIuEC2p
Xqp7HsJ3jqiWWrVVGd29Bm1gcdSqJnTFmklsQCiDqGMRfSlpumxJ4Rg6i0bhx9IVcvaxTeUMflM3
x8F96y24sADsq55xQV2uWUZBdFE9Lzw4MaosFKFON9KSQ+rg/FooUasLnjTNxMTYCK3X3SGisVIp
qiiX0c8d4BNDspBLghh9GheQtM0+5eHSu8gBNSC/P/Uoo1pHft1Qm/ucD2YT+fcZrF4fi9rrrIO0
8vIRDvBJOsd++9+RMq+ICZ6djF8xLgpwmBXmBJ78WUi4pic84B3ChNXdIklTMW78TV2A9X0ku0QF
P+Bab6OtWsFh8/qIBziANBD22gurCq/AR74yiG4brdU81dw+A9YPhXvniYwc17F+VLrI/Yzj9Mso
Axvpd2qotyFpcLBFyIfzdR7A9hpp80+ZmLqae2OJa/NN2jn6O9+GqMXK/olIAe9XVszahycluRrI
mL/7MjQhnuyhURHuYnUTmr46oRMjOw3RV6u2+erDp6y3bK/dWWK1CwXidDgVUeeoF1URPybMYLWn
OlRDFbR8O4LwlYf0Yf3uA0YjjyBxSFq1ph6RG/gQpD7GXrOKJh50BuuquVnomE9nTW9e2M6aFHun
bnMVFNe4AaoGflp/MEJvcBzVpXQg1+1pgEJNqITM6rXsp+pDqEsNXcXO8OdIxEN9fXh2ymUaieNN
gNm2FNwBCeioOkJc5O782bHoqKDVhdUWOXhiiREjBHC6C/D3CeQVwOv8UH54IPZCoebjr7FcB9/J
R5oH0Bn8HgdzCDmSKrDIr9+2wjGgQWsy5KnkwmSSsYeV5uqerAfNL5SMgswhXmbsys1uEETUjzpg
ulPaNjJolZlkV9EvUWKkQpG88eCPLbCgmitySoCIllCSEd7LqURrEgWCWtxdH3GKrSaQQBCWXO2N
X6iiRxEJJNEb7T193l6FXXMfZ2JkBKvGF/rUiIWStM36Hl49c90lI3DQtqw6pcXBPdd0vKGEuFqX
2cfRZP4+vdC5UIdhETr2NQM7Y0j825hZV92LN+aPV+eyNWzQkorWqLcK8wYDov9cSTXztA5vNKlM
YMiAC6z1jC8gnr5QUX8OmhjU0DxTe32NCvUjVoOUl6qtZWqj0Sj25IdsmRL09GZifgzCBgx9wOzs
do2DkCqazWHzeJn55eJq7uRagt188HCAqmOinAVEE0Ui6HJFecupN3a7uGzhXHNsIiamrogJTlDI
afWti+nx53LJCO8lvTxaXhHaUrOtzRImhPJQZ3qHk8VRlEZN9xAT7oxqlg+gB3PjgJTwHT1AyZ8Z
45P+E1wxObyzSSNTqFtindy/SEj+X3Tgw5DDkF5AzkaZkoA7fWPuFbvYR1xuGLiPvTp+sW2WpP/J
QTIGXEuaKIuQVkFzRkPrn34E0wo/J3aOgTSqpy0mrmTDEPpVlgksOxXJ9Jkb2ZW9UZZqi48Pp6xa
jxwSt46c07boQKFfHHGunBc2dROgN9kKxo18oGwR9j4BOgHoXLJnqTcSETE6040W/mC63v9mk9Il
O6HswBQ8OjT1kNID+1cm8b/uLE7t/WYH8y090J8ZFPtk/oOB5upgjMeCNWveKmIOxnV093ugYiN/
G0+mSJ7EX8e18sFWYJi7/Cnvi0bSCr7LxJGux2CNDAflqmkTqn7OCRyGgFTAeSRs9nBfx8ReJu0D
XUtNP4MojSRIjuz1+TBUsqKQTYLDgUWDMitkV+RNfwk/f0ibJWuY3aXBaQ0ERd5hqn4JqgbT55ww
ZL8dFDxMu4vQVidqg0uoAK1Ne4K2QeupdPS5JxSeXDQtPhZ1OBTYarHoZQBTbKT3IXp3dkSrpemb
So4TFgmUelUnwArAAP0OSia9EAmG9RhUFpfx13+884gKrZvqoBYZHphdrgHE4AGwq0obEUOhf6y1
WNYk8TOHJUawd17MbIpXabAh7a6oXi+fztJeZWiJlrZU1MLz1euLFHHQGig643v2ReHRCfZwQ/vr
ZuVs5tLLeCST9iA5rIRtGSeuncnKUzkSqc7XCWO5jcFyvAsP0zLAqy1IXFtTrGlEwR/YnW0fX7OX
tJ3djkv98CHHD0XLfZntJqhhcb7t6HemEtbwRnGuQGRgKXa0ek+zY6yF7pF0v3NK4qk/BzbqvYLz
3QNKXXX33GBC+dAFRt1hHQAyXP/WE1z7voSkUTscWZWCbPdGabG00dW7L7OjkY1NgGtsEoUhQC0J
CF4HYCPvnTX2U9xvd/RPYilJ7Sbv1Vz9MwLtCfDM3CSa2XHv1FoIjyY/tom/IppQWeZSrob2WRc4
AS1pgfC/rRhYHL6Uc8pmFIOgdbX41ybPpFFP6ZAGEqvmDrUev9sAagDhJn7ad63VQj1xK3GgFihR
c94vnQIW4TxJegAzniNKB7GKv2yaxkiudIJbW3HHKrU0gVHbOuTW7+jKTqGYGCIbphQlZWO71mFW
2dV4lsw/QwG0NW9MExbgZNtR8XmQ0NNMiGJBcWWWUGqw9zwM5QI2044hLp48R8FI3A4HPblEiBzF
i0w1GzcKj8MhN6ocVR/8t62TllHUqzADvGbYs9vP+LXhFtx8HAJWNF69qb6Z6SHT2YDYZ51pbN3Q
oO5iXFjE0iCDAAd5m3EONz87UxdK/Fzq7HRiKu2Lc3HElynk+BtA/kKrMRw0xyLvM1dJLCp1D8Zn
1/ulTTmoBYVUEMxUWSRwHOyFLZTFUAglg32e20T8YrPwYDM/4NEuyrnaQXnC3HPx7KwJFDQlmnHc
VbJgeDO+PFrfAfafk084M6tGTGhvE7jEblrRYdvfER0jGBvcfTimqFIE4iEB1Hxj7UGjBi61U4LO
ARfL8klx3TyQo1H+Bx7GOdPnWgcc+c3rIQUvDznbrRhlt+t+3s/aYzqOycxF10Ou+4LnkKOympIV
VmnZG3ywrOT0nF7Y8q2rr8jGXM5yJWqcjRCFT1/Bv4hLY0POo80kjh+8eQ80HQE50INlwKrv1u1l
yjcFj8KTb3gqFo9RztdkbsVW8URJ1nOBgZoiuzYBLFT+qtgkDIedWX27kkVtvON6uzl7JYcMK/Lw
RXqFzQiKlsCQ8FOSmxROi9zCAoh9iV4/b7VYnO5mg1FCC9Jm3L7/zlCDEUBFVfexhD9lDk2bMPQj
EesIrivDnutKdgkuFcqEKZ6T+kXo+DcWVjH4N4ILSF4z243CfCBEhlOKZzsmUO4p+55Md/rsV5Jp
ACeA7vX1x7oUEef4vJcqIXt5boIHevsCRfUvJzv8EWfjQQk1GhD0YhFZMiQbIUAZbZ85lq3k+XuS
DCXArkbSQv+Q87E2II8VaRVd/+DyYJf/eO4rDvrXgzd2X1Iz3dyGuv6qfEMzQD87uC+lW05B6+0a
xX90XXjH89dg2RXfM8a2bm2Hk1sgT8ZzolpU4ONmISBGiqAg0qjEMsVN72aVSFXivK+S612686so
PQ6pwXFB6opHAsRpCGXb6gtOq7a+le4Q8DxXiE2+4u140BBTj7IAYvyHo2P6Kql1sNtN6NBHrBQ3
03lj8lj4Ye9s5nOWlZrcSE0uUXTPnMQXhiOGsTKGqU3ytqO4wt9ZgKMNH03ATNY1OYmV0ClLphNf
r6XVyWZBgOuoMY7hnUbj/UDmhM+F7zYs4IsMqSvrUF61+5lB0CPb22LDncxbp2Qop1V7DflBeq7r
loFsM3rGVdrCFIvqQ0w6+xqY9LWsDrm4Bi0lSkZoWQQMiCCTP8PR0FaocfkHSfwPUedQpgBNmMO+
hvGTgYkpZv//xKZc+D3IfK2PW5rVv2SO0jSc5deRf4TF8l4k/en5tfNwnxK9+thRLekDjzcW0Rs9
E/sNAF7MbjlWeS4f7OlrR3qLOLnvxj6mehNoNxdADWQ2AJ8GuA/xqy50behgk/aMzgY9Z3FYvmlo
ctIRQjkK1kwuTRJD7lSnQAR7jvtXyP333CP+7GYhY3hsVOJo757ctH3PrUW/7eFcWiSZDr9s0C8H
JW7TYn1GIpUEiS55vAKWizoN4094II83OjUtVW9appNkfdydiij8hIkri0NVtdvUgP8Zzcr03Rqs
0Zr7qqJ0a/m3UhCAav+Dy3wzB0hLYiO3GKli14yAdechfJARbvYRnM0CAIIy6/7GOpx/67ivdZK6
48hBm8nKUPM3JQd80lir2WSfr0+t9GyjWGzhh3pEIcALbH9uXTkLQZO4b8qLEiXn8QHntG4QxoT1
yjzaUFKCpvqLXAE5h2iQUseI7HS4JFkhLG2bx9horl7UIPsnvV2FPS3lswv2NHGFCOSfsVcaJ8Iq
q9xUCxLUoDtRTcfQdcZZ/sIiZ/O3YQoAuYVcGsSxKCNDJppGL5hUskUSQhRQoWhRvw1/eIQLeLqv
NC1yrAkvWC0Q4RdCFqSY0RpkhZMiXX1Gg9aVkTegWEqsYJgs5nhOUNygDLsQnyTUIwyzGXWN3xkx
RKYmz4Pb9sTTu22Mb5JWMjx7XpMrlBvt0HcCWhD/gM7VOzz6RYo7VQ/rsU+NpWZdUI9R/KcJdK/z
F3h7++GikROZY/kaUfhZtQsvC/A1L1klUaYGZmbVHaC3nFZ38R131TinxtZdECbaOpvWGjjunwgN
M1hFq1wG9hHuLPqQDI1538hW6B8NyKnzqlH3+VKxOGnFUJsvJutEp7vfATVGvcw7270Q8vex8fcI
ia+MZt0cyQleQr0CQ8rEqjuPpR5gKik9ieBB1aOq1go/Gx3kN+eBIDqI1X75aIbSx20k0HQ9F3xH
fDRf8YXrt9f6Bx1ebNsCI4GVVOGJftm+/fG4kzIgePHjJD669PrsM0mMxCL8aKdU/nQJhnzdMPHx
0xdFffOVQEye4r6ancpcEO2cnDv7O+bSmeQMX2DQajyxjsRg6SipAoNtnb7F+3y6CnxEvouaRHFb
MSMzsT659xOC61ucIFzPD+cFZXc7yLjAa1677UESmiOFpRaZCkb3GSw9uyOE37Z48UFoYCIDTxv7
xjXkMhyBCDtam4ZcJNfoJ4L4++BWgVz4ayX4k5YRszVLG89xUz6EihA/JUBx5cyr4i9PJWnT1YaS
o02eApJnNPL9ZbuhtLAvMXrTS87l1w7roTCy6d1bTtC+O13qlAOSlK6Nv+Fz5sfG1Fy2mX+arE64
A+/dKlAbOtORngCv8fzgBpX5QBnloHEvFCSCM9Kx5w/u4GudvvOVOgfzREGqCaxm2i4t35Pt9fbQ
L1dnvmV66m2jfYf+YunbsqsLJ8CWsYmNOfYb5lBsyh3UgD4+dX0pM7qK8QGvhrvHIqK3Xg43j4dt
0T5re6V/frKHBxNQEZRWy37hteF11/LvcICMMXCAFprRBpMnj9pAZRNPWxjH9CxTM6lmqB4uGKoS
TejKekcgtcuxpDsodnHLLHUzpByH0ALXYOed9Q+UsRctawNXMv3vcQdL+z7irx+CzqUsVq9MM92H
foAXy9h4XXuDreQJq+l2fgM3yWuo118cB0UdvLyfjv9mbLZC6v/HKhSQ2l1wZxIPAGVK8rIt77vx
wYlnUkzEs9jq6h4ymGvXRucPUVmamxvkAF/ooK23casE1ojVPtLDsJbMCeC6Of1qbzzVDxQ5sO10
9ClJvGPFo/YfeI5JfZtqw5jDAXSbEgqJp6e1QEnVoeC/wqjN8Y0tHkIwZZUB6Wl64FQemUwY8L++
koDQM710gCjmCouYhnUJGcFYgtEugn/BAWzeOVfyr+wPmKmnTp8d0dxtD05EAn2O1K333VoJ8cFc
MKS9oGCTcaXUzblHazrrM8yMvcXW3qo9GqdM0u8anZrxkagOVTu5tG9zDVDo9GpXLgywiOQ4qT+h
r3mRMHsCwd44Xix4dCu9p9MPDi5yZNvHus5sc/WOfmpe4NGSo5tKlvQsGZb3ETAU5YBjC4aMyIKI
eoRn3BRuY7+B2vOa56C9A2xkWDt4r0d557f/jdoWT5Gjrjz+bC30i+AY16mFUUjtyyTy2okKzkwM
eyBJqYJJsoYqcazlL5pwQ0R1KOPggQFKAYE4GIwjBLAq+/LChDjscAF2QUmsh9bMbNDkr6VwnOqD
ODafu7lkfSYl2azh6SkarVpPhpedXGodHHAqhi7iAksfPAhjHvoZRXAQUKbmvOfc+8Fk1BHLLelm
/M3BLVp6AKLhETzWc6jM6ADl/ibDGRl4/joRWHKseMOZI06TbLIaq3Y4wuYPOTMsNLOLN1RwC1KB
iBtPYWPHSxan4L7DPhUTg+DGcx6VNVF9hP5ceuyqd2ikR0+r0cYYYstPJwO8aMVOPjug/spiSjag
GwBnVppmzUjuxUK/cfjf+JDMedSZPlgnVbQw5yuj419bg9jaCq89QipTodHt0vhevviksk3SfDEZ
D9V5G3/Hl+8DunN0KXMCHdSKbHktFRt61syKgm4B5E57THsI/7K3x5KNcisDGHeeepCYxi014KhC
lmlNvGrQ0CkwzuRYC82NdY0sqIh0yaS5STqPLL69D68d1u+XuNyi6o1di8iciWx/IUC/d4scXrCI
OqbvqAE9y+yMTUBntE2c5hOsbj8aeJKviP1J4qg24dGy7KknTsaaDKloz7Xe5w32H13HMoyaKX1V
m8JbB3bbfaqTIExSYy9a8VBoKZ+Ls//9wqnqxDSewLJmv/2YAfMj3gRKCOJp4BFjJPSlS0DAXeGN
EJE1tP7cmNWeEvDrQCI5RmgXtZp19XjG+nj/WVdagV0euB2xZfyHO9h6qSjIQ3OjZyTNzJ3lYATH
CBv/7hD8ARoskmCZ15wwv6roykQw8mJE5XvvOOyLP6rP2Ssf5I9PCW/RgrmwptPZXISPD7SLgGV1
ztDUSlmRg11RiZg/RTYd8AVUXDE43xTNECuWGyioy+bHcUnIx+itjbBBHB+eO8pyvIxNq4iIg3yA
CDqwRblZbB8VgcEXDdAfNUHAZeZyb2eozPhH7QzrPZZXW9fH8G/U62cccO0JtKlGwjDJo6U8kLYL
dr98TfuyFO3xVZqCjTLI8CmDp3UtRd5v5+25eUPjBJl/or+slWPhDneqrDkp76OY3GIgN3L+bGJU
wMmk7PnFaDMq0z9LUx4iHlTasZEwqolQM4n1rwyhfE77HufVOyv0uPZwE7ABLp9hvVny3Glsy9vA
oN/dx3jV3Ay2K9lKVF6C6xPQwmaeR1Ok+5yGF1/r3jI0oJFWhJw8nexZ35PKLwYJx+Qy/lSWKR4c
AKhMGNEEAmpHC4hIOC5KgWJlo3mnNKs1QW5fO6zriq/Tzx+f2oaSAr/d/uOEZD+WWSa/0vhOg/pG
DZBsK/VrMRAeebpTVt4r5j8wa5wJEQHtYhHQUKnvO1eX8L6mvIiUdwNwsVlWjN/+T7hRNN7szASQ
PSRYEgqnMWuaVChBsQDrjWPRDSmTQjM5qRT36mJpP5EMnDpgn0t4sVJuNIFFFrNUjs1vEdq3cv22
RJpcQ7InV1xBMJHVoXJ7J1D0C/rxWKh9XVJjtlDEokoTTb+ZoyNTzcqScFtlUQcJyteKyUg/eQT3
zUkC0xLiU5rnLQgcFiAJMt9bzLBIMS87C697gxRyOPpad33I34G4ssu0Htl/OI09ND+cAZJcTGQg
AHVGokmtTa7HE86ZAgetd5ozS7oUKW2LE9m7ON71wax6UkCoeMDQJlng1Sec0yWEDsAqCwtrp5EB
jLJehd0IV8zvv1XRkDknT0Q47jto8guqUDunzXeC3xhdKUEcoSYMHSwFfxBORamdk8DAcpj3vA0V
5r2bWIXecr99BXZH+yJ18rajvZbUMaprdu0uwrf3e5mWHpwscYFPodJvIw==
`protect end_protected

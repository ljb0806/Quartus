-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1DFfSQ+ajh/nWqX34hQuLlUwswHpoue8TEG4usFXHvniEPmYl3y9O7PAeC6B+owKeO3QLmQcviBI
Fnhfl6exsWH7mvgrD2GCJBKsEEIrkA5t2Yjd1jAwPxg9ZiYXGj1lnE5RbbpN3mEkIdHLuU/i+aWE
vQJEhzVnRUpBj+K9IEANbGU35fFpJ2UpMgCjnVFG5gSlZzVFFrhek9MaLoPDYsk4ynPwnMPG+ABo
Dy5DD90KLnn0VB7oLbS+TObM2s4Bp1vk+UMRd7XOt1cDSOrBLT7hJXyUL96/uLGMteb4JfDniVfM
VPX6R4q10MaA/j4KGf5vOgqYq56eIJRY8vvbng==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
7EydbeqSmcdfd0pDqA9s5UUSweXNyH7y7j05s76SJNWN4WNWLXT69AssUmkXJrSH7mJNWsPpi+P3
AImymhW6N8kyt53adzYd57iw6grvjbCfgAawHduQylYMz0tcZevC5o85gHoFx5DhOU9k4vc3WLPt
dyB3o3wtR9fukk9TBD8pY71ZQFD6x1z7ibiHsmdk7qO0r/ms28ClEQxtuE8/QjLTZxpu5Trx8NAK
q0Xx+8Vlp5IwZAtdbbHybPu8d/qxkk7lB6yPvEMRMqO/svW3u1wiJ64eBq0WwRGKLFjwXeSHFaXI
meDpqHBqpOIEGYGjRHVowVTqlLpE/2YyAkaJfiSaWDVALsnRATXlsc6tGwdxViEyenVTDuhCQVve
+SD9MeGHLswP1NepzccxoOa/p8yZt5JTyDUR8NLzAH0S0hgJPQqDzgbtBfNAltDMxcQoHL4+HTNT
RLahPT7jehqwnNGobZZ2OT1tOuzXADA4czxeU2MuLXKUl8GqCKYyBLjo9NoOZEAuGd2bLwaJur62
d9jAxpvFmXuAJvr2vQrDkUFH05M/OOl+DIn1ROrwJKToCRYAeTw0r8sxWaIMz7XUVyQ1zfIBX7FL
6iUkgYWE+7lgO5Y/+ZlrIoiDVc62TZhOxK9Cw1B5wT9sDLbpHEnunhlM0lHHfgIuMgwAY2zUaF0g
7hUnR63sEI5PC3871VAS5sSsZlbGDdwMQk0Y/UsPzLI2CQb11/5SV/BIFJNEDKcajYARCaeVY2b/
aP3Plk+yAGpm+GBT9ZRFJULrj9Gz7bOrRvHvyF0zPG7udsR48YHOSDoUbDJQwFTaMDvg7jj7Sxeu
1YwbMq6ZXbfrckfY+su0eqtaSWetJtOeB6wtPBVfoZmmneaYRMc0fbMj10f1WTDOCADcFU3RzZTm
n7ubxb8ejk4pMIfHuYay4fjMJBGV2HeYEpKN5kpkpygUO88/YMQVaq6+skwxM4/szHVdnnxzXhAh
lOyI1QcI0yunzvgZZALV9Iczqa+VgkRy04sD3rExqY18gGdheWPzlBTmJFz1qYGYvejp9JSrgn8P
icfVKZdbZNz9+VrpbS4qatk53wGP9QaYieIXijnvW1njbpHxijQtff7D8Wu5bhx1Gdo9ZaorXiM4
hu/1IYfpoTybIeT3Ky8vEdfyxAvjFFfy76C6DqFF4rzcebnRiL5waMovsw7wi0+y+wAruLH4vH9s
xq/aejHunirf2aDY6VIydZLCKhxFcJTfe1DJBAfoEM+iK9JD7CY6jZp4wWqN0I+riEyH+J08Yqi7
s6Az9Y4Jr0qhK/20JdGKUboaGaxEYXOBXtONnVVNPReB8XNvpfrQm+L3m+OM3BBZYCIxrDLmS50c
VpnA2LAQHD4IHlujprtJ7YKCw+SdpGuEKl9jn7Bq4FQs9Kk0GjwkNbWTzrixbxsQZVsrCdNm/v+/
IwaRdr/qoVYnoC1kVyuGA/X/KPZnvuDjzik6lCWRgpJdRVpFE1wx/zPnmKtkFlZcKgPhmtwNm4e/
h03ASFi2RRH9CO+a4zn9MDV3vSwXKV2cOmRl6AaYVTE77L1BOTLzM6HdKLo8/jmgDqYgiErZEtGA
uJIiQe9aC3UWWj+kEu1RKrn4qnjLC/dwA3TU+Ul8B5AcrQu5/X9/yUQz2VpjT79MjP01x7rcw0R6
R3PrmtgQS1lUXgwRMS253lTl4rpwdzQdAy/U7OhcNNl26DMpXmWtVYHbvpzVoqTrtognWsxrf1Zp
Q4PAzTEBxo3VEogcNSzrGqOfKbnd64AK/H2UTCGUJtWNhgCkuxbGThneXU2Estexpn/ASlHMe9u6
hWSp01Y2tA6HScIsKWaaSkbSIGG5XUDndHfGPXBpKm5Mfsm+lubzxagEFRHKTsrSNoq0+o9I8v21
Jn4RDexCH1StNDSFZAy6HAiS4qAukljEoXIpd6yC+ovJzgAsHUV2vsp9H9sLFFeUYZNnLe/1W+Pn
vpGpSIz27gIro+awZ7v3TaETiOI4UgEIiwLKO64BMuIqD7liROvdM8LokoCjOOPrW+KTLFe1Xh58
UabUAapxLqKGC1hOA6Y3tyrAaxnIi2ckMQdRhhFujPEv/e9ovDf8JoEVC4RvEeb6s/yPOwpr9KHd
Lgf0wHdHx07FaG2t+j4y4TzaxiKBtrIWJN2DeOTqtQHzfwgP1Zt24aTSqBBg5nqlvf0eWUxa8HW5
VVbDM+R/Nd9vJ8Oxfc0v/WpWXVe4xdoOv0JmfW2SkcZPAfbhPA1NFsBZNKcTC5GepWv0V+ebZFjC
EnVLw0Zt9pE7+B9zyBjqqHPMoNHdtYYBe/r6AKdGLPnpX6Eq4QAwVcOg10hMCq3MBvu/2Uf6sFjX
jLqpAvxwwQfExJnxsZBYwZUJWs8tgSRtmgHr3p6JlrKx/p38amTV57Ho3rhcMkhI5FLPlZOuA5hr
YRvK5EUjt+cPx4coAOiCR6uSBbhObdzBfTVDn/xK1JrVj8lgSVKYOaL+8RqxVbaF+YLQOEtTRA50
SXEkRaw1w8BOfuKO0rctKcuRlju0Xge1OP4m4h+Z7SSrZ9ZMWKpMihoA8nR6lEmBgcyUCkuT0bB8
bnx3TrUcK/w/R/h9cZVvNyjuzgWQ3E0ODqU2NMIqZjTsQ5E0fZWesO8xEy5Rm9u80jjkmLL3xUrp
Sb+GgzQ8esWhFAi5lNozWqOmK5GfxXXMm9GXxa7LLiLkMgxvo+ZXzfrL6xrNwTW/8Nn9wYkEHE8v
hwCulh5+MV2F+GRRF59bIANEkVQ7Txb5ZItkR1v40JhINyZ3bNDpJS/Exoq/UuJqKnsAZAlz2T8t
CVm0BhE7oBkhibETvXvL7azYptdLDOIlorg3x4YanLUjEdr8HYycPKeFJgir3LlWD6VFP8bklE1o
O+O5SJMrpo2gPHVJkC9TSq7qDu+4E+Sm/Er+e5jJrAhF/nk2vMcuP/xcPM40BJewIk/sUVGa4Xhm
YP/Ud2XTnR4wVfseS6eoWt5cDHYUHjweO86OgVV1mKdgN8C/JTmqejiqmHwHaqgX7sLV0Jvti+FM
Cu4BxEJnX7H8I0hN4ce40DVb8W6eQZ+crwKT156KoFmmR8gpHmTQVVArdgfDirWYgJf3Urocr4kS
Q2w7+MQB7xPYE1WyVvxDBj64hfDI0Vv0oHYOs3d3AQHPq8hA7OrkTcBCohvYWFnxjOvywGvBpTvn
m/PJtdP5elSPTEVxPkzLfIebzFh387p4J0MASJTGDNLzNmDGjSLmo/gi1e+X33inXZKLSjS7xXsB
tUUws4ZEoVIpalJVQC9Gh1FWBx7tXoxMz+UYMRpF7YV1R6W3tsWLrx4oRTwETwH+c+SDuFwk2fmA
n92Ra6RduGK6SWKZMVpttc8YCD2238wSyVWN90pxNrL8wWUL7aM1mGjP2wEWuJ1+x90m3resU+Hx
A/sW2vcN/7xvMTaxw6EaaxvDtlUim0x8pkHm0UfZe9MXsjmAyzZPrfJINNI2MqpQE0ObxYz8tRHz
HXTbnFuTqAh6ruamZTAZeXjXD514SBcx0JJEV1qp7DE3MYGg0pTR5kbpN4rIM8opEn82+TpjlNDN
wSRPkLTqAvOCDTripb04QpTAJLr3ZJWL21xOTMDOw8fNlFdLGUwMcCcUBiajJtI4KcRp709+l2JJ
6Zcnl3uhEPDrQL3mwMeQNVCREt8blQv66WTtc8j0odRMkFs+I3Tgk7tyWEYwBUmKSEI77bx8Udk5
idfOXzZz/YnUJh/1uG8eSS1Dhq/JcmOvzjZvL6J9c+F9UGoiq8SdOYtHxh5hHnCorEFVRgT80X0u
tN7B8OpWq8jF+NcfGiv7fvVO1VC+L62KJ9TS2z4hSXWwC5RHW8pAYmeywdzfSGc9bf/uQIuXXJ1i
2wUJZNutfPbWGtDraIGkX75zscTeyrotgqi2eSJ35SuUhqW0BctxvhZEmeNZBvoN53NrNH9pO1jV
tDx/Bs4yifdMlYDCHzeafRLYs96T9SDzYzyURwctdmEiY9No2Odjf069xPos0qEkD1LjI9MlUux7
7FAalKSVg6aSdjm2txfRgZxWZ9cef5g6KPOxQYm1Yfkp4cIdWQE9hp4jeVYe0r26wN+y+U1DKA+b
0wRrC4xOCyCwrvpHljsidTnL1MXRQR3o34FrvWkPPuN6OPwVnbFV6Yv81WkR2o7bYGl6GvzHAiKX
9KW+zc/DQsjIGABbRVQanFUpmwEknpWifwxMBa19novzrgkRp44i4EuKMpyDDB6vQiVMFQAlkV4A
qQDAlNTm1kGgDNZHt2+heFmnloMhVhSrRvrppHwus70mqXbf3ezngFRfv5sLiCPtV++Kguodjd+C
BWDxFechFJWWd8nWqPlaBBtS5n+voNE8+40IzH/sjp/Qq5T6UvdxnK7xuCKbLreHnUfQJKmyufn2
TW3H88Q4RYCmNGE/Ichp2XANO+V3oJnBT9N55ag5n7Lb8drO04A1WL9C/d8VIrTbPeLVxLXQ8NUo
LteafNY2LgOGl71IT5/2lnQ8C8DRvxlNBoE4ekZn4ReHzWQI37zQE4Ydv9BlcxWSZOZjlg34TxS5
ptuztNlMHf2Lj90bb8FUwK51QhPEczSST7AVVapfj6SkNhoYWlboajSEk0jp4iiqB6oH78l5oC+I
GkCopNhPOQMeyRwXlflv9lQb/QpihWzAOEDTQM1sF7cny8uPJ6jcbpaeyd2xoDOCb46i4RybGYXc
efY6COVobQ153okqugE2RYb95D1BY4gCPjlxTqTMRyKGvFkVeStM3Soce8e8+0xr1ZI0jzHHbPBo
dtDykLEQwQiwhfeerL8e8O0RQG8ij06RLMXcIfBmWGBadd4bz63CxWYMQW5lcZUBfN6eyoFgekeO
LtpwPV2W7inYeh9LSWomL973/Cobg6rzjWU3hqwEW7NvKnChXz3w47JH03/ANni5TybpUCFc2T3t
e6clAKMmxX+bW8leoBNDna66msrPyvvMOZNFwebXPopwnXJ+U/c+qixLv5lxOg97sbMWRJZ2vCTo
DT5fSRa+z9hfDSx+kxaMbS0F5VlcWp/JTeVXpUXrasD+2m2U1cANaLmKj3Ral48eOc9oTbNsdwBD
T3njABfG7kNhtQhP1i4oSZgsq2HsD99n/dKvLGw3GiANxujrafb+JnWxNTZqJEWhD0qBde0yGGDM
ktTp9woPNYIwcMJiXqd7Q6MziJiV8htqZ1cWsZFWMJc7isXGtF24iUJ+eEr+A0V535CVKlmCVk5v
6DxKH650ajpE55BOziK39tclQ40gDL9VTQzr3vxzHEW4NN9x4I+QiOalNJ/LP4BQSKNXMaDOzdD2
8nj9C2si5HLf0YxgyU0TfrI9rpvAr2sMJP7vri+vlb09SwPoAXk38nA/XTiBqzRf1SRgJdS4z3TO
2MW6HvHkY6TY9LgBLUzdo4GgPtr4A00t97696yQblN1wsaiPFbbykakiZ3tVdkzF0vhFI5y8PpRP
0SIDrSAqfjeLRnXUpqwIyXhkzTtIiiFABcJ6hPu9SkAkQ+IG6Wm2Z3fQ57wrJkgSoDLK+GERt+g3
h2nq3fOfj6cXC5WyIqMROxgd8edTSLAUWvtyrU3cFXWQVqMKrHwSQha34s8AKTYubsuURnjksJd9
ibAHMLUfTV+NQYb7qaFjgSVUE9UBFfibSDMZrlimsDEyGazJVwYWUKsxGiiaUW55mhrM2DeycM8r
Fqq4PI2ry46aiABNfEBR+EQ/QlsOnYKsNJfiyikfzFX87Y+WAXP8KEv+Cy7AG8Btt3V3OTFlV+X1
t7KOGFc77W0TgQ0HgzCA6RMicg6uSmIto+22fVI2rEU3bQaxzjnMsunibRxxYskUCZTg9pxkh49t
kImqxDzYPOGdQY4cbUtGULi+18uJZpk0fnq/YWxPuOD/6Ixdv/Qnqg9Lf1yXnG+RBT/T5Ojby6xz
c2oqWN3v+ZZzFVjxXGV1WvW/uD7Fh9NhGM14k0iOVvbYzUfm8RrjhoTPZ903PxSSJbCz8XEXTiCP
VHQCBbK/oJw0XRoYWjy3Y3OCE8e1nNzFrQVd8RHcSe9vRHOFUdGmNYJwDPjIWdJTXtA2nnFyf0Hi
Snq48JPcnh7GN+fdhNrXXQ5A+BfkFaZz2tHLvVtCMe6OkGFSnlsXPTWvgLfvVyx4gGzzncSTXYAY
8jE3ZsLRggAc/St/JPDWAhHd/llbCbPBEpkPYr8riBwXrLYftnDrljuH48qKMhGiyMQOmaCQ7vsz
jGacyzfVWqbUymCLm9VAwtPSt2vM6k3pUwWTQCPXI7oqpW4oACDnZaFCeVxh/wtjdcVEUjdKrBJr
msktlosh9lXwyssaqRxkehgDrIzn1tYjoGBGrR9rb7VRY6iJYH3DQuSFU8Z9R1IDCpxOIGPI9hw+
8bgw5yz+lM88j3iGoAhwC7uHQZjg66/oCazMXVEXA387WIF1iFwvzEO8CDftfnouh1Us7bfsMdZx
2fwI8K3sKqH7fso7ZGzIh9ON29NW/qQrtyC9bQUD3dUG2/d5H6/yak0gw19VmpREJi2qgmhoLaTw
PjpR4PuGxjM4+VTUjfEiHJjBG8/dOKr3agojPpGBXhW1RX7ixNBjf9zY+VW1MSLc/fcbUC/FkwV9
dUZhVFInyuvyF1kkf6GlqRg6jN3kXaW/MgAV2qfTsVLTc7dlrw/U45Meifde/SM6UD5Xe51PzrWV
qyUeTjkStNDnqrccoqrqbN3RNHrlgQFzJgDgowxhPhGlqWNw8oX5y3+rUEn7rTCHDP3bmzd4IxLE
K//WPIgp5i85ZXgazBvyG3VzzentaS+DyGMK7ah1ZflgHoaKhqzFDC2WkejePg4kHhSgdlLduTj+
kBBnqz34LS6W0AZNdpn1LKDUWPM5+ErIipgxa8yLgMY2jXD4X7yqs7QPNkmvccwn1aBMfNjrRx3s
D0YYFuCclrehdnpu8CIvwPlWYNdlL2L5Y1uWQQ+gbVU55BySZPFVYidL62WXUKB0oBf+LOn8s5hP
eBWf+bhuPegxNaE+vVQHzuvD3yWFbHaZFJdzGHzVXLSM27c+0rKT8uoG7X25ThagOGRPrGv23xaN
DHE003TYgTVhyExMfeNbb7xep7Cx+ByuoeMzGFXOigAafzjKCuIFiNVrl0Nye3m3zBHx655PqRe1
jUjj4ZT9WA8n9wCbs0VGx9d4mgcbEl2WhEt+Fr0jzbT+Qp6nio/ajVU7/1wtV9kdf/3EfR294Wb6
1ZMWoQzC3T6dVOvb5bfguNsvDoxDE96Bo51xI0aKxEBtAmY9zobvnCLypKlkXaIT3q+KkYHilAu2
/3CC1sEWiuYN4xff39lZ6hc4tTCLwWMIfpFgRpED2qeiiv316n8txwK4nU/Wfa9ICQWJxbrL4JaH
CCQJrxh3koo/0KVazRBsPF6/FFIPnKmJih/5zNSmXgqeXbiCkavMHQ5zwzShJRRwtxJu3roEBV9i
uUZpSm83VWR3CroR4lcNmS47jr5hsah+bbET3XD7mIHMn7JjAyEMceRxshEM0LG+l2gsjQKPHoDF
raF30ktLsViwGewKxr3gRpLQtpFoICJVcOy+xJR7kyz74eE1HRNYTJCCm/KDQdawwHKv7msI5ZaY
6ySjokA8UiZEwaBAMCjDPssuppjxScQ2QHeK8JxDG1AOvL43aKgvLr9HT+bz6rO6hcx3ulzzCIWf
tgtZ3mlEA3YsiprTZ0nanMptFmNJSkpyGXKoM4y0Y4lOBAQbMAvxW+RTYSXwzORxCUOuQQncM9rz
eFdS+4KIqJlE2Lg+Fw9aK4fEOCWnHmJkTqFXwUarq95oyjJEdgo3FqMvc74iSRI4KRjtlNfv05Hn
1yQ16NqLIXx7YITXiRke5WZutI0FJZIm9cZdItPsmaE1E7uclKUGheTuvYFMnPcGE2+TS3/MvK4h
fFcGo/+drOnipA93HeQxtIqusj8qS4ZN6VWzMKYmbbMlgyRKM65vJxfOxY0s1+dS/kW4WdDIdFj1
qjckZ8Sno3+swxO98nW5ObdOoy5AVI+VD9aHCeeiBJygtRSf+0yBbL4JfLUw1DEHn/Wgn7R/3QA0
I6BGqzTAYHlfSPf6vKfa3+hS2M4MaRmwMdo8VCLOWql+EsEmIxTPxnzVek2ISgxCdbvdJA/c1aDo
RDY1vmV9TGwoF6q9JlND0jknLZGX37o2u78NbY/C+2DzbHIGBAXT0ieYEBLnncsAX9UoFFuhn0U8
FlvVZOn/A8Y1pPOnbWDSPBS3neerDr9MZq0uzKGGxmYFe6+mbSgLd4MgjA/AtuXPGGIDgz8wfwX5
H55KWbPdNr0fvgzKGS7HCG6Glu1vLU+hDLz3H1S6DXt9pu5n6fp4QEgiGhMDCdR2Ipkkz/ORAmlQ
ETo3bUGrug/jCScYo/P3MmFQxUuiWMyNFWzd6uXER+h5W6uoE/6yZodpif5XUXoswGu+WpgxtCYh
tRy/H0vkJ0lwo/T/JiiGfenLkXTqGhwchzCFMRJA8DyMbLzz/VfG+2eKiNqhcO6KcpRrkGsfZl7I
ZQaRwGyg2Xzaa+1+9KChWXTgZLlZVnT0P0KZ9FUodWnFI7Qx3mZgzJ+BV5aGHYNm2bgAI8ItKo/A
laXAxFjhfybMfYs/mOkPxxgR3Mdacrhr8G+1gZjSSvoFBZst1YoZhe5/Cn8WobgQyoSvlBErcSMW
7NS5nFqEBPU75cCXDKxgkUPJh0ZrVApBkJEIazsNwdPRtUc61TbUpAdFPaypmOTSptmvL5c17rjc
mckYYGYVSf+h48d5KRtcP3Bwhac8EuubFqc9GJgb27zgqT6oySLJr0d9zIhry7m2GVA6HPLSm6zs
PYMpDiCw/CvlCg6KxvDSPu3Qwu4X/Pq8wTOijxyntICyS6c28OJkkHzs+zw7TymOZm/D/Hri5Quw
0q+WnJBJhSpW7vJHk4w3qpiYgfnOsuOkWGgB+X2uNWGLIF6gCuTj7KqNKgX6Cko3D+un4Aw1xA2p
iUdy5ci/wORNIxOU9RQ2FzaKvjWY+ERlRiUSVJMreHJGoNqBmyQy30h4xYLmIGduDlCG5/CN0p9c
1E2/l2ikRFM1emUMa+ppHtOnIHxpLWwFYc89/tTle1B04xpxS9ElDJXloSwHrfHKG3bKK9tmyLtM
y5vy6vhyaaO4zcVTqugMv5KS8Y8/W74/552NwsD1nN3r9NW1ziYhM/b9t50SJyiWEjlPHuWbf7yj
V7TVa5CjK6IPpIVVMZuN/b4NBLCnk0tLaff4Gm466Xit6xFsyJviyYfPcT4teCGiA/46E4i7/IfE
zFXaNpr3Y72gUFXH096un9fKTAz5ysUPvpWGBPqtjV6eQxguuwrZpvGL1FPfwCLZDXGGv46Im+Ti
0YQAATgZai7GmyY49mBcPh0SGg0aMz3gHHF+tpP1/pd4jJpzrmpIPVQ1nV8hg3UahREK0RFnjPAW
P0sVph0UndBzp+bwj7mOg9udgRxMmrDMBja6RNite5B1lAPB2BRvHXlgbll7iZ26SDClsb8Uab3k
+6lK1newR2ILbHm1RbgMnT5W3YFO+mJxDBYaKR9zhXkzsjymoFSi6WvOED/Nm44PVJOSKVvn8xbG
GbCVoLWKs83+jEqk0N47InsQ3K3lsq1GY+m4k9xc1iv1VsOhBYULciGpq6SO7QCrB8pC9O3K9sNw
2DcoMyMHpvVBRm8wh2AiliDLx5UaGUt1oSOz8QJkIu/ulz0+a1v5maJ8xCBrazmZfnaKnA1jLSK4
dwtmNGF/GQZgdXvbkcYuxuIddRITMDIvf3XOxqDUVA9UnkIo+fc++qwu8h0SIA4T9Cmfjoe9I25F
GlzqsLfXZjsPY4HtU6pUz7hCf/pqeskhN6fFTHN/xJpVSRt7JeRGkPN/VkFag9yvuvh/XUVAWH2A
Xxcf6RG4tgmIowAyESa2myKA20R35nOAIECx+URxCWz3cRhcLzHqFqgrvNLfb0oYO4x2kXQUtnnv
8BxoOS9PnrBfZq95NuG4cZyVlSX7NABJXHirkzpcJTsou47Ruk4CgUlO1HvX6wkf6780ZrYWzP1o
g9qry4h67V9ZeiM70GixAbZDHMxvZQdQf8z9qz77xh787MRCh7JSryPr7SuP95LUL/IG+SLwsGsJ
cuL7Huibd7Z7droNNgqd78gixfsm9enTjvn1PQq6JB+mIOT+At2pstQOQEfILQHn4vX7A4WUI8Go
ZQnqctpwbV7jbO+tUxMP1iAknpUsnfaJF/vgvyjlduWsXvb2FaZN86g/aC3Am3a7j0bMgPriITBJ
BhdqClpkCa2u1DHpyI0qsijBBBopPGVkXmTmnoOJpHam8KmmYAsAjZ5E14oYNBak8Y5XGgOY2zYN
5DgNImiJpl29zmCa9a/JqUbECXVoC/Pr3iQIy0agWH+UABJvYpABbA/w5qNnAqDUJdnKIoOsV29E
dGBCRG1dWrXiQtiJd2wtp/hVN9uQUCDdlRY3k6GheFtLf49YWiYqLtwjWIxndbZ5sMXidWgVucMV
jPcQ5lCzO2Us4VlabskJyyh1giGYQ9uCk6byME513d5u6KUmzbeRRrcU5+MyXwyJ7Uf6zTrmuPSq
qyed4tP/R7mneqap2oMlcfIDzn2zNguyEXK45MqPltIh1rFI6/q3OgZxdB7bnemKhPR/ryE7+4vH
ClZF6AQsWQRSHk7WpnyOSFSMKoD1p6HGGqAobUk6n8I5iRAvbvJXIj6fNRqMKP8p4h00iqmA2LDt
SanQUnVA+9gE9Vq+aNTDc0vgceYjkI1cNw9MUGhWNKH3zDq53W01tpBLHuip0PThUIgNyXjdUIlU
Sy48/KBHLY090SCXwPtqB+oM/zeyiu4DrnvC2mo/lbcSWi2gqUTbiCL/ICt6som1UEP6pPdMdtO9
CMBDvSaOJzrsg9oAdVnHMaUscI4HGCbNualMoPD0a8bQSjVKa7v+0t7ukl17YYHuEBOWgOP8+bjn
2JSSnl6TcowVfpYPnUqgXvoFGAp3GU72PFv8OtzuUzH96bbGs+AIaS8/29Q+JoZDT9bAFl8awLxw
NfUSs9y89ca9KJSELrLv25FdG8jUvn9Z4qB0uT6sKjZZcr8t15lEBosYgC2RS6ErM+F8Uh2A4tMp
7ZxKkLOONgMavdL+7BquFw3bt/oRtchBg0DTvV4sbGtKtWPOs2yf8gtnrxdPJAavFrVJBEhB7ZEF
Ym3cIRlzODFxKQZvic0jEI1khgdeEjpyTZjOJDz8VRQ3iDF6Za5Kni9Ir8DeBeSsINhDCKZ7QZms
kXLubbnt0AEDencX9V1D/aSN/N676NXdtIM9cPlB0O69mo5F1SuUVyr7k4mXX8eLO2Kc5a1s3f7y
XGFoOdQVIKFNkCO9gXGEEDutOBlvnJJSRjBStVQ0gVdhzUTx1LyOuFgmxYBSnk/w8tNR+Anjis7y
5/HkJV8C8NnoKLZ5b3sLEBDPOdqXzChmDuwpWMuBewKTV6zXrEO09JldvqMLmroVBPNZXJL/Nun8
rIz6pZqkQHuyv7gc8zuXh6e2/UsJnD6NlUEudZhuf65L1p/aZhM5tR6s8C00m2nna9gx2JMwYX11
iAdPMOxmVAoEgSr4ro32hR+GXJv+OxTLxcaNaacoiuHZpEH30SbgrqcOkz6USYueikFg0lmyZGlG
2onezIEQwiU2Ho7UAXODjBB0tS/eh+wDib2Z07/iX8QDyCjVfOvSGtN9Cc/YQoMQ1THQSsCk+tmr
+KinNhQWwOfL8ktwd+pIkXAsTHbsLPKXIG8bDMDLcUoFFDUTjiSUQiLo/0o5NphUGN8PXms3OeFR
+qG+/gvvu4WNd6E+ddYhE/dlj+F87oTGTpReMGA9vq9jS9OQ2eC9xl3xuTK/DbQvCN0e45fRWBuC
6AzJ721NHkkYWa+QfSHa5CA5ATsi0xRT1nUrQcADePGBcSH9QB0+/SOHorVB1CpWfbBBcRSU3hhe
80foi84NZ8t/YavP9L44VfuWVIRxRNMH8pBxu9A5gMZAQE6ZQhCbmEAeUcwXJdykfztpFgz/jV30
R2QX1DhN4UqNM/M2qLUqKC4ST6xSmuP3uQDMibiKh0Zq3aT/NR61SnY15qQl94XReytc2n8Ow4xP
pHfqSouvAOUW/APGCiZutqhnVkShw/msEPl2lt6TRaVTP7TMxF+nEJVcUeAff8yE1IZa9NpW77qa
l4pSH1uWw15CZyAhfkVqLadxDV9TBS5Ck6841JMRsgJnGllatNpQdD/Q9L4XrNVU12KnaYL4Jr8s
c5xAUX3SLNV7MXCO5LkuBFEJCsW4kZ3p49OXXSoOjO9QWfaf+h5c6/AdHRqoE91Ro8GIi/ulHoyS
c+PHO+dEYOgHvS5BSZcUDPZ6HjUTJIxge3p1ec/tyDC4FDSyaTg293F4nvrgrqLlisXx2fUZYnp0
a8FeOoe/QKE3yZmjko/neScRSB2YKZii9O0PvRii0ZGJQMy0GGw7x2z08sc4+lHj4MDHzcUk/w+t
ucSyyXYly39b6PNjXfskzOOQinDqADLiTLyhUkG96kjYq7QE57M4jfejKTLe0jXvR0sUZm+VFLc5
cVLS8xYVzHRRTfXPvZ/TeLqWkolYeMedi1McvT3iAo/Zf0RT/23bl8/uADp2SLctPNV0w/8molMI
y5mj7aoGOfD9O3QH3Tm6Av4r36J+jJo9SUi3Lc2dM1uW298smO04ZvvdS3wuHlDuBas7f9Wt9i21
gAxmB3YUdTw6aGAUXK1Po2M02YjShMInxEkFphkNxwy2K+dIr/JWhLynpf+j2KTmITpCcZilvzNa
K+90vog/qtssWKBX91XD8i3nhr8co9h3SBP3KW2/7qiqDo0ReS7bQfiqytGiE6axvZghfTY2+NEA
GGMyT2qzFB1WT5KlbQxDYRfnp+0miOW09zeOrNrPxOG+yTliLH7G8xQNCqTLR7tYfzf2c9N0pUgk
kM4w4v2Nz3h5RjtNQwLqoBDJfBMIw0jfs6HmFRAerv8qY3+b3QL2xKIFZGBRUFKQ6uFrv66SE5Jy
hohZoiydjv2bixPFUWajhtFLmhIBhvx2H6Q4+NCV+mIaEUQoCqmaNdIqnNpWqmq6mmx9Irt1qcxd
jYNgxpJ5efNBmav6hzuA3UTurNNYjXwrkdohPafyolnmf0aGqwA+ZP6G6GVKdLoazOk/pfYAVXue
qi7eGLBHyf1n3kAOEpEhERsM6uo+6rHEauYIhRtRUPjSN50CmAdqGsrQ3BErdeeMYMf+i/hk3D4B
rI8o4fVk8xEXUNl5UigsQzeVlBQl6nRrvKKfunkej0gdEKBd66WYI+TwZ5AEJhqSDt5zpKAkN2x9
BYbNE0OxtD5fNAVYvwtPnVHLCqNGjMeVwrarK7twajQ1PhK9ijdRS/SRKvOyvcDMdICT8uYQn9fn
CxDqxjKrtC8rSns7tWCGkKlxMBYRZ5e6fBX+kjATY/9c4gdMOoneXOjI/bbIwtEJAlps7Gu94npr
z6yHYhnIBbBILT0EEm0dRETYIRcjDu03bymT89Y6IpLXfZz7Vdxs46BaoKEg5VKwk457097u9mvJ
Jlw2ACgRyNG7X4wj9BCXhvFDaXXGw+qHzskyB3LXL8smg/fZFA/7aGkCu+jI4QkUsO4shQEqzk/M
zaSqVWaIFSliQQB4p6o39FCQIgkIOss8MBAYUQ9VU5EK9R7jw7pPp/inAEL2+JNUnlJ4IdD/ItUu
dvzuAeecSDTUcnmLY/f7K3LRa69HE0kZrCR0a8h6dwbOjHrRs9s5o096Kvx8aybA2AZYl6Bk5QpK
hk7QsZeCrmiZ3NuCcGK2LbHA8NVnaVSZ3JsCE3fLho1iSY/E3SKjdIa1CrTWUEg9gPKpbkt0Zx3v
xW+lsLq97CuZafWVbGI1AywMnwSPfGfzT8zCXrnoQvUNJckWW6b4M0aTHSuddCPF5HYIH+kUWodh
OaNTK/MZimhaKT/lrxdn0WqStb3mUfzmImlFWWewd3T4hwvGhMD3wzuc0D+n+zFMh4cI+EWOa9Ll
U5Ulc2s2nu6tIYthdYe5EiWaUkTrKucWGnnlPtLzlKwxFB0+AARADhIQpJs/PnA622Z3an0PbU5/
aN9PJuoUJlS55D937irGZLk5PMR6e3qcM+gb0CY588b5oMOdtCvJ+GQAD4mJJ+E=
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��Y�H�EB�Fo��M#�_����`; �1�����-:Ć!%n2��"����]�9!r��@Tg��i�5��F�g���΀``Д��[X�R�4X7�(�=����_eF&fn�gzn�
6wV&����Mqp�-s������G
˰s�@u\>��ۗTi�\mR���N
Wcq_ ��y�T�p2-/��{Mӡ��P��g�yD�Q�B�tWt-����6=V�@[PEk[m1�e�VB����ZΟ�#��*�R5��b,n�_��e_W�=#B��R��D)'��n������z<�
귣
 �R�^y�b�mƮ���P~������w|�0��\����G.�MZ��Ŕs �e�����/��
	_D �	_0nǈ;B��0;6s��.]p�gO���4�6v <��-�qy����Q�z���_h��/|?��{��V��0��	��o'z �bw�L�S#L�ίci�w7�	(��P�K����8'Z
�3qi��Q���PGݵ3��{X�k��ق�C�"� w��G�j�=��7��->'���`,��%��.�`.���^�Q]��<�T�;�X���^�Y����A���\�9VPG\|m���� Mw[�����bު^/3�b��ד~�z{t�ܧ����)K���Y��'�u�zŪ�R�ޭ8.gJCMi��(n��]�p�V���֮T�h�|�zM��C.�nY���-,���Rp��ٴL�X�u�h�$��?|����G6,�{�#W������0-����g��Nhg�7jnR:ß�*��q��S���'��n����oK	�Sn|�0����|������B�e�4 {�H7�e#�M���MW}���"�*nn��v��h?1o�޼�V����N.�MG|�8�o�� #Pn�']C��9S�*Ž߆H��	Q���ܤ�c�*���6�펇��}�����|v�&�_0�K��p����t+�A[>}5�w�[Q� �P�b���е��5�nYW��GR��3ϒ�5z��^��D�����Ԧ��P/��	��ߏ�':���5g/yy��bէ^7j���f[O?����4�:G�{h�qyjU��Zk�yu��c��UT5 �C�(����}GV����9�<�o���}��B��n�� 
��5,3	ɯ��)�H$s��.���s�_��-�U��U��Q��%	j� י��*��!	M\����)��@���5�tJ��6`g�'��萍:{��[h�>\O֨L�5}��F5�ѧS��+5��=�Q�cХ��b��m������52����%0][̉�`JH�{�c�nf�c!%bO`�&<N�O�%Fx���q4���gY�
�;���/Z:���K�z�)G ��+�/r�X���6�hT0G�(����S������}�+e�"S�|a��`Ω�c���)[�u	y��^v�����;��
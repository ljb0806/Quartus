��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`�����T;�x��Zg���)U�b����\C�]ȧ�n�ig���uWg����Gb��i>������o"V�SdsR����r�x�����5�%[x�
�e`J��:������D��%�֯qd�����D}`��н6a�_�	�ͯ�m�B�jpG�zy��b:�1v�cn��H���G�#T���n��-:��L�L�;Ha͆{���{~F���pJNG���&�P�>ҿ7�Hefv��po�ڐ1��R����J�䬝|�-�|���/���'O���l/��Tp�i��7Z��Zx-~�P\`J�{*c]��RȾ����%�T��I����$:y_����_>k��R|�!KXEɁ+��J %��:v���5I��k��뱌qe����j����}ת0_��ŦhK�FzC��Wt��7�-�Pm�!)\U0�4����<f)!@�)��Q�.��{l3#��lF�%��*����E���-�6�||څ�:���� ���[�e�+���.Z��kE���F*��t�A���/�h����(ё=n��=+�y�D�+��q\�HP0h9��Am
[5o:t��/��6��6�Kצ�?�d3�%���/X��|ƌ`�@�zz�R�Y�!h?c��v2F�"ac�U	����\J*:���R(F�� ����X��`���>�͞9�����z��g�:}�q��o�JŁ�$DM�10�c:Y�Ch�gC"����1C���������Q�������\g��1��OՈ!�㏥�"x9^�6�O�c����e�&-:�%�>�z8I����
~
�l38C@��������N����32!�u��$�p8I�S*��E��7.�8u�02[����<�-O8��`>�d~�6�(��2���d�+�S�g�Z�8�8��}���i�M.�%��:��_�����S gK�s|��������8~��&	�>H���ηt�x����4,	A����Z�J\�f�6*�@>9Աi��t�&���s`
W@șE�ʠ��^<�?�c�!�i0o?[��K�u�ZXw�E�]Tp_H����Y�W'�<��n��3ʫ�8��B!vB�I y��N��q�&I^taɁD��������'��h�V�B׬�|�B-=x�37)�ɀ;:��U��Ke�x�CrA�,.��6����|HO���Gs�S2O��|?%`�'�v�^�@�TG^h�����u�偭M��P$�x�`����aC�\Ic��@�N�} "V$���LFcG�!hu� 6lS%��R�%�i��qj9�*�e�{2��� B�O�����R���^��&
��}3�j&�n��L��.�����Sg��A籅W���w"���ő]�x�J�x@	z% �:g)�ߢ~nrU� �t���߁J)��2��[��2��������n(���(��O���9诒$r^:���#,�N#M���[l NވS���_� }���!�;.Y�k�4�Q+���J���ȫ灻)_{3�� \�E1Rh�a:\� D�`�D�ܱ�dZ)	�؞�:{o�`��b��?�e�No\9��k�q���m*B��#��Y�3�� �b��J�k��=�IB;����
���Gz Y'��wY��b�������{�逃"�����WA��#g�Wym2��$�a�y�4���cT�ܕ���C���zS(�	qi��@�f�g����!Z��q�HE��U?O� &��|$�OY�ZD�9������Z3`z��aA���u nb��v�Jb~Y�ls19�3D��t}��"��4�kf�%bъ�WM�^��I��@�J}c�&K��N����4z_�`�r56��f$w���%�j�?M-Z�@
�DFwuН�xq��Ӯ�ؼx��,��/���t���4C�ql!�	�'��6Q,�7���� �'7BZ��]j�g�2d�?�t�����=�V�p�fr��Eތ�J4A�m�5��᠟����I�x_;!��a�w80N�5�E�l�J�h�uL��N�-�����w.og�I2����8�_<J��iU.҅�u�6���/2e��wAiĻ���,C,A���)`L#*�R��|��B*�^]����cv��x������V�r�����c]v�!����\��K(��6��]J��6̔t0����+^q��˦�dQ
_�X'�����Z0R=�,��'���(�����ϻ���^�՘�S�,�ii�;uxz���it��������N.�=�9 ��QB��ܢ9�������P`
[L #!����DE�ܛ'9p_
�&њr��$��ȷ!�/t ;���F�����9�	dL,g��2��Fs����D��ަ��By�q"��ߡ(c���#ދc�=m( ծ��Eg������UfKrO�i֤}AAy���w�r�.��:7��<�� �k�	Ѓ��G�]�ԅT���F�����ܩ�-����"`���6X�7��D�D�/R�[#��Odf�y�	�d�[�M�(��K�����}�
Wp����0U�"���E��&�a�(5�j( bZ`������\W��T8\����w�f�f�&�4~�zL�Wp�@,Jd���&8�ә��7e<Ho[(׺��N�����:M���$�b��2�2
�12���}f@:��?�pX����ر�bUM�9?ĶF&ׁH��͘��pFS�w��X�R���N��Jt\���b��U�����(���Q��j��5�E���X���
$��;�`3��;حX��R�Rx�b����3Xf�?��v�"4P 5�z�ͤ�}V���mRQb�qބ*w�U������,�3�q(���h����>m�ȓ4��'B��2t�^�T�C���|�`k��c\���a| ��eMzJkb'�,��i,�8��~��q4�a#���e5�I��Y�n��Q{��9n�`�_5_����b3 �c���ϴ|ڠ[��g��&.1�ty����c�#m�܄t���+�蒀FUp?�F��
߿}QTQ�*LuQ �Tk6(��*S=���9�'s�lc�Z��o�!�J�0�־�G�'>֏濹�l�Ĵ	��a��X�rV�Bx�Z�:�b:��4�	��N�p�� 'qSDGk��rķqHb5� ����'Qw!?�4K!p�>��vϟ�C .�e��;
��L�"�8#�X\AL���uAS�������q&Z�r�k�L7=��=Q����QZf�X�H
�Q<.o��}��B�q�&1�����d
:U�v� ���efSؾ����H&B8��(�����y�?���e��ǆ����+�m�� %M�6���D]'S���c�>�5Sԉ����9|1�B�o��#ų�c�_�^@��>27�!���Hf.E-��L@��E��b�A�G�Xt����ŵ�s�G�.�"��$(m�c�".���ژ97w*�!����|/�����Z�5�� �e,S��V�K7/��v�؄��aM>NP�z�Am���*n	�e�Q�+6My||r?��R*���,�l�k~4�е�+
�:�����B��o����H�U!��y�Sx����[���I_�dz7~%��#��䥜Q�c�I�*�����	E���E����5Ԫ�{�(���.��j�rn6r���y5	ĩף#���ٗ)#��ch�%�k�T��n��N)�h��$q�_���`5����	�<����G5��y��U:�^$E�k�1�!�FW�/
Q}���"��7u���F><4�ȌVw��Bur�.x�!,�h�L+���@���C/�}m��o�#�9L�G�b Yl#Lan�x���KcE������~�+#끫�ִ�9hÁP�R�1��W�<��U�	d��I74�v<#3�/@-�yr����م��cʷ,�ϸ#m=���,�@�ʑ*� �c�O�����)B�αO>�mN �[����������˄##_l֢?b�B}�E���n�J�pK8�S��J��0�Tw�q��4��!��m]1tm(��!Ŭl����)6��U�������A�A����������Hj����0����𰥒>�o�CDQ�?æk����׷ #�mH-5(�G#�8d�^�T��\���K�\�U8gRc�w7GO��H��	�%P�T Ȗ�T�ק�#WiZ��e�Q!���C����:�R�C��Ф��;U|���vߘ%)_x15�,�����[���M�ɄA�\�&��;�f-�����A�bg��s�ƨ���Q�<�%�h����k]#ٜ�F[y�j�ڧ�4,�#|�/P��@��du�XF����G��HC� S�%�g�^J�g�`o��a	��U��X�� _fj�o�po��&�[�+J7�`��R�'�K�)Y]y>?'/��	U�c����(��Q\�: ��}�'��U�p�\F�nq,��A���������]�:����ߏ�&F��D��C� 7��3~��7��~$�;l�׸jy&y.2�<�Z)^�>�F�-��4�L�2�c��7�l�=T?�D�^�e�q�)p�^�`"93B�dV�iص��V���P���'⿶�%�����2�Œ�)Kxa9z�,oD
�T_�	�k^y��4��ևv,7U[KS��/Ϥ��]������|	������*�ܧ!*��w��6��Me"�U��0�H�����¯u8a�d�m�S��5I�g"@r�C�cżpݔq��?'����R{��T0�*�P�N�[�S���%�v�P�ᯗ7}��v-�b����b�x	�B���'�(vJ�J��+�6�j{�w�Q�L<l�i�O���Pils�φ�6s���v�����AȘ'�&�&�z������ ��^��(�q('w���l�}glc���À�-�x�U=�oO�gB�7��.��	���-K��6�U�K�"�ېED�r{>�	efV�U��j���rT�@y��6)-��Բk����]���M���O�Њ"�x}�a%Hq�6� ��k	4c�M��(��8�漣V�%�a�$��q�tizq\I���Q�x��>.�0��,f��)~n���zBCZ ��L�'3�a�%�s�l�)�|%w՟ ��c��\��g�*!~�by�J�1�{B���ۢ��)K'I�	�P�������#�*�}}�}�V����-Ȋp���ݫچ��?�20�l�{��e6qd��u�E#�6�C���Ѭ��M+o�k��� ��a X����fh�9畗[��|o���X�Bcr��e�"i���	���{��q�J�����*P@*8�����
�4��`�|nhJ�{@,��Q5�Ұ��a'L�"9EN� �W��0k��*�_�=��:v��`&��(z�z+�*řTjaj8����8Y*U���8��?%�7/j-��jL����c~�M&�ڀ��g@My�<�V���_���KS��{�1��SZn{B��$ɉB=([��w6M����ɕ
Q�܊o?��*/ĺJ\d%/p�����]ٔ�d����~���L��{x�'���Eɐ$��� �ꯔ�"��dY� /4L��b�й��j�B�2�e�P�����1�"�7ٓ�I��ixU� ��;9�#��͝^���T�̫�Z'4����C@�Rc�抒�>�ED�.F�ۤ؞��% Hv�nڑ������������n�3 �Ҥ-��1RDq/t/�5R�w��{ߵnX���a�[�r5G�*:�s��i(ݿ_�V�¯�E���c�&/)��׽Gw)QW��F�}	3`G�
�Ś�}g��}R~~�Z~�:a��0��� ��{'�}�������p׾�@2��)q���ZZ:���E6��3�e���Ε�ac��KBx�

,�b�s��AY�v;`S'¤�+;X졠r�L���b2�����z�&�#CE�\�U/���s�P�qB+B�*��Tz���q�>bM���$9���ƞ� 
��t͒��J�a[�8aҚ[w�ڗ�����v�3�:7ւh=[O�����������`�W�������P%a���T�%P�O�0ݫ\V�!�1�u9�䟁�*e�8��s9����-�����g��g\(���+�~[m�Lh��LGl��$�?w725;�?O�{h>t]�;���ӏ�����#/�'v,��1ڻP�~��Mx�\m�enI�ζ��֐����	�*
��vm��p�f�m�=���o,�y�ֈ��5��"�Vr��,����
�L#0�"�����@-���q'����\��2����ַ�7�+H=Ȑ��?�Wo�g^���N����I6�| ���{k�W?��i�u^��uB�u҄�ڡ�5xy��b��S�JP)(R,�5��xB:I^��i&8��)�}�����r">Rdi��9@�2Q¿��Q*����ok_q���ij��MD��i����$��>B������#fx V�s����G�%�j��u��븶Ԡ�|��&}��]jW�E�	�!�^� ��iv�.D�D;5R� ����z�g`�T^��6Vo���6!��s �EϨo�ؔ�^�
�e��I	|�_#J#!���I �7f�H��C��Y	��<�=�n�^f������h�(���
>��k���^��/���_-��TvHm_���KB%�Kk �����c�E̵���ڽYl�#f;�w����wbPLF?���'�Y@�����YJ�m	�Y��,��5�ש��R�7�&��4+�ˍj�ԑ��~�
������V�*�K}Ԕ�AOOc����5�\֖�v�X�/ď�D���"L$׿-2@���Iɿ�Q��P�&�[�U�:IUn������΃gކ�٨ �v+�r1ь=�0�3i�=����Ͱ,t�#����#��?�cB�&�[8�|���6s��%�m�E7�_�ڶ�휿f#�nf^^�?㴺��l��E^*0�2��'|E�W;�����c���{�R
Y�K	���� �S��k9�n2���I,�ҋ�cxU������j�V�a�VR5z��dk�WK�Zͫ�W�Ю��F�M ��2"��fh�yz�wG%�NqdY���;�����q��d���1YK���T����]�%HUP�Mo�yٟa�ge�IllW��i��Za�~��GX��6)��^�|�����=�뗸:0�0�)k�Uk�?�e�:P�jT�w���`�L7%�yAF����N�RM�y���,�yi+o�8�-�L���z+��:c����)sf͜i�O4�UĨɆ�W.S�.��o��_뉼p!X�"��2�δc%9ښC��m�3���}��KW��ֻ�<��EW�A�hfF�N�hO 1�Q�+8�������{��R�|��v^m�Q���^O�E�Q��]�s}2��K����؅�6;���֨�#�g�a#P�JS
aG����
�lP�`k��L����@R�bIe՘M�����_y ����R(�(�����2����oB�4:��K����(F��Z떋����BmD��Lj����6֭���%��/���X��2�^� h�b�._�I��<4������s�"��8k�rwŪ��&��9��su�"�FB\A"�s�\�����&W�>�����Bs���u�r����������
�ݵ���z�~������ 9����T��un=�ݎx|E 2�o�P�s|!��L�vԖT��P��;���� "�37��v��v���CĪn�V�،�Q�'�N�=`�fԂ��C���f�}Z ����ml�x�Jb6�6�єU'Ey��8�����ٖ��P���=rP��ܠ����[|�k~��I�kR@V�e�5�N�f�@��^X�/#�!�e�����
[��l_��-΢���1�
������0���HP�9[������f�<�G(OVS��{�Y(�V�f�v(�ʦ�� ��O��!�_�[���^��|��tZ �U��͐�p+�s��P�(����t��u{ێ#�fcõlM[7�..���	f��)@P��*��	:i)#-N� Յ���YE���bA@Y��;g~
���-$�{ׄŜ��D�m:�Db�TT�P���X��
�2�{'�7#�x�൛Ս�s���5F��Xk)�uO�Џ�.@4`3���T����ǔ�����qi�u���MϔN2���[�X��'頬	/E�����J�i�J������a��3�_�0}7�oD��SE@�D�IyKc9$HS�3ܑàǄ>A>���0e)�.�u�h�!�uD���Ö��^��g�* 2n	�$��b�ȹ���UQ��\�̉ڿ���<7(�����
�})�߾"C��qRP���Or'j5���Նs9��������Hn��@��(�x<�r��,Qa���}�M�\���F:��v���`�4�/O9�H�k��7z�T�пM�8�ԧ�ـ��ӓe����*���(0BDB� ��d�����	l�^�ǜA��Ơ��(���y$ܽ��f�̋�	FN���7R#},�iRA�(l����A��xǺ����`�����l�סh{�+@R�� r֬�^�[S�/����󧧔a�v$���1V%�����i��13��-ii�2��ayV�^e�m����i�I�_�a���տ�k�
��Tt���A��$2[2p�ʽ�z�ŹR��W�(ڮt:,#�`�f���00�����]6Z��0�f2M��*W����Xb2�Y�'z��)�ɍ</�Hb�)�}�M{���J��:�j)��W�,43��I����7�ל�`
�ع7w��cG=�MI�ϭ����Hay�ȇ��8���`{�i� ���9�4L�[a!�)���%h�K�ݿtrcF�v�wb���o$~Q������Ʌ��V�zp��i/+�փ�$	���inë��/�x�X�ϊ�  ��U 5Z���P�N��T����X=mN�����n�o�SL>���k�|��|�P�1P��ɵq�;H7�a��ܐ��l�������a$�&�*�c+��H��";W�X��AC�h(� f1V�#_����>)$\t�&�ŵ��H_:n߄:���TY��_�Z���U�9o���D�2�*�?;�k�_������<ͥU��%����1����6�5�̞�?���=�DF�mz:;B�&��V�h�B�%)/^C�0��<����+���1�c�	�/l]XT�����+�N�`��1,)R�p��mӏ�-��:;lb1��GW�;Y�Xq]�S��3}�dT���Dj�_?���+K-�=ӻ���K���u�og���G�
�֏�KG'�d��0v�[]�����v|����}%�ޕ�m��4	L�"���Ff}�ع�P��#��A�v�~��F�jc�;����X�C�p���r`Z$͋7c����7��gU����B�'����ܔ2]Sֹv�	jˆ�)��:'b��cU�ǂ�E%��G������-={O!"�dy��:�{d�_չԩH��-)\���<7��#�jOx�B���ӭU�\* eE���&�{���cE���`9fO>���UEFU�Y�H��s��2��!@�1��W�Н�b��$�s����a�GdĊ�\��=��A�b��d4R��#,��gQ���DQ���D:q{VJi��O6���Ϲ~}j(a�"��@NuC1��I����hf�ٻG�F��8J��CP2ч����%�CB`@�ʻY�\�@M/�/����K'����K}A�X�� nc���޲��;s��7v.�̝`4rNߝ1/�\��נ���n��~!��<���Z#���Oo�(�MP �{"�)j[����Tb峒��]���|�Vj�L<�4��#���p'H��hi�S7)�	{d�%�*侷?X�cV��I�TO}��~-�{��JT�l���ύT���tO��6d�@�A�73֏�W)�66�����hפ�}�m��$�*�)3D�:���t�l��*�7z_t�'>q��U���.K�yȼ����M�*容��AJ5~�8�}TҸ�[#���(��1O�JaL΃����{K��c
�1�N��P	��	'����c��*�p<ht���m�M*e�KK�3�'��Y��E����KO%Poy��<JC���.ڀ4�=>��o�4d�6����/RZ̕�	�*I~L�1����l��c��>��ۼ�1�UHLy��e���ĔӍ�c���ɀ�MVi����'�Hք��#��yB$r ��a �
��(M��3�~gf޻�H���*�nW��m��ua�r�W��3
1��eеL8���/��J)��p��fmI���g?���;�Dw;V�Ye���| qze����I3V���	_�LG��N�5�%���J?�yo��?-hp��tGH?.9Bt��鸋�n���U����.��@A��-��ٍW�Q=���R���kA��:Ix1�oD��XEbhE0�Rl�`�~�_0�9N�5��x��`'�	qqv ?h-�����Ţ&g��]x���8$
Kt�����+�߬1�[9WÚ�0����;�� k�`�Ɣ�U��W����5C	T�����y� �B���6�t`!2�����8���p̦��5gǜo��	)�a�p�'j�
�&��J���~���1� ?.Z���n@줔3y��!�z�N�|�vP6r_�	\tjS<��e�Y�i�oݻz�6)���j�	:����'���!M��[��;�L�7Kr$��U��p��m�B(]Y�<��h=@?��g�rК����⇲n_L'��K�a규��7mCAl��X^k.�2k�����2�b��`�s���V�%˥V�ko �3w�CF��*X��bqa�6X��=�de�4Ǫ��9��D�Ũ�q����;�^��hj�.��������3J����؄|�V��l��T����g!�c�.A�������R@Cq��P��>e)|%䱭>�Ly��~*:�.�']��e��R�G�-�MR��TP���%h2�E��z��pWƊ��_C�Px�ܾf������f$��J�����>ؾ�!���q�������|�BD��q��p�x�>+uNw�Y�h< �d�8=C��𻷁K�[ �������p��u���`n��pt����`���y/h��b���^��ť86C Q�W���1,C����ژ)ы�Y0��r�&@���Qo?0i�1xhW�(��������%bw��	#�������������4"k2�"~�tbOf�t4Цi���'HmS����?y� ig�+}��5U6��ê�:�؇a�G��h�,��;6�-9�Pd�l�M���_�n���C�0�͓U[�ʆ�d���n?��t]�i�<(�v�yV�o�Z��A����V���QU9oڣ��͌%��^���ީg�K"H0�]paW�y�jY�dr��P��7Sk!Z4��.��]M:s�}m�v���k[z�>Ϝ��\R�j�Vx�\�sQ�7�����⍵��ix}Y�\j��@2����7��r5���s����s�A]�<��Aߘ��wa!��w�d$����S�_	1FX�z.�ΛN�E�cP/h�4X�I�E8�=��p�`�t�?'��U�`�[8����P^j�8���Hc�|ǁ���g��<]�Ur�Sd�}{�E��$����_ዷ�Fk�-�2�@?;np��5f1�p�x?�'�t"X��YF�D���Y����wV~V\
�	�3Z���c�rE��6ϯ�on�VZ�x�!~dE�k1�P�1�jM!	X���rSS�N�	*�Hy�25��) �8QVǔ=��e��;E�]����.}��!jqv��b�$�W���Kƴ����L�d�k���
���(o�$��3"���5T^,�4sh_7w�DT�gsN�:�����0�:Rd�/otu�r�?Ȳ e�K.;Ke��K}d�|q!�X&�<4V3dA;]?��8������«�,lC��9�빃q2���(����[�'-ph��^�Ǐ�ܑ\v��z	̪�0M�x_�}�G1��xc���Ι���� `��*���2P�M����h�$.و�X�h=	Ø������T���QĎ"�R�y>�7W��c5����q�+���x��b��
Cۋ)�����^��tQ#�h�mƂK�@�4��߉YL�pA;���o� ��`<�4���'�+,�0��-�3<n[=�釪^�s���3��2��y]�%)GES��#������/AE�C?�|�id�|_G���~�K1ΒI?m�t\���1V�j�����9ږf*��B������F��`6tJSlL;,����mƌZ6��L���j�r�x���O4�n���c����oh.���*��f��뷑�D����_��~=�� ���Sr���.U�����g�-n�C�i�ѩF���Qf�n����@�AE��Y��uL���2�⓳� V�[D~ ݿ��!����e�	0�H�uwN[�OQ;�A��EE�y���b	���Q����@nѪ�Jf�߶:hn�V�A8d7����4�B��Ն]&�
aX��Dr'�d�jVx�e���s�_6��}�	c|;��a	���;���r��Q*��x��@��[e��s']�O�����-ƞ�YΣ�x����`y�)�fr���#I/0��ȕ����x>��?�&�%2��c�̳5�5�Nꬹ��PJQ���P�N �uZ�U�s�c��3�r��������R03�A�(�/њ7 ����ڤ��>v�0$Qv4���p��|�z
65@z�����g-;�#���\n��cw���q��e��g�<���6��7u��Թ=E)+.�@�	�j_ֲ|���hxl��� v(�9�|Y0d�!pױUS2w����.�c��8W�e���@�x�tC�:�9���z��d�v�/����>�s��0�tމ)s���{if4��&/���8h���������p�,�V���w��&�rs8���JQ�ۋ��i��SEcY�̌��2�HȄox�g���M�_Q�R�!\/�f�Y
��� 0�]�~�B�)��9�?�d3�0e˖����d���*��p ���iL#��u�~���<�1��ʚ���Z/ ���+C}x+AN�ҀS֮)}}i�M�Op6�O]���?,�D�Ps����d�E�7;�=n�F�[�y��
0 ����i7��pX+Lm8V	��x���{<d���v��g5��E�=��<�(*�M�.y�*�i�T��ŷ�^*�/KS]j��=��v���U�{����'$?������>���j�%ޙ����cK���Nqs���9�bBy�a�n���?U�r��RPkW���/��J=��?І� n���k��_�S���(_Ԝ_#���&�Q��uf?��b|�]v�㬢�����#�Xm���I<{dJtk�yAԛ�����������d᠀��5B� F��?N��%r-�~�g\|�*�ܣ�t��_�SĎ�Ǉ�~�(�o��E�]z�36K�$�O˵�^��>�=�LM�ie��J��\R��g|m����gh���o���������
nU���	;�e�xi>G�螧H�	l��^h'��V���V^�����SP/�M-3�=!~�a��+�Gj�ӓ%<�Ȩ*���th�����]/�,�6\i�E��O+�1����j�+T�į�B�Ok���@9$瘬���Q��d���\�8d��L��������wr6�5u���3m@%���3�ğ��ɘ�nA���<")b��| �D<�{����=�!7��ڜ����aoE�BC+Zc(0!�M`s:,��ob?��X��؅@���xD�:V���2����.~�X~�!F��N9`���*1�Q�z��%]iQ��E�&(�.	$Ĝ�dg���N��x����j���t�H�4��$�à��z�s٘4�}���S%�g�bY�c�V��-.}1�p��A*2������Gnz����L�Fk;�Mm�A�6x����֬�J��Q�	�E�Z��3����b7P@h��ި��u������/zB��v�X��b�P&�]����V�����c��������7��8�?l�u��v�� 3��Y�|��m���?�����y��gr�X=�}$G�i��d��3�wc���G��$��g��e��KE:�� ���(��K��p�aP�J�Dq��b�l���N�D��ر��aȎ1�}�ӹ{p��>�U�0/���*��F��﫭W���,T�R�s��H+�bE��8�N�wa;�Q.Ah}��S�S���a�d@�~lX�E�-T�vw"c��4\<� ��;�$-��`^G����4�u�NmP�'�^ �rԤ��|O��ϱW��0��Y���թ��!'	�K��O�xR"�Xi�4>�R��U���E��ȹ����P���V���9KT���x�UM�^ŝ�3|d�$�:�](W�����(�z��(�}�����n�\�1��%�����c�\���=3��;@�'��ty|�z �^а��_�8����7�slFE�T՚h��n�����Dm�y8�J߂x�
���^7�k]���g�ZvN3��k�;ر-�쐑>����n�M�@4,o*d�U宽��}�j.+�&*l��%���S	����&a{�s�d����%�
�ˤe�
��0:3f �R��c6r��
�7^_�(f�I�z�"{��ߞj5��j�K3[�L��+�kC/Ɖ�M}4�u>r�a�QܶD׵�����M��ͪ���vk����3�Y9+����l����;�Jь�s����ѡd}al�ț
�[���BC�b�4ӓo��lqo�?�&�h��
9m�9{��y.���ʹqM�So��܍���8 	��RLپm-X���\ �;ۇ�G�W.��M\����ާc�{���/8D�2*ќ���Z�z,
�X�@S�z؁W�c�������r<��u��3[q�}q��u�ĔgY ��BnA�o�j�ZT��qn�l}R`���cR/v5������$v'r~�^u L�N�U��IF�Fu��(�F���/�"�h�5���l`������h��k	A��s��5��0�����ʥgp�Å�e7�$�U|/O��)%  �ï(�m�Ό)���I�R���h��*U��"gq���L�@.�DW�^d*�k?:׆*9жZl5Т+���Q�o�F�����7o�PL{����%�/�����M���jP�1,��ؘ!�!"h
N���ĕD�wAN��5�<�R	�$2*kX�q���J|J�������!e�";��]X�㈋�+���}����[�I�X�z�UJ�4�m��w�w����hV8�k����d�����!������NԦ�� �;kׯ�KIc��V���Q3AO� _q���h��MC�>�..��y�t����j�9Vc)��vdL������d��2U�3��{P�ͱ#�C���a�V-�l�8Zn�hP,֐f�����~z�Í�^J����q+|��ꨙ��a/��zٙt���ߡ�K2Ʋ��q�7�D}Nkp�J���
�Ѹ@JB��4f_�e�D������ז2�MSFv�M�˩t��TL >4��^LY
�!>@�R0��{7�cSWW7ai�}�yC�m��!&�U���'�����g62� V�&��)��`���ubu`�a�L�♥��-�5^^�D�CQ|�Fr0v �k�����t��"r�Ď�Z�b�Z���M�:*Y�e��P3��tx���J�q ���(�M��e@(/^�9�jH7�dM1��ې��/\��5V������<��g2���@7����>��U�j��Ꚓ���ѝ+k�T�v��.�V��c��p��n〗��9��6�Xb4��Y���L��:�& ����w��6���D��ԫ���yW���9S�7̊T�h�c�x�ꤐ�(H6ht�tPbg*�l�5�|���ha�S���(�$�ѻ�XF��v�kPå7�	��T�i��+�G����fx��Oa䶈&lg<�Ǉ�8k�ʟ�l	��-�7Cv" {W��a"y�0��oST#���{�1��ih�s�cU��b��u{�[Ρ�^�ϊ��Uo�gѫ1S����IG���e���k4}��ܚ�	�	����9̌�O��s)�+���>���h��V�bmR���.0�:�2<�°㼢�""mM@��3�����c��ۇP��Eb��g��Ǳ��iU~�>����p�J�����N����=&���Wʣ�nE�����$�j���R����nQ@?LT�m�9jL�o��~�+��76�hji��(�����(��w~�����8$���ᨑ�r� ��+�k+����EJH�"t5���-ydoP�ԡ����u�F(�|Q���|��(��^7��M����)IE[c���%�5n�0�ց�m����̦�4�1�7�W<1��7�]�*�X�ȿ&2��ZƮN���Ƌ9e��#�w"b2�(�RQ���A:%쾑-V#f(G_$*sJ�� o"gp��)��g�A�$�`�i���S'�k01�UU9���� ,W�4<V�d̗H��~�n�H�>p=�n ����t~d�a�Ho{]�;H`��+Fel��_ֳ%*��9�pz������������]�~nĴ�O:(���GK���E�:� �>=R����<,4����a���+N�$��N,�:�
tѠyľ�T�M&��Yȭ�/�냟�[�G�(y��ަ	;�����bKO:v#�ZL���{�����kc������ކ� %u�;b�1�ʺ
�B(��}l��Л5���%��>@tA_�S3�X���:�u��^]��j�H�Nc�T/h�{L3��R���\@����?�I}ƲzI�:�0��kJwi�r�rE�E��	T����k�Q�g�UO�B̥d^kڵ9��P)�����x ����d���I[Vd.RD\.������K-�i��oܤ�)�-�Ş��೐�׵&s�.t�����ExZh�9k�F�Ƚ�r d�d����\�r���ڄֈr~T>�����כi�&��	�"��k�t����]A�"����7�y$bz��dG|��� #��-��9���w�>���Q: C����q��.1k�wV�t��E���_���_��@���/r/�9�k/�zy���B<?O�yݽf�e)����]�-�]jY�i�x7�:2Z�2��i=y��&z�I�qǂ�n��
\�ĢCP��NM�f��h-���\z�V�������ɼ��<�{�� b�Z.�-��~'�茥�ʑ0�2�q��JVM�MB�Y=�y/�?��I^���lu�=!��Po�=�<ej��3�!g��)�>պ�2�+�^���`��Iٸd��a��z���%�#�Rr��l{���[�3�1&���`�\FC%3������*oh�NM)/��Z�<ʥ������q(�F��y݉��8��@^p�eQb�;�� �q����K�W�`�F�̼E/\�� �opj1Pjh�ԑ&�iW�9 �m3_�79J�Ȍ��t�{����������+���}�LQ�L�՘���Xd�;�g�hS��5{�Ζ��&��b%�=|�O�?J�D�@#p�e�4m����6�_y����6-E�`� �j�,��Y$o�յ��A%�:|W-�A�����r��\G^����f
�V����]@q3ȓ��*��G��Fɺ����S���DBE)U���0��n��g[n�*�*�v�z��j�[���Eh�2�N�!b:)�pv	1�G�#A���	�:K}��`���Z���ߵ��.�TL�+�p}�|�c��3�cd�1��-� I�1\�<������%UB�H2ţ��#��'WΏa�y��Ľ��nc�޿�N�4�J�g_�	]90�/]4	�l�VmD�!�ו9��~����|�p����Z��/���m�r���p8�5��tB];4�Mއ��D�he[�0_��Y	��c{%3� w��S��U�e�ά�L�`��ۑuŵ���K�H(A�4�� ��u�T�'�:j��0G_�Q"�D8<��������T�Y�ƽY�˞Ar3�vs��we��������`���
���-�)s o�����!��%�g�?R�/��8���Jn�v7)yCsFw�}}������Wl]�Ս��QF)LL�@S�K�*/Ho;�� ��[Cv����r��c��-��#���!d��G�����߽�q�s���?��om��&^�&�;A9ə���L�YOw� ��M��5}5�'���B���*;���e3#f�}b��	�O�돐.=<yL� Y�~��|�)�]_��/1
�V�6�u�y���c�L�Z!6B����z�N�C9�_G-4j�lw��|<h$��3��V�SfX�����`��Jڹg���(��]��ܢ��o�tݻ�G��o����ӖM��|�]7�75EPЊ[��8W���w�g���k�X@��5��=i*��[���(��b��[8�:ҥS����>ݴ7���f�����+r�ŎR�l,�B���ic��=��lU0/m�U��ӊAu�0��Tߎ�[_��}��ٳ��-�mX�2����oˈOh�q9n�;$�(�3(�Z��>q�O�6����9�t��� D)�8T��c38������fis���R� �]��n�]�gƪX����Q:Q���$�='�4��n(N[KG����J��ҿ��`v�ob�Br�|�� d�Q�ۢ���) �7o_�勤�f��e�1���7�?ՖB}+�Ҋ�z�ZQ��v��M�uk�[Z�X�KXi��z�2~"��*�_&2�������H�d����8���o����(^����v(����f@i�n�~�\P�c�s�ՃQ6�)�fp�b���)9��y�?^�Se�B�k� �M� O�49AΫ/|`�ކ�����e8*y�W�X���d�ÞBb����� �h-dWM�j&���ɶ��Gi��)n�IlERV���0J�Sܹ�� �\���,�fYRFh��[��ĸi�b�w���ٍ+��1釞����8��`�m�5h�[/�M=��hϸ�Ěp���PF�9��6DS5�����Pl�����oϖ�齎N���'Ȯ�L�Ե�4�ⲹy�?5.@o�[ץ�qy�ߴ6RNT�`)�  MALK�[��3�
��;\�!��q�Z2�~V���C#�
��%�@'k�{�p�+���Z�_���*�o��U���D�Z��$YH"�U��%u:����Ժ�\��iL�������z��I*{.cD,�X#ʧw��yv|bų�$I��,���h��[F0��@��n~V�,��m'Ƽ���T�y���/�����ǳR��4�>i�v�H[-�O�.�Xa|���]�L_���r$/	}U)5nyb���(��/[ؠ��9+g���R
�+z�?e�O�,��?M �q���;�X�{4v��
glV.i�&�j�>���)���x$�������g��	�� ����C����!�'П�!�n�ğ��p�K���i��OM�@_^"��"{eN(��.o|�_���ξ��F�y��GޟڨK�5A�f�E���@���t�S�:�8y�pk��Yg�.C�!�푆b��k��q����m5�Vĩ~���wY�.դ�(���n]5|�^����mbF�[G�h{��|��"���frnT�K&��zM+ ַ�R�C<�����Z��� Fh�Y��g3�`LE�F��Z�/�0{�����2Y�JXblҳ�	D���# ����Hk���o_�/b���B��O7�!�/�@����}�d00�%�B&'z9����.�@�����Z��3N�����$�Bf�Ri�2
|S�y�R3����ްE4���	v�O2�����{����@N��	�
�����)��V�x��ӹ�a��$|�	�T���о�x>����s�A�]Rt�o�w���[���g��bGK� �!gBN%n��j-P%T%R�?��p��t�Z���Z�wV&|o��GY��P�g$���2u{F���jAA�aZ�m�]cϧ^ﶬO��iXSD���P��`ʻ���c+�d�S3�m8zČ1џlr�'�cR�����i�5�0�c߸�hS��2�����ڤ���b#`0��O
HX���<&�τ���j�(Le��"�隼w[���i(����)n�YK5��j��L����uL�����@�D:��y��Үɑ6+w|�;��l4	�,а\dȂ�2��Y\:�N�&����|ң�D����`L_�{$�qsA�%X�����,� ���Ӄ �vRT��tI�ԡ�!ӁR��~E�|��ڴ-q跡����.�k�ղzV�<"!if�<짝?��&�r�%�0k{QJ.F�Y9�"n��CB!>�R1��Lx��5�_�"�^r���y�Jh45/x����ˍ�1KMˡ�ю'��
5�V��Df��{k�]� �m�������e.q
�~��������:�S�$��nRH~��e��X��A�8�]&A�[.(�w�u�����0Lp��?{�we�89s�@_��V�a��$�:tX}#�$G���A�>a��q=+��^�}�'7f���<�yQ��q�n�D_j��L)O�#.�F��~<Y�ř��R�~�n�jy�ss~�y�?����p~�B��<�]��̹k�%;�&��`ELO�+M�Z�z�NYd��ҞP��9 G���Vw�t�類��$4H��iҌ)��(~8����i��no�4�i�p���NH��X��Q���*���S�s�+t�yU��ޘhj��XM�2�����x�P@N� j{T�d����} G��>�ڷ�B���(q:�M��P^GQ���wfW�;���@��_q����i4�	�̗cPC�c+I�U���O����J|����ʏ��k�$"�7>گ�A�Z����)Ef}=������T��C=u3��l$B���r�����fR�Қ���/��'OEy�*��&��#zk9��7��R� S���������wՐ��Ǘ6%
�F�4����.� �_@�Fe��lN-酯B�H��o3?p��5�v��#Uap`����ش9\gNA&3���Z���?��S�!��1(~njU���Jy�u�B�IQ�{)EHE{&��L)Ʋ�\�}���ǟ䂛8\9r��U
�� mm��Ⳃk����ֽ�ry�º��0w�|U��涺��k)G�!�Kxߙ%KjA�7kjc��l�~\A��?�}�M$�ja��us���I�w�x��Л�2�+�F��6&t����?J/�?*��J����� l��Դ�_����F=]Vul7kaY�4����o��������&#6�<?��(br��ݯ������d�|i��YKU=?W�6bm`wɂ��N�Mc#��/��I8Np�� `����uTY����,/pM���*9:m��z���=����T��wP{2t�R����\܁��h;���Jat��'I�>sw�'�q�}>Aj�q�8���E1��m�7N婮2"�WZ�������v�A�J�*�����9U(�Se�T ���D2Y�\G�ku�sp�o��Kn)�UԾ{	�=4��_К}��u�@v���Gw1����Vr4A�.���uV ���6�y�\��Ƒp���Ό��g�:?9r�i�#g��s�l��Ӻ]\�%[U������bo�.by8B�2w�u1'{ԆX6���kw-!��K�d��`��)��WGUfi���:_s���/��Ա�Y{Ҷ7�qO�v7z@� ��m.�C�y֕����<���2�C�\��@6nhq���D��Kl����O���X%w� ����߶��b�P��%L�9?yr��IeAÙ�.��6��%�L^����a?V�	<ڹհ/�7nr�x��J�=S���#NB�H��=s<�ݥ �?m��_�Q�ŬN0Eg0�⫘�'��<����Œns�%*���M��T����ww�K�\��o����x�fA���������y����0���v .��6܃hg2�D�~�����ňo�ѐ)��`v�Tk���S �G�	a���,�m�y'���H;+�<k!s�S	ٲ|j�u�vm�{�bpˬP�4_m�6�58/x=:��Kv�V̅
��K#g��q��󺢀�v�:���y�$�U�A��ی���ʶ��O` �_���[=��Ğ�4z8Fb��#��<���p���.o}���ϲ�^@EN���a�Q"*a���Z�G&�S�-�vq$���d�`�!;��C�Z�'|e���h�^���[�؇/��aP������ؓ���h��̟��;?�ϟ	o��%.��_*d����a6�Q�*tz#n���8$l��Dt���"W�
c6`y����k�f���8j�q��r4���d����D��jt���]� �Q=U9�ԣ�2��<�p�i�x(-i�p�D�����HEw��ĭr�=�)�[���o�ܘ~����f�P�������&rQ�
��,���:/�9�2<�
qZ�
�8I���6~4�9� �wjI�3r=����L����A���,Q�X	rG�a'���Uʧ�'�9�|��� ���G�4��|y����5_��*m#
a2��oZ�E��&��������Cwc:�R���׷�(p�$�y��o9���6�eo
�)bY]¢h��h�����yT����w�7Éΐ������>P��
*�����'� �b2'������89kOcU#�(W�Z�̃��߈c�8&yz�B��F���[`����|��!(��,��
��O�a�X�r���L��)�Iҍ��T]����X�y�ʓ��hnD�7\�8����x����z& Zg��������ѩ7���>8X��/B�07�z*�޲	��9�R��W���?˅xi\����Q�Y�
/�ߝj[;h̅{j�v���h��[�ᰞ'�wM����B�����
�=�mg�V��j���QWu�F�N�t1ai*��g�uk\J�s��w�Si^Ѷ����3��ͯ���m�/on��|�؃g��E���Ev���Kgk���G{�Ǔ�[��Nn��[�r���mH�i�9�G����y�>���G��t��g*.��Ee�Э��ee*0����+������&��f��8k1����al%���[D���s���c6����TO]��,	�$xdb!����$��uAbKb4�ϒה�U��7�A1B@S!=���,b~W
�%�"�iF���������
�ƑT�����%���=~,��c���$���Q3VL�I�Ȗ����E	fL�{J���JU``Ĺӝ�#p�8��mf�#�X
<�{��D�bu�7�Ob�����j7�[8?,�s�HH��(��X?s;f��3�ӫHQ(D�y�Jt�iupW��t	�@=�"{�\���G�=�J�0��!�˔�?΀X�.�L}���8�ϠʚXbM�=�z�l_,Q���d`iZ�Iשo+�:�M��"a���(���ŎFip^��17?�"�A��S��tk�N���@r�|��x��)�DpS�Qk���%�tR$�������p}׫�f.�m�٠t�52���Ag?��jஒ���-���
�vW������!_��.���u[�64������Mc���e�/�)��r/�� f��1�2]�"؆�������SP[ h�@>�kR�nJ��*I��m�oe��T�_�9�MWI�#z䫱�D��8���*��̐��(h�O3s��>��Zg���=�(o��2�N�I��r�94��A�=7-�5�D�B�3{���CSs��i�zm�Ѱ*\��� x�Q/�(�fv��; �����x��>�Ow�hN�T�Z��g��U5����;�{���~��֔�}�eR߁��v�-8p� Vg��W���a<Oh%�Y��S��/��P�-XC�������r�G����A`Rc��"��@)�9��a��I�n�!?���h팓�R�.V:Q8�OD�v�f�~"��0�P'�ZMl�������bm��!�#ıj�vy�7
>xd�]<���%V���w�,���`J	�1�ə����-E $c�5#��<�u��!˖���%�o�tXQ�ws��3�����G�UA����S���4�\��:���3Fi|��'dK��\��"������1�;�O��T�vO#*Eu����V4-5�>�S��a���қ�x��nȊK ]'.�(;]��-H�D�!������O�tx���@�>b���2�MLd��z�g����L��U�婻�[���L\�«��A�YQ�r[;��L��l�����wQ
������<�#;�צ.��e��}Y�ʣ��T�A̢=y��'CZ�R79���O��o/b�e�� ����˾1��2���1 Ws{�"���O-<�j^2���m����i��P:�c}	��r����8���J����W����� ����� u@D�*J0��L<�\���E�!n��M�o,�[�����c��Hٯ�5���pi~u��(�J�/7W;C��ʷh�F�uF,�ʗ������d�Q%�ɦ���AD(���9�>�c�"�p����G�r���c��ߡ2Y�c������[:��|4�8aͶ�d�:�O]����a`ڢiL$Y��#��z|gV��Z��B�.T��0�I���&?+��-PO��+�@�5�R�&�8!O�����l�g�k!Q�-\�{��Q��e���u?�&��
{)�'��|j�y�;��[�<��:
v&Fbrt�����r�V�eҬ[�nUۖ缆�D)������`��^�~�N �U�s�%�\�F�r��T��;{Ǘ;tc����;�=��qzP������Uy�HhǶd �M�į,I[+�_ǾN�C�1�*����竢�I��Kg����^E�1:��sn�z`m\G��P!W�~9� �6�?Wc����Z���Â����j��WV��:p�"�2�p��@g�F�&$]|f��s`��_Q�Ф��0�lȸH9�� F/���$�c���}	M6�f�vgl���
a�F�y���+3�/��S�?y��^�-׽��x���������갵��/f&ś H߳?�t6����I~u�X�ZEI�.�>"܂��X9�nZ$"�Ph��w�0���T�����&�����^�:��}�OF,n����~���:�=Ԧ�0Z�����i9��#��{8;vl�G4�u�h)2�Q�9��J�_�+H�q<�[��D����;��7���Iˋ��m��G� O��3B�	r����-\������M�����%Jj��y����������&V�c*���*�� �v�� E���c_bg�0: �  Km�I� [>���`b���=�N!��(co�p|�?z��S�2׺�G�4؋�^UJ(<�&iy&��^!�1�p�v3v�f�=���r#���u[dxs��]�,�}�&�#�9�</Qp��[��]����M����g��Y$\�Ծ�m�e8�N}W���π/W�3dX�'T����S��t�ϵn��ت���"��CS��������ϗ4!��eeei�շ�E��k�������Cf���%sF�#[^�!UGd�e�a �q������@K!Jz_8,�Q�4�4��IƵ��=f�%�j�M=�sނ�����Sv
-w�
�E���-�}���a]L����`�)'K�,�8�;Pw8RBr���l�q����8Ņ�	��gS��@�n�W�U�>m9b���Մ�!�J�[�c8���;F��Hk�^�Xg�W�`�?*�G�QW%n����o.@�4-WRA�*��1K� �����yuW^k�Ը����?�t�X�A�JC�F���p�N5y�X��Ã�Il�����(2�������2xw����x9n�=�����:r�]趚��D��%��¸��t
B��Fє�/:���X�*[#jcL����:j����aa����.�^����Ow�2qӥq:/.!/���4��?a��Q/p�\�5~���8��D :���i�K�����/�e��1�	2�?���0?R��	G!]���x��ۺ9J�2����H�<#���,	d�� �c;����I��5��k�GL����
�7*��8����*��`�����?�y�p�mNK����u�1�U62I�X�ڃ�ڃ��ƘUE���<�K��@�~�o�ʉ0����26}��v<��dc��Q��$HF!Jt��h�]���Nd�Ur�ꚇ�>�} /��mu��+�.�xLvb�1���_߀��ES^��Y8���h��@wR5�y������͛+��S1Sk�ׁ�_c�|S�m�y���ة�٣AM^Yj�SB: �t�h'}���GՖ�#�7y�-���<0��4(�y��!���
$�ρ�/����F�/�k!}���
^(aFl�H��u��N%ɥ�����
�Q�baa�x	ۃ�Ǉ+C6I�yg�&J��$�I��A����n���"�xA4F1�W�_X�]���c������T���^Y}���u�>	X��đk0tq/�S�O��"��;H��t/�ˬ �l?����`����f���w�[ޜ�*Hv<� [s�6�����T��N� ��*��|]0�6 ��a����cλ�)�|��V���vsi@��M�2r�H"F�u/�^�y��L����(�>!]KvˌͶ$d1��`�"))w/T3��M\v�rHF���>�W�%Q�V�����/�v�y�
�+�aU"�>�'h[U�uE�ז�,�p�[�p�
�j�"�֙�?a'$�<|j�f5]���PN�Jռ���&����H��鈆�\�ީWN2���g��/����%��~��'�!���Mc�%�ks-o���JX,�\rbbp<1�"-��J��	�OUy>����P��O���xr~ۏ���C������)�ܭ��ѲLmFO��ISo�;�������o�nPF;!�%�y�'�tˡ���ߛ`Bl�)s��Ħn#0A4�!�j��ۇ��O��Y�^><��,��b6b�جz�љfIW�/*�7����܃�ʠ�����d�yާ���O�AZ3��s-T�"} s>���Z�@Cn��:�ڲ*�K�!'pŝt�+o�kZ@N����ؕ�O;Y5\Qh�p<��{=�*�M�҈;�Zcn9�jZm���D���Bֺa�;i߂�.���=�n_.},�ϓ�k��� �ʋ��8��L���oL�}"�;��X!������v��ӄ��Y6�a͚AF+i��D�F~�pw�M�֟JfrQ"C~�FX1`��d��\Ĵp����Z�����3�h��1�VArS)�IH#����������)��p��0�MT�����p�-Y� )�q>�7^w�<��	����Q8C���q���o]t9Oig�!mE2�q�
����S�dt��UE6̊x�wW��v�(�Q�S�����;����)���"��@���օJ��UJy�1o�\��R�GQ���[�>��л�3F �W�v򲖉O.��p"�R��f2���{�,k2����P�gR����;�juV#W���.
���|V�m��>��~�gMi%h����"��Cq��n����1c�Hx���:.؁�t���c�X�k��g��P�ДO���!�c9CjP���D�1�J�ל$iDECJ뛲�?��*�g�d��n�бy��M�5e>]��Ը �}�|yE�ai{�?S�&i��|VΒ���Φ�W��tC���uM�`fPc�5���L�[|��Y��A'W<Q�g��xЏ#ù���R�>������
����\��-��A0�;�]�!�2wDG}��[�X�9]�-��f+]�mM_�P���o��PԦ���>�q���識nWM���y��v�`�V�Z.+��yeB+��G��(!!3�
��x}!A�L�ɺ�mD����A�q���c���9����E�{�t�k�C�WC>Й��X�t�"���-�3�^�䶞A|=�d��?7Z�a׾$�\c�eqT����ظ�,�𬮤�,|�Q�'�f���cٯ�y2!n�
��N��'_5xP˛qކ�PN&�eɓH�4.`�L�r�~#_μ�r���2��q��uR���z=���N|�~q�#�X�|���ɢ�P0j@��x田M�BT�_?�>��i(�L��w]|KP#������;�R��Z����4iʐ�n�׬�9I����θ�Q��A�F�
�6�kN+��<Z|^Sl�M!lj;إ(��E�7$N�Z�Fz	�}V�H�l)��f�bnXy�e���\O��=�&'|Ѻni	T��#��ә�����À��`ފd��$���i�I%��K�+�7%%�sP���g.�0�1������l�k�/�,YY��9�ֱ�ME��0XI��vJ��^�4�2��yEў��7�|�&V
V֐$��Q� ��:(�
�yMDh��6�9�!�5�:wP�ZVt�>��爿��B���{�di��څ�ގ��K���lKpL�C�K1P��l�%6�E^�3�c��d�G�!yVi�	�b=���kRFI�I$œ~ݘ�J�'5"��۞]Dh�S�J!IR{tZ���+�5����yk�}"�6�tU�P/ֹ�Ҷ�2B&U�H#A	���n^N��#�2��=�]Y��W�mO;���u�rc�*1/��6�O��sV�� *��j4�ډ��\/ղp>��K5�)�n��hb�!�xw�ߔ�7�ҷ�|N�Hg�T��[cq.�V-�E��Ɨ�`l�:m�z�ki)F������`T���*6���-��طo��C���\rJ<�(P�≢������ڂZ�^���;_J����aeL��%���͢��0�t�P��>��4ΰw�����1[6V(pb?��k���t����!��<3} 0]L�h!�=�N�9��u:�5s ��������t^���8+���/�6�W�v(D���D?{ HLgSo�s9�KQ� ��P�C/�2ޡ���?�g��3V�2��	,.7���~�r��Sܬ��Е���~B� �W��z؄�1rc���8���a��J  ��}�mА�H,��"�����
�)��G`��颙l�6���'h�J�+yd�O���-�+�"�j�@:��#����ʂAp�#�›�l�g"�+����LE ������h��r��@#��9�pڋ��js��opތ��'�(�Ts�:X/�}�6�)�j�4�F�:��#&��v�8����ًRw���[�0|����꣐��R�M�s����"�)V^P����J���7M�D������R|%�̈yz�H��[�.��9H��w\�Ar�{�97_��,g���I�כ�B�*b(ױ�r3�����X�fB"��lHJJ�V�Cx�.�j���������m�Ln��QW֪R�Lc8GV���`�afP��Y3�ϠO���Ӕ�Hd��( e�x��ʪq�D�Y������c����]b$����-��FIWWWWDhP,/FKW�X��%�⣕�~q-z��Ң�;�J
'z�4��k/��.�s�V��{����'��|�r�7H�]`	j�*(~�Ȩ�T|\���<MOX�~�x4R⋴F�+&2���ү���?���>������
�V�@������Kp��37�m�𐈗w��܉�P����)�З�ɮ�ģ^�� 3�w��Q4ʼ��duS/����J�Q�9�w�	�����@"��[@jA8�+fЂ�8�/��ѨS`�tQ�q�|�~,t��(-ş?�|�f��T����P^��9��ݣX4�Lb9���<������8��bg�&m+u���?�g�,�`(2��,�Xdu��ZWs��Ȏ�L@���QYЛ�ğt;(.T:�G:��ݲ���a��7cg㼧v�В#�K��[�E�_3��i���+�Ʉ�4T����hb_��ц��t�m�����R�E/�"s�i�w��O�(�s�Γ�Y�]�L
d��yQ�B�2J����*���,Q����,{-i�>��gU����\��M���Ծ^����?oPY�-z��&;�^�������?����8UH�Y^�$AX0�j��t�}]>\�7�b���2�7ɹc�;/�^꘬٪%�Y�����!����<5/җ�]�~�q4���I��!ȃ��7J�A��|Da�֘�k��������4�$�Y�p��`�?>A�鎎�"�Dk�tB����) �W��aV! ��u�! ����xq,/�I)F�5������F���m<�9�~���B�x^fK,�n�i&ސ���h!�&���f�_S��(�w
�rCtf*)�>a0�uMh�1%�GIf�ܡ�Þ�H�b�6�.�XR���}��q�S���v�5Ք�py���v���$�pj�RG5�t���jAh<�%W(��]���Zm��ԋ#z�U.�M�=������v��M�oQ��Á�hO���X�i�|�R/��jgA�)�PA�&��]7q�:�����=��b���o���@;mҰ�6���2Ps����/#�?-l�e���el���2[�ⴊ�S��W���3���{��6%��H���S]ƖB>�ݎ����
g�8S���_�"O���S�D�4jT���<���`8�́D|鮘8�<�E�����2��s����W�vq
��Ǟ��S?G�<3��F#��j�bۖ�\c9>^R�V���ϴO�&Z���4b�M�B���{�N��s�{�_��"K���a��3�k�t�o�k��l��I�
�C�Ꮚ�����Y)��Q����1	�e9L`h�1��/��Hqgf�������ǿM�\�X��o�������5�4���SMR��>U��k{a���oj�1Tϟܷlq�v�K��h���.�����������C� Q��2�ғˤ���c���8d���s5�V~ZW��О�pt{A�P�젥DDp�*%Y�.�ʰz4*JA|)���)Ro�l�Ѱ-�wD#˴?Sb�ͣ}�k���M����S��o�QȖ%Y�3[����a��qr�揃59�\b�^YG�3�,�=_8�}�9�`�bRu�����s����/q��ͦ	B��ʻd�O��؝]�Vj3�l��	�U�ڃ^�4��&9���5�&�|2��\�醠c��7k����� ������ft-xi�ʱ.��m��C����0x$|�66r�g2B�>g� ��|����el���!�� Y1�v&:)���	V�3��.��0��k��5ƒ��<�6��;`+�G(�����*�6�R��~g����w�G"dwH�(ƨmFV�	��������Tf��g/�}v琳d�-���2��ּ"1e�1}J6h����ύk?v0=)�$3�՟]�I���U��Y(4�B��Qd��v���Dͷ�RO��	�Z�g�5���ຆ��Ǘb����T����u}n������u�~�1�Hv���"Ce�H���(ܙ�4�k��~zI()Z�`$��?Hyȃ�q�s[�QT,C�ʕە� Biv������C���\�j�CY�nNr�n&5�B��)�@�t2�W,��	���C��l��׫� ;!�5��j<�\�kˎ�6x�Y#�=�Ʋ>�)j0�
;M,%��YSh�K� �-4Ɇ�R��&�\K	c�s��{��L���$��2�أ�JT�{�2�kލ[���%��`��R�p���I ��[��F9n����L��U��c�d͵L�ƆĳfX�hݥ������ح8^K#S���l��O�?'�T��N�=�`K;~�ֺ:�.����w��n6
��&���j���=ՖӅ1��*?"1�F�"����$����ㄆM�a���fYo� �L�&�v�J�lg,�S�0Ω��&�:z%������ �˗���6�'ZA�	kV	��7:�qb�H�T�DR��G�j�eHϽ���9A����gxQ�G���' ~���n�/.�)�[Xc����!c�ʜ�j�l@z�X�O�N��B�ޅd"��sDb�%NH�E��O�&��w���BMK·�*���rz>�sH�͚x$۵��u��o��d+��ֶ�	�o-Q�Ku�'��0�[���4ݍS'wWW#B8g�'��{���?����y�9�������n߲�=)��O@�Qz!cEɌ�#?��!Ar��}(v�?b�a�˰&�j8��#��;�L�^Y���:��L��6��n�f�}�U2�,%D��c5/�z��t����Z�CZ̾2��E$ʋ�X���,~6\St<O�y0����o;$sȿxK����s�{�������̆��B6�%ك{2j�⤁��.�'��ٌdoi���CQ�e�N�#�pD'�,��.���o�O� ��Tr�Տ`��1:�:�h+I���6a�v���D��h��1RB�0�H"��7���u�+NZ�i{�[q����K�!<��+�rq�&_3;�L�|�`�כg\�f������O�Z��߭�v]vD�l�E�m�����
��ҸG-�Y�9V?�I��?
t�gBo��E+�����
(B�9��g�-"F���/~äi]���s��q�_>ob�-��k��<��b�M}�����7\0!D���X���;����I|�G��<c��_��O���!��s63V1l����P*��CG�;�a���0e���Ti�9�͗��gh�EW6^�*���G�s�֟HHK��|E�a901_���?4�׆��6���V=[UmA3W�fL�#�E��:˿��'[�F´L�n��?�/.�<���4�6��^��F�|�R���6�-Z7�d��dhF�C��� ;�̩_�lK)���
,�jֲF����O,���������V7=3�#,�T̈�H	�ޣ��5���2��Z�.���4Y�](�����A3{��b؝=x�־Pw{�|N�L!0R����� ����<e��ds<f(���s�Y��i1���؉a�E����8�X��f}�-�3"�:���ݴ
�zT��VRCF����a�G�_R��w��.WiNVO�~�ˎ��-e9l����{�5"��$T�C�	�:3��=ɋ�M��9\�&�>��pgG�-�t"�*�����:���/�y�w��1��'t��(���HT$��p˫f�xx�qR��δ[�b�(�ɨ��Օ�q�H\�O�E^ouB1�е�s8�a懇��+>-lN��	��"G{4u�����3R\U�����.��W�BߙT)��|_b_�n�JE�)� ����jQz˼*�)(z4/����z?�G�\��;\jb\	ڒ�T��>�����y��f������m�R��D�+9����;�V^��� =E;jP[~ڪ�Z��&g�5_��#��ΑUϐ�T4j���Ӣ���	����Yݼ�����[�@-rM�]."x����P����[��z���Q��1��M�%���{��F��P9�\��WI�
#ĈE���_�0?��>���C�r�����](�lz��M���й�m���	�}|���ᔨ{��G�^��ٯ���L|F���pJ6������Ɏ��0	8]���E�RQe\gKP���]$J��C,��\a#}�i���?1ᨎf4�rp�yd?��o�w��BX���,>е�u�;�{�$j���T��9_X\��$Gv�����{��˳�p�|��Ju���7)JMC��E�tj�*����k�����ŝ�(���ݞTݸf�u;NWpy۟^���T�!�����u����"�Xn\������S6����\��m�ʪ��9=�}q���6�mT�鐔L�����LO���A'���2�N'Y4��`A�.(Jq8�A�7�PT������Z�1��9&`��u�����4B;V��?��[	e ߏWM����N�Kבϴ�nCbdu�y^2��c�p��{y.5"��Yh���A"ï0@�W�fl�Ѝ�9Z�fq��g�zJqF_�yI �5i�n{3�щ�lL�PܙVVt�e�PŅ]�C�J" :$��fwy�Ղ��/%[_T%sf7/��q��W�o�a��e�:��Y�&���_4"�bgZ �>H�٫3���� ���SNX�d���͛_��-H��IE��r����瓹�y�Vt"�p��:�W��!��iz�`u	רs@f1��$���1�nU���n���` ��4���>��	��	|c	����Bq5~:8V�H 5^<$^���ı`�9����iJ��ň|g�z]�n���s>��D�r2�sI��e* A�>�Bv�G�y^mz<���Cs:?7�k�]R��;�d�A��ܺ��0���f��� v?V�F��E-d�\o��7���W��/�)�_��c6;�+�y6q�Z��z3��Q��p
�9'�N��`S��L�g��V�����.��g3��%�ǃ�`�ps�����9��A�{�����[p�.`�\��u~���W���7~W���A�јDY8�d�{4G\�����B��K���ls�Ƕ���<��&VG��GT��C��;J�v����G�G�&.������1�`A�on冯�+����0�?�C�W.�	������7�O�_�}���V��8�� � ���k�بO�
�`��n���r_�k� 7	.9���ֲ7��sR��q#fV6e�Э-I8�Q����V�'�����5Ф܄�h����]/�*�yD����������	�^;��4�=H\�l y�ߏ�;�n���Ga@
Hה���W!/�� ��8�z_z݁�k�waE~\ΐ�TG�<�A}d'5#�T�����p�/�u	�:b�z�>b�ɲ��X�L�������ff�ً��}�J�A?	���9��-����p����a�@�;M$�G��Z�Z�'�����ʕ�8��`(���$� �����/����8Y����LYi��1w��AT��k��G4R���C�WoAL���*[@B�brOY��ms����S~c�SL9�bDwZ����4���������n�;�=��2z$��
g���^Z����PAS���/R��]�촿��}�����c��̂�(ĥD�E�^���[��3���@��!<?��w���{;=P�o_�ݐ��.���9QY�<$����F"��z����V����K��	_ 
�8�씘U9.��PbW��7q�?	�.�b���?GҰ�������BQ�8�8�V��(�c�c�T���J�o6ʤ�P��>����t�)d���h�=�TWʈ�c�V�t��}�;ɷ��__�T$���n-k�mz؟N�X*���T2l�7�{���X��\����H�)Z�U�����?C;�)���ߒH�7��aS�þ>a#%"�H�t2C\?�X�#��y�t$���l���H�����k��CXPi�ϕ�A|Q���8�wm1~4�|�3kN�@�t�� dxK�d� 
��x���B	(���1��@r�Ϸf���/�aw���r( �To��W�^/�1��"�uWp\�4�s#�O}s���2ܲ�s��Wq~D6n�n�}�y�A��T���7zȶ�&9]��+d�n#�!q~�	��.$\�^B-/��v�_`e�͍��f���bX�����}�H (��̼y�%���%y�.�lwm[����p<g�o�E��sڬ2yӒ����;��u�$��#=�V`=]qc��*�XL�̐���-�zm�z�|q�A�6���9J����G��M`Vߝ�	>M�E~�ͿV�+#�zo��BQk8�<3�����Z�C{�uwz큛����-Cw~2v��TP0��W��כ�eSǒ$ͣP�����Y�����ħӿ�ux�@����}�k=��2"ǆGf�y�g���R	�	sX���E�W��n�����1mA���V�� 9�4[���Wj�}u� ����a�x�LNs Ẃ`uk8�%� ��x�[��F��g�1nX��g�X,o���bo��h��fVB�2��yU�!�z��������fG�(�aB=�^�pZ�8�]ĉ�λ�=��v<��&��R��q��o_�U�oT��(��-����r&�>]9��O�.��Y3��"���"ʅP��1�)�/�?�a�Ah������HMݪ;4{vo���U|�C�	�i��@��a�CA����>%���L�1�@�E�|��yB��f�F�O�t�l�;1Xnd�Z6'U ���Qk��x�Z����Թ)j�ֳ�� ������禾Y+m?x��W��I��an(�G�6�v(@s�ξ�.n�S��|�9� (�b�#*���Y�t�'�ׇ�p��F�ޥ�T/�l��TACu	CR�*~s�����|��IpRS�y`�����-��㻍J�,7c��@�q����#��6¶���r��X~����s�w!b�sq���Ll�z�e4��0bI#��������n1AyHkY"��N�g�[��ޕT��(B�j5�n���2]P2C���v�}���m� , h�7T�8�1p�%���tV��ܼG��g8U_�3��ئ"ˠ�S\�4%�.M�n����z�\��m�Qt	�E�]^�]��@�~�+VP"qȈ��%L&�!�y=3�ԒU����e`�Vs<��X���ߜE) �o��U|��"�^ne�����Z�}���_:�%1�w��bSJ�����B��M�u�E��F�	�JP�X�T������5��+����@BVt�#�|y��qu�T��&|�5�c�l��J��09�h�h�ISj����� ��A]�@��޷�'B�����d.�[!�ȵC��SN��)�}�����7]��;�J̺op~e���u�?Ҹ6]�������:͋d��am�8qI dZ�I��C�t���B0}����[�����q�R�P~Tbt�sv��4�qU��	�5VtRfR8�t�K���lA[[-�?+�8vں�+�i2��&.U��<�ֵ�Nc�.��.w���f��k��c�h�� ���J�_�C>�P�����y�����'�H�)5��s^�)����TC����a�%�U��售�N�Ly̺�������ځ.1"�����?���J��zeQ��~�@oP��<�d�����Ia�������[�F/���mO+-K�򨂕����hV�D�v�
�~~�Ї�d��o�ۡͻ
umuh�ۄ��"*C��=s1���O/�Ӭ�#�;u�kMJ��E($H��$x�/G�ƨ�as����0��S�L���~T.E�ߡe,Qě[�F\{�����;жj�����-wl+*�f*B[Myf| �IQ���D����M4)V;�I�M,ߠV]�Y�?�I�{5<��&�� �pW�ۢl΁i���3�����o�'P�lqu ���a&V�����u����8�=+	�3]/s});@�G�ʗþ�ߋ����H�FfLMnl JI�]��;X5�9vjG�-A��L�Ѝ�@��LO�WB��Tq������Y��=>']|����.�k�9�1��* ��d�'�����8����^x�}ҟ�/kN��� A��5�[Z~%sPV�~�������l-h���.M���伨��z�=�[;��h���KTT��ԾK7�e��»j�>,EEG���YF�A|��*ۭmh��1�Ȃ`/Ge�S��{
�}yY/p�˦)c��И��/�un�_�����z�����D�ӀF+�^.�wH��96.	���tcF��};�j�"H]�C�mx�Q�����cB�{��^*1�xq
I� �
��Ġ��Ў*<FBhX���Aݢ���>2�U'o����k�B�"O��Y%��@���f�M�+
X��,&S��n�����l���X���#د��ٞy�W�d��G�=ƁT�{z�R�a���_w���d��Xĳ��_��`@�S�����S���iyLx��6b�V�1�S��q�c���ki�6��]�~�'sͷS�J���)ȏ�Lu3����5�o���	�#����g�G����r1Ȁk�� 1tp���%T���+��x�̖Є֎�ۗ<̋\ �!�]�q�FC!�M�S����JB�l$�v����`Z�:�\����	?��@����k���s��#�ߓ7�r8S��5	��|�&S�9#N���������V>a�M�Jr�?մ����5�7�,Y__��������蟫� >�7���|L=��T�3����!���4�����uu�����Ycw�R��Z�������(nw��]�\B�|3�G�c����ǾE���M}R�>Է�555�������͎p��_u���]TR�t�U����[EU�"CM--���X��[�����)r�`+K��_�4a���4�� ��ZF*AS�2;}�X�K�ĥ�"�(��%� ���Q���7�-n�q���(���`*��}<�������S�ÈU`��FNo�Ɓ�q��!5�rmq0��M5o��t͝��[_�p��\��M�(��\��m&b�ʐG8�޳�x,C�pxޱsU9�#��_���k��E�5����۞�~v ��OxV��D�Lx �����@!�J�1�b+5�_�}���rm#�2���`�p]@�C>۶`k;�$���E8/:c=�l��.�>�?d#��|ٳ�j��)����<�?����`�:[}���>��*��"�ҳn�_FT1[~蚨 qa�!�{�xq�Xm>}�Щ���D����t���9 �r��.ZJ&0'4��3�
ӿX�x�Ɲ���B*��b�&�����{a�n��;C��n`=; 8Y���-sg�����Em�QF��#�ݠ��syw{k�|k�1͘iכ|���N����/Q9���ğ*1�u��C��"�Y�<�V[r�}Lc�٬����"�p^A�7��8��6[�'���p���w��"��P?�	��S �$�$iH[Ne�ccTQ8���u;��y��K�Q7�98��3�T+$�W��M��N����LWC��eX�j<i�:;��0�>}���m`I�Q����.:���ƞ�WB]�"|1�be�4�"�P��~��q��Hr�0�]Qj9�2��f�oς�'_y%�x�n�ųv���^'�^�e��̬�l��]$ml��u�&�<nR�m̥܍V��$i��c����S�ܯ5�2�\�/IV�����C�!|��$�l���^��+��,n��a�*Q� ���-{�O�˘��L��:7����{�J4����w;A7O�y���I�d�WJҍ��O�M:F#p�t�~b��=���^�TB��Įɗ���Un�<b��:��D�)�v�����H�f�:ZJ�nw��Ы�>��%B ����K&Z���[F��;'�/���C��2�����cm�fWsJ�:�y֬-�{s�7&���FEr���sL"���Mm8V+0� o�	O2T���/�<���^�A��ԜaFJ;�$׈N��gk��U1�qR�"�׹:���B��V��]\Hٯ�7%c)��� j��w����~j(r�ER@�g��ūeX��}0F��hk<t+�K�*�)e�_%7�,�'��|��6���S���O�n����s���R����`�UTuW�%B�]�
<�(�U��a�m ��&uŔ	v@vE�]�����S����,�����F� 2|��V���w�cG�:�5�P��3�Ab�]Fb]S*Co���>�A��Ce'`&�:���	[ӹ�ia�8>�-�<�~k�d>L�S~f��e���4�WLuR��Z��گ6�_��Ⅵ���o�%2ʏ������B� ��cS��q�gR�~�;�	D=����B��y�x��c��k���V��=ŗ��_"m�8��t?׎��%'a�ղ-����wV-�tXJ���=�����**���۞���k�Y���{i���HN�=nu����:����c�j��/��U�\��n=�ȾyK� f'@h�0�5�|�X[`�L�J�j�Kc_9R{�9�R�W;�����?�����6�>��VEZ6������!�4���J�"��6l��Ɗn�7aa���JO>�M�!ހc�4��[OeK�|�&r��C���:й�M���t9H�������&V���55��/�ۉ�v�u�Q$u�a�m���K������/?-Vg�n�/Z��yaR�(���e���A��`�דf��
=�)H'Ѡ��]䡹z�����S�z�AywgVy��� n�V��n�.a9lŢ>�MXQIvn
�$e�2q�?��t��\�&c=�ǘ~�#/����+�����7P���o�O���p���1�}z����շn"A1FJ_��h�\G��v�Z��5��e3�7��*�]���miH(#�'[�bv�l�U��]yc��W�������/�<-���%����+�{Jey0	`�WQ�6�<�t߿�9}�@Oo{6���m����(,�jl�>༖:��T�yb�3��TK��S�}te�`ja`���W�e�K �ʛ�cQ��6ݲl���x���,�F�Ѧq��8�jyF�k(�EaS�����3/��9K�u�p �`��q�Z�Ӛ���m������)��=�h����~e�P5�o�0-*������g"1m�d����#��R���:�Rj'E�ȗ��u��F�˄��^N�:1��1pK���#���	�
I����E��+J�T���i
�C�+�H��{t[T[ٚ��)��o���,���P���EQk�gB�����G�����*��d<����D���FO�&������SCG~$X��G�t��8>8�b)R�-��)XO(ADS(����b���("�%s��,��8�n�?���e�cgg^tQݿ�����ws��l�Q&'?�[IKn,~}��r�F�5���f�yi@�v���>�2t�LD�s�O�g������K'�ȟT;|?�/i�������|Q����na��%NEp���%^'��.�K-�P\e�N�h!�{+U�q�����`��O��Y�\o��n7CPC�����%�ނ{ֿHQ��M�5����ޠ^��7�(ռ�s�����""�\�E@��g E���gB�� �.�g��׃_k��?����g�2���������I�ؤ-�K���(@��DK�e�v�#�A�\������r�G0o�CC4D	naR�*�#��\p���Ne��ˌ
*�ե�IBW�0^ŏ����AҨ��짘k�z�G<��3�1Ba�nn�����T�����=�+.�#R�	^I�Rͳ��!���X�F�?��ω}��v�t!{,p\$�9����=Gl��8��F~��.��yj��;6�/'��@���R<g/~u*�[�����]F��i���'*�.�x:�E�[^�n ���V��r��/��d��
�H�(�{>��	ʗ;� �Ι��j0�����T�{�2KHq@�l_�=#V'&�h*ᕲ�~@��[K{,��Ԯ1��X��tɞR��?"��'�]m�;��;U'�l�D�GSn$�Kt<�G�l3�����<�d�#ª�
~�h�乧[��^B�g>u�������gmK�M�1���)}�]ь����|�*U�ڏ�u#2AA��D���<��������hF�y?hH�V�5��O��:�����Bbj��oSh��&AX��UGтu���&q䱷���6g#��1��^�5��ܽ]���0Z�;P�J
�FP�
��d���k��ߝz]�ELmg� �h�<,�#�M��U�Qi�1Gh�mC�^yS�v���ZV��q{�m�ǂ�j��h�G��vO@�ǳ{���t@��X�����R 鋴8�oP�l='W�B�R{?Ck|�Hz�5�#I�ȇ,�D�ec抨�)��x��2d����ֽ�9
jxs=��� 8*,lf~{���̅�0_"�F�BFk�<$q�ο�'�Ƌ]�� َ*�д��D[�a���ǀSv1�2��:"���¤y	�9�:�+�����1����W�Nv�X�\�֌{/t�Q+ڠ�d1LI2�`DO���7�Y���Cw(«w:$!��H�ڞ�T�{>��~aZ�R"��ay�T�=E��ƶ�~Ю��V�ݧ��6*���A@CT��c*���Eu��MC���lA��ч�3,��	:��� ̖d�@	3b���%y�����Qe�9z�kV�S��O�hSp��Ê�X�i&M�����[,�sX�[���`���-$�Ű,���_>�.> ��Q�6�uB��� 	Y]=-�8<��Tw����bԮ
[(��wᣞ��S�Q������()V��y����H'Pc�����$���S�I72K�zpk\ΣVZȋ�=R��x�=�k����9��m\��F��l������M
&�ƎO��$�j��IUW�^�B�?��i*����DY��?m}aXָW��S�B��T��`<����
j�:T\�%�)o�杆|�`��9��k'̃l���oET� E��L\T��ڶ^W�T�9q�l�
��c�,lx�6V`*'{ǣd��IBĎ	��e�'
��[��$�`�4(��ld���q{ЈJ%G���+�,�u
��A%�l�ILZb� Q6�xGy��,~�y�q���k(I1�����, �v�����{�+�!���
K����JMoھ�H�e��{Xn��عax�����<C�!�o$:直Zý��T�p�U�xP���bw���g榬7�:��z ?����K 3�������,v'z�&��\�.1z�`��q��;G��CT2��gI�}#X�C֙�x
��<!2q-�X�U��~MG!���!�I��M,Z{APtgy,P|�il��Iة� g�ۦo�O��r�W�*8Y9�S�������I��~q4���'�߱$t/��/~I�K\M�?�s��@az�aj��P��$l��,"7��1�6u_�e�nN�f#���Fh�z�q�/d���"���8��kh~24t�z�vL��)�hUΕ���^_���m�@�![�y�S8��n'�KN!L�����p s����;p�n��+N�i5���z�Ad�r���ɡCP��6�և���<�r�v������r���Ϫ�S�>�0��DM�!�;^����rō�Tೊ�����O� y�APF�Q�����'bܸ�X�\�K�&����TV�L�БZ$�b��"k���p\v���G&��c�J%A@m :q����:61� f�&��$��"���*?1'6A�}���ׯ���zODn�����U�1N��LyGRe��Q�m���0y[��XL��<����YlL�S;i/甾�j�QH�3�_��w^S[�|(S�L���1�P�L )�r 
�W�5	M�E�%hfA���:�uG�-�]S"�{�2������v7BͶ�;�c�4��߄>b:�]����q<���JnR\�{��\h:��=D�[]�,�)��,���.Dّ�M0y��`�_h�ݙV{Ȼ�����á3]#�oXC	%��J鼑,����N�qC!`�0o����(�e�g��\�N����Se��]`��F�'�;u��]��" ��?<�>�������j�;)3@����F�EY��Dh�3׉�^����~��r[|�%*f�	n�;�����WH7�RnEL��ޜ�욕)̔�9������"ϤeJ��5��`���ӱC�=�0����;�� L���I��U=t����꓋�w�0:O�&�-�$���?J-Mku�7��R�tt��)������ �XKy�v:���h10��Q�Y��A�JD� ;$i�L6��:�z�ia1A�&e��:�R?a&��P�Ǒ����Z���c]+��2�Z��~�Ȫ��\�Ή*��!۠i��K���@_�K'1�fd힦b4m4�}����9�g�dV\�^�߱���n�fYU�|��Zү�t�%#?��{fS$a���^�G��-�5����p�;2�s��l_mBnл�?����`�V��6�W =U Y�՗(�!�]��\&q\�U��[����9Էv���~m
:#�;W4nUg���?��%�GL	�v��?�+ �邑{r2V��s8���#��p�A�7�mF0�P�˅������]�9B�_�E�i5�8�����E �YT��GF�^����7|���Q�!��	~�%̥7�h��Ԁ��1�zc���Pl5�u�d���z��Y����'*�*�켌=;�`˶�N��1���odK����D�h?���n��	���M����-
͐Ծ��'����<��|�\ںWz��@S�/_ �#����O�V�<����񪼴LRG��HHܕ�m�\��o6&�Lg���5�d&��^9��)�*��������Bw�����m�`�z��<����)�m���M
Ӱ��O�pV瀷)D��js�c�d`���zɦ��#ekOw7eYF�ϸ�U͡N��/3>\��gE�6ˆ/\W.�6�Z�e�)�U���K
A�N�4�+�\{LN�]AR<�����7�p��`O.{�?�_w�E��6�:����U��3n�Zq�l���
o�"��ߝ �4|���sH�����+@i��T�y�� ����Pl<lK^,�PiEd���׻��x��R���gr[}����d����Ƹ
<Y��jʓ�*���U�V\�j�z�Ps�!�W:�`��9&���*�)_�n;��,�NȪS/پ����3�,̯�ן}b2;���C�5<��)6�T��R7ze�<o�SϘ���KKu8�Mbl����έtʇUoK���P����e=�{�7��&S��5�����~�D�(0L�C@���G� �}gSOX#�U�"+�X."�F�HC�	���
��Pbu�2EL���c���4��Ck�r�O;oKz�����-�Z>��������%_p��p�b���	��Y�[9��P���=���}8)1�C9����s��w��i���.��*0j��l*�M�#0�Z��.�Z�w�mn���V�N.k�F��m]�joѢ�Dc���o��9�[�-[)�x�ƒ�_��m8;/:v��|�X#�ŗM�
��1
v>�y}��h "ߗ��LbLo���_7���m�)^���_��H��\�+�;2�OX>5� �P��2� `@��:DP_���p�|��P��r���&�:��!lRdʴ��zQԾ@��`$	��`_Rl��*e=��;B#�u@5�c�&JѾՋ����&��}��2E����h�qF�S]�Ʋ{ra=��Zc��\��ɲ����<��!�2y���t�f�v>H��8|R	�Ѣ�"�<�l=΢� ���B�u�r�3�C9+D��/�A��E3�vi�0���Qj�Ep��
$��H�I���7Ln�H+�?�;@-벅�*�x��ZJҢ��B���nZ���*V�x��9���g3c#�׾~�'&��X�X�g�Xu��ir�x6���w�p�"��kX��^��֬���
SY1��?/V���j����n��}�rq���<��_���d��M�T��%�ŉ���wI� �͕���YD�,N/G��l��y�h34��.\�]���DN6��qVڪH4��;�h�=7_��}���)�(�0@��]P�����#�@���,Jr#m���K΅e4�Q_C�;�8z`��<�^��.��z+:g��;�y�s�ĥ S��\���I4��Vx����2W�򥽝޲�鱼�2����w�^���ə�s��$%�m�Ұ*�A��!BӾ�͘w2UF�a�T�ڹ�@�������U�Eh]T�Ȳ�^Mb�\hJ�+(��Y��є�5��N�!��<U'5�ϓ�Ϯ�����a)Y��Iņ� �B�y�?�8�1n9k(D)�t�Z�->$�r}T�����ݳ�sA�K�!� 'ak�p '��7�v�\��ʺ�����X����v�%���L?fٺ\��px�s3Qq���3�	���6Ga�8��8�Z�D�f��z�:V�L�T�=�f�*�KZ셥����q�]X�� `�����Q��Nu�Y�j������DX-�g��&��?E.�_W�蕹��j�HP�@�Xț�W.\Zx��̚0xn�VW�h/�����z�^�'�`�M���	���*e��N.5���|�i,�������N�]ph���;G�k� 7�1y�����1��9�O҃q����m����*�����*rӘG�9���#�������h�ߊ�N#�\�WPG���f=���H��qg����!��y��t��V�FƮ�p�g��M�D�lJ���+T�h�ޢ�Թ�}?ԉ�گ�YV��"��g
�X����m�o�/=���p/~<q@�31�`��2A5�)��R�X�![%����Ӣ��&����n�;Kd�&����@v�&{�s��P�׳�C;��m
d�.�؉?ŗl_X!m�Ջ�S�x�GRK�l98Ni���VxޭD�cS��<LSⴘԽo���+E���<�&����O"
�vl�7Ա�1��F�<+]Y�_��>�x��q��1�%M���$���/������^��Q���~NW-����%;�q���l-7Gh���Ʉ�9W��%�\i����%
74o���V�ϓ�X�7e�R?��F�������-G.�"���bAW�j�³Dո�I���8A�=�uX@�Su�*��Pʂ���ͽ	�7�Skhb��|���&Iĳ�ʛADB��߹t"S d"D]_��3"�w/jқ��y!�M;[Qi
� �͙�a\��x����+lJ�t�[Ƚ4����*�6W�V�&��vV�BxE��.#�ܹ%'�ON�&�{���!7��J�eo

�bv�}��e�F�9�_:7D��B�ۋ���4B�$4ym�a��{��t�87��X�!'��� ��Uq&�zV��W���}r��>]B܉}�aˎ040��(:'Wq�`�+3*��"s��	���n�Z�B#G���	q>`p��~af��Ǔ"��
�.y8�)���X��3nw(w=ٴ�9w�������=�\Фaa��Q�R�v�얅ό�sg��4�x`��Y��m^�*��F��_��Ļp��a)���l8�����d*�t��]�yE�:���ʠ���$��2����^#�ԓ��������8�k���K�`����Z�*���@�3�}_A��#`.�������#[���X��愋��4S��r�?P8Ն��Hcy�gc���
�͉�{�tЀ9,�'j��d�r'd�������j'���Y�Y�֟*0x�X��d�Q)�	������րꤥ��9��>�1���1@X�F�Pr�!S�;�߯�Ե��{j�_0�;�W�L�e��1(�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�t��y�[��Gϊ��1�H(w���-xk?O�"��d�\�SϤ�犂�c�'T��%�S�PC�Į
��i��	e(:�Cc�4I�.�o&﷡mw�&���HHJ9�����֧~�(�\��w/�K`�n�����zκf�.��*�P��`���Y���X�rӊ�����=h����lts Bѧ�)�
T:-���0��3E��G;u>��}
�~΀&v�c���U�Fޅ�(�M�8S�HҢ9���6l��
�:��b���ߗ]k6:��*<�
���
y��)���b����)���p�3���c+B7 h�����|�b��� �w�p�R^�j5�pL�8�%ec sl�	���r���}$b��	`�ڸ&�uq2�<���exi\r��7'�{*:��'�9u�cUS��Y}������«|\L�>���8t�ǖ�'.�UXaT�p<�d�V��X�#�&s,����u�m�������U\đB���4p�<��k�1g!�c{IW�/��	(�tj.�4��R�����^��/�6�quZ��W�-��1�ƫ��XG���V�]{�_r\G���)#��u�,�L�0-p�\��q�ۆ���B�Pi<^tA�m�jʾQ�-gc� t������Ś��~h�tf���&Jil��m��������ǲg���g�!:R���\�����D��E0Wo�v@�S秹�MD��]�c��B�@�dM0�`\F-� ��3���x�<H��r�	��рȊ˳�[Rp��_7���c�N�����yЊ�\#�z��S�}3
�Z�����=�t��f��7��!sn��842�Ja�Ǻ��7\�X1�-7��u���C�7$<��X��o:�!�.���Q��U+��E6�Zb-�l.h_���l��B�ߓ��&��dBt���I�YWb�U�@9��ߒ� '>E��*ߠn4S��z��+~�b�����E�e'd�uKS�)�:�c~�6��~�.k̉d�B!�PN<�����r�jı���[���H���7�ft1��%X(�f�ǔX��l�j�vy9t~'x+O􊣖t�����%ݒ��=J(���ek>Q��IRI���Tsq�[[����uCU���TȜ���,��)��\4�x��rͯ!��?�W�,W# ��� 5��r+��W��eY��%��&��ǡ�PI%�g`Y��1^B9�N�3��p��v3#J�]���BJ�lk���/7D��@���䈊x�M]d8F�v�c?ZF�����y �_jRw�'r���8 f�`��$�jM�!Eʷ��Υt%�)1����[���1��ao8���<LI��w�\��s��ݬ4UEdKS���� �*e��9�8�a��'6�P�����c�2�.�fAߍI����ET\B<0*�������}�~��]�5����x�dD	cG�!�8�{@*kN|?�®S��硽]�X�?���Q��{���P��\��D��[y��c/��ٝ�L�b�#�ɓ	i��56W��5�-\ ��WGw����b��m�<���ID#�8�F�<$���opW��׶�Bz�/�v��$(r���Q��"�$]䲽��8�P��\/��bQC����3�Q1xV�������C����	^V~ �E"Q�u���o^���̋�r�/q�0��Q��tl� G,U�*ި���&�I�&Ht
�Y��$Z��|;��$U���$�ι&�0�(Z��4����AxH�O`�	EޠR�I�w�� ��Y6m�7�)d��V��Z9p���ӣ�����Պɤ�F|lDt��"��B��l�CN�7�WiWi͛���ϬL�Qcd2�^o]�b�d�'2�X��rӯst8]��ŋ�άCU5��Q�x��F8`�ĵ؂���!�x[���20��r���@��S���8/�V0�����2S���ڭ�z�?2!�����>�F4S�U�TG�dg~�0�ۮ#'z^J�����^�Ť"4�ڲ�vq�|�ܼ-�:�������'γR��5��I���O�+_N���/ɧ���6�I����/ �H��ڪ�ldG��N�'���GD���8���xJ䴿i})9����D�~�7��	*¥��Pj.�<0w�|���1�/��mC�Abp�`�%����	Z�j2�N��YŚo��7��3 ��HR
�ׄ��a0����y�4Z����6}���r����a`5�-�7	���v��]���VD��"Z/ꞾC.M�4��x�a5ET����I������TD�M����j�R��*�IK��t{b,��epԕʱt$G�U��٫���GD�Rb�M$�*���G���!&( t
�T?��A����O�e����,W=e����h���ݨ��/'�"���q}u�O��
AY> �-!(EI���f�*5̓��*�����P˴Oſ(��*�N+���h[hy�C9�����Г��J~�1x;��g����р��%�V��
:�R��[BVxUF82�z��_CK8v!���Ŀ����C^��2>ɑ�k=K�3����d���������M�[����m��NKԎ������A���m���h굛[Hű��xv�y���O��Fy�'������8u���q��F-Vߨu���/h����[؈��x9�n�+�ɉ�w"�/��{,��d��\���R��K�|��Q�!oم��.=���8s�!u����бi�c5�}Q6�h�
`k�ݫ�ܵW݊A5D��t3P�k��4GrâK0����Ÿ_C?�����+m����Ŵ�qW��bTdc��~L��:�W����OgFS�fج��ž�D7���b�M$*�(lW�.Ì���>����t,�bO��c�e}h�!�o|=`�����:��Ma�H�To'Əo�}/r������ _ο�
Ћ���?�2ZjP�{�/��7eh��'������ܯP��;--�e���o%��;p�ýJ"�F�0p��؇�O�ej�%�1q!�!
�}�{24bv툱���$��'�+�ec�Wdƌ��o������tNx�����S	�R����}�%�?�҂g~C5Bc��<��o�h�SZfo�2�JŊ��,� y�iu�䋨���7׼얄@A%�H$e��� �Z@��h2���W��A�y$@`�
˾��C���*`H�M�~�*�sKk�(��\��S3�$�Wz�Ģ
��)v�	��Ϭ���zc�׋����r�G�8dkm؁���Z/hG,��%?C<b�`�����}LDlD��5��;��C�bM<��[��A�����XZ�H_��\�8���Jg��U�Z��F��:�ZP�Nz-8�����sJ$鹕�!�I灓���Ρ(>����f�83������&��u����GT�k��b���H��}�����J��jNB'�Q��h��P@��@��'�W#��ӵo"�:�^���~�}W��������/&p�6������T5�U�<.1� |�'�}�-�i�p<LǺw�|�>q�e3S���<�r�8��k�g���ŀ����f]��]@��2o�*|15G���p����i�g���i��na�>��_[2���� W2ENX�X~l L�e�S�B�KrY�	��)�?8�|� �\�k�{$k �e�����u��%j*���i���I�J���	U7�%�Fc��;(։c���\�&��󔨱�[�~8�����ۏ��vs���'�%��oE'�`�c��t���K;E��+m�׫�Xʟ�Fx;���4P�f�l�>��='�Q�c��k2��+��c�/��G2@]�~rZ{�m�FOX}�*Eu:U\��.��Q�.8icN	���Y��|����R+f��CxnʍL�["������r��a+�Z����TD8��Lk���~��P����>�� ��:7\��� �4��G���`�B<��m��W.�Q�\��c0}�"�bHO�1��Y%�ɫA��E	�Y�%D��;��"���9��)�S�r��ֺ�Sm~�J�����c-_�k�G�m���T���{�E��z�z�ё�)�ӡ^m�r�$t���)�L�A,a��{��y`:�
b�y/H�ih�o�O�!u���A5qv��F�.�%y�Wi����|k:��_�ܿR�f������LIx�hD�)���4�sQBo@��揠S�<<A���$�a��ۢ���O��g-�Jf����#55��%�l���������~Lg�VP}��^j^�~�&8F:����i���3����>��_R�L]��3�z���H(���8P�m'��Z�����c�a�ܬ�9����"Ʈ�b:���B����>�Y���DW��� (!���}��@V�rxb (o�r�tRy�NZBͳ.j���Ce[��e�՜y��������jݭ��$�q��u%��h�ژ�_'$�����L1�^��. �O|�l�ޡ�<3�Q�l�5�傸���){�$\H��۵c��i�;N��6�9u����8�y���V�?ێx8�2��#o��MS�É�-�Z�?W�"�J3���=c�U���V3�|p�IWN6�%[:�������$�w�Ƒ�t���T؝I�6�k.CF�y�]�+�M%^��95)���oV{&�d����KQ6
#�6q���o��S����|�c_�G��l�Mb�p��A�mQ�'��o��׀�$�H��sj��:8���a�N�9pJ!�d�eAB���9���v�/2�pȿ��\�Y�o��&�l�d�
��0�Z��]����#��v�E  UƷ�7*�+�a}��)��Z�aaP�Ag����Q�()�����%�ޖ�'�x�ّA��ti�\{|���v㵮h�Oa��i9���]��9�yZz�z��~���Pد�>�M�p���>|4��#����Ї�����,�ۤGߏ��pO'w��t��	3�?"�t�tr$�"Ӹ�����Q��4_!�l'�7��6L��0>!�D6{o��<�X�����`&������c�{�#��7���������� ��I.��H�Q���`����
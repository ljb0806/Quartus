-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DI1JVVQFMywncNV6zE0cIOwr9uvV/1jJvkXsJRSNHrIXi0vLb5Rxa9crxVMmQoCibqefNn9U+xJd
yXwtOD+MSet2fchX7uYEGiCLMQyKHdz8THykwNUjUwLOVPAnGyRs+UeUDiNtxJeq52uzUXhdw/4V
NhCEJxBFB+r370yM0B2MTAyZuNEPXw5lyZZ+Q+baeYjFPN5xbq/V1Irk68TgrjfELPyjEjwOnxYl
iTRmfP5SsP5N8sph9Wkr7l4Wuip80AydUKYpnEx8VNk0UB1j6KpT2DVmgcd2zmmuiFRFFOoDmO+/
gHyB5U1t8R5ZbOY3oce+0cUDuo5koUWjiVCeeQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 90624)
`protect data_block
eIm9Ldj0rlIhNBwoO0OIa2wM+eYxfl+9aqD49fUwGUBUt8u7/lV5e/WiuCWgsv2hi7byo+duyyAk
NW3ntfHVUBinNjxbhnP4ShduaHFIhetuPu+M/rqdivWwUyVV7M/MMXuLARy3Hf7FIZGFGNPoS7Nq
adWznpawkENqEIMQlXGziF30bpxbwVlV23InczuIH7rov7/YxP3WSZyKjj0bT8BrVygj9tNupGse
sQ5LsTi27cb9PN24J+1vDM5w/8cV9+hcFo5IT/pJDRIHt7kvPJt1qLbmQQUu/W22pv7ENozxbqQ2
Ny4iESxUB7H0zQm8MMeIrc66NwWHFCmLvzHZEkl/XEGckYmKcjh9IAN0OhYPC3SIkiaSb9PBuOBC
8jIJq3rNzvvENYuCTjTSNZ7pL1Y0rkkiTNs64koCEfgSYlx6yoY6FpMhCKJwqJBsfwBAAM3kyuRD
ySHSdIGXsTUTE1knKEhbv0lPpjWLXwg/CvyZvuohu+hhjhkiKOkozFP713bZIDZhiNe/seo+dqWl
hT3HTAQtKT/2awIv/k5FsneC8i9cy50N18GV3YDwGL5XFmhynqlqfCAgBc+zz0aK0SZcrU2a9dsX
dIkVuy9wiruNX/Jb4XY6fui84ZYxAyH6MDEB5uc6GbtWW1PJ1vgUnFLBcKbKjzUDz5B0eC2S2V8C
mLKNMoUrpV1AVNkwZSr64FHKLxEVxPFjkBSS978OoXQ52tOmo3wnubihNhC/Ffp0brs+ELSu7IIq
f4xEWvaiY9tXeUYKclBi2MZ3mbYA/dZzj7GKpg1YTqi5fiOEjZwy85xTPFMoHABnsIbL0rVIJ5bu
3xLWdV8Xm4biG0wgG9tu2iZ524A1KSvE6+3gGJW5vtTHXBSTmenO5V8Xgfpy6VloeUaXvy4UlutZ
VP/SkEKtBb3tvK84aPu3X0mgnlDhs/i6eRRV87huu8YzjsyTEWKKcrgzTDwO6k6OuRgov24tYuo3
q85bmIX8D5gWZFpHX618WSysxDhnWwpbkmnv93xPz1YdckFZj6icPBExmhYnZUeK8Qg25WYIjG0z
usLP6XsM8SK9uohO4zEm2pZQL6XhATX20n6wh9qQMzB8eQ+N0JBWUjehr2Xa4X3nncNJPmCXOtpG
nM15n+VXwO0M24pSmoGdfzkL5FzsiBNPKPCykz9vNW3M3EBSx4Eg68q2fXmkinEU6zYCdDi/PFKC
qhaDChzVri8qKWgD9xZ/RhXpyPTm4TeTjOqJXmaR65DHuRVp1AVVUmorPFbrFxXsuAAvMqvLF7a8
EqlquXeMaqLxFgNQugsxqi4O8J5Kwa/kNLABUxTiapr75fYZpdTgIg81zZOsPVQDBUZXLveen94z
+/SbQ74WxZCB0BefunD9uztZIUADpkov31QP3yrBo3OfXOBmOOnVUvnPqJw3p0GMcREiiFIY9HFH
ne1NUL5E9t5XcZ9DC1HD7o0efIbPc1UUa5MztnUPuf2EpMxnhU9hvg+5pj9ky7Ty7SFbMt8euz4y
LX4kW/vis7ZeMwku+wi4Pol+6eTl6FMo2Sz/hn8paa3+DFedZqFho2QaFXVqNNdJDLkc3aEixHwe
iYvK6KX5TgCvkT6oE0i2Dqx5b7ILvlZQundpuX2WZasY1D+9kmQvSV7CJJw6e4vgjrSVhjmZaX6W
Zk/6Y/e2bOmmOv0Fz01V9K1O2Pxp2GKJbC+pxIRO7eyCVsWwTlNjegML/Vn/5EEBO2J9eJdRVqEj
Wf1M9A5cK7z7suycTHiGG51s5GInxew1D4pW8Eim4D7iPnbewuHaRESbn8U/12Rj7KspRbYlxYOU
USyuL8jRS+Jyjyq/FwXWusdmNjxwCewtYBJEb8nUK7RczLuze2dMOA/8BdC1SmtOy14O3uZodJGP
uvQ10TlXWUfjFqYT1jrVZ8lKBj3/xOZ2LkRMQtoM8YZfMbDXomWDUCAs/TR1nMpINIXfOccc4XnR
NWCETsb+BdiZI4YcHAJ/e838ZVKwWeZHezfLUBqSWQaYqsDQu3IvmTRxx/ITLZ+ziQ1TybSukWx0
2NkukTFpRYJPzdfSN13uwe6QFRkxNj1p54R3s52zF09kk32DTp5XMpG4tXDAg0TGG16oSL0MJxjX
nsRs49ZxjIrddPM2sNkfSU5+sPTxP2AZEZyoLw6GRTDLrSFRlo45pFyPFUgi2fnMq0tCVn2PWbjl
4YoQ1tiEWLLr/hsYzaokyxyTcfbq9k1XSRYHReY8wWvV6Vh6W7A8g/bHndJmm0gkiqrYvpOcaulN
GyG5nuOqJd25I16//ZOysjlRdLeFrxQjGYixM4GxLbSLQrtQZUNXpu2YO63nchrI7EnqY7fVniIR
iBCvE/5VGVgj1zIx8PQKlT5TEEyEsTlAqGAXFww90RkJeTVRuzRmYZBDqZA9er0v5j/ncwYbBlez
TZxFal0yKBQbWkEmgDF8L/5brkT1M7ZGMc+xoI/jTTwtTsicP2UeoTzC3260YhTpbcGJQ6hCUHgf
C4wY0qM/CsiGBL6z8phmw2DI5dJSI3Cct+2p72SjYhJ1MK38GLV7djEnevUquiYdiqNi7Viri5zp
StW72tnSeQaxkp238OJCbe/GGT9Ben+3doEQcsqWeEihh01F+ovaTzcbsoR6Ord13FdpjwpnODQi
bAbxDzK9jSDmoN9o/uKRFw9z7c1cN8OisheGm6gQPFPjofTMIO2Fmr/cJJC79uPYKGlAz+W5m+3q
Bw3sMxrgO6pAlHHFzdb/XVhAcKgJMs7sKwh8DCv4sug76jugkprRiYM2p/FYB76vc4LDIfOwlMLC
xzZTy6IkzyJchYDZly7S1yudhWkeapYJT6r60sYvlsj49aVT76P2H1ybBZW96Nn7MrnV7S5k7HGt
ADo313KbI4PfPttTykMP+T/alPN6+5jf7NNhh/kOrZ6Mw0iGQgRPFC5XfnKwxgedciH4uwRWntIm
qUf3Opi4anz/GXyMmZIeBrvJDRAxWDy+xKrb4olMdEvnoqgnfCVLwtYQhM48mQemJSzXLq6BF6QD
tlkQ0xcR6fMRFy9aJfgNgaxenUItUcRs5cfs3ZYPEONQFQLnM4gBW/MkXU2b/mpO8wLHEo9jQiCz
abHubl7UBn4pF3dWTWopHbf70L/brBTKuhhpuxUKTcl9feD4/80RbWAuxR4T7BciaUrmuZEA2MWt
FlQfkPNymeemmWxpxsvMsVm4cICY8QwT1bK1ttxL2taBmD7SvoyWC/kcw/0EPPSgPz5sV0w7f7y/
SXRWv1kMappgwash6hK9S9h2hCOrno3FYkhyHwyfZH3B9WvGYADRRBERnY4r0u4DbOpQw8ltRa0v
Ot/zePz+mV8/b51m7iQDqtmszd9jPqKJYv6hWWM85FdL/Bs7gARtUguTElwwUgfDV0oP81CaCPwU
HEhQJdEe7XJQ+ZWcBtyDE7RDz89byG8Zo3nKwUOXU46K38tjC8yYPZhuzSFPk3Po9eyIgSelVbPQ
noXQqF4k1fSn3kFROztJCoup+JJpbixk/kjISQQSC+OVFnBArogJtlb/8T7J1jzhLzp61rMCWt8y
FiZatGBOgybh+v4SOBOzq8wFPELmUQKImwrgFjHkoQdHhBHwMskIQAKNYLvDALgHcQoWisa2H2X2
csmXcLl7lcsKvtEohCeGSKsk4rYIxKJxhdlSfU+yrY8WAl11M2TsYJcTFWP11PLbE0RiT9CFB84A
HTElKzBbNkE00y8YbFp5j2QL+C3vDnNrvU1bx6MpIDQpLVQoILlJRFE1iz53ujAoFVlWXIAnEIAb
83nfBFNLeRiXDaPl3rg3mu3Zzo8EoZK1r9YK3rgLaIDOuPvoH1fzDzMHSz63YjInr6OXlfaz71+d
L6UZA2LsKe6T8pGtJIUBf8MIKyKv3nwapQmZ60r+BN7h4zafhhncDSo+TOq3i96uwiz7RSYVbbwS
PfLC3jvhJG/wiDIYne5+oGhTHhsWib4u3bxXwPtPZooNy4H9bAry0FTnlxvBQjo5laWjcBjivi1p
w5EEJHmieJsufEHBEdYBR4gH+CA+wYPCbGd0D72OjvDvvlc6r05zQa0xWwd5Iuow3q5WSnQJtpc8
TEfST+LWnr0J2AMu2N91dy7JZjo0pSNzq8wRHCC5QZ3aKVr/2gI+yVDNOsavEKT7E4QyVRuH1+8y
FDEtmQBGvu9u/zvApVkgGPCKO/WHFV5BvhH+Aj1HCzUcp6qmkCsJKvScdij5tQYtPdnxmiGjWv24
zcEUjLuEC44DhOcZdU95O4hHmePBUUf2VoYG6AdJEbmiPq8VOW6ooU2s94A0VxgASLSiVPcHBHFn
wfh1WpXmBGEyJm/hK2UgWjZqJiMugvzoxlmPpypl7YFTIIpQFKgTWuleQpTAbdnEfhfdwjVoghw1
mlELD0QxwsBx1I8bRBn3jcon+z8isccnI/yxuqVLj/OdJlNVg+N5XY8RokYCTXzIdxOy3jZQVHaD
U73/sDFuMYCgnH7IijIznvvbWyABTqZQcvhrSGfzx25H0EW4IyAJm27oKBogqbyy6voKkiRTvrSr
Ril5aBYthoLt7pg68mWdJEHWDPkGhKRsM5X18l1Fuc0kNIGzC+T1+ZoK9BNRTh3yNSq4tGLzsByl
ftIWvTYHPS5hPkoghc3TGLQDK8xw/bGkcEhZJr8LOk+RWEkA2DHdbaKc95HWgreJNT1IYORf8Ua+
fs2Gs4ZMPrOZbNEMHUjiYcqwB5iJCuQ/SPqR2K9RZ6O99ah2ZUBN2MoNeyi2EDyN1V67dogNCo2t
XzAZHc/BDKYjjYmOYkn9nJw+cZPZBz6VGGt/lJNqsVfRzGDnSMidC5W1JN2jRSyDKYtybF0u9OUo
W18VExyjAKuibuGDgS68Ze3hVlmAnR1PrruYDqtWaL9UF122dyVI+J3YdLkntpXvyhcZx8DLOdh+
61R1yGyAZ/WPAe7G6WvvpB/tDNQtvlQfyvCYjdXKQqkkmQScmBW/z50glVxYhW7W48KnXaYORnm9
I0cx1ZwlRM7nPVn4Lt39RYD6691Jm062cVb91ISFjvJYykIZLNrv++f9yDnlwlOkQy/BIHRQHHip
HR8Iz1yAFam8Q7Zm/FvJHmC2UalyGP3VOdHO00UzFG5IEpSB9pZZVrSohQWKIOr7TTKy1sVIXXa0
gX4K+v/cX2S5zpIoDuBpbF65fQ/AsoeAMSd6yaGKRMBP3j7hvAd5rFlOp6waj1SVsdCNyZCfVxfR
nDoCazQvkOMNkS2VMHFXNUr2TVFEYQFS49nEzFkK0a3xTZS9R5MMQeCGOCcuKiK6Ui5k18Y0+cZF
BPBQUmcMo2XBNdw/50j6x5ncVKdJ2/PSpD2KmUALPJqFUHmHNiV+ux9tF0RWOuDpjwX17C1X5+Vf
DysY2udJ0WWjDo3iO5KjzCegscDo8w80STtWblU00SAa5KznPr6+y9ctbJ5pcOKDOKJkMsJi17tl
0FkxAxsBjCyXkUR9aY4Rg7dv/2n6hEmBIrhXNyJTVcXqj3Zw+nqH/kQj0kBnfvuoLLTsieRdeSlh
D7jQJuPgvjTPNctVhkmEVolL6QxVmGdfNgaXVJaydsu9CCMTaEiA09ssIyqyX3+FzLCCjgjNUY9S
eKwVnJppTFam83U/uC37MLrNlZevvfwygc0ox2rfeRnEbVvkXrZbnMZowHWA/XLKP4UvRAcSQpSu
VyIdWn6WVZU87yPZIsrsDXY++WCNK6GH2LleB6krn2kqDrzx6VaMj7IkGP9ws4aoU0o4P9DYkIRd
yz7G3222K+abndMDAPsdXI8Gbt+YiU+eSW58dCvphlmVruNjUpkDbQRiXicyYgjPaK/JCeZTH3U3
/z1SujAt2tjpuEcVu1IpHCMCbRMJalsygmeAC/M4vM2fZBuTfGiSPq3VGs0qMmZsiz2EORIM+98R
zc5SmeW3oboeux1FBCkA3ox3wFiPMVEv/mH8k7RMW99M5IPxwPl7jnnXna+5mVRU0vsUN52sZfSV
iPbXeDziHfA4UJ+znQ1JQVOw5596BwHf15krux/cGjCJCUVgDxRb6mvfNft4HavWJrSy2N8hQV66
3LZD269f7n5PSIJ4pfsWclqhtAuhOWhvwzr05upufAmgsydd51JAXiSZiKLazHX8k/VoOwtiPZdC
nxC3uIl8VYxFgoqRCE/3OPljHw8sDD2vs8KGKT+fQFzdLVHGsypVGH+4pZ77vLCLgKzyKV83B+S6
XKFD5WvJGgzzcWth8ne0/vYWYSJ4RxTovYotalGSvTZAIAkc9Ov9pgbOIwak0Y6zZ+LYj6VqeLNb
b7awVL04p6FjiA01D4klJS8b8G9ytL5F2SlwY2AlHDzcUUYRdfkCSuhmF5x7GY4c/Fiv+1hcEv8s
dYu31okt0JhZ+Ekcw1mOlD+ncMJumqaDOtBi4t1mVJysk4K9nnEI244oV2WwanbImnHfH6DF4sQ2
TRhGKoyVevQtw7U1e6o2bYLLcPaO6p5p5JOMgV5R9p/GQjAfS72jgqVpTvnxq5DXvhEKagpAW4PA
yjaGyug4sKpVql/LjZ5e+nrssi127D54Zr1fw2r5wxXZfnSTPkpolpNiG654QrjEHlsZZfZET+VD
1TomYkAaaUSHq/GLPvsFt4BXKKuuOr6sjp5SFHodvazvfwkHObeGicykwsw2eycQPgCcBV9ahbjk
XwratCVBLG88iV6e8g8ZRvQvLGRTG8XcR8MzWfiIIm6zkh9L//otH9OE/krJjVyGZEFJhROOxLQX
dwgsaV4xDkHMZ4MtFQgTmvICxXQ0e5WW4WxXiFRLA/X7CqQcfMfu5WAmpZzrwY0omX+Z4YxmHDWg
mtn+3aMrYph4wqaOpMRwLhxpafaPTxo1BNeb3wbJbnFazpYt1LSL5bYpFLMpVbdubTj0x3DQZ0n2
wdN1L3AU0BzjPNZMkT2kj7ki3XWTb5seTv8LCydhl2wj1/gXEPJ+Es8IvRgHRaOhqhgssFD69aZM
T8ArqLsKE7Igp9haT5lLK/s20sphIeem/r3ZZAMHrD8nIVazT1dbDhbFYRcqqSZQ3/zh+88L4nMV
wqAy3vVKj7oC3plnt0l3e9Qub8h2o/L3hMMdr+zQda4aSc1H//cZNfsHHyt9O9IuveKER51ZJho8
dFnNcyvI89OsQ0JAn5fl4oQe6jLRPrhboMwZkbJW61ElBssa9tIARyAqtIY5VPKa1ypHtO4cC6cy
06If56tG9JqspZ8xolYI46Yt2ly0YjYJbu5esm80JG7x0GYgABI6f8RA4JV860udKCl+K0cjX+II
ioN0xKHlvADVTP0HH1PcWQzd8aZwgMbTRqMKRH2kb68F9wJaLNZilDoz9VYaArM6YJajP3ElbBcL
M8c2AfAqGKomip1qj5r+WXH5bXYZlsfJBR7sdT0hDutgmnSqYYvbnWjW9ymGQi5N34orcV0vOF6+
UrYY2rgTdcWDc6zwutQG9M+o4jgT1URVdRd/vrDx2gvqbhhMeiRnsg1mjzzRmdqVnKif3lIrPOWn
cnPgPGjP7vbMg/5F/2gD1fOdbeNZ3Ky3hdeanFJsyBJok3g6Z+XhfvU/stxfRKLPUgJqf4X00Ywt
B+X534cRT15gE+td9jtNwV0358nZFr5L+zJJiJbBrJonEy7eXXU5w08kGIx0GOBPMS5ur52JkH1Q
UfwKqXLgzam1g1GRqE5Do0fPSUdFd0wzSiKG0oQVUVvtPLjz02ZCwB0askkYid62TLclXkNwKzNd
uxXULyBf6dWFIZjfOINo1utJZNnpjkIJG/RO0jjqKykrcaP2IG5b/0+GXSRkae9FzygC87GY/UZf
LhA5wGylnlo4VImnKj98rbeFKVeAkAkqDAizIv68Urq6/hsP3eKSfPaJl/XyKxlmgMFa+TZPD1mE
jW7G9z3huRp9BagZn+CMdyDROI6NfHiL/vb6u0eFmGJvCRnMqOF2Set6EeYpcAvuw4D81+JouDo8
8jVtQJgbD/tI2m397VaHrL21QZSctsg4c9Cf61iPQs6gU7GXju/txRgEBDlmtEmR8tuglCDMVxsX
RT1GIgnpjd10TrD2/TylfqT1bxtx7wRdxTrm8mLanfkfpYj5UMim/I/THRyhkt9Oo5uyz4HU0sWV
uF0l3Gkixy7zMCLMg5jbNNqd1Dot0UP8yHVZw2IQAfeS2eg3BnLdFMvZiVHLfT8dtCQWpgwa4qOI
N5hPmI3GwZR2zcGW9f7yhYYdE2LRz/CtLQblKmXEK9gt3l6UpXHpz8GOMlCDDuRAyG73253dklVw
N77EUz8DuEKBcY30Tj62WOwEN0A//C8/UCWyvWOEcQl+5p4/NGHiHCSVYDZocpGSkpt+XQWKmdBO
CT2WDiJb8ckPHJ8h/Tf7VenyI86iYeKNU/8G1Eolk5Otkj8MJw9SA0fVAD76TjmmyZiCb7P2sSKw
l4QnAqc25L1VhIxAJ+VOPS2dJ+pK4r6d0Gq4HN94iMQjFgl0McmBIgJ5f/bqApfSfecn3NbH7ppH
33Nq0muFiKUewcN3rGBK7ahtJl7rwt+YKu1HIi0U5pVL9N5rQfSMmSz8cvmHIhyBdFrFj3x/0KMZ
yUFVEVWyRpDhcYxyk3VEwJ/lqIJQrTlNvSXRDrBBQGegEebG4Ue8ALlBL4JlKqgyNa4ErV6QJ7Y7
0+W3Oao69w0eSAPpXnNKdJ7SdtlFxxB9KNATrAkHxSSqJPrPo9cTPy52MSRIRIyCL3xIhBYjf1Ip
NOSMRb4i1OQVMpXqln55nZbX1umS9yHEC/r5hRps180crjujqoXADmm745Sk9HgsEn8iVdjLgohO
DDYkPMBKuPtpczKqRUzX4seT3HgdeqxMnSA0GbETDlO5lZ5F5FXkhibjMkxXweESoP1FJO28gqXQ
auPNV613VePe0Vd18nLDuUo9TOX1nR8bCQ+ptjg5rMcSRMFXspbaN+b00WbXw3sgUpNkFtunAdFm
ZIAOUW6x/sMK50asc9NXf3A1k899Xjj9OB3nXWA6hCVTCe0r2PSmDVg71rX1KRdCvXnRiZLRWpue
2O56L7U0MiggA5ANxz3gz1l/IoF2tMehe2B24UdMgJwGLwoebnjv0oWwEksuAgH2Ep031Z+AJ7Fd
r0w/Kkih09qB/YHJeGFCdPQ7BTO10+Ezw/kHni10xtrj5Gs8DTLoW6h4N5FaP/P61YCpyQJ5eMZK
DCZ3L5G0wqLJcoLO+wGeE05KDaFbOFjloMHH2D+iuDuWCBfYBpnRCqajK6E0ion1Owx4lUZc3LcP
Uhm9KKBEvo+zjjpZ/bM/S5b/qGVzZzeEBfMpxuiNusKrMVfGtOuH86TuTENfTYOR4zyXXW3XLTtP
BNe80oT1GWOUAoAaSkBl62Cy6fWaCrKo/3t8zW7eXxc0P+7r8OTsSG7ZY2M9uhKJIOP8i9LrXiCg
+jYExM2m2yYcv4z+jUTJjjdZbJfNdQnqruUT4yqaNhWgKHMqUO16wgD/xeWlWHw/pvQecyI93i6t
fvua30XERO0Ky4r7QGlUjFcg1P5F8SdB8xDt2ynJjf5OhpjjuFtA2AhEiPJuECEJnBExALxi+1he
QNvNOxhSQXxI/yxIORwSXKI7k2DzK+/kvskwNCGfFKxSBe2NbclgkXXHqkGD0NO1xG4TWLIEWUKD
l/ihIgLcpv85xjbaJHSF4IsbZDHmkklITtP/ojQI/5db54wt8mt2xe1NBSm1TzdBu8tTqYSQKOeL
JKxqvpHHRQLspuqt+N8J8qsH/lhLNCKB/C/XJidFLk5BMRw87Vtttjwr/M+nVTxSH5+HY4iZwhUQ
VXoIc+ygMIJqFcF/4UDBOQuu0hG2RyTPtSN2hMimpNQgl4PqRJWnYe+iVOeiH9rRGKjAOWZqk95G
wLQWoryAkipgKkZFfDVNf0OHJXj8VbNHndPg+PYzLesvJdrLhvRQ+Qov3O72zdGQGr8k9xn6VPbR
KUsyhcDjzGBPTCSDGlTRZjY1yWX0JhXcR1D5lhY0zKZJiUvOSxNumbrzhHQBgt9sma6pqP9dUGV6
QZyMpHXqhgxm1jGiBPq7v+GsT/spsvji0DuWkoK5rTpFkB6WXQ8TTLslr1Fz1bmQD6BJ8wRZgOaS
04wzj5ReRt0uFoZSg4eIY5Q0qY6OZzFFtXO0i8M1p4ZfqRM7cpodbTmHQ3ZHX6RMSg9UcyETYYMT
CcDDjXeZAbirCYGc+jOR0oM7o3gUahrM7cyA4pznc05wkFHzg3Ld/C9cwtI3bCUSaAr/VMCpHJ5u
DEgdZ2Qdi02xlNqaiGjF9KnOrBajsE437Llf0FMhlg75z2mE2nLE/I6MQiRxUp29lQpyMKoGDwkq
P5NpUAzPjbahVkaa37BgBiSGWrxgd1LUJoegLXwdbmBrdwdEZJHrxkvic+0i6Hil9F52LF+cMrOP
TWAla3jk+ZifCN0JJxD0JKFEwFKzHZxBbDjQeQ1lggx8TqNT4CQ1Ok5wnJK/kGveAli4OUbAx46a
iQgSvp0yY+qg0x0DwerRBMXeMsOou4ULjgJzoHTzUX2QRKoCaZsn1AbGZhK57s73r5XyriQKKlbn
uKoB9Sbx6BdJ+c3mauCX0KDYVmjZ++Z4AJujyaWXdwVk9RDXQN57644dGj7ak4t5oQfCvIYwJWzs
Ttr1AGjXaVpbtMLrOA0sQwbBn/71sP/+bHfs/F5YgdXK/yLXpSUSGk+qKTnwTMHp4V6eN51bTXXI
4GITwdBv0/+ccLulkHZUIhtS5D45ZMyxIJDRfxK8SqBD+tsIGXN6r39mJ/0uix9jGbYsh2qUVdFY
ZuTNuWEbKN5kjXKBZhE5FntHWScxcstGxIThKa+GUkbCPuWiOjjSyH1f4o0N0U4J+NzH4M1f5SKK
hqMgnfJgQHWbFglywEbEoYFVZESkqBg+DfvjezpXDVsxvsGquZhy1FixMdOA36gqVuvlsbGUFa6r
+J6YXAUOPBDWoP8OynU41oiUj1/5+0lgJmKBL89ogCNCa95jBQZ8z8GWjVaonmsaHsVFhd2NKArX
vuf88Gjk53AFiProsSc9jOxWKA3S7E6WVfzoh76PYtJ3yRQTOCJW+A074NjsxY57AhkSdL3naruG
/3jvQtANRp6hesHSS1vfgn94hdnyWKW/qY1ouvA0aPYhT9eUkhZc39HPSuTJMOo1z5hZ7qEsDugw
hndFTwiyScrF6F8FIONSssuy48iRSk1h0trGkz9CLbzbEel2SZP4hsh5u7utYCnGmxSAyENiWkUy
7WOGXQK6TR6Vr4f5odYwpsELrVM9LT98uUPktcxQx47MRAF/GPrUMEOOIvb8/H7bZ1WBa0gRU7mi
33C/HOLIpSWAuMn+eBSZRhCjBWBRuX568P38HxTYJz7rL9k0SBfSgGDTgbzviVFA5IPonEc7/6MK
Eg24LgLW3NVN7N3Mkiq0IsJz3G/XscFEROjHZH6V3or+AjbtpkQU3Gh1ZKKF1d51j9/k1fXmvpGQ
86zlVROanmh14pAcMyQN8WjcZRAn7z+yzsQAY0RxOC5418jHCUphps63xATDg578DEoTSvU3M3h5
/bi9faTY1w45Zpq9+1TXtDyYXOB8GFOEqhdx4BdNNLPHX+Xpp6Wr1KPAbIkZB9IAfjv4IKdKHnxc
nBaBdFIfWwdp29fuc2xPGvOEFJX4vzxRwFVSTE4pnZpTI/jTTEWmT42f0S3iP7wnX/ZxCHQ7XNa6
hGoyypJ4Y1EPoX5TfIyspe5saDcPBn/+aI56UO5xGtw2U4PZVu9bOjSuHoxDf9nMgv3eYsJAPqir
2pAbtJ7SmUye+8VPrXi9ywYI+NYZ494od7qLvHutNiZBO5NLo+4rTaPn/Hb5E7xIzSDnDQYaWJo+
0AerDZOFVJo98TzSyIJtuawlfZskKEMpvJgSRiDtIqvN+SitPvK597aL3AK4FI77z3r2m26XZ4Yu
brbpB4KUTnh2nZrjmepgLqkbu9Yh2q5A+62Yw4WefdtNI1OVnQbF6U886jmGXXzRpP9oZyrJ9KHS
ksty7KLTgsbNbe0qaaKUrzoXq4NNUuWAzZbe+ECIxxgLaA7WXRfJ+UDbDNudF0m1fcAgbmBQ26U2
7Yeorq2HIHZ4EH/TAI1bhFWg+GmUZtRoFKK4MKW0IFlndlzEOu7QiigdwQqeiiTkGrULQaiO17yX
P5x3Sxw5pqBmuC/ZoYFwG8UADMtkbxzscC5ViMWsveeAf70vYuoDmRP731EibHvFAuNeN6lKrS8/
3q635I17KyW06usrSjMB4CDi4cOTPrPR0EFl9lcVs5g24rhMbbglZ6S3OwAQZ2zGtWmP3hozKu4T
UHuEPD62dk/Bry4SnOeb/o8j6lUNPKFJN0+gOMDTVJY6nVWjZVJApAtiRQyL2KofMeAQOnwGZ1w9
JpDt3+Z50HrqbAwNnK2RBiXw8gSpsZLxhKH8NNYY7dEu3ERcgDL6kOv8FOeZ966WncRUjVGVulkC
1TJ0S6yPgrPszosVhre4xz9P4fn0YdPQ0Cpwp1dPWQDcHsEWtqDcP+0m0/d9xeO+v//x1IW5HcKq
usJ/vi2cld+sQitMYRfG4Ag/M/pjI/hVazD59+AXrow5yuI6BIcK5BS2K4m9MCLKkIHo6n++60gu
/IRsV/IxR7SEJtSUMFTHw9hUG/xER5iUDRQA+WsftsJGFrwBgTwoE4hd2z2U0s8t/AZrGNt452qG
4vPaOvb08HL2Wu7MRfG4c/XwsqabFyP/7T7eEXcF5cYNmPi9XSXzLN2dyq6X+Pfrr/eYw2IiYdn1
MMlfIm6Ov/mVGenc3QWQAZkfh4rLepvLrvKFMqkVXOuL+HT02EmDXTLYc5nAcMGebhDsVx/ghKNV
EgvJJ+8N18DMWFY3q3OQUHE2JPUm9EHQciuzlgA7P3LL6lzaSeR/c3zMwE27NW07FnAaIUWDX9YX
sLcBKgvq3YpReGhtc2+B95EK+EktG+6t1nbe+hujzluQqI4GJ3coPb2FFnBl8RqHq+W+C3aqlIJn
/ApqcwcCY7hedx+bvBPLxOSVBN90bU9p5B9x3xZuo13M0ynkitzqKVQ5zRfgyzUaEVjKdUT7l42P
Ziz3a4kV9RMcV/y9OPwihtNKdeIopNerv5c8RBIkGGDBbY6N8LW1ey70QcMHE/5gS9M0U+/qLR+p
nxbyPTb9Dhf+zqh5+oFcdlO2uRxll+APplbaCTlgfWbL3F1wwHPymsIq1Vr7o4hukCRPiZ8jy4+a
vKwXjpdoWBaW8yyVvwVbaVwIKIVRX4n7ExloTYcX94sBt0DC7vRq+/qoXdpyYZmFlGTRjQAh5oqw
l3CSzdbDjD26QoczN0qSpRPPlGxxlEGxFWMcYuMc8IStGHY8qHm0JyZNx0QmhKlZ1XQXgNSR6ZzL
AyZAhUEMvdKB6VqOpHNDaIPzUIrSLDtlQVpIm1HPvDXxakM0C+D2/8drX0HCXw+TzOnPVYFc53B8
k/hzvzS7+lWFHWzaxY1GNlqbLc9/UQcrvk2TMl9ew7cVJM2XpuaQn35P8mYLo08nocA9uIIE4Ly9
p0iNtwS+4c4EwC72NDh6mOoRUKvy6vGkER62kX95JWRtZZCy9FzwPDDwEqemZsb1Qm3OQde2Htls
RjtN2FO7+xMM1SFJYirzrqWOQ15AYKw1o1cQK368MYsSIrcSIxNd24/TB7YbHAEQQaZr7EP+cRXc
b/dvW+IBiy4h5zQu7GhAY5avmAxbyJ8DAYGTqE1T7QAODX+8vGI/SUH7M+ws2r5v3NzgVACkj+bo
r6cxO5ikDTnWVf6C01zomR2h0Xem+sMHOkjo0TZwuIhZkgu00kWaWoJUthI7xVwAr653lUXREFks
rj2h+BtyKItET8yVlLJkBPJh/tverwCFmIKn5/9R6imTqXRZGO8+lUWh1LaA9u5RZIPpoHNphKt4
bRQIb4fZxJub7WPqUkSxgzZUGevj03BHr9rUcq7qFUmXs6ENVv43EVGnTy6jX/gt4FkivxGQcF/i
0PBtI7o5+FubxFym0Pc8qocoZpL2QNkav+O4fpRgaElbSLEWxwshc+j5w/0Nq1GETIysg6+8DlKh
4KohrGHDhV1Dtw1A8/flwJ9Zs0q8Pd9DJDcMlcp6HjnJTXaw1QN6DEHiPclMjN6ROqjsX0/KZs0t
VPiCPQM9rJCRFtGwAyxszCAW3Y3KSEdWs8JrkEi86FmWJWb94Dmi2oJ0keZydxbvVQK2bq+XseQV
0zSX4xW37O2llbU0d7Ifs7th31OFoYgB7z39Nw3LzzMmjqorvWwAE7E2E7MXTWiTKDQOtvvKq+o4
/BPl6UE9d47J9xl0lrEpofryzNZTQZQQBM+88115bOLgC1m4kszKzHunXW6s2zP86LzBwvdLmzhb
mK9XTjNww8+QrNdEnnitukUvZuEWUjo9WJZJe3Yt0T2GLb3ct3D8EUguTrZh9df7yTK7BiWO54cI
Jyo+t8IEE3s3in4CPK1l4F6l2Jt2crSc7n26GQhnpruwRyxDOG4UPYvzJBUYx+IRfEY/OnfRRYgW
xcz6xGeZLCnKeP9c8a7ooCWIPqeS8zdZ1Bc1Y3vwh2SQ/anYMq83MgiA7XUbfeD/fwMAg931thHB
DfUaAmVfva1zbISPyf4alavae8Ye1yAx8zZwcI+lzYjNCAKyCuLKmHAzlUHu1Q0MAQNwhXCaW7tU
1Ev+w7Um908ChW5PfN/FMrhV+NxVU9hW4PhuQDnZ6ORABtZg9Qd+uBWIzfL03gjpX6i6t4R1wz5T
qzGbDjeKhciemWJDhNn9cXaQW7yzj4Vog+CKNEBLVkHAgckZpIJRx+VlZqUp5HXi9wVlbT+iv7Lg
Ag6iCz/C1FiSEIJf3ivrLVl+KfE3sUAa5kwhKgAc5lz+Cc8eRDfWreckinsVn3wjKFR0dU9XGdFz
U76E2HCDY4y1T27/Q3ULc3XAxaeDvV3jH3DCCI4gtiTTSl/GIDYJxMOXgqWg2jMcXRjktLHXhswg
6T2YKNZlAPEHbNSZHP8f+E58xqJ5BrMhWBx8LifDyd7gNMqIcinlvRhokZI24l/osUqAnJC4Ziau
hJXXqh4e1ldWVXJZ1Zgerhl2/Z5JdjDAp3vp6J6TTpJun4N+QCb0CyWf3vBBed2ZipTnL01qTNZj
0wtPRcQWxIKN+bJ9mcJ/4DGOmrgnkcEuAsRVoWfXKKCupGwfqcLmP0WNs7dqUI5IzuDYEtAB+M6A
Jf0XKfcb+dg69GKcgmmct68VvZ0NYhu3pYw2FwO2qthPqb6UAcOd7ft/v+O7NNi7en0UtVGuJcwW
J2wdaz8QBbj5RJnOnM4GqIxDCsmGu6R3J6p15mxhOgTuZQ3PsuTm8TtI5CdK9KnViG+n5p3o5289
adguse+b4U3oA6uApn2ckRl4ZYTqLebh5qEyZXKBhsHSbh/z6uHY+jC4zwHDPpaVrLJ0TDfWP1WD
ACktmlF5s32XUEXSvLE+tPJ/YohWen1rL4MzYorX9SZdetD4JHHbf4tLiq/rqoHadAZ5e5S64iFC
ZIpJxzG/lZJHim28e79pKGpRa7H9ZUWXmgU7vIUTKDJpCcwdqegH/8NeidWE2SldEa9DkmLtSjJj
/BjWTiXoHOq24Kc7bdvGFTF8Y93ZMJeF4keuGU+Dp/FVR/sGBodWDW0Nal4Vg73KJqb9xXEc3imu
b9iPiLRHBEiD7M3CgzTlGj8J/0yUR6j25ZYi3dJwyQaafpBQeRs0DOHbi5E+ceDjqfH0BP6Ofe3r
XtJUZo1W4n9OVJGTFuIyC1YcuwfK3NDnlOuxpmLK8sbwNl4vaiwhqBWzAcauHmdIq+ID0d9Hfwht
1HXv0pxITLbeHXIdb/Zx6IunGwI06QGPXLQpDLVg9FseQHINbwtBetofzZ1ajOuy4FLPGSm7OspW
Zv6Cq0OKqtNy2xrAO/6wFTDZH5Ip8QTXwXUImWQPg7ofWWjjNSkEKsFfU2dekRvoNMqjTFRzT91X
9KPmYt86vA2HRwpUA3cfFrUHX1TrBZbJwGP2RXZNPyd3HcjEB52mbPneYBXeWuzVo21ESRiilvWh
YxP15L3eANXIATUWA27IFRwr+0rmLCKmrdvCM6T2oEdz22KxtA4keZf7W96KpTRpOSI+5brZNaVy
TNPEERYScejrO9bisW5ymmFbSL4tuNIndbTh0KOJE27YRiBgV13vh0NfsjRty0IalDmnO78/lki4
h2evRPvze3qBVL37QONRMgibaEIrqiN9pmzT6KG6aydplLGf9CE5bRkDS+3LOl4NCzsxE8I+Iyri
hvfMi9gQ7+fKGqrSFwFhRSyY9w13ZXdemE491Zf0x48GtP0WDAOWZ+LT7maR0eaC8CaPamHJlvgg
f76laiygngOsra2x3TXydOGSh++xnJr/kkci9dltGfNKbdDZZbrIA1ctR8NG8jsFQ0iwv/iV6I/7
xfOV6gkjznSRGMsFdzz5qKx2L5qUvvUAzQQqjhyCIuvoSASKdbJyy3bSdTAQ/W/e5/BTL2s2o+/d
5fgnEMglNipEGMh0E4a1inWd23JjiyPhyrlNKdMkYqsaXyNZ7CEIZtPn+vTg6R2eawDrIZvCBmAV
En3IqTaY7rjmaIxyzKgJC6tO9/GuUep3DAz6WP+a5S0NuHkUSS3TdV2hnuAPu4cyp/v5duHhoH+m
MlVCjj5mYnUc1HM3xqwJMoyH6me0C11B5IppugqpLJuGbcmMZL11uYW0yAP6FZ9vtaciRgXlOc2D
RF3pW3ss24ZQcdsIBEm1QK5BLjszLde/LysTwIQOQfza2O9jTjYMCkvj9gNxsvsG4U1nEtP1EQ+6
KS0pZ4HXdbjE5RVqwq0ETtLFMVoVXXGYUN3fWqU7HOkx84Epc9CRW2g/XWa3A7NNt7HoAmIoO+Te
CZANIWcuudGprOvQL9roTbRHr139UJCcL6/dQyWI0MJNfcliQAemzdpjJM8gQTQyItYFuIUJDhjT
R3mMPrKurothov3awieyv/KEeCmU0LJwnEagrxKOV8LpPjef5WzjAc46lYRrs/Lcm3BbTWoBulhq
0NJJPg7QAHXci3z0DZz5uEVP+yS4AYPC5cdS+mfbn1yLbfQzHLy76P7+0cHIiP3XT4fWfpZ3bj9L
v58RVga6Un5fzoxSRPBcSwf4ZAhUJtWRwRItIFHGGDXPntxYn8ujvnP9UzMV8tBbZPrkYgkn940t
45xyca2tFzpJnbJWZOSo/5y2N40n0FncVyVj4ln02AnC20usfI5RBp2YZzl7s5X0sakFG916oVH7
yqUIBDkKDQTghBz+EKpR14TovXvWXkQB2WZ4nWNUpOAWZptcdL0OIrozb2eZHzwPenJExkm0ND8M
mG6J3YRvY/6MTZZZmDzIws1bRf+0FSj7foc490rjttTBDpQD3O2FdGAaknHVpI6oQn5galiKXZ/+
8V+JFPQIUB7lbGojrjA5yxCzLI8FjW+8qcogqus2/z8OHxeVJMYgFal5d975ikz5IYtVip//2N8c
7+E5+5HE0RN2TPdegZARXCsee3IvEnNY0oVfsotmUl80UGl9tX5r5My9AYTPy1cMXxPLjunLUoQE
kACxP2HCk4TSsfdISwsbpkojAKdGdeLbA5y3z9gfhrAXkCf7/KGD/p4xaT3E2yEvhL8YJc1pEXPF
Op3iL0+H5q9S+RMCN47vuB27PkC+nLtd+0PbGFO6U+cjh+E5Xon/ZYUWfjwlcPWvfXLrhsVBhVhJ
YJuFN7jh4PTsUc0Qcx8Rr97oMSFiEMq6wP2OcMtd6PGLDkOXHxlMZ1vWez/vkswIJKdCoU3fmQB9
la1Y12ZuhMItszaW7XUMx+Erp3S/kuPrQAtbeDBXOjqcOVGdKf6r0fKUFaPc1G09zt5M0dotiAB6
y8aQP8+o9wqAjeXfQdFg4ujkqPvpQqnJzIhK3CEq+CScCMLLNyu1SHpCE8dDqVrkqOriNEUmz5UF
c3OUhxYitKvWLwf0t6jFP/HMUofmtYcv7YX0wuM8q/oS34bWIXzQSxG03uT+OIh4Dmyd5ulPQvR3
iOnCFT0e6KEXstE8Y6MIWgWpU+kJjt6oZlEm0Dx4RbkZf/vpdOV//d+WMJSfqbYKTZL0flv5JD1U
BlM9un6bkf+uu92Ss62Lj+RcM9ptxbbmDmhWjjVrpm9mABUeTbselx4DoSU5pX1/L8tlnu+PpAh7
u9ev2DKG761d1mQ+E/F+2hyJlHlPXl4CLlUtnK2DQMGLvAKzPKguw88XtcuzbpNBGGPsq8WL82rO
qSrIthPSLyNT1sHwiJmmryZXSLyR/JVfUxDacM1wDKuF3bUrD4qzgbiRSf6mojhVnCM1rOzZ1lEV
bolNXHE3HOhO5JlJBXX1x6MQTMGERVXqCjaLKNPL9JfvbOS7/HzHyDRukwvzWPM4BGTuy/YMAEa/
OOf+eqTl+DLYUdDzl8BPU1x7L8DbSGQQnURK0dxbEQcFnCB9gIQASD+JPGut4giwSSSPPI7mHF1J
fV0dCRf5coIPmo3NUFIAXrPjfAS7IQU9CV52xa8GUi+zVZKGyyUe96WgmH1biJjLPnWEd6w1LMu3
Wyc8QSvtSmEi6/CqqmW+tfRf6JEpxAThECIhKcOZHcBXdhjQKUpI21HE8mhGbX1cM6k+Cdxb/JIy
PSHNQf7jJqonznPz37AVrIbHj/iHdLM4KzkKc2eu26zYo3jfoheURJ1//iLGc2xpSof1KOLfI97q
nCHuSJpAwrBP33uBowOk16O5Y7bIlDVQewTRAd2gZAzv+JSZZMzIZ60kdZd5oKTbxMSumSpyJ/6R
BYwPtbcXXCKmxSlOJSYiVyhrH3naoGLn2GNu7TVyRhPl5TY+sZLlzJrEby3nUNf4hVrbxWzx5ZNx
2NUy7XBgIt5XQUKfRMwpNPrboPKX3mDk1qmZaAJQ9M5/HbP8nhAVsiW8XRMAhDGkBNkzktjEIikH
x5p9pjvQtZyX1rcyyk+FHoUFfZYmF3jDZwPS57gOFWPAUmi02TKtwjsV3g3/bZryycipfBRtHAQE
dOQkXRRV3NsSbM5iTvgozZNuK+ARnqqO/dvhLn0OGTH5c+zm+GFdwYlZ/XNzSN2TAefPI6PWeuZo
JtKBZEx/X83XsZIHQGGs92IYCiS4NuPsvUuCFuTmIkidSs1VjX28FBPY59BAFSY0ZNQDBnDqHXqe
3hkiWKi/QzjijSIjA2ssBUw8E6zfzKKS0v0L38Llu2A3s+KAGWjl0+1+Dp6euVMnWLkdGPkj0y7l
MGpJSL0KBfBOUGsve0NWMyom/zgmJ1NsXs2I53CuAhg5mA6eBTEp2Q0inRQKM80jALY331y9Twf6
/0RBVvnLSI1h4kezvPHUosgeuZHFOMxVG4rPV4xNYht4xmhex/3sUkOINO0i+BflXH4/rUxRO3Wu
O/bbb3r36CWzy0SaktwQdGXdh745eNSQY+f7yWC+gh3ievc+CxX6Y+0ehqQ8gtmTxgOPXjQmt47x
BHEoO5L8Kaei4ckFDzErQJ8k8/ZQW6tMFWDm6CW9TCaP/e4w5n9fF6fDHj/nEf1Gl0/A9FredhXk
o9YNbF+vuLQ+FVF0zHU21opvNPX06LpmrtruW8bVxmAJtf25S9fkozbjzLcUJ60/1C0HEm7PGvGo
rTC3oFWJ2q/+P8670DszAchCIjN81n4ulqQM8sokrPMjmqLJdz8SMSTyEO2zUdtJqCeKx5wcjEBm
By+xdmEfR8tbV0p9BZVAZFRy3MJlyOYC396IjYMvFrDBokQBnNYklKltyRwSV4pH0YlKd6vOBUly
mugtl0q/7QZ83UX2s/PaZ+CkFiHC5KPD7Gtc642dg9kiLrcDKY+TGvavOawhFcn8PMbt6Wx2yY1h
8pjZK/lG4tQ5JaSE7McgZSEfJhlRzsqlQpU+mFfoL+plfy8IcbXRNpDI2ybAdA+UIVTF0M9xe2QO
qPD3hPj1/1uUFmLeTn+N0WuNYKNmg4WYlwyzbc8OrLZbKzKU47Y+ysvfVIxya1MxggatCzsUX4Za
rodSYt1bdOVZ7pZW75DXKRwleigmHMCOu2VBsKC8LRfttPKz/KR3/il2yXf5AykEcGKCEwjpRExc
IXW2fEEQ/RmJQeOnGYrrXBIK/H56EMwPg/A4scarSDW4SeqRnpuy0JBOXptqAudfjwnO2KQCKr/g
24PCJFtEhmr4/D+z9qbvdq+Ts9WddcCevGsiFhFvBGhdPFEZ+/JATU7oZrGhT4PmDNK+UQV/oIa/
tRpOYQ+CbZVLKKWHChtV0KJc7QkNbqnl+NEuorlDs7vk6T2qZaOqTNDrxE6DCOk+kNY2BedL+PMo
t9RxM7BUXWRVOVsa80Fp9YT/dK+Amw5aDTBz8WsqBaNT2NkjfT/wmMvF+tZONmFLlVfmcYG2qAe0
eldg9bWckVbWlk6WXCtY5p5TgS9GALvVGKGu7NoL/2wC84P8N4v5RMPjUU09RS0rENFj/rhb8vPd
HF4WGP4sO9c8aAyE7o25u64hfrjretjHUJa5JiVy6/Vm9g8DBmcqpgTJibDj1ks51Rxa6wCh1wIL
Atq18GlRm1UzZ7r4yJJc6Thr87VA1kxvZCqZk+F8c8155O00d9ZvulKVrdoG7h0j3bdGI6O/oGE5
Fy05OA4Wv15LYTDKootszhUUlzMGJAPz6ik1M62rWdiiEnOY7Qo4zn+v+9MS5DMIoVpS2Li1JsHe
dpvll/lrMxAY5FylqSTaCNYUjDcqgeXvM6YKUt4qwdyLIQUm/IEItHB3kkWq7T7GE9UFhtuM3gQ2
KDs3yQWhuZ3wnBhf2KRVdBgUpAVArkuEboDwCd8RozA5zscd9mST+sxDbaYKaI3cHhv6Yng88rMk
/v/xbzcRLZvzYhn4fNuPLoSX3HPc+j4k/AwaRpV1iDXnHUBeoePVEJlcTADxxeKiM3mLBTbYZvJ8
Vh7EPjYucNiDie8BjRHhD6HOoq2jRnwti6IxGmIYxzSCJAh7eFGX/xcghOfaJvmNsZNraveXKJmz
9aK9clYRh8EyGw3imb5h+7xgXdSduGa5oAoHuaxUSTY7eFA8irAWo+KtRGVGlzwBz940vXWm4N8H
I60N92I4CyWwnMqfbI1L7UErBygQBlj3plYhwyfW4PJFUdnQs4NzeMJkRvj7ZCmU/GZJPTrBt2Cw
Ec7icmHRCTcz6Y1KTaacY0iF8xRGzeLgKjRgRnr3uGemCL0+uJLefb1qEeqesIWYsroKpoTL7oDj
lufv/xCK4Wqfy3OpcvBeQM01meGIlgnnZA5HCNfwGqbEhP381dTTG44zNDa8Kv5ezNwCnjlI6RD7
F6rw0ML+PfpxGF8kpBoxEqZWO0nuxO0gHAZTBc+Vp7bb6WOLLzZE6NomkGq7i1uCAqvuLoVrVSq1
uPLvV5GKI5BBObmgyOWPsz2e1S/UHh6anNG5kJ/NuUSxuF4XxPVNroe/7wu/5WuMloqUs5d/VH7L
nOZT5qIjB4SIN1DxCGSfIJm7kSOshMYpZtXXFbEITAqWqFzzJaybKCxLal5R3cIKPo4e4NgFbn5a
y9/b1fo7wYCcZiGLGpz5Qlav0nNbnWUY+kWLTm5QPBr4V74C+CeYQJCGjPBA+n2fXiqznjagZOb3
ZG4J+zgDXMbMjNrbRWnhQCh/9LsjF5Pa6KoIm1tT1H/u/BKveVytbEq4QhU49AlMGU/4i8zlPq7R
ZYp0PzC6wswloenp8V8UBln8IJucflvf2YZGoQHnhMvVvDFe/v2wPzHOxPkCGbZ+UCY3YQQNUG4I
yKbMh0+X3K9YMQlN/u88ziHF+t9YZIDvqR+63zEDpRLyuWikv3mRw7cylA56kuoAXfJ1KN3WXKOt
HMef259CI0fgnQicot7ygYE5uAiJHZlW6mnknQCGNiolnQnyG2BWqb0nqo3Lwx9GI5E829KGpzLt
bHqcykc/5CsdOoocZq+Pol96m00ad4JIq6Xi/yQvB8dFJzu6XvLGsrJgyICSU39eXc08k5jujUMB
LzTjAdx5WBjijNXweCFu9Xj7+RGONCtnsTdlcRzp7u4iT0bHKcuYx359M8lIu+2hOjHHNTltXAQ6
WBpmb1jmc8TZlejZ11UwQ0Sfr/gzry0BOM7ZryBQ3yeWbUJOlmusRIs0fSeHrZL9ELHPZvurI3bt
nNCKa6FEHSwGm2uym5H8K55fTqwjocq08muPQ/RwVIZsp23LFTGSBhb0cwMa1R7s/VCiBd62sXVF
4UPCd90prhk/2/HS4olweDuRE92mJpf3us/mQPYRCc0eZGySRK1RzQprpPehTzr2ByHY1VTXwq4G
ht3IiEI/2iTeHTt0s/Qagnl8kpSMvc5/NW+Yzj0sfyYBvYJ9/fSV0WrZl4mnNZpcXI30RhQ2DBAa
SfGElUf/T6JzrNVllaPLcAyru2S/9jjhArdogTZETTqKGw2Nopkrw3b153mrDEx0TGofEUNVjOIt
5LRTnONPbVCQ8MgXMlYYrj4aqFOFEaBJm4cJFDi+Qdj+ahCibUjNkk9tdCemr+qRG2fyk92PQv9F
zg3rE9HQ7SiTbFuowrhJ/yX3NyZGIutSm3zKYv8YN+qalxa95/GK8OAFhTn1HY75JsbieAfXQd4T
Ne93zHmmW67lQeB2hYjlKKigF0b04AEkVYTOKKr3LI4uT2pKGetOqEsG+fch53HJLePLSZzHwSYW
/3dGFtwdgKCSblllASfR1Y033nu5lUUUMqQ/6cYueRZWxlCqOtkvYUvbM8EKbUsJ6l1xOneFyUjH
xemfcL7+60Nd7gaMWVysD2xUo877ua1N/lZ1jRrXCFbqNop89q1eraNsj8jz1Z9qavqt213CJL0G
9PNGfWjKnDsR1VNkcan+ixMLTSHT5IdF9mjTSWnYDjvCNyGvbny/S/QSRC0Z2U85WvD7XxFIq9y3
Y2ZxAHB6FR5IwhqnKQNyOMXIBhu4ayKnX3cRUO5qum1/DopIKg/hxPHZCXWVlqOkOproev5Dxp4F
swTHPZwS0vpgLerXkNo3/aXfU3yv9YhV3Vv2vhPlNDBSCmiPODZDt5iKJg9gwRAdj73/qkYO1im8
cCUrCpLekdg4IJKdtN0ZY2qtc286PmLYPGlIkXbG0YZGC9I4RbOH/Dg8UjrotrbYr5hn3Z7e7685
zZQzlv8qJ8weEqK8/QvHYl+06DUrmHQnKlIeIDKZ9PgYQaUz0vXA+C4niVE3f3RYXwNzwDKVA8Hc
cLuavkYWfr6yNJldSSxRKf12y62CnT1gMOYuGhysiK8AS6DqUk0sa+bN+1kEpm+dSSdj5p/krPJD
aX+7tO7U1vQP+k7yV46L2hnSiK+AWmF1V3XlSjde6gQkXhCCDy13Q6ukFE8T/92gn7FCV/PAlWcN
XPkaGaN947cuItOdhkE14R6XQy1XPhWnoKoPIemRpbaTAxO0laTnIP49HR1sv2AhFLVTZiiru8zp
LBceBQb6Z0JRe2kk1HvsDL7zBuxdo9xYdo1oQyMGiYL6MoXAuOI6FyMglPqbX+tB9l9entaseWJl
EqdkeEFvNdeb3dmyHQ3lQb4JfcNxOYLKF6cmCji1bhFowhAhx77tYPSL99y/FraPqxwkWaZ4GAew
TeidWvvxm4xO96PMkP0wneizx1dxZxXHFAJqbpYUFR6cE3Ye9Bn/kLNWiEtDTPcVqOwP3Spjg2p6
AqcSdEUlJJcCPCGZvdlu/M7jkxqB3Mke9IrjZyQpq/7BrTqlb2rsdI6F908hlIPeb2CIclNSJUEe
MW86rvR+76BhCFI80Lp5A6MSRRSMsS4RGibo1xZVSCZxhxLb+w6TqPguz0nLyfIJ09NGH35i/LZy
T6jVy4bId+1+1fWzyg1YCYCP22wyobHt67AC9EE2RnZstTRQOWTjWN34Pe3fUXl3lzNEk8yCBaXz
ig/vMJNqoupaApatFZZXlI0pUIdxWq1hvOOgqXn4IbsjawTC+ogPW5rexmsmYWRADpVNlhIP43WQ
9IO/6braeolm6RWQps9jU/5XvlbVKpvou9ar9G9clbCpdNwiqvo1e1vYuwIWib3RdGfLmGdQWiTn
FSmcVCkF2MGAewDG6J9JddoCeOuhQ7PYD1XF0k/X/yrMM/ykwFXcLRLm/3zR7OiiNII+ecI/9Hsi
wgL/fVtVmRkJyiW42NgWrncCM6Es1A9ZGbsmhvLMuuatLCCdsk9Ex4n5kGqmVr1d8m+Ondd4tG7I
cQEUKP9cP6Q2AQOl9s8nMv6DxXRq8iChTLC+fZkf/TDgYeSvTn67SVZKG2iNlGyZJ0f2fqoz4qIK
3lLvxhjG9ffN0PbzYWMxfUQIFu9E2eyFfZgTPAK5CTo0DsxIZvucHgMWsMaE3q5oRyMF/QS/0qna
H9+l+nDDQsuGMyyrxaRItYVINa2KM0ecx20YAKmCagwwTJLvwt0PKWQqIEywIJkpskhAdaHvHkQu
az5ljm6u7muwv2VpjXLc7MJlANhUm4sKKcxMPK45A/9UL4DmRP0qo3npQVNBn1QGjFFDxeoZzcoW
vKJ8nnl+SvBe1xOPjCGivzU6XEpb04JC1NbFE6QLg05SC5MlXAKiAbfWMWD/7I2TF2oNBb9X78zG
mUJ2nQOHPJEzxyAy2gFhbNfPJh/TzpAcnUNSS1lSiaQM48/oKI9shwm7yT+Cg0hYHt2bQNjn6dmc
MHGzaH4+/alwrly+bpKNwzPs1OktgvFX5rHtDYzgFW/d+1B6xuvreoj1a7deQKfXkkwBfDDqKfAW
IMauB4T0yipuzdkbWUF7uKUk6f0FIpuKvzNshW9fLZHT4zoiMr7HA8d1n/yKaR75vL1f5eWS9qch
DK+9mjS1hZj/YyRamDRrVWF4aw/fI/1839ItlExc26CTpJ3VzeaJPdyG4Ge5dWLnaZug3yrba+2p
LodyfvJ2L48EgTtKmjsiOZixYDv2ZWF1kYQRsIDI5EVZKJ2M5aPuOOMfGSmQNaMi80S8XpCf2nET
1Ukczqk1NlO1IQZ2VgTETCicevp6xF6jXrHhpoXRCKg4piB7dm9zNIzYBmjGQ+dEPFal8iFlcl3T
v+jkwQM1tKsDxe061V1Zfqy7ZTMW9wGzBwHx/2aX6ULQX77Mf7ToUD9sej/Hn6TZW2JZaYBlFWzA
T8rpWVCRUjv+V4a2DIH3cqKwbrKjsXw9cVryIO0Cmus2I4Aechhka56qZ5o/z9bz2nz32zu08qDN
femVl3QuGXLVRSLrCoZiw99L9GxYX3p2p/g9SGZFdXWyWYy9pyN0w965wmyn/wcFHa7JzmD+suI0
VKDByzK5LPfvD0CcbDoGXU8ilPjYTJmTjpwMMHanQeF59SP4cBXpqrq3/ihZ9YepXzJymwSgkpDD
dN9rsEFG1UpqicDTxWQvOFcQLDCUzIK7TFbymKgCRKWXXl9uo1S8vCcFV/dWTOMuup95HYMMEkt7
TiIPfOhdaDcxQtT0vKD0EQVw77QHDjW6N+W+nS9GA8t6cHVOFpbueGAwQhXjTD9PoG93mSm1wItI
tg4p04yUBQQIKTBSv06nRf7d93VHB9Z+O+IukaTVSPkteoatAmDqOyE4Nk2IYY1YfKMQlP/6ySTa
OhfZPZGLW5nWQxYeBkjm25Bb17lL3k/UcNLupKYEWW9Y1LL20L/hoVAfJDIucnGabKfNvvs8DEUt
TLBnLpRfHSXnGMd+I1SmOoROpSWVvsEMDvNL/6s2zTz91LeKTKCFm/YHlYLdkraLGYmJ7kV+ujPe
DHeAIquALH3XowkJ3rB3uoyhxa7+YbyWNGbBfRIPZgYDbVqOsvxFAcn766iJddCyrJbazw0cxfvc
uR4bdzNGdwAqMfqaKqU/SjQVEJ6cLJ0RfC84n983ktGQoMrcRsZQDbGiSzBkorVMAkPCN7PbP5yP
mygY1PmDLnyF/SMLxo44HKNW3YHwjYhx/6m3xwz8ZSPY4QiR+5tiCe0n8pWqyslea48wOanTiEO+
44zmt2vWYI6VDHLgbAdAPtwt3YoQA9Qic0cj1YSkcBrqOCl6+L7i3MKHvmhOvdyWVjHN/T1uajp+
a0/nvV2iNJXItlyJurrvPXgldQryfUNFIcJUwU+FG5eKhpZVemLYIMRuAf0SL518yFuawfjbuI3M
zcGtzmdPNZjP0sgiWj8ewB1mNR8DzifTOlbkq7HSKdNVB/bKX1DEFSferuwO2ei/zZ+TkbGUcyEF
qUTACpghrYKl4AB//tKTeOyfeYkjuJpAhYAQCmTC9s36nr7yvNVNqVeo4vDtjQlv2IXE9TK0bDk2
d+WhSPqni8GAERY2DrUNxjLJb+g4/lKWWw/hEFqCCHALEc4rVgbdQ7y/H3u/fZUk7EhCVr0Ly7EJ
dUHFaISTuiFo28qPwoJlXlObLs9kSYLaE0wsUHkWi0NtglU1WO9vWU7tQKk8AP+r2DNuT+qXGgUy
yInHeEgbwzRGg1XjLHxvAWcTV22pR6XXknIgaLNGZg+o34m/tEqPvZ9DCwSgGu7y+A2GNA8U9Rga
DHK4wucbTDVxreTszj2hU8q/RhNkrJXOWVRNobX0yhANpfGYQSihu5Q8tZo1RkOkOlCSEjcwkw1r
z79UGRKU7LWP9vjxttVTtOogKI7gwdbZ6/jabf5tuhVxE5QAM4tlpXA2mr/FnxagfEbjxdqcEJHo
wT/2LUbTnrZ9l01PckF2BDycFHQl2+273er1WzFhFV3VYMF/wzzXMgQetfdHBoK+SaM9dIsvnLWP
zWU9Q3zvY43CxzsZsCp0h/HOe58epzInckt9N1kyKnibGm7fYCENhy4MN+5tM41ZWontZppBZ9tX
Cm8Z63UmHiepWnxdILZ42sXCwtqq+5MiX09dWzCtdi+u5KkIR4dhL8vDdO1TyCXPwRkAyVIG/se3
+QGIb2vOqeI/rycLnIvidab9EnguAupwAKSx1fguRjgQFI976ZkUiswkDYZ0jReswW51ucxXQ3hE
u+sYfkA+047k62Cf/B3C6Qks9k33t+uMqJ056pEyNxgHZe+W/JLzDvlrov2XYcs8k6ESQHXO3iou
z/DpNMhgBikLE3I4GJku8ogjl9R2ICLvXeZ4X5VmjeaNo1RQjNP75XMp8ntvNRQ3ZWQGCnKS+LaC
cvfRqlFIfIwwHmTLsDjhdzX3kC+uhxbIFJ5RS2Es4tNKZYB+k+k/LWLeRjLSo+Nu2vJPneckIXVO
6h7Nyz6Rlx0oEj7yyrdUBWC6LdyyuLLgQQSSrizXKj0k+p4qZgobhFetvRFkmveklJASCVXaH6Rv
SRGEirST2qKazNXJbegCAJUatfbn0H9b+bCn5oIQO+Py6rN/1vOcdYuHLsjW2k0XMvEDX2efrzBw
wCYfraTTjUuF5/K2UxM9dPmnhKK4q9RuT2ZXYw9SUYjHslsim32pnT/0tdTUaC73dTJlwG8EE7gs
QHS1xL+TS5UcZbQr3vbGXBmQMNC2Uyu6loOK3onXWXz+jgyXbJ6vBfWUtBeLYLzN5uEK/9iYh3kf
5trvm79SkbWDD8g/eWjPCexaSBvivTjGv+uycLAt9enqabVQHXjmekXyxXOlVVKG1YwKNY1xdWIf
QPDqIqsXUfwWuUZ8AcA3Iy4bfY4Kwo4Gr5mHdYQ4KIZgBRbzWwUCrkkO+X6WfJaHUafz2f+t8969
bxe8ql4bNwQIWOa9ixtezV8lUgUGrRQ0xzVoBndw+Y/1jCz/T5cUxVTdy5abcS9eQtZxPQJvPmG+
hdhMgbkblYdlc08hKdglycLWtJaFsiIGxP38N+sAJS0PIYG1FEzGo33IMmboLw6Ufu9B4HFbu+eE
CFbIIT4L0XuhAOMMT+EFJQDZoN4oHSR+No7Opl1zxExHp4REcYmBFMNKWn56Dp+8tWYF9HQ+ItyC
yCBFi5KKioOfTi4Ls8U/Blrm80eNGixKFJaFB02RuwTDjI0EJ3N7m5gNnf3/mInSmiUE0qBU6drS
CEEjjWwwDPEKF4twtfaS5o7tfrzFrnRfBXHXQPG+/JJK5gpL33VSTXg/D7XhqP840px8XsFdx1yt
I+4OcDu/Houz1Gu4X1UiADurfwdrdxpOtrN7FfdO5qGXpyjfHjqxb2ROV+qb6Y5CrrZQlFBPwtiT
dW286Wnr/DTDdEuB/h1LSbxfvEacjUf2ARGjRA2juaFKj6L1f8YNxAeO9xTyC/bnkTy5t8mK0VJp
yULT4jM0MW1dykukHZf5L8akbSdhDiQbCDCJQQ1JXBLPaqZZ/zpVPFXYUmwQ/NaK1pDZyNnkQDMt
y5O75QOf3TdlQmGxDM0OVn7I5IhYDVKTpRZFFXRuFnrfrtDJnUoUcyFUwp+kKH+cfEKrrK1KJxXm
mYyF4si/I6QxdjGnW8+eCf3SS+SD7MNrrHXvFr07xMSHzaauQakByUhcoJO4NDAoML5Nk0Weqt8M
SpZNZEief5a3hlrKHw4naBlzEZfU8JetDoVPAJib3RTbD9KnNyW4Fz1FO8mGMQQbcnxRU7P1t/FN
lYH2A4QcpBVaIulVKwlqzNdVeNz14HRONxYRhzO7oFjcdEx1Xf7e/uj+EtuGsnW/UmkE61HXmcG4
N76U1uV/HCOcMHJt/kvUhXjzBcjNaZSn0p0cHaMwuJoYKmKBs30iJs/gqmMcH4xVg01ZopAhPj4Y
chXk0th7h0QIL5y5Q4NnkVQRmpc2eiknf080eKZIYg+qQhtjONn0SIrqAYdDToolngqKO1GL038S
Vpr3BHQOOJrY5Rcpl2nLmqhnq2Dl+oMU/tKq3kaTKf22W+ZKP68/2CyidxdNNfP5VkYCBIqzOyrx
eYH1CYHmMD5MfPrB6/DEUPK2ZsgJwUMjgpGjkybB7UPXgIbyqV2jus1neBPsIFURIxpT7t+NBRlr
mYtQadnYUDOPgdMK7676R9h4UoW6RlvOoE3j9GnIShRpNwghll7cjqRnCrS0VFtCee1tRdgIvYOp
0UjHjVxRmjlyfWxpuZCk/j4AOyvM29lbr7zUm+ip5mOf8caWkYgpq/QEUf1CpHUqrcKec8e3uszX
iKxqOvqtPeHzAtt8BkcgyTsYkO8IUcioXurusyRuit6DzTl92zycwxC8kAJb/S/VePeep8ZTc553
ol4zV372XSx8Lm/2mdrBj/94WAAxjrjjFXWGvG4Lbx3V6w8qUWJ4TP9AbYKAop3CHqExSSvAGpda
1caSfMOUqyunaGu6Ru0FJMk3c27xuSsHH/jJ2jRIISQHqF6cwX6PDVHKmvy8gmHmqmzpUPEQPLmZ
Z4cwEDjIlj0QvU3ECGOBmUo1csF0mBTPVBBf8PkICSP9xqd8+SEbZr5uz6QFeVcUpScGwZowJQig
IBSIYxduFJeSIeLrrn5IzRXq83VBdOlxVQpEsEYAqwr5B2EzTi7UPqRHoTCxEjaZSaez/ePyfZRr
Kbl8LpocMw+XBgl3vYwraalliTTXRf3K9hX03A/nwp+SO31xm16ip7ucR0g1zOMBZgdnHjAImnOX
/pslnUCeiMLM8Qy5eWdqQng38NSUrgPPYchDQE8uajlfplsX7Xmj81eXSM1oWCrFC0DiGERBqve2
/WthZORNA5KMjXJZXSI9cKov7kqBi10T2RcRphTrIXli4nkGGhWyXuTwD9U6mRbQHzhxM+ymFnS8
SVlF5aLKtVG+e4qzwCrtdw463UjnJB8Dr+x8m1oiG00xLmy7bzd+cQ8KlUVCRDxd5IrVskGDYf5k
8AeuZ73cuxDltDYmmmCRbXIHxpKcVx0P1RswvvVRNTQ3Wz4UG9+PQbycCMWCN57xgoGVI1HFutVM
mAbjrJDcUcV1T7qfDWLGf4xhNCdzqnMFSRGFENT9AL5MFKdj98ZWIUNzGkdYyKBaGg9kRY+9rtpc
UmmohfFswlYS3LxnLQ60mOQyKB0j62srXMu9aMqtquiMIrsXknsh1EvzrkBDxBsJKEg69WqNKg3d
Vr0HznsG4Kf8LVr/zsLi84gGraLPt31xsfFmyg5YuVKa0YxduS+tCJxNmAv0YLpgBpYwoanhSp+y
s+nr0h9DK1vVjC1t7+bsycjgKt9uVCvAprWjD6Ga0p8cAUpahejn0HIuT1NtdCpUZox3bKJYpDOl
UjlxAqOMucarGRw+D/dZerM2AjCPy3XCcitiqyt4C9yMp3IwyqY2gvRv6i6qFfvwuUOwTf7kvjoV
MwWlsmJymUN6N4T3YaAMtg5I2wk4fSo9uzBk0Gr57FrjSD5CZXOjYrrXXPDKCv+VVT97d8pND5j+
yE7OZQaXSjBUn8/s0EgZ4uNjYIFCB7w8P3u+0leR8mP0NRvN75zaW4F60YQXpMMYkAi1f8+m2Any
+SwFutLnoVvXvockleaFl5ck4qrDvbhMZYrjrdRoBQ3Ym9GoDpYK71+vGHlBaC+skUoX7A3Ky817
7sAXiDtLyrUDQv1n1WDhcyerkNZxASj3VKPYxHoUGa3MUeBDMCAjG4AWmg63CsS/TKXTq/VFicpz
a4kvkz1zQYACljonlz1AeuRJUdM8adb4NpMODjbFuIHbj7/eLkg0TlFAp4Q8l9B0MDGh3FElKQQH
IrPhx8BkrtbEulqJF9FMHYsd1KcnZnucUHfg//sMKiq3d/+pfnA4wRcRwtGTUwQhJL+1YSYH2BKr
9hxfZSeVM7Y6KxNe6ssUHDAopTlBq74ORoTSCB2aA4UznVvITtJM4eQlP/bHEyqDJH+hR3QYMPL/
Lf0wOBKaZC9UldnCXP29ZrvjYj63382R9bTQC3JH5M0RlDsWEKW3+AC5LRLZmyRG5mP2S3uHUaeJ
Z57AN6Xk91X1iVFaZiltliYocYpvhmLZNgee2+7S7AHJdPWYnM77nmKN5gTT/qsL8Ijp/VzqmUgH
9HvT9ZRGabb83AoG9QW0Sx78TgcPWzkFToM2PvuE4OvuPnmRM5FAUH7OdNk6NRRTXsbmkOyAfMgZ
8MSanYl0V5JKGbb/RKCK8Bt2j+McIcROippE7b/YXzW2Q3wzBF8SkHe4XpTI12dbxBSyF7il3wox
zk9Mw5KAmaZezJLB5GSWzI469yBM+SP/oliKKf49nW4scyy77r8dvBjRsmdmpzRvyFINfmyvmBnm
CxJquLj/ElrTZ7cLwHuFkBXCaP9EV0tTWwxbMKSrB9/QE9yBpcyKQTAiLlvEUqO6sE2oMUflsYQs
OSoGyOVs8HSnejS6cj4NnQyQzeVsR4tid1xNRItWS1VpJyuRUjgcHoZd9Eb07Ojwrp02Mr2Cvyn9
qDEGgwsqjj0EdAymTKwYxlZMwZtjbmu9hmdMcr8YK52R4v1xTyhrydyjIuKU5Q2liMTBy+UCtWA4
h555bdgxQ69W8z8B2apbw6+awRyoEKVHHWp0v2w5hQiQaJy4rbm1y3uiRwY/xmNwL11C0r00WNgU
6YJB+GnUIAXiP9gL/633Q/KXlbKpHoO+e/9IHdrd26BX/JQdc8zuwJlh4+X0M9cmp08KzghsBVA9
/67fYzxR3Sxk4RkafsG8vMQv2Vi7frGIfprxAGynLZqi32k4C6eBS9DVBlVFAQrNnRwXd7GORcJ1
EkhSYqvSCwaPsllf3SxMcTnf59zFBr8sCgVz5OzLX1YdWUg4WsTcNvaFM+UcptrjTgSnUez7hPwc
ZHjTp7WK9bGucpI5tCSK0Cy/b8lyRaEh+nFyBkGF0QED56mLyWAbkXfLUcqpH9/d/LYKMJ2WOGEQ
It4rzd77AdoKPz1p3Yl7mj5388f/5TEyqK78FHeEy67pAvOLH5pJ9qACxgjBQuRuczRT3lRu1awt
TMcZeiWZL1/B6rkOZ7xfYwJbXlK52Z0HcP8FNgy7uNTp0TNdB1P9FA2HCXiuNOYpPXHaiYFACa0T
G7MgKu3V0RfNa7QOGzOEZleIyCbMSEA5SOmSRdHA/7UQNGIjdDLUkFUHIK1u2UdmBTlD/OktPGik
izj9ftbIK5QLDikYl94/WmX9mbH1h4XDsMsk7jRhWteCCqadR7K5cSZjomS5a/zxo1eRWkh6A/S0
2mET+UZpYCDOcj3m7pe5FHB9c/YgE6B3T8ebJOnjfPwKpOx1hun2LFYdGNMUb+XO+QDefJTQh1Z8
NcnqLKsnVZZ9JQ+L3ls2xsRfZLfcfN/zkemo34SyP7Lnjj1WYT4d1n+lkB8Ra7Mk41h8haKhezhl
Tx63FVhNyLp/gF0ZbQpJsUh1ceiOs0F3BKuLIbGzKMmmxKKd9ntjzgpNrNubLZuYg/6lfDHDNy4+
LoUEp0CG944UaPEpEozgUurVUO9MrHSPrUi/ToGI7FAiQ1C+gFKTOgWyE0D6ybkyR12JyO2hzz+u
yf84Zlwi7BbahlRTTl6BjC6bW3mNjOWC4eWBFmgKdOvgI2RC2FxkmruOqvfOp/w65QO0sc3fJbFO
djrIoyL57xlyE6zmPKv9YveCw/WZIoUFCtCu8i8yLAtApAtzoDpw2bgLlH9egUkODhIqVqmxd5uR
VHhejIIoL34ajmpdYAStGupL+8KwdIZepocxk8yD7NnJnLr8gZp9WB/Xip9GfQnenw9YljqHIMiy
a57UtEYT0cAkpPwcOFKD2spkVnfGGIhXQXTsiJg97dbE1okggQIWutgPXQM6cu5R1T5rhaeE8A2l
dUq+mWePede7kkxnbbQKl7+mOhbU0Ttxu5VIVB7EH9TTPVMp8EYazA7s964bYZYgtdfTDmaCJ11Q
NTs8Wyh6pJZp96JswXQkuf2n+0F8+tFGc2sBwL61JiuX8gTC2BOrnBkKFHDQ680q0OAtuIR9DMQM
42+MbkHKGSTlFUptN1Mxr/cwY/1P/Odbdy07Ft+GyKr2i9/RzbyhYB4Ghch3n30wW7Df0wiSDcHr
ZweCie4ofFWACjWBdRdghQcFFbQYZE5QKnPSmSbg/9lj23bsv9CrdRsu5l3U74iIfM+tnGWEFX02
ktHvItimjC+1FUupu+UXewP77N92BlGqukb1B3sMPtTaU+GzJfUOmxwfTVL1dTwrl3F5Y4GMLDbM
bvlKVC5nGvRb+hUxvbxJUKwPZabAoXE/VMnhc4Qolmw/fL+u75H6bhPbLDX0nGtpIjXqjFijpc9D
i9Tts73mA5MLH2DL2MQLDaw/3ztXFkRfAX0cYWMUkWhHJIKsH0o5sL7+g94BO6L5LgfkS20+sCRf
Xe+v8L25+ZkJjFEJ39fYlSjpq7+miRve9M209NwmR1c81NF/GRKgud1iH5U7axVf9vFYeCFN0xAg
vAnzBi3sz3AYnEdzJYCfCjzjNio88L8meFx20FSSWD0AOA3NJ2AKXvFW10GD7yT+bEhfPD3yGpFh
g+boSZVh+MnN0biOaLwgOCDA8s5FhQBcHnkg/+NAlBYpfYskjIuYZxSkWKU2f7BjIGNcZ+dLyTgz
+xvD1RYjjjJJwJ3t6DCrjL4FeFISX82Q3s2ng79WQOT5uvsUAOfo5S3lNXkYiecKyOn2rgGEFLjj
1uUZAirxS5vTSPpedA6Kom1cutRQ6zc/WhpFgKTo2an2KOvCBRs++dsxGGsEk5flkIOJ5wr1+IAZ
pd/cf+2HfxqeFEP1VuYfvQJZGz9kMp4XmpBLLVFGIum599O7MR6ai8yk8s2Hx59doIbhq/LK3UNb
ceruqMBIplJh8dDY5dKbgU8FTk8i8fvuQDu1MUcUauP7BcFi9fLfpmINp9lWJs9Ss9M+OWU/Z9lg
WT8H+DE0Pk5A/JCWYQQ6OE0wC4WvYYBdnXQ82ZWjr/4YjVlcDoatrsQGqw/ILlZhpX0T7fNELi12
hYn26YSTjYK5/gJkImXwkPllpuf8YrdgnWmXU06gbHpaK6Ysm074PKvA5Zb9vNwjLUmczFiV2p0O
hLUDlvJHnM2S6VAU9N3VNW4+qKER0XyJQAvxx3Bdb3f1y16Nir97bcbMc3Qu35GJboFUF6QaeaF3
Ws0pJLeLLc3M9lxIpX/uixn0/mWBxdRxVAZ1WDkXbYEgkWDUuclNFrM2vBfUlQnYjuEsgnF6pkgi
n8tOna5fSJuhYhDb2wQYdmAJlDisNCo3mlMApmYUYK72xx7f7SvZvrgpTxj8jtwfRFAUPM6I8I10
oXMTixM3zpLA2EVICGrgiZXi9daB7H8MzyNm47pxpPmb/pL31GeOn7fAru1lTcM8xgQ1rRvmSq3d
Y9sBcmP1WyLGFAP5NG3NkqGSz5WaD08Utsy/JwKXirO/Uw8jDNYiPt7N8OpYKNpN/x2Alxkj6vQ+
DOgwV7fWym8lzQKrb+mfxzNb2uZLAB+8f3S9+HWVyGT8zk5jk6eJ/o6UOqU5aemTA7TRpG/zL/DM
R35wUHHl3I3t0Zwxy5zd/Xb3pOxgAc+24WgNh196WJN0SVvD2GbhIMOXyj/byHKCcukhh3WW2WrS
+c26SuXpC/i7nZZo+IhujrRAGeQ+rHPQakOk1+ZG2gskQu1ccIX1AidrxTe6uAagvmOZT6D08Usr
dpK+cyzeysCwu0GkUj5WqAclXPv9r+aXJLWfmpRzHnGZopAPGzdfne4sfLOLad4DPuRwv1YGijnQ
wsaxoKh0HYXMrid59L7kCr8ddB0qEb0mWZ1paYTldOGnzEwkz0EGVznGEAq6TBuCZIhECWgOvm1m
SAxXfYJY4B4JdYes4LhI8el+y0x1e3RACTea1GTPYcynX34C7sm7BFk3CsjXqrGtv5jWfYqRMCEG
HFJ5UrZlHoM07JlEZrDYYBSDELr/QhTkXM05IlPLOIthE+zK/+NxIcmOpd0JIDHIGCT8zi1isMA3
E3iSzjYgfDAu8VMMBBx3rqxYuTLBuI25GvV95cHCmwUhxaowbAVRQyRwtv3nKZV+vBIqOsbnF3/f
/XMq5L6jzXC1kP6yNJjAlTggRzrSpe8KPM9AL+QjfQ6td3BV5R7aT7EzHMTY2xwydPvnQYV70HCn
wINkW2mIlsiZSlRwyC1ESBKNTZuFbEQSSI8DbhLaxPyd99xssi1TXWfjVNFbiWK0BJ3pTLE7l4G3
ja4QwfnuEBOMp0C8v/rHAMKA7r5GYdZN6Ft81o6uXJLtN7XoBh5e0KcJMz2QGIrGp/wl+QLTh8Z1
D7kzvgGIiAUxoHvzi7jtfnMomeZ6NZlpOAvIQiIFRcMnd/FdskxBALeVxofRiPht3txG7zWXnTA8
e7foW+KreLFFG3z421kE4w4jtSnlu2HgN/sGrE559BZk+xQG96Js01Bo/JYAfMh1BfsBzDeuLdGD
QTKhEuzRWX7cIFHamY9pUqbb45rh5AUZanw77qLNTUEL/0xOrcD9Nb8a9BcnTlFOLwa3wILh/ATO
sorwTOnvKJpFfjH/7b++sWO6m7NLv1kH7X1brCcX6wLiOYSPd/T9cL3f1DNUlpWxkZQAJCkXUlCp
tDz4nK6vM0DpJ9q5znSl5MxHvLD7LVdDpLMkgtgWyxCORrq86NRuJdY7JkTAU5igJWO8XTuYryJ2
e67WCXC39IUaopD73wXkhiRNIJjc6nqsy4cf1DgtaXUGPwEdrtG271HuqnJzPP/a9N2ySaf5NNyu
l0mNJ0tKJTnFXSgNkvB1cpAfbVXxmf2dmPPbkJc9yAu5NVVNBPodGKv0KVuvg1ehO5Skk4HIucdr
9K8wMT1H0VRYDqy8vcn+vghFb8e+GMXo1mNouHQxtHhXvT+qcgVDM9pQh4IsevrhWwtc89D3GKLk
0C542RHRkeYl9hV8ebYzVgmcLAYXiIxciQbuQmYKXieIqapKfpb9HfbeuXUY2krNZoerzsZgMcSd
03g/PV1UAtDEJdEs+YFEqRXaib0A+4wi+eycPI9YGwvGZGrx4i4Me5yUVIi8pcjQq+g5bJgT5A9r
djQL0ckrp3BZ48WzDFz6ZGCOK1xsql77nFDCJPKzM9AuzFYTNcynntkpIEpT+z++q7etTEOXgNW4
JjJAK0QLmShffp9vckg2ngFZxC5YDdRLc9OWProQKTuVCIsoWJ7FR0gpu7zAfW0/27a4hoCKhmQS
Us/E2uWJbcCgQ3T/8AQgFfsbn1kL6VxAxbYHkRWBlkJ7VP41Uaefkouj/3tZ0tCYjq2uGNO+SISp
1XF5fK9nNyFZl1AjwdINt0/V1ILuhC8vcjrbZG5khUHaLecwv9UsIrG/ASg9/nIPgkj80BlQCbx0
djle3bnLSnNS1O8lsOpaxRuSVKc4Ok7khkzdBTa41ygtxYpfYq4xhN8pjWDfW8W2ZqN+Z0z/Mbsy
nMCkr4V28bYqGMQRmxjunHnHQ3LX8vvOdY206Gu6DaGrIdExmWzvUxEaJNCHwQ7/V87EjlpfkLW2
hFk/hwiuXwZxBVtvU/o+FTV9O1GLI6ZNCf9kHscx2eVXOkZRasevLlkE+EC0gsjDdV47RZw3fU9e
qS/Kg4R3xUZ1J7wiap5zFDQWyYraRf+K7b15aSaPYFqQ5SxiKY0KdfcljVk4TbVvcN4rPSt3KYeT
1U7bq8BLw1lRL92r7d/KGxnzx3JchW8ZmcA6N0hI+pQQ8onVjHwqwriMiYa/tg8OO3eoo1mFcwsg
hF8mLDALiRBaROv3nQKl6ndDVGt5JsUN5lIulvCOJKK9pDUc2LeyRF896+Ibge1Cd0p3vkmCnj5r
JdVIlHTuCAX+s9IXbvWijN3gbGlhYL80eqvkC8BJWQ8IEI92/uQMsm56tObOiXeY5PgmsPimUojG
kXqp1Reeq2v28Qcv2oMS3+/LpfD00OEr2+5LlGxqNvOec2ieWWaK1RwKXz8Xxv7JoIzm/uCeIt8c
3PRLMiXw6zolArnTjLT0gwypUelDT2a39byTvdbRzgaEnY3p/3HpVq9C0d+UhiYuuniHe+JPuupd
qRgNy7eEntfHwros/OkS5knytjeuNleEFZw3R7dTaU6Wpug5lMvSEJmmeUXYjqcrd6H9A4im6lcs
SQHwEUANy90np+aumogLt+W2Tjy9l4nIsfjkr50Pj4SeWtXkj6ykvStta7Oa1Ws3bj2KKBlbeBJu
VewZ9XRW/IYxL86kfP5MF7toSqZhghGKSdPmWRqYhNHjDdjvsAzaOIznXaObCK45Sj+AN9VohTlO
PmPugVFbMAKA2RT5tbpz1rBkioXsDWYp70rLyA89nd5aYV0Tn7LNZoSiDzSUO5Jf7V9oaAL0ZoTU
uohF0My9rqj6rG3pU01cn1/FvdM1QDkX3ocyBacvWAp6FDFlnGcGwNRjcov15k39dnCdPRFEFyID
YtIq1HltK3wt2hV1VMCOVCifHSOUdL218zYMz0GZw2JaMTnM+Induoeo2Ib4LEwrmfB/EWXGANO4
yQdLi4XNND3HLuHRgYhuqszwWEqq52o0qVEEklhbQ1ySekzmd1yuczqkxPbNGJPuNsXXcQtM0Q3Z
EyDAQBE7di+AzVIeQ+gGxYE4F+ECs3e3lWne9ekcRt2DuqA+BJjmbVtZyDfqD/bFGJ7dKjB3hHDd
9BxGebFChY0MPaBekgyE/diidn8GAE8aOfApio/sGsvEf/TxCHSoAN10rEKr+zuwrjFNcmJh0TN1
XI552rAC+kHzNgKzgvj8iaQBOFV3530CaplAYd46OoRIXJ5yoL5nexl5sD5Ri3pWkJ/O2nQ6PEBQ
vieFTJJiKoC3FdEDMiLyzlA378qaO77jglxXtsQ+KEhSCuSGD0tJiTO4Q75eVtHgpaGUDWlJ0xxh
bJIiudZDeDjMGgrmwPZP0bUUpgE8d3bkcYH5oYmOqDSyugcLc9VlPzoQlcrWd6kmHIHk916Ng9NQ
i/xSojqaWW5LshlunWTlwhNEpcdXlwfx3BrIjDEymrDDX/AtathVUw59j2C+JZ4T4ddSPv0y5qdE
6tUAh/A3HUeQxnCf9miIySoBeIXMBvubFgAnY7WOwL0waKF3yNFyfEDrszZOAi3/nZbusf0KEYcF
Fws62pGhPqcEPCgyWVcoBWDGaSwF7tvx6ZlN05I5wAPhiDWAJm4cEE27NiUJtmd2Hn9GBIWpZ0jY
+G6Woy44Q+fwPjroGuMOrIf5O0Vxf2QONeMmhpMfRIJkiZFQilM48CztAss4Id+MKJD0ZDsFl3H1
3lneoVgRqwqV9Gc3Y1yKXzed7oClfd+lkI+lTbflbyivJ7iuTF8AcfFK3QQ4ka0KdaY2aH9IDGug
QeYeuE8jQyLp05/75cs2Yvu1mXzLJjDeBIpwe4XBzbRM0oSN/KmVYgxaGKPFU/i5byfnVeZpcK59
nL+yYn2sJswjYTwjEN8rnrCETvsF3SBpk5CwltWKi+yRHCOmC5xusCYVfj3Bmn/Z02PSN7ZmckRs
noRwIuTi5j7D95QpziBqFSl+GE0whQSYqY6y3b03BqHBkjtvmhxqcUE65dxXA1T//uGk+MKpB5pH
R9eGqmd8jwrPAVXLr+xwQ+i43lOFP6WjCeNqWKian/kF9CEb3dwJeHIPOv0RVp9pbVwK1rZi76TV
eSQgrrs63O58Rn0IREoXEG+binPZmoHKysjHt7zvlyKCgHna7B4mgmTBhpMK98J8bWP3nho3gxWX
zbE70yJMrmdDSVDzece1x3qYaBbw2T/T3Q2hsjuveIpX+t1ptZkpo3BnoQThUKpsWXU04rW1x54v
Oo7tpUkiKXf4LyC7Wm7NoqhKWkwaAC/B4Qs0waRRIoI48+z3tcD8R6atecprgvBdYj1V7UltJ8Gi
aBDCfmal80/VEc14zoeKPS+kcuDic0UHGQZFyRKQbY+R94XQ164BRlW2uAGsF1LYhJPcQ1qodYjR
UslWs+0z6sOi2PBRoO9d+IFh0ra4dZbp8b8eAQpbofhGz/yk3hV/WVs7nzits2NC4mPAFqzmPQZf
OFrY25vDr/VdMIx59Wz0LlWlQ1q/Vtf7fnTMdQJJt0k5U1xaqHA1M0sJUf6zW3nyXpTP3qDrWdQv
L3gZdfjSP8LbiFEATdA0SQPvqOMLGZXl3MJAuWhmlq3MGAd7Bnz7nOm5MgxPC4weCrFAhtMKcRfk
1v4TjIj2WLLphWVfJxv0XCJ+LSdhqzZR3HlW4sHAkxwNPViLEdddPHjP+Y3vISkwONpLVeDYEtdP
1faolzhH738j1B5UDUQIl3LbJ1vozlSpJ4+2hMPKVIBZuovIY0BH6SHMIg0quLz2do+64/ThQAGw
5LtnAE2Ht6RXOYE8zjkr/M8vEk5GOuIUvn6GCNcA8pbSvzS629Wf/oVKnwld1A/JzHFEI2dyTHDH
YZmWWypZzqCRBH/QA9qvfRcMPiRSUng3fdWbuBnAk2Gaxrae4SmWvbAahktbCXTwcYgg8+CxPHgC
EFSdn/5LfgiYR5cVNSgCJ/Y44z6TA1YTHO9paAbi/TadH4jxoMchFru3HWTq7WtAcMv1D/Pk+AEI
KtMOLXhIJ3S6FgAXDCk78iwR8MborrPMIM5WcYtzfigwGph2QWiQzILFai1jYCAcGFsRTRhxy6Io
yiv1cRzv+AN8N9EFM74i+oMm/lYR8ez3ZFgvKGANZ/q51w4EPcbT61ic7G1j4GxSDA5d832Cyids
Q3Gfe0f6xEN3wi/Zm4gIfzIQBZ5vLtnukiATihB059o4t4Tq2dSlH08H2YwSva7+p1aJ3Lu7Oqvs
WetwxHwP/FrpGtZh1/CV7zsgo5Gj5plrs4rLvNOCWbXxetw1oC2cvwBdJvgoQBK3fmqD45/h2VwO
RC8yCeIZUqqY2vFwMjNYWaI4UlG4Xs8A+Qfh1Zo5Mt0dp+vI4nA2xlI5gbLVZBhqy52LfusF6/5U
+fpJXKgbyZaLkRNornclCiVroflT+ziV7c3BURW+M/5qg7HNfRXxF1KgEnx7yBpIWr+6r0B5JwfG
5bTTmIJWw0eMP1OnkUMlb3WN5lbQOAYFr8MsBaNCd8KG+EDYgCtAAIYpEuo8RM65Cmxcy6IvwTWG
uclIF2VmNvUVqCCOIl4fKmtG8zWK2kqdTLxaHI/ypLL5xf8jiEBGkn/0d6n2jDMav9cNfcss38SN
603RQP9YdQ8NuOQGO3qt20bgApEF9pALDOHaujp+RKOh4dy8Z+QJ3w0HAGVKr95S6OfjRbVGD8/s
YwqJScOdTWmfWjELjEKtEV+HargjGVkGblmk+IZyG/XZtSrJxVZE6KaaQDUPwDKkPCGFmyuT7jZy
l2f4YxHjAUbJePibVC4k9SXa/t4httCRx56rwmmW4N2Cnzl4EXU11Q/3W+5FsWW6f+DxKRwWjMNR
+zL5NMci20ByKlRQUM9W0Oc9TfA23IQXBYlv6WfJaQdGSeXC6EHW9Gswf3xq8VuBhdxIph64AdHw
l2VVh1LYkeiYtk6ScodfYsUHVnoprURkvpcGGuUVU+Xfh0p7PEN1rGdB5yU7FTdoD69Mv57hJxKL
OZMQclllElNiGC221h8Wp/LkyU/5Qp9KjqQlar1JWB0aZ45M3l4pN5MHCxOmqRvD6WatwNPjuvDA
+ATTDZIBbJUk/j3brc89aCf77s1zd3rZxKvRtt/VXkzUzzPrZ1l9rMUe8lTmd3vpUOQajT7qqsVj
G8QUvUz6AEVy+yUr0/l2/R0xZeCWhYqO/WSitkWt/p26onC5X/MmdUZRSos0158eH2Ci1BryNSyB
yvQagGfOgUrJODaCflzmBJk9IfkI3eDN887mlXCwfNOQqpKsOXXowCSnz0GEY0IfJV1Bjl4lrdoJ
0vxTe66VVVXmv3JKjWXrltsFE3vgqJ8bakjDq+esvVH2CZDh9eUD4gLSpR+fTA0Udm/bxcTI48w/
PN1XmgmBkhsd6OmP5GvHgpMne1F21pKSlkGh3kt3G8n7ak9Mh5afZrkAySATA01NsbQrFOYcskZV
rLwBDdQ4tBz0ZRc9KBct210DioLq0qkF0LsGGjHE+DeKXU00s2P0rIumcVhMi7ZrbGgVc0HTv4HY
rkJi222RqQCMYkd5KSjNnhMCL9hl5APJwWPeffT8sFwuKwWiKcaBLzmVUlPg5KQSKTl29MksnAYU
ge1PBeaij7Y11U3hIgsJbFFzn2NGRwvciEFUuwXbtZzhJfBl85TWJZJFK0GaoG/3f94YhBToAktj
k3Q0qqTIos9wmYOp/PgtV9FfljOCrb3+VgsNYdDc0XKNkVWPnzdinrtbKkzZzehXKFn/bOr59Qcz
eGR9AZEFfusld/3u1l0fFOj/os9ysKsBububAGda2+cTv+OL+68yDQFctj2HtijgaOUnR8RID3YI
ohg9Qh88tge/2b4sn4YSRV1/6iG2MyFF9YSzuVE0KpaIQl20vlNBi2H1CP3NiXINkZQtxMG239WI
edgT8Bx/CmSp1HeOPYfy47kkePr8PF/xTadGGlIt0ODVUl9kv8r6VaLmi03iExU4w7K4metviqX2
skUvJQ/SxddlpkJpiOn2Z0WhRgRB69VGBqSQs4JNo9XtH0NHmhMfSpyCkBQFBz3nTfiNwLxuF4XJ
cU1K0AM/dI6VjuFZLrDTG+easw4IREVcZ+3ggeRuRnjDQu/UGO9NSZtu/ejJrq5gB1rUOYyIsKol
u6ZSTvHTkd7BE1T8s6NWPSL/g+CDDgASQPOxQ1tYJqVJaSy+u8gUXk1nV0HNbOWJRZDWgNwgvb3G
r3iZXf6Wzlea86EuQJ+qrg271Di01C0p1M3YWxsHQHW3dJjMWZ1uOBcgNaMa4I/uqAa4jPS1y0RU
Rqx9u5TpoOfoWZY5k3X//NBUebZC0LQ20mVIA6CcwRuYFG3PbYX9sPAhRs0DjZbqy0uR3w0hEDHn
k6Kh1jNm38/INbF0IEl6jgy28yzH5MA4nqs5maSCBXrLzZ2+tVLKCnqeZX9LVWoxw6kkSwdowP4r
XeioGLw4pULAigc0XIDU/clRGDh2xV3HOFoj+IAyCy2m/O95uab0Nh4eV5KIUMrIIcowtj1LawH2
y8XJQ66Y2ETPtssbOm0ZK/yAl3Ib3+HP++EN87UUWvsiDCEgDjGO55X4xfFP/A2TOpoThAMzZwMX
0pcPV7Xdhx/QQ3xwHJ2dmDVyVeA1PAatWos7hY8whRsfeJgDyxd20/FnkEBhNvUQo8r8oCP4W5Mc
crAkh0N0JQJ+/nay0gMmgs4ekq+khIzeVBxpl0qObIJNEjI9f4aWN7U2DiqluH2JcD9bb2KJuNF9
ckNPaAdw8JbD5O30qOuHg7/MxcFKFcpPVdL2Yk4Lg3YcJlMnrrCCKBeW17/u68GY6w5zsdz+TTIk
qpEr4fymuc3uL1AnfkZw31QeWie+iblj547ogQnUZV5TuXC0iP299gg2957G5oX7i9j9EC63zL/o
AUZlCsoYvFl49wTwQcgWyUlKg7PQdnYy1JgWJ3HV2fyDVmTp2de8ElrK7F3FS67kI9W+OLVpaJCM
U5ufIGpgXztyF4cB9t6T734GzX1JQSDMe9hTubIJkOR3mGz3cjrxo101cLDPdWe5EZ0I9olGbeG6
E5SBAOJGCKWP9ojheeEPQoo+qqvtT2ScaH0Mnn6tYV8TtPFB3bt4QmQcZGhOU4HPVVyqnDCQuhHw
N882tx3kLRbBV8bBtexN0XTD7LZYfmYg7bpxHz3RNwz57axVNM7nbkQHm9RLmpY+N/G+70ZuDLtU
IORzXZ0HLq/53fL1ghqExsu7gbTG0amYYzJw2iB6LbjaUMRtJBkM3OC8dRYa+5fGLMh33SpzfVo6
QAOrhox5y/G7XxO44UJvg14Kj0UQb0VUVRoR32j2UABCQHC9OpBBiD8dVBoNV2dXtMDR9M79ApUs
3grStJp1jobhGHTb8BW/uKNoWdX8H8o2ESV8wJHHuufri7pkgAIgMHPUXFnpL1bw+McxT3yhXAh1
6Be+OqBam6R2yiIftvtNIS7dReaQ08x2q8IE9i11Pb9UJLez0gIIbPCwCf7qo/hv3HcWmVoH6S2Z
3eMFoFyyLL2TYzg7SXQCTZX4SvZWuIy+oQICBCpuofpNzeuNS4VPAgMryNcOkJ6jzgnHvR9VtK5W
UGKOX8za+xChVrUW5RMrsqkbWjBImsWw/CHjzvM4EEEchFro797zWfx6EfHobKzqojSvY9+R7R5f
/a6Jyb9JnUs4OCwj4Gk6nUT9ktGi45TKXp4YZfWc3RJKk3mfmtusaiN27m+CFCTpZs0nCsWc9BqZ
f0jm2AoQ6tSB/441ZX+WdKDY+XqiNnPATuNirIirmTcd2wfjLkUuN/ry355og09abmOiMOrDgzIx
/Jd7esoNmqaA1wiGepRQe1G0AdRueEFVeMfyMgqtYLJ1uD3uCORsky3MgSPOUwchpEZJ1DyAxDQS
SZVeyhPSCwLdzTlohp/xdnZEIEkgYbOhg2jC02TSszd7m9Y2nja2oBNaNUF36Pkul71p0XyX88oR
TqYjkzlBuPo4rvg5zCEmvZ4P/A06T9XipA/BN0/p8a1QJwgoXEm7Ufrc+BKBqxyQ4wqaG9MNdDuD
t2PDw8E4ya+Jd7SDM/GDW5SNx9U2JNDXwEP6cLQ0RWioT8hepOQQU5lHTFXmwtwy4Iga4SkqNQJJ
jDs3Gi/ZIolt4STdKagZHHjBDK1qTRnue+CZtClhJ3NGDjioxjblLkmiDX9DUjAeW5GTL7ZNfrN7
MDBss9m5ZmU2JRFlHKla7YDx+e14rlW9hnzM5o1+waCOiZo+PDmosSLXp3Vp48E2GxBAkOAXIbU2
dB8K9E6sIBHkEznCc2UTHld/x9zfldDsFw+7dRTGnKKcwmDPA0MBwjmqAnNgbBJkdJGPodR39mbe
uPo3s40to4PEMmgbVwo/9xNPGj70pIfRdZvHVCq45V+mVY3kLXlnJOJfplAfGXytWEBhlSaqBqfC
BTjhhb0H4CSZG+2OHVNaKvyszJlBkLB4Kh8ZizIrkCQs/+K7A1gN3+86lcOAd/AiXDREuU3xtw0g
aPGQFUjDWIpx+bC35CjASJ4Guhqe7nfbfVI28zaLJiTDZG7oJi+mCRrRGmwY737SeUdocunsYjqP
zzo5GXaIvTiBOHjhUgZbAkZa8IqJvFpkfU70DkuaLwmgMT3a4a3DK/zytlduF2EvWW1SBNH0/d/m
q20eStXGHPxmiTc5HwS2U+AR2q2UgvdBiU85hYlbW5aR/mES6eR3de1RexpNLWuPZF7xpy+i1zRk
B216fCHIPUGC6MPpdPlhJ3aK/FwzrKZxeMANu+bzNtcrdASZ+qjw/Ecwt8aV+DvlJOxxNHc+7tBs
iQ+gv/xAUvZgBNJnJ4HyEzo/FT0hbYmXXsY+CIXIpGuT+PKCogWMcxqCUs1qeAsjBbM8ed6m1CqD
lkTUo/RH8sQ8biC00Mf6IsntsVVZvwy82yYZjBjd1aM51/qxHbq13wBlOElol8s6FMhiWP4sDspm
bmYYZ2AS81DrTRUk7+P4r+Sjd/zdMd1FWS2AR+Q4WUm3xSUwc5MFfhwDYQeBuihskVd+qeWwPfv3
PHBQKCzqV2v+YmDD2i0cnP2dNJ4XZvGAPP0/5iHeRiD9c1KV0ShL12PPT15vF7O1jqt/Qvnubf8o
pCqdaiHhyUBVekqSMBm/l+Wf8t2Z5gkeDP3ZRnLpeXnYup2acccGch8nP60BPFWdzxV8mJgmKNte
qCSV9uak5WRZQWALTh51c08R9dGozvNKJAbAC13h0urXbn8EV5dizi1p4XItdfIBjIFY69m5XY0S
bKvetVr3nvhu5oH6HnP0HdbkBQrmFsJxptvWQi3t+g55S+lejxRPYeIYddctX2qdFgZoyC/IUBO2
q1Kk27RCfDZhPHxxF0E1MBAO6DX0DD3rDL/DEF3VQ8IcdUAK/3lh0YJ2XBzJc9R6QXM0x7NcB+Pz
WugA912PY8rSHVF6GBSV2/ugaUe84fg/EfjgWaBIYVkwafXzd/irXjDYXfrgi1pEHQFsJjafvQnU
0QQkjv70nP9PkcjHA5sppWb7wQ5wxZWJcmroZ51GM8ORfnks3JKXJgQKlv3PGz+vLLXK9gF5rJ0b
a12WfHjGcfRZMdLvc8imjkSUVPq1yrgNWpClWff3M3KxHkIsNq+5ZWLRdXFj7y5JIUj/1ptL80Pg
VpOsIwpgQpHTzlPFBygPIN7nuYr6WaClxCsGrJLU7lZfxpl3c32k/RVDAb065yx/XR7WmWqt/XEt
QuSuNHtN/fQsKGF0cRho+P2Vahw+RoVWXtO2u324HXypvWRkCcQ5iWdtQquyKF0gRpBzUSkvMC/o
PhhPezwkpJJPKYhzTj4dHRBWzRkp46mOZdcmZiZ6PnfDUSdGAHk6C9NlI14IQrL9QrBz5rs4PKM3
Pmgq8Y/+jnMsaCm1GJ2G2axh64uDRsfJklGOTGAgvv1fHlJSGfWupaMpmW0lssHlBMdfO36ANDKz
F3VoBPXYcG7sfK4qnx7LFsU4fGoEHejYUsBpnn5gq3iS+lkmQablMCsmaGQjaH573SReG+1HOCKC
gpeEZ/8JW2CzM34mOF/EOPLFdSEuwmMBNdWimCY8YKf3iHluR9CloCEcfpysc5mmc/I+WGW8RKcv
mWAWzm4WXlAV0SMP0jxSV12Ws1+nVCO3mijsqsauW1uhIPzBH/oq/B/Hosd0AOo1yFc4ENfOGswC
9mKh0lCqvXE+t6I81n5zA+hSRxyEwaUphCnv+wnlwjiGdde2sRg7+Enyg4aYQCVgqLHXWfr7BpUc
VtgWMbsFDvaZAXwGEFGnn+piqLdEDFkc9AkGqaTXi4nnRMiaxQeGVG7rLp9ukeCEXC4cdQD2Rbml
4DR66G5/eDgioggft3A/gbfP7pjaZMqZqpfGR7SYE30pCdpe4GUgS7uHCvoRsanEPBLKXR1PqBwp
3Cqw2ysS1pNKEbfoArEVbVaZWPUtoRC057ix9xFv0mEOQ05wvSNcw/ZJtE+J3DkhXJ+2KwQM56Ed
GOW7lNo5WnE/UNgFzL3CLKHCSvaS3Zoybddyxgrfl+P1KiEqzzM0rREt14NaA+i/AjsilZlcY8gf
EtsyZexJ5yFhGx4bgWHSmmqOcHnN3I9GQewwtz/gYCKgVDMHhVN+1Q1E6FTraquMSs6QXybofytI
RuT4nzME5QcCsMPqJfvkjzYr+to8JXUJmmK3ICw+6c6guu0UtJHUP6HytlewW3GaDWSZc83Y4L0z
0EXeM9FjEBdXrqlJntOjGUl/TIb7QkizDfNGe01v6jA8wY0JYDII9Wg+3srJzPZEq5J2j03S9wtO
g2sFJEFy1bNdSMhyGqL+GuXQJ8NgdeHRUe80gm6eycuTPH+O0RhrRjT7W4UarW3A4cOurZVfoP95
oJ4R8kxbRBf5XDmj+MPMegvck5/K2P8nZZxaje8x+ruBqVa2ZVW1VCMICV0F80YVY67/csL8rHnm
6IPK34K3y9fWMnoK6DI3rhDNPOs0BA1/MHstGw+zuDF+9WWMIyQ1p5GmnDaSc9jV6+IctgSt0Sde
2FXiT3kTYAFDCLRhuw8SmfQAtgaR6BQtkQUU+VmajzeDrM7F2FCChpCpJzHm2VYn/6W4GjdaJ25e
L9xcmnL38ig5NNxK0ygnFhAtaTGn0TjhObH8fsoczIlKj3HUo6eSg6ksGx2YoPSqzPx0BQW+YZb1
vVkyKZx4KF37u752+lvAj+YD0UvvIrCoZ7O3xZTIbhNZyrVBRH1BwUcDZgP2ogu9dmh+N3a6n5LD
VQD6GyEAtMUK2xNqAsenEGT+LL9nOp+mDt9Y8Zq0Rn6v4lELspoqOb5D6zYmdqU466XuRftTuUVo
Uk8+ckTi5PT6i+ougKde2SDocT6hg+vrqqD5th73A2vkp8aVQyH5/ESE2eGUvuRZkb5o/uYDfGOo
Yij891cLcoYMLbuPAe2o39iaAz1L/gFKpeSJQqkDgCn4SDbsTvF3frGeMYFkg3DO/mctU3M6H1M8
G5krxTao7pUnoqABjnKpICPe9tpMDn3rO27VKdL61uETmTKiw9+aeuwADiAZ2LMw+8Vz9Tw5YXSE
417NlSBu/+97C573swv9pD6PPKN+M2xyHC9NsGyAmz/B5VZCQHk5biLek9F2LNlrkCOIUQbPAa66
Bdm58+hsznenkz7Fvb6OzELVdG2ZiINBZMAVJm4EpDGcf+rBhZM0BPBvQjCBDK8+utX61mboRAMf
rpOBGieZI4l2/AsHqLfNfQaaVXoyDKNcRLFQNdILxHjNtdTXKPVChjCybNDbC6SXMyOPGLuc7+qV
P/ExyVeAPjxdKRA0bw5qLjWysEYr7K0HBzbYr6aFRMvOGPuls6oFFY2HYc3ozLscqjAVdQueLQ0u
L7D8mOVHofE6opj3/PFj3maJp+VCTsqORsVrDFLUEeEgnClAToQdtU2u8D3Bj925+vgXlTr0GLUa
+noFGdcDu0YwxMN/58fwiBiSUZd7FPrx3loCfyAL8gYWaa1LmgFpPKiscjHESnRObmMqt/lcdoNf
qqH0xZsppVk2/wq23Qp4Y9dwZkzxM1ChIupZWyYFTPtZedNreD1brhUcBYY4w5h1kYB9qQwcROcO
NWnU99Yepmva3R9F0Wt7NFKt/YowNznytQCEJxiJXdbak8rhmIAIlHTmfFbu4871JllqJCv6JKeu
o8B3VVuEZQh3jRBHu+cznsvVncAuLoaimD5XP/Ll26DnNLrAI8IPKvxOYUFtaMjWF9K4k/X3Z/XU
YYcnL7JKU3VxRe1sjZUJcZoKKh45wzIr9/7d3SQS9wt+6P7cfsxn6uGSKakR0Q4SOqyhcnx9Z68U
vCLm3Xp/CISTcXmPZpAwAP9Kh2jHC2t6gAg1QragmPDoF5c4a0TVWUmyuTH5YhaP9xLtGbWb3RBd
6H7oxALGjcLTteiXz58bBqeJccIoo2htulNnYEf7dKu08NcOowk4e0sKy/y3hydlG3g6VcrJSYRg
aizV2K53LO6hnqM1cldMmFLPtsf7QJ++LCUdrRLnexqm3/Vj7oKge4b0exiBQqyWOjdVRSP7JWOU
IjvL+iQulkj763ScNWQE2d2o5vff0f6slUJPJL0mpmDWPUug9Gi7OWuCYNtI8XLgK1mnikqckyvb
/pVJVJE6f4SXhaDvae72Gqa5rj1+Qr7COzqqLabHsZyyKQEj+X0M9mfJYwH136TNZX/ODQCC+h2G
Ina6++7/AqlWroDqAcaPFzUpd3vDWYTz7XLOnMA88Zxhu7xFQPiDDTq49GvFnheSEiueKhHlObxF
Gdt67BNdo5R5W6i84jh1aAQjPKRCeISWuklKPqgYZtIqHb0ElZCicx8dLUw2bcjZQjCYunW7OgVT
32buhMCHVgm0Abj1AcbOD6kM5QXt/T7vvhkaqYOBdVTDocijYNh6Ni/ma8WgMqxYyD+wz7pxXNEJ
RE+C1/AvS3fvSXFlBndILVqkNgHTEFbpeEllW+R2acM6wzY9OuELRVyOPuhF/mLRODbj7ZTXotEE
wUMJSXHLXpF2KXUuAg3iyolhUWJGaUUb+BfTCASw2FI5sDbutdPbeqTpuH7c6gSSviBSYdTYEE/f
Pf93+0CY03dEmxzjXeCiAqvuKsMMbjgprunfdzrH9GMvortiqwvsiSRLZNLjuLS4zBjKAkVBv05T
4bbncjkwLdkf0bqDvYrw1OmSMoQUfi7394TxfLvam6f2lKrf1B5l6o8YA+6amrFgo9GArVQg01vo
eQ+1EI4VhutGO6aUXTgOT0KIBH51u07ECtKN7pSKe63bO5S2Rjn9IQemH8LPzKffcrFt9SleFGN0
EJYg1qihfjSwul3sXlWM97+LtZAf+pNanx6s/mOkaKbez2H4KrkvJFT3aOE5f8PJUX5qkr3coSKW
qypepOpG00iFiXtBokageHWwbaG8wx18dNeExZING6CYJ9zEv7AcQtU5hvTuQH3Iij/WXXr7CYuA
m+fgxaSr0PuGhlbYBgh4fhh/C2ydWaYIbzN8fYrkGuc3Iey9B0VOOOhTuDSvrP7XWmT3G3j9NK7I
wDTpg7s4N90eqfb9avX90pGQWnkhvR+tsQTdDEOtj3F7aheOTOEDzmhiBzR8MM5pa/Pa2pOgppJD
GAbLyfc2q/beOfWiFDjimCowGUevCQbZe6hrMd98bHcWAi4Rjomoc1i72aidtMZNA2pX37zrMwh/
Q1ElCGS4cgi9g+TUbo/jzTjz9YaY7zcX4BjCh3XL0uPrlZvGYhW1gTLWILiQnygdy9bd3yo2B01S
q8aXoiRqTTtW6c3eXpbCJZ6/Ye7pTrXYzgTMBOqYh1ZDJ+jFzCUjHp603smMQ6Hy/A6cHJtxUTgD
b2rfO2cmg29lzydwuUQ5vgtibIbulKv8eCGhSsJldjekm9nGbpArOkafroHeb0GhQ/CH/GqUu+I/
Jq3mj/yaAuhQ08njSBy0I/YrcXfe41tl5BlE6IKcjeZu7zbPTC/phA0B6HIEC2kJZK5BpLiNSMhH
xSwSlMbxZ1mlNVMu1/VnA1bBWRjoP1dMFElM1H0dcJPPZcMm52cbBv9+1MaT/RiM5vYnBSQx0CD/
SCvuhvkTrlrlZxnnApnf7Q/CmvaG8ATmkdr1jNL1nKFFAuNHvGZbkNCMWybaWnx9JWkDhOHWBLlI
NfD/FSO90QNEZPvF+wG1L4S2743Je70OmeInc08JXqonUcIoboBiGciyu0M5PtSC+Loeld6uG18U
SJ5fCCRRoUKpytrXZrKPHwwJpS3SjKqNYjGGGPjnIYJZNt9E0RSCWbiMCptLu3mn2JWY8MDfMOIB
RC4gHmAutCc8kGJ7ZgRF1pmNcjzsJ5OdnwwD0akVh8GMwKYHV3jX0B44Q1hw4TeCNPp/5hoUAi2C
G32bSpJrKlnfnDpD13VzXswBYS/qGVouKWNhA5REMY1gNi3APwTfE55c81+9kB0FgiRTUIMHV4S3
UUWyCYLcwl2PKYsvkIfOzbUNkLwOqXmYbTtSIjXH97Dc1m0bJCuGvwjANMcF3r546LxwLiPYfr2s
2ZiSROxrHfuA/jqJNfRKyLXrFW5ZM66kCoaDT6iMj78wugjAfW4yxWAcxM7uo/nqXsNnSmKI9B1Q
ANzZwQ/GAoko+gzShYcYUi2D3vaYyfIhNj36n7GbxstGLj050ng6NFMaxqMQWNF7rEYltjM//YF2
P+daemGmlvmqxlNc79sV+yvtb0pxnOSEOyGWLaiDRJXEDfsJbnpa2knIcu1LeJ4kmyySpK9EgRNV
+76ZnqGnH1lu5CFcEjx0+a8CF+vdbAQow506g8IXy8+VxUDxRNLg5gyb9Puq/ZPfaszhgRYr/xsI
zUJRby6LBiSE0Sfv+jmr7urXV3W4DnaMyAaUG/sA0wZXIFJ/090x58jq7LljO30aPV1vcAj6ZDbd
+mleZplQlSVwc9HULOj5G7XUdhl/GemVRHn3WegRRLDVCdwGhiZfz6U92d0WtngVPgt+6eCUeQhs
eSZtZvU4C40zK8X4B3m/FRlILxg5BrEzLjcy4gmz+d9tVwa93OqNWF/SCZI/Tg+xMgtzM9iUn5I2
aPV4UhbRaYcjiwsMy1X3AKg2J/k8JZJTbJ6WeQ9KLWjeeQ9SaOvMThRLpXJhLEGI3SnuFbBwfVt+
0/ltkDmDJoTksDICha4qzumg6VzS4zrkm3rN90/i6c0KFGp2WWxC0oO0QB3o0t6ixPHW8JuqvFsw
PwkmKTt9BJy8MMCDIzY8R2RKrZO2+KKXt9oTTXziC7k0SjAs5/1OZ70RDCXBbU0RAMqurC2MBvAZ
X8xd1nmSmgFh61yiwLJQvI+YBwu53eW0i/zkiUzcXB6Lj6hPWBrhTiB7Hjjd2W9/KlgABTE7jyjD
P0LNmyqNwCuNYw4XiJ4SuSeOzA5xxrT42wW0n9XTtmN28tcliqQvJtrtv6MBGxhqxuRsF6qTq8A5
8TYOeFPUCjouIcNyXN4weeN3fBqZAJEJhtgXku0K+yvXrvsnSxvgyQMF9zdq+XpPFMLHntj34UCU
lvdiz4a6aJlWEQ4k2ciZhyJ8cNKwV/EQ+qKUPBL9q+okFRhPDNF27Rr/VyMSFeXlNjEmlhKQmTYC
xjjoHYd4Ahc2g60OMuowIukHy4ouk5Y3SgwzOjCFGQ3iXOfIBU6AZ8EXXMh6mTFfbstH7pDSSm43
5qQ7W3mEfmOvKEPxgk1U9ubXA61n4Z2K+Zwn/N8PkhNFKIbAo/TZeR89z+prsc4wAdPNA2LppEcN
BqldMAFJ3y0LLiq4XmGsozW9LXwA7ZNjGHMshUgKoSJNKWWXWeJo6ruZnkzJ1QpVomNC2vBA+vRk
UgaFlxxm8HDYDKAwe75zk1DBSVeVc8Pj+E0dbndHmVQLDQasdD7d1vKZfHRuh2h1JSJDzG6GrRzI
BFsvW6KjwE4/Uc2yLfkUznnU6uGp5NN0h2LmAUwYTPAUpxJ6txPskF9ufyWVKSDRWPHP0kPzF4fQ
BhKuXXIaNMcBpp86IV0ff8FjVeDWUh73iM2whZQkDp98Imvvbasy1RTb+FyIAyX/ps7nNPvxRnU9
woYamtENhg9xVzUPJTiY4iR4v5loDTme3XnQofsvRYi71h4efU3mUltObYoT6gyHnNMFNnKN4Ty0
i2ZR1FbDOMemwHA6jdjzrHtVgoyKt6MgyfE1/ANeh3Q0R0vYZoojtZaO+zbqNiHRkL6+ZB/O3PFH
ohEh9J9ptvb6vbcZiV2sbYydjPKgRcF82UQv5PmUPqZvfePzayxGuh+/96fNvJwWX2yur/EpnjvC
QxXEt2V7eP0YUIxcjkED14MpW9zisyjh0XKvxQou1VZw2PFEhjMLqMEOhwT9uq10ZjHL7tnaj60R
0ghqN4AEwCwciaOf+dhWlWGaevQwByiR8+LS0gKhkmi/11PPKcrLlkx5i6tRNoLiyyj5Q343X21X
D8NgOyKpGS9yrlX93mBrwuBev/Hu3/w4R6yN7lMnkkbsdkhPRavK1o/nCz7bBFhML9f0kKjSrZr6
yOPNkM0tg8+ZLwBX8jK9n5xqd++SG2eLqQpDdQP3PRac3BvLZnsDWqlecXQ86rJsWfhCO9f+JpLT
VnenglbZDyXZ6qApZN0+6Ll/JQ/s0iefPG9f3CwkQpqe/CRGu3WVExIMrdC8WVQwey7ki4Q9pVcD
cBmT0FzQxKQE1sOihelBZWD66V/Mjbxah9+ID1MEkyILJWk3KeCdUPCg6gJEPdCSCnrNv/jWT4CK
wwY+x0+HP5ob9VAtP1dtHqPzY1fJS3bD+2/250Af01SaRczCAOIWVh3n5h2tTd8frDJ58LzEnmCE
0/c1tvM8qHb1PxS1/LNr121LTVWoVGs79LH6e9xQzUfEgnpuePpEX6IpxZ50QHfSxjJw7tRMNPkk
j14uwBpvzYF0g9LhSM6z7rTynw4Q/otGNgupaAisJl238gkiCgYMpxcDx0ra5uH6baqKiyJGOpKj
CoQZhaixK1Fs1w+j9YBBESJ0XXviM4MiDa8b4d1tjWhX6oaw8C8ingwbeEJIanoOwmwMIR6ok4sF
Q8jxsRMI7xHwVtH8UWpD/8ZZQ47yZwhR7Pi2amvhAeiYG2NsXaTC29aPT3fvc0Ioej3noiWe86Zt
cJy5bRazn8aUz8RE6hMvG6o5Epe9+ArnnUkARPmtAS9/e6RtCxokBUKQH4pJ/WC4x4x8KchB+1lY
Ggj9blp4+3IV45eLxVt3EBk4ghqGYp55SQjFszU9ahzH4d8L6G1IlKSDr2HsB3JNrby5VB9Jda/e
enIcAuY/xgb75QXl/DGKWaVNDy10sg/gjRUvU55RCJg2XYsnZwe0Hy3bEbsi7Tnb28n0l8GLzVIS
smGsfbLaPN324fXuU/9Fir65aTX1cS/gaLcuaLP+xw74RnmMQbNdafBSh9iZnkJd07nq4UgPglMY
J116/KGwt2UyEnpVkWks+s4VJW2iJxj2ZtKcb40F2+tWHmVVN5EfxemB+i0YbRWsgcQfb57hETzY
23YgAFaVTHEYkT2PLuXXlx0IasoF/7ZWryg9ZkUPL1ei4l9QDy7rNdnJF0qwc2ZHkp8bEJ72SipF
CFtPemoByq6tHrnoMa+VEYmL2/pOrittzs/XZWPPzfdmQ8D4Rv0IQjS0Af6RSvjjwo3ZhFDNHxDm
U48LQva4IzSBrELFIaPxJc/yG+XB0LFBCj4uVNQZ7sllUMtgNz0Gkj+ZnraFtbYQTagkl+2FucDE
OvajuwdI9DlhVRGsoJquVklgpTRhFENlIuGvgd4AT50gkXbGH5m4+0V6J73eWcL18fKHqp1cAI++
yFoT7dEp0Bvs/j5Yx4GxOr0ZpQzV7D5MLGHSf6D3e2q2+9W5GzPQn69t01vvYbob3vBT/AjHs7tQ
IKg34gUGGifMmUJrVoBqSS9PhChgRjoCTkeeRJuTiZyB0t8l8MQKB8Oj8QAGTqXNXPnQipCihqoE
K7lWIpW0WFo8WT0YTlX7e3rKtE0WvYorlhBHmkrUB3AXrTzjoDWnPuzVenmpyYoGKd5Qt1ffWgac
TaoZrzt76+qmo3+Gbv0LbeZ8VuC7/y0ymOcHmjFOeIM/99A20rweggW4uuU98HjfmyMZNFUbAZMK
peZfvs8s4wF/cKG8A2MWM0A5iCCfruHSKjSTLzn5eurdrDRT+DR4gHVReiD24I6chgTueOwsH410
P/cHvE80A0ydkFB6yMvt82vjDFz3tdRksN6gy269jgDFvyg3VAM+iN7IcEZZaUDmVveej/Gm8ihB
Y2P2+i+gVmoOour74txQ+FSFjby00ZJptTwWljTwxiVk9XuGjmfC7sPfOgRmRBGceG+XZAwtpkgY
mb6taDzlLcSHU2V4D7TGnjrwp/dSUHlf2Q+8r3P/7IfbOOTMVQe+pSkYu1fIVb4KKIT0MnaedIPn
7G7tlzJbcjtzEGmtwGCXg561g88/2mZj1xypeQHgJQVZjOEtQdCR233SgYd70lnj1Vo7MWy6mRtB
/dkQxurA9PL5Lj+2FY8JFfMx0fDyZJSeYt8cOqmQuHT6YE73lKVQ3NyYt8SMXdQpSIG+ihoC1xu+
gf2lLXcrLebuMhVK+aGlZSxbMLRJ/I18EFx/aCft5lkoM4QKh3MjnEvgIO9C9h7WovmgKbucPrQ3
Q7MZ9PLNTpa59AK7nfy2+JB4BbV9mxYKaxWb0guyHM80wH3m+5xTc78QMrddc0qNUMS62fFrks36
IIrBoecPLLx7YGv/9V+Cm6xXdzRfOQX8vkwDWevH7tkoySXjQpFPXDnkBxeDti6Z9RWwXs5fOK8D
uh8XjnCoaiVpUxicXXVkrD32PvpHEFnkQyjZOOolC0h30bF8nIs9uyBS3M8ikx9YLslrSFHAGSP9
ZF7E9mUt8OfRHuSrDDPrsX3ZZgfK2QTSEhNqqPoYuVZGUcuycSNov9ka0m9SAk/sc/ilrs0y8l/8
2QPuhFyrVvPL+DNPFTVEcjtbaENUTRPgCYcBumb/OzS1G0K4kAaCFVlbZbk9oeUbD5Tg6yPyri6/
EfvHeSHHseuNu9qZc3fqaRvywa4RINRGw6+UUHwFOakkXr0mAOP3bfEtJzIQVlKts1CApGRgOdVp
Y0CEpX/CMb0mXA9Uc/3/BlcLdPWH7NEvmpGIM3bSMdaoAmb+3oijQ28nnC4gQnznMCV2tjSjSaOX
f+do9Qs2hDskTnsdO6b4Rf1E3FMrM5diH5fcovR/KSX1n5OewTqTyVbSYeNcqohIUQbxVOU5aYga
ogJiLSdfBAmL43K6khriFIjyQeC9/dsAYMnHtWrknhvzNE4qG+ctnhtLpPhOY+O6FIPYjvOsLBco
bE09pl5n1+TDShqNuLzC19D7+Fg4CMDk+524p60G/1c6HnHGszrnnh5BAITBc0qu5KNpYDiK7aAz
PgjgHGoxpbYr1vpheX7IYebBwewNfGO5hPVi5KBN5GCyE9DOI4ZNsLg5FLQuegmNsSHAM9TdE2q+
wJ6CqWuRppIugeiO7265KLGAlBpV0/Vl7/O+iRDlWntmP9QeTl8TfVzweLsyLG5v2CkZPjGaVPmk
JdR+qNwf9CR3nAF2iA6JW6oNxaeGl+C1d7SLRxyVf/PVxsn1eXe6MfLJcWc4Uy2mPQcQ6AHL/SLJ
nyvK6VCgiq091GH0PJRQAyGjl/UIycjVW0UhgMM91OYRLxh5wlfGXuLiQYVwg/IyMlVEbkB9DA6Q
Kr5ukPB1UDDiFnoFwWdQr9kRPAILRX3eTYyIsU7n28BSN01F36fbwv+u+rOS0wrmIiw+5tzW4Swv
iSQxMJOcC5bCLiRgttpO7b+z6ZJ2/bnA0weiZK+D+Jfui5T81kacctON71UbPva3SXCiDhReu3Ol
S8qRZWgAdEaYe1aFTfwjA+15kGapgpcomyzxkM00pcMRSsGUjWLyUw8qH4Nw1jPKF0aodciCzH+8
ZHWGqAIM1dR/4ior22bgOu43m38JCjtZWKZvb1NE1j6l8l+YDtKQ6VNFsOkC/X95puVxwH6ReWJ9
JDNCeQoN3BvdwNkxIu+dbrrAVaPUTGue/h06NxTQj/y1v08mMBur/j+TAuKqRO1jmqQfnGSrCC4s
pvB/jfOrvnU9bd4SQcxhu9Q9kx4OvTva17yZilLtaoIPGj4jPDMJLN78iXk1MgPNnFdI4R3Jh/WC
/kmIYpwvKGg+Apt3ugFi2T9rENjs0fl+rCRg3CSphBGy2codNF4oXpvbF42kVe2/tkEpjNuhuaSA
m9soM4pQDhUNaK9Ab5NmjfKhljyvAyuL6G6LGWzksui+SJoxOo9ZgV8HDzpN7xS8Te4JKDY5FoRm
YQtPBexL8WR6L6Pti1hUVTETAYEgAE7BbZJWtzATk00CsmMWNFFGM/f23PlLLXI3zB8S3azUazUr
Y4V7YScLcs9TwXg1mVhMdmV/hCSJADNzkW86UmEMm43Q5kYaIJ8xOzGaYzxUO7bQyVY5EWQz5L3P
1TqDi+oTVt9xCxxKMaQMo0iVwOILSlbWLI8mzuhvqCmYSw4KomuoqdOJB7ftwabMqxZGRhTPrmAg
jpHGCI85S8h3NGjReIPpVue7a1cmWWGnIEbf7pSqFJdg59JPIAcAbVQ07v/nbfndsj7WmecNAv35
IkNGpu8aXSwnON9vKFQilelCdNKP/A/HRiA6T6g5nflfrCxW9ebcAXMPgAB3jwvccOncp3jHr5eM
zSfz6L7R7oIhgo98renAvVVm4RIBLQNeJJFpC671zpHcgVE7xJ04ha6F2W+j2r+kGmi21N+DLHaL
DV7YR3yx3NGhvC66k9MFjzhNB7DqoqhIUG1u86uBvrq2GNvQr4NPWXO3Vv7Vv1pHu9oDu29zyfzT
7fBxJyQ/IRrJkka4LZSF+5rj41k6xR+Ci+G2dtf4pjM6ccITEc5bx2g65gJC5MHYRlamiu5/p98c
vZgCjEMl4uLb88ZSpxlbYuCh4g/QjrEpUxBmm7YzZMC1qcR2W3q4bp30YlyXEAZ5kxrb58nyHXGK
BUTXhmltf1J90Gap2ylf2uUwC1KiEcPJC5YIuJe18Y0t23Eq1p5TeogSEhrkPlfO/L4uZ65UsSfv
2WxXxXcgn7VvDhzsSnS8gAgw5QEvE7B8xwKm/NEkFXe9VXhzO/JSb9BH9vRD7djrzMk4RfpyxNRf
JT+XhUl6KNwclXMGA/WrvLIzsInnjRAv+mCFhyugX0YhWxcMCAg9Xdjec2uaqb+OvN7Z1uXpf823
mk3tVAyprMSQcQ7sfB2XeseGuMBGqd6nHUKdJf1Ul4lrekF71hzXipEkYVDiaCeXaYoj1Nm6uIk/
0ChILKcuHYN2qRgis2u/p3d6U8DtQLU3Z0/Er0QhsHSA/8F0fiKcA4m9QBhf8E3ImURZqEge7eMj
9mODYkDpZHyWHRbXy0OepPz24pF0lwljrKPEaFBBZlbS52agwyTfjyG7JfbsjkVmkKnMfCoo4+HR
qKLjziPM+3+IkoRJ/24mbuu0+utJXjmq9eOUMGegoGYs6cuWeEEmjXer1J5+ksPrKTDKv3c/2Eld
dUhTVZb2o01ytWaR1Wtx7JlXIhVOGhG2P1ZnvzdadMQe8L5WCB1u1QoRwaUqAqoeEIptdOtUkaUu
3AzzD1loS5kHXUBXxBOaP7Uy6yXXh6RB6EWG2kBi+ztHHnvGW0zVXtVPHCRL/+j2vTuIR9FN9FL1
N0AtqNw5z0U+V5Kmj3qqQCXc+mzlY1aOzFW75amBGoVXaHdC2J0fSEzqDlxkR/CATaVag4PZ77j9
sgfoGZFGK3gtNe7Sg50ae8kHhDlYQDpn8uMGbc+My6ZtxWIYQhWHkjEh0DXB7HJwF/yKgvhpz/3g
Y2BPpRbM/oI7zvtE46EozDYvQDqHJlH5raBClIXMzrKh1RX3lW9KBYywKGgrkshcnfhHdDoN9wYV
ZHy9FofL3f3FWvCYf5YhGq+Gd0gMhez9tVcYx8pgAGZ44magiLntNyB9G8nK62O2S59kF9TyT4rB
jTHbvuIt+C7MvQfJfAM9NjYDoshHk2lsC3FBYqqJ2h7nB4nAlwUMRKaUyiBw3fSg8mXF/iT9KItx
0jh3dLOIxRiUtzKm4ha7jeZV0aZrWIeVQPGITjmdl8OuGkdShh2ieGp9X1IazowwShJe4CNHFeUO
ePIvkfMTqJgHQLKyUV2XkOhaxPzaXhj8CY77hXGEILdyL7+g8hO8ai5FwE1FVd8dFGL8vvt9442w
U1V5FDXT853i3+87OISWYrscFFRs09+/oiMWGFBtvNUoDAPJDFE2JNjjubkQQZjZSyHZifda9C+G
e8Ow0gY0HnF1yCl6q3WKsBl4spWhGcipffZJIwmv4OHpdA4d9jRa8JwG63fx0oTQdHjewE1IFy4b
r/2UpmoAtVQhfiKuqMCrmRv5TilrfW8VZesNISzv5AacvviYyQnoJbpTw3pkMGxMSr/9Ql5D1Hs7
ao03Gbq6RJDk5pxyyB5iW7tg/lNRxF0a2n4ReYFWMni4b4EV3NYucDwQpumLPD139MqttW69/UWG
nfYCtE0g5MLuWaP73joywTjQq1Vu7TfvFlyq67XQ1k6hDF0gxYp88+5sAO6/biQ5ZvxYC24pVQ5q
VGj6m7WA0zbQp5iJHvB3pp2YnjEbgJ2KpxEYXY9DvsEQWQWy5hNN4MAE5TVgt4WAGeQmWyivFE/1
P8OjrhrhYHaPCJt21emEqD8lMJi4KbaBxmjhKJzB/iDZUqvEh5l0VHhv9G5g+/Y1eIfZT3BpmqPL
GF43jtel6sx5iv0qJSljPrMSKHeLXNhmQUu6JzxTZUEM5yc9c8GTke5gqIIMFBcjELjPI5mB8xWU
HWWSlryD2mwStCiMFx6LqMxuFlCcKgyGEFXyxaBMmYWSK/eDQDOEGn5saEcqngbhMf9zrHbpMMnh
FkmSvkV4yZfrlLW9yzVWeLnf7500qsBW65LkOSFIEAvis4QU5kn2hy4OTZIOK8jSAzFnHO94+kIS
/2sFKC5IMX0desO2gTC/cWwlNkvlwl/vuwAbxnyO8NG9JKlcFZ7Kx+aVA6dfC+5hlm/tOXi7fIRA
6eklh35YjTyvMmaqhSW6w7AMWwty3tMDlmsI1XGIEOx+duTWkEl3gHoayczyi300rw5X9IvRB2Tw
dHjpFBCapgoMJFu0I4O8Y4uOxBLp6VF8hOf4hT3fIqQAo2M3H+pXG8jBzXRuPHyqsy4r3SYv7Uwi
3mNppVCfxeZ3rvpZLGUDAM+9AGE2d+3BhbM9q4yD/+UxDfAK8mNG/F46xI3xRpBGpgvoRYg6W1P+
S3oXQudxTkaa77WV43D5mrWreQ21Gu0Pma9duXoOLT/ylHNUbrogtCxLDaZhiPpUNJ8tP36yDYBt
9DbtK++FbmaQfgYUarb1cBMIvnWTfkoRabZgut24PpbcG3WVkPahaUpzeSf/v5QIYgpyIF2xWuCA
KdP9NPJYGqEEaXWLcc2Hq5n1XK0+btlIpThipZOn8Bb0TEE+836fepOXMkcJBJmQNYS8SXu/ftT4
QGxlWSF6/NEs6pwDNE1pRcykHpUq141nQSKEwS5ikm9dWfxp56hEsBGI/3et9d0aie7gfGoj8sWz
X2upWiLlTkEN2AWDjxHlONRWZnLgULy5iC/ljpf3mbCEJfQWzl9ZQ9xx1LenJGbeeYpV3UhkQPwY
1fS8SN6TbnTFMOiLoK/phd7P19hzsM4RvSfWcHuIeiMotLxzvL5K461H9p87KH5Rx7h315mnKisV
1+7kNtZJKtQ7HyjSqGemdAerMt+xpXFpIY7Rgwo3pfWnYAtGR/lrZhtn79eRNR9OzJ0uYwc3k1aF
y9yxumtAhtuVze7xkJvazugS2IS0B9RXxBVpR9Ms5VbaKWZ03iJHWgZwe6iFLWelKzCipffSIXTe
bnqzqbGT36N05m5r0HRNt761YUB0BPzv+ao5CzD9lyH1SkA1PDbZR+dYGtLWfsI+SWQ5MsOGjv4e
iXWn2BXh992DJo1nlGteg3zkXTVMdrJcGLAfgnK8HkIFxapJvStAI7wdz3TdXaXn59J3kf4RE3U3
6dBHHSc3/LSZk7oROweiVo5UM/DpPNIyD+DJmxCVkIlz8PCU36CtCd54Fko7hcw/xu6DsyYHLO0z
ifayT34Dp0UV40IScWOUvBdvqpYY1o5JG4V3KTgIBCqkAqjYvmjva3BtkW17uhZWVr3HFtUwT13z
FjyRPLhNhVfvRGW1Xtzl4vze96tNEBjEbBF5cADyiP6mXMYUUR/l/xEXToagUzWnKSqGK/2e6gGv
GA6vFFcrxfMQrKoYQNw0PJOcqZnT5Bbwgb61QeYx7nlbCQpAfq9GgQAxbeP+6bGD1BMvzvqXLCTB
PVmtpsLauFFG+Gai6R5tgFsTvHW7Fa90rNTNXAmAWT+G2/aOOMNMl1Wq5XhOdf/2SN7EPjgds0N9
vYfjHFVTybUGVlT4nmtWFgI3wF22i+h5VGWxmBWPY/cAcvhGkEAL15RujwB0gZ3nCwiHgoKqF08H
xoD7nUInv6WVbvjbQVwx4oBbyhcdkzulYrYHgkQSYh2UojOEUpqnO6QjF88hrt6lyEhkH95O8KXM
2QZtvtI9rEqcscby/P/3HrEx4WUGU3/fJBf70qop/LYTeJa3qhPpwaHnTQMl8mcGuJB+GGIRyVYh
4ner4rJ3GkTTX2DcZwJgQ4ZbdzVVYaHoKqz4Wa3uRZDygId6tFI/JqiCIt9ofFRAkUrNPbqEyhZo
pCHYTfEubWuXezEhC7/GbWHFIzHMXrSMP3Z7ISn9P/6sG9LT1TEXcMC7625/9uc+KA4hQ2wLvlus
ykHnmS3ksOoPA4ukDSdoHbEHoU6B52sq5Ktizdr/OTj414K8lY3ZvlJHROafgDlQP/HEWXVHh7VI
ZxnIR0KpH6mefGJOuuTa5+1Os0p7lev54bOfPlAfsBijpRa9+aWIyna4HgOLOFc/O10LCEIBIBbO
H5t/WEJqrNLNgN+sVyc1po4tzCtO0F/VH83lM3AGPQsmdhbGXDcvM8XsOOu8DM0GMbwdrNBMLQbS
o+ymLFO0BzqwG06qG8SLhQl7+DxLYXBkIX0Y1J2OzWszELkwqEk15JNLnlLQeaILYHAyLl/6Zmrq
1Ntb8BCKVOmm6jo7wEvmm+lKCDUorp7nq03dFWMH7DlW99+1H6Ms5QYzdhuywzK+SmwLcVGfRJkN
DcViE56JFcTymawRJ38D0ro+UYhwZDnq3DvaJfEbPEigjhvq6ZI+TFget6wu3+bhdbMwp0+/Ziyd
74IONuT127ppYnZ6g4vQITSmLPfJ6G8E58UaD264OzxeuP+BtlBaAvO64A/3XKrqRt5kvrWaGs2e
TPBv6NRdlgRTn+Z2M09jUJiQFoppTn4/VKPU2nCgPm0d5b7rYj7Y8zOSIH3raKDkhfmVoxNOP0lK
3Qeyzzl9d2TLH1W2S5sKgtGeFVZl09T/pj64mJ2XxLp0kzkf9lBn0B1CtiS+35AdB9tnBCshgsUw
/SAbEjKZmeJbZCOPiyCQ4kpztiVl9ODwu/VPtbsmGg+xopNPuHCy0ABmnXdfEHQ4A4JJS28rXGnP
7mfKcOQOz0Za9GTlm7f69MysOK8IhlPlM/fsdvuM4tWYRgz/Ex1refiwAjU5YdkUAdWviWU0MSth
xcFaciRtv+TPd6ZLeZ2pqM8KsxNuA4DqR/IXK0z3mEYNJXsw9zFtagPnWcm7bGvx0ktEz8tDn9PA
EUN5KoSXENUE/qaaWsese/FAI1Cgt9hTwwd82YaWVrv9KbjHMtHBB6ysX48sBDesJ6vK6AEcny5c
jSgCiO4lTIbd12da+reSelNcJ2oHqLK2n5R88xID78dGSUQYNKO6ZBOiPgCOZBO5WuMNkSWWHd2l
7IFTdhySqhalD25K2yiYaC2FfO9dJJ23GJtknZRHiEYuvFtgEeL26bnj4xxY8Pi+tbt/lgsDWIH0
NVrBgNwRTiDbP/UNemlDwQpKZzRRlxLmoN++vGyTuTcxqkjnfTCb3riqYeXzjrwRTjzivyYoQUsH
Tb43Sv1Nq0L7+juK9nyGyndeEmhFLYFSxo7KPR2Nk83y8HpC/Z7KpnioxveNfrouuY7H9d4DA9Tt
V6AOlVjt6tYqXci5/wbOegurkP/M7K5N3HE3ATGRG6b/q87nCvPPtb/DEnpNkqh9Ik3A5lzf/ZTz
+WbyJwREQCsVBZg94i3ZDF2y6WaWKl62qC4VC/VoaJDP3fSKhyVyO+QLQId8IGiW/R66CH3kQXGW
gZAUHj+S97Gz8ylPE2GzPKSIW7MA5+2gmWpfocDIvjyZWqMb9R1eCUlmc24S95+FGXGsjgc+/L28
MRVYhATogyYjJ+lFzEv+ZxfmOfHvyaDwGNhDouQJ7icE3K/UrC1evnG6OlnV1VW0V5HNcqCmIyew
0FnOZdIvwM29+0MmVoVEnkNyKhh3IvdWieBBn4h5tKSUfYJFExEcvMm8FX8lC5WQ+ymFel9IE9ba
HR4PVW26ygkj05FYRFwSv7ZyD2Dg/u35H3zr773eKMwPljkkuO+NzRC0PWnpx3V+n1hkqfDmELiA
TPckqiiKDBSKZW62mJxjlKFj0nsydgvBjf+LQwu/LxeiFmn6vsFki5A+ssqiGw/d6f/dufkbNhAt
Wig5v6tLbh/8Jy5azkW2M7WzlgA4/BgkJna1qtjQ8+Gj2S0gnroY8ox/LC4shjfJ7Tueg/iqEfil
FggEA18C2llN+RmvUjjn8EhH/UVSmPUMQ02Vb8HnexUgQ1CaEBHV5lfD/vBNH2AQZTpeumaF0I9A
7C4YoAgZPEV5E1ZAAhv2bsTRgDBvGYjpoQdzLmk5rfSYo+Hj+NxSVn6X7oGTXhZl8heXaWarppdX
eXLAwGN/ldhLVlR/uNCkSxU0quNCg8eE7C3qzZyuUkuC8Fy3Dn019QOhj6HjHtd1wuoNgFtO3Fui
hARHQYWfq4+8xdL6p58xBO6Q/DrlWa7WvnVs6X493BHdrorwPWovvoPuLGK+pqbt11OLLKs0fzn/
hiIQf3iUoQ6Z6YpY9SClSa99A6+ORCwvepm4+UVLZp/GKfMr+g/8pWlSJarEDmgSzbqFEJ2EbN1j
NdcR/4zL2TtOfLbHI0JSQop2oo8ASkAx5DizXFmWngH7IRbPCArwORBPH3Vwcf0SNFxVwfAp22wt
8VDy+iKikDlGHJefsh3SWvlJ0j3h+Xe+9EDyb9EuoqKBh/JK+lldynpk1DbODxGUWBrEV+07YLe0
QZR8TA+b7YME0VggDLVcfWuitrlnJd7vu05umuwjGBqR24tY6A1KgjC/wjGy8Nh8PPGnbPb4ZTgb
eHcM6axl0czI1Qnu4euPShxMggMPat7elbq5ramb+X4VV9H4ifPpwQOCneW4/t28PNlP50tOQdZm
7zl29EdI7QFTfuY2ejX3ObwN/xbYUhKSxl6jy1B/TcEPjSH7ZnIPcUoz5WdddsrI6W/ooDedy6K8
J4ghk7rKf5ly5vrN1t/A5iddr15GrRHa+1CK/Sjwy16An7J0Sis2lbBbYyllhnnp1V1v0S9bNBKF
yHO/IVcyJ77x3LsLzSI2Fk8AwD74NT/UAHe1L9jSGMP32YiSn1CSvu1BjVLiKDqtxyI33KNwuI5k
78+5symRw9AJk4iBwm0gGkVEX3N2OVwZnP2wc0DoYmKSjfxJ/IC0LXWeepqmp5PKJZumkYcKDhHa
bf8OkDrWVJFjLrpZE5bjE1zcpcgxqw1sUE1hq9hux51i1Hb8L7VcMREOEgEak3zBuEWSb9j+F08u
VCKr935yPzxy5dXwDU0QXhqYHjTiYJq4JVsCTObbBKo/jHkf6LykKr4mac9Vsvft0yqnY6RRMRQG
uYBc9LRTCqXPUsnuVrmwcMImApAITkuJK/V2xNPKEcBcmjFRO8rVXyuxzlCMmkNTxHQGTurt1z78
B3ndsb6CK5dkeZtEcy6GuzObibS/u1F+7OKwTdSiFJyk2SYKYFHTJS+uuqCxrwtXZM9kkQ1PEZRj
/l0fPjWP2cJeETJRtjEJ/vw89UxNAqZuqPbijQc4BkN5+yJUtWpe+FftqrDuAvxv5ZAktKeIgfMx
y3r7UMIbmrQ0XqDrk53rgAh3yyPNc/t40xwun2tZwmeagiAiJ+taWQesHD/2nZxO9tmPAvnIPbei
P0Bjzu96Sxp+65CipBFla66gAvEQ22frJPmLDX0ixVI6gIcT+CQXyDwVm7CRg6+Ru3D3dFJBilgL
/a+9rkOGJpQ1rpxtNmbaCBdV+JRAgcKwHB8fGj3BA7D4zeFpzdxs5QNvexUV+CbtWSthxpF4etop
tdRMo3U0EGBXp5/3dm/O9xutgDdJkUb7aP+MXteXBVHKZ2lxQqGSAK4q1a4MpjQDi1Hmf3/CiWF+
Mm1HHGtCWCBkLzPdhlFIaIyYeNOv3v6ph+cVYAyS1lh9hKRaLIhvl6XL7KMAgc23dcXy1uLzwwAJ
z0wOlCErtLAJchehhvVuCxlZ+gQTmygYR1/Xl59BN0wB/BIwRd8s811zJitGhcMiJJs4NcZ+H8k/
wU36OcmfqRbGyh0rhcPYOUlDnioQV0sssHQxllqeo4i9ruORRTkS9ryU4nfVAjgViC+bxvdJFapg
VKZk2s27ws5nWYaCWVXGrKYpmRCQO3r3SbaD+Dp69UrF4gdUFgSPNfrr1h9VrRom0Fx7g9TCGoPs
eosXx8kIscY/qMXYoGop3ceV9zhoEbnBM9f509o3bXLD4UyQrJl6iGW+GF0YitzH2E7S6dy/4nbn
+J1MQsVGybTzMhPc2hE0aiEVSofY6VAOXVEItfSy6/Fuw5QotQlq/C25YwAKMESsGcgo0kjhSNni
Y1yfwer8+M0CiQHaGtVK0esmLej8MGOJPqFtaNkXkcxyuaxcMiXOtsPsRfOYG9yIh8gQ39fBmNFe
DoSwTJ6AddKyPeAX8AMwZCTNmFdtNO9WdSOPIDWWS902EqYyrXfFDO5D85Y5UY8SXKA99bdKNdcI
fAj+5H3BBCtCaicY1X8brKVQswjQJ1Jci4z90XEaOmAOKHPAapZFEKZMndcTSv2UYNknKUS+rhrJ
YnoOjCdeKRHHuX+yMiSoQlxWeQN7rCouuXYkDpWQQXASa4GZfKsQ2YqoL88W9CISqoGPnRyg4Oc6
WyZTydGIXcEKJoXeW3Sl/k/YzH6YmY4xrTnaMStw9NkhauZeunchWMEDB/4dJxjYRg+n4NfrRG6M
aF4rSSgtPkawegNsWZGGUGFlmpasIUAVEW4++9gYl3qHLHHx/MXAgp76KivUA3fs+2VlUswS884C
P9k0/GbyyUGUNpiZ1xhpcbmsEmIByggzTFvr1s5dZs9U9ugHmxm2VYjeF33o+PLqkFVWhPY2bE/g
s5Dr9nzB2a0cD3zkYXDScyw7pGF6aayUmHbcDlmVCDRdyW8SEY9hZu0fioYwsqA0IUyH59rjxF17
cbcVEtQ+LC4VWUhUQkGcIIptvmO63qt1RM4xBOWYFh4YNEHB4i7R/zIrviTYqy318DAsn9c3NLmH
xt2uWvlqSaJAdsHYk0/8Cjvp2F4E1lU/b/sGZxS8x8VyziomWshBCOGarUrC1tvTRcyM0gfGKTam
WRkN2cjb2wbraHaAjT3TASlu9vRt7gJiEL2gCh4aYrCa6Kc2B+9Y/6ick8O2T6Nsz2eEWMxyRu0Z
NANF7mJod39usiZZxduimdfH3FQRzElYCK3Rk7WljME/dI3UYyYrFtLSCQzmz6cIhyW3nL/jhjLN
st0y+oH9rM59qIuET4Dek0ojrbLC0qZ6r1yQHOE3TB0LWX/h7j5uEK09Kbq+tNqVP5xYqfjtBGKJ
TEzEChN1BsNfDaoJ6FCrumn8jpu0rDbvXpg55XSS4IW61l9c44EdGe5LPHKIQS4YBLJeLiNBDY0b
p2DMlvQPdsqfW19gZAzyqD9KauJMJYrOKZ/g32HYmZJB2dUwcS7M9Gf2KvVtGM7liatTntxol0cW
7VTcPPkiHXyI0ptJ6N8N2nBZCQZ3KFQ9uXdXaA7wfzv7wxMxku058N5frZXNtUmk7mzD62jKPuYu
iaT7Rcv5Qn5ivXyD0yJ5hs7TnWESgqaYM2DPIk2EJpfzxUHE/7ArNh/hmBEJKTvpEWF0oeO27PAF
rIZvMiQi0Sil4azljpQMRY9vMTxn6NWtWIu9rhSK/zfHzZpneNrMCc+5gj3v0zXUO+DIKr2MysDv
QYPbPO8Ibq32paU5/L8BSXe2jUhl7c0YTKUMztMnkZes+QFI2GPu4dpRFmWYRFVE6YPtjyQ28zrj
noUuQMiVSpFbgBR7tWdlJJ3c3zhh71hPf/a4TSZDkSFDEtl0Lse8LTiwyazgg9Mg8a1vkDo+fjrt
7EPrb3St/w+C9y1ztJ7/S4HusdYQ1/8mlkeAuPSo2ysEUlijEGqLP+yGNGSTPspvJmyRaJyJRgVq
6+gt61EQlNAtXFJGk1ambogVXRsrn1lXzQTevgpyjIu8KoRNsg2D4D1fhU6SYs7n94Ux/CX4Iia8
/L6C+Ytr/4HaqQMwZ/OSPTUV7NeAxNI0zRQPz0o01IBdfc1t0ZfBRB1M5pW6YV/ddqYpfHekUa72
wZP1ibY2Rj+rPh0sWSgdPx3Frvhqz7FOLJ2fwdwWYe27J/tI5g/93qMpCCoaNBPscZCj5d2n2U6B
IzX34qXSHwjet/vXi404CMxq7DSdDy2F7JcdEPsJGB94itcqGNdzC7pJpqerkMlls5JRW5NbzKt6
NRBL/4j0Mcre0l43YUX9eU0r2IrOzbhplQn6nmBT9k7/hUIa+grqmDToJ0KsOCmPO64d1ueAHhxq
quhl8pWCfcM2OvinO4xkb5jnIN0fPRPDYch1a9YxegH3hSLVp7isLWAZpPUsmxVcMNOpYhCcsvaT
XRlwx4PX9XwWoNxZjQMic8StmKOPb4M0j5R3xUrso9gSesCJzEEjVQoPEfANBiVT4OjWFFB9CHJF
x7zQZv3mtYKwllipkqWNPef7+OxrdBRbshJsDaypallODThtxf0+cilcKJ1U/tzBYGaQlE5Xl8zq
JcW3clcEtnriAbbyGx4r826oykwEMHcecVfPj3cXmAUqQRCadghTl8MfzqNW56OXB0Epj1hFoSTa
sLVwjKQ+Xea8uIkpMVfaTkNpsF1m4arB2v6YrK5HZ7wSGmf2+unZ4xtGwj/KbIhpy2kZSiyWWx5Z
sX5v9puoJzgJHOf4QSPyEj36WGbJw7G0jkP/mvBh40yvprd8eXNqdBDxxrwoUiF9so9SmBK2KAxT
CCYZGWC7npBHRjPhAgGvZSRSrAsb6MUES/uW2QhKVCVb3k0sNcqWlggcnNuaEVY+EV702cb5tYSP
Lv8IhpglFTcHu7jP4cqO47cY9rKN7K8nH+CTdECt1CwQlnAXc7ZB9nyRkmrtUr9G47CNNZ6qyCfs
Sbzy6wGHBo7mEgOA2L/pAK1QnQb8sEJW6G9PwhaEpN8CIy75s6jbI6xENv0Lp591P5Hqg/4B2Mcu
r/HeP3tfzNKxf4cauvo6qLEwTUs6XS+VBO57OB1Ji70D0ep6cGuj+1PVD9Reih7ihIn2Ykn+yc11
aZN1v2CxvYaH0M2yDz9RM5K+C4T4ClOwxnQH+DHlEYYx89KJS/KtG7HRUaKk1yckYR0amXV97Yh9
bSB5T5FsVamE0FBTnoI6S/LuGjUKjVteUrHjtiLjL0P+cCN/XSk1I8ISTeLbEQCn5e82o2ANAs4Z
GG62vxdIYfLZPcBbzBRfpNE92/JWnWSiF2kTACDk4JIHrizIBDXD+5w4S3HulQfYz/9xY2MqGgQm
XoqmY21XYuGCrW0GG49/DlTI74Q5G9tM8HzBWroF17MA5Ufu3SwINh+hqQAkGIeaCeoEkIqrI3z1
E0+I3rUtLS7dAu9JZOVeeEkdip99Lxoc2UaoeTzTi9l9ipI7QlpwIKIvhecapqtylK83j5TMvMre
ZNP6b1P09CcxRdgnv209OYDkaZ78pzrC3cnaqwSZ4wW+BnXY7FEEkqnCGoQ9DIWoHy91+j9Yvx/B
RW2SDFUQdb+5Lsh4nhvmuq/GnfcXGtT9s7m1IzWCKuEcun/cdzvCCkJvMffdKK6kznk1b0dweI+b
EIOgMsji9HEYGve20+CThjTy2dRQ2hJIP+y9XynzozNgiB5XoRU3UbHRmvgCMPkPwrc24JtT5LwJ
EXfIadUp90vWt66coDERZ+P4i0MTiMt/Yto9dnM2HV9TkTjVpbPC564oAMo/Tj75y9tHtIY5cqUb
vEsssv+8WPQguvqCImKrCNgs1ktKrbTbq7wJDDfC8lncm6cwHhqAyojZ4qHE95cuU+BTg8FEKLFP
WTbVJexzG+pqHimep+8eIrBbG5acnMOnk5W9coJyvQXmgiknyT9uWX5jBbu0xy78LlMY12NHjoyC
T/iPgzqflckogkB12ADK7rcNjlPtb56LV21gNQ4sgiDIvl3xklyBz7gGpUKVn7pjAnwXQM+Po9DZ
EL5CvzC8Km5zeY6TXcg3+1rTW4zX8qEH5IDAbRDKttw1SUW14w30+sg2D/+iucLb6MLpT+uv37us
SUDjuTJ/C55cYWrA9t5im+7JPBs/plJQUfv/RtKpH8yXixxFEhMWByOgqRYG76B1LxjbfkHyRzNA
GgZ3LZUYRRSTNUXcmgxsR4MYfBdn/FXm+jlr0xgknYH8JcPWx+BX1nsbhVoB5V+IhuRpg9dLHQvF
AEH3i83BCnKKd7JhDTFpyyBlMsC6Jj8ZFoMubJKmibby7ZNivQzLYHTUglz3z+i9ni0MMPDDUt1E
8tKfMP4mzT5tNwWwG9R0VffQcZhslK/bQPOv6k+SWZ1nIo11LLLMDG5xuQW1M3zt15zpwGv00n+T
JrDWc4O4b3kkaM0X4dC5UHPq+SRALYjoz22s/oKGc3TlMMxIzxeyzYxzVtcaqLB/VNMuhVDbe3ot
3TpthAxuXoF2mYV0hDp0/+xAaIk4QjIlqC052Noc2Fy10SR+LGDovrq17xXY1NWddLuUbxC+UFMX
RsLybK9ix2h1a7er21q71dehw8TsbVJkxlwVPuxGWLQ94tuqrX5vDHpNOBFdCNgEKmZK5Ut8kq6+
iDVoY3kx8YBV8tiUqLBvRe3pmDnN1MHUzDGzk7rB5+z3APxuNnFYf7ooeFBKbMvFp3lXGFPwp+Ak
4Vn5mK/wFQwOrXY2Rv3lXTwaQ+S4akArgy5jYOL6FKLqMT5i4O+VSWnPMVGhIuIKIlBCimqKRsMb
R84cxKGsBSHxzq9Xe5j51GIYObiLYlfSVcL0rmOxUbj9B1fznoY+vSITOmJLiNMcLT4DwcpdKNRm
7rzZca/PD5eJwgD/CUiBKHBnRE9dKvh68Br3NRirU+EfOXMBLyjTSdysEjjE5nINMGCluQtnKZRk
mT7RJadEvjLYwKNr6BWoHH7B5RIxpYls7Uy6pqVNotSNewOtNQhjA7MUK83yS3ES/vZcuhXyFpS9
uCknLuef/+y0YjHM/LHJ0+XCv7niPYxDIvbKRZ9flDVOMrM8bABUfpFuY43XVaE105t0A4s0bDEN
Dt5qe8uhqocGSjKn2fktPEsyimzPDIHjXerKWmE7Lsed6HXvRwsrEgQINnu+Y9ce3xhsourPMj3Q
ZlPQ9tiYCVVhmt53Fve1+BAOxd4fAWjI82U+jzB0PSVIMLw0Z9I0vpD+GiKzrnZ3BbFE5NOH+iy1
xmNJSLXb0s0f9IeOf+qUe1CZIPW725ukGW3Rhcgrg7pPImOUlW/g0jS1nVhd8nE3jt6Mtz2pga8L
clcY4S6numZVmlGNkegoDC23S/S0CAH9j16l9mlLIiw0yCkitOUsuj0hr/36nQUGao/6mmZ+S4Ko
1MlwcIti7NQ+ziG2kEPp8EIoyie4Sb/9+J1lYgKR+p5Stv+fo2ASiBDBtooAu2sXVDRvZtShz5pR
GJEVwHxXWCst4Ox5JLTFvZK/6abB9NRoUqGpuxVblEIiklxZN27cBOhJlVfkd855YM1k//rFK7Iu
KoliJ5G7nWFOXGynMIVOJA3aPeZNW2Y7tmzIVK8fAav+1mmVAjTxCash6oSqVHlKL73msGdOuJWM
2mYd0kJtr2vqBJwhWkAe4lKIJeRRwN4DvJHkHzpUbmz7CAodECC/ld4J7+zSg0AF/rQCGDFl/of4
ITRcBFd7uw0ylhfGoP28LhVGfgQQAkTTG31aTtoiZpftKGjjT9m+Hd+ypRvoxj0y1UJtOCHGkK96
nbvzL8nk3BwZuNz5e54fM42YmJZb8R3A4iIkJ2bQf4hpVUPK8AFvjCMygABv2O/kMs2oQ/OetmMM
g61vLO0r+Yl3VOBFVd6Txe9xk8wRmdj3Iha2HfoNC1ctHzGMVqWSJP6Fz9L+1vO3eThHA+BbdMJ5
u/TtKyceAkYPDgh7gAphahYCjtHo/9n/WCRdGl7Cyikq9kE0OWEt9U7oDtsz7dwty/JA2STB9dIj
blPSgWTUuaQ+38aVuyj3mGOzprJbfFQljKHtKbKeq/08+FKkdb8DbhxaKB3lvNy5zZSjqteoJfdO
lPR33s552so4S+c6gK+Xn755dow78zzKmuTrAU7YdK9CUudVlHM0PABZPaCf5DNSk/03+WKNQ56L
QXl/LTqZ600lum3TPuz+SPFg7vCUa46z94ugqVg0cEg/AWuQ3Jkf0AW5BzokkSFV173Vt/kq5Sq1
Hc1XTkiPMBCFQ2tGiTjmnSBcGJO/iuFUIic0/bx/b1A0IwWiam5TmufmxTzjg/4tNZYDoRjUgcBy
57NFEMmUdkcigKuvIT4/w1H3I9EaaoL4zSDLjW5vmFUhZVhdg97xHt8IpOZ+KhNTPEfmgNM0IIc9
d+Y3fHLp+7Z2bg8VC2KaFgxFU4rJuf3zi53L62jG/BYZQPcMWnW5lbsPnP/9E9xp6h3y01gfDCxs
fg8nYepjFcGUCU1waEhaVFe8FI9wBXlysc4MMhRzciDchj9aq4Mio0KsUIIgpYM2q05ZN3e8EiJ5
K27MU81gvAIGQWjt7uzIfz1JtqR0oYlMceK0lV+jTBd6SjhBZy1KCKO4tiFXjJod+SZuqjTDagKn
RNpNL16bFYYWZaOzM0z5xVCFLC5b7hjXIp7jZu1GV0sksCl0gJZSk7lJ+kPUIUuhevK3EVjpj1U6
Bt9Ad1JizBrB3eER7u2HeECVqNV5iqPREVmPmIt1fnJW56tioXcXUHwfZJT1El4mzJrtOtG0qWvF
lIPcvpBCJuwzYSmIxmyXRj6jceoxNlosiYWB3SFeWPwMnAi70LOnhrYqVNvTLbgfWtLBY66XIHBl
O4vhlhAPEgeItHEpedrYaOWr7CScUCcdlnsPdLHt9UA10WE9u5MOd2U6D0rq8bdtjLgSeb4JNn7/
NyugKo8INIxQ75QuzA2lNU53q8Bf3gFjf3gW9pX0BIUsBK7DaCDvCxPbdq0vc1MQf5HF1v6Db461
sGEIoeO2B5Voe1/fIHEh+u2IsXCwO0sOncYeMnooTaXws3uJhz5gHZOB1mbewvwOMa8ttkWNqCNU
wRIvICav8r0fWg/KybFFwqp+vBlKT4c+Q0amwuGu3nSuxbEWL175Wleo3msvr0TTrSkCowfSq5G6
mdZ7VElj1n3t0Wj/OUxLPzgXI8GD1xQZ4jLbJS7vt4b1hIDYd/BE8FxJNR9RaxxTgmEsZp5B4FeM
eL81SikOsK222gy1umraMYvuOEIfIgH0Yo6mXwhl1Zj5iP4Uxm9RM9KPjE5xuyHhA0bTN4K/Znfh
0aCDrK2OBr36huRvgVg8JumT93HDscKVyZq21yu76nrVEpQm4iNlgBHmklY9ETURnM7YcGkjk4ae
8gAHVjuSwsVwN3RGeGSq44o012y1lJqnumNjxm3cIHEHZgbDdVRva1yUAd6j54jxx4sRWXuaUGJs
FhuJczF4vbpgJxsQRo48UV7gBuExvanamOP34CSMXaFjQwI39CHX8obLCH77qUQNj7BuAxArHya3
2vGZEteSuHeCz7GCslTEbQ4CX6BZHCBqQhcbkbfPmLti94wUEREVoI98BjVnrAa2nRifMMahNSAW
TMzUfRUZNFs0IiHHefh/IG/WtoHJLgocZAqkU+sY2Hl/RjXHDy/trXtNeWsAeGV8l8ma6KQFrj8A
K38GKOKhjMLb2KsEfumyiK5KD2qUUrVN9d86i4p+xJQ+evxH0P0CEVIehwbJWVT2MHNhmU2fCGh1
+EZhC2W1XGjSNK0MNPxjl+0U79wc/hkXcPyFS75conL1EA1dFrH2SaqVaVhVBS6Vnk/IX4EPT6uE
pmpXo0jOD8K0XjFYaN2apG+gCROm7WlXP2vHj7JsLaiA+vofRrP70AXkjYoNbIuOjWvIA+seFE3y
YlINaYpJc8a/ykT+YvW+XUhbGjpaphN0VlQmVGoPgQbXSqYeS+ucLEIeM0lqy+hVSqC2aHYglyDY
48oeJCVYZHLUBEtZoqjH3fExj3lYQnlvgk2CynuSLWX85bxeLjDYyB15JVk7YNq9Y6UDBCN4RxMj
/XD1JnslfQhVYrVIpHim2p44vK2IDNSHXXeyHo81Rce905SM4vlCnagjXZBaLOMfJ54tcX2qVUDj
IVF/6k8WII0LHYLQP+apSZEx+qy/5KDd6+q6ETyNosmW4bXSRNYDE6iNOeTpd4Vg+GV6BOTGHys5
R5ELlgTpvi0E8h3XZ/dwYLlgq9+BNwVbJD6s47/RhwZvIf0Y6wX0VpYd23UlKUNq1/yCE83E5TlW
PE+ZsbOJp0Rp7nSGwyRThqjOLQNZ/3G9JSe0sIBObRUQgEqO+GfnYV/Ue9tdV39bepNVDnJEb1k+
b7622db/Rk0SYY1XImEf7iC5K6vgh75lFz4AROsNV83FBCEVjMt2SPYrvKK4GqXL7q2JNDzIpZdQ
jxEMt/u0QbmBMeHqvH3ECZ/sLliF5TiPXPXffXG1L4pgZSedy4IX+6+TZU+1y7m1UdwKQelllh1u
S/5duZJV1Cpg7FRCNwzakek5tK1M+cMDOo2SiKlPYq7ebOGZf3iLF9smdOQiWS8Qwrb2lIVabFJY
t66FmQDsNBaTsb3POgjiCOrPRXZqr3/dr95vRYS0pgTq5dj9cXmtPiLI+GTgZhswmp+7qaO9ksd1
oTWrRt88Pr7dIj7qm/pqdLS6OWf+r7M67pbIaTkOsPj38CKQA1/vl3PN2AZ4dblG90zVB3v0QpkE
W6QDwR7Q7u6a/f+qQ4VW9mZumFNksdsZ3z+C/ezH8SWI2ZewjqAhMNIJ9zS1DIl3HU6wvFDFYQaQ
PVC6BEZ7HntDvYzvLavt2KOMKFtDSL588CnMQVFTJQFtbJ7FLAXJ3YGL+wR4FxRBFk0EJKN2n6IW
fUDABbycUNvBjA25FIqqDl6tuVRVDDMZ6B98L/491lS3XeqXj7NoERlGBV9tu9QgXKtx5b2Tasrv
yW9qUI1JeSTqvswnqExrl7I0fudYreTh9SeMwH8S6+e09r8Y17TgwUBqnejEndGARogswUVIIOiz
2NwjOwkFKB2PR4VA1xQYBIEONalAvntZvQH71G5NYiseG+ySjIbQEYbp0ZprPGdDUGK19ECvmFgc
BqH5U960nf1hAti2lwcgycuqc77F4uwYOOzyM3M21aPdQ/PvhDLRm6Tysmtvl83Lm1ACRPjF0H/Z
YRi3VPH+1CMT199uQP0imk9DwOCf1gNFss5COLpNY35Lkmmc4VPzy4Oa2u7OFNQsxTe5110p8LrG
YHkfmh8ogzhKfSJKbonWZAspGDtbi79cFlWAFNldz4D08CdPsgj3rEi4r64rkrZDz5hLx539Lbgy
yEhXSUszIRCzT0LN3slm2/ZB2cUSMXqSkJme7zahDL3qGV9YtESfpU5+pPRcEbUeGmGeKHazWrm6
cxitqy3P4GvOG/h14RJtnt1T1HUCVglI6VBhQhFVRCVEUg4nUP3lK6Xa+iFQVRrydeZfx7QrfN40
YT9mhcOScyqfmT4kHmgWKVuIj27TRwCw2owGLWB3glWcLBdAMof/NnX5OchlOWtva25N8gCqPG4Y
0QnkyzeYr4pR2FNr7tvbHKE6vmJPwvmNk1NcVg7cFlgAzkJKAla0XkdrNsc43D7uRbYdqJ/CRenc
RpbhfC4IF8wYNCLDiBGgQvdA6agqdQRk8syBZQMGuMk9oSbB4mIxnARmhfY9qcN28Xf29yJ96ha+
orxQfc6OooUBmTkNtJXAdL2zR97B9qVAgmg5Suqpd2pJZgAYcqo09rQMT/fkdctlejR6yw1irn07
XsyNYTo7iNL+dO3UX+Qes3Ef/QaWxC8MTX2n6j0WMva09soiEMrMlUDRssYLFb9m+94uh/ps8aS8
tmszAEXZz6mZBopkWTRuxEU7E7NLen8AxgQcRYdGwUmALTlkVkw7hIbnLy2QjKiHzyLXNI9CzKhM
l6Ldd6rvKjtOyJSWN29SM/ThxaBh56vAjbRopdF61luZduDz50wC+5m8aBdUalP54ZMy9BWY8U22
bkpEuDxJEdKSbABfHusMheS1ikstVgmxWwYbbey7nLe//EEGK5OxJraMYFkehn3a2cFVko5v/hsm
hSyXBLhOXfOcgGIqMOS0r3Qrc1cL1rmFwdjahtRyrWR/YiQ+HVkLUJJauOC7KWrHo5ak8yhLguBb
uAuuxn9IFSVu1CUmkTcp/aIWSuXcm6++X3JYaSid7QuEDfByflqR6+Z2p+739SRdXEZmxqaLfFrT
J4fXi2wwNTWj7um6/JkvaZP47zf+cQ7KMWugvTch1j4Hk/OAp8CYApj/qm35oxudTiulRkqOC888
6RfUzAucEcbL3LQz8S1HMZ2FNbHfW1QWGzo2ElQ0MwRKceprVi0InxVVy4XmoPfQjW5Tap2NH5Vn
m7tECagJ8FmjPh50w4pxdyQR9UPov69KZbshwodMLd/cczOzYpxxSwQqZcH17MLOYxTFlPxOlP3t
LawgjA2NsK/56KdBXUNlL0xyCsqOYrJ1KSxKgpfKL/+ZELq1OiU30pzYZkGVmKAAwwZ3Y2DnFHvl
bKZe8shQQJUEPviy8iqZJZLNflyDPSF09g+lKx4oXxMnJUkXiMLMhSS7nMNL47udxebZblycSyg3
FIx2LP/rHBo34v4aFypSzirYZ+Z9XIkSosyEgmVtk+K/5WX/ivMDJmeXPnllXs/HYI7JzBc4qRXB
16tAPC0DpOXTtX/F4/xSN1dhBcKQ7N1/7Euo8uZTymqghkFygYKI7BYsiW3vz2T75PjV3uNLV0ix
7SU250TVVxNm9Ea+txUgGuTp1GbzBxRkzah1cjEqR7ln/XVfQlEbJKkka32mVfeA/UukFMNCytQT
GS6qH1liHFbI4UdXUn6+NZ6t02YykYOFuYbx1Uc0znMAdF5cHXPoagwzonHvnT6Ega+KSVMZHCTa
DM5tfHkivqvU+jEmeszaSs9rWu1lacwYn9xrLdVuR7QE20DmsvuV0plSqXSfR3fGIeEhmkPsNQlQ
4c/UMNqB6KBWTfYzTraciRTxzhfVgSGyTHSozIfOAHdFQcD8f2ubRus591uswl0BIM5WG54tziEr
Eu9cnSBbT0m06vYhsN6e8QczmKgHDolFYSqjDSh+VECJgkLpZjxolFoSVejhZY7GemWTvkbgE9Jf
i6y9sYGAOTo1C8Q3igkTzyA+mx+lAyYqMKaz+DNMg3hwEPXMtoZlFBXwjNxviFYLY3JkhrdYC9Tl
G7sYh1gjXHr6SVk7UDUUWCMtLF0YATJS7MwqVdx0JalLnPAv9H9Lbt071M+4wEh1vtD7xOSn3i8o
e36n60sJ8ilv31B00CWuTAhauMTKFdfPlKRP3ud78pqt04SpwKFqdLkBohK/WXytmavS4/eQyWhm
pFMvi+5OtyOYPqYBwTcUcZwFfTmO5FUlbdwnSiD4BAlXi71VEdZwUTEdCWEXriT8A9xzhun3Seld
PFhIY87z6wu6XHuZ6J+EGsm/qV9HmANmxEeBFnezPoETaPVOpgAXIWpVwaHjTvGEARu1BD6sKedK
6O1BX1xpHkcMNKlrpgssnsBH/qHjHN2yTprztikmx0yozdI0vxwDXb/Y69Uica4+qBFVKwuNxCJJ
HOYf1ZgWWRJTU0jl46MJ5vNj2h2E2tw8htAPoUMXaaST37vjqiPxU6tWuQ9RBb4JmdezeqEzShqR
Frrz5J4sMWAXsyTD3+o5BN7J9Lw9RPdpHPnBkzCK91i/uchT1yRMCor0I+RsdMw4OK7GcSDMEOM8
Pa7P/87fWZE3AW/UYwvnLNJT+4ikm/XLQteUz6QPQhA/ZvlOfV7I1Ygw+tlXI1AvZYxb1t/5ou/H
mlnqRVhHw808MbNCSnNm7b4piqyelx6vEHyN75BICjm2N7M9o3ERXU6cMmUUcQ+5aTR9Wd9lJ0Vd
o6FY3BstUwjK5nYCFVwrc6Ispk5dDNbwoGiJECLZ2HsTWMoE50Kso0Y6Q6ZNn7gpehmXzP8y6vrF
vcU6Cjk6OwxgR8ZB5iLMYMrp6Cs7hKYFOjWKDeP5vYGOplFIMl/fIkQ8ZUtRvV4UDt6xOUEK8nwt
2VMTTmB/wJ+U8iqQFRDFbf0pgtHKZFp/8cbYVZAWh7I/53U0ehTVUhNHmwV5NRgMnAPWTJHqK4LN
zfgZC3HrkxcJorDMtsdAcuEN9YsT8diqmgmfjldGyi3RCJ4JusiBc+aPui3Ekrb42cS5DDD8RrRY
faJmPqiP+Ecipfk75FLlbPonwaiOfyiP/76CewalLnZCZgrZCjAWN8BVj6PFzEEqZp/ssFDmC/mS
c+yX/Yuck17hYhisKI2hhTAbEAJh7ryIb9RPT5imUIbnraYgBe9rSzkRAPuZZlxLWZQX79lnr6TO
XzrFbfrzNccCzSAv55dMhwPNsFIql4RIbIlk6dM6dql9tSFq8Y2m03RztlZrQdKFwd5RYugWkrlr
b53c3CdV5EvnewsVRjnWhkCr/AkLcVYKqqpXCrmh9cApevdVNYB1W03PkZLFkITq7HlIJ8YyAusx
jMuB6OrjsIORQiOWc6nl3YmjH5/9U2ZvabtG8E+aLqgpvCnFiIgCfJ7fQSJp6qeUleOOqGisE0YI
fWDbzNxxMx3PrZ2PJ+lJ68SrdX9sM6OUU4uXqqgpNafoPnIK9nPiXNfhfaAZ2w8opeMQLZvkbzOs
9hPXFeWHAqTi6NnZXWFYDTdT2KaYI40ARrJEdIQH5DDSXreT9+Qm/EclKyPmIwKkdNc7MXw+MdOk
9qTiR+dYBDtmmO+JdOHXeJ94a+siJgBfWYI+DO/mofl3seekV3J5+HBe0jbogBx6gn94gsbfBliU
TYwrkMqZZ9xq1HD374e//qJrBYoQ6gnCJ/PAFdnuyHuEispDOpE38hOKAFLiF5J9A0jcR12zEubN
xOwy9vnGPAzUtj7KjS0FcyCu4um66w1JOFzC5aJCSNk3IIb+rc9im2Fkxq/bSdK+1flQIQNmSeV4
y8N/Vz71OD4xdD3ji6COcTIGsymA8YPHBM4c8yopkAYTCgOZB7+5vNyPEMmIGpb2JF34pbBdjZYH
1n4bDy0QaPtIT0SW3scoOHQdlMloqOjJe1jQ5BSvr4ZUXXv5kQRaK08awaNO/0qVoKKpwXXqU60J
zC8fcG6cWgtXgel+t6xbHOjRHH7tMdUOgm//O4hMebVpakHHcff1YVikF+fN/qLZX/Rxpu7PBBwj
ti3rXOqujT0WVCqHnM9eeK4n3qjIInsDGNnr6JLlWyOcZxTrKRjOr6cSy9zT3u+d/+jiRtUvbRgf
x51YbMoRFAFXJ3Oh6sQgf+bomUj424IINpwxXk97xameky6wnJ8fPtdojidoA9FozPR8AZHWBIzl
3dUH+OL6EbOjw50Vux0SWEg4jYHj9HaBFPhsO5BbPcw6vmKuzOHBUv9Lff85xpvW/SOJX2xFkiR5
H5kumfZPXxRof3FlnoPNXlJql8YgEUga06K2pV9RVRogCMD+b+wXQSRVZLOD+myZKI0M/hQXeeHu
vU+6QxLGhGabG4OHIDtbfJk/UbGBwAt7+ebEpA4QU/oS6H0Dk3gJYsKD/hNw6ez53J6161N0yJt+
U19nba/Vi6HJ97/z9OeuBnjXgTtybAaotiHWqlJrp32LJNs5y7s0RJIEW30yIQ8bYWAb30c6YKPZ
de18HDJiWSw65dt4fKv5+w60CCSQ+99+AKTkNb/AR0AkFxFlFoEBi0eLRO+6YAgHMdUFt08sZz2D
88WzxtLlE8231lzpakJuGdOZ84EvzNMLF3xADoTEZH1hBU/SYEoJvp6Hc0vihp/00xWLHZZmlXFc
JkYDcwB/j/FEl3+O5rlV6CzlqdB7HkaRxlTyR8/uAnIH6Oq8BckWh6jfJyP4pxvHybO2O0LgY5oE
0hms1tiLwp+URr6jD01HOlKJuY/nMUctvmT9p30IQlL12mJen+LGSvNPOml0Poipl7eVeBhDw8WC
uXpnFrfyXLcf4ZPbPxtAbdhjCl989dN0uy11makYwLkBYCDMm46kDvKnlNLb2HPT87gx9qU6nF/I
WP5/5DWo5vmnEeCjkHRXO9qF9jnBRnTXGpvcv2viaPGRaGtawEBvpuTHOd7MFV8sdogxWrYtr18G
t9x9uRZcKXmbKiaTvv6hRLu1b3JTklafzijDmFA0MGyvLkltaqeNUIZayDQZXBLfZnJ+Et6P/iPQ
NF5LKkyhg27AYqnnE8bjNdNQ+6JvzUyIOQH0G2iJy96NhfwMvxN4vwoQiUebTplFUc1tQ0joCM4U
AkBYsxlivHhI5DM9S3AV8J5G0f2LMsh67hbUT/IHpyAHVkngQQMIFqzVEYk1BLl7CuDu91Rk+jCU
iC1mjW7++mAWCnLSWDBM0RqcnfGmRMTv7x+B5hxf73HLg49HT9SVBVW1qq6fO4BtgEtcrLsW3PLp
1GOwWagafUKB5BZS/aQkPYcR33bcm4VY4dIIGSa24pOTBwwEeXba6FaLUqTVwZMOQxm2/+DtuuVd
TGWiIPA5k7YqPhKxf4+Acb3TthmuoH6RQcPz8gWJZ7vlt1lLzxWQW9u+BYGBFvAYMSVNJYCCxG/j
63FAZKdNFGrDUQCEATjwJO+xfvvxUq7GVvBbLx/3hvK94PJxZruclqrq4UI0JbuSlo/IAI2aZjG1
DId3c/NjIDM+WyjgVAQ2cw88sUK+prYiuoJ+Gsly2JXX2HQQOluyf9DnKitFbMLUAYhRbqUzQYyL
meXhtzaId+QuJ4VsHlIvDQXXjYsUGaYxAzcPMnynbZP1HlBa2fSSagjdX5UIE46lA0aHVCBEwf11
1lFaCUOtu6l/9nJVg4qYyOAs1VcYpf7JGu4EqW4+rS1pJxq2qDUEO6pLcPK+sfAPppe9GmPUPjny
vsjpdVU8V9KmxB9kUd3UR5/lhyokNStAIH1pIMAX1cDdiuUQxLOhvAnsAlqVt36n7p+9rd2qMYSE
QTvVL7ybkZ0o0ISKlim7s7gyRBoS/3LwwZWM/HfqPPE0g9K/0n22ky/cxaN2Jf8Xp0p05En1+kSD
nC4NZ6E+x0UVNryG5boTnGkh78HQ0f1RTczXmwPCYWaaKiKVTJfUblBRtA0nfgL09xUJIDrwuA3i
Uf8Y/E6kSZ9mk6q3fy2LilqdeiDg7AlO2k2fDOCGfUJBoRHbtoSzUiMdELbUCWVcCXp8ATfwMDlQ
VYUaJZWkEk171C35cDX+oLFQFRRjn6Yrt5hYUrmUMc9gi6N5f+HFJ24jtT2KvM5QTPaXo2fIuRmG
pJTydWiPrtiM12bAuTujcvyQsQ8yPp1sX24QLzP8R5Y/l+7H8nbDemhEsMHIlrxlAhxoeekvHluW
8Yh/bnP4yHUJTHS0Vlo6S4XCPJ0gz4zEyp7LY6xudcIEmDA353mmjLgTkhojXPgEScjQTZhHHBYQ
N7hFPMXvgvTUnSNXIIJXkZ495GAhRaw/CCt5AcSjKdtVVsCh3U1k+oeXuO8W2JfO674OLRn9KjlF
x3UGoNMCdXpMrGBQ5kMhEiBxUCBUb24b4Sid9z0DtgAZt9c2iRY/JLBeL6Pkr3bg67q8xjjlpcqG
FkZV/LjtsXU9jttODj0OU/0gRV6GbGc76TkaN+1FEDstKdpil2USTkC5To6OO6uXS7ASwR0v6PTH
rcgA62NWL6i/Jc2o77z6K+OtIQlnFD4G/pWxKAOgWbO0wmlqbWcM4rMMJqDt0jlnEX4UKmmhu3LR
N5VoWegoQOdflGfFFCMqp4/6AlSRl/KwQt3J/FDZhU8KaG/1POVp+6+XAKRCXSr1sUEYnxzIIlf4
gDb75e+Ynv0Brkf/WTi71t4QvX3mJwzt7Mg+X30afEZJdA6PRK1pn5/rREVT8NEXFaEGit5MXZUu
RNXs0YKcjseLkUzAAkHgbbC6CVNi78n2zz3vo7TmwNrhdcLvAVE2VyuzKZivFIxEgpTBwqcWA5kK
Oz/qUKThg4WIac++rHyRPrVHHJ891JTKmKQO9G7MUTQCXZI3wPZGxDOjYlr+rqX6gjH1uYcw3aFG
DIlS8QHX7k99amfKA7AmQA41T4JbSDV0dXVO2xcnoaddFLQCE5nI1KLFigv+Lhhh17yz2GxhBR5C
MILyihc+6KS3H62bSyoVA8fJqLSSkkrwNqgbGpKGIlLQdyegLteZj7F7s2DZvhWKyNzecqjxFRGR
dgpIDGXLGkOtQcgf9PrnAwvtX8m0/ASlJpBbT+oqSpgAz7n5OWhGZG2geKhiaY2j1rCfV9Szubcx
Z7WjNm0UbrE32EJBJHP1F9815fT7kblU2pK5zf6y+z3hQ7i3CK2ffJRYFy7NTiz1IIjaaDMTBqC5
yxUgb5AbHa9d1nva1ox00Km8I9Ey1fONfkOX14o5IUeuoxrXJtViLKu3y/cbFHPSSAt09lsj27iI
nCn27rKKbMtSZqiDeoym4GQYLNpBWR3pNB6V8bqIqt8VOY7dhWdOAU+gxSH0oAORpexJWvBqFIK9
ZjxVExyoMJKDc4CQouJD30eY0IZn0a9u0BbyJlbPnnXwTwNwSV1c1Cvts5R5OMNZCtZzrjFShLI5
wjqelPWMNvjlS7c+g9NI+VbFJfLv8SFFJwROv8qSngygGXmY4u9i5rS4QcnbyONgB2jYtLizroM2
g/D4t+FHMBWMyMyEWY+9EyFweIM0bjTeOb4mXjnQ9XBnCErpvoraZrpzih3nlKqNClA6jSRnLA4V
2xsYCPwLMfKP3+V+cj9OyJaWPByrJ0Mg2knpIzWOAtH7NmGF4HAQe+tBqgUdtZNF64rkFd9oeXwZ
45wwHl3L5uVo6M8pD4tsExcV9YJgcfQuD8RGNhtSc/zmWn44xfLQw1a3vHnorubTeISHieivAAXm
bIvlSTXog5wI5TAE0dfJgsqIzWt5Sr6QDHb0v7Zyc3qR3vwx69unBAzWDGnvLx9dvgpea3KbaYT5
fm3SnJYDqOixK5yC21E5T77izy3W7jSfiOjVa23tRKTW+vTV0VJQrjod6mnXhU4xOojXoqc5/jSJ
pdg1FNbx09T/6qmOmYABEPNZcYCn4ntox0kwPFUC2DoCs1uIOLI91zcZem3YlXXICS2nQ25ohgtk
bBNVmn0wMiDgKhRcNhEH/zNcsME40WG21m9DfFt79zbDs+90HH5mJHb2Nx1kYJCu5r5+Pg0szEIL
ncx/R+v4WhL0jI6JFVgChb9N7F9EZU3+C6XJ4cS02DebfBVvAuogMtC3MzJ3JYjhJAqomS15b8q8
6nWFlPIXDYzFc1q66T2tl61ZsPMtJ4MLhwpMYK/mz5d5ahVQzlM7c8HdUgpSd0F7GeLQdAohxH4B
RzGSysW3YJ05BeQUTpgO5yhF22mKPfNtHVFP+x2jgIk+2lpIGMnGMHCU2pFBbtQdBFvK/tuuMGjb
tlf3xmGa/TJYXlFh9rmNkepfvUypR/6x+a47OM2KAjWQau7ZuTvfoQV/TFjTviLyb6hn6iQal3Jl
o36gJbi56s8iB7G/ap0qrtTRMIuuTR8P/BMh7wfAPBI9wnGZve3axJ6dBi6wEN+pUObWmsQ23Ihq
ikTOeKvO1QRPmDhRYsr6CNb/lbUL4TGOX/Mlk6xnkXMu962JAtAgBc4sB88aEFZ+PFF3G6F6dnaY
NM8S0CAED67ki0hyfHAthycokvNjafeLiEeA9sHjGw3Uj1+v+CS/EZ8Xr4SIepQbuSFQ3cYWblmH
VS9orbyvC9eiWmV3WbGJ7dqU5RJVISIBTph9jNw9D8MKHUVVlXBGMqJayc8VTX+UYy5DXZJTSdmM
MRVhNUebpb5ffgol5QlTTQ2NtXedSWY4USVszt/EdETb5YNdagQwtKan23SIuJ90+MmxT0XRt3Yi
AG7GwhGchH260MSW4YjYKVT/WuMXFF/7UNG3vO2bWa4BZlYp+mHrm6HhSpMENOP+IErCvtwsWKFB
rdnWuS4ukd2SFKz3n/JFVn2wzxtp9ow1izWCmacDE+5DmNN7P5vOulE/h+PtQM4Wa5h7CYVewUoe
HsQF/qthfjtZSngGBFLL8p/IWJ9DmckXLDDuoiIyhm4FlOaXSFHnavDohTaTdsdrC3oPuB1LgXqB
MWXbISXBMIk867X9CTDTh5ylUiAfnSE6ZAelfAfDu/6H6GQPYRUAEzmedC6OwqXvHSAxrTiDkd+v
i2VfElDYrKYb3rPOZZ1AD/YvkYnmnK1mYfxreCBfQkHiIztJvS8xR1qWwb3wmJkqfAOU15fQ/M64
/bkDCdYfkr5t9xvZkNNTVCKW/EU+RwsA9jpO9TmjFxhbnPjHv7lm+bZHXjNR1jQ5qVhbnLgIS/8g
E3kc1HsgAvREyPd/QCImb78Egnyi76crMP/wuCS5+/5DwPUHEzUcJuDkYJNAWwXBcSRn3ubH9jmr
5lNxZusm7c7zl2U4InOD62aMDltRoEeTUbDaZEyac2y/hXcd30s55cKB8TBGhxNcqUHxJhs/OaV0
Um4pQiX7E4sdKUonacUYDCJUzh7yPQXr8IFH6ZaXlFbdM1HLGbZxeIac3jGu2eKG1E9yM3AD0hJF
cmIuZGuCmhTV1m5e5cAy+YRdh0mzUnBzXfzbmAEraVrXtObXfXGEaYLIRYY1QVxuIJ+KtkCXa+n1
vsy91NoojzZSoAl8yYzRnUfv7+aIiPXU1SLiWionjBtwA0xa1j14TLLkwAuUAKiSD0pgjRGf2R64
ne6UKuAZrhhW5uTMjxudbqhOYBQP5rboD3imgL3K5yqj3hUe7S7r6JQxYqCX0+JPh9VDuA8HiT/L
Z0pt5WoznufKeGxTZ21dvPj4aXUtKArv6R7HMG+ghEC0YZFT/gkqOcqclkKq7h9kq2YDOah1TBw3
N7lBU4VC5IM2Of3hE/3zuMl8ehaoZnKNicEaSuqBeuwwS+2FD+dyLZ5eO4nJyUtngJSnYWbQXCln
Kt8sB9pmYG5R+/j0Ei8jDtbEB7wYM6jIb/2szC3A8LnzrRU6/oxVYmqNXutN526d5rMAWEme0TV+
KsZzwvzXV0XNw1ZzB92DTBn/5i9cVbiO/bcATrWnBDoGmPt5xnzkNeMtZpv0xsfoZCUw1KBhYDbJ
+7PlifxDK+vDb0tH7QPSC7zb1pzcFrb3zT4Rs7OqZCuVRUVFDYHiXuwZhdsixLTV2tzWIjY7EXsb
j4irRdQi1UQMiXgGmPlLhu3h6i86eoxY2BbasMJGnqTgXVs6ptCdisdjH05T1N8/8SO9BQ1n1YBW
OYsbSi9FhVy4HuR9xnregEOV6q5Jp4w3o3QIW8SPyAMvx0LKzSk2Ym4x8lotLgZEaUeBfbfsBFSP
4wPhg3XqpRaJ9xRPP7Qgt6Ihp4xLKXQx3XW37IHkfyIKf3T0gkTUPeNujnXPLv+2yX9QoGFZ7aMo
NwVbbq0W3N7xMeMIuQ2ocEr7cH2SNEuayOeiObz/Oon3QWX3BjhYnpWx+DtzWzj3wgrnoDe6Inqq
aMrc1hXYaVFNu5jg4K5f+74s6aQKqJZok6kA3NLI5hS/bwjelfJTt4R63Ul7zm2HI4ZZ6NGIdstM
/uKG7VMIBgf5L4rjsp4yRYml5zO/JF7Klf0FRJq/OLnDhTrJMCutj/VyJ0BDHEgUPU3iGfvK7pIc
3Nbh4TXCrNH7QIlSqy/3quzI+1kZhxYBF5dBZ8pQhfL/1RE6q/ylXYN1OItX5oevf9ocMJvHmDsQ
D6FiMzoyZ2fm9WPYZsT2FGx9MPS/GTm3ELOFijAVk3QKtz3wlEqX28DvphNv9L12cKXvdrh0UJtE
y0b/ttErsGYJeYw7GlOIBuFeNhKziGBHwAjKvRFlLaPj2UjLOgLpzMj5oYbCWfIE0J76UrjgXbcb
o6eYGiG7t5ccocruGvsDArGkbscBKusjJuDz+NESEg+ufUsQ04rbw/pMwONbKkMl8KJHnIfl1t7Y
HMVm+Ta9NFC1/eBJfVrfL6O66DRNlCjM+bmfkEkhFp8OR1sj/FuXJmsKThZvgx4J4psba2CXep/4
v2G53akq+Lqh2evYnuJw3gctgn84S0V3KYCHJtKjslauyhI5nmJkh+iR3NHnwrCsLp+mzcVe2+cH
v9OrsnYoluqyxrkoJWNouuOENdqTLdp1X577VjyAge8/tuPkc4gcmWqKuB5Z+T1Kk1J9DJ+WCSuX
x7MfwrlDuE18ZQWDq5QRZ09URkSTExXCTHrS1s94zIXUjQoTQ1nP6Ev+wr1Iy9FWVxgurSeITwfj
gc734EQYlbHs0pcdNGhfWEH6HQacm/7OZ0gH/TC7YEEu1rTUnpsEd7/vtRj8iIU+6NN1LJegZHnr
O8hpyio8nObRSrJ7Nm2ZyFDRowe5pRM08fHqsVCrfew+tJdufMOcK9hdZZbEB2O9ZihmmNHMhpeQ
IXZfN0zGyeY4pt0Gzbq4SQckWZrL2sSKd2xAWMoVRy5J8xDkEPQJE86D/fLjg8O2lMCfY/c0X9gA
Ky8K8sqJ33JVMd+e2Kwko8eJf65Zpl6hsyR0XrBktV8Qf9ErmXXEfy49sAoU4d7bNG7lKq7x5wvv
IRoJ2PAHk22dj3vSWGxwrmocTyXYKCTaLHbw0vY4E0bRTqyEyeODK936KPIe1jRmdOy9fBBa2bd1
odaweRlUZ7uGUx3t+cHLfBFs1J8cYJNoRYvGUPDiET0MBHDFTfQ5zkD+l0ALXx5A+/FIwLNqGavg
4KdDGqZ/hQj9qzj5emT5i+x3VuMSGLtM7BagdUzN2A8/1PT26ZhWVdpEZ4+6RW20ksxagdsuOolW
2V1Ac1eycmtkoIOHHZ8ng4huSdPDpXWTxIJxIyuHJ9MyQGGDo9mUpyvrGmwejq2qUpK2Jg56B9wJ
IdDtJWZoaw81h9SgDgNR3Sz2E5eJlJ7qAxyWQiUzIH/Olu7yQB5U3tUingXDl9W8T/T0XCw3kTaI
Ll/yrmkAeDxpbdxxTLHxicea+kL3PUso/o41LZ7WCuFZCswTOta6Eox6Se83N4tKOMKvbFvqmV+p
9i2EpPjoyimEaVzOEOPyZ7IPKxs6dZj25wEd0mFYKKjus9JCtCkUA3I83LNVrrjjF9pKd3Kk7poL
oBG1bwFOt1WUDFz1ieddV3hCgvLYLtduhX/oATjdsZ+PN/q9m5+tzG7uiElcLNsy4XKv8ajUkDWN
xtmMkj4x2wnavnGw4jPODY7aMC1oY4x2X3SEC7KesnfmoNqpcTMX+OKXREUfd+hEUSATwpTGAAdv
oSXEBRcNuu9HF/LQuVccx4tB5Uj5ij1Ac9o5nCv9x4MrR6Zyc9d1k8bAAlZT72L/MzDo88E6bWtB
kBhrjBFrVJF0km5sHGI+2e9r4OTNCcn5O9kK+E76qInTeGMC0cwGTr5xfUliQSqOZ2AJ2QD5pPZ0
eCjazDA3oec6zl0IWkAx6KYrMqoeLPJXtI01hhL0CBhcEN4Agba51tnSPQinKmfEtiC/uZmeaNvH
ovAjslJPv4wXDbRansgff433YOYiLfgh+vb0M1o643N5Dkgzmkj3ca50VGCjKopOX1KpM/3Siz7g
6oqEnUQdNKsGC88XPPtY+f13ekZUZWlUqr82aQLSeWM+MAjqX2IKAc9MlA6GyUvRYZiw1Wvhzfb5
ROViT8B273SXX6KmdkSF9zNJqY5Uz3tvpe9u5Cwa82buU5CQvydSLA14LuizArhNdGSv5DHdnNHy
+fq2kAsiQ8zapyOqpt3NjwVSFCvCl0/Ff0xhj97Def1BY3VOENCvMSUKkT7giBtU9sQaWHcU6np3
8QPFahOiy70f/q9WBa6sKFzfnn8kakChFlMC9YmVbuSw/Ijo16Y4eKLCPf5KhvZw16Goj/jtJj4X
nqANW8XFM6X2g3Nsx5OZ6TkQ8ywIRFsX/VTPWo2yQsIBJDf+cYKAZLgPmQm/Q6dBz7SKFsSloWG8
x+B2Us0diiAURP5kRXJ060SoMCr0iGmPzB7Io7ORj42DUK4OTZ7ArHwcM1hAw0RGWZpyxEx/5lRR
BKBrZpcvEmbLXpVNkaH9pHiT0SVdZ1QmAe9t4YbNeLXHvd4rnypX5V9ilQdlkhBXccRSjQgN+IvU
wys4CaSUMl9mZDXiaySmZWkky6O0WFZiS+E2iuUVrljthBVEiwb5i8ni0oHSZALNZf8CA66WT0k3
4i2IRd4OPd37oEAQ8bHgaitkpWWt7bXjVARF6g4Q5rWM/jTtn2H1hK/nV/wP2xUNbGwdcjOsjqud
rRPqfGIRp3CCNpSi1R3AuC3s9kITEd0vTTzJJ5PpFHl2I+M75ImzOAcJTlEi2dnyV47LFX8bwiLQ
OmcFGJQJYWJhtceRtX20B9duFNGcmsndROgk/HiFhrisggJKzgXcRgoeZMfkgL9QdeK+NNXoqLU0
iWM0SKJISTAHlPYsqGgiqUnVJ9rZ99fCYCa/DlqOvMqyz3hEkT9hGZevi3S1ikGUtMraFJm6+6Wm
0AXM08a8OD+do6Nc0NhsO2LUwAzpB3N6TZWhu1yGY8K0gph0E3CSUKeUTzCeeIU2QDSS1IJ/1UDu
4S8GWy+gKcNL6u8QMXhjECB79rco2tDPl2Z4UAhkzsuVxb+q3bqhBJEJp9htBn0Qe58zCi5qxMux
v9jClpcUilry9Ua8Q9rkdx7phMMtsag4mHFr6kTQyilnvnUSfaD75Ptlh/qeg/iisZDtE1+gram1
yNWBBiEpCGb+h8o4pxLSHxJW6QIOJiTRCb02b9IKgCkUE61heFJVTnNiCfzJ0Lr07Si9oZmgCVVQ
16OvUI9Zzbcy31h6p04OgE/wBt8plI0cENRcIul0mkYwlVK7CAYr77x0fqHjRHKYHUX/foyZPnmb
Nig6No6CA+ZVBgG8RH1+g3BITZ+BEW5VvNFK1NyTNLpVocD6lMgRc3BPA6WVCBo0JCMqJNwL8PBZ
gxtmp/HY6bjrJT82iSqX+ovTh3bp8CmeW3y/Q+tx56rUwwlMks5IaTjnBbSQnLONR9rwQq7qL62R
5yHfb825hzlh8hsKkwj7+AXMmgc/9LgKi+8enE38omktUu71cSVT2DG3ueRRA4u0flwPppxurHlz
ZugoKASx6NGV5N22KK/17/z4gM4MPyzxNayLK3SHvKEPZs15fq5iXXPNncbKSWRB65JthJafGrKJ
zbIJe4HtTCXi6kthi8LCU0E1lYHBxwSVn+yhlfPGAsIWARbL8NFNlG2QPAcW/osIMPuhpC2OQ5R+
QnaSIud4wEx9bRpzoAaLIh2TrZYMKEbNadvhm0J1F1zL257bkstG+3dlw+E0fz7H38fHSddF6TNi
n2aWyo+cvAdMVffJZ8ULOWH/Hrhd+r00z66wzB1d95x5dp9tS3+jFIpPxoMxN7y4mgHXvTNUK6ig
ci4julL7TZlO/S9DEC/0XGg07ahG6O42DE6OG9r59IK+GTxkEazS8e+yb2wJx8FdBEUEA9lGYM1r
91L5Et6jqGb5fYRxVvbcbx0xxeKwaJeyoi0IgUtbjj66B3sg44Xbe8/9CKqx+p9w5rChKEVsWsZy
okpn3QMb0zBhpbR/vdMZBxeeJAN++f1zXnXDy0YxS9N/tZZqY9bdVrj4X+1+wfOrVfohSWXw9YmA
oml5B47Ln247vt1Jhr7NW1Ig3eArsFAXK22vT9kl6Dk5cLMyanUFd+DBgEkGIAZtopnM47utlPaI
FtaIF/jYJwMPacl0ziXQvy2yuSP8v/VFhDq5Jh0VQI/87MoUT4BfZGDEwu5iYtDzcRm5XxzmB04N
guKpx4NkHGxlAfKUW5taYf8dKyryYOk5yu4vX48J65gwsR2qbe7FqHBm9rpZlpr/rY4RTbDsRZYU
4X8+MrrXr8tZjVo72nSHWZntbLqOLiRquiE6HODqPboKqJM5Rk0TrI782FwaKYB4Ifn1IKRBN9aS
3+5sVayZHk8EhZgVErgRB7DW8aoE86b7AD9SjyG6N05vmrTx9y4SvlBavVKEuuN2dkjuAwNC3t63
4L/i7Q5ywbNSpJFZv3HlwYItjjgzfB4wKwP0/ZBmPVw1Grc0jMUoLiGhjel5XtZvT/PMecMVdFQX
bjCVijzYvtjsu4D8zf+JlqHRvHM/hAAJ/7At0vDkBTCxtyr0Z/ey23TZMqwQ05Wue/M5y06y4ZXn
3nqnWjrTKTefQT4cIB1n8lBlPs+Q2uOsnqRS7TIzxwY+6bMKK1NHK8glGsfIf+TxbiP6+V/wcnts
O8fxpR586weafeApdDth1lM02mK0eMkPM3qbyhbu+2sSCRozpE9C4X5oBjA7T3EpqrojifXmfCEx
v0VWaw0to8n/66aq9CrNE5xtHIB8FPvML5+JGQ+jZB30dD6L1R/0xDMFgLzjsZ1mKtYTIAWLQZat
uVS5v1J0KLtblEMBb14dNZZNn1RvNdTR8oqGecuHvusxmNVxevHoJ7/8dOLYNEB0PaIwgJ+nP92y
3JAoYyfNhatoEDww6W2YBcW0wNGm3hF0dIci2COLRHcxxmGn9JWVLY+cBmwVls+hrkmGx3NZtr9+
e4Gwl1ls6kSqv5J6THtUcxms6BfqCevqEVWJNZa0/DqU9V3D0qAOKUL1UduHqZvA0j/Tw55cRSYl
uL/zJTgdClfSEOXBlvA2DymaLaao9bv3bOl1qpURUTpVZ9V7eDzvK75q/TtEJ7PXznTs0p63ot17
WFniLjIWFIaKyE6K3E/ZHSeH4O2q5KQnCNN8DkxIQc9YSwFxdeOj5Ln5Q7bBb0/10Lf2ASaw3QQw
QT1jFWl7PJxF6ioLC+xHX0lslELs2Etj0tcrwcIUAwlG97Qi6KSOCVjhMLz7I23jOudYXp3opFxt
ctvcRhpQi4tNzuyIXitCViKu+QaRhP7nna0NyuarbnLSonhN5KE9JSFqxMps2uRr4nNmFlRRui3l
MkntxXOyM7EX5nmEne6GgEuSargZ8zKG9//YOuB1CCzUji9m6CaZmsGEBJF1TeSLAUpdHFHO5c5l
XxvNgtH5kR3q9FJwOdzum3ekcQdCGPhjTX0XNPK0fIo1dsVmwcSXq9cLyrTVyG4FwVtUjvIwuvqM
mIjqZeom9yH4+/p1yBlAQha+hpzqvZIm7/0k6DThtktvtkF3l5d7VS52DOCQQPrqaqulXgGpPw3z
Qs8HAnSS1Nou1XW3UvrmtqqjhiYrn5pXalWvxk56yRojb/jZksIabAwxC2bRB+IFN1tYbo7Cqi0i
x6eNvT5h4irUuLNZaW4126RMV5DbdRgLiL7Wrf1XxShkk9XdqOCyb7uj17T5Y1AEcMEU1YJrd65j
Lm7QbwNEEDeh40ystJ4ML32sq6rhA1FCU0IuDzcD8JwwaXqC3NLvyPEDqxfK95DG5ExCfQJZ/SUg
ems0ZneH13iojzJ97x6xh+2hFlPd0qBmqO0IHJ1ycNyX3urXJQK5j60TeT2Q19kJF7gLiq2QCbuD
QYAZIBdhHS0OwDVN37CqBVA1Zj96QINlz5FYrub0obBr+0zU9tQQNMaQ7b+CdYjTBxMPWy0I1agJ
hyIjldJMWsE2PIsNnyGznJ8Q8rjwzOWGxTsjRpZ+ELYYVpzJqwqVcmtA0j7jFnryXfB+E035Wu07
TY+Q40cVJTfHuKVP+sGgoexEzBIx9jwh92E9l6M9/UBQexMSq48q1RJ3Jrnkan2vbs+gIBbL0+P3
NhCX04hplrwTr7rBS6/mg3k+QLx5p4MmonP1WBHVk781WSGYqRxnzRAYHgvy9lbgi7bMgfZusiMd
4EWmojMgMseu+iKdioFElNITpjaOzQcHx8SaMCD+S5Xvrp/52ZdRKO3j4NTeDwyFNOus3syZ4wCy
4PmSYrruxSRjGLej2r4txSvFhV1Pj6IX7JoTnatqSbgjSMmeXLpqBFziYmiBOsxbYUOWhmB2HlLP
j793yjL9iJnRsGF+sWDXA5Lw49ivyQ6AaPXoU3x7rQVHJpNlHQgi0ITqbo+fZN23LYAjiNAFpOC8
JOrOm9YZZCgCMRL1u8PMvq400TgmJC3bl4B3TrqvduVqsAo4vVXUUVETN3Jn1GPuXkGXA/Y3NKkk
JaALBanlQaHZgUg4oIWJPtmieB2SKWFBw/jDzj8K6AMiGp25m19zh4Zy1mMRD3lWoVjMMMDfzU08
iVHlu+r+inATbxQgJ3Fz+z7NWf+2vm+royWD9sUo5w0tNp0Y8az1SylS2Y+2w6PCNkd3E+D5WDDd
yJkJRn+2vXMqU+kSPOiWFj1qTGnEdLaOTZu75wXvilxsCOQR8KcAZNDDZ1W9xy2MRecIML9Tsh7P
waaO/ymgrWmQIm0kdlFEOE8mKfSf0aU89Bjb20DH1NCZKYbyeIeFP4AbgQk9rPpiAKHJ6RUx9nQs
aGiSlDPW+f84CfBi9YJuqGa+z946Bko0oDgx6Z3jkT2dzlbCC2Ihj1S4+3b1w4S7WlIBu7YvZzlw
A+WTARaHCkUItN34daQDm6l05qNpNSxYOJkPkgJeI93f9PpTX/3ThMb4iy6Fed0Dm8QUbRx5DQ0u
vNWBMTp47LE063xy7aD0pnNGK5EUuLj1pn5UF/Ln+KgatJfKQ02lFy+eZ9GqSnLfGlBGNyEZjzKB
tPR7IIe5qswYDqiVQ44e/ibYe4SNWbOrNQhFGX/qbBcGajhXbAvMHiEo0kk2T0badoMjiM0tDEVv
3zv/ZApyll/EVuNajLlwTFPvi0AkEwe7NZG7PiZ0U05AjmTQGpT2RLD9KNTKVcXgHIC0MuELi94C
MiAHUYmEYP6mrmrs8VJnejKFvKpehKrpJ0cbYvatNEQExB/5ryaSi6Xduc0+aJgys+ZPKgl0f6yh
WLvCanNR7y5i92GbDTXGsvfu/W6NaHplDTAOelRMQi/TLABf6yFAdYxH216P3A3zk+hMLlNxegjG
uRsbNmpvynMyRf17q9Qts3l8n9bEDY8NbCKuHtzEFGYtGO2bs9kxvANrbHNc/zeaAWhdF8xFntrm
CddKYhr7xARcvdMC5jpdw45ztgOVocPhgx/tX50tEaPY8tpUnsW30RzWZhhevXfJFFkXKbY+FPTe
p6G49aQzHnefzGB8ZAuh3SmF6SrcxReXLdeHOhAnNyV0LN6mHk6AtuZM5JioCfQDx5S3tnCBDOy2
cnyNlJXkBZQi9pszIQ36LMtb26lPm313IaUpn01fcJTNCmVe9yTH3u73y8nF4RUTqJ+zaLhZ+twY
IKeBtbwQkZFTUiNOwDdthN8wsC3eaIBLfS8XhhVA1+DmY+DYoWnyX0b5mPXarcLCG1+WG1/FvywM
FyWwd4CGefn0vn8eXUklN6Ujx8k5/slnohhzsd0Iaxh16bogt4iOGV7898MlWMiu95cFziBEg5Uf
EtwoE0sd67ilSkodqMYOaKrGZLJ0E8XKWMZs4NA5OTIIrPPNP4FjZatHiA+7WXUJ97S/CfklBdXU
/r0rhY75ghPSTmtihHDxcQqRg+27d5gRCCawUbJNSwQW9IUoyZSbbHDu41V/wY0xYqyOu/i4TgOL
dkKgS6/we7YxH4a/I7ROWaP0LhwpY2idYb0kiaa79xhJuqCJpNMe7/dHCUY2Nxn48+RU8DL5BA/1
+tl3dnfZcGYXBV8mxPrBBeqYqYKJZt0LX82EcDF7UouKvIipjhFmeobSj8r2ZXvxzbUquRGdWKCH
v1LObS4e8VeCkNJGSLra44qye/MDIdPowZ/gnXymzrup11WoxSlbWuf4uq5HkNVt2ttZVauB+Z36
U88M8KgHKTEDOkH5vnHrfQruWgUNpMAzDSBjJGPL+v+Oo8wc4IQot64rPxIjhWAjafuhNj/kq4oy
1NaYcHqL5ggdlx0QXdEw5XCB3ltUCCoR97fIP2BSOf9oo//xB6C13u/mx3O6Pd5qwMg71ZZ8YNKj
8FFWSCl57tB2Nv+RKreIWefEITzkN7zxIUbT7sM08rhXXGnCdmlZHf3aIcv+Kdih22HlJ10tHzJD
0vs/b8f0xziTrvKd9J17hl2HuXhksDgF2LC+THI5javM6O0ZgsLPU6EixPWVCbyRce1/4Xt3SRDq
0Q/FqEiOKEmGIUDLT5u15vCATPsMeTcO32nBnCAJJrSQHDne47K5n3pJ7igXL3d1xI7k35ft0vgT
rTn1wazPqhLQbu2QK/Nx5i2MuEBzh1BAID9yZABmMI/9NA1Ry2ZA4MYnoJ0Y4YlaBzCyf2SX8k6W
IV+vgXOa2H1NcrNW+he827AFWLc1UN2DUEHchqWw++dKl7Ug9sICF/dZcS8ANXWTeqEi9a7X7KLn
ar+As8kuoVAePafAiLyw1RQOWFz/254alk4mRm3UgYgvKKOqgaEpWNdpCO5puwDuiYdTw4mxyncR
GggUfC9QwA7/dxW2Pt+yIFmqRlD1OE9sGDJo7Ji3qn0vfqMLlE3QoKGXBFRDX2Gg/MCAyTLVqwAH
ADLHzRwhyc/AT3CAv4nD2/oJBOaisjgjJrGx2Td2P4HzLH7KyOSoXjRUjM0kSLErBqtL2ui9tMv6
WuyxJ2BVLEfWf6JA8vtRMoq8BX/fv14AMK3QmAPjYNelP55vkvC/jp0R5Ju74dx/SNYdpsqTaljo
0a9F906616FcFEqw1EffSa49Ty8T+U7m14E/HavHyEfQbF0Lc9i5BN25mLJwhAbMLeJ6AtrYMEG5
yK7KUVySjOxFHsSX10bDuBsDMpGXT/ZpRQcDLHQ43hrLa5gMkNyF2eNCESrrpWqc5GcfOa496Ivx
2C2M6fl6rq5O/c8e62GpZzmvjwuxAfoebvcqBO4afCPFibol6OTVpY+KItPgnsYG4439ZRS9cmCA
uEgPinupHc+xnd+TtTDa9iQtzxkdprXkdTFqOAtNZjD8kT37bxDRfCLQmYDJPLTcPYMRGI/NDM+p
HKByYQ595j7I9n1yzYW1kwBruTFNVQZC3KiLYsvQluh+gJr0HRl0FFIXdb3BViwjkrxLtzsCuz7h
BcQVgod4cZ6NCvcBpste67vwWuHTIaubJCRauAc6XkzkqFw3S8YHhsLCFceXrsxoAMoQ2PhAMvX7
0h3JDmnK4hlTQ8vht4egrwgvvqEOXPHfPnCN59lGTX0rxQBAt2CM+VeDC8NlvooBsIiPAlnJSwuo
50kicOgrfBHMqoOhCenvuU99obDCUcr9N7JLNk3/rxoa9gwaOtJlRRruiS0+wZeJvI1FRAHK8poE
l8OxQyPPEgbsHRz0zRkbydSKZm5EbOrIwHyOAJePRJJbojCIaVDAKgar8uDvE1yhW6qMDQSF58bF
yblW1t2Ljd6suKFoddQ+PGpm2ksXFhjhJOjj2wulUwwE06gm1kBsP+6MkZ/oNP0rEG82AD9NuX2Y
TloaVhtvxySFoNzt127SnkUZUuz9986FFYfoJE929TQ+cLvPPHqbYGug2eulVx0CjsidxPO52bHW
fGz5+NKP6s+HeDus+rfoh7Osvn6pDhS1CTpdKuvwZnw/RIkSAuRowIGTsxOuLz+eZxQmY94xtS8Y
oNmdeT5yfKErz/BaId8nnzKcpr1Cm89AYiPSpQkUVRpLjs0VuL8v0DB+4cR3JkD91VDVki/lWzbY
LtxMh+J4oHXxg3S9ySfMOaEXsP+yjvWKZp7bJXjjxLgIZWU0rDCS78gFxRw3BnXOju2ZKtb0Mpmf
SCAoiJXVfNWMBToDdn398gOHKG0mYPca3xmHPX4Q/yGqWE9SDyykvvi1jJkMa+pwL/kzcYPeDdGI
gOumDfiCgkSKiQxtnoXC9jOahCPSHF1yvCVc4nauZSCmMmI7WJvzxPw55vpYBguFV6iBOcLRqKm5
eUZIbHz4A7L3tQc8WXlpEphx8PmCfPEd7sTwrTYzU+7oQLdes/66wH00wg3ztkUQOdisXa2EMFoe
aNHbgfkQ/JDYb2kHTilIE2QEfCEYd0nWD9f90kilVUMIPgoy1t01aa5paB0Ii1Pdvc5ADM3NwDXS
nK7fdepZckLpcK4KIv6aNG8ztp8NYbwZgmDthSkFA1TV5s2U6sgRb+hM/0KdaUtYJB3PEoA0+QKV
E6Yzl0afMtc/FekB8o1QlLclDJk1GYGBMFuO4WHY6LLmoWEj+XU/KfmYSkGpVh72xComZUn834fu
6REwYGNuKsNg3I7Szv/LNoYaLqpkE0ZZHmqhaImU2Uo97AneTDxYAvq/odaWdm95HjYgLK6j59ch
w26l9Hr7+7yVvAyuQOEwmvpc+0sh+hs+hslz8cUBgCiKJu95ikqDwZDdecAwp6Zd4IPzu/wjKtUf
mWqJVORJWg7u8XF4zDOHy1o3JLZlMiUi70QOeMCNJw++kbbQAgPHfLoq6AwvLclGp6zSwFCkkgvE
GJgkUuwth5H95iWWtOWYkuuozo9t7OCPcxUCUWUXLy4wFufC7gl+124Pf+A1la5vTsLZkwb3LyWa
DbCPQUVMCXicaV3elj6C+fffKKAXNvDhg0cnRPJPuSDF4C8lZqoQJ8BImh3VQEYs8LpdI3cezzN7
ClSfMgdlr2Y6GG3q4MU59cb6F/sS+2QmsRfIvzKJyoSuYd9KxUp3ipls2jKZG2XEDlxmbHoCIwa3
4E/LkE0hgWf+a3TEc6C24Um7JWIjZdcHll/1fRDdhv+zZV0MO7TH4TqAk0uccelt3OoZd6bE40oW
rAeNXhoCzCvtg5GD7lgJt3I2b1f7DjHdR+A0FSA2yTsTSlO0hOg0awFO6zkEBmqrgdJ8wtECHo+S
CprC7qTKN3Ub7gpTdcNLXKhUOlOfBJS6lYRCMxe+ATMDq48gaLRWfPSWx+DDRRS1ihhp61gc8+Kh
PzTjNQcVkzwajqAydJuUeupaerF2CdRZUs5oYW07EYCdOtQpJVq/C9Y/Z7Bfq0kcQyAmvr8ENAVd
Kekyv15VWr+Wb3uPMeGuIR2ICpfqGLJSiGKkoB7rJJnPYBhu4+Pjrk70G3EUkOb3DGCcqZRAZLGg
HRq+iHMda82BXEFlH0QuZcb2m+qOZfvMsb72nLYSeif/xUKDJ8KoW7jrBjjnTQqKotGfvopQzcpV
FslR/zOpsl+fm3qOME0ya3GTclpxofLdLdPAfLlgViF4EP6i/99h0uIKYumEwtG70SmAx6Bm0vji
+mUoB7JS/fErNqdWOvtcf3L/NCkGlMkuI58lvE7kPnmayidtr9/gg7RB9QqNEmu7XTLiDDAupLVl
egkjQJx4ufqrgM81RxOPZi7+zs4+D2TfrXLR/J7Hj538ES/KLUzTdgrNdiVSoRmAgBJN6JSXsyhl
rEbFKPcAxaVeay71GLrzpSLF3i8H2avpqtjpgGm/ug4XUxOssp/ysBWhTWM4AjIHr15sxjXgd7KS
dO0glGxCsSQt7jkGFTodlA5kXLQ1h6FapZzwyA3ypgzPPnp0pZqaVP7CQqz4G4GxxqSWW0j3dHU9
8QMWXtbDANbWq3c73Q/iiQZu+2Gj7J7/80nqgZKypexYRrBv0mfO59QZkElZpLWpSga8pqBV9FPN
/CVuLCYIWrIhE8KSLZOD9U1oXPATidt4z0YT++eOrrJLBez/kZJdEGXG5QcKUssmNpPWQi6RcT0F
LurUvJv1KoOTGIcu5RthCb2ZrJkmmhZj5Oiks+ilG3WVhedqfDK2+qjMsOkBbP7P4SgWM1710inp
+6F/koqyxi0KA33D9A8kFjhkOV/G4lgawsWDImmetELbbeDNa48gdHABNy2Ds7CavrK8KoZKJ7H/
TWFjrdleAAwRBnh0FzJYiU1Wifw2YcrQxXm6wkiOXwJ7elO1p4VpXkOKS8Mdoi/0iamiemiP3XuR
VemZdbWFrgGB/8uT5BfdqNZvLHQXA3Vzr8+CLCj/V4M3XLLNcFEcWyvAw837gqx0C/lMhcMgiUBI
gtHVEVR82hf+q5uZ82MF+ScO5EhSjHUkfcNirGe5VfZG2bCJ+F8Jd1fEby273nQ4IwZ9NhyBWmiG
QFsHjy9kZdhRnJIQP36n9uOMKBp0A1G+gbrYDgJVq/unNTV7ZznCaYHYZ+/c8QUPB0/RgKZarE0i
WpQRoMXuiErGEkho4Y2FNunTGmjIHprvb1P4nMBGU4LYZXs8hVLcW6PlDpsXG0R3t+S0D0Bbif+6
mSaLpa0KMU/6zU9pzEqYkipUjlXh1Vsf599psWv1XJiq3WCHSSFSC/6IUdHxqnd4MEyLtZpBqnUJ
F/voOHV/oWeAoRtIuUeKGF1z3lQyBgue9fS1ybKUcRLY5XvsmZa8EJPzJj6JrqbizQp5NjQAqPC7
sdzOCrxmtc7FFWht21o4InJARSG3flKmL81BVUhDgTbY8ZjfGYCpiu0J3p7Cn7mGEY38ODFyYGZ4
bGCojeZexSq16f2XBNiqEiYNdSCy9+ywSIdXru17l64mDxdI1SdbPq4ZUe1S42dCmzad8625cG5Y
ITQKgb9mz/cIc1SX/eMRuhDDLiMKSpA8PLqOko1tAFTDI0pTc5F/zYxcRBH9WssYYaI/7xXwYelv
4LFcJ07xgd5IY7AXxT7xhkccKz/KV3UAG2MgYSZLFBnz6SDz5WCUDizt9tSqkndYtQg4EF43adtZ
7gZkPwr9hDb7Hep89a6pbXTcccj1JKuJaEnmcjWZCZ3LCkMyd5atCThQzHHaX27n1jGJ4cXSUUKS
WD5+0XN7WlVRJUVWWq3b2sLCecHvMwNOMpH/SKBNkkzAYCWJu60mJnWFF0ABIXQSwU+OiobKUGJl
vhCgoohmoIFpHieLA9/+R0TEu0nK/+e4blUbAeMlq3oVcX57SP5zp+8Ci4yZIaTRr3iC2MVPWOa7
wxq2tv8BVxLSv1R6U7PpqZ8SR16VnybwA9rYcowOPrtHw5neoD6oyVlNM+8vYpm6/sUiDVgGA5CT
/Z/0+kVVpU5oOeMCHENmtEQjIJUDFFntcPzsDUg3UhzGLYQLd8s3hSwbCpTLLBEMOM7Cb3IWbmhp
0Ls4jgsITmDtjbOC4N4Q/VAkGZ4g4jGaGOEOnq8O6wvGDZv4GNdMky3YIKvp6ZWr2sajC+5WPxX+
RJMd55+scOgqkY7kCEfczIcrX75MCpTVolrfRH1BD54wlYov3rHJyYZzKFdObW7e0z/FQmYW0oYh
BP6VYqzCnmvYzwp52lzZ1qeBQB8BLjiC6IDFRB3zOk3z5nuFBypabWw5DFXqA7D8hr8PYkAdQTZL
+QCX1sOX1QFMYv2czD9EHiYiwB6BVbGwWcQ6CqYw6SSg4MKcNNM6+5U4+Q4m/01ueCBCht1Vv4fd
4F/yiy+LKvQ8mNviUm7C6cuZThnW0UGVnYSxnMlsLSBXe3+4HV/I8lrFPbjaZZZLWMdMAoblhRD+
W+aB40+MfxdrZF0TYhNMykA4/ZTTO0JwXZHC5RVK1e6tEOrB76GMk36g0mKgfqwzOdSzXrl0ru3f
anFrtXgCUmSPKV+pVS0azsYgdsLAbw/el7Ji43RdX93+uczAg42PRbUFnfau139x5hCuc/z57DmY
s7dRwqj30ojz/Zutbpj3dJpX7jlglgbmJsSIcpppceDXgGhyrt/+BlTa/587CdIp7de5p4TDpNZK
SS/0/VPfigktmimISHAqYIcxtSCcHVKmEZqC2RcUjRxoCuQQIhn/MgIuDLqWhEhZmn8YfTh/9nly
rHwyuzlEY6c65oK8tKof5wK3Q6n2VD3Bp6R3pLEaeS52lEEKYUmACsmrCP7VvWb5CoNBGSTdu/vf
hS63uzjAMCu6gySdFiAf89XfxXxokDKe8/Dy7qvUST3G7MXGjmC7/OFyV83L3lWp3OLnayDTyKp0
t3pbRRdujq7/Q7j+NPXs/KTEKYei4NjbfD+ZymTk0xBoJUC7BF/lkmpLLnrLBApBGzgfqsfIdPcz
EE2AI8BaS4jQu2pD5bLejNce4Xz2/OJV+Bs57UhZ+kZG22/KESbz/p3QydeRiwYNRc+rK+ybXKWJ
0U2sXpMLaZ+DwMB/u0udo9wLKrw8f0551O+F+7tr+mVrLlqV6g+inhuQsSW3cqYBWWFd6xwaLNHU
pSBuy8hFGWiIUQaPkP0eQPIZzQFdm1Yd4gutxQeZf3EUqZw++D/uSQ3H65ia6CD8h3NMNqpsFWbt
D4w0I4Iuf6GmkznJMkNUHQtl9pFS0f0RtRBuQHEXrSmTl/TfwcQOwQdI+YmIg4QXQY24YgMmi0K3
o9xNJjA5bKpce58rtYW+3Z9ZR/HxaGrPsXF7VIYOiwoT83MEPcalyFHLNTPqU+ZMeMifG8bzdjIC
QZHKZ+MC/63peu116WOdeD1BFuopgGht/v5jys7CGD9e83ZDhv6ESzLOCYcWHN1UkY8Ls6b5wLco
W8Zu1tQZm2Ilii+EcFNrRFWnwI5ymu5OYbLAggAocouTtYqzW6CKSW4yYyWKkjSxxMmzD0bzgQk4
+zrbSf9QjpMHCOmXZ8EJrVtkaeyQMfTcqzEN43xVvZx0XL5F3jeszvS//PrMgdRFOzmvce54IwCA
NijmPvfDBoHEqLMNLXRDBPXcdsaUR2eoMD7rz4iFxpvI+/JUcS7yvSr8dg4qO3BgvbTgC0VVz0Nr
9Ok3L/8DAC85R1L1pV3BhyDtF4xlo5TRocqRbXYPhcQzLvO0sBwvyCWeo6cnZDA6V95T/awzgPGX
q5AczFnvw6TtBIeMBHV9/bvZf8lCy3JWTxzCF/r1RJnkMp33ckZBARzB/HcR79+e0c1V9GsC7yxQ
AUHi+CHc8R7gTKDDwrSvv8TBe7fvsfwif565EjQ2rxCAmtdCCvmwdaPQZhRkLnlHsTdGz0mTKWa/
td53pjBM4HSZnj5zgeKoGYkxiae7sE/Oto7T5EophqPcwix1Z2ym4cKvs7yPo2sh9afLVacBJtYz
kzjyZ5R4MPCYJbXUgU2/bCeiHEpa1uPEWl6F/MsD4weICSNE/Akv6vCg76QgkuDOv4AVGPLgJV/5
Ye+o3sYxgBeZ9fLMGZTu5ONxOt2ZaQxdCRbGnQ5H3aEmrSbjSWq0BmvmSnpvQQQIIyo/HVdgrGId
zPenYxr9RuXyqfxfB2p8HasUPyXy2Kbs3H3k46jxrZOVjx+f+yqdW8r9X4gJtr+nPcDVpu8j+cAt
2klUdOJ2EXUvNZZauvkho57DSNLdd7tCiOFR8DbAVZIYVePAGx8rU7ZVFDAqvWBaPdtMtWWL+r+M
9ZmtqM95t6RjXAtfwjR8upBBqZYEksq52PO5SxUHWUV8mmJU9cBrFLWHFGVEI4Pcl7whBawab7Lf
3hMnKyNGW2CCTNyMq+Ldctoyt8YtV5VFdiUYLagpd3TzvzEcOdVOZ3YZZlxQYtTlCDToc7U41+Ph
huCHu/yVD9FlHHOUYeyLzwOcp+rWseLj475CLRgNz/k/zypvp5UFygtNUoti5zHZE41X8PEifDE6
hAPunIjwqUFEja4Emx5v7KOcAm5iI/NZFdZ1Byp2fON6sx0GJ0m9dzqZFwM8fK4ir/xmE6MKnZON
9Vi0QPfsfoXtNXlT3maBMWslyj/5kccgR91VDjScdl8jrI/+VB0+7tB7DbQ+pcASPl+S2Wz+tm9q
OVnisdxnybpE9EVYUjnkk/AqRi9Itil59P6dQcJCoD0UZE2tptck00WQODKFoUlUhItlDyszLdXe
/+5lp6lf994bzHvW/hKhkSeeb4Z9iQM2HXzAXd+sesEaRX0GSCBcBa9evkSvZ3eR/zyVu4DknlRR
oJm74VT8Zjc1IzF8g4WfvAzbICj45/ud34Wq1QTvD17Pz/QI7YtXKRwk+tQkiSYf7Dz/10F2U2tq
U56+jwX8VmnZb356dkjIyxGfsYQ17FFuobDv+2Dwb5HnYyfBwCSVobKz+yV/5n17GhMXQOagt83e
MuYN5t++/IdvJnwMrKmLPXLyGxrQy3+PsF2c8fNGGXDtnVFYUXSi/fTEs7iXhxeODNqO/AH4D5LA
LMdAVMknXx2J//ET5zykYk98LgDLgKeSQS2snY0Vw9bE0E0YxPqwN3QZ5A15bMHUqab7MZCl0eEZ
D7dkiwdlnLuZAVKVIgBPWuupB0A1GFV7AkDeV10O5OXzrsQ0MPx/zslWLAcX0GZiIHtgBPBE781e
osBiK+fpjgXfzirOCveiMx1v3dCAWg1iWyjthjrIFfavBRyiu6ztFhp3zxCYQeY+ARPzYAAuSPNH
WeHEdDaZXUbX7TyecdOmSKuLRMi+axzsFuWzicV1W9eqxNIBx1foPspGO0XXDtQtz7JM0epgSfMi
ubSMtbT3mm2j46mmh8Qujag9TGd4KUO3imWMAuRhuZO/epMapyEm2DatDhQvOcJhW09/nxBz6aRx
IUab5peY4BKEj3/bwGfTvXWS1uSEi9Rk3sWqPBpNKagec6z/y2uhxbBuvSnWzpfB62NtYohZwvdd
MOAHC3iA8zZWmLyjvlZAII45AnAdmiW601kwo57iem1hdKxPEkwU6rkI1qk9D75PxgxtQ4o5sg8W
F1GWJPZaHm8Ottm8dmudAfdwDBOyytHsYiCKssfw8J9UT4X0f935iaXMhQK2O6VkqXyTj/OGaqOn
AIbaPRjTYpzYXkJzCwHD61A6FcnJpF79pjpicg2hPzsl20cNAM07tofTAQvZfsgRQS/qySMwc3V0
hTU6veCqq624b7+9kcpcAYHm9+WJSyDCNlOf7jU0Bgok94Eh1uLU6feuc82AdEtWMV+3977Fpkb/
MrefPrNNjBGgQfpmCQh0fK+VHYYoxFEJVBAMjzZzIucLUZHfhxNK/+E6XPJxHFASnz3CCTXuAtaF
pcN3KJ6UelCTtDglxcTb5DLpe17q3xYjjDgv5AUGkmGglNBkwoHp44FLotHjm26hKf2/EEUCMZ94
ptzMXuaJCh15ZNarxumE2hKESyVAep32vrlJZdLAVPbiL1o1UD0ywNClD16X1r40DJOWtfVtVQ6s
aR9AhEJtKsZoI4MIT1Fu6bBWZHJ/o0Tb4lBHwoKCrAvGBwPyLtHE6AqUMKMrna3JNVG1arRaKUQR
R2FRaGq0xuOx7fOiHH1dnNWxoMnwbhhoBXfhlEhXEBqWZxK9zO5CVOBdjSUDOrdl6MBMGg4DqRSK
eLOrDqc/k0zVxmGwobRsuEO0q5154BGX6Epw7tTAc0MvzFhlKefoiV3IvvnsTknJ4EPTGUEw3sIG
6jzQMzdtepp661Rx907cmRycpyu9Ges+9Lgzt1Qn0yt15O+mGp/0OTw+vsfGj5wFgmVaT2xc2wgT
JkvICu5+1cvKO4O1FN56ztOyiIf8Pwi0rSAU3Ig6qpzIFwgQaIbujA/BlXWZHV40c+PKJ7nf7xWV
0kHXesSm+ZpLWZFf/avsBTfEBYto2C/3Agg8jycwusa8jxd4KljAEVIOnclQ8xKjqjOocNfM2Rag
GU8DdFRnmlZcsruq+nGkElEztwQT0ZG5KFc8T5mBjKmyCj+CfvFfOsRwu//jEtlmNtQ6ueQM0PX2
WC8jBY+1SAFtB8gwBoEvFtNG2f9AEBnh4w4diu6OFROvc6XxiieUvi97lnVED7fMG5FPhoTlqTZv
0hm1HC6OzDG2yUQcSJx9BJeZOkxSg8cKt8OTTqqwr85lEpw6ZXxlU/wiA8mgLuhrdhGfY2JO0O5f
k31+nZBFPlJCCB83noImKUqn6WzLOHIhyJc/9WH0Q5uEXWdj8zpb3kTx4Ao01DhCrDVcxL/pQYga
XuT4fXb6mbSERhY4zRiaPJ+6xXxT+896K38JufHidip3EP8Q7xYoVSqqSTusPKD5dx92n/BYAaYS
6ulVsamd+N5K4/I64wY5Qoo8shPt+dWedlzX7X6OHACmbF/DR3ENjHQkTiqAC70zAfle0gyIfrag
yMVfxpBeYnZK1hCz2+k1KWFP/ue7XODzvnwCRRDKgF7bi0S+xXg3mQhJLtFbF71FVlY6dTT8CO6W
Ah0fyhY2afq+P1IJ6Gpu+uJdwESOoqjBDif/MxGzXSHWyBcigOrzp/xqTZjwqcpBdc2xixke+DhA
x5bYIYwq44q3yCi27zobBOZF4HSRf2dkn79kcJx/wTiQG9zieJWd06v7GOM3Q19aTTUs4i64yV46
ijT2EEIkZ1/nEacOfoQNEf9qcqv4NDdBZ6N/m7arH4YcSzwtPScZx4rEU/OUi9mU7HMVe1MqLkZk
pM51T0yZFgsQIlON14STJ3FAgXeMiOTAAY05UqbOqwXhCzvQck83pV6AmrfeDmfgf45CwBm9RJQe
44habqNhPDoIROke5dBwckJpGGUsCNTY2iLVYS++qYYibP0y02t0zd3ukqNsZO9GlJDFlDuKTIyb
AqnoiECk4Iy/mVWp8ytdghaLs+N+kepq/xbUeb6m999QOTiDqzODAxRARraz5csNgNN3Ppd/FwZ1
PEmwnri9DYvNAi78FYpEkPxSY1WCO0Eg6xbfMR204GALRP0XOroxaaIMpaCwpX5+ZOENij8bnytT
UWVn/+9Gx9cwTuQ2FHgmHDcrtcdndotXdQOUF9r25r92phru4+F0JZB98aeb3JSC/Ybx2j4w7Zie
Eca64xsO8YQdUrj0YxLBGGxEs1DA+1k3H9Sv5qF71bSs0D7BPnvQhzN3nIFM/8JGH5LrGkgCBebR
ia1bEWU/yQ9m+xnVEWivgbApy1qIlyEUbD5dGi0GgQIRERMzQqgCrYJBg6WHpR6rYPGCAWUIkmr2
WNknUFBalFpXTogOiLHI3jLmt01kfUfyIfn/DZcOlDO15UP9MW5aOrA68ryzEhSxbmVQuxYZ519h
d5a+bxJ8GoRQAnfiAOuoEUxAHbkzOteFD74Wl1NtHIzncyPRoqsaqMyb+DaZ17gLZI6MmYEENGwT
2xtlEJ6idQRR6Eu6knvl2WnV7k27njUMMxbLTrbCfG8AfAbhxB34r6751OEKgHhbrmvuc7A+G6U9
FP+T1Faz++tmHYofS4veaRMXPqccZ8HiI0lc4aQoppzLtbcNKOOsGZMlLq69LE8v1YbXvMYIH2M1
2CgkYaRIE6kUjjWc4CwS2NXFj/X2hNoz4wqOnE2XIYGvaBdUeJDrqG8/U5kcQHQ40zVabecSDFv0
4fXH9ybIRm9BArTSPME+yRkWPTTAHKXNxitBTQKwYRIFNxppeDvtNJVz9DDu8EJns0BQYd5uTQhQ
NJhDmPJ/sHKFM9cfG7JRRKPLCmTULrm07dJfSDhawmXe90orsx5emtk/fl/SSKZJRBGXLj72uB7Y
P1ipqHVwvTEoTNbeY+kt/OucYm+TizyNfATBAT0y+8GLStIUQmNbyfadXLegL9zN8uVn/w2f87v+
qdc3ZCd6lPNKGzJB+UkpsOJzqf5YF4NDytkTg0OSycUdEF3b+E18xdNTowHaiPDajAtvu0puz4tn
eYJl4c+2sGfb4zVB9hbqIJz/klu0SCJenhIJuh8AQbdAekiyeCpoIk8nlPLTPoZNanFqou8BDRYX
I4gqHb0qiy3IAIAOWgCdH175jOXFuu2p+ZRZr5oGa2C8iD5Ee6BIrS4Trnnmgd4EonmqoYKfNx6P
wbPh8H18Gg3mAqCbseYnmcBPy5npiNLk18AqgnQwTjS/DswxDUzBnSGaFPOcn6sOuSWg3Jul3a3q
PEVc4gGcYQ0TckjSxFa8WbwvFM+HUHKTf4U284uG13cFvsXSxsbVYA8LbgaNrhqbBNR5Cu28OEY0
0DHCCIuSHQ7KNQVTSHoWZJ+6Ur0ysnbNhfHqUHguGwSEbZgQCPsU58zlJmFOTB+e5buxUltifdbY
qgSaS/OeSxMlpordkKxe+E60IxtnX9T9unRgFwThoFmMSsPA6PVbVCRXnVXJh+Xoa8ZI5xGSyX17
0YK1B+aQoT2F/6/S9jAyJgfbxXdd8CUSX9pnSE67zCYUnxYsrEnUvBozIvaZuaPi64s4TzUD5aih
zlNNoMYuZyeBfRkOjK1EpRJhjaEj+zzu5GOBVkEAWegsarxXqncyTLWy+YvX+/Oohr7ABMPCaS/C
pCj/IESYB9EDJEvIQfRTMy03cHPMEE/UyHu8bsHTD/9cfDrJlZgUI14GBEGycBy4bHomCHBtloZe
V2tsEiV1j3WzVC0M+PrWxpjr7KYkqT8w7oNj/lED2CQ/B++eJ2TysZexO9IhKhfic0U9aaOdOBAP
pn+pfccjF4Wg8ShFfAzv8neqHyIccx6p+5m4xmBzbIH3c8kTxj7wRhgB+DgwUfffqEc1sAjiLCdj
HkBeuK81Z6Y2Kb6SiQYwHktgnqONOCpIJzj+ZOIRXqICCqD4PD2bBAKy3/GQrmBCY1JgWEntPXio
kFr3wU8TTnDXgt73mlAi8try90CExMnvKbJtk2yXtOfOm1f00PwGT3JHg4t4dzMdKnAYaPYlg9Kz
ZkNam8kfB15iQ1D3zLLCAdQneg9W68lhaBAHzVbUkkhQugOTHaX5Mt5e0b2olP8e4cMnPK6FNAAD
CKnIHSLViHnozqs1n2964EYQcbwN8vK3gwr0DUy39mYxijkfAOCs+SpIqLG3ZcQcuRD0Sw7OWCV0
i/NWCrz7PXf5sFtZZOm8h0QEkCXqtjezO/jIwPoJBKgnyXPt5GEhedKaZemcOSl5edjkRkjJ/WLi
BFI6zLuU0x/lduHGSX16uq46om+n/mmBq6j+oDblXZ3p+RxD8EgyOKQUIHWCkQL42cOCggOkzo4j
BvN3I9MMPiZ0yMms2bOTBB/1GMUVq1/CZL3RkAVkFXWL5DifZRqcnngjfW0GYA3hus6EtJ+Ade7y
GwiBEA0y8ietEd24l9Yp9LWDiYI9qsMGEbpo7+jvyr0O6YSXeVcaMwPK/Pr6NTj0MqZvv3wVnaJ1
FvAf4fODQpoAaNPjdGilt2h2u6IfTWUK1wHOc/Lw4em8GcGJfjKbLjNQ/3Lr4RBHA5ckGJjzsdU0
cEnzm7hx9M6MQwXVu204dSmAH+MJzZJ9YXYpbmc92i7JGhww9vBsmqjCMSXkP6UZgYtbX+tR4/Ui
KaWdm/uAwevvFtoTU7ykPybrHkycIWERKewTfhFcGPMdd5vnuvlC4q0KxxGDHLegcXFoRSyTYDfq
KQLGF74GZnDqPi3WFBb+iknlzUH+qdq3r4NVLPQ0GkYCjCaioIdeZYyQKaLUJXLiLZIBr0h9LywS
rTHCW5vI5dMU+6CLowROIn2LM2aXnoHKR6xvCQVNynn5bf5j6DvS2w7LchUpVBTe96CX2WU+G9cx
zsfyNApuWsOsZKcuK55zAH2NBtUsFNhYV/ZPHqYus7ykwuzz1qi8MPXv2pk3BORb5+j/RnllHQD1
AZElIgxUmqx8QtkyDSXPVlDYCvz3LjGBDgn5HjZyWRhZ2tPXzyAGo7KRvbM+VVB8UHBH8WT3Dc7e
f3xL4X3mROsLvZuIKt+7gXthUSNnqlhvbLuVzN1uTC6jokW1vv42KLyYXan1SoCauvvw/8zKFrwF
BZOyr1eFyuAF/tDlrulP8MkJk6Xk/0yyLIGtErVI0TIo8c43B8HlILYn83RYkcJYYK4BCgAyVYYd
QQ3CETSc5AXclhiFBVge+nQS8TSbpLFkSjJjcukTQ7CzbA15COwyRi+I9rwPuaXoah9qgP2NcMps
F9zVO92nBTqm9B4BecROCHELxDNraMVYF4/V5l8S60L7G9loBLyq+8ucPPEBuiyKVxMG68RN+MPS
VDm/HnleHrAlvRN0wgBhxsQBGbYzAJNRBROqcdavaLD2na+UtvBwuoybigzBEiOyS3oBuirlTc8/
YikjjXq+1L4b137dO77S8Cp1OsHSkaaPcFnXijC+I2holRGMiyj3XL23Bqaw11UfZnjVU11mNb+k
cyZ3660DHhwsd/vjBO0zuKi5ni3bOkIF9GWFCpH/l8a+JM5Ur8ONeYqQ8eXuf9mV3Bsuqk8rabC/
fxFY7YW5GdVlXQuEnuHdu8lXv5ckb5mUdmfExrF8LKbstvpx1kcSdtgh8nPANy28E6u2/5OOObJ/
VkI5kFJZsShvkTbUcFbIKLJ7rSSkdAyXlqMh7aKdW+Dr07IHwH+ZNJfJelYLIjDr4zvPNTmDIlE7
m1JR3yuCoazSqYxtyRUTVeQfpPIfoPxbsqO74Mx7vsm+GbDhxZyfPdJlwfGw6sNL7kw+Abkmjwon
W+zjxIGvjLPhuY1gQ7v0rVRumZ9AIJFvHc6n5I5axhB4fbbMLom7skQe4fPsyBeAI60ZRBH+ohzK
2dlZi5nL7tYV5mVcZ1ET7CFgsr4pH7HdMBpEUhO6Yo9rsmqigAYYgSBuCekQlzJBbmSkGx6snzYS
n5PHgDXHnkfW2fFYRPnPM8sSDYHN5GGOGHfxPxNPcNWt2EgcAlAgBv4OwxZRtUPkjCUv9J8RddAq
anmIaN7CYcLRP3/8tEcG8TFfdIOd4Y70THnSVPxD/Ax6uAo9DjvbvDQ7sqSdzTGjyGmuZ49J+nBK
Gx7X7UTS6/oG3UzlnbfU71tP0bYjGx7+I2EzZVdn1Ed3EYdj98pOeWWvbB3727iTEzMg8CA/ogSc
gHdqsR1mD4wwpusT2YQp5etzOJ5TPzvo9l42LG7li/EBnH2/f1GTWx8A7viOFOY5uJH3XdPHYkGa
wvm5jOClwttmBH1AqWratEd/jdmTQNzfQs+z1z8cnNtdVeNzRv6kF+amGUgHQneXwVddbMUaMZib
Kni38GUsMWiuyfECvOI0FJ3dNLoN0mQKiuNXy4izCkGsczCex90XOv1fxnCN+iJ6DFfVae21ww26
uKt6xRWCVnlc0v5kEfuaqwVCUzvBnHTb+gdiBO7z+11PgaGxu8o8BEqnUqIq54C0zgtJecm+lfsq
u2nT5y0+S96jQONaKXamW9QBrnYmWmlUNOhmq1LhtMCnAI0TQSz/cj5LgoaEMBN+B8fZ9rVqx8so
UaEZdRT7QI+P9V7hFtcnreSChVgto1hd7UyBE++K851Q0LayqkHjyyoLQjbAm7TQ6m1u3Mft8vFr
Uoc9rWRVtBRCoh+eaafSsfUF2+T+sPJoy7a6d9C63C+2M+8o2GAM2paDcRkANb3mat080r2bIe7Z
8uFtv7YjtLvI7vf/ZLU2trZ3Q7eJEkSH957R/E4omErR1f9+9GyJ09xIxZ44DcFskuX1Ru/GzTy9
1z/rz/U/gmB9Ona9zuKINcNbEhD58HtiJubCXnMgk8TR7KHy9taHYoyM+B85F/peirx6YssE+ueh
XiFdAEJswcdcOpe6+/LIHpTvpfiWTNdOLTxVSYApKhWJv2wYKl1s3bu5DZtNr38OhZowuvN9sd3t
JfMtUg8TYwRZGX38ZNfvLc0IQ7E4jzCYCTdzn0uW6mvmQUvv1uSHJ9Z6cS4JsW3+ALQYHDuoFY2I
WdaPuXiPZ71vQ2azQwTlIZBgMZ6tLSNYfmKYG0javptNH7l4x3C360s11q5flFO5V5hrmCyPMgBw
E452G2BQk8htLjozwiam30jqpAs6OAmwKaDaBmJm/ElWiwUKVkZKVEh18CGB3nY5Ln/9BcFANIL9
Mx+7W3HxE/zitjngfI84RUQy54BhzZCf6A2gOYO3coPL6lvGjV5jqhGRug/wRWBrsOpIAHCDkJgo
9G1e5DhcTSJi6bDDfnFn/HILWHC6Hq6UfMkF7WhJKLPixk+Nu7ck0UHxuTfwu80SStdJI6dQ4Xj3
QRTtKjYB3MPRL4QyjAqEjf+S6FLDvWbfzIkavYTflvn+sYlzvl13FPqVZSMFqW9q+tmdzMxdA3eI
5Td+uGw0QTpYmyd3XdDIX8h2Eojcc0pCs6V37d5gyoOspPUsg+QkMa5ogZh6kcN9D/Ib1iB9xRsb
LpjgzFtbpZ9DGNHiOXtJ0DCOv52FmnulAp9zNuSc+6Wf1kymYgu7li5EFAD0nbYzh862Pklll6QO
uVa6SPunpdsRe0Zj/7cQvIQQrcwSC6+Y+RVz5t75w0rJuxysL01tOzsVBjX7t53OctHo8B/msuL6
uOn2w+zyuxAQXHHcRRRdOeLk0Syh+03ANRKM0VZ2EyNTMc94rWS8pmeV+v1hO6NX9WUQjako3yVP
dlixVAk9wZhGfJ+E9Oqoyxohw7oH3mc3BGktM1jxQ0COJQM9y4MjaBFVG7osag9WSLdhKKLERT3b
13rWvPrGtog0wSWz+zVy47nmZb3JfxBABMyX3PbsU6fKU83WvPUBpbAa19QZGAo/Rrn2ooiD1J0r
VbQoxGJxXijwpFfkTaHMBdsFTcyiTWCzInWef09rlVHnxA+rei2m3am+WJEZFYa41nzKKQ/0ytUB
GyPdSx++5buJ9A94DA3rVGP2iVh2XnuKe7fLrAAWYK0yG0XJr44I+0TbEWuECgj/4ybPKx51bvR6
UM4AJo2wVxrPPhvGum03rnMmNBbIo3j7tJwZHkq5VsXuSBBL3QFCaFjmL1UOyLuRsEIsDGySDT5V
O51bSjF4m0pw3hGQjPVOY+ulxZvfbWDOeWoP32/MvUqpg+vApQJjF75dkzG/O+vIltPOYpfa+Rib
Rl1ykX9GJbJXnZbBChpimmsmP214ekM+x3Q2GKPwUVrct8OtAcZL7JA8IpT15YKGJdnPAb+TByFJ
c6MIeK65xRfVVAyYAQsSLBEqZX4ZFbsXXMX372p+pY2QYf4GGfEMMqR9uHpke1r9ujyJ5nL5HGIH
ghZMe5bHeWEfz0FjqG5PBLK5ohg/GAZO2Q2KGfkRpu5DeyfGGG9FKZs6jEKLSyViWjSNGW0bpheE
6NUQxRInFdmQI6fwIDREJ6FeRRbQjMn6RbX7OcJbW6GxZK/y90Ws9xa2l5SfhZOEFTZWOmX+r+BX
9vDoR1FoA1i4jrlyZ4it9YgPplVO7dbm1GaXluQbWT5ksKt0nDxmgyvxP8L3zWtyWb8mq+AYewoP
LSgjZ44KGX3jaTDsy6bOroykCMwmky+zXKUT80JXNMyLhDNPQ6DbEdHniNBovlS2FkiCKjupnkfs
mwWpLuA+tefj1QhzfpRLTx+5e9sZPzcHbPa49uA3pNRHz20PNBH5IXaovoelXksRAEsnwjVb6Qph
bdjcrymzmkZ81W2GyyNDTCiqvY6bXsBx63ykruDE/3SCHgrMXOfWhmonwLHWL/4HGDrJjYQdw8Da
8N03f9Y5k5FMK5Ph4LxmJCjDyA4GZnsDFh0JRuevnspuBLiqG+0xrSmKU7rlX33eUNBWAQ0H03YX
tXSkOtfs9pas8HEVNYlebJFOmQutZ6+L/57TD/wTzlleBl89kdf8ZPLwsNDb+GFtmD8umnEngM92
N+alk+iUA4NDWxqHlNxbWOvhXBCRyOulmwdNhLVxOg5ygH+FMl9U2WXOPK50Z0HVueY7Qje7nBRr
016DjHeFjKxJd4Td99GhAA4PYizDDAedCP8RUU+3GtRRSu47W/RHDqSicFBho3qZq63u2eY/nckm
dC2ZbwbNrw5wuqnaHZ2xbwf8fScJbAuWn6PsFdSANLn1yyTiXbIOWO8pD9Q/OEgp54ynvuMEObPF
PzWkI21G4MtEy+gBNsQ2nRnAKB3DWYyI1NKlyKiOUFSKEwJK5QhvD8UfEXQHz8u9Ka8Q8M0iZN60
DwHfmF/e7+ulrn+SU7Y8b+eX99oTsmA2upxRFx2sogW9UsQ84DesFHzoohI2GIYdpaGllZDOPZYn
zolzKbmT8oP/kKwIZvc+Hj7aC9Ak6Znyq84rPdoscjQSj2ZB7DJPIE+jcIy1n5E8piGUNZEd1TFZ
uw0nvg6OJ2in4nQhtrRrVv4X+gGq50qf976lx3Ov9iJHC407fdxZrsz8HSErPQUiSDRmRfB2ILNr
NNjDRegTGO4iIHnuNe0eF9HeSoGKeQsk50tEzqAX7t22kJJHVbDXzFydSvhW8pu4y9lxS2HcJJ8I
zrYbis6YPhZTOiIQSiZYkrPyrMkCNyNoQdc/UZ9nWzBFJdZ4+NXaOSpExgGcH23RNL/+fGTsAQQ4
Bic2QAdhZpGC/cbSZzezwmMq7viyHK6uhKco7lcqVScWMTOA4kDciV0D11qwdgORofHCJtQGhiBQ
44g3busQDLsBti0BFHOLCGc+jrIEn1D7Jn+m7L01Q1NqBQoNREDiSiBYIt3Ejt6Z7VMeydh3wIvJ
H2gbexPF670QXtYYpTrqi5EsMHkEZmdwJYmJhSoVuDOxkfeMke3OYRd5EpyeoOTZ1FL7cAsDfFgb
5W4J/aC6ru1/6+GSOxeyhM2X9t0/jXSX8te1zydFH6pLwTmLP3epfqR8ezuufOuLB8QrGLDQnHz8
B9izZZjrvx8Q3I/Ng5FmMPebu0nlM4Akhv+IyJOKgH2Q3282nww/UAJFnrftg/IXGTKJPIkWikkr
CG0QlLAUHgnZzMOp577UQUzxVOgX+UiFC3AmndZPcyWj7AFA8RevvIH84d8yizdQEmpYnNpGCn76
PaiA9pGzt4Uxpizvx8JfDeH4tXPM0+VgPaGzCjjuhgcgrFjkplzjozyrNDeuz3j9U+0oZpu8PpW4
/jlBGDUYqA5PZjCskKzE0SewvnV+rlyELY4A23sIr9IcyfT5dhxZK7nv8kTuFdafHLeQibMMVotN
GBWbCTYO/gDG/+/SHUqbGpzRSM/yuqrF3SrexAMenmoLOHZGc21ahIrLXHoKewGnPMriITdSCiO7
hxLV4ksxsGxIxoFZ5JIh+38Xeb9vanyZyuX6Ty4bmZeeR7lOB2JCTngR+1D1/DLxv8rqbafWMLH2
uIDyuB2/sjU3fuAYiqywBvhb8pkWIu1w3nEkvZwhglKcQr/R+EkooCrM5RtAIh/14Ew9q6kfaHxJ
MGnFWEMKbgYS3LvmiHelAAyXA8KQ1uCPRBZDfHwRMuaCzmFuwjC7NwyXaEqG4ZA9vRs56tBDWuCT
EzqGXe8JL81qV4FgxP6tE/ry71+upy39QM1SRYetBjxou2nmFM65QtNpAN8F2ZcGWNnMHkLzTLeP
JXhz2pFV55XWcE8STGMM6skp1YQejncwjWKcHmkUKLRoqfgZUF1Zn5k+Nkbd+KiWb35NBWf2QQWo
yyLvdo+Iv7dXpNhVZYF/beql/MdWKZL8BEC1SqvuZlJiEaRovuPAFUsYTnVjzlWwtoR8KKPRQTR1
GmuH+XNeDB/simEphkIyPn3Gro5riPKG5mpURG4db1BT0axBgUbOXw90qguWcXrtINhfxfB5sWK9
jteewbnx+FtsHKkn49EJIDA+4wDPVcSopfwijZ2K5IgNtdeYMNUFRGiuMtQvTV30PT2VD1DPI8Vc
rgI2zYpzo00bfSGaBmg8o35J+harOeadLji4s3ior7AiEgm7NDthbfDj+a0f8B+iB+fZWeKGilKL
qqY/0w9WhvIlw7tiDTM4RVB9jy1K3rCf2TSveMyo9jfuBtlpgpz12kKbZohpyCJ7rxzpNF5qG66F
HnF5D8dxXsasUUfuSBPr0qhX3vijNCetXIIfXb+YXFjl6XYLQFOIdVTZjNVjJfm0ziTyoIQdHFsK
7F/1B6qK3KKD41NZFz5K3beVvjlTiwb48IZJWdrRN892oNc/5lK4klbkGbIfDmJKrvC21R6eWSlV
QYFthTvGwVLjEXGKglxE1LXUT+rZDTgLg+UkRjUXZfvJc8IlKbrEyJjv5h941h0M44PouCaE+ksz
Ndcao5+X948jM3Q03EHxa0j37g76UamNnyJVIF9Xuo6d1ArUWZllFYRVgEmvUaPbZkoBgjXkDmjc
mgK1m3LEu0g8KKSZ2upeRzIGbvjFgEYSYvjl9vOcUjPI4w5g1jQJ9ye/s9JVW+HycbrNFD6PzpZg
kD5cB3AVBU7RbPfqYagrItuPS0fdXcNHkx88shVZdu6N0thf+uopz5Ut8K9I8SKgABKbUt0JPXI9
b1dC28adf4JgukfJgsiYVQQ04zmQHrdWEyMpr5wAU9dukb0RjSWd1ny0KpY6RmHiGOZjO8XJ/L7R
1o4t3WRovbOOVxvg5rL/2McmZiLQo2n19Q5pbpDIwVG7K9qKmKeogEVtwWMza0Ag9VIr8RUxCt8Y
CMugs3+ZUg0VVolR1Fuy19opeLVRqJRe2AMnrSse/aEizpCNeJe3bcyGDm+QVcSF3j7OMYg7Zwpv
tf/F2v67/hZJYzCAFFdAKnoMg5V2O7/WO+btegYVJN89ATwpYUsFbUUGTFwsREhAjmsVOxWJ7kAY
cnjWFVqB2ih8n35e2jOqpOoyBOuuk0eaTBoaDl1J3eEAa5ZRIyr5by58S316IZMpIJBESKmAw+M/
oV9bwboKxDZrxo34TGWcR+S85hzyVlYW7Sxjeq+zBXrgJ6sPXpRrILlPTRFjtrbbOYJ8SIBHfw8d
O2BYrI3cQpqqina4DEjEOS+yxGW78k1fbT0qkYwAh/qM4pPLu0i6keuBpAOWoKNq+cqhVSX+PtmQ
Xg7/g5yfvcwX43gimMK71Xr3Tkn6qQKkm6AaQu2RIPWkDL3LeNOqkjmHuHUonmuBFbXsUsuEW5z/
xUHZTH4ijJUJ+fCG4q41LbXShJzp9uqKwHpBYrNs56r2XAbJ+5NdQZfi5t0mIyiQoP97zs8ojWtG
W9a92OUorkXFZmEiiCQKwg7VTJifaIJRmtSVgZxp1p2fcmBaIAfTFYRyUdZ0rrnV+FAPrBb+N5lm
T8iYkRDFhxOgzjvRnkr5I4uIH97S2JTdkAQ0x6Ha1mxXgGWS+OmZf5lIFivGOk8CvmjovHwsF/zb
BJadnaPNlzdD/uoGsAoYWsk9JDmVzBwRCrL1Z0kKowCMpymqNNxjay8u1VPUPHPlu+JvjvUDVTN7
7xv4FL+mj17RIqwQtHbFIT8p6JQg3Fc9dhIiWUW3Pf8puBgeQZv5rDnRC90u3MbkY3814p2McBmF
n5XpocQ+kcdllNV33R4IBvtPD/roKXN2odnUNaPs/u6twXOiwCpV9TKolIF4O7aapDT6Q+pK7Tna
dpowx4JiyE44mxBtVBJRhawS88td+2TDm9d82ay2lCiUzN0i1yRV3e3dArJ53H1VvM+KQjfv1lVs
4FTV35EGqej1dElfHSVLUQBRmhYYQ6MLX/XU0dhv2UwvpCYdhRLjaIjO6tebS6/xZ+JnvA3Kyzo+
8/tQ2TZf+aDDMHoH+uVzq73BfGH6jQeAHHpY5Y2cWDBUH7FfvmNle2m8lydJlpBQwehBz+JFKNbl
zQLmeaRNJJcsUm4gUAOUwKeCKiXZ8cCMlAUNcAPAZPIjTe0BwVFrpSDKp9S/+eKNWgAt8l9pe/U+
zeVY+mLqQqGgX8ZFX0fknoKgkrnNv1vKx1iLd1YWva6hJvZt7i3mZJi5AlZSN6ySVTyITJvjCMl7
0WVHf8k4GfDlm+ogzvQytX8hsqHqWg31FsdTULzcTuXWrSDqENl3YZkGGKIwlXxeqeCLXUbh0KT8
XtNgBekhNZkSHQquOhxhxnpLfTeRjtuP1d+Sn8QzsesRw7DjDjinr0HQzcf4JWlck0B0LvPYBw9X
UPQPBswWQmnycOIrvQap1dR43IoDPE7NuqCItUbpZUaV4SURYb3q19e4FOIccVlI6k5YqvMvYl5k
o/Rj4rcqeL4Mqwny2BHFqfQJX6XZC1thy9ufCR3Ou06TGeRi/ibAmZWznBHDJZ+lJeSdFutAO3lG
v//8WX3zkF0ySYQfYCFFnp/AGQOQbvAzCvAEKC6zM4+qJMQ3HTlSgb9j1QAAVMQ8h4FAqlFbfNO9
g9r+Q9VMu2I87mwBZKe+wWh4ziddqQ4JFMqmgPO7rTRChlDpJN0W9Str5wCAATq3VBDOhqN0bUMK
SoosLdZyWR7NJVATEMSidNOELqLZWSpV9845CiUWVkFvh2/SAgIL1f/udynVegU0fRpYAmvBblBl
J3rj4E7HZYRtRLvxynObfEBd9t6FBoLdu9/iUbdNAwMVo7y23pUyf2TwCupGRKM+Ms33kdIif41b
DMB0LFhdMRmnbPFJsQfYoKt7at1VVC6lOWfostWEXhitkwj5WrXv+Bcei73rImoP/lqUmPsHL9CD
GMDE7V/ENCbIfXrWkF/O1vfh5icQsuk8FzJvLaYcJccsQiVqkgO2kVpj4glOcmrfEQ4aLTMP3QX7
4RtbEtRbfa6umFMzcfUOTVfhjCyBJ5msAbzUcJaTRDQfY7LXo0akhweQyDRXEi1U/7x9WPhqTbQx
iCLtkPxmZfFPZ/DOR/xYRaIsM+cJ9HbZvLIXDL3ZCQYHxGx90mQNo7CR7mPjP/oB4UG9gZxHNDl3
x8bn46lt5wSjTS9XlA0hwPIzEqoYwe2oEs7bkya40fKIsHy7WLm8V8zYtVSWiHLnzPSIcvpi8pdB
0UsTuaFAE9uRrwzOvVQSpu9vO4WulRTiztb48YxqV16CqnYhocrw8PHn5nFqTAUT/xKPLLMiXUH8
G93/KL7gA7usiHZv3wAhFoXhSLtA9aJdot33IcO9RNzonrEajqprGIh+Hp5QFMn5WxxaTgoJLG74
RW/xvjH1eCrsRFafuLaE4SnhytmkmB1LKMlslpgb2YyHp2dIYOrFZrTLSDeplwl7WPD+LIr3Hey1
IZx8UjHs2J1b4HJfouNILT6rcoEBLm+yOFbE3F8mbOk+RfMrr7XdDJ1U93yJVpUR8jluAgEFj7i6
gBoWmVj1TEiAzaAVqfW/3KIEi2KqqS09tSsTbjP9SLLg2OAEPBBoJ/6KjaohsdQ1BZZyumaiq4Ss
MwuxLYxPivDPRh8WkMHt0NQwaczU4fWUsbC7GcZYnBoPmjenyoWkAvanmf8vdfDL4WuSre2FzAAZ
Oi/K/gOnXdO89gCW1bCwat0pIVQpZu+t7QE2DZKyAy/0D4DZk7E0douzVc2uDSg/8Eynlvz9WwwQ
ZFr7W0LOnA9XUKtyTmjpLqqAFAnSDSyCVg22sUWvBJ+EJzCvuKjyOZkAtnFfMGirl1lYOxZcbqWE
xdSXuxM+FVYEKHKJzdMqgwEVPHptQOGaqvXPOnfJQpuEw/ESQ5kkQHdP/7Rl9e/WM9s0GFTkR/cl
Vzh8iXVULOak3UB64who+a4mo0ko+GGA1Fiy31JQA1MW6eTUcERHebbi9Fqh/dH/8VRAGensWXM2
wbP741lg7I8NegQ20gxGywAhopfe0ZP/b2B83mw65CEBcNJGlZxxEAIyBrXKWywZkSkCmrMpOW9M
P7zzvZjk4Ck6XMa8ZLGmhMoGcOgVxjm/G/T8FBMy6Md8FVeQLBkeDOhK+t+oAjBKvjzbJV1kOMPX
Z0MTftHbirma8Dw175K9f6SuTt5BjN2NwQU1BFD1wbzO50ODAh3dApTrhNTIlcTcRHBno/bnTgKm
dGgITEwW2JpQVE50JScEOKaZavuVT6DWyJwURnsvZVal5G+GFyiYzc9HG7IpX3VkWr+JHut+J2D2
KNtqcJyhXgGF1azb7+NZ9usdXMY/M+wabEUhsAQgLSZ7HG0ZwEqnf8KPjnHBN8e02myPjjv/TLF3
2m/d8Qo/fqpSBXjZzxdaxbAja3Xf8OzYSiKTJE0GMJVnLvzWieUfOlOU5vIipaDTLSXSWteyUxIc
F1NnPA1opM7+FqGNfbYuRBI1y8Lckl3xUiL9VgHCvY9sNAJ5znKURt0SSdLxWQGUU5MO85VlXeoH
hl3pVVWHT09aUt4TPLpfnI5KrQpNZMDQkguIhp7R288/anqSLyAuGtty/K4xKxZXY3nAK9C9+y+a
bCHol9TkfwtssBl5w7hnqSAkq/baMdLlaetOqn84feLa6UT+U/o5Vdv8JRfgdJnXM2SSu0HOELQS
zG1V+bNj9t9v9i4bw4jn3c61sq5O7ItTDtoJX/kIopy2SB7Isr2OgeUm7bGRTNsRYTxU6o912luf
UXWsoNRsexzh5EC32YmBJVAQYXhj7JjrymKch9w73okjpaI8IBMfmyeiNR4sYuSBXjpjKuB8aRED
A3NucgKcAs+G/To/5CEhowFBe+LWfw5ObnDOuUx4qH5LDN9OY9X30/Lx6/irixbKkqlAEecmHo55
YfUgCPzWLDyCSjWWqpZEDOnD/C2td5mebrbW5K2JToTraZGRx9QZiaQgvexdCyNs2S67d+PZruYg
JwHosYSPPsoGm1kT//XMhBWvX8r5PnVTd17qK+mthYbJ71DgTKwd8fujYxNpxQPfTy7AsQ6A9pUa
s+mCO/xlITVgP/SJ+h5QVY4JInowfcJcZHq2DCKZsHLI10xefI5URPbXgQnSw1ISVcUdqVbNi/tH
acxQABFDpCAyNCGJV9flLstOMWvvk8+pXXrauY9mbJP995UGA7czOZ5tHMLwMTzl980Of6wyB2dI
hOb7WzrazLS6VLqEn+u8e5XCNmIY0ErZiHoztPbXQ9zZHKXmeaDWcKEt3Pqc+bPY2lgeJdlwJZQ9
csrj6K81j9F9EHE9fprBFih7ZTfnli7mNtDEdqXiBTJ/uigeKEcY5V1cfOo4isNessjnqbXhyawG
LoCwGJcSjF2Lv6qQD4mohNyvz0onK8n+dZPETdZdYXBdJ1/Oz3kSJZ0QwG/LLAGDxW8InEmPkK+j
oqIajfZT4wGXRwm/odVbaZUSaxAwmRgR8+eSq+dBy2UEZQcjoRHej8RISFKiKQ3WjXSqzJDsiaLq
Io9OCmidl4BcPUZXQ76b01BlXbn20QJt3+Ugd89Mg2mpAYGnGrqMmpktik3oa58pthjfoBowKxh8
pBB4NU//mnxp7w+3+yhBIqgO/E88o1EtuVqE25SKaEGhUxDqmh8pMbfmulIpXtBVcfrFlcz5a0Nh
e1gyLvc5/ITRKnDSBJHhHLFG1WfigJJwSDMZMJZ8Yfr/48JyFFELPF7H/64l7akRHrYCDiKoZOgO
htTR1ZW7sOr+SZTR6A6sXdLs8omG3Vy8FmCMcV5Gb/cNpG8vhUUU7RKzLVz17a1kHUj/Ooum+2Pq
fwnVfn31bC61k0Gq9+Kw7bWO7+mU6QzKKwLSh+0+H7+LwmBmMf2dOL6lRjTUxdxWrRs6eQwqW0w6
m8GFfxy+vdxHAAy13FQz2I3LYl6MWxEf7HZ0pmskKiM985bBYmEDrBmI6FHL4OrG9tXN/MbUdOLF
+0IX5RijuCxRsnkWjWP3C3ScQNhh9cH4VUL6a3uGb5lfI5cHclFlACYQeN9AQrTIg2pWSPhn1O8T
u8p+nK9hV7hannLhy53dy8jzpxbhmJ+8Bsr18FLFIh0dThPKgQ5b5OjydpeYHD0CjJvDez+6jr6u
hJHoIEfMxzwpm1G+UOE1L3JJjVRdoTkAeIsl9ex4ErfuN7Dn5Dw9MFeelTBefuLfa3kMO7Jnv/K+
5xqPSW0l1xdUuv3klWxUbbWxY62t0r7K1cS6p/eMp31mSPqFAU/wpAjq/zg/X8TbqC8wqtHWmKZW
HHrlSQtTrngavbnbf0DWWbGmxgx1aiYaf5kyCa7j2Avx4YbTrUhhVs7OAWibAR3i+rlWOEh6BqQK
9spt+aECLMPeY6rMuA6J3MTpcbs3WI+7vsFioYGL13U51VDYK2gEP7w5u92Qv0tNPcqshKeiuqlk
oTDj7v1Ck3r9ECxMGY1ZSn7f6MLDSCahENjg0PCisRjt3P93g1REv5aZf6GFySqt66m3E0dIhPAf
MF2bSxVF45ie3muxzjOYVAYYaoBGdcLxw8uM3OhuwfWt4WS37i1ZQgp3UGb9AK2+2kHgMbzQ7WAJ
3uzYL0cbcE/val1hEy/Kgfc17etbD9lQvUMzXvLLv6RGKyYk7Q2t6aZQag8LXO1jU+vzu80aIhj3
1NVcGjXnsueUC8Ga8rWc7jkMfRk4FebLwVL19qrpu4l1iCkM0fXJ3SbYyl7q3S3Hvw87/rCjgYVo
RpSTi8LMdAX8KOg4rWKD/P/5pO6PdS6FTk64bxRRutmqNbFF3aWQJ0U4tpjnfLstin9HH+ymDyjJ
yRI5Fk8dkzuHFoIftH1tIYMEjuG2zQMGdQz31cYpyxDhdEmPiR/fywV++eRFjzcjCPDxge12PgSP
PZ2+AGlAXpYoF4SUqMRMdqtxxNwdc8BIt4ZDlQR4HIpFuogMgxu1V97ARqJ7SwXwoDy+L9WFSpsq
2UaiQa4IPfKiTzEOPi8Z/Y78tcKaAksnhlNyvR8y55I3cQHfLelEVSGhUldX+GX6VxOszmimsRTZ
Li1VbNSYh0rBwSl+tey/KJ71xhWRiMhufeFunKFMiaG4VUEcY6A66B6U9LO7h7AclNJ7LSz4X2l2
Y9CdpLLTOMRNBz3WmzAqGlQKxXWZTeGQTVG17c2aAmG8C4aXYzxDlOAoNroKWaun1i2CBNyQFhC9
XJOe5mzHs8+46MNEplQ4x2z7f5HFmTh0N7XUPw/4pJSbeoXVaghzzIYo1G/w9xykgucjPsvBF2lE
BNNjtAQoJWJIo1m5HimmVDOhQYIGIr5zgIzsiJfuCm2r9lnXe5Nw2xsdGhbRXVOGDQWWI/0Rj5ov
ygeyyG7SbuOYI2oaVPUK3CQvraNxVFliDwBCsD8/Bf/g3Cl1LBXaia7+2ZxhAQQ4qqswxBrHrPFg
4kYAtRFxSTRBvPADukXz4nQ0AV/UcM96YfZYQZQwjdYj7u5GPeobxoPgER/8n0s+saGF7x76SvEn
wmomjwqag3iCPi/cNk1YEA3IjFZOHV6Ox4pAVexCawSKKF9DJTneas8h2Kx+Mr/PO72M8aPCkF77
4YY2/ayFLVNvpSalbZPsNx2NeMwift9IXg1ReCKJHzAzI4HtHF16du/cVkjbqVwfIrAt4+3bOAWX
vRFHou7XbVN8i7bdAGQHlCExj2cTzl3ZD42Z1VDPfH3SqoYbsyRx+Dl+LaIxW03sqvIU9Nlr7l8C
OEeqz8QDn5hKhRb3ky02E4vICnO+ZtSJIDi8T316+tWLl4vr57o9zeOotvBVG5Yu5NUWgQNC547E
MHthSsfy08T7nXquhp4QEp9J3OmtyZzA8dDZ5OeUU47P6GheGJKDK9YlkpbeHbt5HjY1zYU4hTbf
FJ77mIRd7ZgzyBxXBWvg8PL624MX5LQ6mEW4c7dp7qp99bS0wa/EfxCU4+62lx9sIwrZglh/UZN5
PvZrSvcWA9oIzkpA3Aomih9o19O3eNARHuFJgjWdaNLoLeY1xjN/yf9/5rEqK74oM8F39+lk/pwG
+unZLCLa30TMsMO8spIdAnVhpqNlniNjsXQGjRfqBVAq9AK8UVduMInp/lKVVpQf1cysysHwme2+
KrL0hvUcUqOl5CpToR1iapD1MwGJDri7ZlFph0wTNMyNKBrrVYK0u2dWSWvbiyJOb8T2mI6gKJTT
glCQpzviqpXKKlRgeNOocodofGWSmQeSZc274T8cYFhSA/TySnVsA1J+qOxiQQQ0WVfxWH78JUdf
beIHHZ5WXGeKcC17TZOnw6ZGxBPhiB5qrmM2mCz6s56RX1GuF33bDStsRHK0AO9gf1BuGPxGfNTb
yMCSsleU+OiU44pHS385W7gIFt7xDqvuKh8ZqlLpJpRmD18ikL89d1+WFien4ORrUHJHKa3D+B/T
sUwBfi205arjjatJj+ILnh5q3dc+sMkCnfIGW8DXsHkeFFjb9/4k/f7hdkNar/o+2jSqWeE075Oi
5PC+SjJziECbLyc1gB52TJ2EBbYlpQTpXzdVSv/YAHdaJeb8Nzl3RteIwaJ6MZ9PIbA46he8kl7A
HGQYpoWGWQ+t8dQmeT9NnSus+XIhesYJbnweyC9AaAZ2gRPpVCBCpebWkKW+YQ7pI1O86DQxscyk
RqPMGsZ+E5MLo7qUQ2Pwc27+34Ayfx7tQXKkgbeQqp0eE8PfXf3mWGkB+YpH91i2ZnsR78vGd4hf
ATerPsY4Hh3rJ3d+OSWQIs1qq/rTexWK0Uvi7H1bo5oaEoK3ALPywmKIejCUpxoAEmXvv0A21kcY
m2hZTXJr8RAjqg3ARLXSL86YTbKv8rTjyUhgXnkapQMTTaRZ9t+Y9Sm/amciRjV2UKyLyQQjexWG
pi1aLB+KFzrh6Y1xGI6dznmUzzeh+ebVJxBgjV3L2pRWYWsIbKIAHNoms7t6rgA+F6gGMnJXNMVK
e5/9KjhzBV2oGneTQgM+8KQeXmB94SwK4F8YgO83UOhlxckUzt/cpN3dXh7iGpEeVNov2umrJnK4
atMFxPwMEYlymnNnu7W7FVJbAX3fZXS/IMI/pB+QF6hGmqW5odLv16ilIoGy8mctNlDpdauFFfqj
BnhKZfakTQjkqwwfiBhKjojXR7VA6Z7x6R8zV2OyfeyrFEbpqczJpyuZoaJCgYxIFowS+NSZwpGH
HobT5+wmOx0cSLFe44aYIff6duQtizh89z3O593q8Xn7++JgK8AsqyznFy1WvTMUePGxhv3lXRmw
bRdfgVE1QOeRdHUUORs3+D7KRP/U8Dw4FCY0prah0QYJKkEAwNzdQVs6oMVMEoj3cU/jalwzqNda
k0osP9GiG1WZHkwb1hD9zZF6Px8p5sB0WH9ioXdynovVtCn+cTUq8YinqRR08AkXWP56S2qasZNW
CeDEFEhRW3cNByiPFMuY/OoS1ACa66iOF2nZyI3lIH1GrHHrldRuHqOk7TMof9HuopxeGwEtlQL0
7/cvoBOvP2y9Z7AVHdjw9Pz4eKiPpGkXKoKkTHSQIRWe9bIG4MucTic+PIfplaeyYErqsbOhkuRM
5OHEgyMDF7vx2RKYkTEExW+Aim2HV0bMjsgtGBI4F2ZkXLusW/N51mv56XuaHuih3HUENjAwfr63
htCX3xPxyPbwn03pIH/ZfFMi5p75KRwWVYrgPe+7GWvOkHw5EDTScBLakLyv1f3h566aXI7I0wFj
kZENTKHASl28AwFDas4yQDl60EuZhHRb4p4z1fZZq9ystIWmOOoZIPyDVDGMOxH4tITgebg1H3tP
w7PduzCwwJuxS04DYGUeok6JeYhUSzrYZq5TV9e8jbY0fr2hibRKqimyBXPGrRVtektgFIeSv0YP
iNC38DwNFrGURvNaeb15APIErw9/2yylNF6HVIg2E7mS9QP3ph2IgksGyeIpAhs+GkwQB1ORenym
PDaYGrwS2c73TnqsxyadwIkScej7INl/Xofl5wmQ8eEp2R563Q5vZJAbJCIX105yZzH2EEpeCCBC
anAiyVZyd10+4pAFqGC2DZMoQ2TVJvAnYbuD634OQFV5hCBR44az0+isCcr75MzEf3WRdqW5nQ3Z
5Y/w3QhOmapKsa9MTVsppAVLs8ZGrpP1W+0a8t5kV0slmCy/4gWT7XwFosdmJQrynl91PnZbB9Fl
cQ1Rf2RG0dyafmTasUYH3aR+1oCw/N3AYsODQbtTkCfYr9RBwX2hfs3p663/ZvsPfxuEDqGHhAdF
ES5mLTsn+rFcAIXM+EQ9Q3no50MzxRXe4GlJNCMr7dKGG21FLzO3Y1Z50IicdVZX/dO7+hg9KKHI
5q1Yk3w1njgakDGTKVXfSywdjNw5URtewaHzLzGF0zIpLNwj6NWS6Bv20DRMcGPOM8Y/
`protect end_protected

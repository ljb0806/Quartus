-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WM3PSV07C2P17Ib42/OT8Q1j5BCIyHEl9HcRu50+I0NZOz1AEfPlT3sFnowk8vV6UWBt783N9QlZ
k4mjk8leLmYAwYxMyKErzGJg2F6ZLcHl0kC32TlLMRA9EZk0mIZkrw32qcWzG0QU+UDEVOfqP6Ja
GTE2ssF1mnkbkjRYxGgdShkyF0RTGEDMZMLV6FjUojfzQV65vzH/gOUiwAPfEzq4tKgNFcpsSNOB
SXZEYDNNv2hHUXoGdtZcNc04XprdsD3KGD6Ls6Smwa7AjO/+th18SpTS1Vo4FFyKZjxHy0DLZftV
pvCQ1GYJ+afbnARU9GXsHVg9GZGX9/6WtXTHyg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9728)
`protect data_block
4Cvm5ykyOJQjE4JnrckubY3cODYahInj0vOOVzfIoy6Zpxye9idcaGZbOoQAJdmUXN6+CvVVLrAJ
CYsgp9FDgqSVFDM97UnlY1c8E3z+sx8L38yWarBlrYUEMG4Edqqxrx/pWzZQ3aiXkUlFygNx6UQY
Wl4oXGyBrC9RrhY9GSQLQjY9CS5BbqmDO9WxnzptxtrDMUat9TgGqOeGzaMcr+lxDEH5OiCL/o5w
PKwApaI/1NkDcwQCtOfZ2tVBPeD79WrxeYfYTZ3+qqWZuFt7IJqhG4kWr6h/y0BT7XLMy+7gUbKO
zX2hlqXnD8f0xeFohDhouYG03FDTZ1v8WPeN7md2Ed/fUUJ5xqce9SbRlzGJIn1UtixusPwSqlzp
2L91EDSTBjBqvLlwLn/YDIDFriFrlFmDy9lN8t6eotcx4XReWdNZa0awf2ynV5XTprQIXmAeZVh9
rnSie6FpfOXhPLkTpn6RA2m14XMSXn+/kUUVgYHLE/+dlbXLcD3Lq8SDjV+j0+amSM/07pUvp2Y9
PzbJy1fTD1w3Gg2U2Rl0Q5DlqfX9wuwnYju56Jysw2W1s799TyGDCL9HEMcblASXL/dvND6EAX4w
XqLH1Ew3gcnX7z4vmnBeDS3cDvApqvEH9FqjkdVUulosU7YsDuhf9AruQ976kX+Y7iA+wAPnMj53
2OAyIn9wfZGV9A8XW3L3DZYveD4id6pSgGbL8gKpk23sxhECeV6s4SBBOTE0vH5KFZdACu6+xAtx
/trNcxJNvYvYfu6YWGyX26WwZFFtiMLiHVKU1pduLgr52p2lFdWhAPCah0r1+hd+bj2d7kuBg9dD
Q8E29WEg7SLqnmlareJlvmO+3CnAnW9QfBPGdettVB7jraYqQVbZDVlh9YLBxcLGqk4M2U4xHlUw
SByLHXM23Rp++JI0oyz9mOCdFbFn+9aEh0lHcuSUTx0TpPQOrZk3Txl9poZQBteem7vm2K/+wV1n
i1qoHWfuUi2Gw25jjCbmibBT94oho11SluFdgW695qzAGcAVGdjbgInAYcZgHHw3bdtkUyucnCCJ
y2qfn+BjHBmXssX5jctc52e7eNlrWcl/uOCg/y99iqJH0nkcV6kgmHNI1bsOEHgdiketsBoPVoNC
9/2PbHqSHkcHhqgUMxJERlCJxZxGrTpyCEhcpqQznN9cKqbf71dRsKEikhdXnc4pfX5XPguHLZCC
xq1QhzUtdsx7ACQrCIKfGoR0gMh6w4i0LCn1AnOeIuxWu1u970ZPj4hqlSa40o7+WWUr2LhWLPT3
fowtkoCmylAv/C95lmHT7JI2fpPN9A4hFB7ISE/sew7cx3bJloa2B6dV3aFJoGlS1+NV36wdavx+
PH8eug/CDiGVdrblNyABFJDhsb9qZoo0z3hFKItZNQyY8LxCr/7opYLbPRb2a9zv5yhqNbtcq143
m5QoYzQaUahQK/WnmAnqOraJ79n4GHJQ7p6wcj3zGMhdbxJtuE9WtvP9kj56kDA6LvW0ki0HPS7M
gUHXwLIHXHj0oZg7iN0HcvKtl8aJGupBib4S6Ghl/oCZ49vtS8MxJpOAN+fkUBgZ1+M9g7UD4Qlf
al8Qu1hmp2qXaGnvEvBOllHFOY1JxulpB4YAg1aqzfLyxDRQrN1mzxYoy8ZwLvw43EXWEyyxQfWy
wyEIQf3eqaozZ5HHOTHzaXXxOCrdkCeCA54JUGCkAiVYYT2ZGc9uVrl+v2IyvazukGIlGRLLYVJW
BNl1LVQB+ReAE1CJEZn5hAUrVx2cc8RlFRjCufCGxu4wmIfr/NShP6imoRJk39zWAonId1A10vpd
DR/jEuDLX4KFs9dDXWD30JtBcLIIy125hMCwe852IfP1c2gKr/+zDE2sHZxaAedVewxDmYV8YQ9g
8wtUbGqfDEUct59IevV3WjpO6IQXLua4EV26DSiN58VCPsesq8+OUsmmcr/xwjFgdysZwi5a6DDe
BG3DMYe67T1GWJLf4F0tXp1TVgpL+YvAAQygvPG6KEdPi3iKXHLQ8CVrYqq7mn8IGl3tfK5pIG3n
c6mo/rywx9DV2vlMic8EHVuPyjghy3qqIoxf1ULVytRifuEAsvvao+dEc9Nc22moeUY9i+wQYLy7
SqYZIvQqtQWeZPAh8ERn3gag+VmJVIfA3KdeJhhNefb2qBONsLldXBFI7ldQoGxyK2prQnxfDYWo
hbkdMyKs7v1WG7StAlwVhoP0UZMbPpXxM3uYH+7p+hZfUCeAUewhB1+xEePUFe0VyS2wZBoXQDJT
ybEpdktqLbHkMWeVUOtGN3Mq34h6U26QvOLc9XvgEL4USmwueNSZwiXdJIl8ka6IqxGLnJzCHF84
rjAqtCjR9e9C2UeYZ0zkiJPaYn2EtOh8I+srPMVqvZRNsqki0HZcp4gjVEyFZe1SeUTIrFpWqwp8
0VJfwmZAeZAObNdC9JkTL0hzONjpnlS4+7g4AGnwCto6QgjPVeik7GDqE82OtDXn76ROIBt6Xhzw
S2fxh7TbaXYZ/MXadcB4Kg1GmLndlE9KEqwVqvEI5qRxtC9DzlRnF+J9R1r5nH6FfxJIqG+qeFdM
AinhhNiVWbve1XUXNtARFRmOVNTTMH0F6dDPvayGeEykTeHKjraruf1siOl66X5xviUeXwUQNBkt
GfrGRpq1SzduL9dY9K3+COC7aLFZJ/pmUOo3EckiH5T3MSwG+OQynu4mGkddciTXvaXt7EUm4Bie
QKhFvztDyq7BcbpC1ND1jESElVnAtrFaVupO92CClCAfw5sBSlN2eSgMoMrFNFMWJ2BEH0edDI5b
G74OMJwh1/1pEQpfSGWaJ7EC6CB9FPECzaiVr0miTyR8cniyLxyO/rM9jrDRAQvn4mL08rWdKc8u
Ecp58P91cn+4niqJe3uNKb+u4JDNCUHI9lxGJysUAQ1YbQDN94kaZ8wj+50sC9LzCr7Pkidz3e93
UfsDV/W7c8iLCq9si016NgYjd7vz6T0BgAufGTYCmCmPQpWYvS8//ja30jQ895GmkECKYyb96R7e
j0FxHJYwrSxqmNY52XMHP9xv60JIv68LsUCjFAGyNCQiQOt44c6YJjvdDRn8hHM7nnqiJjSJibag
buJd/iL1JNtNIOOcElomg0gW0Z6YMfB7mpHaJPHsz97pbmlh6lx6GMQXvbXKDWGC8e1dEO2SJwkR
ZaHtilGz6qwZXRFJ6rHbOjQA7rtAL/l4VM3aQDhktpfY1WLRTFcYcgpwGW4pUznYLML5We66kTGK
Q/b4+ofBbCizWbzjTGjlkbrBtS7FVhve4aDpM7Sg5ju1IOBq681WEEZG5B21LMSGXKYv8tlAkjPf
bKKEEVB5U8fli8rvljkyujqzzJAJZoVWChhNLIEFEJciNw2zr4Dd3D7JID0Q6tGRWmLzcKDIFNIf
/5vZ9Iea2XlyUeBzOEqKjihDtCKpCpmgiN+EDRLo6wsAYyV52WZzVlypDCIslpiZMglkI6RFdQ3A
oAxWPLS5J8JPP4cJ584g81PykD5o8JBLov9NvIg030hgQxrPFYOc3tyQI7sj22aZgpn35O81NTip
a9j4y7MD9P5bM9arxk5EJdpQ+LCh/uZl3RgoOxDECN4Y3sEckt/DSYHcKpowGNmKkiDXcQxzCFyn
bHR/ngcDM5juzhu9qUD2DzzndnezmCIdO2rAtMinZKc5w438LU1ieJ9qM2evPAT7ELR9fLvW04zu
JfE4JIe6QZz8wX3aA+/Kbwg8vi1A9zlEJP741cqUC0Te+UhJLG+eLVDvz0nHTrOO7mITcSNFRnGZ
1NSZ5t8w6+zCH4ur5L9AdKw4771CjPJjgJHHJCT3Umkdc7zmdxflFkJttMlYvzHALZ3mw52vKzmd
5RArbmtE6ROTBQNSBb3jDmZt4piOnuBWyIkPT4rN82cmo8GBSMFUT9b8FKldN0Rc/pFIPWojJcIC
b6sWdKV72nfYZ7Ahf3511yI3hcgsDs1eAZKfRfK12IvE8x2fB6XJDqTFDslyA4XXSULnKCmqLdZ+
EjFm1SvBNPuDl2/AJWCsVzpnCibYKqUrZo8eO/iu/ksFvnrV+CWyqAvwyYPS0JQTaWi39G7ADujA
Jdgr3mV6/sFbtPib/bWVH5NWZtzQMCnVVPz+eaPi00hLW/g0MNYZkl+CrQsgfPy2BKMVFL0vxw4Y
K2cDkss0G1gUQDn6xmotdNzQyx9repEJHJcptscyMbS+fSZ/Cb6hSFbxyPUrdWb4ygYUQcfSXbp/
NJbHemz4/KiPD/KVZaMPlacCoP1ckDcSnEv2GZYIU5dkxxCJ/UON2/oKrdAF82PGWbT3lqsJrCVn
FeBFGM9AlDLbnoAUE+zxaak8ENiD7k+ShPy+GCDBbjT8CXWYiYyX5RlOeayj0nirnAKFpgbmECgc
EUlU8AytJixzMF/Hh1MknWz51FQDnyLrJaIS5Sl2BJ7e+GxYgJUP4a0wOfs1YsulpVJb4qyqTolB
YNIQjv5hRnPZMtI8W1jW18s2JkO5GZYTW5qkEwZJC4JUwZjF5IBN7obK1hxxTbgeFh9koJUOouhq
NSGYnlahdBg/GmM/DupFtWas1syDNTFD36jvLc16cgqCR/C7qe1gngEhOxojb2QJ7k8tTcb+XDOt
jW8yuRcyp4tfvoDLk9t5JpWiJ8eyLTj3t4fL/njK2siAuv+JuSnoKF6N2MgSEBLqV4YnWkl6EO3u
Z07fUihokOXWTMSNGuEcNZiTtfa9hSBeOLaqSPMYFNp6N9ttdQt7w0YEgm7WzDbFbWu05vQeHnXu
ABP9zK2yWMorZXeP4IZSvRVgMhIoco2C4pxl5vM+eQlq5pEInV93rgvApiRfFYmjslGvLcu1TV2W
+LTuyhW338WUHc+I0yeKyxuHWpyhvskcYP0oFd0taw24+fnhFqW0aD5QtMcneJ9UJ7ctjzt3VNMQ
vBa9Iw8//p3AAcsWzVXGYG3HrQpwDEDIm+ARcb3ggONPndhMRTZBSQvx60cHm08mldVJb878Ghh/
xGEqenVN694O9nYIxLTNNDPiZs05Ec10YJjiG9aMtnK272/OOYIV2nAByi0PfGgZY/yhP2RzBitj
sUqy2thma8k8K16OiNTnPRJmdjueSDw/b21ijN1OywAG5auKjcvECs1VQBz5OXe8Md5L9nccS94h
VQNmyQb+gbnuzExypBx6QBSX7sRqKCRwnuTFNdZAySGjTDMM+8Tt95VwtvJj1mEYV3WU/70i0BnW
spKRmyyHsXnPRc6ZeYOqp9OZhqXtayXGs2GWye8B/U9HDpoAZht2lQPkedOtjahJg37Q3M3t+S8U
SD4hNNBIRXOrtgJ7njkqofrZxWsfI8PKbXgkk6vNAZIjSSifsHYRe5QDPOGEuu2rjzsfEoZSg5yC
4YxfP1eyZJ7cXG3um0cEg4/+JxiI+aWXdHjXohemiBrmpVzZI2ef6Nl+X3m7KX6wOZxs6JEXZlv1
9gR/DTpmypTJhKqIUTeMvlJTPPHWD7Z3K0Y3XGK1FY1SJ2gjN05xB5cnnbgS61lpe6IOr2+uGhAB
Qf6QXPNrvprXYZ3KhR+6qeLzBuBQnfVE4z5z2HlYfh/r7iavEnSIybDitQ1Le54X/ROr6rm65Ih+
uPh137S4U2/mZ8Ax5SagGKbArzD1MZm3nDYgg6ul4PXDqTmlynmD0NypT73zthuGBl2XbY1FwVMG
o0LoTtnOJWwZWeKepb+TdkBKtPto4hDFeoZyHaIenKvF7N6Rf1mP2fHsIoyx3sG4zkLSUmE6koNO
jroScjPggSRYZK7s0C7JicEicpTK4XkE4LMw9OoEN/Z8ytMxqlvNVFwJqCj7pRpMyai+r2KxZI6o
xKI5Rk3jRA1lzt1cOiQkwJcfo+U5t29y1s4YgbYoW37HhTJbK6tmHNxBLf7VTWgX7LBxCNt62OS8
D9zjPdvcpNL9dajXhO7KtHnTXAdq2oQBnAjljFxiTu/oLA/O3ReokVxVWrqqdZhfYJKaiqy+YurB
UQvLwNskNdbfj1gMweGus1wOcNlrwTQ61HDfULEq8xM6fle6SNHPFfH0Su2NwOMSoga/wlSRkFjp
tCUBPrQ10uzvecqPkD9jPC9e/XeBYCV96RkTVu5yDXjTI3vFQTudeIPCJgJrnvm42r6t2ULoC55c
DqhMD8MzIpUnaKMSkoWeLIoAmE31IfhUktdNpUfOJWvw8MMcVrQLrb++96/MytBEJSo14HOrlzuY
UNW+imgvsJmt3e8XLClj41hqnOm4TjalZmZ8iGs9oPWndtCoCdgjlu8/+bSrzzfPZFEGff1b7IlR
oldHGyHuXFNORZOLbbSWQnA4kBE637RfIfB59J88PaLdoajM57MuI8mG/I0caG3rRJmvW/w43TQa
LuLAS9tHQB5Ywm3PMfe59qFVOKpvYmtjSFAMA7THxXzhSlqjMyYJ9WVLaPrmMlVjOMEPiQIWvZ6C
rAS6M2MVfhlCf8POhxkNXy18zvUQW6MAG0sgJfOjSte5XR5318xs6jcT56N1PUXTDj5Ab7IIfY2y
LtvXhKaoKBub6lkmowSusQvKRDLSegyq4sNM2vPnbIx/2RvV6REPTNRH1i+Ho/plcwGeFZeMYLzf
EgYuKvWux0s8Adrj7zNKIUVzdN6WIp1ckqJ6qSflJ9JvfgfJ+obKdiWVf9ytxovxiPq//WlJTBpy
0AxcHv/Nt2HNJ5gvMLhJu3XYcAphX0V7S4G+0tqLONs7lBJG2BTiSZUA/BP/XFsxVNeGTlLigM2y
Gdzm1JXuqpsKWQzbGoN1nndFzzy+OQFurrOtO6JbyKeeGq9XisU2eYnDtsM8zvoBhfQkGdaJZjXM
VXw4z8Op4x+YoYiZGkZ1oJMkoYHnUPSlqdociuRLgFvVzTtoC/2sVtsgeJmCN5brJ3VdFV5yA0xQ
GcjqYZ595RZoaAJUr1hlWQzk5KORwEzOtUARN3KJth3y+ZbqAKyT1fUe5YEBtcmT38DIiFQERIJE
YfJ93e1BpzUQ8gh97YqSIVUqJ4vDQq5xes+yibyisgT83KlBatZn40+dKfxdHxrPLUx/P3olOimY
GT5d3laM6L+w9UhSNaI8MXWg5GFLXMbfZffmqBqPCV8dWqADzqyZmoFFkOS7sFwGHRO0Im58Osf5
bBkAqaLz3qumPT83Mw2rlZYAOKKohAgRioFQdLjw5WK3hEGT2lngmxzwLpXIPYdjJGpDMdujJV+p
k68/sHNY8XkK/Pnw5Ad+IAQv1OpOIHOWBi+QTXS5k2AFc7RZk+tGTZPMq9tTgvyCLNcHkeN58Vaq
Gl4dW5aPv/aE4SWx4Ai7ijPcBPA4nClEik8Yy03O4tw7pzIU+2XxUmAMgfmNJRm1JPG/FoaIWTeu
74KuFELEfBs3SE4Sx0Wh7Kpu1Jr74d15wTrg5AdsR4oQhKQ19ipatnCqB+o7VZGVJO/fJP4ugxnU
EFpdQldhN7/t15eR4ze4uWAYVHOjAG90b0R6z3xZN77khNawxLofDnn7Oyy6zPMXtmfuWu9q+pQN
T8ssTR6acvARz+F+vTtI1A4yQSM0OZVsjPvFGBceVGeQHRlAgmy0AvB7OvzvwSrPiCuOdSuM/v6j
WcEC2B85mZ+2X1iuCkfWewt5VV+oezAeid6WHE8gtEFgUtE5x69sVgkUaIUdy9Xerysz3cH9uAR/
vPkXyazF2vZW9i+Ho3Xe7pDxxEfvF17E6pNmzbnj/Aums6/XouW6YXW5uRImYVNPnjhXJccpF24s
dHlIOHfLtFxaHpEp6oHyIZ+0TA9Ecq532lJ83IahrrVbwyRc1pseac89Yjfb+i7GlfGTlzIgaVES
8vf0a9AmzLDaLcXCU/TpwxDZgC4huXAaVVqEPEWYhoTh1ShUvBTIlLPM04TXxADBSQXpocyUVdzE
n0t5j2Vzl8zUsVR9ytenY8cAqanFSa47bklwTYhgFtNWUnYA+RA+AUkub9zwCg1PDluXps4Ptdyr
0CpJUc20AC87zomwdlhDsE+9BNb9qbuxjJga6wGkwhKsGHzfToVonaDlOW440TrAAhukL3wFrGOm
hyI5+Nz0FEcxC3oAg7y/uqWQ2Mznx7m0zm9kt/snDLZzxqHQVshcTMC5D5I93/xfyU3y5UzXiKHT
CWBKBFXuYmdRtP3yaeFJcXKlrbi2Yt4DN67K4pozBkpiPtudo87Hxs0ZDE6nq4Q7MOsVTJHqnklq
EEDn7FdXY1AduHEO61akH1/1jc7IqIoa6CTTXvgMX3cYuRTS4HczaS5Z25MgSmWDWXb0zEcED5l4
rb/izVTy8SfCjpCl/e/uTrTg5eL7v/I5Ec3E60SUGPT96Hx/iZqnhaLdwZfosmKq5S9XtHAzSNTA
CB8whN78Jhvg1NJt9D6WJGmhAPOeN4+WwOBqkZyQp0ihVifRcxPt3Or3hJ4+XvgH54804I4L/tnX
nyaqs62H7Rhlf2UC5jxDkli7w3w4NRGVfP3IqwdCB2b8gJ05WiLTYgBMbZcvO9EWiXZHrDmM6seT
KchOPIB+FWVniXpc70clzfnDNzvdOyotDKnG1a4p9DqEvVE4zx6C3w0uWdO6STfEpZKdoS9cn8o6
ykTLLt/A5LfZu5SRyi1DbwQ4QcEue/8E9ZINRsRT7Pv+E7SZC4Y0jLJEx75OdHAvJ/tgduB8Xb63
Y6nZdLzsmVCASL/piJz24m+qEYQMu2ud4DARl5NHdZzUAN6LVyX4PiujDdxOP6eA80BDALpQLxcC
5QVmkJwp+cj3H1hHah3U8c8/m6pEFua55CYoXqXurKz9wpjEVFtE/M6btSA/hVCQu1JFX6HFq3vv
UJILBg8iw6cHceF0WIckPf40tKqrmRfjw7uviDmm3XWWmL2U/5bcHPkGfcP63l2bD1Mrc5NZb0K7
4v2PJ2wVWABH9GwvQ7SsJmekSjYBl5ZLqKw9U7gUGgbapSX+AOcaeNcEYqzGRjxss3G406jtZOTq
rpD8unIgSixGkBfl8j195y083WVYOdmkkEG566IK7htAmrhIxOUNa0RnrKcW5etszy5y5ypmPhgn
mjEoIbYEwSp5D/z6qbgt9Rz6673piM6xYjBgDkEE0jiMMFgTWj1ftLukuzXMdfPF3ge4asKSKBbd
qlwzaJ/FFSA72EeEEMegrop/r0MBWyNJ7ytsocJsxChzpta4NI2dAwzcE/IDvPgRckOkFsQ+fuJ5
6/q0a8zePhddRUk+/Oi3Qu0pN1ch0XqHDUYYK49mJvMcFrlrIAvU+VMZG5kYM7c46wCvYBnEiphp
SclgVlK63byYxzPcNJ2MR8KwS2+/hzSkrMWrztVnTV9GYyhYbckqz6QP56//jkNKzbY6cOIgry1E
gcJjJedHlQ8NNk9c7YmG8x/LauYI46mUDSj0sgjo0ZGgcR0ChhT6bmJkb4JLKfQ/d0qimlWN03tJ
JKxzNWkGwrITkMkvJF8UzfJ6YOTnA7bJ2MPm43njtyxXuqATN9BJ/BpHwBAsY06mX9EPL9JttRmu
s0F0O5mGzFTCreJ6jDz37o3obm+wWELfjpz4keUqecQsrWe+IOvEAyZ9NuivCIyBsZv5n0w2IzUD
UCwggcRwCQ2M0CIyA2w9in42hN00nM4wt7uNGf45hVO6047wU5Idc5NYQeS6WV4dRnxrZz5XnbE+
KV2QD4XSgs1AMIfVByx+9ZSNSzczOKIGn3vTXl8vnVYG83sbYo4Rz6HmnaY7nKWqqeR1EAajQ0Ye
D6l4DBx5jAkLeTK221BPnZcA/LrnNf+CajmV0p1j6DLgpTOhzO8Ffx9qX3p0YbhkCCnpwuJ1Eyem
Q78qsJpcTXNYPgluniF6VaK+auRZFt/pbMs7UQZlH8VZH3VEqzhYk0k+Za7obKh6p9n7HuH9bxbP
1/gP5aJx62X7ye/k8ZDUwuvs6wGlQLQdd7KwJAV5i1xjLR5kA2g2Uu3tc5Dkr83udSeHb1dFoez+
6ptSvKTwKyItZWeV+2oTaVUAy88JMzgfhjaBvrGfxNP6eYDPtrGt2PyU2nDiQ4DzNN/8rG9OkF+L
OyZaGLU/QDMnBS7sCU0jzbKtHXQALpThiC45wOZC+hr6LnVXBZqAZtD+rYW7dO72b0k1Ea7DiSPg
+8O5TD5bGzsDfb5BB00trXKMPqpekALW+7Bih2Hxgycu/oDRtIzvSVIcfH/XNLZVf4u1y/ASuyBY
LBggm872ZJ1UX7Gj/kEVdepUOC1RjcimjTXVlVenHeKRWazmD2Qh20uXU4EgPsdOuFvDjho3O+9b
eMANfm82S8zTLTkRPg3vlVfoDddJVRNOoXC7g/mEvyXucOagOCYlQNpmKCnD6iK6HHslZPBuj2l4
d1U2gUtcgNczawDtCxuBqhPDJDBdWrI23siUApuSNUkrCkvCyendetvUmvVsqGaRlI/Q5vF2HlRI
m2DN2GhSC9+eBGDT6QJEbj05rxK0uVFUUOFC9lt2jpDx2tSsBUuyOLfBeEZShJQDTK5sqIsUt9sG
Tk61dPDbKlWQIN+j9X8HGmV2Asp38OxTQOeeLFPi1YbkDPq19TBg797DJwnie2RktSyDbD5Gimbr
6QnoMe/qITYdCYKo9a9YxNxmBm3jzPywZN+2tduNLKzmr3dvvFTnGAoSsxv3Eeb474ElucQvaf1/
kZ+KwqwujRbeA4Yko+0R0BGeb7rBVHlteRVxsoRbksqPN53AN4Y6gBdu5LLEIPy0JZUMfng3O2zA
xef6Jvz9CLqdlBx/dClOVEn7I0D4N2iVTdb3qpfAfnU1+TSJ8rjRzAPvI5lalWwCLEdp+kkwYeKl
Axso+RSFoHgacjgX5blqURzUxVsfG2KTIzlV+Eyy7DJ6+JV1s4rsHSp5am6g+wL3h/uz3gUa8oeI
PQbihLucp2eU+gTki4FBfd8fPJuTlGnY3zT+rgrgsuz/RCmGgmar57X7/sdtL5YPUdZUerUsGpK0
+Vntn82cG6/GppSzYoSZ96J0xm7fYNI5HcHcra41VEUXN9P+uB5FJlrYfqXoDb2VBPTf8tLlhIq2
htYJ83QTrjJiaEkRufiR8MwQqF4DbhVzpme8VfHd/kZiu1JutGZuvIWlijADWFfrzSrpYcC8OJKe
x+2IlKZozpBqgsLv4ECLw3APO4HkDAg+C1lkm6bqhTtxSFObK+C5dC5T+7KGZ6I4WVNXrqBwidVv
X5/Cib1igv6PNJOJbKAlOeCACXNoPt6lQBhJzSPMExtVcIUaedQCmCw/CcECFC51M/Gk+U+Pmo1r
l0w2Z9Z56zhuuB9hByns87N16hHzMS/R9dy+r2ajE6waxUdMojarYwgdUBS4Z8YBtlD6hWVAgsEZ
SfiAdWbIYN3vyDj818KJzufiCmofLn2CozEYdELR0qMLVS/JsOv2hRUlVEGXt1lfgrvnSds66KL6
k4h3gaIYKtCN/aO05VaLvR4PBnqu0nhSFN0flTWeGLgH/lHkUQcTZexdwJBBoGwxpGgzu6zxLEjC
ap77FGv+frMTswD7QWjqf7KRXzm073C5Ztf4ZovFgE1OFciSNmfbDDn2e/OnMTOnlkFcbvOx3XSQ
PBSyMTGUl0vGwPG8BlA/GzDzluTn9gIrgj7ZqlrInkV6vR/y4/ftw0S7Rn7zob5EF4TE0SaI7Xc+
d3CH+wziE3KLI1sB76V+FrlYjHg+c79YIc1dakcM6zqaJku/dI70Nya74qw86+eRqDPl0FvNLbMZ
cL4gnRE7ME0vK3MoTNGEZIeURjv+4sCo/xCD3CZiaEdsKLB0rFcihl15sxKiBTitBMsFI8S5U/7C
vw+DXKDETbXF7Av1T2xa/Y+jPPyIm3Msj5Lxxo01hHyKq7ayIc9S7QYDZXEv0MkdaRcSzmGW/nPc
Zlo3yWVTEowTs48NAgzgU2O6WEUXlLe4sIA+41YAnQzHjTrUjnethMdyUWvRtuReJWaFEtJ52i/9
cWtOHKSbXCkc5k4+vrxxh3iqw8YpfhiuLlu5zZeFxC3AFSrKHCatCarws375mxYIkLd0h8ydKyMf
Gyc49a1hgfXWPcgUckh1m2MRq06WnsRONDdzT/N70JPn5C+uGz/aYA80JOgS8MnYTUewHD4X6SQU
zXuP7kqSDn5L//hQ1vnEIhgodQw6B8fYtWRsVyRzwbV3CLRw5qNyeVZPexMhe4KDvsp0pbIJj6sT
rpLe2tOTFxEb6+gapX01k66z3JhY6j5+w4yVUWru5FClc28rmsIWW2OmUpuersvsUUbeZVDKAtmG
AvPS5+fIr6hcJ9RImRTQ+cw3trQCI7I6/JB0rY+H9OHbIoUQoV2p4DG94NQgX5TdPu8zanV1jNDl
9eM5IAvRYlClX5ed3VwCg1Be0dFZNy+T8lIxrXGg5y4D2hBoIxyLhN39LSMDDz5WEeY+vM2crKb6
EHyjem5Ss8Ste89ncM9CclciaGdGERmRjnUj8C3Q7pI1irx63t0JjdxFCIll9kzhNa+6+01YbV3O
IbbxDFZSqfStKblTMalYcIUhXMX+I6XoXr87M9Td4BjR4kE1MiCQQgPqqWYzypv8ZMYJ8Yb2EMLI
O3kUj0N++OIisgqnhHh6+/mkdeoVSC6/eSUaMrDcDjlhU1Wb4TsbXQR3j0cNiPIuA0N6bSzwGuwA
GmEiTnwdk5LYuanmzFnBpQ+n+spuShVYbn7aju+RgE0Fqnhaazy36LJKe/o7czf09h/8meJmHRE/
XcDNkz1zCQ2RkChVGunuO+RLkPBdF0IET1QjnDbarM9thm9qWehuJWg7DKQaATfwXYJHpOpu/JzG
uK7aRtrf1T6jYzypp3Wq9oTeTE/OanADrt8cn7vl8dlLkbgXp3pg5OfPlTLV9cJslpBW16pFW1Uv
3MUSy50MXzR26KoKP/SSemfjEzRrozODn7W5NW3+qRfhsn2opprALOXM0t1PN4O/rbVz7BOJ6/Hi
CtjMgTbEt3wiqNNbrikwipSMwOc3vhZHcU93jQCDprUnNiiAIAQ=
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DEw/ZqQkhyuORutGHhs22F3dMmzBWNL6qymyrMcdLf/BGvc0yGSaK+FExqVQezSH8o+8OVlJ1nfG
ho7a2l1Z7J9epoD/sBk7fJaZzR1J1Uxy0qOIttMuKax0BkggbO/AfwWorNtED4ipyxXhR85vckJ2
YuQN9rZSx+MRimj4gNkt5ecMYFaSKFBkItWlqZOqjXZvmBsBgcKvQamY9HvzwonYG7dCD0WgM6bY
GGhqHEWgkxb6iFdT1qz+Va8e44Ue9NdcQMSJICztXwNmdGsX1N+r78aOhpsM4HyDd6TGT17/VQbU
18y4mxQBwHXTN7bBG5ejJMpG50KWhuTX/VAEWA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114656)
`protect data_block
+zRph4L5Zj6VHcdm0hZM532AErchuCzBV8y0szSWS+0/VjopJV4APV9JanWsgvL8mI8XeDe1O8GI
XNip44TRUtZiIkw4lId9TR2++jkX4CZwql1AFDBS6zh2LBRl8S6R67ApUAL0Y3DXbQJi3hBNL0lY
e/qDyo8dyq3HX5kgqCffRE+Y7nyuafKqJ6d4NlSLCpyj17ob3xZUR3e66qtdFAxEq0FJCjPIbNS/
d/h4PVYsepjrQsmop9sueStHxl/NKYCEgLnzevGKUAsDzGm/Bp1+qQ1q4vFzc7ZTLAcGtft4OB6Z
kEASh/F+bL/oLderOoNNNfsUVhMwdtB7S0gERUYfkGgNqx98PWJk9iFHBi6fu9N4h9j+EBTLZHUe
nAruyKufH32etctaLGhRMShGYVWe/tgTfMTfpZ+32VhNGdhN7de0vOEGYfIKFhkmxqJN4uHlfQEZ
lHTHA3zX/YwcJkNLhzKjS7oEkGEdNCS5YiRGCTlFz+hZsO7Vzvdt29BrpQA0CiC6f/hasZtwbdq0
Qa9iA6/+cfLpKcKjKKcR7GMeYmFl9k2mNZRcCCEQEI31RMEIZmGj1JcIUdhatz5VfpFtgkxllE8c
8vny+dK9XhrhVPdt7SzgHSuk3OrKAX1zstEasuZIfN7pMr74Bvk+HXGNDXkXZEr+IKCZWQGgsT7G
amf0mzOQMVdaFUCk2IkxA35DjP9vxF1UvaAkKL+Tyw6or7UeAauMeXrL+wNrZnrgs99sDSpoQ7Br
8aaknI9XP4CK2iT132sZiWsUBFetrvgqm9m3V691UQKOqVqfpaqZyJS8zkJX/B78lIf9bd+PGXVr
Egdr0YLae10iuvLiV9Qji6PMRcRlkdPl4qGV5X3o0Bq57y7uVarYrNe/4LXhOwBLTa0MlqMNliw/
yMfdoEPyyr74u0vO66aBq0K2QLTLbpPRIbKtfuwpK8q5b3EQgTSmwfRcwDVwAjdH776lCEjlRynI
SwtmnyZ+6Z6G52g/m1uO++1KW0LbzCqp2R0SXMuDpxah1IuSg6BllyLXC68n8ymzP1QnfuMbd0aJ
szu1UrfofwkvNxHuH8QkZjYietyQL8BR6xm3b8XEAeBvALHVKwJQk5nvcSbQr+keI3cLHqL7hufL
F/hlz8DRUKaC1GjhLn/sLDdhfCAH+JaKmqwQXYAOcQvVGUODv6hA1mo/GdRkY6bCeMk//KYLt49Z
UCLaJy8pkvsFAL5IWKOj8A65XBkT6YzK24A4+t/MrbjKMKIko0URvT9FIe/un5fK2Dtk3FOPHlPT
HEyVMR4EIrc2QuB4vENlU4smWwW7VaUUSPUY0KrMk2e5+f/fczvpm+V8rAMffMLwTf1mUxbyAaPG
03/fhJUn0wHOjtBUWnMeQRoEE6hAaGxdQSta7csC+Sw5C5kmG78Cf0lvB5YDaOXCUKq36Z1crVIA
hxfdzHWNuol7dkvyxjkDU7jBVhrZ/rGis7NZ/qGFfuuSNsy/S9s92UEH8LeGjjXbqGy2Pgo3jyPI
BOOVlHgBUZudWCfOvqH1oM5tQGty5b3dj0OezSx9DsNQj/hC4JBJF/yw7I6cXwtEV6WqRnaVwkyI
B7eDjwlaiMrXyIlwQoIWaq3oOdKn5aIxNdxcfGT0KBvbWkXG4HqS7ygTfj/eEcFabLzYpoPm8Nhc
m6nPuBs2oBPh6KkU+SGn5EtPLsEzLeJLkOJcmkmxczC/r9aUFnmbGosQjtYgHSkeDq+k0GlbXK8n
+oPKzMBODGFEiOe5Be8NedK2zp9CvpANJ8AC80zo7Vzomk4myRetssoT/gb0jXA5vcTTn/EGvu+6
w3AFSz0+GHosz9cjh/aG99tr0jY7XGWHLRkebSPBOj5LzHVZ4Fe2O92B4o78XPY8LmgI0B0riFH5
II8DZIZ8C06I+qiDx6DEewfxYZtwLxoUy9bU/t61WGUHEyViN8wc5c0kzuoBYBwvjLHDtN4RGA1+
qwKEkYOpS6dyKz6AVIuEw+7e2atwuKPuxrXrPQ9Fjcpmx7Cr+ENhDKcRmX+tQQ/A6Byyv0Aa3PEW
s7vpMuM7zJIYbFgzNfYmUlY/Emr85Xybl0a3j0dp4owUo7pk4u5L/DSeResk9EHK8PUWv+VzP2pX
UgfDa+aYZRmTEKrplLr0sKqmMK6bN4vBvxZnMwxwdWT9oL8iuW7RS/EMBCMrPPOsPAVQlKUf74Y8
+VAVSOihR2egTgSTCH8ZlwUKcwF8AhLpZw/FdXNY9gnRumtaysZ+sM0h+qIShcnVg/n+RmdH9kU7
CFgzOrX0mMcrQfr8lBRx18JYUhCdrTKKKh7roxAun0xd7WS+m7PodeHxQ5koLFGsW3JsZxh3p1UI
3DyeOuksny+Kx6NK3+rqMK5mPMXRKrO9xMaX+Po2yFdTzwhL8VGg2mEv2IXZdLr+gUleASLzq5C9
IOf6yZ/jZAJuDqKFs4y1JuJWssrAtYURt0dTrjzIaZrPDXgvATunH9zkZcGOz8FQyEf3W0VeN6OE
XAo/cHcTzwy0L+PwDxYY7roZtDbDQ92vu0HU9hBSO33+c34YGSS+PqU5BLssvsZqIrqWQXFIdZj6
3d1M7IjL68Mq3aM/xvwYf535764cdrKV6spglYWS3dEqlcggKkArdE1FomZ1uuTJRwne30TMqSaA
1wBm0HjepgeD1qIXdcMY2MziFIChChT+4NDq7vsV2p60DbEEbPvBJqmN936tvzSSyCoSmkZLDNaE
paWwO0LAVTPuhiYJ14LSf0NQf9HXdsbfmbB+2hJ9Pwzs/g5VWIFBGpqAV+8gOnkAnIF/8n06Cdc4
1a6jMk2VyD9rF05/FhvCwtIf65Te8u6emVvOttWHxKPbEiyUcV/l6ollF5UNaeTMU8t3WBHSNl2V
T3/DZ4YM8bV8r/dt8Wj/adtQVlOhlcOZvMyQxj3NIOAyAlim0zXeTzFiAzDjf+R7j1EBhE2FuVSp
gV8tlyMry8Gudoc899BbzgYnJD52EWkALJOLh/v+N87OK2pV5ftT6Bd/Na8c91A+6b8I5JEUyD+t
swdAxi48BC1wM0geapla0tyXMClXamAuprFikQybzILOH0nLE1dfoAfcoYn7Cfnr8FSCLo5ib/9e
UiCZEfkJQAp9JeX9We8MPwZ2EkUMbI1QNtJNqS9yCJQveR5sYqylakMdr9xuizvY4zgLS7Id8dgR
phn0QFKb7ar+IDDDehF15MT4LXmD0YEi1C/yAm33sRffk0sPLJCY/DqOHo/boo/v5uOfR9W+QgoY
p4UuM4eTjnIFcrvkf4ohBX/kbAwtN/xdZBF1kKTnHGcdNZfsws4k99BU7cxtLZCm7cAw2lYIG0IN
TFs/6e+r4gAemYetVNEPX3D0uFh+blBsaP13DD0+QNXEXBv9QPfIIlOoj691l28HTt3RG1z+t3mr
Xp77DlQoNwvVcJotlQRLeALWxzSlmXAmDC56btbcyb6+D9U2IAWoDLcASb+WURlQoGolsm96tpe7
/lVI/j/RyAUwtEPMcCHaQ7EBQzOuVCCe00ASo6WCeOXc/jnjGRDECV/guU/vsAGEk+43vc2oLAJQ
WtBrMiUhELBzinb2jc+vtGcxOsdX+ZCYFZV3ZN0AGejy/UfJZ/URSt2zknoZlOJWN+9l1i+SdsAK
xIK1j12ZNHLKtZxdn2tsYxo9FTPvm/N+F423XfM/A9glQaHPm3XjhPoyuNQhO0CvF1fHRCTiWxKv
wKqNLEGoq0FxiAM1HmUAPiNQGFIm/ge3A7iZd5UwTH5Q/WBQP6MibDM1q53/4jp/8CcYKH1UCLjY
6VWuwL4BEFA/A/rmb2uOkYE3e0RJLi+Z6qip2bXOJYQ9ERrZEHJXqzicUVL4CsPrfRGsed218C8F
sZQL75cx8zsUC9mWdktUTizJQVJCIWltbc4wAxe+eLtpznvgBLOTcXpgqKOWi4x04Po5CRonWfLV
aiW/QGso6SLZcOdLJp+e6kHixHgwxVAkifzV1WNKkd56ikD3vyAZfb8OwlZJsxg/Pj6i4MpBeX5o
g6eUQqJnVXFztdGXruxFAu7LfQNj7hICYv/USI2mK5Kr5bWvTRsVbqZYQdTYCX6yQqnB1J+XWMo3
5JtPtURHQe0PmonhKehiZBgcHLfKsMVx/K0DBVf1AA7VAg36zIBEBjEZCMn8iQbyUAxCVvPE5n1O
FYMMQex7R3itmeXQUf6b3K6zPj0DycVEx8oI/Wn1B5xtb1VvykLreMRJbbV4F9rGhcsg/N28UHj2
WUqP1BeivTxKHBDUtNIuam40ifGzJ+Z8dERsGN1XzEnxinU0xP3uwSXpVLWirfx2rnonF1BywnFO
NWNFcxWuaPwwrxNGckggwxr8AJZStVZxiEEs12q2yW/hfOP20ewW/D2ta5axS5Vv6jHyeC6xjm2l
nideXWM6ytKW4T3mXvVz9VtWdxGwe8aELvgl0qUfOT/5hEK3vKQCZWtwNqrO6V6q/23CmjJBOvDe
8gleb+mQWmXY0RqqGbb48gXGMotlJcaNjpDpa9JhyNX54aqcZcSslDdga2LEWZYIGGwkLucEPGw4
Jj4qatheKE9K9TvddYQoXrQ8SkYmk4/CYjI6D3wvFgyAztZHyA1rlKDQvfLtS+RTVCY9Z2PhQeuX
vUqs4n5RfOF90pDi9bhZXFI3SQYYmT/lwedN4Yce8asktM7HxqRF1mivW346mhju1/necJCMPX1g
EWXJetUodS5qp8/RpzC801htzsQpuPFNjXrGzOl+tDhqKCQ9gmX72AGA570rguH9ZvGVlOTDCLIE
ULofreapeoi+NpJQXkXsnqO+1JOwvSEoLnnfBSd6O39eAJuGSbIdNHaOL3ofQxmfb1DquoBB0S2p
P5BhyVC59c+r2gAnoYqpzkoPCxv/iD0kcZi/jtfrcgOr53BU3amDZaOzrz96e1EJNEhmRozcvJfz
z8kdbsRbPmAIcOQrbMzFav0m6sl8h1Vr9ZIHi7ODls2EWu/jvCY/Z9/hfUsTDZlNa9rRU7ojF0iL
ZOAZvbbeY8/Lxw2ERsi3izjo8REWulEFiPbhNe23VEfvdpT6FToXl8/xx0n1F2iY/La65hADSwYQ
2ue8o5Eqerxd7jde+dhwQ4PFtC2WCg0XlxSEHv7OF/0VFGShYNv4x/fHmNcIrY0aiwzMb361/PWV
LKJXyKJQwg5A/QO8Fx+oBL9SrYiWzyTRc1WhOlGsY3Jfc0QGrYJyD3KM6Uczn37mpLq+nK+mBg7M
2oaamOurBjQJy69SSXDlpbr6/3ZOCFXvHiRnrzL3Yvg6vV/R/O5BDzR39lyOYAMHkbE2i0DEqS52
CAxqdTDTjjUKbVVdlBVyQPI3C2IWa1+K9FnK5/0CnCmuDcjspFItxJ5avwFNCZFatsC9AK8t0hFh
ztBpM/XP6G9mV+Nudus9cQWpuAMAcWfE/fxEdNhpwlUEA+u2g51J/b6azX2Q2nShyhCURZ+Mc/Xv
60bAoxhz87+gZzk2pyBlUaoG5uQJh8u6Vavz5zoTvtFd00Y7gY96ThWaR42ZlAmH59pApty95iUy
gCRpKZfCb7Umg22c7p2I6kh/E9fNZ4OO4T4MIdsmR/rfG667zTGXW0J7YsTF7Gapds1GU/s6L++C
db6jbxjEMyUx0BR6ozAr9mBfGl+jn+OTfpCs9ycE+3DneT4iK8Zxkl+qX0SKIM2apC43hH1cbYvy
ArZMrNoPYdwfQxAAXzKXhrswXrpgn7nlpZlfZKBjq+TUmEvimEC60tiMTjjQ/UzrYB0titQ2feXq
G+RRSNDosAK7jWsOdIt5qMpKW99zYPdvilyepU/dfYmc1x7B9DmdNQpZgMbTM6+q9NHa5xqOSGTu
mz03bGhcO7I8UjlORlLfw3TdXS2ILbDO1w+KyD9n/Ua5uMkpTSZRxPWCBy+Nv2aJWAd0wTlspQUu
0al2kZ9Kj4Effu6agOTvURsX0dI3F9MTkFmgJSJwXSr8GkO0X+uas8aobw2F1Yjes2vcMfwAhzW0
7hhqpz87zJ7YrzOcXeulL/laAiuDk2YsdpcpZtVGCbcWpHBhV/ZwTJQ2hIW0QwLi97i0cDCvq9hm
2gnz9YR4ytvTBsUIpKJvlRdq0iUjzGLoYCH7dZ1+FTfBopSUNgZDk+xtjfc7qxaJT8jtOAgf77+l
vmpSTPtiCkMBbb3CX2Fp36jYNkKYN0oBwph+Bpqo7DzRoRLtAP6aD7OzLWV0BCtfWcJn5vLUak/m
HRcAG2JdzO22zJoEujxIVHK7ARNGIVaeRNjm5C8tv29ujzCbspD4nRxb+Fyi1Iyor9t/mX1BAI+8
79KEOQCiFLJmdQO/zCAd65UHTVKwXz+37ockKOha/2YYe/JzKM6aY8JnMwi7uz1uNfkgIAN+KO1F
Ol1mj67S0lPdeuCwRWojbspxMp3OZzm77IP3JU5wiq8o1aoyPVuW/Um0dkfkreN8FFhdIuSmGokz
W7K5MQrlx/3G9K6zKHVj3TsTqJhaRIrI67gYtKqoQY53jE+8gbMFIWokKQfR8KTTfbAVVqkelcoq
/QesFdc1vwG09Lb3aCznIXovCp1hsiWMpJSehE9y1U9hzeBx3GWohKFBfooij0+1a1LAFQrP7Xkp
vUmSw0Qh4wzvqk38m+b6Uk9vST2GgvxnEOYiahXKXXCt2Pjbq70fP4PDw+KSFzifS83k+rUHu1Zk
pE+v4dUe7lHEPQGg0uJqBjgBwIrfsTFx2iaBpjZ8L3P12APq1NAMdPqPvlzqxzJMIljSjQDRCzZY
jykZ0FrCXEM3I1F6wjvtQmrm7x6H94gaHQgdarAlUhfl27W94daIsZ5Bg5fDaR+XHnwh/sJ/adun
e1SRfjT45cFvEZyaRGU+Z94augIi76hlgA+Z3JYz5X5bs+pb5qfx/kS/ibinFCRpMzUtkhoGwEtF
F/HaZ8VlQXGsRyHN5APDvFV0JA+4e5vA7xwE7IfWevhA1V0k+0rsSsDX2VTJo1fQt1+l2jl39pUm
Akn3gJ6Xw7riUQm9v9HXOwISFw0Xag0UVfPprTeq87vbNtfwPxGkl6JM7NM+nyAnUpEc4wQ2Vfxn
5A7bnF91dstoeOGNFNJtYkOhZY/RsPSL3dGCbxmQrRR7bjjfaE4hhJVUX1iF93rBio0G05uPg0xo
XqZyIQbY0yPFq7jsRt+exe/oYmDCTcPB5pHUOJxxY+TYwPb4qSRh/DR7Mdoy7yHi8ZAg8FZql3Ff
kvtQ+sxHd4PiS+fKcrYvZygPiscUIhUp+vsRc4VE7Uldh4BucVcfzCpek2yrhZ0d/FYkAUD2HHUa
GNOcMAutZO9/Xvg1yt6t8bvtZ/Cu6R/CMHskpJEttcvDvAQvsVrf3awuKZbcJg3C23MaIyxKNEub
oUSo3W0hnYIGorZGsHfSWvcIypll3xQFHo5Qs429tpzD+RcQ6Bx/5/vA6HbpbN2yqqPHTXABwB9w
oWISkue1uRD4I8APoaYijHk0kQ3w0mSGq2AJwZ+F/hnmDsXFMhkb1jimUuzVRvMJ45ZsNwDPH5KT
sTobF7br+SdD9W7coHtZXHc9l71Rcz/1Jw6oYanMD4qIB21gRwWplJU31vJv51ujfLddjJCqnxo5
RxDDiWf080Yxnvr1cT6uAHD5RB4lmuWdqmlOA6ipNHyiz+5rKb7hw7jSyqK3bCabBD9NchLIKnWQ
sntleag1cXYVVCg2FY5m72e3V2Rk9OLxF3O+1FWtnzE2iGNRxuEI9BxvDjRSL8wcA6j2t4llTfYV
i8gC4olQ4o5jJ70RXWQuS3sIhWwH5fCRg4RyKxa/n+IfdQ62wJwKkB30ES7bDnbsh8M4O+kRXM3h
u3/eMohh0U6OKcPq8sfx/LQ5lYKhWs18f0QDlZtCT7xGi37cGgno+im7u4wRxNcz0hAhoiJSrWuU
Es3G7m6UQCG96nSIhixZELcJrBO3rH6+a4HmF32NawKIAmRZ07crEyict3mU7A+whAuH8ZaVNikU
307LKRDW+5IA5F2/doijJJP9HnEUaB63iJ/KS0CtpvW5arAOz22zBG6xv2fsjTbTnYp9ZiClMvpD
jnQJ8m/zM8ehhVKlFV96blOODMpIZMyVvAVs5YvTRsGQEFrzcbIV3CUuYpWsh8LwTgpFbPjt/jja
h8tIL3mKJZdRV0nY+KnXR++QZrlkKvpv1TGPrc8EhfIJoqGhVEC7/Mtf4W4CSH9jY+K/WlLYXNyy
DD3NdxiOQdQm9sibidOvWfgvyk4YGEsWxl7yA1DM2aoeeuH4FUjh4cmY9ncJgs1N10EroXIf5xal
ehAmpJg0Sn3o43ftArAY502NmZvFzdgWJIQ6JLpG04MMrIJArztVo4XpaTAj/2CUfVN1ybqSaHJJ
cPH19f71K3oQ+hr1eApvv/A0zviacN5nrP8MvdPhD80PrtIU1VX32FLT4W0EJq0GGrrN7PJVY32Y
AIWi192yINal5SzwY5j2bNXWX5T7zpi7yPy0wv4nOkjgAZTp7oBNvvvQUfxwLoBCsWOMkK8mFTii
nl1UpjUcyY5A5jwZS5V9A67l4W5yUBUxK49uL3EIbELx2JAopYuEc4AqDkuT/gFrZs/qA3GlFDhs
IdRZZeQN/vIcJIFOQRBeg69uboaWHA9VTDhlArSEgZs4Vmfnq2qAzsbS7IuPJlKPme6284kfnRFh
/bQNfAkmr0IjqtH5k/2pe4/SoBJHM6WqyQl9jGcbSCewRYgSwoaHNtOC8rGv+6ESVTaZ1GIOYtfv
Z7DTX6yyfJOgySuXZlOHiBcq/cIqq40t6RhivWJPEqVkEumrTPGH11BOufKG8f6yJj5MHdzsrmDR
mdVbC+2N53ASxdZB5xlUTa2UyQ22BbZQVriL6A3Xj0Grs18zGrZaqXveWrD36FaLEuappyc2uNq3
fgXXFhNkkKAckP/UC4+yuar9gl6pzHVYE32JEr3Dfh6ytiksE7j5MPzpPpj6gzKDKtjfv1ChKsrQ
rca026ulbLLO62Dg1/CkSl3xaGX4pCbQgcp8ngmBcfJayDSKtVAKmickO/RR8F+dJzHu7HcbmjEv
R02gmx2dR2PD/UMCp86glDNfzTr2c9TCzmveFMzuAs4F129h8C54nOsl3NiiO7Cazo9JIGlywMZc
IK4wGbHHmBJTrn4UzerXPzbS/8x0NuPDZeAscxBBoKx9r4wcSRZA1YHGRH/7j6wIWt6+/sBqBWiS
9GRHP7L0sR46VvKiv1KBJ58Bm3bUgZ3nGNEGxn5yJTuZCj8upsUf5MGm5Sa+ZH+o/KGoJ8wJcXYW
CWbWNGAjoATHCewAAzB2HFZHWnIFMziKIG8YvMOzc3Pm1DcDS25bj9lkm8ml6om5aO2RHjjkx3pe
euwdAe9Y6i7Y+i44Ahlt3F6+Da91Tr7kITDhHsYfi7UNmukZ6JI+a4shhzoFe2g8A8M43mIqD4nt
UFulbDTfiDR83Vt53zsXohc3vptYHAWpj4qMaTdglH8Qh58HQPwOm3LhEmexc/yBT1TaeCjR0c4A
468Qvt30I+34D8W05bk40Sltaz23BrMR4HCzfClsJQZLmJnyOmflgXxpCESaLoFF1eye3WKrVmCM
VjSOtnwyOd61mnAZxnlE89aCXCjcSyMX6hiOFgalbIRhJ+9uSMGBT/kPltTwxQl/fcyz2BYWz4ed
ewRn1y3EyO1CZ7PaZeeDx7y48Mh0NUvp3X1IX2qaRwgnJtS4/+GMVKk/YG2NQ7Hcalde5s56JYWy
ooHplPtQyd3VB2MFNr/V2BUNu37x7CXxNRWIPTigWFQOuuhQeLy8QPu4ktQzLAsS0r5QD4ZbQTax
g9Fo61kBpw/eCKvVs7Pen3wBxKNyeAhDA57C3+bZyx3mIKbQgEvcvk18CQLwYMTreLY/8+Gh/ufC
uOAKdbp96H/Ni0FcS5w593ERQGCeEZZTVHDx98STsBm+18GAcy1tkuuvSsLIm9HpLRus4p1F4R3L
IHa8chENwcPEIaHN1YA6o2muLmTpC9IIhGB0y1L2lmnNpTR+CYWSCsnHc2baWA0MJCWony3OvPhN
wmb91nUXyKCUXWstE52orwmbMN4rKBpA6pc9lAkBbCB256ee98VOvpLpDHQ3ybtSbytl1ihem+6o
nIhkXDVHEW+9D4wFWq3SBWjqxPGsu6rjkGhbr7oMEZMGJ2g0a8MJmlcIqoNvfIi4r351PsJu0F8h
B3LYcmRCZzm9D+2DLrUzlRJepkar5Ydr4hEAs18je71YsEkD6xJJa9n3LWgIFL5QKlan+Er/Yofr
cePwOyqCpkwrHrTfz/GbHPTjk5fJxKzCVzQzW2Fcd7kSEwsEey0Ga74FoytAMBlmNRt3kw8gno9o
A3sx4mG/MQ93+uI/1nrhMgSWxBv8TidQpQkSOhoNVJLd/xejUpYwmNAfTUg4BzxJpD2HcNjzn3hc
eGRgZOj8WXEykT5MFxkAcPejS0jjzcF5KqUJ079sr5WsnKaObHUkfcH3DYRmnEBzSF7eUIWkyoPL
fMBUuS96hrLkSKwcTaeHJJWChwoP59XjkjBh/TclO1sQfq2mY9jsPFxvYmnWRj1v7Gs6xrN1Fb4t
lm/VGcORLNjJIKuaY3nksq/A4HnTp7QmHJBDP0rWbDO2tirn+vOZFBDV0ZH1fUrN8uPf+bfk3SAj
C9zMpHxv846I73b4rZ8hqnBkFjEJ/ovhdKhgNyVPmHbC0jfBFv3oIPqbLh37DjireH+7ZNFNDbJ6
fu1/3xqlSZsrodM/c2jPVA6G8hz4GH9tm3uG71wwxZId9CgCQlbGuvatAqMHZVrh5jmzixH3Fs59
N6PQQyvulUBxijTJYubMP8FYqaeuuoTKxSktnt9nDEfFLsfdOGQh6uJfFPjE42/3NmmP0efbwkma
1mmUpltC9PBS1WzuiKDC0LX9+mNn8IvPUSu3QxhMkQbrQLE7KSJImnlbbpVzL9AZP8gw7HLLyJac
/yKlpBjc0jp8APF1ApAyYiTd4uA0Ra4HK1OMCgYnULwBr97cMc1hOt1JhVDkq7CpU1VacoeWKBlU
6Vl1bZDf3bEMtyDeZOJ6V4YZOY9VN4J0JQj6T9UN4mVJxjhUvQ3l29cCpjtSE+JYWSumA7iRPnS+
pE1kbGisIxtoFKutYvC4sYZsIgUIf4M7bPo3J6dfTWDuBeGf3ZBGCm8SrdzRpEyxJUMnAAtYgfyg
zUOD59c5PLTVjKkgHSH/OOEZDP14Izydt+zebJOJ7BmuIYrRUq8TZO5MmWo7Zdv9h5UMrgsaZNOO
O/cG810ROeWf8FctdQRPhdNPHvNzPR5KJaz0wu5WrZjZSZ+uTh2pBuIF+8kliqIhSZWGvsC2OR4G
fKBJ1nWzNpBFJnpQCXWtXhs5rwzGG7nwJ0E+vI0yZ3ViFQHm3Itv9GeShKffag0wkF18YxbvshEG
66MTbM06yGkeff4Nj1fcKfIosOtMYTzQ/mD/6IQMKbwGaQHj5V5mgSUHo5p8GArC7qm9yQ8Fjml2
SmNY5GyT5lZ+O/D0Y9MP9yNGm1VFNbLkdiWQUEZn5YLFXZDsjpAW/Hxl2rgFNeQyBhP0gGRX9M5c
/kEGZ1Tuhq0ebkqVfBKK9Rs7KftxaANX2YFdmFqZ6AhbnPO+h0sTzbQR9aSBjVudzV0HgmiJyPkA
S2JbRWJ3v/3wl9/yX1/HVjq5w58OLrEiE9dVxx9yFo9rA6rxCK0o+YfSOddoUtH6VsBMEsjs10Jd
SEIZBbaR4JZfVJzv5a32WXbIPw7/cM5jE1DBYwXN4db/fO1oLvyFSQCeBBpBYILoXQsyUnvu6eCR
8QQzHVV3Cl4k/n6b6Dg3TEtpcKFK/PI2diRlRiKHwE49+rBrywS+6gW3S3m1xyLdIkVdY286e3eT
3D99GRxtUwKCFU+s+LWrGH5jM1uHP+G2qNHXr6JXbrWFwg6aAd6HqXJJn4ZfNu9yihSYPBwEE1Ur
JQcKc/vCBjG39asuUV+Icjf0d19JpA/59XrHxfmrGWwW2wmBQAnR90MUqFiROU57pye/HjkmTXzY
lbS223IPIXjI9R5PzOro+kiJA9YTnmI2bLWAzKad3snArDBQdKPssTPpfd0FHVEi6qtq7AQOR8tO
TONvckZapLJ1zZxQT4/kuxg8MjkFaWh3tmS3O0S8wEpuB3TsY+2zoaI1d71OCA5fY/BtZgELBgbg
G/Kyf+weX9+2w0FEB9gL0E0y0ZKdRLLWSjxT84Tem42cgwtHfjuqsI8u2HZ2hOKcFTlzDKxBPoaU
HVePLzziK3uZ+qUeWvlvxLFnr0b2BkeNdFpxKRWn32+adqgYiQs7jbaf+nBzfVSptNDXUfOHwf24
qoWldYNKh1Ss8DT5ROQrn9Kh0OSI2YlMv1o1nHSJ3f2+x5m2EECcNu+lLbpEixHeXBM2gz8DegCe
rFpUyyamccOX/0oLGCj9D2DSKbbEOf5U/7tyJU2FmmGXYkl4sDxMYgi2uGWnWXiMkX7b+YM5df+B
iSg/8OB+FxIsmrD3Kn4IcLZ/GoZFxqFYPw5bCBdPHs95nuivRSlxAmvV4bVbKRbZCsqjFCSt3LVx
3EFjB8n+jQo6M1H8BZf/XBqu5AhSOSnQISo2JVwZhwnJJGblkuAL570K68NikCoMvC46w3shCMWb
rxuibdguQsINJ86Pjjv2FygKXR8rn2E34FxO9enmpjy5qmzTrz0L+Vy4ghd18K+QiIVbSIMC+fcd
eEJfka05cfoAbWUc5nrYuJH65E+SVSKIA5LrDEMcavr7LNArkngVMpKh04dJMZD67xxXturCnW8I
fCK4mq5U4bWh/7DxPkoJI1p+t+Vc3OPU1pziDPr5oTaie/YqwNIqGRUmB0PjJAn6EcMbvp9qQIc1
1FjdBKeuhdh9p8f1JIgdG5swVkYmB63PX6mph8r5J+YHcQViunN9AFOmGWtMJAvHLAqEFhjUh10e
k00rK8hzGc9OBg4ks/UJJWmIf+6Gj59EXXD1/O6B1EaP17B9OLyopepKppQKYdl2leegiJaZZI1h
hfpCSt4L1DGvR0C7aeXvu1llmXButRzjcmN9IJzNOrlbihXMdUUU9uOIYMFfIUm1sdCB6qU+cwts
/9VsnsmlWKpwb66bq9MX46AhFfBmKx48+TxiChg6rAhWATuAHekxP208qpwF5HuPBbYcdI4qQkM4
X57wFQfyGEw0gp+NN8UjWN/RGoLbqrUoa2uKJ+rJHyLW+pHC+soB3kX2x+nau92nANwrAV7QETTv
8/2U8QiASodmaHzclkMx7FPdfk/I+G8EEiE+ND0R+Ez6rHZ+cbbBdlL67co6z0SWSVvIfy1zQhrB
4MO3V7QiiMOSyP9mJDwm6WyXzE51YcQ1VhVqPbzHmo6Z4wi26unFrV4Lml8HZn0jCrR/qctGgXwb
0rA8hgjMgtWkdNh6pNh2XqyFUaGzWc6MMufHFvWd2tRwDSUla35peCqcLb62cIji0xqEjNJwN6FG
XjD0SmYWAUzJsgJwqK+QZW5dN0k/Ee6o6QlNdTlCOwKEqHAHVHytR2jRwVdDMfUjui0pYapNhCev
+GzUTuFfnc95nxg8m3ED+mcm21W2mIn6UuWdMbRGVNgcC5PvO/FXAO2ok6vl5bS5BzVoXWqCogsj
diCBviZ9rccPu+1tPm04sNJDShUTseS7CjfOrFT1r09lvEad0aGR4QXgaZOPhVBfznoKaiEqNK/c
LrdOe0KBFzS1So/0EyvqFyOIGP1Cbhkh8GUGTDsOUI0s9ImUujD3+yejuO5tORAM6nUuKbK1P2ce
W/UxUCvHRwL/WnYHdX5+O71v1vPEJtER/gbD0A4rFE/h+WhpePWLW5R509eqZYMwMsmtVgByRR3V
VtRIcXdoFs/JoMwMqfRveCUClChBH0gvr2RDn7/yF67AQ4Fs2wSN4g3hSKowfvtwKKHnKo3GDXGC
em5JHGW8YLlJSvalG9ks+uzPfRZ0F3IsXFBRTi1gs5BuezlXHk0mT9eNSm6ECSx3+O5LSNd4QvZS
flAeYEds6YqWfGQZvhcs3bLsLV6RUEhpqlfkOYHpK8xdVkmeNDAQ1cCLk+aTaGqh8myCiKyhepFG
/3ftvbGzYzUhYtrDZtDnL4NIs0BCTiv3gpgsiKU7vSaVNyUg/eNAcnkq30q5hOe/D1FNsZ07d7hn
tkNuYi+1u0JOCh2IsBc57Q6+8yGQmVFCb4BqLm5I+o4MuFwN2L7PM7x/FwcNgqTHIwei2LO6WRc3
TF9nOwoEP4KfKyrsNxWU13Dxr0VycgOOTE/U8SsAgZhTvYS/tvnJ8yGQDF94Le4sAhv35o9SQSfB
M5Sku1ij5aWthzNjd3ed7RXWjitDexMc5wCIJIhNsEExUps0Dwskq+RsFexcis0HMoN7LH4QQ8ya
2/ufosKevG84pnNvLBduli7e/GJTSwiHge5sbgcc4iBbA8gijUp6w1MJqCvdNY+tCgjVn8k726cM
wB38JQeUV7lUxgPBnp4HLwsxiFYeYBZ67CXRL3VzXc1Y1cFzCrRRuQXY54ltuBtooQBKIJ6W1brS
Z190n/i7PvugCPJ9u4C6bdO9TWfc5Vmip3SC2Xtu5/WlTMbS4HNi5rD0HCEGf9Z7j0UCsly7WVqt
cZ5cRjMRdyHow540H4C7/XTG/RxwyYbBe7KEN21DapqkOnNxBwYbfHmqRxntMoQ/aWxvV6WrGEim
P8ItL+SBwM/+NxewxCPDi5dJHZJFU8/U66d4R6FBLx2+NweJp4BaZbr1gZ0K/U5viOIaLqoTD8/E
2x1VeegOZ31I7JRJoZw670XPZMedIQKGJsL9a914KZywRXkCmQ7GaOEo1z+AhKp0FI29FQ/0dDCH
ytZ53yEqn9wTd8gjy9IIWdql5u7EXC8OaLt1uqUIbNlUPuQ4KUryoAyK3HAtnEepGeNk4cuf8C6e
IIIywAJ5FeyPFEPvkfJtOu0Est/WQ/rcIFI3GL402uLTGDeO75ISJKsqUgBC491GSBPtWxS56rJM
EfMetHSKE/NTIGyPDByp4PnWdOf0sv3DlPCfDayeM2E7gIKEPWi1N82YEiWieu2NxhRp94ZbWtsy
FvmZHyoafIdr1UGuDN/fbYfGtoJ5mSF5/PUz++w/xXI3FbNSuQs4INDrLw1xva5SXXt3r3GHvO3X
RJ0PBBKkcRDWl5ijf2YP6SrJixkKVUp6E2rWV+j/bPVW/67Kq/S88KZwNBPLHmbcVOl0pWN/Abq9
+1j3rnNkoweiJ380c8Yw0f+CG1XyRYWMiYmaey99p3ZoF3LXo7Dra4wdW9unuoYyShZfkxU5NTW6
b2la1s2zR0nEDzcde0vgAjOslfuZR3aRN6AjoYRuzGThBixO+Pf7fHNDQEW1nHKmqss4PjwiTq3Y
63RhC5eXTK7azFvdoxpHKHncx/fkwa4VeV3YdOjXlFptn7TZd6AAXBQQS6ba26LUJ7I9JojoxSiF
KDRt8gQXSTDnQkGtdCTdL3u1PqGN6dCPJa7EDEcGFXRZr4VGNugyR1i53DZ42dSUb2nQ/BCedzYv
mfIasLh+wiDraV3a4ZT6JTQyQJDNrUlRTw/xRrdzrIMy7T4Ka2BHQskfamF54cxqZlKi5RLEsdtp
KLPB9eROMwXm3RFilu3YZQCBoAd8aZ3V/blwmgWTIVtssfupjXCV28Y8QytfkvgmLmCqhIbcBjDk
lLFRgLVGLYIL7dSuziy93GvlhGNwJtgNmiJ9FCxNofkY3FtdSNxkDB+aRFYRlsh96qLqbPf+A5WA
+tmyeX27mvMCVZ1rF4s6A9a9e9ygZ4lsf6OS4exu5Ckh7ABBj5bxIipLEEo/HUWpVKJAllaEZ+iX
A/5c8ffh5fPqZd4P83HDML10gCb68WLkNIHFRFKLvALdV8x4GRl+QZEC4Y3hGsC9aElfX97Lq100
g/MQMAv4TujnM7Rb9Cd9Ksk3WaGkb6vNH3avIiYBds3Sgnq/2jPciDQG15z1sQFfgneDjC5/X29k
LlZ4dcdu+wncfLOfazF4Kty5fO7QWI/aYri/AbjGpCQX5qq0FWqYaTFNYmYgz6+1SD0O9RvrIWZ9
UKWUzsXTqcUPK4aGmvh1dAMbtT2NNe/X2uItU+ppNZr/rjzjuDasQRrjOivrgqbPqDvMsJf/gbpC
lH0T77ncuMDK07gxA3bnh9cKj7QWrJUSiCnp9RGnmbVvhkDDCuf3Ci20OZENXW8xCEZz48pPUQ4M
wWB9EmAU9dxHPewz5hSq2ySPvz7jTS6jiD98JYhKPyWoLUsI7N9ph68CW7lyfLMkOlnvaJYBETfk
vjkbQ2Ae6S4Zmk8oAWD60atkVF6XcPgiS3PcSkrFXQ1oGFkIU4z7GdZw0dciJrCHoTrmObgQ3LbW
dk2IXgDNfLiJzR3Lp0Mc2MoHlGu/C/wqNNvcVN2+leXuoBKv02+Gi+AfF8pyvhjmjzCg5peAU6+7
1gUbHgpx2EqfV/s3h18dTu3zRl+GH7qz660SK7iyedSUJC4asB8QfLwujB8l2/DI0GQkAGzD64GU
ZnEN0mtN0uBoqmIPq1eEWPpXcMBl1Mt1hhjFUaB34XLrMA4WYt2+LOlmc+0PuPjuZaus0gv7AT23
FUrUwjlhS45ri4fftd3yEPwk6f8V6UzXt8eDG0qh1iZc7Wd4U1VwwbhB8tbzo/6+pKqiDyRzVV9U
38MLjvTKCUb5eolZcqib1tG8T4fVZRjKDlAKwsJk7yFu+EZniRaJlLG2KWMQ+oqwBA4Mw2/FE/64
aYEQ8PpMq5vMAJ3WL0HNZDwpXoWCV3IU1aX75kpJkO2RmJGbInqXUOzSmgrHbNdZd8BeAqwuKkSe
gshIyFpd5Hll0UEVWl2hSANt3QCxgz05Q9f4QXSlx3zxPuxCr9SV37H7i0QrATX7ILRfYth0wZ66
GyasCNLj+ShUKvQgWSv9yZg4d4hqaXhh8CCSHAzDitAWCP5U9fXZJ+/uUiC5K88yFzEdfH5wGMmx
Lmt/ABSWPwW9rpog8Lr+uvuDvu5LCRrLKxwHV2PMePpgn57mALzzH5E/2lQzOGgfPT1E+FiNgNjO
OVi6rVhKEg8lcSeteLU8wXZNQMxKCM2hBsxOF2AJh+Fw1uvY7TyF/c1C1sw2n2P+1XvJyoQdkGy/
/YkkSxr4FawsGCvhbBwXNDgC2+qr/8rbOyrfK3rvqWNx6fsXhAv1fmS6kVqLTIlncFELOYCCioj7
8/RbsBLzR5b3nEWxSuiGqPtmX8TrBHTh/K4tUr2gj6KMd9E0SB3CZscujSDAPWAO6tyy7x8NcobK
Bo9a+qL9uJyrUk+6GXEggRyvEOUX7mFdeZV00fOIBkoFoFx6xRZ8udmECCsxltt5AQC+ZJScK8/Q
erjgmsFNiwCX0SbknbrZ1UYJZ00sjLKA3TvYo7ZrGtbQ1XslNSmsLeMVsKIlryOdxoeUqZlCyc+n
FQ80TRTRKddPovNfSGLv7R+Jtw39ztVbLjdqnNRFl2FFhStpLwk1tdjaJAS1rUAtgR/FE8VmMrF1
9z0o35gL4qBv5yHf3xVyzYb3LMi4Z6Nmr7/uTzw4p7i2ZH1hMocdJGJTqk+Dpaw7nhNRHl6Lw6GZ
RvdrY6EMx3YZrzwvys3ULJzO+vX0yOz3vnOJSb1uaaXrP0VJFwJL9hY/uhB1FNU+snSwjyS1QXIT
opBLhJGvGKFAzz9j8NI3qWboBcg0zvG9G1e2+yLPFmymeAS6TuGbjymhKbtKGRe2OciP3MAgO/e0
yrnlGAuTjTISQIDLESbzH4cQRiUnJq/2mgxx3BgXtU8POd4tOpJVK9enkvhPM2xMFlR8QU+F+qy4
pEor8emGJHH5TinaV0C5PolKSUEY4rbVLzVcPZ7zydPbwBuGYWuASGcM3NkYPfW0AxUifIEo6ojr
/sEAYuSwATkJA8rV1GsbRxCDgBR3E91oferWxoLp2qwIT2EE0kr6gthcOithxCjHQPUEIOAfjWRN
OG+qHDB6vXkMbNLyZ0IoR+NWHgFmklsPXQMa0KyCV91Kr4/fLz9/NyaPhhBV2DnCeRp5lbt7Vq1W
2iyWvjc/YtkjT9aAOKaKSakrtXS46ug+IAHQfXjsWnFQ1fGe7rVR3yX/SnGT1yJlE1LbuzFtEHXX
/Pe0w8hxYEYwrRkmSj253v0yhvwAtb97x3NTyacdr0chQNf9c/YJcJYk41xNtaIqIvLmWGmYrE6p
qDdbLT8MFbZz7Nh5nWACQ5ssflNghZFRoKRveO4vRAMWq8ROqEezyM5Ua+tcXuSYjqVFrBtxvNJq
x6LJ3ntvAacrm7Xn3g4WJg3jKgqjIKkHNrXEhKIolLUhVs4ucWw4+Bdp0zS7AKVYov6dTvE0btRY
CHiTa0jfZWfjF/v3kTI6e4ec+r3hOj30m+yzS+L76Hg+U4nvnI35QzPFwYc4fLMOs2nuVdWjfCsz
PduoKZ0cEu8Vb/fiPL4F3g1P9R5rVHr0rh+UQHesiSK8+VoQ+0REaSR94gtLK24ngypoBgxQwDVI
qcGCtn1KUf3s5MV47F2WDa47FhL4IPdBDMWYj4I9fH1A1D/YGXWdE7TrfUrCCJNUALFxP1ZWW3Cj
BggWg0DshrzHbmE01k+5EQJQ0uD4bygpb4mjNyliSBC8JTtsMl9I/rUZdT5eCsmXoJQ/W6LpZnAl
jrzVKO+kadWfNXaHF4dLBDgkirpx4tPEtqguXMSaLpuydJVV0unyG3ex62DiI7l/h7ZIg2CdzkKw
oIkKXUhpyvKjwyPK5SOOOSxOgl5IaAY3QjVIV4yr29t1U66ndxgM4vc1dqshvJow2wr5I//JN5np
bKkC0g7MLy5HBOhkqES6RX5eK+SPHCT25P0TmXyarJE3FFoJvmbPq0qXEEumRf8A8jFkLBsz1t5q
IS+0NSgMWXaOHStZAilTbEWSvQjn2vLEv4Vy1zpYtf6POPGJ+hp+hen+tcxO2a4Ob3NmD6cAR3nV
BRhQ3B4Xd/4v4sZiQQz4A+euRI2vpRFvorvkrlvKRnEA7BNjK1ZO8TUBGXDwAqPaDNX9qSIxRWSU
u6V+xbXf5dtEgHN3pWdFzPgb306iN2J7zTMFrcEyTF7f8yWLmQmHV0/T2n/UfXHdjSeY15V2q06Q
urAhLrB19IJaaQjSXuLf3CkD+o4TC8qtae4HnRUclBOIkfhdw3nyTC4hLn0tXrxsCMNJY4m7vJog
MJgqiGyHlkOwUr/480FcPHeX+GC/qg/9ibSdYvG6o8nb0GK8Hp6uXUGz5cuQmGNLwFZ6Vq1EleRl
QIlarKXFMYQ1xZ9zEyQKgr4vZR96+HciDMONKd1zF55KejhdNm30AmhnY5D9P45/WeKVEx2vkS09
fjFRgKxryVfPY7jtHzb4vc0TQdGwBg/cXu+H0zQxAYtnMmOm8WZJgKPgIkaevJRFPfJ1mBNl67T5
pPzIXONsVdbWsWwP0c/6Tx4D22TqxARm050tGnaLnpgPPqKxt7gBV9HflSlsfrijFbQPUgHu4UFw
FxWEiTfhvqXZryVcSXBdnYi54aKkv/MgvU4JQKvsnJqOqR+GmP4pH5uz8+sDvip/8oQ2EwmzX/B/
zbifL7apoPfYE/LV8QrPqZYPkHN5jLfJ8Ig9aSux03vr2tmsey1t5O6YUVLzUfl69mt42mhfTUkA
+C/8StBKVYsHN478xQesvfCoV0zkWRinyUGxlbj+qe9u/bwM0QaraMJq4qeaVduI+4TiP7lb+jhO
k+ZUwzSnUPDtlMY+taxpmbStwJzSx0pIEqYSAmmExWiOxe7+3AESh1bv+Yl7d+rHqZeRQZukHTNi
Bmeize1UOhxXoVcyRl7lOv/Yter3oP7tQiAbhhPQR7hIhWDqmalAvULegmHaiyqLF1KizsZZPsBr
TO5243JuPvcPF7cbt8M2F8w/eXwHKFjk2g3G3aiAYGdbcRxmzvSsn+K/Ogfxg7LFyenCCzTgwzvq
65dpQ46UOnrIrNqKYgIpaL9WhJKmB9H8NtYzucHBz7L8tKWY+SBumWRytJKrGBb7gRTkojGeefT2
cq4XaABfqUATtmBsV5zE7r7LX6Il0j9OL0kFPIycgEN57zeteCtnwX5I+Q2r9s4W0n7ygK7C0QCb
YRZBHqxOZ3yKEMuOlk1zEPnUYNnGyuT5Ur5YI5jYxiQ7nP2/3uicPe663c0qXmztHKVvSt0zWPym
d/7MvHCh7AEZnWKl6czwffeMMKTq3uja2ln8Cgp9eqv3OYMlEHjxq0YOa/dTmMH9siLpTBH4o0aD
fzgzbBtLlbzIvEhahe7/2Jyp6OwffSipX3ZSuDf97VMVr8+8vKi4j4D/pNGRLCJxURuyymhR+N3n
Ox/yLLaj8+Lm95f12CiRfkTGUEdQVwG9XuBz+iPdxs4JYRSVWyCOrcgDnQzV0R12Mm/PUVqBwxNW
IIGO55GYEbcmlc9T2fyhSQ4rJq1F31KLpT1wS0PsXWku7HHehCR1a8ujicv11u0GtHT3Nne0+STV
rr+nHN1u59EnpZDyEKCl8jTteoDwcryZeDs0kanRHcK4vJ4rlgi+r+xcMRfXT/krnsVWb5BCs7of
vEukE4OsYcX+HT6qlfrNkqAHt8xNf7XqlMyG6h2JGn/gBnFXYFtOXWNYNa5x8nLN5xqG9VR8y3wO
VMimAjoxyaNKithf9ntnMiJvjuSmpiL2N1yuu/K7wZEGLe4Zsw7dH5BXdGlrmtFYZnO3ZlBWy/+d
tqOBox/TTwOehjIRdy+TuhxC2dDSBAkoW7+NbXa5AfS5SHZhuqDiPIUJKqxFgSqjGntLTAgQY/2g
Gig6q9L2NacQ0MgA/nS6xq0o+8GusrFXBS5hE/cMuFCo/w2avuPJhvO37ELMSa0cXOizTZaiivgT
vZgs3Fj68ekXkSI23qhjoIVXUUASMWjwrtd79Rp2JZpkp2BowMq8Xj12b7fRp5z8ivL0NnEbxGUr
k+84llugAIR2U7RAkI65kfj8DNYT74OV6YNvPmS7tTJb/mpFxV7etXcG6cimcPMqGtTeYoEqAdJs
sRY12M4bSlpd43io/S/QXhsFbxb+o565lWM3IprZuXIGfS5CQmXuJgHQZQtVfcQ6g1+W8q2rCMB4
skYSRSe3RbcQL0bBFfcpcsb0CJGrVOpuuFVVZKMtQIUg1EHJTroOVCRqNpW+/xkfn43Uo7EsUppQ
7r0s3x63fneIbuXGCveHhOY3m/ikreNaki+2DaNaXpb13lcCYnlZp6s0DNTTvE5ZakE3VGSTQg5U
lVuMI8MMPlCwhQtkef4m28YwtfeK2QF7YaexqhPBv5m5elJ2bGvZjGA11wtx9IJTtqcc7DAADmyd
ADmigk3+8iaK+vAqdKB3R75mt6oxZMPq2XoMZ1RXHAMqJP1KaQD8bAjE16FWLmso0fX3IlY6WFbM
RayGmvq/glBk3H673wheVoUukIX72AJkbbuoTBMLPhKKDdxlt1x1YZJgLxMUSD2/ZAVB22W5BX0w
8E1iGYMlJWuRAT3CRd35gn+T3Rew5qDjvg9YOrAQvozzkhx0+cqhTVVTCJGrTxmBWyKJa5wiL9pl
0kwFrwvIqHKrq9d9YROiOXu5zdknyyJ4uAtYCjrQOdrEV1byYhwp4G6v2RfWnXmUztsXeQeweVEg
gfCt5waQg9GqTTLCNidxmOSnGzqMMMRTnAF/f673CpIDxc2+F/JXon1a28t0gqkZZ9jQag++qe+f
spGWHm+H+1QN6hX3923YuXOKWM4oxkvFkYgWdOvjUjR8KiHwka7xNv9F1P7yFNk1hsZQSBXHB/of
/utukiTFZin4Hhv4UST8z2osTEKuSaXRHMYw2L6w35L8MAKZ8JxDvBfafE7S+3UI3s4Fwp7E8+T4
G1GoB3XGBGM4+QV3fHm6vXiZHJG1zLOyP89ZZx91W3XO0GEXaIAHMkCms/L0BYEvQvD46A0H2VX6
Kua6epnHcYO51HtJTGshjSLQyTwDydkh2PMSjXp1oJA6ENDbPRxZYJGtMsHZKaT39PKs9zEWac2e
kE9el19OCCxzROWnGOmfx/Ut+BoXnKH6GKXOzPpwzMcFDOYIV2g9FpYDPDJsEmeuMOb+Hg1Ap4B2
Ie57BfVcCmbFYbQDPktclQKshF4+N3byFWNQm2TaZVZibwTltrpCSDkyQ41lBBRQtGngvBGV9vPg
nIaIflpkbBxinlGhpB8CvMA8U0z03E3PI3GIdkLr1445PZg9yy97mW4Yd7lCVMAgYUK/x6Ho2eAK
NyjhC+ZAaswIDD+iQ2MlRUIncNFzr8ody7EV8UAUlnYFDYoQm1z+XT/E5d6El0SIEGe6eVSQ2+2q
s5M5P9Ys4VEP8rB5S3VZGXxkaxdfngfmPNkV0mqoMEPFshsGs5wdZtYMqNFG28Mf7Fp6zJzyh/Ns
U7kPzASuUhVumDGqaltO1UnnqH81HFz0k9bFh2p0zj88jwln+/uHvsBETSuecHuU28PPb8pRWjLU
UGYSiHqwffh7t329tm46Qi2/E8UDv4Ei9fFJrX3Yfgqv/5xt9nKZ48Xgx/ahd891hh54keHrGXVR
DTsAddWhaMUYohYTpeudphbpe7REXFQ1nZpsCJTxBnBJd/36FM8W2ZiE3U5pV6AdHZyQyMw2Mijh
2mCTsXGmTiXoBGiC1yd/7tx90Ev4pK651DmzVnz4folbQgkuDbeYcqXEtke1tulqKAQ1M9xl76SZ
1ndyYLUyf6ni19HIZWO21Q44jdHuQTWLOBceDBBbxgR6r0G0un51Phww0t+cWwRbXcW2H6VISl9y
nCxqNm4VR7ogfY6JeegokfhmvY2MG9xclR9DqcqDSLRSpucF8ixio4VPUwiqUoEOVE+MekPQr9Fg
3W0GIHIs+m0kWEc8EhntEfZvD/BQvQapF0S4bxc/HMxDmR1AiaFDrzLprZaXf2VCFujxtudiWvf3
rnLTS8YXRXxmAwYD5WMNZGEhFTb9jiUZtKdUaG2BzmbrygDlSsgViLf+GMNgwueLpr5jPfHuWqIY
hRmGA7EkrxkNY/mpFkLt3WkY7YqsDsh5tz4QOj8LiBfNJB7bdBhlXG3A0wCGmDuZZflNxKDu6T6A
VbENQBfeh8pb1rLXNKeej2gUjRyHpsMLNsQgGltKOHPDAnQCCxwuI0TPVmZzOpgHxpVgRGW/pkAF
J4Q6z4KBs94w77w7kQfVEJqTV7GQMupLxBw47VSNU99HEFgzs++qxkmnXyEnjsGnZt+WPBBvNjf1
IQb8bD9xlVh79aV+5pmJzuu5IMj02D03/tLyKtU9spNdK1T576Ey84fDhP+lGcfDIyASnT6ZXysG
7gtcLj3COSHKfEdfMKA+DoPZxAK+U0m8YyS0SLTVAgSZMCJgi85CQ7hfWtbuzJ1YWpcP/90KHmqQ
Y1ZWkbLMa9Myf9jWYoraUZIcwR4vnu4uTIXMmM5XJKc2mAYDcWoWeZxOHHz2yXl0S7Hx3qqDb/OO
F8CI0e3bYQAXusj+hN3sNVREnvjRypy+xIAPKCKA7ursvKWqx5DWr1So3hrX5STfW12azGGGyolX
pCnT9jnJhm5a8aqAMkVZAwWOWuB9Ia0EEpxwNVLvtzfT8Hy+EUG7KB9AMe2/h992HAUEvPAF2VJo
aGiJV/T2D7aD27KT0mSeFJxdkS++wrQnryrR3MxkWe+1z0C63UOqXlf6XeniSKCdKwWWXG5csmhL
pXovQCoj67lssRqoGRY3U4j4cfW8R+XfIeKttYqPJVlyfOG3kgpEZZrGt0QGF5k8N+BTKSw6i1xS
zU1sqjkTKtZgZO74wtErkx8grszj9oSTAD5iggOb85/6pxs7jor4EvLuZ0dkmdzNZXdRW+DMcpd4
BdDpzN0fH9iL0SJvYk+0mXxEPYEpuC2RV1oT5iFo8yMKOuO37xykAIWeKzKYxJK5CWp01Y0A+F+s
oyvST8MbnX+wK4GYq6s2oq+KdWnxyGtQiof982GFv/clx1lCika3IdueihUwZhSslJEvjCFWL4OP
HOHdXiS9Aq6Od9DUC8EvVccjUuoUgnKDgRNZ/8cBkvA610ptUbExzbfuoLzKg0xiL7LKBndRR8ws
DE7XK9uROe3E3cf1foKpJfW/KF8Bk5yV64hNeyXFPG/8XmFwKwbYgQ2ZP2HX7OgXK/a29B8s9yrs
KKpo+lEnm0aGQgDnEh2xkGNbzE1PBgQKsUfh8vSKIhf1zRQqoPU3IqPow9gz2RW2Tj2288HbwZYz
GRnv2sLm3OrBw8hGzVhQHNT00BTwnzTc4hgoA7UBskHPDsZsx5wb7lfLmGvxBHKLRPnYf668KMbY
KCBVaonzQtFIHAqZTRZjILf9l3YHuSDM3ik+LXTyyDHjWIiowuZ9IXmOQirXUIyfOTkWrMqND0VF
FZFZ24UCvJ749bguoHscRvbvx+Wy4KOki/FV53+gWbyyYo4ycmb+PkHCm1jQfmZd3do30pZd/Fse
gxkYmQtSnJZzBNwGsJWQ+BHE0EaD8d7TvLZgm4OQ+hwXok7FogCT6ot5LCOVGn4YSctc+vaVS9ZC
pCZYZ5XwTouL+by43Uog2Rx3dqOyBudX5SG5xmT4SlXGhaLAkviLw9XtaZ5IaQWsoMtGsT1mnYfo
qGedAw69eccxBjrIJprWhSve9KjtWCnbl5m0QH/Tee+7oRvm257zVClvc+ZKvhaXu4MD5FKxM/2X
ya3/MQytUxnS30BdYQsy1+6zUN/63MQbXnF1PgH83nlaLNbOWWBhMpflFSJ+DaWm0THg1adbtZCe
4wHcUJIFTvQCUeqgXwo+lx16Fv0h8xDt5M+u8c1ztRQosRKdHGVQlqelqZn1H1tzfWemVvYc6BIh
dfPQ6ISJdejy1eODIvC3QI87uyJuTVvtx7s4mVg4/oUexXfyfwkGf80bzsz/uE7ma4pmQbWoyLJr
jzzMq+k89YCxZUZIVWrG8IfcE9KLFPw1hloHztj6IeRtzSs4rPKF+IxvSBTVjoCXzper1wa6CNeG
GuscHuMa7ah+GoLorf+lwgZziJU1484UvOMczTsL6iXpfODvyCYI9NOIn8Feqx4JsDzfi9qqGUb1
j8KbkHBQF9k4d+KRfPM1cur0GxTAJzAEHIICUXA9Frr2GJYKbJ4H6BANW3LgORJJ0b+Ksij+pPiA
rjUB78bP39XaOmIjeClXpeJTXiNAHFfKOxo04RAF3jCYIy0WvrAdX6makHRXX+hpkrB03BU3ipjo
H5KgoU6huVPOyZ6nNDEbWwjidFOx6kOLc3rONRsBqHOWYuNKF5jX0IN0VJ9hucq+Wj6LZK4AZ0RC
Y4JgRb8JC9i/F7cPb8XX7mjZmDvmejPz9kwQrLiQ63NP6XnsODCTK0KGXyAyz0NTyRiFXpSVeR97
UFfhyVttHiDSOcodCGsxgsAqscObVxnH/S0njok5OzENvtiTiieYsUzlAVRncs6vSBTuL5G9G7xn
nTjVeEwJGzfvoatVe2FFMhUX5R7jP3FIdtdQ7gx5nzglQYeV+jBJB/+hdlklxCOBsLeNPXs+dmMM
pngxDMwo5oY/0eR1KVluH2Poh6K/Kp8Z35XZqyWf+lOzz/ncchwtNEp5wWYpfeoAO+cZTeikiBa+
5R3maF6pb1gfNnCvAjmWJ+xLWjeeAiKR8xdn4M5dE84d4yViFHvwn2iSuHWVsfXkXs14S6EYE9mj
/dKZ9ZhZe8XsAKYW0/icrRnOoUUcYg6Tu3C1crqsnsMtWiejUMn5VDDAXDcvPQq/Kg6pP/MDA53T
QbAVXAdbvruTZn7b3oParYNXFemPcgdIYQmyvIYT4fzxXbplAzc4cRLnPeSgcg3nBrG4wkjZIRCP
a4zer59Nbca2X92SxkrwEAeU8PKe9BdKaNs0Cu0jAjS/mxn0PqC4eh3XHvtGWzlYNyaH7+jylzAb
vabpKRs2oOS05a2FQrkdCO8882YPdqxsfJZsnql9gIhvnfGOc9bl4EU137sWTdWbnfONanB1Joru
JNAuIHKcSodcZbEw5KA2LXTfmq6JNVk1OW5tzy+Zp5yj0d1S0G2haoDkVzKfyOURLkIFC8dzQQ6y
AwhFDnJ6hV20SYaXMpyEmhCUVEPgxAMix7p1CuHCxURh+439SX7Bj5Mc3H0EdJmSYpTHljLXkjCj
NTlmdSMj7sZWP6Gx6sf/9Befao4EsMRaMbQ+r0Ddsq2KWsln3vcXlX2tymCKRxl9UHZS9LX8FNAQ
pa8yOSwMWAypG6oIH6a0p9EQmmv5qfSYz5ClikbGMiQAmGDJEjPL/LL1BszVZ8vRX/O7NW4Wyxwa
+GMuYivETf4qdskgr+4AbYXtEu715l/soCk9NGNEKselRbqekCeWlZmrEKm5uFT62v/qu+lru0++
tv6bk5KQ6QqR9NvIp5RrN88HoBUoYfTUE0Pkilv9pSb75MTjGTnxa1ewBFD2coH8IgZGq2sdWIgq
y6q1lmZmjrldAbGmmVLc+abDGGLBigl2dhpvpiPJG1Z4o4YTDf7P0v6nRA3GjfrnO2OyEpaRqnuC
lylvBUjJRbGicaQu8UtaN1Dvrt27x5IMefQJmUEc8qEu3I3g0yDNKNd7gAEmyoXvKSXyZZRPDUJz
TOeQ4B3aFHRgVxFucOzZs5pOS8QO30I1hh7fJssYxACAf2x5bx/f8TIS/4LAw92y+tNAWedzFLWh
Ka+6mUOLXnva+hWHgEpTc+idFHHvkbgpfn0uCon+Uft8UT68Z74BUT+VzDArJoCnr1A5OtmOXvjP
Sj3Wn09dBl7s/zQrypgJU8mb8Fcb89qyC0nc+wPWYJ3PH1BmwacTzqlpDPB4IJPuC5H6/1D4jUDU
c4wpKfUJtzoE4fg4/TQpMFcCFNOutA5kxQPfoft9cX0r/M2X4FZeI2hR6WWNLaLqZ+ua5UuExBzH
r1y+GW/Kv1+wZRGEUKE4u7NBQsVkf9IQZhqxs5Mlai5Qp9sNiFHmndfwhdx4dXYt72VdDchTWh6e
0WICiVhoFqGe5/7hRjZ1wQjKwvwL9E3AD0PaQOY3oNqomH1fShARCF4QqO1ZF3NuGyHJW/TxKlO/
YviD3GERk9MfjavYpOZN2SisAS8nLgbYQyu+s7fcnseVRSQ3JH3hSC4e9Wq3OPafh7koaOXKZKqk
7518y8ueLYWvO9ZLdAMdWhdFyF3ZIeaVUtQVwe4GH1srUFurH1V3KC04nK12Maeyfl9E2wKtKkb5
C0segIYgw1x7h/DR1igRNKcGpv0VChjM5oFKZ3sl+pIi+SDg/w1tPnuBFTzgmIGT0JJEj/B4nuxN
WjQdewgyhB4H1l3ZbW3DTViAJf9Vr9N6Us6i3EA0TRUArJrbaUIvWTicLZlsU1i+OTNKuHPHyB/9
D/N/NV7XYerKkyI7HcuvpF7sXFrKFyXy2Cg0c8b0T5Jwa1SnEhN0V/FzumvvyaroLxbPGvNzwgDl
8/nYr7feErLy9NATXmShxPZ+mjddtJwZUWVEhYpAjdZBJjrDFpPYzYDX3BB7qL62Fz0YN49pZz9Y
0S+nQCxyUvW2chtdztSOcHvgqzOAzPDRe8r1ZAe+lrE33FXuw9ylx0hX/aSKZd+NWCBmJVjApH6F
t7Q/aJ5qvhNWIutT4dLCtTeFx6jQMttbmlfTy7SEZuXH1lDPFydLVC7cJaQSBRFBOqOEJdLgwnjG
3wKtm/qNvNBmx77AxjOHKjDGHKsrksjpzGmglVaf7B31wwMDA0MulbDWSGqD5Pq7Qqkn6f+GhuB+
dkJHZJp0qRjRgrc72j5Ob/B/uq7Y0eEdStmixMZi5sfJEQs4QRSIccoaZl08IWdKYj2Md8l7CuRc
R6tVyrmBL/O8ssM8FOLwXC7vgGfanRcLWGTNLgTnDwzkCfr61Jy3ZPJzZW9YgfN0uxW3mqazEqXc
nZ8Uy9UCoCLY+33pT6HnOguFbRsv+gSHSqiJAq5hP08NP3uH1Tup1ilbXpaLHTeTd5ig321kjc0u
LaqqvDyUxIzBJR4nCdRgWyEdzV9Vn1lWAjPdTFLDmf6O36gZLWDvZv+yPJRXW/8wamRQK4e+rMhB
+akgZZ1PkvnUCpHsaw0Ep3pt4B6FYORffjuKhIzfeMQ8WGVu4rgn/doyZ5TVqvbMgKvt/Y24vToR
eCNhEeQ7y5oo/Amn0Q7kPxMgOziAn9f0/XzaZkDEyCAeq+vjXX5ClinNinsucKn4hmrSRviiRGGw
B1Tu8BtZRmGdxR0Q5Sl4a3EUCCd+EKxl2pVNPaZ9CYP9QmFwUElAyFQJVBGJB7KSTCXW7Sqen+yh
nLSMYzWeYkmrVUoqXm0+8oktUSR8Kg6U8It0WMVMN1otucGNBcBr3dS04NnBProfsJ4YB6GyW2Mb
4ChqoMabWLU73LpS0GY3ENKo0Hrz7W1FQle5NTpYUFnJ+lRfNo1SCrA3kHsZHPvc6AYTVIIfOFIi
XC4QxEyjzUMcsWLRGy5MQsU6gJcZ4jTTg8kfGvfAgomx2KIao/KiG/2t+TMTGgFO4VpvsJfYz6DT
c1upLyjEUNM0W2y5+GjvHQrYsUAj9UG936tDZ1YUUtqfzL5V0nrmXKwcG4x8koiesETJPr00rsyI
RewhpJReH8onXktlUhTOMfmBUZnKnS+50kIAjPNp9izzWwXTF1ofWjJ8BPCFDrrXeqp5fyDgsY1c
9EBOrSAYW0A8giNHQoP0OG0n4wMwjn42pvjkMxfa9ZvJAkS9Yvd863sa8xdVFkyRqGgjaFPRtxEn
IGMIOWVXA9hOHwGqRXKfIfJhW9zn4aheJMYN7LDU/DGWItMd4k+6K9BQyr7mYXbXB4z7xgWZjTeg
BW7osPn0Km1qDVWek1ACx/HNR3LYMVGo+Ebkv/d5/gp++lyk5pZ2tuXOvA9vuTctlYA9GnzHdKpw
hD6jw987W0lo3PBNuNbeiqY1akVraeGWs123qR86pqr8FHYW3ispLI+h65cOMpzJzYO+SU2lU5+I
BIXFAR7Db4z5JenSX55vyWaHPtifTHfpAyIdhydXh1bzMguW5NESrtH3B8d82kPFAiHyfbPFN2wv
Jg8Cku23vonNP3IaCnC2QbMnYu6TtP0QkY8G2avOwTRp761/PjANB+uKID69y8rt3O2rB7e9l7kH
W4AA3gHsPaFQ1VuObiTC4WvmX5SvGwC01j87KcDm8TlYkVwyr2EoqFsATy7PASGl1hSrLB1EA3/b
n9Xu9QpcYf6iWilo3985mScgDEWZAe+M7K9BNi4mDcrGVkNMeYXM++wwkEsim5ULB0rIZj0CowQ8
dEW+ZJL1II2IoJM2IPxwMn6phA0/Xx3J9k8nAi76lVu21nROeh1rl9l4HyPCa7T5dVSmfOkVbf/d
H9mxor/i8XgQ12GuVC5eyDtUNkRJx46vN8tVzK3H3335xNOBTSSoaQR5T/WDQC1Fv0LEupqoMt2S
KlMtWAF0PeQ67VbFmZWnoFBMLLWjRRDHEMoVLrJdvlOxB6wNFZla/J0ItI54AW09iJAWzu6mMQRy
S4DwzaMPmsqrfnuAvSY7bzNJtaBhJThfGuEFpilcFbPNXKD6uyKtkDY6C/yuj/HxWa/bdNzr7c8+
BkuARuXA0bn4xk19up3RKczUC9mOYIvBKAYzrknwnUF6gz5Ba6CIfOulraplQBGG+y3D82C5r0QV
yoT3l/j6Jmwi9lqnfLTdq46s6mbxaRu5mfMT9xWqyo4BLWyhOjv7Ey27Spkzh5zbU5cv6p9INBsK
A7zuhvyUPFn7IuVl1DVCNHMZqW9p+24ZjrHYuvR7wmCyiMJAe38WdYuBAgK3zNptDYX+cNvA+p7k
HpfYz91aDGMzJ9iHeGUG5WLgLgx981X5eIBLU5kiahaIqHvmD7eGRn+uqgT7P4c1HbJMqCWtCEvm
345Fub4fC86WkfEVLgPlaKXm4jeXd9xTr31tsPpTx+cqn21TFFLmFUQTUcmOQUqLM0gClgcWUVeg
PuvxmHpnpeanYj+PF6OL6fqven41CwKr5O96Qe/AZTffH00BcodjZ7CQGkCGHVCl3XdMonMOTlYS
JNVijvWaA2RB6CrXqrJMdmZVYp30u5gg1GeS9tJSNJJgSoLWzx8BAFg8deNZ8NPMYMf7ikPfPtKe
QtkmrXBKAnJYFpNjkt+LIwNH9uuqDpT+9ImfrjxBG/4POHJd64ypKqIBQe9iRy/dpW7mO1yFuqhF
ETsVFnTkbPY0+Zsu9ckKDLYVCWNNrZvGzh7JImGv/BBdE4Fayf4Ab5AGrAVLK44Kg2b1H1Mw14kF
X2GpVqJOPCf+Pv/D06cWZK0KcDtodo1AQh5un+xbJQfo1DaweyWw5QOAQVo9rO9a+R6OCJ8Hv7qh
H2CThHIOS27gT7khaWoKDpRZccNpwiiXo0zqpeQnlFTCRnp+n5LwxeKggBz/zGrlGC5uQQs1YKDJ
KI0iKqNlXKAF96cT8miDb4cQaeKY5NE1bW42pgQsWbAnD4vmINgF1g9C0LaPqiwTiJHy+QZHVVMA
xdQ9Q6sIHReBhXc1OQLaZG/uVNkcFXAmxQN4KghSSPv7KASj6qpc6Q48w69DzAampwBVMN4vGNhF
9fM9+s0209rm7Ye/18JnIY8LbnQa2cjfD2kgbnTjIqFH8fPLekmcQe3AVmCr6yQRHAhj4iieW+N6
vf2Qchm471sAbP4bBZCQxlDbgR4kTnjUlcLi5h4hOBnUU1DWID3AyT5OzPhQKmm8nLeUWRITE9Bu
6O6VD2vYBPFknj9eTJ+Bw2kwyUnXcbT2olUGERYIn3kr8AVPq6JGISjjQaIYgA7APHRvKtihdM7Y
bn7z5enLugenez+82pLKX5NBd0MOdTrgV90HwpWvBWNNx07qSg2z6jNLCnsOczRaOFvipIU3D4U9
3JsphrjcV9myO3uQvOpuMHtQ50MAp6PLyDUBoPtWxxGe5INdXp5z40nlT2Yfny3ik8zQyQbUtXqz
1L31oVQ/c9jOOaauaPzlRBaocQ6kpAG4NR6iEP6DB9CZrZXSUWOjAkLt64PwL9JdRKPN6Z6nGTTC
GhaIjoJA3PklN3IVpNaYwZuUC6NPSNQvGtc81QCPgV2usYUp9x6lnS+XTH+MuNdYrwBjHvoXzY6a
4rdfCcrX9+FFVMrBpKzSVQFATRkzxKdgxHjNtuRgp9jV8MydAxxgM6h7/OqCUPH9z6J6/wMeGeLZ
A0VAAtKBRlwZEACpJY7fTboROuWoqwUVd3my/7vflIceH2uROxZt5WZhsJIoMjCL7GkruCHwUzMB
TgiY0evFZsElQSKBW0VOdD5lXG3blWSB76gDEQQ/sR3Ndig50yDS1N5x1w7RwavJfr9RZrO7PbDQ
PLfIbWpGU06ARcB28kbnSFoedJULzbW2Mwlrnq8WBRNAb0+1WOP3KZrf4nsUe873XrH5z4N12Alo
q5tzISRT33nYVo8TBfTcQ+IKeKH2gLWtFjoJNxHLAVMO/FjcI5LcVT0YwLVtt90BEPD+e4ycun7y
ACeW42vbAygo0f2myiH/Iabdd7XS03sHiiXBY/6jJSwlcLqwBKWMr0ztKL2xyLkH4CBNJVR1sOGn
3M8jAlSjYZ75zEWLDCtYuRnWtvoie31h6YDwNOg4pCxwFKeTpl4XS00+W1+L4uGA2tnC7Yai/NrW
ztbA8qxKK25GTBv4lctnaH5SRQMnab6PtQ5yDKLo+TCVvcipWpPFMcgLocCt5QCvGHP+TxGtSehf
tYa6YZhdCuwtal3c/kpYizVyUkcFqxX+20fa0lWNuIgvfn4WQFhIxprmkVhEEMKO6pACKBbNq3w3
ItvqB+ezK/pzYSIIt7fyNCNBoaKdeem6XJ0cyTVtv6TMmRtbK1BjAZBXNrWwZVSf9NOD9UnbYQep
oIXPsEC4KjpfaYHx3K24pfDX6Oj5LY3+XG+w8cUpcJBVZjhAuCztN7nDY7vEROmP7hVXkeXVXW2m
aGapZ2HAWiGyXmi6XoYJly8vZo+ZS7B7scnMLwOBHB3/AoV0IoNV6pwRZHv9E+7kxGO+Phds2vLQ
EO531+mCp/VWb5nZJbRvTf8Oj226bZmYHSnZ+fxhl8j5vHWh0HbWi8R7GR+V905TesRMe0NmUTxI
lNzCrN9gGqSoL5dMqMnTEitaHoqbB3+Pb5zoLO11s6W1hU45k6vTZSvVtqPm+cQ7UswKKzAlCkxJ
yhBExBVyhQM6k1vJ6xPU5z5ghHXHpixx8Dh2lkkA2vMf9H/tNVq1ouLvpDXalR5JGu7PuzlVcSiH
KUk63g3YfS+/CAfG0v3EJbg42NC555HSjCGISL624MuHMFQXmivXi8YG6glZhcy6ienuWobYIn+o
87yR1eRfbX2ds13UxjE6ohrlKmJlZawZbnZCUOla0kDR9iQMrLRDZ3ZWMqrbAyvfTgy2HNFGdcgq
l05D0gRktaxOFT2/Z7lURGGKD59YLtmPrV2+G27fc9b57t8up9ta0nmae0xU9C3RFfOLUh7kdEEY
zksnAg+QElag88T1d/I67SY+czEcznfUHUJP2Qwev5XzS76zxK0NdNoCUOGSzU2QiNNGuLwfhjRl
4309yH26E8O9oDZffPH4C2qP8hRehZbqQirPMJxoQZd0b8R/i7AuKsyC0zoUaEv37W7h+jGvsrlF
zpLw+TWvRoW7EyOTJEn1tgBkUyBwgJYh2C31ZbJ2hRU9IqEZUNEgeOIfa6AD6vC5rdHVX9tJmaYq
szyf2FcoExArlHOWKU7Egi/qconWJ+ASMkAPfnbmuF7gDrV86f9K1iFHIB0k9AoBZgqprPN+GFqI
rH24+nQlMSYFm5AslB38Axoe/mtN6LbAhXMpymEggGdZs0A3aoJ91nGpBF9/G+sjz0UiZ6Z2VeMk
Q4QcabQ1/cUGJJVMXU9Nftf+wSIps0HJidoo41kVzF2Fj3z+YNnMXBfh39HaDNtSMZRBIXkxrjMF
8T5NtBLA0O7lLNc/f8xkP6BiGl1r98yFP6OPlOGNXXk8WGGPi/taHl7U9Fy8Z2pdh97ddCUF/jT+
xYiivSJDkgaqUTBWnLtaV3Tw9W1iM24lnANBKJCiCcmxV6UrHx2FLwDROAvy9rha0qTTZ3WRgQt9
k6pHzWk31GVLxXxNKg1IMs3QhEnfeQuK1kZpts67DHtCL+P2kqSNX6AzhzHqrMmXUVqZzb+ASH2l
pKo6VeGDgxmG1d5FQCOX/bFKrAYqRf//4Jh+sqok+la+XxVaLW1wvh1Nhk0dMYOGZo2EqzUAFKdd
8K7JGl3QPNx4UTMcYc3y1Q+SwDFzN2zgc0fpBB3kqoUdWegFXOWEVjPz5EwFKTU3huRTvHbgmPZ8
cuIH0QvFdjD0W8C0x6AggsQRGXJqVUSQX9tJ8FymPR6OEXX3Eo8o2nEc5pjq76FAE3k23hjCWm0/
zTFHHz9Knz8xyg1hI/4f7LYus9D8t/FWPu5yhT5oA2tUCohi+fBLh5QUfemiIuM26pd1b4uf4UTr
unPOoA84id2Jkr1Ibz7YY66y2gh+IRqPVBsSN5/PpeZCNBGt2fSqr/6B9WCdTSkHlGT2J3M1Y1nL
GZpVZgTL1qxWB2XNGYC5W5lAn3ADbYUS3qCScX++1JeU1BaU/AHxd1/nOjMtiabl/4/FlCEUGSvX
iYcbu/eLojWhE5MWOitPqfR4wpTVDOhbPI8vbX9RSAwSPFiVZVbf1xer5fQhjjF6/ABKNhgtUVqr
agZwoVHB2OoGLDpnRPEe6baewTFFTFn+Hzg9BiPTTg0vmJOFUK33Baws5zbjL/PsxyyLESbA/qeH
BBP56MLMyb5VFpMgJVZf2ZCOrxpnC5gkcpY0zCKaMSQJAeqBM49Mq8zO2y2Yt93tbIv1YL4QBztI
qtkrsswh55XlmCgYHHx2oBaQ917Bv+Cuvb8HzLxtSajdRHFX86pyzFtuxnxmQbdcsyE42rw0Y/uc
v89pSft4HyEQdu+gNGiy9LfDSGdh+B0OJiu1nmfBEv8TE624SM0Dh9MwojNnzpjtekLwwn19QQnD
A/fOEOsoUwi0Ft1GXxw31+uaRHLQ2dukO1zoXCAGzcsXwxNcrfPrsll7SiK0pIka7VpHAnpmI445
zSlJnoelF0WuWyC3Wf0ssJLPZPzWgJ875czkQKj5nTVZ2S/lPMqBFtha3wPGd9C/qZ8bwU6WjMZ+
tUreCPH29xZtQsLalIK1JVlnIwBbR9hp0WdAeO0R7ufOeGlbLCXD0rxk+0L1IlfaiecDJiz0vIOU
Dk+non6z+n+P8GtezC9tp/Im6B9MgvwmzYy6AxBdHPe2MpdP1rqszwojSopqSLKUVnndWcb9ibPa
+T+ehhCBSnMYn8Pk9wSq8ZzFrwnQ64UA9Er5yD/b2QX//cnw1Lo9N6ti9r+UWXskNzxwV0xBrDfJ
2I1e/FGtLG0aMFKc6ute5WqguRhBIskb/BDlmHmzK+ioeNkLvPtzs0Cyws2meH/nX7vuJOZ5EV6Y
7M6Rn1CRPKHTIbknJADl66526jgzWo7ZxWS6YFV/AI0gOYzE4GKTPWZ7+ScC2/MsbgvdpYNxM5Ph
m7+Sa3gn2LrprDReuh7QgZZT6b5UQxRmF5gxe+jxnTyK3HDgjWNrMOgGOJiL6ddnMyAUfzWAEkNK
u9XOSRx9nxfb7eeXr00PJw19CCVeBRAKItweUg+bv9KKZ5UX3hZ52Akstz6QTwOxZDkhkwHbiUly
d1CbwtZlvqszmWUerV+zdViu5DXAH30/9fM6XWokAHcaPj0rM1oKNkPHJ1cpWSc7D4imFcfAs+fp
IbXHhZiJg/2ZRzOkGsHsHrKiTYG/JMEeviaFV0A79NOHqfVVM/sFayS/DPShsj7AdWwlqHanDSGy
FLqs+pyMBjA6v1M1x0M3H82Fh4Y9h9TelzNyu5QuOB4PTSHmYTnxLDLsbR7OBhayJ6bkZ/gTGqN3
93cpT+uDOqQKjcZsu1B3iy5jQcd7LNf1ROFYQH1U1apAbEOOaYhrPEsxqms+sQB8TP0Cis5dM476
GQeq9DiJmUI4rU4UhqBB+tn6Ie9FGxV7eVwCItalkUluSNLdiBc2J0r6/3nb418r2/Ee3t9GOxCm
I/VUfcANE1xd+JfuK0rfSWR7iCd1So1mRV2n5haiByw9ey0MSFDkrrgh5E1SizaXu7csfSp3uuY5
ajyoKMmfeNYU2eefMPJ0QqeEO8LBICS+sqB02ngVpnaZlLb3Q0Twa+XBagcoEriLBqxP23o2gqIC
8fh/s2YNOIKvgdtiIwPiY8ZIGrGz/JsZyZ/CxLhEduF+EnTK2L8RQGKHY+B7QTzYZ52jzzrYyxT6
lCStnZwzO2W79F2iyXpJenIKbIBjo1elV6qQHxBfTOB/CUNJ03f+a97yk89UP2XcJq7BeoYioBK6
YRXrYwxV4wb9eG0VtIXtnMXtCeBYqPwv6kaRZgnXDs+gojRUVc4bYSDpypu+TWGiHwVfMG7fpfIF
pwpQiPC/8RKfWE4TV+mu29u+GanJFNr9DHJmqarZMvT8QsIpyGEErIWAjUOHyn60KQlWoTrsx4gv
Iys5ytBZoLcivwE6q96fuQ4oVmsNXK5CmIQ3awQTz1urgukSiV8MblNPyB4PB5QOpZvBIVOdjG+4
nQUNGF+9NNO424m6NBDBJbkUULia5p6bvyf3AGVSZiUc/lQ+7ZcRBkYWMYjakmn5rHaF96CdlNmy
tQZpP09NqYKG721mbf6ba3Zd2/Rp4ejqdw0WBUEpL0evz0TItlbyFmBMa7zaVQcgBQXfAv9hs8M1
WCgx4+7b7l3VxEkHj4mORZIGCnimsqDv4yUE73kTPxXUTfcUY5e/5rmJaS4vHOcuxDLA6sp17SR2
0mCQlgOa1fN1yZnIfeKHjtz39MMYUQuLL5mR6OZWjQgKCPpYbP3urLqZSp2MuzPZdcy3nZkmOh/4
nQcFtWUU76AHgv9G84y8twiKTx4vVEsvrTTKjHqVlvkB5JcbiF3zaLfJnV20ripoU0z6+hdsoHEL
drMEQD8sdZk3mGVVL5HvVAKSTs76t48wCXg2gDf65hNG73w0Swk7UC0h3HXlJgtbAQMYByVTxiWC
idVl/j6xrUKIL1Fgo30pOT6oWA5xn2afAWKVW5AGlUOHFXFUFhJZSjFRcg/8M373zmxh1qYKP9k7
ALmJa8W0pj7aY+Yi9dD8dqxVNWI068RzSdit4lz8Gnp1Wqr/C3xqF6r8EqKDFjNBBIfe5CnyOk7/
cEZErqfUX8PLzyrU/7OF6wHK+Yv0UbqaQSIqTC/GbBkUo+0uoiKJ2C0QdlAt8oNNQTr2WwRcmc7R
05XJ8UYjtx5Xo962/7qrZjqRzb93Dz/77YneiRrxidtuuNEasLFxwy06vU/LO5iouNr+7HXur5Vl
/avE+Z1hyuDoYtxPCwmHNrtf4eYtQNo+7ReOcADbim7l9CuXORU6IsQf1HuAihR8skn8TVxwj61b
fo8vATcEoQESFrMr5E1JLlFApfyx6AnY1RC8VdcKR1VNcLGCyjm66ArOpVVKjyFg3J8EoVLFdibA
25AJ68YUWBVYF9B9leaoBoGixG5KVUoJUuYVMjxyZID8N5Cgi4RPltHywkma8uMM0O0Zx5jWwbEP
fJOJbGS6rhJ3pyZ6khtwWKxbR2B+cz0OeDyVj0T7TXay4N0PzBxTyt3K4UfeOPGanMJr4lJvooFh
nsUYPut5Bsm1ieuwAl/SbAhl2+CqzxcWPA7JFcI3CFixCJ2Usm84qtowuD2ns9xPMBcFZoQDJHps
C3QP0gMQC6iNGfDToB/jZNN4UrX1wdMQPRgXOt4sDZCe1JXtvy5RjBQBfqc0/KKePP6A4xLKOnbs
8ryfD6DJGIxLGhK35NXaK8q9SrWHaisG+ThzqTJCKcA+X3rWV//ifGwExhcoJ9vernzO9N8dKAte
ZmSgdg/FaVlzSrfpo5ENezbgO/s2xe5brxE++n3V/EjaKINj2qWwM3nc+nywCHj9sEfOOmdl0eVf
jf/MCz4OwJ12rOc4PvfH7hTjB3lKHLlSsxKyi/7luJHpEx+vdmgoDGJAXUL876Kwl1yM814Lrlzz
RmKkzTiZ7XLqTLa1GPif+E64O9NUsnobHLaHYRFQ0RPT8Foi1qnsXy+ccRJAwKXkgwA2rZeAxvlR
xGAvNf3ubDdi9ZK8BXc6+FSjeQwRWN/DwN8RXXIoBE+30PYHnb8sRCAwBiS77B9QgUbz7HOO9RDq
1on+eWlMX/4F3gdA3rgiCzP9Vf1k6Ef1oh4fB7iG2RFSf6KjHNzk6BBautze75u0/TVDZl6pnrKi
B5ajXuHxisk000TJIBwKz9gD6I5GjBavEK+pCZI4akWXW9t+FCxcKRsLLlIToX3joJmBYKCYaA+U
LKHOzkT9pMovmovNEutoD6sGpFeGu3N9HzYyymEpKgL7jd0CUAstYayZ8MW/YQSbq+tkntItpoaK
p7L9DiiBMXmRbaLY2mFfWR1CDg9TBASkgLehbNOfh4wCGD1S560Q/vGtzi8fdndWuBO7qQGQw96/
3K7vBVdQhOcj9aTP2Y8NT6xJIBAfL5x1stl582wGygqfvPlGX2SfF8Pm/ZKDoUybevp6jT4xJThP
cuQuV3cvhqR+Wekfo33042EVKupjxPqi3Je22XOW8BoWVR08SaGasvr/orqZuIABR81/pB9SuwAK
Z+Z8c3rUC8mcJQztCasMr1uPX+IhccqaNtj7T9IbsJmKiomH6CajyIo94+P823LCG/1WZnOcv7SC
hsi5jjr4OI3AfxETpdIVQqxcKxdnQS8Ws/SzeGPKFzYE0bP6346TtdOHkh3kl2JJzY0IJO90LQ61
p4HPdGwnDWQ/7Mv/9DV3lu8vuO7dPf2OFqHmLKDe/0xgYhKT1CcFaeDg0r7yaxrPUnT+L21zJmL+
a40num0XOyRWKLwAU/hDTm+oephfv1bY4t8l0JmkdSF69HuoqC94HYJL+6vfERQf20WqpVt2bFTD
EdEugf5vAkXsG3rtfnwsfnL2FNQtOIyiU5VApwb34BSUW7PdU/dhxx0aMoTeGp8eBOm8hm0DUGUI
IzEcrgoZ8mEXftJ0VuMXGEUuL+ZZvMsrExKNuntIjG7PdFkfjCtkMPEzkfCzjenVtTPMC27DPfti
9Fh+PUVJrG4Q/Yd5Bma8K+XVp854q3h+2kusbLvDh8rBJyTwfjbpO1wkYO31gxdbIRhTTkQ6KM0K
oJEMJ6oWNcbenkPK1flY6E1kxrEAkCSgVY4kaO0lga16NhZvOVPoirAevBJfgOZP/vEEhOErB6+R
uItirGYIlUbHGkswsoeKud2jYoEu7aba456a2tB12yJvkBgIBycAd7SCBa9oGn4ojgRIbBw2jCEx
5dIzsg9JGMzRX5nis0FocP5Wrk1ix9/uZTn9CA/G15K1KOIYkBRj8jYrMe2oueFG28h/5tcYCrv8
Qs276BHXk514X7yj7/qP1wmJob+DWuDa661Tep/S8QVxUMab0JmfzE6E/KLCVPtZTGpajiann4Fz
QcnWbzUD6W4yBYCmGaIxAmsuK1d9akHk7nYfG90GL89eUF61+7wVsTUiIoVXHfeFytUN5IX1K9Kk
I/5EdJdHhY0Hn8bc5mjrEHtD5HveOw2WAjYQ2tDLttiKnsidn29KUU9ps/1cVdPgobfMCIupzspJ
whDV1RfI1xwja+7XKJDWRhUb/tpE/LYDwo6Qy9xM6OLCeCW+ua2Gwvl+4MHxunQhk/6Z2+ArVUv7
BZ0t7k4xbbVt53QMLysnnEx+owBLTb11PgPZmcAq97WZV7gIt6w72XPY8gEEl8Kk1chjy+90Vd3s
8myRD3VIJFJuh4qmU4epERmvZzcoin36QNbnr+1Js6tBKQEb+gIbWxygiVA3ENucDh7QEHbw8Ws9
TKLNP9PXJBDcNx3pMixgiBG8eAH7UtRkId96qta2IGyEMLIkf0E8/hOcSQcBCc7MLTVnoBaat8qh
YEhEar2Bq8juJLbp+VfFJmOyhp2w1yLmvDH8g4D/W+PjeXC41upZF/sW5VqMgm5wcHIq73Jpr3pB
X2tud59iIg8TQkT17BqHsFv+TryzyOnxCqOe2nzze55wOkCYokzSBh4TWlvsoVflbDFbg36YS5wF
eroLBGUPndWgrr6TB0gxV2n0Dc7jSckkJbNaRp6WqG736AhYdSyUSq4WXLoAMpoQMl0Ik13f/nzE
3e7QmbwqKPW431lqJzGjnFy83iJN6kgIqmYhQeWkxbpu1Xl1GFt5r8d/v5BUrkzaKPAWInO0NHUG
bSrPr0YcmosDD5cmz/31nyRKNtVFeZlQAPIjYu2wmpBgTSY6mSHXSgHdEfVVqzNLdhiykv8xYriy
dTaCBJ+igHpXDUKmANdsVW4OrURgJX+iBVlt7matNDGNNyn/kkmHYRfbSW4H14r7N8U3G6pyWikb
8DUizpi4R3HKBq3qK9VRnEJ7u3qLvjd4CKaEwXxpCbHraEfhfPYZqH4JfOlrsl9Lcn9P9u3GD8dp
ueJf6h1kGEcvXYC83UFrYJKxXeMf+y+4yrY/nI1DtWDhHSOTJGQPvYsCyJ1b8gqc1jZiX3HrLhjZ
YmBE9elD7UJEMIYEoP14LIQUh+pblRMR5FQxfGWbpKRQT6z5d3bKIOwpt7pgwEq/vx4K0K6T3np5
YDru/P+14IafQXL1yKdA3ENGPh0vHVhGGJiibILby23JpJyTvdrGKHQoUz5QHzc+OCDb5x3vy2XV
UNYrbjcrpNS2xCte45C/RR6j68R7ijI25jG1MeB1uBtG994uL4+tPpPRpK7EljMEqk3a13zX8fJR
U/o3UmAujH2qjNI16MFV6qrcePH59pZ35oSX2+yIf1DgAu6P6CkBTEioBHwsUPaTr4+9i3wjptpL
2Cu9D65SpveBZa9yM7Iafk9TPNMaquTsZKvPcuM2ukTH4ZFSp8zKxqF6e9Z07CPX0SWcDHq9UHwG
CDSz39QQSjutDfO7CA7oOwAzIdWv+Umj+HmGJHl4wOqbAzfxEg35Mmg1OjA7NYBpKrD3AYokIzpx
Tiu0/iwSuyVIADGNzVHkFUxANjhgNTcsltt2RPVki9bayfCnbMFieXGSpdT5Zp49mQ40/VInhI6x
C/bGWE5/WhtcfvI2kl2EerK1rqgmOzpGRvTbItuD2oB9ecOWNXUY/KPIborOoEXp58ikgqNPf1Bo
RTtZdddLrdY9GZsSRbYW9Yzdy+tvxir3CD4JGt0QvAUDfnqh6cpfsXhJfhPlW0astIB5PvJ2VHTa
8GIx/5gGi+e9g8MTSh4Ij2gnIOoedLV0SItSqmpJ+vkZ8++AwP9Fbpky21EYchwKGnW51D2Q9bjd
MiHg5upMzqRJ6J4KuLTANKTII+g2K7uJ1ejee5kvWkOA+k4VDaTfkjP6CzuX/SuoZjZM4vDEgnFN
VUgrPQb9cqfXnU7Xu3puGI7PyERyZDKVFBrqN6xUrYhfa+y85Sam1V2uT95jpsjTQmNScWx65AcG
SUCGnlkTCb4eIUZslHzeFYH5HpQma24r8zLezwarBE5m2baXZ6ZZSHjVQlbXv3G7k7IPgyNi3WZ1
NpjRkVl4i2ceanNP9703D2Xxo2V9cdME3x22naQvMLelgtZFcSW9f6FV+92pZCmyul46SoLJekAr
6T5SKGH8g+xUqoblgjRQgZcP/FCq6nial5T0HguYd0wqrmS9hf4pr2B0u+v4bm3yr8NlIgPlmu54
rzDMvCOLEnbIM83671vhwmrTmvalkw5rQy9TmNVpbMcmKkFiZF4vq+CHnKzUP34K4eHFxXTfbAaL
EoyCfTOy8wOwYeGYm9ewiCHaNY7hBorETBq02lvlhnnPYAEv4jkvFKhNmFeN7RVTsR1ccRIH3Apc
J78ieFqmf2ochhf1WRDdMYMo/CU6TMcgZ/TPtfAFDA5j3vG4ThhaRHljs6G3hOcSvzTWuLKQdPUQ
E7xPy9TM7cv26rCjzAY3sZlgNoL0kLHx4dsYhyHeBzIzMwT01HpP5gfJwloZZcpYxf2zmkXLA053
sVf8mZ1JHdlWYCK+a0VVWzoHukPzjq3csijY1fGqc5zqw9gnrj4p0Fl/gb5ya2kj8ZSLnM8OJFEC
G5WxytYyRoMgPpxhALV1VjDLaZHjniKeuDIp105Q+1zHzNIFrpM0taVjrdrwsmTcPwCm/9fruMn6
H97d4ykLOy/3nesCrTcPNXHQCn8YZ/Eb+d7cpQujj0nxCtwwucLP2t8e0ZnGBfOfJ2O0wLNfodQg
mNfigFt59LJynwhQDvf+B78Hdrhu8R5sAtlv9ZtQr/RuTtnlaxiO0kB8U2axDosqqvZaYYtlAO5p
aBL7Hx/BQkd6rcYPGxm0elNS2u6q2WCN3nw0OMCl1Oy84hrFULEloelgwnD+g+AC8rKad/qi+RrM
j8DgDiLgTowNaty3cxkgMP9Ex+9Pylw4DVmpzz3PRIeJjmuXWbcVlafX3F4tK3okyKGBFrhOvkM3
Eh7YWE3Yl5zO1W1TTWbU3ycA7Mzf30WLqIOPn6Su5Sv6IUTJCPrw7rdmsWdP9fdqBA0rvHOYM24G
No0xEF01JbaMlhu3lgVH4lylC8CpSlnGu8W0yJs9Mx4Qpqc5Rf169aL/YdtLCyEYg7NnowNUKxPc
TzykN+xfjVkZVV5rzz+F6YsFTkTA/WPIaAbzyWPXNHnooLL+rISiK1sEWBSvfQSinh6+b0FHLVmE
7D+WQPomMUb5yaFg3B952mW8WQDYQWC9KnYU4OHwLtnvpeF64I/tbPj9wQhfjYUN2+y/eycBJe5I
09FgWEe3vDngjY5IYnqd+gxDta8Om+ruTIoBak27HGhVzbBotL9wY09mqQO4Sf1TGGJuO3W0iI10
ECVdkGmtCp88XAsb/rMu11oQjfwz8s1rTrtDjqL4FfdIxLvHmIGvDXPlL3pjw5SdZIrP2Hx8nzY2
F1EVRKEytoleTVzQ6ss5y71/N9qEFXyxXBRK9/U49kJlyyiEf2XwB870XUvlPXa7dIgeYfHmO+LT
1QwuRi3GmzEsIekfCNwsttU02uidUd60eBjrA0auyv3wzBRNxPTnC1LDcBdL3KJLVOzpfoXi1q+s
IukZkafaByErbFeheUZTx3gHp/w7RNpzDuPFbcpKLLnJb+UlAFZG7k0XHr4M0yaIEEQ+bvYZcWIT
z0fb/yhXL+BoTPbrJrlc5PX0k6TfWvjW4SEjv+VxKcYI4uRju7m5My/CrBbV9wpmU/uTN04wxkLj
mZ2qs+q3dvluHFaJwasm4VS9LD63LZMFI4Qi/Py1CXEZtKSlLbE2BXRLSXc67iJ/WuidLhv9oTuF
ClNZaAz9hsrv45uWcUYErlxiXDbt2JcnAjOLYnldgxgEnArCx1cV+7ecqqPfhDPdwqHaJ6v1aqES
xyw0ZjoqeGd18DpHpjPg9M7XEjgreYIMwdW0LC+DdpufjHMbyf/JId+60FtlPtMJ3xUqpj6MAsR6
wYrWH62AK9cnrY4Spwue8EziBFKWSN195xgXo6W1xV7XJrdqSmCx9gloqoYLEen2igGvxPmA1lRU
KMpwkOtKKxdbdWHFYvzNBMPcXo37R2lyaDQ6NXzyfGYMcndf+KTJmfQrioDDBWvES7Zx71nmZ4bx
VL2TzdCufHG03zwMuYlOxntd8LSa2hN17BI3EHKJtHD7eSZRfQ/g7ziF3G30bfZrBd4zgpOpmxJX
UGqdONdLTcvTKqCit3pg+NWaN76bxeb0vXZHM3NW6Lp69hyq/LBs63f4g5ExDVNvgRiLttxYPoN4
bpz2iznr8vjfAEGmaF1sfgOIhLJd7Ikrou8zoaF4HLq0i6MHBAjUFEIBZSIblC+AJzM47mvDxG3d
+O6CfoUZfxVcxQsQ9IbARAE/czoIgBYLTSOrj8u9DgRsQuX9kXUrfavFF9ed5WKUBugWFeQriCvO
9P2pOhsPQvTJ5e/fMUKA7TuFLGrPN/uFT1tO8pTUEdJX3ol5YJDXflY4phSCx3h9WSzMz0A1MjWk
dfbY7gUFbaArSw6GqWda4chkASA7Nt4zlERADLiElR/bfh/bCgq0IoTdzVwlskYTfW8jvQuyDEfo
CtLO4EHHegERBFLEcvGlqOVtGThCq9vHFBvwZeWk+O/Diq+t8JuE8vsW39uVgs2puI9LjARu0045
ViroHwp6rAR0xrDhBNeK5EROGgOEEy/2WHECI89hm2XlrWgtA1QGw5icfF7Y+uJgFEY9hju8b5xy
AARDkNtH+7x4fO1jKoVmM/XoYrjCUheg1Pj1OqxC+xvelwmq1Z8ErWfzlnXfeh63uB6FJ70JGvT+
BDEMoUafZ6drkNveqTiHxA21esBAI1kfXTF8MYSgK1foAAiQAS7koi4YL2+d2kQqb21yL+bNo91q
/ZLM6WSsk42kzjKMdocBYd/osty0Hz8rlpF7wK4IK0RtIGdq/hEV24HlW5HSLixwDjM6ZoPXrYvR
c4+mFLw0hKX4HblozPIu84FQOs8/GKCeE4YymT0xiIDedDYwYKwMhKqTsylk14AL1nw1udIUlZWd
ZQNmNY3g3Wl7381pPrXu0NA1G54VUxKieNPAg0k/umJYxe21IwqLfhExCLDLrxNEinPRAj6Eeg6d
6C3kRU4UByulBs786/u1RPIYOXoA8QeMgiJdrdD09SvVoxiFVWNGspAqSsZu6L0q9FhFIlFJa5NO
Rqfp3jd9FaNCh5l+bmoA8xVpFCe05zPV/VOEQqE2NEasCni3zRqXeJKgUGWU11ouvDNWwP7pdAhz
5kjzRImNwkBq4XqnavGEc3luZEKtVUMg0rpexrZ7bg4cAb0BlUud1WRqEGjX+1gD99Ck6+oPig8Z
orjCAJBWZlpLTxAJfarynwFl285ceNxFPFqvoBrzJxzqhprzbwmsGr0YrzVMfPvZIQAG5T4EL9eA
JHpNyVN3vWX5uKvycf6txBb4O7c5BT5f9Mkfvxnl4BmILvVd2u4Hp9VpYZD4Sr1ecWm+vp6s1YvE
3MU1w6JxYyaPIBFDtxrwaeDAE6nQ5RdGkHa9ysRHMAsAgUpxw7MdEVZ4qjNAwSdSbPg3Z1v5J+xO
aBHidT0mVOrl9O8vG6LIaD5RLs8pnmfYL4dOcjEitw9dcT7ARtWxxOQhtPHRyvWuRF95D1Ut8loQ
H6nEn4EYorXW0Z6MVmOCNebG7vpJoemNxhsqponHRe3rvYLfCvTpywvDxupkVd9AIL2SV1nfmYb1
/GhKGnJx6MITm0EUw3+o7lvwr4TSHzWJc/eCMnc+7DJOJdKhMKe6h/+sXTRhftYzy0Db+Z+daL8Z
OLCqefoV8VoL3cUJEwkvqssJQrIyWaqNL6gMYzJ6V1NGYPTa0ZdN3aTDO58XtmBuaMAIcIvw1ugu
5u9KniuESmqchQ5MbswURfD3hU/9P5ahunGPW6AV1tafg1kAenQLjQbhp8zHuDkLMD3jlI+C0BIf
vaP2pqqucZVvSvLDiPx2WkJvG4ew6tuvuQyoGPcHMjDrzGLtpf+82qVPsKA01YPRThNudJKyPgKK
XOfHBhbK20mZtjT0HFba7aTKUfhZz56waRbQXCD6QCFNWyFU6vZxE+dUcs147Jb16EzeM0s8lZJK
HrJ3CTJ7El2WKbmmjlrDZgmZzFZDW7ZNZarCg/EiqeVeTYQHg2FGbyv8qsojkDWwcijJzV/hoxq3
fo20t1LjjyZafUpWEDgywLzCgiH6yxF648UqBDYrED0VqXo0TdAJOOkTjgrcgFdPcAlbDPy9k2y4
q13WkgrytFePaqKIXkiGUhBBKws0Qgr95J1vziKUn65UODQDG7aVQtg8EMJHujZ94sOX7PL5N4Sw
KzOE9SevhEllpfhxHyZIr9QvKafGdzPbmv3qjFefd8RGqjgbcFgy6Tpn4Jzo+/ayVO+BYi1KJ41N
rQxS10s1jsEq0WEAkgdLzjBIzYpAqH1Z8c5s17Odo5GelcPL9wzDY5WoTZ7Eczb9DfAdQqZJqh4O
q5FpNSkZIvXd+lBIsI3We0Js+d008A+PBiy1sV2T65qbXn/7Hrh5Oqx7C0jF/dqy75j9alRsJemo
O5UmuZ+xYbpR7GX1HHunO60zGUjKwjr4EVvy1bnH4cMj1KgstEnDriKNVjfuDL+aiOWWX5zRPvgW
+5JkqIwUih3Y6paKZbb6aCq1DbcuZQ7c6UsvvXr2/RWwV1KUNyoane8lLYOunk3bxxNRMsE6jOTG
O1f49nrSL1BBku806dmluu5UIwBl0Dy2hTdC6XIkUuHby2wgKksO1eugP0mUZ7gutSTHGSfa6wDg
GGOqyMSGkjADG6CQLmQty/cmsC+w8bKW4BaR5jDAlY6kLthE2V4JKN5CHzAT5CNAva7WbCjTCYD/
jy1/19clwopd9C7h22reh7lR+mQBPFR9+xHCGHWvQ6HXHDeguywoYQC+1SYKFMZQf2vyWT0fVeR9
oVNZ4IxoaxDt/Zq/L5q838/UK8NTM4fDIC7a1kY9ASvc/hf8EQlqB6Az6zVPc7xVQcq+oVHMmeWS
KThBCrvnKnlY4az+evHxYBfNJpxrGfVK+6hGdaduH8t6xqEcqAjd0wK175+yGw/9jpjrOQBt18rM
FxryFApmX9AQ0+IwEN+ODEQkWBVBJWB7/oaNupf98+lT0yXyxCVWyLUSiTTrD915dzPxpfL8lUHF
Rd4F3Cgk4rmAM1NHBF+M1wgTKm9hqt55lPSLw6Mj+02VcFR5wfACOmgAFOoA/FZxffcx7jyiktE/
hCAFpukdCZPdUYS/dvI8B4Ckfs0TffGI4pjC+LKdctKRtp9n0+fsToull0gNIySZ+OLpspj7yfs2
VyESCLcfHvn6NY7bnuOB4+gkwAPJttDCXbk/kCRGYIAhVdb9Iv4Used+CWBcAnq93ByLCnawYTQn
QKb7FmTDO2SnnAVwqyyttn8X97GjFurusOrYZTyfVsEJB0VTN9e90GNUdNguh/90H/Nx1rK1mkse
8LC31MBdUr+TMskLS8BB3FIvygti4m3V03z85hFz+MRpCPVeJHkBIsDY781VvJVCGcjMH7lPSMY2
4bOWHArABd6Ficj/mswelduVN/DCK0/Ht/dBc/MTYIbgM8tl6NJldAUl+9STotJzPgVga45UJWcr
w5fVS4hMX+wMjWWMVx0sMJQ9936sVoNejIbStY9OHJUiO2NW5Q9H3KxzQ57xgeWCdzzhBXSTP3bE
FlkThak4CD07TRd6CMlT5BKAnFWRgIkhvA92RgdaKmmYBM8Xn2mSHv+hmF4KY8A7VnVaHGto2RMH
NjXI9KqATPQKTDu9PsN/UtXJZvIbTKuPe2AC/CNcOUUvWY4imJhGQqhiPXZzoXzSLhjC9rBRMhog
fu5y+tddYB9Uvi7mjOxnHsJvk+I/bb0ikrHRqK+EnKLRi310kpCmRwnjV0MxdVG+A4aVQJsn5Ipn
ZgBpnCE53oqULCXoav4k5vrO3kj2bQiBAcOJsEzaGvJw2gk/uhZiDEAX0tAtEERVzXUap3mAGvgB
Q741/ztfF9cSj0YGH6ojq8hz0v6x85LosCN4KWSxm6frUbfx6aTAq9171zCA9DVBXKyfpjajN1dn
GX7jKQHd5KwjCWc0sHdM656yVI1tDWQ/OpWeYNA8vZS3ldbEf0G5hoNYjSIGIPusV9fBAd4Rq04Q
Zfnh8R1xQuDm6vipBvmtqpUtrsaWHEeqJ5PHNK9xEN2rqoa7MzO2tkXtztNUHaZ9qE+/FQuuWHOD
dp6dkVXTEtd1+LKsn8gOuewWcF7/E72sVZDv0tj2XlwvwJrlvHMGx8IMj9hmJZ8n4BokZ75YGuV7
/7gLX/FudDVHdfoF/Zdj063ddb09WR511XpGOFJIIrRd10q3GTu9LMcAlVajX/2JbPRNdP4BHk/F
UM5WJ7sL/T5Vnytsx7z36qEL0e/9p4UKF1WV5Wqu0tGpr0UhDrMAtYvDrrI16UDZL3i2nEqp1mFc
mOwRyDB1YHo3IvOib2Csxh3DZ1w3VXe1Hh6vyf8klQYmMEAJmbGummwTSSWd9C3z04yISaDb4/Gu
MwOFwdHrny4d3/8rAY1knLeEeOffBx9iPaY52hqo9xS4cW6tSpBAbgVzRmjhDpXm+95UYh1lb8oN
o49ljPRUO/FxMow7micXe2C0iFkrssMz1wtPT9qEC7oCubQUjVoeNMJ0MsBOHHtEkYRlW528GacJ
aLYtDMJwYjPPzRQpB+I17LAA0GBYMb5eGcEiiMAk/xZ8ncYa4zlX6k61RMbrQ+eBFCvIB3Wh+20F
Oo4iQUBDyKZQP7/1G5lAWrbvS/WKf3ptqhVht6/DJ+rh4WHfvJXLvn5CpP5lHCfzo/FekaXK1AxY
Cd6TVFD9fqqpW+cgs2LQr4JMiQFQLTa7gOq5FP35ySx9Q2AiaF01Jlw+FndeBfHJthaEjPXiMwAA
ZodLe+4ReXcqwWMOUYv40+i+GVxhjQaVPBgGXKTNUi+CL2xqrpsC0OTwt7IzBML5dCyrPIN/2xuR
h1afJRq1n1ZNy/LJpRNAggdv6A6hwpztt5XnD7SgQ07u+R2V6FRtb2CaCmlkFWkFneIkrxdoDnYB
8fsHDaLa5KE/D2OMkT6UiloQZtMQ3VzJgyom6fAJaibCx0+Q8C6zvzrTQwNqIBZ5Kwz8LzfS0Ag0
XFmmig/0MRTblZ0BBtYda5Cx0lXtQ9cSN17cVJfQ5dLaRQ+xe644ff7h4hZSCpkWtUI8COv4lR3x
CAMnyLvH6ZFCKQgfyAC4ZRroQd8Po1HfQ1vYqlYQUW0q4lVvEanaJ5RidZzUaPbPmeBx0l5+NeAf
kzGyuGr0K8MaATod7NRD2AiuV9r/sn9M+zuSKGTCH5qnj2JhI+OGG3SNOV19dTk2RDthWmkHsZqe
ebm1LTMbnhOnEeAcM132vtBaLEmPUnfAFlQkmYpPauUI3LDuKWujv/6Jl/MCqBwsM41gOW4BIHcK
ys/6HVIvUfQlBngvET5YQe/hufDjg5sjTtY/unwa3Q3c4KoIdh7asKzY/XfU28ZJd+4sfkIrg1jQ
Ukz5cEEDzdQYZANsZ1WsWItygOk2kOHs+1VhMRWooedtZZ5csNF+YTpoCtAd2Ceed45bdPtaFGa6
TiUQQ0ECgnzMMSj5SHqDKENHuN1U1amPDbJccT/TWfb/03H2Fxv2eYMYpbndkD0vTpKWYXSWWoRV
ME15nyAu0bMa6WUibMHKyq/sMYAoOH2p2dYGgFGwBoorl9mXw2AoX960l23rC6iKvFYXmIVff7Gs
lAAiXnLVBsHD7VIbllRhiimIsn8P/Fk9c2dJGYzWirDkSTuAulLVzwqa5PANxS+NbdzBd3tjGQf+
A7VqqDAJCUogus7rzTo2D3mVIeycbplU5tN43nX+X9mwA0B+tVSwHr0jJmMDO2DyYADWpaTok+Jd
r/ddUW6sONluBIBNqu/PiR/bnCPF95eW2cGGDTf5S6KCG5P2dfKijwve5MuYxtQLvXyH0xVSnH/U
71o8zA8g8I2jAap0LuKcGMFKoZ9Cp3Ii13Wlr6DItRq5HmebZnf7ZiHrOFFytPMBAmQzaAcoSDXz
LZu4/aVHjz2GjAyuHtxTs0ZUxJQB2FJxIX0HupNCgyN4JsMLXQBntLZSWhSvJfrzme2DP1huMNtG
dtIli8U7jk6MfPbkJSuVg91WFnkyIpWt90DdtdnlUVj3F+h4yTmViEA7/N3mpYWbadU7pn5RVtOY
J2LrMCLtI0EwaZujDnVzmfa57hjEiCLe5V06EVMA6Ip6A9pcrophYd+eNFJhR55zmn4cHdok4v2Y
meztrep6N6hDTYKtTEQPrIIoGb/IhfzQhOtE+hVaI1CX69gZif/7MJ0xJMN7676h/1wjf1w+2TAF
NxtxV9rSYOFh6TkuYSYiuMORXrJkKXsy5k/n612sBMEAlYVvDRphc2XSjkBpyX6hrRhTfCHChqbH
MRVoeX08A10vFHiS3ZAv87c9yhDpaHU2frQelXBVOMpKQRKyeFgTII2iIJ6VLvurtNzqoiubepoh
RGrjtHxrWm9miSJqjwMoSH46Y3pmedp6Eh4k6gpkY2JZstGRAmyEkib4YT1NPxTnPel+DRHu1JB+
O4b8f7r5sGnySCZqLAaHs80BM57auZxjv7y1LNWOAzIn5UTXnmJAn/oLTi8vshszc3WtYGUDHHGL
oIw/oPWkru1RBSgmdfpxPKBxNPan6+T0GHWOZ1oStD9b/MI+5wgs8dUZVAIH5taBIdVaiEFMXmcn
aoUk/+6WN/GFuoxH+u8mM3BoOFKJ72Ck+7DsWYMK2SJ3nFV/prDdfmy7Hsmj/8b5EfUbYfV5T6xO
wO4s3I3xJaM2rnALERGUs7LxD3O6FPDSZga+ND5koZHBwWc4cG4O3j/SdE6hgsbwANBwDzrD+KAC
JP3JTQFANbHgwS8RCTovRzoFqblkVzwxppXhkJg7mFtlgNL1pHOEdwVFC0k9ihNOCwcRXTSUhtiS
YkkZszwiXQ6kmGb0VeJbPXMRVgiBG0NJ1juwxQkeLf98590T5hLQd4SMjiMJ4P5365BrQ7Hn0JAj
+/oRqhExJ2f/SwQeyNCrwea5eoD5mu4tN7oIWLTwOU6RJJjh2xBqd56QIBUxKhOoKNKKrYlmmpET
ZqGOLMHz7zl+Y1mcCkxB6hlnuiHgM2hgP9DSNF60KRBCkPqFPh/LuMYrTu4mpvqV4+/ibQcWCjPI
rX3+6G3xiqXqCzjwbAhHibu1Hi0st3e5WOAU0yzFhX0aAY/b9gEwpnP7PAxa/mf7jZxDmzWPdaEV
MoN1EhOhQVU05te9yrqfxW1YO2YKrnKCI2cw/cXznhllDoWg2JDXM1iBmPRGRGd6AYXA75r8aQhm
Qd6KPPncrws0e+dv9D0ycZ2f1tOyayEM/JOZE3OFuB+3LE+7n5F+73LlfLzmENPlgsEJ5VzHt+id
KnIaHo1wSw6WSWo8YKQdfayOaAS0s2htHOK+GvqpM8XP7ybPdKy4CckV6dwrVtOSJBnr0FdA4gQE
tPaV5EvQ2TYhpm8IQv9sLtDv8XeLDoiXxdfo5KoZ6WUT6b7AMt7a0SgqJRsQXGQxjxOwbsr5IL5K
yhqQ2zZdehU5mptI9fw+Vq2u1zQIMv9nmnG9Zvcq73fLHKfm186IsU5Ke1CTWpvbG+G61OIl9JXx
pFSYgZHwkvHDzEopwyt+to/ZM+uBGJf/uPl0xeA75mZbB5KxSYVevUkKUSjvFgubTp9Q/OSV33Tx
hTq+Q8TRtbTUJXyDTv/TxNneYQW6BMI7DRy1f4ucATi7E8FGa0kZaA/e6O/vjvTcPWaSD/Q1o30r
4sM0vHnRNvl+/YH88PURNKvcbJDrKDA4G4kVvlGGnLOWB0edJSkFOREbPRVskq/K/i+ltpYYjbxr
shMkVLjB2UzkPLEe6sBtxD1TDuZ7WPaRIT4hlmCZRef+DKyEcOu40qNa4iMjcxZBpvNwXjYLOeqy
oR0hpy8YLa7Khp0e4a72l4SeCSfzMJM66AqCvM/ygc8RCL1NfnMDVPfzLuN+qCGGjHjKxSeAG6gv
130xccdHcGkgUdMnOAVC+OmwzdbZjfi9qOubYNWpQReb3uuH4aSGrFyrlLaFmZKVJpNPgIELIqbI
u9R+EiHM3DxrbapGSVa5Lxx81O9ZdIXNUao9DRH+C/CD75xpwJ4eZirfXigi6Bvba4nsNsrdAZ36
yToL7ABqYAmXuhUoatY0mhPU/7zMMx/7L/2a4MyPLyO1EokCP4zgpqbpOQ2DGAZPZbk8u3a4+K3H
YEoEOIdNZu0Xpv5baV5st5cqcqITAsFlGLC2ilFtV5XHnJV+w6BofwLRhEJ7TnQEk2EgtJByj/X2
AXZhFzdHUYjS79m/JrW0fD8i9N5Mw05+iyKmgPVuxoA229rkfdOEL8J4gknGMm4dc7aczKF6T1YT
9yLPvyPGJDqE3LjFNJTGyTvn+TGpsDvC3wZyXsQRtFfVw1LJxBkeMwrmQsb7V253W6MGp9o7J9fn
glSaulmkouP0sJbFsqLUamr6Y9oXPSbmRrBZGQzK+FdR85YR4VpQuTqMbk9xq7UU4SKu3FRJr/bQ
57zfIFulwAoG7eey2PC5Qr8nVaKRVL99O16Gx4r4JYtVOFTto1XF0YW75siR9lC81mX0c5gbhMVO
C21AWUnYCptbVYbjdtuv2UkTwYXV6wnO8/56Q2HSqYbwR8u1UVAuoN3aIU7vLygvRedm4uB/ww5C
3ekhimvyICEH4Y+qS3n6hSa3JUm6CQ3pdiT1CzqlOeXjl0iFACM7bwtc48i7GKM9iomJsDsJF+O3
mdzWzEgLxpnqaMfhaF6bs67f++W7zQ2MlRYWq25BNJnn8ycC0JodXlJukKUUOaKwjHMB8AJYCh+C
ucxABG4CqbaBudz75+5uC4j6jkBUWL/WvAU/uD/llbXa0pwUpeTNaetlE2kryrFdaj/sLJQ83IpA
MCA+vB1KYwhsqoKEGa962Dpm0lUQbzewY753TyinA9v443wRSjNV1kPWZvfMou8TDTH8hFStoVkJ
TBK4NoAuapeVdbt0CZCt06RR92zyNtjNnql8NbRNC+9I3HAzdCDGJDZml3uHuaq8WdqYnGoDaX6/
t9sJrIyBTJ7GmlpzdPNxnmsfBkeNzhUgzhH9uKkPBgI1b/yWKyTVwHRd6Z2uBBhJaHQI6ITGQX2H
UNDbGBrnXpXQGxaVBX3G4ZFS7dvsVqY4j9dWfBivTxqrmTJuxScPZRgWBs4YIX0zh5XE1LT9NVil
01vOelKI3h2sVUE5FBT1YhGaMjU1TO+gWmAfvBL7GQXD1/w5f+bs/v/kPUFKbQ+tXMe5iktKg2su
+kigOYojOI+HS4tRkHuDvHPETzxTs2CpzPG9PdgcAHEkLdS+KaG0I8PsH1GwrqaT+OYLoVpLn6Re
OTGssdwMpGjmQWf/0L/37GLUY1DeGqTxqyp5Hkna84BiKraRXxntiuKhNmgkIR7M7WuewCAYTisl
pm00vNPzmhC2Iu+SthzJqXRZdm+YQXOlEkvvJ6zai1J1fqLT1yHPyOlDcLka6ghB/jFDX4xX96Vu
HBy0+L7bvWyEtLDTMVz7rySUsfhNI9ybKZ0308btlTmAts5KQyN5CUioe5T5STZyQz2nXByJ/Tnu
Paksm84jVtO+ZwsLIT2Qlteqzhre4QNLKrT6fP0eRlg2EtPv3DOanTZAT+gbs0KonDlYrp3RQ08J
UtLkl0VC2s/tJF1qHkA0449V8//BBGXXIipN7J71RWgPUwPUl3PrXUT0qtDFbNrn1/d1ZR8pQGlg
w5jWKNPHH90DvDALpL7sLj14+yrk86EQamNhT/2UuNWjfK2uq3sqhBLdNKUUx09D81fYREHLfFqr
PgX56/cuKE77bGLQQ1FjAbiEb+5QQpukoOZpPiEmybA3ERs/ygGBT4mpHJ06DW/OASKZIT4ma2o0
XOPig13l/OfQ2WDj1GxUDa0h/46zZ3yurRkm+3EsyWb8GQXPFuF4HuEIH63WK4jVZJWPQ/tADSFQ
zzfpPdW+05ZCTPiCRvNXNLS3Tepv3M1EIdrcfcVw4Nl2V1ib0veCu3PU/y3HFNzfgHyjSBDpAUA+
UFfVmLqVqsK7ukZkpdz8Mp9mWYoJX4P2cybyXTOYH7TfmDLhXLDmvdCKv68xsCEPOB6gFxHTb9B3
0bfkONFWNLXzaXDtSetRhevYqQm+P+JGYaR2kGksrvVJbwCWcl5azbG/oAfOdDuzmvS779tvHHgu
GdblnWSXSbsOuhP/LvYavizlyInx/8LsmN8iWxTe43/ZHatR6xzTFJIooTiT9+Q0emFYkmEc+fkP
waPVoObBatLMDRAEnRZQiXD3xzi06alvvmh7XNf1+lk+3As5fqj4bO3Lylc+SyM1pQrsywph2nSk
qqiFxsxizhOfABohhv9GcteFV59pEdcSXPrXB/G8ens+QRMD1LhNfDLqbHmJIxpk5kCywJxuTDVV
8Tu7yJrZLUSb/jqYTviDNCeEl/zNBZhiGMNSAlrhTjbS1OCgW1KvhgarkOU31gSebYcmQYpnZHiQ
iDzOgzTjWQHgSBanjj3DBhsn5IPrZkaPbyy4N/0bjFaZZ2ljE/BB2fNV5Am0c+/oq2gcrYIw72MS
BGMqePB7ptAG747srYhBpJcSuhmnZQNVGofbIc3hwtDA/OA3tsMHhuxK523of4LEMfDJIxjqrHRb
QjBJ4Oq9opsGdwptOa8cLbEbsRB3CXuJXO7IMDBNZJL2CyeO8kP0xcf3uH9ZbdTQa5cEIOsZQanx
mn1pK/FXW2dgBdbqWW8xFkSiLpx6Tn60fQ75LtR1Xdhg+/EhKeIm3wksq65zn/7UFVS/6DyLXmdO
7y8NkHD1beBLnJA7P3WQhRoF2R5MsmljSIRFtkYl8+tX1bbF28RsVcsD8XMpiKAs/czl7TrkG0Vg
/Vvjn+ljyRYJmgE0okXt5vvKFfo3VbG02iy0neyi12uDIFzcaeem+0YazTDbhjcqckpwYwpGazbG
q5ZW+7JboLakB7DmPQXt1Hh0fDoB69zRagJFaJvL41p285IF7ylQhW1JbIfhg12228M2pgk3n5vP
JY6jnEA8vFKS8d08l5Or8KaV5TrzjoTGzeJJA6ZkWQlGmIxddX5l78gDZrJYrDXaPWLi78XOxpwP
YYLfQnIUnvBplHeH3DUmQkT7XX1TqaiFiSsqKq1JiNq4ersOMVLd38Zfu6kh67AZR5O3USRpUzwG
FfKfyyGEGGTUB3kyA456r0uJgKJCPX24UIBsQhc+oYVxeIDCtdVWBmNgegsAkjDLQQgrVA7ZwrzF
2vvDun/SzzCQVzQdfTX9H9RjzYZGv/dJhbY/BgAUWhxPMHEA+RhScioifvovdFRbAPktAKtbjfqS
0a4/u9i4BtiU2jRCb/WGEhvkRwTLQ5ee21aQYvtdgxK8wpdX2bwnw207TidOmEkkmUtXkw78m0oM
l4x5N18gsG6VGi6IHqHVIbR1yICO9z4e4OD88R7p2DxJ38WTlg1YeVKgP6x1PJH/zMJx3DJufbhd
lFbxpwbyEy+BlSuKaUPcGivw+rIf9QQBB1IpksKTVLjENAKLeSg2s0P1iKUpyNmnz1bjrdzSYByH
2QgTU6SYfQL93wFx1yAVhdqozEizvqMaF7/AsnqtU7r+wCbK4fxst2/rZWDY7JUW9d//4OZeSPmR
HUfVrUZgoRUeOCYOqScqyg1WQhhgMXko6FhS7RQ7zgB2ilyO0U+uVA/aOIoKntFMD91LyMaoH64I
e0CNP/bTTJvfC/LWNZ/GNWTpbWityBZYSmMade+vqxoTJ2CkUPeP6LNunAkytcLhsnuMMgNkSZIx
mcJ258NwTifQV06rx3w7ydaXlGJMhf2n+VKaFTly3/HT+RoXBvvDk5YbumsfZKpNY1jyUo0eb/zf
8UsQopk0+FS++Xfcb1O6Uhz00uVAhMO85ybLKPawYPPxt4MIy58SbBdMOGxG+pctz7mbrezMUHgO
qTdKpQtfxWwk0yWyvs3nnmGAcaqKWl6GyFgChM00vyByD4Ucz1+2EdY8RfrM/FrYHsxm8a6JVYxq
jIvJmfJiwkrcOpX/h7XYiqYT6hJ23iuHoIgWKayuxZhuDhZ9ZrfH7R9G3CHI8x287q45Iv34xeZH
EHs5OJvlttEJfSfZNZ8GyUuOHuQX4Whj/MkBwcDSa5eLrifRwSClGpxfjAj3qfKzLwffBC2L6gRG
s7xBMGHwr0Y+B/hbhlDnEEO0HPgncoCbjZlq3bftnw6rFOIhPAzNiBUbD41CTn1AciUfuwYJHqQY
r+xI9IjK1N4wvoot1eOfFhWkUHJvO0TqWPL0inewAhTXesRlTsnYAPpKMZUroDnzwD/3uPkIscgd
85+aQ8XE8tmjUW99XQvpGwwp7687JKeuzZ8AonqmBZfUbJlYTrLQM9FNw/cWe/oa8l0qDc8NeurC
0PhaAJCkuSvCIGQ41I9Wyw6UXzFjiiMeWyUUBgfmTKOER3mxhs7P0S1Gm3AxxGrxRZ6RlpMNWbqX
p8qreM1Ryzpts27xfW9qN9KSxV6f+CtfTTAt+dpNY8umO9toR0mcGVCQnGszqItlF+uUoxHbZ1st
J3TIxf/9wyvcmXsCGAnaXUNmGImKCVKnXW7QIw6TV3kXdCzNRIqWMKI4HoVKgO2KGl0W3RrOL4dL
V8Dp3T4QiMhi7gD5Z1/fs1df2u321/8FISpqzxVf8DuuNllI85k7tGBxGkW9EU4ly8sSeRymXKLx
0ctWd5lZxQi1e/qLz1Wd2RoGg3ooFocBrn9fgqb0t85FVl9V26CaVZi9aU6SMAVzYJjbGDxKLDn1
koFfy2EggRUV9ULRYD4GioaqrR+94wnrTRcpHo1NUhV9L1ad9aF4WkZVpBVywF944MPeU5CwxFBa
b7REHHDU20kQLAgce/s4sNcHnDmBkDigbtE8D2ANmB8s9uKXNp3yRJWgAoMc3BD4VXAe47MvwAra
0JMrMV6loHHulzw98A0Q6clERQDZI12bx18bBIJ5tx1zCZYaXISOyfVLINWnsAhS8RjoRgQsYt3s
LR2src+CcQMSoDBKO48yqPeteDYYju2Rx2Gi+xvM8GJwInEKA01pkXbm1nfcjJ6bHMkHV+uE06JU
ua277EiA1P9/9FGhMfGllQauEvlRX3OC/VQcALn08HS5IovtKHX5AXQ8SrmvM7SyuvFr/7mj2OJT
yhgQhU9AHNoKApLw9ckWpoFXvfi7Ia8B6onukDUOyQBBxaHsp+cPvJyehF79/Eci48OPyWYuE4hr
O3w+MVnod0BPXtKgBJM3fcDQJ63hejWptYw5LVOWdAEizPbgUkM+x93UfMihhd9+vakzWbqXBpLM
NWopH/+5+60B7Zgco4ogETbc9gFNWGfYQnB3SDlU6otzjIG5DdfjKePmmvY55vuqoAL4AFNlhdBM
K8rcVHZ7ol2rxGDKeGeXkQrWLD0+SLCLvdLCJlA+np22jUopz0Q9sS4IxenOlOA/Z4tgJdrZ2cOE
8RodFMXbLd6XImlt/QstvdXUn3IFzWhbntw7k/Ri7c7vpLbyI6707djDOvwXpI1L9kPE/OHc1uJC
b82WO3lIUzpHGFDJoeEME5evroMfUinZtFVnp4Ey7BG3w9Nw71oZjvuPFRnlzmZvWSWIzapF70ub
NrCdCmCazRcUb083E+2aNvqpltx6Vz9Wp1fZXj2AATz5/zYdpKfIbC9W6GEswjMVaooi8JxJ2zJU
vRv9Oxvz9vxyTUmnDO3xCxo/Vs09BqD+vLNwHiVcfH+HgqhXueoaBgkZnrYMTMYV/YFqQwdDc5Tx
dH9OFyp7Bew8PyUOc6Uk1yiOxPG3RFIQPvTOYxqs3VhkQ3eArGHwBQQb8wt+Ff+445LB9Ny2mch0
2vAtsjSs1G9u/SKwWDwDc6B2aMVD/Hf/FJEIgd5lc4mJt2GpUaSZmrIse0k7m/JAS+3+qDEKxjeq
H2+ySW1IdxzCt1jUlOGgVg0uS3If1DuZncyEOPbkkrrzgQTKL7rYHpK2XFg9Vx0feg21hJHDzK2M
w+180U7flHqITvmVEDqYrrAR8GSgKpwIAMZbZszSFUAtrobq87yBjInkNrqZ/DCkUeGyeG5L4sFC
PfxzdW0PGaJX3H45iECubJeyb70QuhoaMNQWN7apaaqgCDrmbmKdwZ59AOoPEP+uzGGIEnGMhwda
B2KirQjNux53/BB3/FC6wxTue5HRzCeOxsZxHUFeZDNbrkgBotti/QdLGZ27+MdGnNOxeOBtF02U
XlLqlc6pc4Jn5oae6BTNsmqbxbcR3uTMr6AzRm3Il7l5cvThi6DKom8GjG+TESb4InP227GTzCJD
LDFzTvE1Hi23W14svFpZvMVjAH36QDWFb4ZWNt0rDoMoKlzx23dXaMgDSvCwS/f7umi4z/3h0Nl9
/AXxw9GynBp78W+6gct1nD3GXW25WzJ7dIx58bQy1OLNMzb59DNdGut6gc3nApwdgQV/Qn7TLPZ0
2mSr0SOYXFxr2rDoFnmphSIzjC+o6CSfrhIZ6WIw8NMTzVFI5RuPNlUj7+vfHZtteF82ibcupvN3
CsD7N1Jg/0qwBtPw0AI1EcNlPgplFZf0EAuX1H45jqd8gpgu72BMZ8YL9caxTm0zMUFsyJsekJCf
zan1mQl6Kdr6bpIXTlWSEo4TS6hiVtvcESX5Ifl0N474vtelo2Tskwi1htWytb05/X0VPLhNc4Gx
XYEV6vnO80v/QCG+EyWoZG5NpCGuk0Nh5IbJUIC01Hs979I6pJm3FKj7Q9Yo49JD+fmulTLu7zz9
uaZSe+mGvqXgNcOtjBbh9Bk/YHWLN6OVQgE9k/6SiOVw62glVrnkZoX/c+O99UoVIYXnQu37kkib
5IqlolrGIqgBb3QjqAq1ElxiSgY9K1TJuyOCMGIQeyGW4uNrH4ChGJ5Z4P9gLAkrn+skLLPJPDYP
WH9QRU+6LZxX6CkM2FkKV2+RbGWCRa2ZWZDGHE9NVfg++xoeSIWySTJsoR2VajO5QCSRXd9QaS1T
XorF9483wtbbeOhrJ4QfjIzAwm+QuRFAEmjSb0hRY3DYGtjaRme4eHJgrXEDOTk3u5sST4Gfn3Io
Dx1IJW1elp8/aWrsYWNOzlFyOenqqyjGguJjt43NvVHqejjiBzXEtjeWsszxjUuvJgsHeyEba7n/
B0s4kwPSzoWiydd/bmPwXharv4vBBPVFDe3ifohGq/VNJ8Q47G6ck17O78EfO02HACNL56kdbjAq
t35AAF5rQTbju1twlY8/rchIeuyhMkKkNu1qTz0ArLek3JA3ws2bDESIuFG5QHWInx/RbqvPL56v
pm0aZ1iFlznmz6+09vWqCf/2bCqzaooZzxCkKUwAcrR21XrDND7pSxtgagrZGgSORSK4M/P35X2e
WIobGYTtO0j1Ysgd0HWzUu29a5Rl5ZEh+Kpzz9YENpOoD63kn9YBwVkmqlUomaIV3iHEFBT7OkAl
MFrOhnz+grZDZC8ug/6pEiQi9t/XmTnVkIw927kWs827v56DaMbScqiuDJKNIxpF69ZuMDezZtRZ
iM/iwr1V+xfp8tCKZYtS/1GyhpidW7xFsZjhTgHzD5dRJVJh/BCzlNJa1VxcAxxeb5nD5aLMPtAK
DIfiU/W0VTAfBJ+sVL//Usda08kR7bO83xrteZWluwMcpUHN2e37pfMqf81uSyWyzmuWE1SVj2Kz
AM/31My6kcZhd3sZqyNYJjb57aB61PAOyMdQweg/ZqSK8Tnur3inL3Br9a3IYUNnOndO4rGkRDtS
T5HpErGK9ZeDgd8UiaKX7T4cOBExS8A+FIqRsJS7VznkaVM2L8OYyTscT03iqe3IR2n/g1GILHsh
jhftVNSIjpz8Mcx5ZzsQWAL2aIPb/8S0+XbbkKozgIUMRTHTZ9Z+BppaNiCCLLyIpVJFNzNiGdgA
j0BZaEH+mG2G5oXqNUWzLFMwxJ9CLS6/E5/KhgHW0ppFjH5QhmTt0+g/IMNZkfKeq4mpc3LX10OI
X37207xYf6k20XnBey3XuVEb9+FRL3Pu0ahh2I8+75ukLYjxeXFyx/1zlk0uHZpfT9bNxyAlWrpG
Hkj5piwpUKsTADE9PPocUTcpsGZknHQ5WzjinTjUCddfAklhVgHEIY/qnXXVR87/nlW1EPnoQFSq
jg5K473x7Rt5OTCHkL7V/YnsW33RTeMwTRNlzFYn83dfUG+eEYU9QTWm8/t6gv8ma5s6acPIQ0/7
xbnEKzTdQIWEO55FbyQAz6AIMe2t0miGbqL6MqaNqfZLqbWvEvswPRLDj+tBXb/9qlTaIkuj6f5i
yo3rvvmD1cs6YxPnTxYTFJNJasBoAaDBrKq/dRQQOmu9pSahdRK+gf0vbg67V/pY95umDIsrjoSk
S+POy6IeTrIfjBy1qOtA3di9s6JHdmC9g2tY0T+F81C0Kxs5ZzuTn8W+XwvCs23GJmRshpLsDYUy
4usM5FQX5Ms2pnSp9RKfvDDzQRATHtn+EFUxRrpBZy5y8a7fym03ITaAxlv+iHSNqaksUafLT/PL
oyd69v0KD3/4/Hvs+AQu2nrcbDh34eKPhpuAckXRSz9jgj5lDaIm7rPeX4xBTpQ03rKGzjX+coBO
n0nFZ5I12NqYhpjTZglvq8AWNZr2ps6HWsB0R7b9soVypO+viDpUaRviW7DaMfAmS6ioYporMNzH
gDoWhrDpJyQVztymWbpnKWp6KergdkbDWRK+UJ0yE0f24MF5164oauacT9MV9dIPzBJtNtQEskpN
cQbHBEjgBZYLsaE7TERxnfqBY1KOli9bVCWkHRxIhNMMPVfNpROGhDRshp2YRWsI7uQJGLic4FZ0
5pHUcnWzFoNBzpg9fvJs3+yUx3+biugpDM72m4X/q/1vFqPtdazMXjAQtyF7LXxDq17TV62NrrEw
O7TTn63iIUgQCBTd2uNcMb7I0s8dao4ctiuKZZ4vh6Umkt+F6PKlzTwdm5vKyRDRU26lYleiVRuc
5GzsA6kvVhrhVy3oRE5rQ8fOlJN8xU8rPjcMd0duvGcfg9v+DMiGpo53EuXss0Ifs2ACR79ClW+0
zul+u5zdOxEtI1hbA+FdyzgLZJV3vdrgLzk4VBD0xCSre+QZvzZ5AGYc17Hm9WT3UfHYHpbxpL9t
CFOBwzfKxXbDsz4HRtpHd2jOGaFnprrrTPryaytxBeMrnT2NEXcsLeAdq8iKim10rFsHfsGylXUi
KZ68tsJGrMrx3p9ffeKFKv6MzS1bbK1elP+Q1qeILBUe8A8btVtKlcvkqYZrmj/sPr0Q8fdWi4nc
p/5uIsK0lB3/hts8LY40tpBFR35cb/JXlW8qN+SL33FOw5YwdBYo78OQSvI54qTXKXrpxAomMXWM
OrayzbeS1qC8D9ED0zqdAJ3ZCMCBTiSwpV9J6ZRanKlMn02qOEEjsT945v+mfPGiPm5kl+L1Ink9
xpPTkBXWQLAxx28TuaLgpAcg26ihZhKbKR6jZCBANVCw8b4gd7NWpHm0DY798IAIIumywjr2IJI2
7oWkMSq5wgtKY6JIYKnU1q3pb8Qhg+esYYOwW+05pngXpr8ISBFLdQg/zi513ALWI0GsXBWuu2eT
qK9QSNRFIyR9hkC7FCr4F3//LXV2TNVs75EtKeTSD8DbV83lEV3hB0TMRxv9n8d5abXtwxuwh9jE
FGUpAy6gbXV8yyAhmi17srkHCilm1xP61k+kg9abDcQr+TEqePw+SF8Ug6PT5kM2/TUgmwZkCeHf
+AG11PV5fq1JsA8WpAbkcVXQrLqxATyVJGSJyNuGZmuuZY3HDM0JseAWvphuZzYSOoLqpfiU+3sr
SVOjt2UlGCUsWUeHrrVMXMNlHqodhFE4e5YUampIHQoj1YAeHTclj0g7nLuHaDuPr4a5rhSP2mUD
RwQakMOHVIjIiN+T/d+U/GkzRwZvUx9AFVjJN4rJJkTMdEJh1t9o23xaGlg3uSO/0bek152oi3vR
BpOsSBGWINMIr1Ok1YQOqLhu2pJzQsRk5L+L2pAN0KtEfv+zU/Rfkoq+mIYRU+Uc4L81wWdTHVv+
IAzDKmu8qX8gNchan+QRgieCOIdc27suGe6cN2IHwmtJ2tz2aAxI/XKS/pK2E+jlajltVwhEWxNn
/lnFwZqTkA2g5CgRjn1gVRq8hVHyAIyTLcJ6ieHgjd7Z+Ry4UeufrK5uRVCtODwht0HXA31oWqm+
1pT3TChVw1NTS7eQliWLW9KQUkXa9tsHTXF9c0PE8YvX58BB3p0JmweXZvitokB1xu4YG2izVEtB
dEBy0VvYUqCJgMGeZ59lPrMLgbG7BXX39nqk3gjXPUg+wdLYfYGw17thusQq4Nk/t2I61DPb1r4W
+KHMO48dL0aHIx6l3wMo2ocYkdf9ywhwgKZNt5uYXzZJsAc3w+nJ5RS8hSyz991ohmEMZeYpEr65
p5PrKoNtYIkBzWkMuIi76CbpFwMI7I1MPt2sJ+OSYPwxRnYcJr5QbtWD+77r9mfodSF6QY6NrmJs
+Sqf7FAwY7YNeh9WpoQM7GTnIMVbN8lLjhJm3evyKE+JHv7TnI3TLQpX5uQPSQ+Q4oOomNVfb35W
OlQZxdq28gMcjJ4YqmvhYBznfpNrBViooRrIHR6XBgEV9zKPrrIC8kA7Cicsc/3UKLTu+JGDOrup
gsh1OuLVrHBlSEHZE9ShxUjSOccR6yybW/XFZi3IB6CCkZNYIx7l7X7DAkd1JnecOLd7IGvkydbq
jhXOIbw6+bPUFUa4HnuflKrCNDOwhhDPCHKVUiXFyrCmxuAAuU64lnVRVttvLYNSPv9vaodtnR4a
pxTgBeeKjzKENLtbFUfst5KJX50HL1XtBOLi2u1UkVwSS+w6SHeykxVWpL0CJX4XCsJYdvsS9/b3
KLxta4eeBRiE0bOzmJqEhqs+HbqmvPHhpiyJHnex+v3lQjdZFqAm7zUMKgmHqZjeEqFI8jdOQsGp
w7u5yCIS+a+IdyyuI31jXu+OFmdYVK5GBb60YIAflaSKMjugfe2LKuYnP5Y8SIiV0mzmK5QwuWFY
7CJFX3WjPP7+1PVduUOQAif/HWICLtuLOeekxGi4Z18CyGzdmQ/zV26Ryu8mlfWCuBAxvKKnBkWK
zOJ8A7eNHD4gJse9yLV2FIyU0LleUBCUkA04z46ZYYe6upyLnukuhFakxNXKpeg0bH3R+LkapKO1
VAlAJMCxGlNCYkMD1UcaGp62QBEC094xdMI1yIMWXw2viPbk1cWQBRZVVm5w6T1GafKRnfE/SLFc
MoSv4sYcAcZagVp8oHvZlGwkscdIxj3Bip9/kPbwyJYj8SYOpvo3BvSBKR/mA0yOm1QERUWm78NQ
P0OQza200Hz7nU8TwnmHX7Dd19LXkj0RNnefXIaOQvjrXcsOAzURw3M7NPHh3jKderfkCJPAQMQe
YlB5mDgo52ygm9Icks3/SgVXYEI7dZM+hACkuXeMKHJaWEUqI6BjN5D+xp9j0tMUdIYC/c0SpMQg
1FOc9vpXWPAbK4cDsT1PxnQSDabwziE5GM6WxqQ36s0/cgRWmJFc0B5Syybn7/OEi18Vx2z1bY0f
PpQhCcJrk2aB9uHwmzgkvXT+tFU4J1lBGAxtXSaHs7Y+2+H36NvGQIXRQB0rhB0uJoP63n2ZZds4
vnivtiZbposAr+Va08cVz+o8CeCDeYWyycpTRqzxmpuueVk2eaUcyJgHocBDjI895a5y7SNf8Pll
QGcQJfQCvOUhfiop05c1jWR759+NPSw6ZdLtND5WAt5eQL0DcX5rNt0yAIDA8Gktjv9JvkHUR8Lm
Ofqj6Wzrz7idNNG6qKHrWF8mVOcNA+lpj/BjSoapR2CxsrTjnn2ZP3ntBNQxEbUJ5+6UHUFuxUuV
t/Y3++kbJbrsFGgkhNvzznt9QddL/5+b7/hvbvRwoRokJBA9zlNMiRtl/yW0EymzRyZ4u5oYP8Hi
zCYsYwIBo3yYSZVREd1Kj7U9ppwv58qgU30c9Q4by0ZsCDmiSBafJkXT34wxPC1po4NeFFQkTs8M
6wddtoYWqU2kQqrBtxGasS98jap93I7pO69X+s4Q7CfNYkxUKZv+DDfyIssFdGu16E8tGhvATO57
w8w+oEleOLgixO0fLzQspORQbiyh45uiQbdAdYiiOF8a+4yr1ur/c8M363/GjOH2syuYCBl7xgpQ
lFqiNVXarCJFRAXkfWIDi3NeIBcBGnUGgisFFaasku+nI3MpEbI9XQKXBdZTGKxmJxyknQSnXJeV
hi8SfDPCeGg+JvcCaZdse1XPg1SaJ5UEm9YWJ7ADA200avaqrJ0F0xe9NK0u0B6N8L57bP6RLRSK
qdGQFu30w/jeaZsmUixr+ROWTFWVdU0tNtiLBSP/CagnY8mO7e1yJsAdHROZRZ8YWXF6vXbq/TaB
UxTCmebiwYM/SFCat/cG/mkM0kLfGBR3J8odtr3AvYg781d0pa+avcSl8IBpnmXtnKYCB/3O6GwG
+fxE1xTY88/4P2BtZNHtF5eXsm3bPvDFvXQ5OSpa0zNqML0iTNnirwdGfnUBVivZSgo+kFAZSV6k
GM0b1mhZzUdFbfnP9PZqaH173tR8nM0Kq72Z2uJVfsftZn6gI9gjX0n+m71WUY7pTAA2CulhAokg
Y0LwCNPXV4sULhtj7rUtBetXDw0JbMtDOxCRICuQ0ITkYH16e3W4iJu/RW8cfrzUyOzAF/4dIi8G
6RxzaJ6/v+RDzrkN+8jaA6z0acIbqI/0AeYOjpAYI10q1KMAiw9jRDXXOPxBuwxOUdFC6zJPOpbz
Z0B3SKUCVSGMXSDZwGY+Ef21RHK2acb+z8oczL/jF3F4dpMLZBK5Y1HhUsJwWsPKaBOBlegijCLa
REKPB5isPBOoio6pMXbOFWv7b/eQd3DqP78LjPoBNcHlILGw00sh5uuVWurH2DxdoUB3ed3fMT6m
3YOVKONZGCb3rkm34OqFNwvVYSyvXGCsfAmPHlpyoZjJtm4T9CZOCQKyg840yjfI+tARNMgYI9QH
ukYNnzkSj5hvwV1k3gbycxh+DE5SkRoHnfwD8OsYNPPRFjtdGryF3HZRWYLlDBbofOm3SVFg1ocj
gqq/KST1Zqm7HttRlgnyTTJC/9Tfj7wkqlgxDdGUgemddBWTEsgOCiAICciqzX25uSyoeiV+rFC2
Fm6Nm5eiPA2SzkQlMGXGL3X3uSs6bViBjOQOwg+I7d8Rst+kUgbYCVkFZSoJ6aW3vDvzyK9SKc8p
K9Libg326f1D05UanKoENKxLjdlIQKXeTXe6EUuG6qoUZxs68R0XbcjBs0+js8jBvtoYFxbwLu3M
0v3fgk2nkZjWpLvl2Vc8alkKWGfxYLtPaX0cK5OKLaulj1CK0ukSMEWuFwRinVfp1h3CTeFljQX6
19FGHweFvzSEB3PVrwQA4nstk2OdvXng8iZLQ5UZWswntshSfKDlRKcjnrShyd9CldgR6qn+jljb
i6fsGP3x4WbJrb4Cr1soNWTh1iDIOU+zC2E0aq3Qc0w3E4/xoU7rWObbj2DkvWlkFoB4Qyxr13ix
h89dkxYiiWOx6mBMM9Hcwb64gAplK2/faReYUNay4PBYS9eQDQQ+E0AVu1a+LFJ/V+xwpws68po1
xhv2mO84Z/XT8X48riRM2RuIGdlLrBh9s4cjS/vmHj7CWCfGBxzhm9QnWk0rkQIKpfS+tBMkXO79
ZwCt/XHdjCvPHLg1LbynCCPOyri8jr3/Lb1w6NglPShHaxTylBqhkQ7Ocli/zriesYpF8tfTmqKc
ZF0wogozWpv8vLbpM+BKM35CjQnkwFoPXCGT09tsI6MAYSJvB3Ewf+Y7y3myL8n1Gn5E2CquxU0I
68qHbnZiJvKhUwlUe+UCu7XuCGhjZh26SeoRC8h2OLxz4bKfiTZLckH78EtKBbqFr/QzPame9eAW
3ZxQM0RMwrm5sL3WRqG/txhtEQB+rFx0bSrfhzkc4FjGIYMPDTzKfLzIJXWSEadZnQ7xdaMlD+Cx
rpWJxypD/WsW0CmPD8y4dBBUBey80TX10rbpqOmLdJH8+RF2+y2Fhqswc34aa2blOqayXKoJql78
rL0DiBFprSaOIXQOgcdMF9KIxiSYFFyH8XILkVGnDTLHi2/tIoQUvZF5KAaMicu2G2C50D/uuPlC
w2MHGP8l0g5omhJsQk6Caf7DBrERwuWbNHjc9fLZr/eHnnHcpemiZsfbnS8Y9UB2T49PYFPjCkd6
JzplqR3CiCGFr8cNE8HMEjrlEQHs5mDCSjvVmFoJ1T7fH7CtrAR5pTs3ujKEn9La0DGNGAwD7/UL
p/hxHsCZw6LcZ1bVCL7hXFGd9JmLOUzA61zNOW0WEgyi6MSKtcdZANMPbGD8x+/peeMJJLXKO7Ap
tEmZsLDKx5Gn/1k9xhdiS57wdfflIiWLjMNdcXkyyANx+hsJcer8JdzzUSRk5N41kqvWQD/0QuMc
nPAsGj81nvdOxi6GM8S6xlyALvXRhvbXZ4rbXht9gVqfq5u8iorIcQP0LYTn9e/ZvhpMcdVNf/Ve
B9/0/yzCUYumDuIngRMMmSnC1FhtK8I/CE1/c6YhTBuWk6h7P5dlyy7VyGxAPLfnsY7UVP+cPuAz
FDLDl4FQSk3JfbfFYtCxsV6f3jOsmMJ9ezrk9U8WD53NfyTlUh/RdNLdZkYGIyYO/UJ5OjV9P5UY
ib1VYLt850qNkWnxMwtbeZVjnGPc+BBTeCBE8bigS0NSyyGswRlK1mQqtmSm76XAhpotiKUkOtix
TSzw5FAwOFAuJLEpsLQt+jEREHo4BWfu6eC2Hm71BJGct8hshGMZ5LDHtAiiWbt+/E9izHFuav02
yDL0xvSFz9NA4BFgBDOSfkvLIuCwzH8P7lbTxhDt39REZtH6AE41u32kH9w8wpSnxTQ+XOjq4Pxj
wWVf2e+3sNeI7ZurR83HOj+lHaQ1jqvQIX6TkPh+6JdkOn4TehChFz1tG8YO1c70vrFjFuZmWNwo
Pnqw0XbT2FkM7DRB3y4iXpcqrbQaWV2n5QRhVuFooQsArnS5YY7l1xRu2H8pb4a+hNaNHZrwQvTI
C85ShTwzmh9gozpuU6wjoIail9MHTkVnPFoowG6NsBilfqrzQMYyHCjHj/ahiLJ6Wkfa3rI17FKm
hwNfNGnpSGid0rH6gyCqdQHhGRgKHqfO1tmKsSQYHHS/2Cv5UYRdXShzmnCShcMYm/xDJ3ziBUyk
28tL0o6X2SB43fJtQzoYtT/+pnQat0SqRfgNVdn4VDG6nO0mB4vWSwxwmn0M8B9frizkN55pBA2P
yuzOUgXYU7bwiQv8fq2M1+H61jSUbYX/TsCNjqrURCVNH588ynBM+jEIekM4/NHD97BDfSnGB5hr
B049mwiTgL3ro5xiaXbCcTyv6M7XvJPm3tnBAeF1sl9zZ0jsjiyMjmUUTxbnfGarVyL8kBfmVf+Y
r86GdysQquiQ0aRAXhmaVzTVu5bwp3dk01w2YuErk7gHdanTMr1D7vqp65SNQs1cb+KFdEeZUEEr
UPVDKTrRCSIptVe5UWftj6BOmBEuzMJCR4tiqJ8PYvoQJp0cRkohFp3iD/B9DnpIq/xrjv2fFTGG
wmtWJpVk93p0p+F+wi1JVljvJ5FaugZRO5QzNlfxL0P6zCd19A6YkKJHq1ZGjXFqRZn5Tj6j2VYH
7gHUFqDc63ixW0zBnlqEkYnNHMdyU5pvg15Vka4Wgc2xDgthrggiCCvTmFh9IK+yB7Mj4NcRicMQ
+aJUtjWetU98rxcr1RJMQzKJdb1PsQBbR9UInlQiAQkaVi+oNFIGseLan1VLz91AaegpHYeG1Pjd
sLIgkmYaDJ5EOwTH6Yti9ML9SBvpTGZI8/bwdKhyVxxwFUenAfyzYck4e9c0Imfr7lpilvjLs1Z9
Pjb97ou6tF5zF4AZYPboEQopF9/tsX1MHsTRo7DNKJ6cWCde0qFcovy96ggCuJUzqTdPh2XXu+hQ
NLxjtzMmhWayz/R0mJOiSj6aQFJdz7W24BMGjc7eTVO6VDz5TS70PZ5oZcn6GClknWvRFfQ+8Gfn
YKidysybP0abuMj+sHpgzZVm4S0YcbYvrvuant68NGiktf8UK33+hAKG8EVNE/7VuSdPoCRguaC7
8bcxiE16pKa7RD2t2E+Z2YWEuKo/L14IeAL1C8YT3xm9XY+NcJJP8EbkmAg7ofItF6qESjrTq1Rn
6lkw6Xh2Ldu3EFi23wfkvh3NWbAE72aS9Pjav88RATg+dP4Gt3cHJ02Astox8qP8UX983jwAUgqa
A21CsBDixubDgzMdORurC6JGAoN576QdF16aUH2/HLqu7T4pI58g4A+tguFX6KOT1TRg1oF3MLom
lst7bwx+s+jzw6uMb7hzBUjSAcmVw9hxMv2Xp7LKN97sd+6kk0Ag7JI+v7Gxo+tqDLMk6GhTAstc
4+C11o8D/a81pfg9XNxOgMBsQAb9U/buHXTd7DiIwQzf+2BAVChSuio4s8vIA3Ig72Nal04SqAqk
Y5ounxlzVKEhJIP8IwiifIsiCtY5FlR5PWRnqf0S/Aj0IfS6TWKhAASvVpuqBLz0foHqDHr+Infb
7/Tnxbkp9rVvYfCnFL3RzMgwr1sCtx3k5mAdI0QeFslp+pwlGichNGMTdKiJZpeQwYOv/J0X0BJT
tu96q09/JGBXMsV0Tf1Cv7la23x6q00M2PcaZ+bgi3vjW4Tmvb9QoiGcsVT5k9k/hD+eFXnwliaE
o3pizKiYx61cgU5q8GGoYGylbPDemjMB3iXbO5qD6UtGrOPOsmoLi03/NMNpVHC9BT8AdCcb1Nlm
qxfXjN41YvhnJ42IB/d7WddcaPzQQtSDQmp6ccul7EPGPRU1YMvGZfRtoqDrh9SYLrCH0YczCtCI
oSCFph9UJgg40GMdiQPqR4KWOUJPjjmVOgOX645TQhgeuv1N+pMQQ5UTtIunP8uKH0srj4xYbKpi
Mu4xZAw7PnKO2cl04oB3/+AlCcWCN+UnlH8PMBgBt98Rj4TXrOxF0WiVliYltcFyGRGg6ab775we
3eSIx9QzbeZU3U2GYYMEHXQm5CDuEv8/vy7nXuyy5lIg8LhY9T7+d6splGaLJVz8JIN1O3m+HRq9
mDCsqtuO3/XDNUgDVNHm4QfdYyILxWGBz4RRlrVMj6BUZ63Ry9q+ICasPh3lhrn6wgEj6O0PMBMj
OVP4G7Ug299Ws8fiNhdSw7H4s49T2xYq+FDVmi84lgLMjexhPdo/+hPYYwdJ6O4G71lWC4iFb/jr
7s4MizGJDzWDODf3Zb+azLYC04I+nzgRLs+q1ejNoUa1tDFcxosZy7Zk3X69+ylOdLlL/mNhFuyA
uYPJQtRvGqt1EG5Xg3xNLpiLBxDjuVQd/8yuqAH7mX5AUOH54y0aT5nzvh2QHNQDI9OZrlnZpSJN
MLkqUf0ZdNF+51F/Ccz0XWYid/yvtp5jmN9884yKTWTyZd8Jia2P4vg5xva9ub1VDg0/SDh0dVj5
YEtN/5VKDyF74EgP1/cgHlrgkWwkgqe5kWovr/MBR7aWhtA3lwRPh7Fm0q2/JWTnOMuwMZwP3cyD
KG9FhPWB1KY0IO8ElQ98gaNTOT7o+/XxbTG1OWdzodFApMoSgKrfjkLPCQRnl5tl3G2zXsikIg/3
ivBVdMHx+9iJoJSqmmjlXsdX4tLHSZx34Jy6ZRFr36cAQv2pd0N3nfDxtSy6uYZzFi2wcUxrBuh5
Ux/DCL6KKVjOO/ZSaqqE6VzheZxiJNclCTDkpOOpR2OlFdIw0WPfLeoqZ+bsZD9uL0Fe/pN8yzaj
oNMVEX+H2I9dhs1Z+6rxWqWrSCGZYR734vSKY24nOk8bFdie8c0Cv9z2gJaYWW5JuP/EYjaWW04T
sreIyUGoiDl/PAo1BRrP6fU4+512oDikoMTKZOohefNBGlsJT3YZ2OU3GJz1Hqsb8edcY5+h6KWL
8WlNptFUxxfwDKbHYVNwP4K6bA5r3s67vzTPTcEA895nGEESjGj35qnN67+akTE6mkiVeH20T/N/
+v9yjtRxTzSCf3TGnVcGrCliDUWxCRN89bHeVgkjrKdjgxCTqxOBEIadlUt474z6PHcmxznNZUQg
4kLvfzpDRR5PTG/9qeoZ3m2iI60oJTxrvvTE86tVv8S+Uz8cl2xgN1Ak1Lcave47IUF9MzrWy/qq
lZLvE69PtgewHngjU32pvgam7Bcwm+EwnxVaO5SO/RPHE+795FPR/oGQsSYfHnIpwnTby97FLnIT
cSC7tOzFYDIa1BBQFk6GnV9RHxUiVgYl0ERINFtBX8aqJ3nsBvh3yVK3vrAPAknYQ5lY0FY+JcTk
KPdwZt4ADVBIIvwFvKhhpww2NDjjRDiVDcB3PA8TkgxVFF6ZArnyLe7BxDC2jpLXz6mi0KEXdSsi
lT4xoShfwQfts7JhVjuZih5muuhN+tylQMKFYmhT20mjMt+4G22Alb2C2sA1VN1ZtsgUsDaKbDte
lgwEs8au4cBs355hNV02k12u6aOnqD5/qL6uz3xlKrXW/t0H8W999W0k4Cr4TrQVQZomZKumSoGE
4q64gPbepAdaydqG3DGSivRAuNNjq82xTIiaydBQutL5/8T89q3GN6yH48EDsegpWs/Lh7na2Mij
6z5CpUl7rgogcuQ7IbJ8kynJsfRwQ2XzKG80Dt9bJVeFeSiCcTbbEBTo2QxH7f3hS9CP6mKWz4HW
MkBn1f9cGs2ma+4XTivfxwuVwCcFUWBgo2fH87vUPg72Y6Vl+lJ+9sohp1CwhP/5pLjUQkVOfsOo
RWBwXGqsV+cu8o0KapXz6nU8sofuz9ZyOYrqsXx34O1oiQ4lONz8/UYoFdZSsVAb3vT+abnSprOZ
47PsgwJt0kd9CqaUPq/pq/qWq/h6iGoKlEViYID4bDIVn23R1+4QzTRQcgTi8Wuz17NOzVrjA1r9
t0ogzyiFF6lBIxVxAFNfXIigDyk8cuExD4wtIq95fROAq/dz4Sb/WsQiJ2QA51Hio0sojRAFRKeX
8glmnu4uPMuRhxCo3dyE7rPdud8WoI0ZR8YGU/mquzT4vhOr/qT12vNJixB64eYbE5zdvbfnbGQx
DAIRAZHR3VD6hL87DSTpsf7GclaSA0F3qTQ5uJFataZB8YZTQpmmTv9eDFrbOEfv6WmzNnPPZHcu
kviUZNYJb2nn+vDdSOuZcGMUykNx5RP9PHny63vG9oP8G0oBBx8h1OvVdmv609VOEXJrJzMjXQ+i
j/ibdEx7kmu+ZNSoQA8NH+mp54ZpYXX3fYP0WR8qm/cSiaP78VHZCMpuAlGVjJTvg5aoW1Ri5UeZ
sicoBUxq388QnDUetvdn2uU5AUdzZZNRJanIp+72FO/K2qd5HoX93lRDy2Rgsy6bFAKy1H9yU8Xx
8poVG1NtlDixG0Q0v3ENy4g1qqpcPsR2y4fHRB7smYfTcWoaJEpHLKcbxAM3mGEeyBFo+Y3YCWPA
cWpqXFhIsDm9pFBd5jfNkBUVqy0t63SNupsqQ13Qou8eZfrG2ibT3ExVUod5ddlhhKAGmxb4g7+X
28MsvgYLg6bdllsYCNTRr/NqKf2KxCKrc/GqFQXInL6kmSXjZFO6hh0HggBmga9WuFqAoTY8AaGD
X3hjJ4+5v+/DPQ23K2QKSm15faag1kZPDcinzwJV2TD/HKbRjLq6ZSYH34EYjw0sHpxYkU2/AeOA
iUzcUkiHjvv10pKVC/c7/DM8jcflYHUlCgZH624ZgJoERV70xUE1u8jxwsiYKdGHt9YXsTErJwlE
S5eGY/BsFMANzA5NinqMYwZ7WGa8nKdGbaAwmxPtpofoqAWiKXovvaqgvHtDJjf3CCb6eIN0DuMv
7ClrhjrRDk5ceLtHVPJd8KCA2oYwN+QK4tExOJOhe7GB61BLaNUkdowOAgQgCE4djZOCcT4nNeF1
zj3oCXNLjfYrwzx40ESZbD4E4+ZfxiW3ZlWSKaNZvu6FvDYIbHRqqi6begXZtZg/ZEGiyQ5FR4z4
OMciy3aURcKU7/EB3rzFgHU5ovfjqthRhBoiL3FVAxJHWoAyfsFmZujn0TbjcA6RV6OUlKl2s3DI
IwIIJ7/Z7p0CquS7zUVOORuKEDjxinxIu2FDaN40unjtZ4U3OxkCX0x0wcsvReWfp5BAcoYnH7v8
1f24zry12eellVwnPN2CO42VegBzI5zt8IVPR1zpfOGixU5DxqoBId30moVkPGyi1NvP4gxeCOyL
j0j5O+KdAEtLkqqc6EH/c9dC0x0rl/8XvBjbcEaXUbUZlBd1UApy24xk67rYEoA5bI0c/rVM+7/x
DUcqNb0NKR1Z999UO7eYKulNdu11bCvp3pARTvpK9Wq7REFI/X5htDtQzuYKcFbydxT9GNk5CnBJ
8VnlMJzhV5pFEQZOp32bW9Ej7y4BarlGI2ZKZZ2MpLTffolAcPYd4s10cq5Tqj7YlgJIAFr5QjLS
qZWKf9314C44X+QsR0c9hzb+TXYVkgXEEqOFq2k7+6dol2HnIPJBbCborHxI4A5w9W3IvnfxSuuP
911ss43Mf/q1ZCxwGgBISLDTb94hEETpqI8jRWDgqDMvNZ1HcrbYt53DBdb0gMg8UgSF5rE5YRID
/1M53KRM536s3N/RBjpelwUTXWfHyFiabLniPjhgLNKy9JC1ajU/avR44CzLYM2DGdRhHLLYYmcx
I5+1XdZr/sPNu5VEd2i+zhVc8hoDwTFSmQeca/6aVnKvFZ6mTmrxBsRQmYw/0Slp54h0312P+Gde
UX80hgQ5gm/Jatx69mUL49GqJTCOqaZ2MurRFYvPCh1kZSdLoApaY9WRIzzAAsij9HsbmvYgT+Ps
NiH3av827saJ5/QX+SUIXvjjqFw5u1OBUOlbKM8Evo1YyTuNJOLEnNBL/aad8KT4Oi8/Xj591NBm
RyQuv04DDBxu1w4xumf8ETphAQ/pO8oD4oQEelEfRParhn5dD/CJ6B+0shtqbMcxM2/H7OmU5Vdi
/BdYFVq/ulITdoHhrW46EnpJJ00yfwrSROOjkUnbe883O4zC3Hxxqt+yZ1eDmaX0RM2X59VDh3oX
u9k42eo2M939IenKzasRjO5YX5PbT4Gy8z571z1PrB2n8hjZIL5g6AEg/MJUUAM0bRY7VBL/ZpQH
lvI5lPjM31dNwhyoc+Dy8JNGMiSX+jq2XGl5VmXTlDGreWfV+u2Mblj7IhHrrF2DE5cgaqxsqG0s
R1vkoEfg9tQ3H6DLgSMGdAr3wlvzHJzkqqcI/SkW9I5GZvlVoXL2QANojKiiVmKwOkwW3Ir0dBRj
ptS+OaSs0LiaE6al7HSMiRuDhhWojEGkJoNwe+BzpMgEXxcWDw/KojcuM+23okScvCHwPpFGNj/j
1GN1jVxPNy2LQf9hogjuUZaS6cRM5GHIdg6ComnYcnMTF3npC2Lcx928MjMMX2nGEIS7YtqjiWMl
oSgG5jOyO7Mv9GnDAoIcV8LuDNPfE0u0eQZ3Eg+W1O2DGuEnJby4mwNfCrN7eGOkgXo1lO6ufvI2
EcUj8Dta2tQwyIfkWb/uEGXrEZ7xnZ6VD1+eDB9ubbxgm2C7Trbn0Gdn90xC3OVqE+BMyzAKOLQj
HvorT5N8IUXMqeEgeWtsclGNAiR9WllG6z31Gdgtmtrpw8eikNuU2msxZodWA5Kts/dC675LWCbO
ux8eAiWwbihcpAnmmY4So6wYYu75vF4s+ThX/cR8+YNYymh9rYUDxA2GvDW6MzvENVby2kx8wg3x
G4TZq8VGg+5QFIujh6V0fEzJDEgDjkWLA6/OdkNfn+rXaOGRLfERVJNKEkZrcZJp6W1ordyTu6yz
xGIthyQn9uRwgu+B2kN0HvdxccMFmQJemjtuAMesI4oPGzzTs2JfbQP3z0QXDOiqFFj/w8E1thq4
K7XmtJm3xZXR+5LBvx/HER82P6VG3CNwMyyjjJXzE7gBYqGWsu5xitR8dluWN5Q+vkTk2QLWGgc2
5whHSV3kCxq2eKVdrdz4BB7o4V/b9sin52MBFSqqs4l5zZNV2qKCibzy0SqRR2tfI4aXWZS49UuY
cBGRdlYIA5dwWB681Z4sKHeyYLvSz33EvGzHKp6aySXJBRLEVqoeum8VBTxMGUmdAyw38jYWCJMm
qRIX2OUyRNszr5+oCRIOaVpxRhVBr8btqyQRJEfgnmupRskmc0ufI6tFPynAXrPsehub6N5devEx
r6wUy34YEa8lPdm/DXrBrcUzWgxZQGwuxNmENzNdUYl/kkRj30SeOdK7FGcjLwq3N/lVUcrW8xmT
3hsqfdLZIO0QrM7cHmIPWgJZHyOICx6exd1cik4jmacMHxfI83OItPjMZzSPVuNwzHwdf9IOJaAJ
m0eZPFF3Ug7GPjvh38IPeMhzfwwF/LsvkvsUMdBLyojYxiyD+XYiAGEQxqOq/u/Wx1yJ68uB24p1
bJ6HcUHcMv9orhXJko0n0+aq2+UGTUvJBcNr29ViauURi2nKxcK3BBkf4w2fwHoFhRmfKIQk/NAE
lFTMhi4gkpDrtOYiJJZZ4v2eEk7JhrPT+L4X/5EUsbUQ4Gj/e4NUm0FWHa/vEYbGlCu37hApEPSj
jTpSLC08qVbkjpTxvk22u/VKvqW0J+zuQOu9t2USrGx/p+veFkHdCiuJiXmqoFNethgoPFYVb2FU
dd0uiTP8oQ+HuSSrmoc8QW3BQwr0T9WVny9JPrTUuJaTdXLHimKhFG0Q9QzTDh5nEBsaAXOZNMcS
x0CwGFahiIjxjx/qpYwL/O7sAJKslKzCI4Nh67kauHPNQGYdrqWcN26isYDuBZT0tYI1lzWUaJ89
gS356kr679mLK6gJCHZSRYRj4Hb8Aa85NYwOSzAFO9WaGjcxCvKDfuduOXCAPevYYF8EHe8xyfEl
wsNCR0IvGPLYjVA0k7CC1+5Cdk8bIPh4odd81VG0SpVxJsQ7BAY5DmwFAe3MIhQ2BIE44bef8F2E
+grhXydTBV0KbIyUjrA7MTsHOaiUDAdVkhk5cAujRze/IEgVJWRfzxEP8l0+gNjLbAAC3LqpkFns
GM08YvCF8adbBeU8dRZbxYn6uQ7dcIWygxrNeks/BX6EGXOf8pKr6LLaien1+XV3zTXMqGanb27v
kyBa3TZJbZTiDeaL73igBLgJF78NauTkMZQJx3nU0hRU6cv9bCRFsIAd8cfglFshGTBM7MV/Qzhn
Uw1yFdYTuGFa6nWtZOzkXh+5JJ6Nwn1HyTbh42KtZMi8sV3ErQYCB5+v0sxl8UNJ4PpjwSchy5JA
7UkGZugY484e4mPeLEUJYvsXotv/SuR9nDmyQeSLaAxZGKmGFOyWx4HLmTcuui08byPNptoQSlQB
vUrE/iA/AWttyUUZFzbOfHQ44OKi48JskhiQhmDZlkt954adHkvc55BuZxk6LIbwu0M2AEYkkft7
MaiO0OX+xmuy5hPKlGM2NeXaQNyhhaOt9R3UVg2yqx63ik8FdWBAt1t3NjrLCwOrsB12RkT5a7cT
i8N+jJ5JVwURkm2Ncfcn2G1z4cIxU5N0nSOLk/I3MZsWfVDMFfgB/q84riO0zB5w98AoorKLivkc
K/JVMDA4AGH7K04bGd1Qo8IjRcTyhscVcLQHkdOxPD7hcsxXpA3Uhufnx72ldExjwwrEHQb515qh
VuKf6ZgGuZjQ0r2S7G6BVDT8zfNnUAiCGmT5nVwyt+DJAb/fDrJzrTQrAij3YlPSg69rLloCu5A7
h6sYfeWAkA/GOIo6CNc9xYvgmemaUQnhwRcnWSJ6lMMH+uF/t6RIJnyASLeqwmQzRSZ4sWgdIsb/
8sLDXa8rACTD06CTP62cHppDEEQdd95oYuK/0QqYQ8XcDUHxSf+EDPyaIppS1ziPBD5e6oUqseKT
MLTUPoDadCU144cbx5qiR/W74WW7HERtYg9MCiiazhpVokzaNzrx7yHC6ARPBodfgnZq3K6EI1E0
gqTXsZvZ+KGV7LG1E0khff0flR3Y9b4JtgGg8YsPHfscploEw1G2809QKPVaMEJS24e1zJrPBawi
oijoeo0eyZKQz1FUj79HEdc0Vp8VLMSwzDyCwfUzCTTEx6kRZtqiuQcbKzDWsh0uHF7TWKAzPciU
5ShPhkWG7z9310xNNpxBc5kcQj5ieQJsY4u/XKAV+jTL3AD3w1lfm2lBBCC40Yh9/31ZUGP77rju
nKdRAgXbamEn+2+ME60dId6S/IEW9/qLTR+w0m+wo3aegNPkJOMY5ByoWmBzxZ3xmYuunNpQnzz4
1WfKbTNk3kzkw385nNJjolcnbMj6RugWEquyzlzObYXdrmttW++riSdNvvvVEVRGWpakfu91FO8p
t8Tfdw//Qq2t04MZkoGDH9tdYEdlFOLtXg2EuN4RfShHQ7Y8pxwia7CmfS6envGfA1Jv8I8MpXQX
LfNOqPiyN3h1Ty6nFacN6IBf11p6w1geUb7suAz7zYlTs6ZW9WEBrg5bq8NXgIGQ8hpBQtFdCT81
HBMAzQn596hz1uocO4JNu9V1rNmqStFxNVDcwMPsaTtMjyp1klnwK+Glm2KlYIfYbhHObrXjr0TY
zMXT7mF7gIzRYzbTidMGLFL03pxNtqXjlXHm0YYO92duEhJhZ/g8DH96ipvVy+JPXhqZU3Dwvz1u
cpESE1mF0Ek6qrrNiCJrTm60wUeR7a+5s+rpMJWswL5HhdOaiy01Dc0muY6nwUT6VQRF4nVk8fY1
eVSULe9W0XgLBNkWe1DDCX4bTWluXTv1ZCTb4e7v7kKzYuOI6gx2L2IZp8xv5n37N+ZJ4pIUFLWD
IAaUu/SHqiWmoQiakznSQj1lc3eF3kK6tC7FqlmV9nLs6ISX96HjQpE3mF/b+tCAg9YRfROvh2zO
YIRsqLHDv2gsznSQXFvQft8mH8RENkX4mcFuj2str1YZW2odKz6931NFh86YHAwLvI77+RBhjpmq
OEO5RtXfxcwsbqrudkYeCSkSGHx+NUKLd3sCqA9Xu9+XELV3LHs+fn/uvDMrCZOtv2jGlkeqzEhp
yKE1HucDjI0jxPTxfBIFbatbjiaepVPdoQNdS8cExPjyP74bfnGelM5/4bHzlXBA6PmafnFwmy6s
3JRP5OGkLEgfpBrh/shsqFZ2AFrwXpzSfJROwGSGDxK5/Y1Oov2oiUNatI7Rz1Q7GfuWLbOOSJKl
As5Qz20b1P4vdYml4819s6xiYPngiIfBFucQH3teYn6tQx0wmHZg9D+ypMbALwTt/8SitTTdm34a
oXXjZjFrlPeJh8lzfO0HyHRQnZhnPQJa2EsCAYDBySpV4/XewqhefqIV5oCSn164KTXmSJmrXeWP
ApMg756ovwEO2+jJAHm+UmTHWKqZyPr1lDrbPGXuAMN2G/Hbzf+u9aa3QRZ89xHMWsUE5p+DKmGN
ctGRQvp1zKeLRwAONKYWa9u1aQIlRMqZPLQbWTa3tw/DALybfbDV6BNgRQKJNAKz7LrvxIraw5Kq
uT4VMJ1CbfgC1ssPi24kPaeuRAS5ITd51jSRNQAAB+yM1CT7JLWnx31O7PrSn9spd6LG0yTtm81K
Wtk/N6LcKUGF/P3H/SJCOt3wPybzVwjhixoD+5zEp30n6exyyrGaquAOCHsh3hGjvnTODKKAQ8JT
O1R1PxiHtZ55t+O13S/NLh/uG+HkZrB2rpovul4O0YkF2mBo92RAP8vNyuAHOKfLTVBHRrFMrWY5
koNZvJ1csH5Jsu2+CsGuUDwi6bUy0vwyB0S5sQSUk7/af0SflHDsNcpKef/i+X1ap6KlYd6LKQO2
BI1uFrRizWlSasd9GgdGhE5mc47Dy8WUWB6nvVHVGcDQDZuq+0sglnFXzfITJ9WfgbORdRwGgtCr
8z6ryjdBouAKpatFYnwLhBcCuKOLMwsKPpjfaafNo0Up04VeE+6aizietn9O96D0z7ng6fhBG2Al
Yfjs/5jScfTDquXzunCRA0zTnOL4wZahpZ19zU1kjlTBNjjmQsU59vX3xQIMPCF7P0PNYxeSDt67
W/81o1PPFGALWATkwhvp/F4OuyUX+lSTTQ+U+25aLvS7LhO/JMb4lezlXjKs1kkNncrGV3huLoFU
DtrRIb9r3g70W99sYtWfb8ugtPbUipI3Q8DjmDnYuVORy3fnzwWqcZavTPW0Cj4QmX4aymmUNokR
6sKpYKfV7HUSyTU0O4V0Yy7y9DjRxqcUuhl/DAWi6OtQoKiUzUcchMytf0aXWlHPxd44JL+zAiUe
XbMSFnP8XJ4ZUiSJBN8m2yLmdNoJbAtCqDmkl9RBTCaO9z7wzHfF2j56lvkFyfekK4IXeL1DNisq
nzGKfb7J+lmj88mjZT2XLyLf0xPPjtGAzyEHsGHsteQihB9N10RSImJQeK3qdW1XH85Q3OtbSUuD
lfuE25L/zEKD+yEUINBR91acjKD5wUdUTW5etcaZ4h8E7TaoBu7sXMd82oHUrBMeE5Q/qFs57zPz
wqujWBCu5FJQBC0pYV0CeJ4SuW3P4RS2w50p2imkdNK1tg+syfj4x1zYdGXCLlajessCrjWqz0qZ
lvB458Y4RD/a2nNBpnoapsyGc3qCbffYSdw0QzQm+hmtrdX24RjfCQB9sR1fQFCSHoKcHWdlgxmc
TQlFwQ3MYRYF64w0FvrWHDGwhiJzpt8nvC6V1DeHezLmchl8embs9NSt9S1w0Dlj+j+KOqAxS4SD
MDS+cL85K2anmuqncHi0+DOUP0v0+o841JNMFyBU1xMd3MvCzFhxYcz0qQ605/IetqI56ClJscXI
NCy5DsCNNbTf9GQwHHLTcPBhqsLzSbqI7OlBQlfRKM7V0Cujhy3eiuPEIAWnjjZRoMORCNd4cC0u
4i6ldRmNa7wjAIs6g7va7GijDVsZfpzB1jqwmPclVLAIoAOIrHpICUntcbl0BOhrfo2cmI+tgpLr
nu2z1HPRwbG3RHdi8Oi/IMH6Ad2HzIGBxU8jJJPIWnntXeUehlL8OK33wkuQUWfr0FyDjtQHv6Is
1Au4xvzW21aQN3x61KkYvBtHoUzbpX7W0fY3qIavBLCKdHOM/zU2Z/jPWygNcuaojeA7s93lDvc3
51dShMeBAmewqJcaLS9E3zFCm1iNL0CfcapLt+/WnGCsklntW2XIKGrxfX6UEGt40kJmh2VK+nOH
oiUKsiTV9UE8R8wBq1K+Ju3SwJGAKq0ZvXTFueSu1qOMxpujmtR85VEaE+A6aGqZ1T7JbUoP+bl6
0q6N8bGxGVxz2a8x4CXDs617U8QPPI3wV2HK0pJ0bAFRDHvbS9ceK2fqoe5c67Y+dP7wU1jbZhr2
cXShVsA2tEHhIJs955tEPRZvYH9ws5bgiLUJo03TjVYxX9CiosYsAYgY6dZPizFxW7qg0CI0LteE
16t0Xr65oKKRUrrLDoDdYy0Q6lHovhgGL1kjE9kTIZzwPbrUo5/VN3lJrjisixsEuXbTUHsiTL87
1PHJ25N0SldMNVhxk8j5MIJS8Wt/cWM6hQNipXPwBvd5P+n6ng0FFxbjCgly4romORhBjNAyaGVx
92iK+yWBLxJEKscuKZu7Yf+z8TqwQpGj+mi84ZIPqUBf0nYfZdGvyRB8tru8lg4Uiltx+Mo9Teo1
E+nF2A8pLkjY32LnTgGR6kD5JliEt5oOjpgNb8vEPVAORB9gcSrEROwQT+bKGATA0N80pVkR0PS9
jMOBUzJsFjLIGFAIn+1sNwu6v/dLHjAG/XVm9MpAWQI8CJ3Yq7vC+CGUEiVmx9sXeQYQQOpYfZiC
XaZcgIDZvXTeVjurYCiZsJuY3YvxM0l9ikZI8Vv7SwANtYxGbfZSQYYp9tHeIs53sg/GVdDdl/3R
gGAQ8gcvtH7gJ+KoZpz1tCt37fiDgU7wrbUigvmq2K/JzZESHctK8eh78Yf6sZZj8JZXCBSvpe+j
V4oSsKZh+F4tUh5E2/+JfybGipasDQu5li16VibdfxgW34WkMOArKM4hKSIa08oS4fPCJThCBm5w
4cUZftQ1Z8x9SD96TD/1EKfIDgk6O8VRcmKxh6DKy0ykm+T2rjeU46uM5DYxndkuP3oSQP/G5QJ8
AvMQ31C12E57IEH3J2GwzMN7psrPPIlol0F9PFuvgyVHg5PjMb1BYkiMaYmvpDFV/fpvrdXwuXot
VUWOzylVE4vsICAZ2KKYSFqf2emJxKL6RhA9x57tG3qG/LTPBh3SESSVKCsVLnP3MeRFsnzLHa3V
dJgjcLsrYeC1gWL5cSrsXGnPvtlKMVU4svOgYiOGmgQ+2MCaImTqyCbCh5NGZYt5RPKDVeJIZX0t
+dsPWtX601Pb5eU87JANzLK0RRfcWt0IKPEhbD+I8tMV1HjDBmAt8sZ3zMJQJVixz1a4Gm7lOO+Y
KlIkMF5K5O0+SEEirkUdVCBw0119laMiAndEPeMGtPGBgFjGr7fGuFr7HNQtCC9pns2UZST7Gtlv
3W63+Qox1WbQ1ztaL5uHv20OxR32OL4EgqT4YgGrK93ti2QCegYt+7P9WgsAHoGScV3TtsKEpTgm
NY1a6FddGMIeTsoQaiLLaxiGONU3s+dsF88iRBVBmgZfNVilRKwdRayIcIH/OYPxRO1i72s4E/dJ
0nRZQZmUw8/Q45SYzGCMcnw3xqMUWI61hzLogq4wU6i+D9cXOzev1Dun2eyaBcZII5epp1+JKCHO
ifQzVX5JpuznxobOnwI6NnLYOaNglOWHTDFcykkAE+V7fei0+z9vZlALQjKEzxA67d7k4ZLN1T11
HyGLmMtuLUs1CVa864b/4u74jeRh1v+k04rO3p0oFFVKee1RjwE+6slWr6W+4BuBaedwCTy+i+Mw
Lr7K4+H8/RKgPdrqX1CB447Oy1iv5DN94xqPq2SPVqV600aH3pphbfOYsKq4IygPzhKX7Bqg91A0
vtfp7z2t2qI+u6rY1nFKjznLlYW/2slwTqE2gjDdTe66pgcmtiBjpGsUKznsp44tUq36JJRmsthQ
N0NWZOsaPc8O2RVmrzU3taH+3aB5mGG/rQjhcZOm3Z8ofAZA58omfhyXoaaf3OHJI3Yxljtvr3Pa
T4XMe2jcHqP4gWcak2riuqVejsQjUexEpO9u+QafcUKIuUZPQeBOjpbwberhGdvud5XU9BFmI8dE
Dyjsk1xjmyONMq2jCko1lz7bJwWENzZs056NPlbvdPTiIBQ6ltF1cnk63aP8gaVD+FhLa1aNSP2G
fFmbdbZisQV9//xC9OOA+fIw2dIPnlbMrtoMsGmZ5XDJwzi5Ncx9ivKM0WV8skFOsAeOXUkQf07P
YWrEj91Y/rEalfjQvgrCkWgYWyy+1L2vo//y3ZoHdD2i2niljwjWAp07000U9XkxfKCWBcuPLUMN
rZ/jLtmhsJA/pUyF1E1eyi46ip5zP4DL5UzBf6w38Z6TT2dDwjEz6SaUjw34LY+khs/pgBwcUnzm
NnuhrkkOLSFd6j7B8kI3IWRJgewoC49zUKG/mUpQk5Jm7fdDjWoRmfxrQUmp47XTX8bdIGDOOVz2
Zx6H2yeqWafv0X8Df5N1EIl25Ab9M/OCYBBSc8nsZFp2Cvu25u//kwVJ2ZIKYRjT0nc2D45ljVVE
aJvbCB2/cg/jEGRu0Vc51eHddTnhFczv6ZS+t0KmMVeZ2zYxZUAcsFXx4I1ZrtAXnOrRw9Ftvq+g
E2S6ncjNAxEK94FSXSXXXeUyjG1HTobgMxEfUJBoq6wRV2OnHu+qpyqHhJmARZSRWJ2PxWI1xFKw
R9I3SNVFf5Q4MsqQMOgGHKxLGugST2e99xGXqro1k2UI0/ZbSomGq8Ta4K1sC4LAlPJWSmFAjqdA
VH7VTy6Va2FG0DSrMaTV7CZPCjaAt0RAZRF/pL6n2Gmywqdpmmx9Po/baMacNGBQaBYwpnpsoH5L
WaIPRpE3sk3pOL/Yiu3ZEbTTW6q3Q3lbPlsL8PKuqqY7Pu+qvsaS4v1Vx/hzhSskjWOi4jP7YfCe
jZWfzNv6O5yqGhGE5LWmMjrXv3k2H9G9SHVCyu8dHc+Pb4VflBwz5wRMmOR3wE7j59+Lp/qf9shR
CkXvRecnHsqN5UF0VGabLHjIqg7U3opOyNptKeui6D8LZQya0osBqqg4B+xcsm7N0JiGjw24Tsg0
cfnm9k+rahF7SpuLTq4gUupqdU60SJkVGSbwN4UaAgpHIHPgsOStm7U/a0AQ8CN3e+CVUwwcXC5h
spkfZpWW+jaHkYFXpd6PJQBEyq3wDx7dnF1mNIYtqAH4c6meBfgacR6MzpIv0vhcFGQdh39ZsZIi
7Kfn6uIWQ9z/A1duAHoJOQ3hVXObWo9wDx6gRAfDh/QoQOVFdOukytvj0IAVccLuc0jYKu3FsgR1
BvjJWVupPJ7tXd053KKXdjmxrEUZSddKYkJiyJFevxvTtu5X/V4xEfTndUqCqN/87zPc+yjgC13t
ptGTa8kpVk9Sgpu0tOdPC0qhPnceP0MJZeNkmOV/TvqTbN/dPh6X9AZHNQPDeYL3OBdLRB8y8tw3
jYDFQ4EoMhXpjmQucNo+kbUKAa6J0GuVxwcf0I+/Vy9OCsCQtBMZCOmTS9WpDEBFTBfszbAa7pmg
Soubzxhezws80V8zJ+XbhqxXG5VSk/fDJ1V4x8rpr3Da557GgP6g+LGUkogY+il456GLDy/ds3Uv
+EeZDpnyxMzgBMWKhiTYp3T9TKSNSKLUT/SMVGHOYUgkqSUp8XFQy9sVSr3gQV3ZRACAqpH7fJR0
1nmL3esU1S6Gkw7HBfipaEnV2ExzUE53W58MYB9y/q6eRjei9mt4W9IaeT2MuaK6PQfIWzmBvJlg
vbz7Tt7AONpkPzUl8omg9tuFlfeh/u3Ohjk6BjWX/YC89wnXjRhYZ2VE5GwvgiP+2tHx9u1ZBn7v
GaRWacNoWraGDZFseNR0nl2AYwgUh/J7ciTnCbmNymqRd9Lzz0dCaovMHhcJS/HfzUbo3WCuY4kz
0ZRmocnm5SzznGPBdU384xEiVNRqY0prLOtnU49TAByUNa9AH+pZL8c9a6TDcaVmkrV1otJoYMSn
svhaQgknZHcIRlpaYwpFiTcjklG2T+R8eEUGVxMHgC2pikDIJ3ulCDRONRg6AxtD/uCtkm83t9uY
eIliSfs3jWqYCMHYLc0jQQhTwDys7YMeWRvp/QDVijEzW05R0mkJhgA5vXGyQg8K+vvLmSrLiw+6
jS8tpc3UM/aKL/SEaE9hDyo+bC5/fzGzEWpEYQ8wMwdeVjWGErvwLJ9JjD8my0qv2/u/RdY0LWFV
zTvDEVK6imFuigjd31xrbJTQ8wl1VCOXHyo4kSQhfhTfAmr+IFqE5oCiHB0F/5yuCZBJU7+RMmTP
r3L0hJAMOedIZaSonbKgteFlDVi2l7i2FR/w3p0mg5BVFLTq0ZH8Hk0DFpFjr0C95KY8MgBDV0jz
OUDwNcCWXJ8J3svrBvOOIuRQPYg1qMyniL/oAE7mftHyA69jxDHsm1tvn9188RZt55fg9KCrhLCj
AYx440nkd50OPtZNWCSgjh3TQkBZsYcUFL+xlpQIa8Qm5FBs1GlRm0HTO5VOowG7TtfLVXINydbb
KphRQeVtM4FWXj1CSLgQ61PKaJtDbaMiVkna9eWk3BblnB7LwbwPugYEqcpR8Y1b1U3qWcPjolwj
SDTcEjnGcYo+vqfWhbCjRrrebZlPrF6y0dOoqGr7/PhXMf8eb2B/xIcxJozdQmFkBC06IF0VjnQe
uEk1JIBGZw1GDjvhaOd44TcH+bxhsWKwmqlcQJ/I/yu51R+q8eJ5k3aZKgRf46ub/X50I0BSWx9M
qhh1EQxt6EZiHN0Uv/S3YYywp8amqDNu51DH3kPKt/IFwQNm+N2mWmP4EUALQnQvctpR0uc7/IYl
ZaJDHRrJwNsDMQQe22wlxgFBJudqhQEemYOa2xeErb9yWYde3obApnQcpwwyRi0Sh0l68rE8OtcQ
nfJLclv53YHjb22327D6YTNguTuDBINNnlZgp4dp+DeSMd1ZwYR0nHDAW+GoziqlQvEN5hzKXkhd
qNYZmuvEwGycOjna9nPqaVoAHqMNlB26codkCKs5ZvC19L0d1mQq27TEGrTCB/2FLRpY06iIou5i
Nii4qHUtlWywKhHYGfqFYVqdKmU4xsTwbGCq00wouut4MIUC+VlPZ7ytxcF3VJpIJENYuarbesQK
WVL2qsXUu3WqAd2SAjo9Bybp/21+fiSm/lXotar8RdrNVGg0xmTFhtuSrrXJ09ppQfc6pAV0eyP3
3MNTOfJyOLm+PSYqLd9mu0mRTx/DPSed+ZQARYTT/WaBgpcIFDxEeSxgyq7NWAR/zoEMznUGbgQx
zgqlUNlRu4pbXeC5djR4ZhU9AIsMJzj6eNhpFGAzjTHvESu4OtZ+JYnOEm81b96rL3u4m1modaIF
rs8Rmki0iUfK2iunZOXr6G6qAB4W4yh36NisBgLQIXSGF4kNFTf+F8kFHaysA0/h4HesgCArN2bf
8QQP4zbxaprYVd0NYqPDIWh1+Ny/VkSGTqVPTkRcSnAz7WYngZ/SvsPxewVR9/rT1TYGvu69rT2J
JucztZodRfyV/BCWzQ9an1XBGiR00ZicZdwXLMHELPnFhMIBIBjSuRBI8SAMdUC96014M09agr7t
fAP/+ixkz8EvlUBhv5s3QcLRD71CunXpaZmTkpEXTDSzY8i5kcIimUraVPQ/kXxGOJFr91scwxzg
8xDio8mreVeR5TR60rhOObJjC4qaupZjIJVOtl9YKQXoTy7byDVdzbItSfX1ietGaU2Z6YFi9iO4
1dVe6XQsQzDqbJqnjqKTHKQ1o/RnzLIdVySZLWv+bG9FCffAARHrYYCO/CQSSOkkn/cFRSOKt2w0
t94HuKS/orBi8HnOpkfLS+7ptwT5lFmAgtHZq8jqYlWeccUgUbb4gm7hCoa//3+5XwHaI8oepm3f
A7kt6DA1R16A3Q8RZuk5WxJvboFqLWv+t0CxuC46qBmGAZYGye6BwWi9mG5Ug0gL8MrI8hbzdD3m
MJ6u9vxAIKDqLSHSrV4jOgUeYtQRlc/U7sGNC50hN3z/Ja4zOCJHCfZ03WK7yYgHdUnqyPuWm4Wc
K1slnYIxaZna78Y5w1srH2wa0Q/Fy3m0hHrKmkn0b0gtYP4T6YQhw50x+9mBjIv0vagNHNaD+nBr
AnisbEKbjnG90vl74VsKm+EvZ8vosVTZDA/mhY1/Cpe/LnGfl4dFrc3iu5+tcle+cM+az4c/0PG2
3UQumwTRKdLam0ivPCLHsLJhGQSAFGDT2J6LnUk+oBETSMPWb+HyO9EbIdPHUgwu6rR+EBMdUSd/
nxiRRI24pYBkC5c1kcWYPV2bPSmcQpDQxEzh34SmeH5K2n1Jsnqhc2ZzGcDNG60dBaEIsjNiIRKA
5EaAHUoObRNKHXU79Xtu1lsr7WhOIrtSCTNiS4PJNvD1mqHdfv33cMsVKAAU3u1lzKx5sDeM9cpA
TOcZO/8nn2ek4SYxj9IbNi6wZqVZpP9iVLO0ZTFt7kCBGTQW1Bjeg1x+GY3c540x27mWgwojAFnq
qVB0dpop2V5GYJ4fYq86HK/JRa+qkLUVk/LcUoL1BBrw79TGvAvNf4NKPKufs1Pfph27UggDQZb0
jMzutZxcUPDPye1BYgXOycmFqJCTZvpMN1U2dtf/pAc6DrTd7396pheT7El+RJ76ItIeNq/3k+QA
JG0eYsNeCkGj+TA4SJVEGuWFL9HEGVjlfFPrX9lTwugcBL1tYOAK9Ct/8kZ5CaJwPcaWUl//Uftd
whLcjCQauogySH6T7yJKZv2ety2rs+4GX49dj1iXYUYsWW1RlVlnqD3DKmH7AhmtDmifQzFNw1TJ
WkDiFQf3EME+ebmqbeXFKoZ/n4kXQ98EYv6X5PEMPXxgQmG7CCNa4JcNc2dh05mU5teoyYFyV3UW
rrtvmLOKaX73cICSihZTf5oSR7XxHcOSseHJtc3tDbcC9k70UNxiU1DgYrzMlUsM9dp8jl9MwoAu
IAzdG1GgWK7YT/2i8svRnQAtzIZgflvVOv7UsusIQhBHNc8eqL9BUwbn5a+Yy+3RHTgOBxxq56Dk
30UUDPd5y3nlWc4zuXnZ1+0mU0VitLWAnLc77yPYz8zPZODVWfSkK9Mmfh/sE6O5zzCTr45BdMC7
3nn75vTBi31ISyIKaSwijPwZgEnV1aCxlx6pKQvFf55zdyAjgaou3nagzdUNI8+Ss3l26Veiqhm3
Idcpy6uWjgNdD8ZXk5LN04bj7+64nbjj4LDXs1lN/tL0tXxHC0FniT6bhZBq5bo001uSL8O5c7je
ec2NBBIzp5yc2Blak1qzPKF4sZhGe0Li8xkvz4Og9Ic0bz4GjEwt8QycCmJ5d1q4zQ2v5dWZgTiU
l8HTHcu9D7trtja6+fQcbQkI+3tUp6y0Fr7f97SGbxt/4LU2IujjSjVC28JzaqB75P5mEj684lOG
vPPZFMTQdQG7GpCoPQ+jkgldAKUeQfd/NIElXrZw2q3EZ1Y6ebSdSiQ41yq6C75m7NBkSFzUmk5P
I4OYR0zH1HQKYbgFIVGShPwk/OX9L41wkCjqLZZ84gauoncOxozhFjJwPIq5m5A9KC2p4oeRO7hy
cSeF5LEJmgp2kuz+lK7mxGFdqi9bIVBKT79+Y4+s19f8hw/hpSMEcYf3+WDKp6ZjBAG7fz0WU1il
HDqt10fSr+rlncWv9k3s8CN17fEMuR4L7MJ57cv8XrkmGpAhNHnoBl/Fix8pHCnH7B2ETqJjYo8x
GQcjIxfOJ9Lr2EBLJINqBhAHCXDnhA0mqkfDNY787zISxoIbAMEizJqTPjDkOWT8/AMtLY0mn/xI
s7Sdkmmq99Osq10AzSrtnPaqNNWLEugFF3HcQ2I2eEiHuBbpv6y3dc+00/Z3aPivqkDzOeIIUXwi
7LUpc0hlXb2MtWC8hQaKRIuOqIxVCPjuivO1saruPWMqqFnpbWIAHJphPXPiU68O7gM0YQjJALe/
KUFi07Ea9Gi6jruagI3yCBMFsaZa7PIlMO3KykantiRzGiEOKoCqbfBCOQ47KZlgn6n4KZxjTTiR
d+F8xAiZGYjE3iT21frwztUE7w8ecWnFek5PuQPKNEn1qzlDzcr0Pq8S+2XefkhHcEHHhsXUR0dF
+SljrQdrLes+mofT6cvtH6D1GFiHHsYwwSc6r0xQYBJXUFnsZ43e08HYVuJ9E2K0e3Pxa97MSysi
2Slg7dhAB1UOF2e/asPk90M5T8wM1CMg75FKaUWinsz6G68Wn1pnJBRRgja5519Ue5TwuNNgBtLv
NA2yHiUshUuuF8ooM/AsYRVIMbwJAaJag/7NpwAPadieoBCqQ7KZSQ+goR64i8EddT82QMQl58Aq
qeNBBUjSgo3ZxtbOrFODTV6EyvUpzBRERgkExVQTsAczysUn/sKksxxAOviZxFI4ywlkAUmXM+EK
2WQi8aO5AsKf2yVpzYtZnHHLVRxRUq+041ve7x9vXpYYfee/Wfw3aAC+M+KyT2Esj7p1DVzFkLPR
YyAevwXP+oWBgYlJVvdD5eF9BpRDHqYGiy50fsh/xhbdzpf2UA1MCoPKVJTB8wISUqIq8In5w00K
r2lakCyPSTo27FCbQqkpyH6zrG0I6+o0AlI/SD+AhzIuNeocnIlp0CtVU+Qr+TdbYimP/w4trW+w
gdbIVTFpHr/Ax1JLHerOLumZOmthBUBQXc5Miaub15OSGrDex30zulgaj9c+a7HPDWttpuliG2UO
dpIHtWyOdqhETigS4yZh5+bk/A7LGZQ0XrAVu2feqsTVEs1pi1RAnP8e/ez77sSRsauzHtSIw3WI
NNKf//Li2YZ3I/AtWfz6Hhq/LiqHDfkmN5QXYRY+BlTVE9qaHmymkF6j5JoCkyMJaIwc8vpZptlt
EUKKRpDNWj4Jb1xHcr6oslpu0TEE/UFgfzrwsUON7tJhYhe1aVtLqzzYhE+oWIOM3oxiBjU6VRO6
vrxDpQnqbFtxWXLDQ8rLvMB8FCg3+3gwX8BfNC8uwt8QIzDUOAXWaEX9tI4GYDVBt+88rX0BTGgS
1ZpmxHjO9Qsz7qTEeeHbWmVxEvjcPvxwb/D/cwvbZ3l4otDtN8pRPJg9DCTizRpruAQXbWG8Nrv8
6eKjLGKGEmeyfr66H994eTsy31Q6QYlzSBzLr81WtceJopIwUXw1ZLGE0/x00o7RvKNP3U1q5Y/n
b3noPlnTkoxMJdWm6y7R3dEhBJt8fYAN5+Jyn+B64v1PcsXG8FVwV/18509kk0Fmto1h72CN5Yje
Re6qRZNBVIy0Q6tbi6EFJZuCD81x4ZKVO5Vlo1JhLhVXxqEzqRvbqDUW83nsqvMBD8cQck8uEE7B
W3a+msd4JmR8gvUZACvo2O2BRj8Ny8NNZuPPI7ZWenkoj3UxoHWHO2DbHE1DjyBxTTSTI7k/a2C3
bPWFLUJoFlKetp+89jFhWQnv9orN+PKN1C5Oj1lydx7rt4fRn+EB3H/R7Cc5InoBetGjGLQY+f7Y
XApGzTU5FqswttoCgUKN3VU7rK21a1pT3VMabqsKjFsT90S0Ot1fkpifI19OpRiQCRTXxR0CXUbL
r0Yn2d0Pt+z3xOTc4BxR/29ELEMg1i1Hyp6mDlt7LyFoA8kxlZryTq5YGZa7ojp51OfCfzgPrPgV
Aa7LB3kNry4p1lw+uR1kZ40PJRyFZmD7pxLOqu8msOlNPl3wJqdtLGcEHe2+ljcNDXYR69FUvDhU
h6yas/K5L9DsNpYD01tQYx4Za5bz2sDR21GEtb3FeKqaPD+TkgPU+IKP1Zynk5Orzsmdwp6gLf5/
veschO2JEScuEEnl9C9qQEzG6vwIUTOzasETYzJHZl1aASzGGodPzd96UOL7JAxmOnlrcL/MRxHe
3KTTY9T9xtTrYdYHfbOppqhDmgqIZQ/B3Q5Sok2GgC4mZVV4e4WIz6Q/zETFNbwOJVm8SmqLWxop
1VXf+Bdh5vYQ9TvR1hu+F6nGuddr2qxISbJpoi61p5VQfmu+IbCU3y8XxXKPjRfPgANNXpv46PLS
n0ohQdNQ+P4rkiUPsQ5A3LtawFTb8wmV4RxCuumqKm9XDo5yEVrEoYYD2+Cx+j2ab25bMQCc9/eS
BaeUwlLh1xEE5cgu6NFH0NSSTBHJzSYAT1/SrebSho/B7a8Vv7hlN33QcjH7VBcI54xcY330LcUV
HjxaFFMWH4+Cg9jhy0QaQWpnnuzmWxd+kpy8gnx0WvAimhD1SKrxbSkO0nnq/aUbU2YUnz6e/s4J
vqsbKZzNL3QHkIWj1IV9RwCK+QRcF4uzjZJ2biqFBIKGVykYYUsnPp25c4/vQRtgT2B2SDCJUsJo
sDWcFEPuCEI2reGwznTTPmD0FGgTj2+JkQmdcyxri29nQOz2Je2L6D83MjWDQS9uxYDR280qPyO8
bVBq1JAQef0QzSmpEo9JqsDueIkcTTRgk9aTVb6iMYH3SkA7UZ8kO4F+12kUaV49egLBHzL9oxDo
5v5cqf7vDw6MR0IF520oB46VIu2Z6PzNnD04GH5lcgmBte0FA55fgWcfTYSuy/zklBJ0N7pjJMfb
uXjQXXmT3/necarSxyT4mkG+G9JO5Q8yvyQs+bv2fIdrHgspYXVOHLOGEScApbPud3fW3b8Z1btc
mveTVr+bRvKRNT4pJZ+ebwbcOv7QlgycW8T2Fw1bAjhlglzFw2T0nroamr50Dbb6FDMbZRTINU3K
oUDq4MYjBLhOgATDMsiymr1dj8+dn955pAklPi6xnsCyxuHVBqRlSy5l+gA3VPpZMGMTy4EqjEiu
L6kSAILYH6z0QHblx9LA8cA4o9iih9KufdoI2xpIaVbGskDkFFTMczZVpL6NhPKnAfNx6GH+9s0K
lGg749ogL/Tk/u7GY30OaSTkK8Ml9aepYqQNeZHcRqycqpVp9wd7WfwfUXMoKyoXQc+/+IffWWAm
TSBLhbEQycLImSMgARJdvczBlxyKgm+zuHmgCEcW88mtwKlr0GwK4GMUOhnHcTbtfyPEL+jg3qU/
D8Em8sK1dU6ecT8+EmfOHB812WE3uFeuIpro5MUIoyedHyY6i4AH7DafnowF5tZ2JaRvX1yLqCCb
h0lpT4sZV1vOjM9cMf9InQ8lfAq5qc5j8dAxYoqlHYqVAo9r9rVdNnHkTIce3DTO2GcEFXyLoR49
gF0fM5bspgLQ3wmnmwPnwRSDEFkk+BZIawUXBQTTI9t6gdh5mAmIix0HtfuPpK1JWLIn79bNbku1
rX1nPa8FR/GnNcyYWGxaOysbtnh3Ff1OEZW0dST3aZMg5wW0L8hLkc36PxFhPRin10O2btXpnliF
hsk/Jz4Ud45QFfUTohAViSVuIih00GKxtCxyUa4aZATDYUHSdTcV5pLccN4Y0v5FKZaiN7xMzpOZ
m04xcNFyrjkqoJoe3wHSD5BLRGODsQw4pPJDe2KyhJ2SQiEmsJfaL90lp6a5Id2rJusNfrqSwdXi
tSGgO4wt1zYhI5hNXctsVr0IVmkFxYuCt0WCNG8+ndLZNLpqetm7WGP+x3YXHAXyivpyItONlWSj
5bTxVLdePmEyFusC7dt60ZMw9OzSu3mzP0BT03gCDTGqmZd181jGT8NKv+PFFsy9BEb1Fce9nFgJ
PJSqAbcyBfGyJTdS8PSHng6W70JL3YYRyRFCcFeTuVIdSVwqYxMSfPOfrUQ6B6H2aL7hsw7GR48k
hPaJ8g8jPgGXPjI0tFR01d1bZnthP+bJnkrE0b+Sfj7kUpJxn7+gox+B9WSIOa0Uqkjetvb+neMt
e8e0GOUJ1uKK/MArFI8nxJC5y16CWMcGngyDYpzttBiRn7GSHJGu9suvJmol04qhAEWsFsDMacZ7
MIVo77EoLcjOl2KPLVgZBsB6rdjmWiNhvdL+2+c4ZmaKGEsP76S7Qibenj/Zo1P3hUSCWaDB0b7h
V+5etcTFRWAooZZvZGcvo9iVuKiPBxS6YVDOiUN1GALXqC4Yo5tTe601kASPA7aM5j0BigUtdPzy
BO+9IPCUVuy/GQbCzf4ydfiBpvcg501lL1lh31IJO1TaFVsNe/gz/361C3480K5STO2aHdg4a5hg
kXmSk0kPn4RyyUIKbDdIayX6OHYmHU+SXv2x27+VNhQNdpIPfl1OhhqPkIR7QRmnw/sbMn3Rce3j
wDV5Ny4mXs0bgKyClsYID1wKDjoJEoXRk1A/QD9DSz0kbClH7DZjVhFL6rwX6WxoL0Ys5QVH79hQ
E4CBRVWfqYimY5yp86cJzll3uPANPsKXSYCHOhvvwycy2NnPyxUQMVSOGDL4lLaTEv4lugDVzr6V
JENMnoZDkMkdXySZrgrQH0GYzBcCoxKb98dFZpWC0sGU3Cmx+d2TmXeTgpSjdxcrhAys6byIq9YF
osRQscLB3bFTsiAT3CHVZ3L42d1yeD5GepEU+ND0bqLSABUI5fcMR6xp26C9ZylUZNBJ7AGKZCvd
wpFFwMbMGLswg1F25c+5Fys+SXkqVliaA97F6lraJ3XXkAthf0zGKWtIh9AcmB23NqSBdTulXT9N
EMRFPFF4pi3nRHF1L8iuC5LDGfdXQ9jR+VZ7GwRtG3/NbRajOU8QFCKzFJtpEV/ncJLm9aCUkGrs
rVyfzneLG4r4eCOVJmQYX+5DamPnoxNGiqj+QzjTQxoilI7zGIhqPSYPDL+JiAoZ1hUdZvd+LFYd
lO/MlqzmlRhdQEevfMBpkM8Y/oZp/i00dNbMapff2W/5o7z0hO+eprpOr3FrtS4tvVxzm7Vqn8vb
OgwmAj1B1g72+T0H7TIZADvSu494x4xFTcpX/3JQJCSSw3MCP+u9XZrJO3aXMhPOZpMbjie1I+UJ
W67CH9ifOnOqWUnl6KfQm+gxK5srJCSLNAzl+rB2x/PrC4eP04HtFGr5cbgHBeU+FTouHbUbZosA
9Wlu2hc4t2koGnWMvVA+i18zaEOgoi9oUM8GNlOOEpNNUByo+GpsuyI5OEw19pdnAu1Hy0+xUqao
RW0TIc8VQOHK6Rk0XUA64gNlBh9NowJFEX5FWVfUGeLobN5/OsmAPZNGQOaqFvo1tTo8ZBatzqZ2
ZZ/oqhn7KAX8s9gd9TetGHVF2WTqeVWSzMdg7I4PN2HuBN48NjOmUlMN3q0EQ1HYf35r/Q6LvBT/
ixwPhI71YjO+URPYPBvuQvCsaXZCcg5RxgMN9mF/xNrMVViHf/eFgqtOeDmk/uLl1E06l2NBs/Mv
bMccM+2lJLHBx218d8Kxq8z9OCVMCnz0VBNsBlIhgnPtoWVDWtxdKRVeylb5sgILSupvIQ0zrocD
iORbsQLFz/rinahOdEKhV7gk+qlZhsBMrdtsYBWeoqSlOb5poMUIzz2R1nj8QeaTZ6ZlIWr9R+g0
icBvHqJMT0XGP+bDS88lVC8WqsAOE+QRDEuv63kAAiXj21jFnBt7t9F44CP5kkX9DCzaNVGZXc6I
inGRmo8iGNivtZK/gMQk4TEduI775AL7T1e6laViX2Y/sj+XW8vaEkfjOKPgtrEO4HGLEmFHdtyL
FEVbc3HrW46yJRy+NaB82249LIKlw//9uDSsHFX9hlN5JA6SSMciuPHY2evegnEnpy12XtJG1Q2i
KesLrWkeLwxQCD/9m+37e2Pn3DPJvsGHdTZc99dfOPWJ3VGK6k2pMljkGdkoG1NvN2WZhNPMGYz7
CvrLoD0XsOSE98ii9UENke/6ym6Fot/kMScorMYXyddEY0jz/9b3AUVVS1L2tJ3Eadp2WlOFR9ZZ
judWZULk1tEJoquPTxuhMYUtsFIrGTjd8bVbx/L6GOhwPmPmFWHAtvOoASLnW8DqynHdPr7Zsduc
XojXcqQHTiA45ApSQ5OMT1YkkeqOKEjaPTljf0qEnHZgU4GLR8VIdX/adbdnmkfpuAUN69PYJDdd
KrpnrTvQDyaaH2UtngZOFk09zDtJk4OAbJQWbOYOZWiWsgaL7SaDBQxrGHapZ9rEeWtfBvVqHRo2
KxZsmbpHbp2BZH+BAQJRAFhBsXpRyFFIZdvFEyXawk7rydYAVlOylNcckGmexIOlt/2hX2GNa8ZB
7ijDhLTv5/H+UHiaQBQhmdpYn7+8Pm1S+Er9ZyI33SxgSPRMIjTNAn6B+WE8DKNK5zQu6M8rfo/R
7fbWKqJerBgHpdAiHIuT9BYYvirVs4O/gVgkj7nP6I5Lfyp8VoG5NIQS3TE1LHSFEwkUraG+ZanM
qY3RewFDt5BWNJjxm0BjxqkDlAuniEP/rAUmBD/aX27qikcvWQx7+aqx77SKds43V7NJrpwdlUzk
z3n/fihhH2Bnjb3k6QqHdTYwJTgqBBqZPoKWjbveODtv9lrVIJLxHP0k//v32fadwmR3Jbrw9B+A
4QxnEzZ8cRI5BHrN4/pyQ/frXxwkwyE+RwohsBHe+qk/L+q5lmsrn7c1hC7jn8rtqYd+JIbQouHx
P7+Q4Iv6w22I07F38f3u/Q/xMeoUlbU4szagch/mEUdWv9nH2jT4mvzeoYhSThhJlF3k/7Rjvs58
UJTyzdreuoKiMJxwTdp49dt8Ci77t/xYPZWx4v8DprFE9byd81GL/XiGEXc+WO0ru8T6Mi9EnPyb
0Em2gNi3NUwkiMIz9ms6DGbX4oEUK4YavRWe3kC0hIKPtIBqamqmSJmOUofCMmaF75weMPpVySml
OfV6+ZzxGok3Crj5OPAaQoEgQmbgKKDjzPCDTHv97CKc/pyVXvNS843eo/UFz/0fGDdfluNeDju3
qcRMNZ8wQWbwGnY/b1r5PyKIZ9x01ePCeFgF8/Bg5roe8tllWq6toqpvivLe2vWepQFX0qqO1FGm
RlX0HZ97oo1bMVsjpqMvFlIHamt+EDgtWuOzzPFn7H9xgmvSPvDlG1DoqBQpamZnRXs8DgiLt5pQ
ZtGfD06N5zaryuYBDKYQWL/izjF5ZZdCcsX2VAoP6Tq+/kDdmz789FatKcHjBZCfWIUOHb/Otz6n
rthNVAUNsWuP+tJ0Tp25x//bOALWYTtNDC15/hJBq3ah0mqUEMBZ1IrGX3Mcr+83amMe4uhk8WnA
RDGNvn6NzDDCeZtuVjmb8CRl5TS+eycIKWwCLRhuRklq/qZZe9fdx+oJcJmBkjLEWdsOHhItOuOE
SLVhksvtfjc2c61SWGTYKGglQ2BDGLb+pVgbVdmumZ3RcJ/p5IswFuXtjtuJ3o1BaUTKZqKO6SpV
ZqkXkusE1fs3Hpr7N5xZfPJ38u1RCae/WhscEalvFAxqqW6t1qPuUnvyxL9cZ52yOd0RNGWsCxoG
andhg8Kxq/Z2GaL3RMC9oD9G3qRwyrchCPAvZWeSVkwjlRKY75VaLbZYTK3Rw5lxraE5bRsiIUGt
89G6cJUeLdjFMiPXv/v0S8ezxHYQHY4vOWq6FH4hBbU5F+eWgBTUV5qb7gkiE1hzz8TRDN1nDHps
w9hbeGqwyxBYPIDhbIFi6+4uOnXxKDp526VrF2DANMwyDDELmL2pY5LGV++WfJ853UM2HpU129SP
kVtqPK/MxPpUCbL/uQd2F2dhiAEPBV9U/bUo3489KifS5beRYiJxohxDDZUdvjpn9Bycq3qWXo2O
2rwOWlt3TVnhwi/geA2m5OayVLqfMvDCLacPu3c7ka+Z3ZpR/1/rBDJORabHDeIL5jFd1t2mq57K
lLQqC6dgpsFlrhIBUkZCYwc35keYaTvYgfSn8yGwGNycKeLimzEcF/EaDGQ9MzJKvcYJch/mLmNA
KaS2dFBgzcp8tcaLExRico1xxXFF4KloOIB6TvuUIg+M5tp8TOGfKB+6JLJ1sSygryKc+I8BDAfJ
Uklkac6Bm1kj5RmDO83jJxtulVBL2bi+DZKuZFFCxEbBbx8hy0ttc4w5H/sxvOIbfuMwiERnf0Bf
FmEMXtOeS/pU9uNqasFgSQPERLjf0E+/a5xiVE/kwSaf5KJuy+vIYMy35YfeWhRFE3fLxx52dBZF
OvnxLH5nn5zX32fhqE3dsZcof004mn1LEshWSDPuMSXIWL98SPm5wprJO8yQVp7UlLH5ahqobbEp
15DG6H/opsP0sLI4s6Dk4LrWRY+FkIbjF776gfeKMbzKAN0xWp9hnQRF9R4YHiVrpcjkIVHKUTHy
o91uxRwCRI4k8pfDSzmL8O3H9lqy6K7DakfZl4vXdzQRLPZ28/PAxcYBWDwFGKAyBAbCZdE6+xp6
lrOIWiNPxTQry97RtmnFo+fMnFbvEO+OJVmEKOcH+1bf4cNkzIvVW5ymotAoHlV6WnLiLP/Yl/BD
Ky/OUnBBuPEeVeZT2jNCQVn7WFjvusGqxWhUBjsNEP1Bl37KGYiPEh+UkkrjJJGSE7v7exF3SBKu
v01n7AAaV5RqP35alDow/ffa8WsZk/9IaB/gZFAImOVnmBDXHNlxYc2HHzpz8N8ea/rXsHLCZnph
n6SMQkcVCSbO4fyoTl3Vex+U5Qi/j391ZQh+w08ji9ZefvkEYKb1rJZUjDvF7sBo6WwrgNHxHJ2+
ObFmB48tCUwQ04cemANyoHc26d+9gOWZnFXSCFz6ieCfftyTtQNQikPfRTErIddvCzHKd9mJAS4e
ZXUt1ZFbe2ZN1iDg72PdmWTZcKnnlD0nMhsV8MSS+b0wcCyYgKUTV7cwva6vVmQBvJn7aSQ6GrdC
fj8UTWny5s+/UXnnnQdX8M22NRTr6Ei/OF1TP9SF6VT6M0DemcdrprzNrV1/SFnYBkJZNCykXYPe
nwQGJGKqt4lANlQ9Lb/B5HY0N0SDCG9Bogy88sdEBUavkg6NZGqOVHKuZ5MBBi2zIXkgxDFTOXmc
AmITUNwt4VONiD2yG0GhSF3qoTrpLHdur1GMKdVqajwFODY5O35VMHywj0uk0j0bFP/HVnhydB/l
IM8FIlKn00tHsG0hr1cq97EX6aMfQuFDx2CcwhNZ6StN1W/t9lM4LuSUYQib4ssVKNfwbdfoTszW
V7BOJv5YIK9dHJL7mgOnD/pHzT8s1etgljoTt6z+qFEyvcny4zHbXuijKuC9tFFRq36G2F86fqdx
H0s5FiBmQ/8k/y5K4aMgGX6V/fk0vvZNC/2rLrckfDu4JRSDOjx2n6ZbH0W12XxuiGkN/WddfMR6
lDwGTqcVU5JzBgjef907+GkYkpONSz0tXCWO2ZUVIBypTFFjqtKFLq+3VktLWi1/YiX95FUqKjSR
jH0NU4XL8smNsmJvh/aXdjPWKy1zwcj6uiF6SwP8RAz8ry0y+1djz8mwkAHppTIgVfAE75Q/yBRt
7b4vlt/O9g3IrAP/r7F1+RUtgMK43Yt50aRn+ULs1T+/Nn1N5i3L315La515doyyiCYq6vFAKVbe
EGl+3hFwtBuGs36L3/Ew9lYlwZhrVZayIPpJP7nPxDb6tsWXoknbbN6FETeDjeQe/wP+CttCN0zK
MuHHozG5+IjuivMeTBFz6wd+71OvP3yl3YsxwYB5hrMgvtkK15AvMQQ2hAefBAcMrB4CzoJpr06U
OSRFZIPP+Tb018lUOwdymoO/uHHhlX0vydhlVO+XK8DNOeaigneL2j4aJOQc8sQmVUHleg5MVi66
5ipfTWk/+P9vmSIjXH7vVnCgMNWBrHai6D73I6I+Gm9/iI81Rusa0gOntcr8Fm2LelhS4z1vaLk5
3yr7/nOQcONvo2yUbU50PTQ+Hn/9tKXvWipA3dFCBOYZnfyuk8vecldKM8myuwWnd8JDG8Nn/HwT
ijVIwDJiBXk35tcj8X7782L3L4zICLDZCfutusWrTFqHR/GRP4zwY43kDtxDz32cdpnyL+OsETnk
s5jgoo7mCRFJ+Vpt32uS/t/IRSQEStgnKa7OZmD7rIIZ1HKgeco57eGz3qy9ILernZyiper0P02X
WV3IqqnWxmTZv9aC/YBwKvZxxoFRtR3mqWFRm6Rn1o517S8jl3gGq/NeKf2KVckNF3Dp4ocnmt6M
Btc+G3ErUB0CBsf8ax3DrK3AeGwAUwJ6A5BWC/hT+3saYliJl8D1XvZN55da9zZ8ZBpD9gaSnMUp
OC07DDwdPzkPT8bt658o6/ufQq2kRiXxOylEmWf8TnRCOWH1q+bKpMRWsVLW3z5HDtjM3mNN9usa
uUQTMYPHoZx1lEx303n9v8jcFaNY5kuXfeEgQyIrOh4GnMZY/Rl5XQUKDQSAKtChpAnrjoMoj0wK
EmQ3DbX1s9KAOvYvb46nJpxB28Dk0sZ/T6hLr9PZAO4pCmk9fiFYp7iXSrQNbcda+aLsNG2UunpW
jWE9adfllNobwseXeLFE7m4m5J9AkSOTjmprsA5zdgHBeECsMD/XPa8I59DpywoSJ1qjPnHjYWM0
UyrkYYqXncOTOik1fIDsLGsZHbgk6JvEpVrjpwYj5FX+IADDwppi7fmFfHb7lV2ZUIx1LFNENfh8
U2QrqvVoJ4MR+dU/CcQx44QbhMrEHUSGfy5hnnMbmb+bIME6uTBRytSUgeP4bv8R0o5wP6DbaDU6
sXYSlATQPyRtm0z3A7uNy2M4EtnPnGjAT8llihzaQ97tXU1dcPppIH88VKY3A57r6RENNjxzBJmC
c846GL6cOxAhAqTh6lHZb2kJTui806pAXGjGfCpk1G5Y1sQiGS/nVwqfQb0VPs9B1dFa720GNYvQ
WTESYzEmCWZm/HA9FE778sqT1/GvYM88Tp4oJrcbP+qEPityDTG0if0ZbnVTwEgBcPwUqtFMA/Db
4GcD1ocIm/wdrIIfe/fY5dqVJCyI5FxjSXsZKyxCMb/yhLiQ6SyiS1TwB7VjIqPsnmansQrDMgpj
iYkjiUUzQWjRoQqes2XwtfFn+HaZmiRYl1QBYyUDidz4PESx2CCUUoP/VZiYJ6rW4XSld8zvge1K
/lsd/o1Ao30HU8i1v/538ShYKF84sbJNzhqNNxrnjps6a2uMwwQpidAqoRdLjE6Rxromgup/Eg0q
Yv+9yhOpGslAvdQsO7rSBmpudPYYbjwuA5ygr8RLAm1BpCKvJ8CVygTHQiRVcjUhT34yBuZJjki8
/Ejr3C3dkgiS0CrrVx4sVwtyWEI8m9N8VI+8TS+93ulJ97h6RK1Pp/NU2Ta67ewvfIANnJgP7IoT
7cknVLrJGvq37fJxn3I7pCfezloEiVaDVwkPXTYKlQia7JNrIDk2qmWwDZoxzmm1WvBhO+simTXJ
jRRl2dyBZcb2/tmRJsoSfnXXOGvd2Ix8jmLNcf6jBtWN4kWRnSyCJ5vi1p6X9J3fhPLJgKAVQQYt
c7LUvAPvlDtZ4aE5gyf2Bf0JAyIbJ/A3CCdAGY7wl+maiNNPBEePX/3g7XCXFYlrfZCuP8OwF+b/
RRAK8g8BZCPv+cD/Uw4WXIdvTBPDwU1wLBS7AnbqS1m4Yti3bW04h6TM50VFPnYFse6Tga2Ekd0t
MS0EBDwytb0WiWl0mM0t191XyW1NEp7if2py2dQYgASNjNFCnUV77vs4ia02C6NQM1zp34hK3U0H
cQmqkKW5muZSDkD0vznoQieFE+fQ5YoghtmBn4moUAWW9QvB6VgcpGLAlCe/bIpCpJP9PxlVxtYN
VOgGeJG2gjiIoD0hR90/4QppmBP69XmxAgd9aqQCfgj+b4sGnBPtUD1XdHde9+phvbABdzLSZWUo
DNhhxqsx3Pa6nUkLOKRrfmFqu0LRNdJNR+w/selGyxP1gykvrhULVTSsnxV7whP63gX6p5eIm2Jb
f6HkVrsNokuZ9hinC8aeIfkKpRumWwjhCCMsUMd6h6o6qtQSE2LbALLK49o7jVlEwqSJhzQYfT+u
3mK6IEJYVPQG6nU4M97FYBNjzcZscxYw6GwgANLs6UUlswVAWOCqDJvb9x4kc+O8MpNFBtlMt6c9
a1JTRSBFRRFBkT7QDdH+OW2zYY8dCF43BnfyO87j77Y572wFvKHFIc9M3JZW0wndPmJ7t12Yutzi
4UIJI1dNUZm77fROIi8KtsmKxBxUPawTcsylRIpLkXv0Jq2vQpn+c9U691HiZKqzmhEDEmBlpSM4
laAckvrm/rQTdndlfinOLv+LKgYlW3oGsdEtEPKRUwdEu+PGLZYkiS3SyoOKSNtJ8NK+/iQslOAv
D7vOHOP57t02KP43GZsC7/+lDEgavmddcYYEKwhpO0V7JZeKwUwumAWaJ3/nKdoV+T3C3PQzS19T
yFJ82Jv/h9GjbOkkkvPJmhWrM3QQAK6+hDQ4ULywlH/jX7fYZrZ97ctyqnBhzdZhNk7cnPJSJq2Q
25W5rSavdIrzBxud7D2k+XATjyCLNq6DGTjoF4zA6A55YllGoE/NDvK8X0Vh0+/t0OIUSl/8qdVn
jXIfIm+KaVOAzpMbYAn0v/hELYjOzHSw63dqctZojvRWG8v6A5vWG3dBafBh/VmdgRt9l55Qo3Mq
PTQqi6OoW+oyTHd1VU5mi6yBE4qjG7rKrJt1opI3/GO/fw/2QwKpjGiQd8Cu/3vR5s3Jmx8dzDtO
t/Jl9EsFoJWv0C6cGFSVorFeAGliNnmWzvcZRlAvhDj5aheqsNzE1rwIjfkuL8OS6ngdaOlBaVV+
YdmbSnqD1ME4VcYpHW1eLnM/B8ow1R1TBnX5coae00exH6hFoMhfXimm1aQFFd7Spt1S+0WkpAsh
41v58Q4n7hUNAb1Xx0WBKda59q3IqismPCrpzsddE0lnjI2KsEJqOGPkS19zanJvOMD//v8/Wkdx
ODSVg0Bgaf3/51inZK8602b2AxYkvMrWjP2eru7bKLKaAgzn5p7ycoYsq5oQxXqxh4PEAlZHIWno
F4MZBWlXdocUMjIzGSKar5zckwbvIFRjBRBTNs8EN3+BJaJoHlqeC1Cav4lePR/yRQhxLs7PoZ9B
ZtQtsLi0CdqqqcJYWznHdvRVs8jSESwKnAMVvABcgiSHIRD7N1hMnVMu0GmAXhDXOts/5ZJiec75
N3nVvKsPgD6s0Vfz/SEMHltrXpYiyCnKYNbkIIoocX3OBUuK1Hww8z0PR/9EPg5vx3A2DpuAVuzu
ulBzx5nK3br6ZFnHslztKw3N/Su6yWv55Dt8T2RGWJ9HFIcG/iaqq2xXcO4twUWXwQv1bFnZy3sp
3x+QyGvbErJlJCmvt6qEfwi8c5t3ZswSnS1ODjomrKX27EoPd17UB2Va6/HWm3T/6nwjQdwUCP1r
YGbwlVo3K17CUyR0dcs0cO53Ur51aYeNh9MzEo6y+egE04dEh7NpYFkImFUSsl7nCEtRp1SgHrGg
mQXrgcxKK7WvLRXNqWe21MnLAzz624+Fyk3V2HRTUeAUVk5tu5nNxCizzUaagyqldHOSqm/K4cVl
eXvtkoAfOmt8U4MztMlkeHctmfYKZ3QOiqXAtYnrz3lheMqFISq5rXOS9P0G8uoSaNP+fxQk0yqA
vpiW3K9mFzzhTBSwv+K7GsG71eGy23tVzw4er3VQAqHvUAnNuUqTkRUghRPt5iHn7Hjnr2NkU9o1
MsERaySojW7vTaYprep+o8/cSrOAroh7yMOc/aAtd/KLOOTHP1LwWaUMwx7zXf4vX0gVexkaFNBb
u7t8wOWbK+DyHytJFOJKBWCyVKWrhZc7EOW7y0xcwrf6C9vepjg+iOHFrz23AcA6popsfTDSqsdn
MottKEX4BzWrswDzroTyTL7bidr3sMt4fEUoMp1i+wsvrjrbFf4IWC1mHQ42xqCHQXrzFe2tb5iW
GFVtVJMFe8jAdIDh+AjxZhvNUb4gXJV/ziFWs4WNHiEMZhK6NIdbi5NXHr8EQfneXvkUhCizFTTu
QTBjVbaJNi+NCC7hC1jTRfM7Jz4cVsJH65BFCR7zNfqWGWcmhUWgwO8a1xWUZf1vgbl+FadQNcDb
9Xe5JU3eD+MbxYXcceDzTkfePicN05uIw6GIip6tC5RDlIRJUu/c0nsHL4VrR5/5PzM82ynSGV/t
RCxIlY4jaTsN3rlsB/jOxETNAr4GQXw/Q8/krElxp58pBJ+eqNbYc/dBMvOfP/GdejUus1smxLG2
owa6o/LwnhYY1nvuG5t+gucuTRohW0+3+awkVklEUGzU41IqmU1gu/3hWs9fmOHw/vNCqv65+RH6
L0V/kbdVZtYdaYt3IqAaiMCt/9jXcx5AtwzkX5DXOHQ5KiMBvLk6qSYGsvE9X9HI2DVO5kulmCmE
gd9OuktSX2HuiyIGU5jCDYSBsyh21Pv2oGU9Gy3K1AwrwHIZISgnmYR1OICdqgi9m582+N9euyET
1DQRLGuZZGk25us/ErgLkQVsHX1u90H3xScjWwKRCqL4n0g9uLUkyyHgzyB2AVYTpVq0LsmTxQv0
YDSAL2HVigmQlezwBclv7Py+BThfLs2CDNh/sVluISzaqzys7A6lXVdzpRtDszBcStsi9lRsuIS/
7y+IwUVm6yDmssGqkoRGfPzZ8O0unA+j5FkEdK3wF9avjsORuH0KEtBPcDvA1LrgrJscrXbe7Kpe
BavUYqZLvW3eN1La4PoIuAdSbTKrBVrD3Qjnp79C9tAq+FmRXHmca6yF6F3/Cp23TmBgQ+6n0kG8
eOtnmatdoeE1SosTqfEjJ4DAk96O8KibLBb1Qh3eg/JIJtbv0c3JSAEKR943uUxWoJ+JDPC7agEG
do1VUCX2MfJvIGe7hNaNsqFh3gr5rSixtCB6fkC3XmFUc1dbtwBTwnf2iv3iKRkiOMVEilqEi8Vl
ApjiM9UvLv5nM6cnSdpiYY/K9QF9i3zk7RBYcY+B2jVpAOiGmc9Y5cuNp1y5LZLciPw65MWlQ07k
B0TsYNbDFlitbuTbyDA5Nz1UGDzrMjzjDf9ZghAMUgL4kErZxJXqZFE3+Cow72j2CwDss8P5zVFd
7lvTTu/ItXHD5JSAbP4KUGHbXIF5qklv177BOkvPYaBoBUnBCpjTtcCqN5BsBDfqYfxL2cKOOCeA
phS/lEn5a8yWaS8gAkmgHmx0XO0e3rnN8CvGedRDIS//EHo5VUTUzE/RCRpB7rXNJvgrzyioit5c
d2Sn/6Dqk3YQzc0w5hkP4qIlJj5d/zrqeY22RO+jBLDsO5nR9IM8R539blTz6WlTPpkc9DuNmu1E
UqxEqdILv3hUVz7NMiuJg52tsKJ//t7RH8+aPw7p+MHIFd2Eg/8mYDbOrqqsZrNBQDMp+MoB/ROB
UgmP1g7hMND2gxYGR9q6F2+LQZS9Gy1c5uFho2nW/pVNQX+BCRqql467bDClMSAxr3+jLbOdTMV+
IPul0OMsbJlz23WyMGNKKk0BGND4nPEZhs+30UUJ3aRxPzuI9ANShy5wwX8JCbjC5tR/RC+bfDZF
K6SXqxvJcFJTviy/5ILTQM0t1mAkquJ5Yg8ySGc4nVq4vOjbQNnyBUVRc7VOmhtirw34TP0jGeCQ
zBGl474BsFvxnIiNUb1GRXTiKjCRFwkwBEgH+qGzNJ/C/tB1KqqEuVNYcMxM1LMRVGjDc2isqUN6
VWHT+0WlK9f1ziDd0Fwg8rwZuVIGmKrNdLa91VVABbvot8QoWt5ooBABtdXIt3ykb9eTiH5PxnGj
/4uKywdvpTl2lFJ9oNP8a39WOX4VrpCrLLUa/947saIaWxQdAeJIOs19MOEd28U71j6yEi7uQ2iT
Tn6BR6kATeT34WGa7MPY2P52alabn21MmH9VPbPenb1+vtFGoSxQ+epPrETTN0Sylq6BBPcpLLNA
idbPYlWxol6uqPAm5AnOUM/LVWs7WpXWtecL6g/dEELqaYsekE5W2dp/6MFvo29d6Zn4g4JokO92
Fg4so900raIk/uzqC+cxOH0N4QVf4uzrdingc4jYk/wOlUC6nlMrwuxgOofRpQ8dM8oUyVclDvMR
o/kHbbDnRPcJNwrI8/4sAdaZA3b2t3fRoMFVkbrUUPxHKNGx4usblcEKdeajvDc+dXwGZNJVc3kz
2R/ug0IdAs7jCxvlydqobkzpfJWGoym5BIW0Aq62w3ZLRXXhqiEiWWQ+8jhTJCugwc27zpnrTiFM
tkjc1q0sw934sOiMex8rmi99rvkbflc31ZeqWH+nCS1aRhGj1p9S8s6t6sfdD7Q8NEW+vgswFZYS
A1YSvvg73gk/Se0bAEBSEdRRGtG40VMPkIRK+u/gimbSOFvgUfqXCh6xk0w8lwvTn2kKPjMSqtRr
Hw7wN5753t7/MOKDzFbpPxCKuI1H3OmkovD1yvazVJxdcxSk+gCba5GAI6oP2jqE7fWZDHlkOvbZ
Wlneinz42Pyo7Z97f0w6ImZDlcz3FSVc6yJBH8qOXTJYTuI5Ny7CKIPodX0yAyUhCi70xqpOO91H
qYvL+fEBSZEYRXTZ2t0lfpwsoyD4S7m4c/5PupCQA+2WPV69UI/Xcdui3wd+EEISHNlBIEefBD4D
VxhYuIcnMy6cJ5AltpA2kcUd+9on53j5goiHGqKAI1nhePIjR4z9wTmEcUFQNvx4yrDRryf53YeR
GOaQ0v2sYspph0xYXCrV0X2BkQqTLEUfLA/0BtgYrUoDg00EvivWXNaBdkFdidIjWR6AQ4n+DbEM
YIDk9yl4WSCdqvfRXvnpqpolfvIwyrW2thTsJbl9L9H+I/FLaA78i9pNsicp2svemyst4x9O9w23
468vpo1IX8FXFLM7STJfdXKlXUCzk+91T/fsHU1CIAJhD6FqeiuERG2EHmcHxY1RkcTNBfQp47iS
cOT/URdNVLdc6di1VbnCy3dSuyJ8kP8HJQd5TP2oZruVE5wgfszOrYp+gT3waKJiNnxz2LHe1bWW
TqCa8+mzRXIwC1o24ygnkJxVIBqVTT2oe+scDH7dEO9Z5E0/rpn9CCboiUK6+QwH45QDSmrb8hj5
mGrwZMBVIaq0cvqjUxZ/lvLiSE13oBZlqI0M8fs8oEu+JpIR8AGx+M9VG05xeNGcBr+QlP9NVQuc
/si3UnMXf507ua7Shj3wP9/s6W4sIMkvM2AvZ+BGeIZghLnb3qNsQQeCfU76QeW+YIWtfMHuX+vo
P3OQy0SR30on8r5/I016nYIjpvX73BU90KfrcCnPZwnkA20WtzJJ5OpTu0U0fi6Ve+hYhDMZ6MpF
JjHqzibVLq5fRj5zfwpa537vMd//Q2OhWnsh34nva/wEamWplBuZlIVneP5PicN8bckXFMbywQ8E
dS3xmNOzowTo4dS2la8aVvHqyiRvwUB1QEI5epU0LTDk0Tav949YKRupt6PRw52cK2NhoDWd2OLj
NXzslb4gZiCM1lAhlUBgxD7OMZvv7CitCq5LbZKrM86V1v/bep0/aBK21zzaPxRcJVPWrleTLqVW
QRIxy/WXSEmv/9+H90+D9ghnfRbVxgVUU6fK6IbFVJ85ZS6WzezZz+s0dwws29dCFZ6ULV1otkhE
4AxIB3LofXi73+AtOH2SVZC7JjaxliNeTPvGFEImHfqTbp93G6xMXYzjdErbuk1J85NP6XkzpvW1
lTrsSsI+KMIhQoQW4n1aPpAJsLbhH4kfA2NkdRaqD8ibTCTxAxCDkFg3KJu/NfsSCHw+Xs7VDdUl
KBcGnGrWCzb9cFmkq6xA17f3Yux+TdAzTWtFKPBe/xea8Xot1mX/Q+VuoN0UPIbBFxYYUM2MuRZF
6DslgaEEzlYFKQci9U7V+dRaCzhfNr67yjgHMooYBoMkvilijYzzkoOfQ8AF04/oN9sDahOQ3xcp
89tZ6rLBsaItAr1/XO8Lr627HDi4DRv498ftkr/Y/xbxhqsKLratuWhvlczPv/52+2qyTiC/EnHY
PjqN6WIQlsso/LHmKADSLNepTDZe1nWKdRm8TyHeGFY+PWRU62HJJXgIPXhChPGcURfricXJTEx6
ClYluKNRoqAXYQ6k0YE/XKtM96AEUJi7fI0d4ZOr89Fd8omoG5JmXPt9yMcsS2PQ6I3F7EqgriVJ
ZlljfeT2nS+91DXsmQ300YaduHyDPXJ83U3wSxhv7gitmv8B6pIy3wZ+5OOjB9bQ4pZDP6sqtOyp
w0e5xVBJfoHhdzGl21JdUiZyYuBE/PTq+TfTudgw4788Av8EUIrVwg+qB0sEY4i9yGwSM6QLNajv
mW4nxVutt+OFXKUIrMlSPCcctVUH4vInpbhPjy2OBXuEtrbI+DiHFRjNc7Kw9r6tXU0S4o8UDm6S
LoHnJdgG6ypss84PuRekG7Tiqy4I+74a0bylHW4RNyIYHji2f+yl8GsHn3PxtCz+QtvbVP0QxSgr
iAy0xQokfZC/NDwggbjL0U6Gn2kVevOyoLHQKFOo86nYzGcqmRk0JlL3i1rEbZSR4L71++5Y82kh
wkxAr1sUh6fLC465xTpn9GmhYckvPyh3J5VvY08n1K3AsxY8gNp5KlHoTMyo/uziWWbjsIjvqMiI
qJ2U/eH/kVa3QV1dQfjYvxwA21zMVFtiO/B5RtBlhBmLHju2iUk6+y7J6dVxbqVupHUr3d39Ee7g
am/iXKWNpajchz0DBYRyZfAM+ZGTv88PB/mzTvEIsCsqZvEpHDKCWXcHigxHWLMFDiLMBnV5AytY
lBPtsIjXEYbtiSrLH05PvHIdyjZharpvGkap4yTXztCHTWLLl8s3ZR16d7rgxxjKYmbWlLX4dEU3
bIuV3gcjX+mHmiq+QUAJ5s7eVQFwGzWwGJjuHG+vRnmPxUK8kPxDCLzPerAp0gL0rv6iGEfzlEW2
+jz0nlBv1xCQG5P2u0arQ4ZtBzL4mN/ZEtl0jNZKK8JupkgcYzCsjGmbXbuPjQdD9p8WllTmgHWX
a41B4jLPRydI+asGdi1v6VvX+d1t36UX/ZKTfW5ze5qm/nT+0A8+qAB4+kMtgseveldmDm8fgyDT
sABCvuFC1gTahQx0jVunKnxLvxDHPTbyGJ+X/EOdqDWq4woGEnBoqzbr77BXq0JFIMgxK0Edw0lq
/rq73KuoTpiQQa41bQiVLqfSGD9nkmpRGbEv/L+LhyuIZKSF32yLwRTfImiWNEho0ONEAqUXz4kn
fh0hhXL1VsAi9aoCLoScGt13YkFd5LZ05Bu+tWywdM9Bayo/bjuxbLxqIYDPS/rmhEx1AhCK0oUD
1oK33yVMkiD8m9G2ozlgkluJa4zZEVqIyX8mjbVg8q0TiMSJWr1qeAqwUSfvPgUm07fQ7ncValR7
FSUTUukLoaeTUlqZbIbGCR5M2+bsDW2hYHpR6kBsG3ifa1S7rj7F2TIKSdGDWQJEKA6y7vIhKJLd
Nkf4Sl6NRUju26Mu7zelmKAN914N2wBI+vvtrMQTw1ngIvwFy5kFU95cgM/JzxovFpS5AKZZGO7F
3MJrimGVmB34UlTFQvUeGWsJvRFBt7Jiwb2WVOyJdLoNjMu0xRZ349ZHdaPT8x9oEqpK+pa7mMJD
gxNxr7I+Hvil0EqYuMFF/dqbI8CzXR9SOw8GPzm0direALRdrVg4Zo34l4o3mCV7Ii5cjCmhdYrt
Yoz2r12Gn5hZqLmn4gH9hOPqiz17u4WtVM8Tixf7x6dFKK/w4D4H8JgWi2j+X34Lda7GU8GTpc8D
skYpvtYIjZ0qgo3Wr54lc9SdHpUKO3ojAM/C34zUFY2Obm8Rk3KcWEivIUiLd/54SSUSBfI5zHlJ
AZVVeJgtYjrRlURdHfPrpnmHtZX21TnbLcHbNKrczoizU/oBuYHV5M/3aSfs6rUlD7TWgNRjNheP
hzXzFuD2P9noZgw6bnik5fLvEL+nfRTM2UOL875Anu+AQ9EowBrRtI407H4QixE1Fzth/+hUF2y0
YMo83LWXNNixXasqpKblQIam82uZBLZTteX9SOWNaCbDR3H4JNt1Gu86Za/1zcsPvtBwspovmMy1
HeAKfvu58wiudHGgH/4Gi8dcYFzDxODiAk85RL5HA1+9YURzZWw+ZdxjH7li/WJDLZcSAWjZ4hHf
KPOZEEUXvyI1JwgYVyTJPElnh7l7y5QL3ekQ/hokoZqbYt/X+xF8JYn3IRk4E+cP8aqCM+Cl/A+w
94vuANy1LumbN+EkQ0t40O9k34Ad3m9ruzS2rUwBxBqlxhi+liY7fDDtH7MPFbcdcAqvdBujytic
ldudQzs8qvGdRMjrKuEkxmKExrKUOI/mBN33htMi+4521+rgmW0YSfv0NHe5icei9RYZwEUplgkV
exRJHZW30SBE6O1C1ZQzX3I62d7ifj8vKiupGgqPhSvGK+OkrBLDCxMGTvPtassVxLTEYiNJeuxS
RMiK0OgSrozBMJ1zLN5ciCh8fW3wPlJ+Nmu6MnvFu/c4KHPYLPdeGnG/d/lX/eSmNgJqhu37de68
sREr2d/N17u9/LPqrqC7lUUvgCmMc/foj+BOblYMSitiGMsAVX6+C+IouXAyB41fosI1/t29Fno/
lbg0ZOFAJ8HGwA6kJzp402nN1Z0xUyYlqkrhocshIf+6BeCRcH3lBDG36bIDP+uw7J9gD6/cDJCl
jEIzsDhOO4+oke1aEfDlWqNgsIEHMM0/vlpTnpDJGpbuZjYNhodSlaoZcIU0mNoaFOcUWondZunO
UJNDm/NLYVAYicAjYqujEJUdSr32bUKrsTXTsbnmFNbuRVFy67YeBSN8r/vmLQ54+afo5FW0pYKs
rvlpq90baNL71xM8ocRacqkYGl44WZvRzwxnHhgVYG/H4vqFvM0so3Kulf9k8oZDiCXqg1DmHqe2
nwXeQdtG3lpKGdExH5Rxraoz6lxYwjKUc77N2nSECEsbTvR7ZFjNvHZU5smNY760F6ZdiMUA9OwC
sEd8F4zqkcvcxPoA4BWjQU7qHgtZetMGu5R40pRiWIAiYftAVjg+wYUVwLLc6aPEqqoWEGdHDSGr
Ys5emzjqGjXJAsLNNIvuyhULrh3aavL/rvlNdrnOPqwUkEP+bWEHpXvGrly6C5WKDTw1oOkTTXY/
Afshg6OHOiinOhM033CtNS6o8N3F6z5BZKtc92/Wtt5nV0mZdsMV7Ff0meZzZxHYS17EFz+bUVV/
OB19W+v3qskBuZA5bTDr3axATZH7oQqG0E5hKW+USFzkqrknghmhEWq5jKgo6APDlZP8pKH6V7LL
vksCe7JwF9twBjbXfek50ywc+u1C3mJA3/6aLNcoO8tYGeiq4JDqUlOJdxDl/d7Xazug/pSfO1Qc
TJU48WlkF1AJmogzGgWFtsOQKDhZduJ54dI9PFV+jkLwuBmqpNEvNf+iyltlqHOoqCbzNC/vKFGs
E9MCxWuuoV2fo77weP+vQiVLfWGgv8XIeT1gB/LmdhwtH6AcAN8Kgdd5oChR3F/UrVy8yBn/c/OJ
tj99hNHo/fSPmLmo9iAzdeEgLBWOj7wRZ+XSOMdKpSsrkQIQJA1fLukBXIZ8nRTK4UXpIFmCDhSK
piSX/XYRA87P3MV+x0zePGc5vr0HcIBarv30BOndSICgjuuqC1zHOSEjJe+VtYI6zbJSYX7SE0uE
T9cREUHTqGiTcYo8E0SCwbAOxsxC2IEfqeKGr4QzP9DH+24LVOILDB8a5K9uFnW3JCKGrAXY9com
/xxv9StU33itpbYfMdHixB5EDYPz3h9gIrR47D1fx1o6YY2P8/uswz2796+d59zuEmJ8ZA+AfYhf
8TcIef8ibzUxu2Jc8wdEak9XvC2UE9P6up9E08CpM4exqiC6Yo2fFrT5CzOCod/N3sobVS2jPoOR
T67YalUhYtq51JhACCiuqZZuzRPzs1sOxtWkCnafdgk0Unf869tKwOr+a6rSsVqMqhG/VOVReAzp
UzG/HoIZcPZWAf64t+YEW+W7WZ8vL51g4W6qZjOiS5iRoiJ2wIJS1K5k82Uwm486MMj8ofeiWo64
4jj5HIHtZDfEdkWvEU3q5UlmjS4ouBtqjdjcSXBxSoH9s3KAKXG+jsZ4PHiAJRmlfxpBO5eW/jha
SItR0mnzSts4F0ea12G6K1Lyc6lQiX94Qb/iDzlAcZMnt+AP9XIrZVpCO/9dvMEFtJv0B76b+M+P
n8wLNgy9yUDCDPLKfeQ8ELqqDfE5Pv0j74ru3kqaQB2elerX5XSQOZH0FWnbpgdUVDvfpbOLiZbZ
UNVFZxwjq5+6w2QFxnizhjmzh4zcQTFxArR7CSle2DR0pK+/E3FRCRgN+Vz70e7S1XR+0ANwODIU
CvMDFRSnMuR1CmkJxByocGiAJ7IGozKAcmCHRmSjtTbiokWCR3HsvsBUjH/gyZaszRN4jAmABWCg
Z0sj6CoarD9Ul/K3igtjy31ZkDX6ogJu7iq+AS4PzLOwX567ooGbTuZ+UieSjcbDt30pOw549Iw5
fZiMA8n8DyCq6pW05Jsra5SiFJx1NRwXtEurF6xXYX2dhFmwbG9glmB4cFfX8UYSaXOAS2nErrgw
O6olfZWDv17NfpSDCxQ09LBxx79//2K5kLOF7aoBmWPN5bfvkpzozMGmeJxlXL0l8oIJ27/oMqqa
j2tUHedCao8djxXBeFHA5HiK1cL7k9DdfDJ6Rmx82wH3lfuwfs3wr+e+Pbpc/8iugl/DnkhYoFd7
zIr9k75gUCSAJ66EoZGnZqn4rf6X1AJQB4E02mOl06Fy7/CfvxBabKCh8ifkV+YRe9bSLGE7ve3C
ylWPC2q6TZ7IeavkiKq0OLA67cYsJfmkJzcYQxWM6ji66dVkrcqileix0O4BHsHz6r+lIHBFuUbC
Moccw+d2rXkqTNanx/SuRttPhWoANkMsx6d8Ozh9Pcr5pq9pYWAtJ/28Q/Ls9D8ANWACgd52KFqR
HLtAzoZaLMrjOwWJBWA9gcaow8aGFYAPNFoXFrV9+Rdl6hF7d+crklQ76Y7JLoed0jylhjNrwfij
zINbWwNE6Q4EqS/sApJ+p0iCR1ieRDudARpUmNmlsBw8P39wmdUFNW0lxYrJeYkutHkjF/L979i0
ElvDkrNviIKy/lMk+CtKQD2jWVGlR0OAzYffxaefK2m7L9a5SGV9ee9Zg18bMEu1FTv+atA9oXQz
qQcgRQ48YhSE98kRdFTfo1zM0XK6IYCt+kMLnzG+qxFhb69+9m95Z1Nt7C1xkEwmha5a93lxZ8zR
oM94AG+0paVSZ90PcK5iyV4QxWGKzqYQTW0ETcE5WYkn4BOBfU5Toks54H1XI53vFrSCfffu8qTB
h0Tp5auj+tOwx2FjVPJb/KMNUR3FH1quIm/7H+LaBLy0X3qrHp17Nh5mGbo/5JNd17ECt3m3NzeV
wWzE6rHKy4V4blM3guLQ+1xFGkkWGxGGIJ4uwSWbEaDz+bPnEkW3iMmidPB8gLz6ycNImRW8ZxFL
dtS686gFzS5jqbg0wzKzlh2dOVbMPTewnqA39RxCKjl8y8Uw55E15WCGkpNMCF53X38rmBGTWy5w
wO+H8/ttfmCN/DJHLJP4YA25zqLgbwIfOfCUcmpdJji3cszrRSimt7zLAyPkwXDUenXhiQas4efu
5KDelDirLUxpODOgldW8mfy0xk2WL3X0wq2jttohnLSFw98LFrRStdUuUcFfJcBZf/59yFXXjZ5r
avJ/YABblcbWLfgGmZ70H/HHlaYOHTM8JP041cul0Gxg2E3atPX7SEgYRXKQh2zGwze59DK0AI42
MbdNbQQybcEUgzmxZ2ZvvGDbprH8MAK50+fRRwLpb5QIcO4n/JCCbIzulXQh6lvZM4UkDhqMEXiG
w+vTQyx+DjDPpWYRgMmMv3o2xdImwWj0SgWDvPaIhQMTGw89nngXoc6imMdNcKSmaO048XVRaNBM
PyPjsB2UU+YqSfNHJdIrGRdwkzT/Q2SpD8vslT8vtcPBjCd08XEqqcW1sfIpWkuJtpBiszT3qj6A
+YmyCfAuBEo6ZyM91jaOulvSJlt+MuHUnbUzUJfKJU4sSigWX7CRBV5lPX1jHheJycs3G1ZNKoXH
1qyR7A6o+MigTvsZoomxMsdmthKmnoNhWcV84vP+v1yX8JJ6NhY73ERnqu84nzrrykaTCzc8PL36
fHgfXdSebYTsMAS2t1snDh9Ya3yiOBYxRHN2q/va3FbBMKq99UNqL90hg7Zl8r+X/37puzDOfwVf
X9hhnHKg/vLNMcYch0csleJyvLrqne9eCBLT3YHdtQBbhN2JrtlBwJClZ7Mv3UNw0W2/8GTNAnNS
UfIph5ShUBwZ8d2EKxEe32GTcoZguMNizv2u2Eob8D9nGBOZnFDhy2SYCNxwx+00bjMN+e733RYd
pZNpSIM+QiAIcPUC6LugB6czzkF+PIYhciIccg98MofAUj44WyW2bQH31twrlCSUKRncOoLK4vN7
w3VdO/IhSTOFdoJSu3dvXjB8V1mRKd+Afjlgs4pYjrFSh/mYpZjp6KRrk0jPcg7J4v8oF5NwfJ1n
4HAJ13IJQLbZp99mAdApP1HAPBJmJM1EViDE7pSPL9kQDMyEDfPSNdxWDAfM/eHVqT+HQlmM0pNl
AOEVzMQtixMg5k05h29TJCRYIhb08mJomVwlUNbfe5p7fDseMZAIL2UA4drMXKFA36l7cG16sCps
zFBxWoo5q06XhAs2YtHYpixKBap+0FcNNMXWL7I1WvQUXMwVYSPWu2PjOhDY5EK7vPXgvo0pAEsD
RLSbqUr8zS1mKF0RRbhalMU0mk4A6z61BxsY2IXNjHKyd8oeTxzfaMynJo4fy2aK5Eu0fu1xQzw/
o7s4pePLw2/xcwKlM/YpOTOf3SMuOd6ZR6QZttXmcBaQn57ZAA1GOCdQaPnb2sKo+8FLouIGP8Sm
2z7qTVA2KGO1ezVCgHP/swIS4WtRC5jmqCYsCLj+LSeTsMa+7H3HpK8sRiZ1tRrg97QuJUEYeVjT
JwPkTliRwdOEnCNEepQOfpQzebkOIuzheRAOBWH0gf/UMz1oLj2jjhapz0fSz49nd/4/A1LRpcuW
YRyLxXFjL0iXPmJdLuPoLdMGQ857cGD8vCmlaD6vREoRns9q/oVYKxeX/hKlTBWm5bpX6mnjnkCk
jhe9l08NM+gzBRp30O0sK7dfsf+gn5MeWvSQEtjd4+QQN1HgnYHOa0XT3yiTr1Qkd8Xr7aVbnz6R
nWY3piaI+D4Ntb+2LyizEFVqH1zIqYXbo7mWGqocIWtrZy3uUuYFkB10iNmmNJNshQP/0U/DBuBT
iXk1syPzD8/xtWGNJn/SySshU1i7YY+lO52drWhlLnNsDvzV8PDK6K2F9wJFxn5Job13FTZl2JpS
Ddp6O3nK1JqCuPGT0t2lEeL+w5qRixSErmXHxXsZs1XcMetpFxWSYunxLLlypwjFJVE//tdcmQTU
MCyiWWyRbo1/lTJbjO2VinnajY2Th/43ilpbtAPL8v2DKczry+HJ1CAJFHmAa/4zAZKLBcrwS8XE
3knGIAxp2sG//fA8AIu6Ok4ICTbgI/K1aKHevyLRPL4HeG9OAM9k3oVf4+SaV7Zeb4cMf+jmeckU
ju826Y1mESsbiybJShA3jINoTSL3k/r+KEM+h4ZIR2A+NeerfIZEN8xOa/x7kGRqsvpRAkgQ+WmF
cfLgJBgfDBbzO/8oe6wjNrt6zQct9NDEKKjhI0l1msLWxlm/o3YrmwMkk2/4cF36uusE6ROXhWVV
UExie2cNBi/yBuQtwMcq6FUE+fBAqkjyIuFRhRsmIV2qEgSufqhhGW1Ir+dsabztAaIJzF8d+G1Y
HyncN5oMTfLqQ8nIHL3laQ5eWzoQ5ks9yR1f8wXtxvhaEqCtnXIPJon/X01tkvhUKxLaVzT21Xv4
G1AILY6AJu9vx9RXTcvp8SflmRXjnbyGCOH1R7W2oR9Ows+nSsC3N5SfujqAb67QV7lH+n3UcaoV
+W9kNZG6VCjrI2DbC5C0LYcHeO1/gO/u4CMtExDM+j//xL1UYrZWs0PWQe87yqe9KoF5RqjnF78W
BTXL+4/SkM4iOT671emIq8kxjuqWN+SRP6rdSgtHp06KlUsnde0QOEwFwNMzoO0d5HIvLFGQazqR
lZCGjZbHj3ZEiNJvvauVA12AgquGvckEnIJ2Dmfq50G+H9MuisusQ/ZOrU/hj2fJOOfgKo9m7Leh
p5YBKYdci3uRlfNwyWAYUEZqlSLf0Gs/MwXqNHptwxVVg4TFGgABcfRGWVVU24tsGaDLl/lVRaKk
0DgnEn7neHlvn/b024cApawqXMj2/vHG0+xxSfvPDkwqQLbEtyTuOdHtwexNqpTUAokByr+2kPuC
IsgY80J/d064iSwP1pb3qaSixZPdDVUw105nZ6hCfc8rKSYfheG33ZmNBAbXB6yXYMT8loNpnY9U
SXTYjuIteEbLULFTWpnxo9QQphlC/BRcXA8lVtEM780s26HZ30RqV8gaCNjEtlr+8mFm5ns0ktH1
uk2WHJKm6c31dmbqGaeG3xBe/yn/78yL/TxxEpb0try/gOXqb67ClJfw9t1IkalzrBO90HNNqjCR
RYeMkK615uG7yvXxcp8KB0/cVe0jrhssYe/gB0CJ38qla/+msNytXc5c0wH1EvO7vblUODfzel4I
A63L81M+Nf+e8bcrjn7XZ13dlVa0fXRBpHETh03sgTcI+iSshuOdOgpYKHl2vemURmrz9EvNdwDh
p16TZqoNAQaZiMv6Fj5pUAbU02tt7u5wHePhZe82RKt8spzqiY34XGGT2jGAno4JNe4hBO9uefE7
X02wS+DoB1C/a+nvInV+cqtZ1gtIrkfRTlml4oF9XSRt0BH+J2wesjPS+M8xruAWIJQPBps4WzdX
xFkkZjUPAdKll0j5WDh45dOVlIrf1tdh7Ea77whJRkF7PTHtleP0pyRoRNfzP/1jdprVavLxfuRm
pF46PCnjt1VwzmOy4r+MGiG4DWYcSn9fgN50g/JSsp4B6wtuTASZtlrq4pgb9y6WjkIPp9f7efbi
J6fCZQBzcXYzA6YzVD2xEEQX+Ez4/rHpI7ERDSn1vXUbr5Jw27vIsjTFGv0Wfv6Ua5udn0Pl8TEw
v2AfEnwZsYcLDXZ7yG4PH4+L6txe8SzDSK+muyW2qdVxVXy4F7T8WSp3LWNEh9emIn+2gk73YOAZ
3CEy1FRPWZBRa1+kboxGmYgyHSnEt6jZLeB2lSzQ8Js57Bl4rrhxqIsut3ckrp7x2QPaw4dgQiVc
BzoqZbj0rmWMfI8eYXwrybxQX8Bedz7ECVe5VIDqF8SCDJAZdN77pDtrwitgIHzSruGqR262bZww
Qkt9/UAlcHAx6EDUwNInFdw9WkVm3u5zLB7pufRte1mLZGJI2v7xFFTjQICNuNLtQmrOjDGRM4w9
cmkrvgY4rVDq9jjevVkwgdSSa5CZUfP+cYkT+u6dt1+JZHXYPVetAgwt9UQ0QAKMhf0UkWSOd9FS
XxakqHmZ9D6548MiUJvzCzr1KfVp/4T42wg+kYZ2TRG5b3t5mjkpuDgT9objMg3KAxb1MNNzGVGB
Swyv5cBUHuRSf4rbFZJm4SYeIupvzsKQoeRJAr+7gZg7POoIbIAV30dyqdq6om51kYXdwpcJHnfh
zskgtPpvUFH6UmCijKSRHad60TK04KOZjbve+nlvV8Cbh/XFjZwpCnZLiSVCWsnttzGCp+hxRhUS
dF6kiQ/01bELbFFbZbWFM23gkTto0flEDbswExwaahsS0FWJ2HJ0AXln6YWxdFHsajEFOTU/mWKY
jq+VMIj2QlSzncBCm/lKFgijspFN2VQSDNJNQ2dzZBqN6OTMOKDr+6L1yd+9NL7cJIdDUexKf0cq
v7sj3bR9p7U5l1NdlecgOsNhitSe9VvVFPE6FN0YGjVtGgCsgSbzcTZT38EE/dOCvzdefo3C9NJ3
ykvefycWUVa9O3WpEEAcaaL5kiwhccbm8dhvcz+1Lt2ut4h8gv6CQg9HaNOrNVHDW/1zTWTYsPB1
5mgNAMKtlpGw8RWV2IhmY5QN1yo9nfIdDmyOmx9CrmNkUH/AXJNQUinRro6JELbEYGJx9YXlQJ8P
wocuLQQhnJEz44/hDxT1y6VdHBcFQptCNxDM6Ef+yyo8B04w1rCSfAbm2PsaQOyJffwqfFB42H4L
aU7ms95tyD01XTP9fUKv6DEp3YG6EEyoXZUkZq6GJnfM9nA5DV+BiUEXVSTHpk8GcX0x2Of8zdQc
UHcM27pPjQPxl7QFlwFbx+P1RwttnNwNjxWEeP4Qb2pS8fyojRWmPkFD1y7rYWUbfSUtGZ9iNTJl
9P/bHYujli6EVHDYqwVJM7UsKVD3IZl/a5vk5+acYs2RaOghXdhVlyrG3zwUnecJ2qDx6gOSXcnD
pqVRcXIdEVpFB6nvquAGW+zIHM1Ydm20WmIUzivt3bzvEr95G1igvpt4ZUgyFljM8AQ/q32qdj3x
l3Qx3pI4FYlmlacq6cmqS3CvWVwYCDtaSRJcr5rIufZCL87F1P8NMqYz9PyV1FgGsgbpW4LkvEQD
fzJjtVXyFqfmQ2Uhgfo2nQ1hoFZJeajitOZEHV8OTPB9tk30xg+mcmfPpOjdzcLKu0jgsTUSFBoM
tQ+Z8DiumXqPr8sY9evs4pz+PHZsv7v4FVycYArFgLd9ysJTi2d3RVFfY4zWLs70Y0YZVtNeNbx/
niUpom154Ckp9u0mXTTCpZpufbUg0dte6SiZYHWxVvZXTs9ueWhSNlPRvXpTLpw1Pxs+BFm7nsoI
KBev6WbgwpOAEHS3c4rxNZDIpRqiQYHGevzV/VJ8f1awxAGJY3hWP1HWNFNjGbogXq0P9PMavwGg
G409EwkP3RSb4PDraWEViduedBdiMeEGo2F4EAZxPPOFXigCEcHRvE2Sygr/BPVzg/YF4HOYka6F
TvsPM3RSZ9dyJTF7bH4/fpC+Fph3reO9T/8c3f6xp/UCXl2RiYKb39/CZnZLD++NUukw6dygX+Sr
E/Guw3gW8aW4/P0RK0w7n1sWvDmPyu7lnDIaXA6H9UG8KMkEv5eLkho6mNeq5kJqIgEGaxuqR2WW
VqhWGpnCizgk9pZWtevPDB3nkAbySQcD0FJIC2PMQS37gK4vRwdQXuAnd1r2eBio6suHr3PHi3v+
NB8OuFciaApI3+xJM6/PWXIO59G33HpGxg9I6dHBrZP/1LZ8wZyfbqry0hIo1jkq4EpTgnQWPi1E
aJgJ2w8Ptmcap+zEoh613Fkj/XznKE1YPkP0s4egoVH1Io9YWyiuZLcD3OzpACORrUqPY3aBTSwO
HbT9H6tJw8Ng/PNtfLY0yo1qhj/uWcWG7CKVMmzArouRhsLrDRChlf5NF/4ODcSo3/o1VjcmqVeS
jijWCBEqtGqvbZCgTdtUXnZTbDLAhEHtINNFUn0SjAvw7g4fyC5QcdEa5K601Y7IGHovq/Bt/CJS
8OTpJjXme5dID4DBpmFap5XXOjaRXgiWFBQhk/KGk2adKUqaZPLZD19FOmBFXT0yqUSN5ecA7k4t
xEuPkhLXN/eh2pEeVoulqA686BA0fweIqlZpIzJ9k9m6hBaSs5apxccCVUVUy4W8InLAbtu4zgFm
q+YAYHmm6tmHJXvGtYtVGwmX8PXsOW/+4y1wTzWOhfMKjl/Qg5mPGNpVuYVIm5Mm0tw82YujwUGW
x+5Svn9P3COwvZnjXvqF0p5JuZS98LY3N/Z7hAS4vJFb5+ovoGwnz9ClU0QUeeZs9mAOEAksJPO6
26eQixKmX3NaeQjYYj4n5qU66qYa+avLQjewQaTY5HYCb2yAruyF8OC2FH+cXWbAlRv7WAv//MiC
b0qVwqN8cfjiwKhA3pb8oMctHs2gy6RhkhLWT5fuU1osQPQHBc1rCrOustgG8jWfet3NVaRF0TWI
munhVGDX52fiuVI2PKta3qPYX/eV6Xwfnanc8k1NW32E/QDJ+qGlAXY2dML9aArAH/Bi0TUat+Oa
SLMvFAHXXUPnt8C1mjsBBsZ/h1bNt7uATfoog93Ce5IaVWD9Xt/AWXZlZCasLoaNAHIJ4LdB94+2
k2RqsBTbktNtAQITvG7pNOEgTvETi8KMR3favHVJs9/RVBvKBLIqyxLsGSOJbfVYgWyaznZEShg+
oAJKS5a6f+VsoPDCRrL4Wp3orb/Teob+p+i+kfB/CGHJfhDxT2ZP33rTWJFE3MxuxduXH2uj57Uy
8CX9GcdtEmw4fsR4lzPshczcTLT5+rxCp4rcVL3T6k3q5ZvUeqdTMtjQo/ZSPsMyL7UZoTLhi4TB
TfFRuhvuhLQZUm2yO8AK48s4ujK7BFP/QwjADE1ui2YC1hu3jWhkDW6ayMK9y0FzptaQQRY1kyfE
BWu+SlYaKObi0Xx9VdZ4t7l39/vQ832oTvbjwBCJmncBap6Xb02D3JjkOHyuN1PeJaTYtZ+Mi7tu
KgpHBcBHeFHc2mJGDZjbmx25gNzbUkBaTrRIF8aIwQHUFM06Kwh4gSThBH00AdGKXrdYRGxV+ujx
aZsIpZg3FjB2BoLDAw103NOTy/OtgIp8HXc5YOJeV0Yc7zdEoNl1mq8MM6vJGVY4whNWg9PXGu0G
pOGNVaaM7o1tYy/JnB6G9NHEQ+73Te0NK49QF004dxRo2SFa+oxgUkhxVCCqSBdmBb/a59q9HZJZ
kAPI6c2QxDZuaLLYCGPC5NAAkoIwHETXTmSTvKNOH6bvPyluM+GrGCwTQKTN+z+lpATPNcDDwizp
rFuJL5RSsFZjLWaN+MU3mWEHncjA/FnZbJE6lePsx1Jrb5FgzOiBm+CjAJ65XTBHu3vI3ypNap4O
/fCHTJdHbwpI8RDMCj3C19WOHREP0U4ppqRFkt/w4TfQiyt5b1/P2l3PLBzcYjfoGoq4R1YK2XRk
afYhga5uHdWFhFIAW3QMexuaErIWXphhk3UJMHT7USKtn7WTBKFlfvTirtevpaEvW/OXyQho18m+
mGh7+1t32OvzFqNc+lTDcMHQgJFP/yxSeeRzFl+VXy8HMSKE9fpSFHbGXw38JVTsFeVHWCoHg44b
e/iayhJURd6owwh63/0fKlrIDMDo7BZp7payMeufFhZFA8FxZsDKXB5aRq7gIw84ivInIv6vkcm4
qalN8KgBS0aFCcwuATWgJ00lbYI9yqA2u9han2h7REsaTHzsVdQ5xZ3OXceGwRk+iCMtuHKkk3oY
3wQrJdjLwH27gQLT7ybfmYg1BNBJagExnK7x2ZbwQzFB7XETT65y4p05ek4nsoIyPJHfYztOyK3e
pvm2nRja5uNdgNm5qFepPCBjW3KcyJtdoDJ15/DmcFuTE300y7dKVimVif56wrLdLN3ZNgxLcBNC
QT8qON7mr1XJaSTtxYGbbTQZlMhsxD1G3CMypQCcAYJ1TdAJ44Q6de+gcD047hiiWldt684kDQBM
0yganXJPeWVbmIE/sJQizDJTKn0RE4tJyks8KMST0Vx+8SAvRnmp6TM8XhiVA6uIlxGDCIpXnXDb
/j43kt/SH7sXOBNoMleinMt3A1GEv6HqfGIHbjpS+AC6SMrWrqT9s9bn6OLuecYoCd44UZywnkMa
Te0wOgMJUunBJYydF15YSv6sgng+Ec0WQPN/OF4wfvXTVckpLQjZawIACdJnk0alkqiEsDsYZC9Q
15oJ9vpe8xiKA7ugTB1L00uQNJffQVuu0rbuvWgKjVkkA3SWCDxd9pOwIuSeNlmMAQTJIXlrosIA
o6qQSTevDiMb6Z+fBir75ipYins/CuH8Wig1sCUja9XtceGm80lSU6VO5hReMNOqoT/8Tt+eBKMM
QLwfUt99cPpR59Qsg1aYNLsg/4P60UZzeoacSR3ZjEtY+JzWJxoysMIBh9o/Kkdkm1vw3qTtpnbS
jbmOJwVLhArDqs1Lt897ydq4dFfOftEUYKFPkgcvwPDu2XA1chtglMGcfuJ3MyWSQ8Y0wv2dRqyR
1TFOEcjo/NS2GkaNaQgxK1p5JDxlMf2JLonP0/QH3rL2NeGVW89VUEJYki5q8OJ1s0gOnog8Pjcy
3v7HE4ZinnHm8AiWM5AsEh6JwlPxC1CP/FekASxQ43Uu0jI0aXimKBn3cXAXk8q3iRVCB7/6AX5p
KFh7IeOo47o6UvUV0w3X7rZKEj4EJ/22SNVo9uVh90/yYfxw21Zf28jYz7EQTSLgxPOafVRyiWZY
VyDtEZxAdq/hA8LU6elAjH2sm/7ukoMjzV0YiNiJPtmGRttmFN8xpVi++cVhD22+cp9zUmZ8TOiR
F3uuPK8bBg9Uh2+SHdaxFsJ3x9AuMq5rw4GE0N/LEY4wCT6vFlDCPPqYb+lD5YJn+NkQxV6mM+Vk
FwUhN5zg9FSEMEgfN+/q2dtNWt1T6l2ZOVauO/17H6bqK5RNAKobhPmPly7dyoiAlIzB+SRaZbQT
H39LKDryLfZ0Q1pncF0EBBasXVtA7w3PNazTCcdNRwUfTLGQOhAtBMMBRFd7HfNectve7wUsX0Cu
qpI9heB0fw9c7DswWV+2NKqx/NdZvFRZnazOWUZR6/CXg+8SHXAwbWE8th36jfZrJmUV1YZY8jPL
Q73xQ2hzQ0LBlfLA1iSrRJmiF2GPApaZ2Yl49sIZ6F44kSGqRyocuncVSfo8gmjGAh03evQW+zam
feuFBUWoXZc87EwAlJzXmwXQW4rwxsZaFgdVt9Yb9rnq4AASS0+LPp5RnuZZIfZLwSOceGnYPXQk
C4M9Vf4SgNhkZJHmITs9MXZNoFo7APpZEdGoCgcEB0EcRGI8G3pLq85FI41P0JW5fuNyL68J6YXJ
OioiG1xJiftevBcHjIXJ+5z0KOwzWajJfr4/6DZFxxeMa9TVLxlp2viifc69ihBWEkd9akzeu9jn
WM68fprryR/1yinRd3U+pQiKq/VTsM7MUX8vy823ro5Zu/FEEqwz8ZZ9z0Pac8KQ2e7fRqQoEHfk
62b065FuwNVVkSO/B2LvQu6VbwvVKOFLgdN6djBmZOZ1nSvuHH99QjFxw/Zhghaz7k2PIJrYQHj2
B+wZvxzxMcAp+pQcPEwtM8SgUZIJhKf6d5F9sReMMDdDuWxtg8Pq1ikOD7mu7NTTn6AbLjktM5r0
GnY7Jm+pCfhQLWmSXyyxuChXPUGoJdSUnHJYlVu+9eb2m/cNZQh+f7boVst1SzKFxHYVAOiYrZQU
OJwKgkmLenjt0wBJsFFP87lcnqOkLfeg5P8id8i5XyDL69/imuQAvDuG03mncSY6l/NdtJrNBQYa
g8bvE58u0Xv2OgIly2FyqoQXzOpmH+xIEQvve399Ajv6DRRavMDLvlLsqHkV0V0x3fTUzCOa3YQB
jdtDDZr8Z8Sxw7WocQIqRGa4xjXWAJG7vF2CCFUWIwHszKVZntCX0yFVIIg4ojRogZnTBH79woCd
YUtulQKyxrsoEkEMraKX/fQ6gZyRHj5QcGa06TrsbfZsoBDqX5nciyDIbOLCaa3T8k7HioF9AbM4
gBTnmQSETnhFzDasUklrGe+RDv3BFD821eVde1tGHgxIFZwLyBsnUd5RMsq9k5jExyuEvY6LCGfB
nSuuoBqcqPvQFAOV82IHb++mkcsBAe7fJ4X2gT3ddPOgZMcPp1gEMNmgCQ1fVbcxkt3q5IixpzAL
zIJEE/UBw5VFhCQmbWThSmOdNzE8VDghdC9V+Vqq+wQPw4fQW8RRsHar0fH9ag08bIvxQPBJ2MOI
hlYifWRDtJT0zG+qztWm66M/brfn3R2rVSL1FBxV5xs5ScoDPNCNQtF0peCpLitjwIPrQrLsG3ca
jhfLv+aslLXTUi+4fKL+5ThNpzXiaG4o+jy3+JUZ2+IUxBuLXMNKHJqAddRDNVgcp/CCbOZXzHjj
kU9vqfVfeU/HbT6R4MP09HvAHwnGox+OdISDk6acpiABh/X2GwB7A9FxNHt4GvI6N/txeANOXuEB
AswK3DS9Wu7eHmounHd6HYa+reQvE+hUo6IoHTCJOd+08CtioQX0PoXbHhqiMW1g//djyjVutMQq
No/UE1eppwzg8prlhBT4R61+2wtYIO/PuYX0kjgJrrREjrP6TW4YSsFI1+kvoXYzyjLXTnCpyMkW
F6C+5JQm2coPAAI3By9mbu8C3J1nFDHfLr8UuM9rZoiIHCZtAgIsj32Qci77734UfoUJBj6Jie3A
QLte9s1GLTEYx9+tum+JZ9WJWTTYCtNi9oBaN3xSzTJ5HTyrKQ7ON4EvA8/4jSY9LUciSbMVZw3N
FkCvfaTL7CmQLLEb7DeO+AcoLZ1TWyv+vWqgNI/83G1PWTTfXyH2RK+HO9mwv4XmoC9chEYXCO8H
sq9jNKR9KZvHhLnYJonV7AP5TJUuMTH1jo75YSOGj+rzbUeBDl8s+5/uzJhpM16viNjMgmcuRu26
oW8ifCy2KSOO0T6gDoUCf+krq33qWctW+x3/q3DD5zLCJ0KR+PUza3dvblfxoSKz/2xmP9/IlPz7
cvwy5lgiMT58Fg2l1ZWekNOTsIeCqTuzLMcdslI8j8JSXY9VFyeRgKxI7S94ZfGp+EMe3ZqLskNW
u1D511ol3zJ//9PqoZ9D1l7MxhgEuqA0KSjXAPG0JQxCIY3cfU41n4ARwoFdATkwNv23wLICULaK
AUJyFQ2wtApHraE+tMyti1HlKXbxbmL7vpGycGSDOuGbwJWDe6yV9PoKgtu8JIbXdTWiYEizXIo9
VOS1FXEpdiv/tqwr/sR+7ME/Fyj90+D37jQlLabWzQGkTDCVzi7v9bAUJQcJki35kY6rLU3jEa5k
PeaP9dGeuUQ+owf5wcNgADC3bXOw/V9LCnOilaqlBr9A//riw6iSjCBe+JGXKE6yVUoliQhM8OBf
odFXvYX3h1PCJabtCSCqwE97HQWATHTLLYZIUqqqYgpQBZse6z8MOLAoYZLlKbi7b19xx7BE7vbd
MOdkI/PP8LJoEkQbddICIAJegbErEXI1DSiQBmJLsfxc/vJpviCsMxUhErrpvb+jhsg4/3XIIA/h
mruEx16Na8PA+O9/Ia92HvtWJXCDCH/V62HJpH53b+mrYXOs05uj3yY7j32otcUJrfsbkU+3iFd6
LsJpFuRwp02j9I1YBIao9bZFITHA3zPSTaCqgHq5vUXkCwgopgQjrSlwr5B+Fiy8uGe+X9OqCBZv
qNkBIc75Nzom/C+51EtSRSwpTdO/7Og/s0V8+p8v4jhTDchV+NLvpafPTZk2/3/YFkiNkq6GHvkC
jGZ/sop9pb6G4mY5hSLSKmp32yCCuKIE4/9avttjzcQwnXdsrDfPYdAsy03DjHZQBsI04cvgyi4P
/GmvQ9/i590/xkiAo9pe+Rda7CbfXTBAj53HtWm1rfENr3/47HLNKyV8s+dSUVJ0oKxKnN/Nrpgb
RyS4eQ9vJ2gfFT7vHfCJ8sPCy0JkXAp2V2vvJ1ZSYTH77d0ga6rHVTtEIWmgST9+ALKY+6JLmO6G
EQMFUaFKLzdgooV5uHnWuFnwNxDNpm8gH9N/Wv5qPfzvP1paliIhbErFPk+0tOWntMKanQoa6Yhn
j+jiNVg2NvuhLzvLWQRoRHG7zrgPoYE7u0mA8YcNSZCdnDiwWWj9RC1LuPN87IvIgacnhkyI0B+Y
6V8Fg4lIndGwa87vFTSltPgwcrk33Vh35JXsGLSjzKsPu8woXv3EMcXibg4DDjFNGT6xC6f+K7MN
Mlx8lnUlkw4ciKHxrZI1DIY1RFzpkMFVseahp5oCl3xKK8vLYVkf4R93bl1H1t10TdvykUKuNRJ9
qeZvJnT1H7H7Mfwz1jHHc2QPLxNqQ1xiGjsN5+eaQ8HEdo+asyiRYgbIff8f385/gQKR9G95JUex
mRnGRwfZjT3BEYWZ+8UeuD1fpHZRPuvP+bop/B7Mj7MBYiu9pdwKY1eFXGD2i2+qkAaMKVSiSzpg
mnfjd2snGpNQP+WmdbEFCr7YL3knqgE7RQlAMOpE6m1za8DdZVf9w2G6LaEouHNrA5ZgI2bzeznJ
7fPabHDikSkMkIO2RyJzzZx8bZe+0YmVqb0qL1qn8sl1u6vAXl/98TcEj2v5vnQ3nU5UEUCr7SUu
+wdqeVRclNLkzWM4asXbZkIarhAexTRsvwZoS3KXWZEjJERBbuad4F2Bah2WoUUGxJyEgFWXEk6k
kbAc9lL148iMrNs/E0pCEDme89dYuQll0301ZYMIOyjhwa7Jq4klYBZX0PlIyzsdo59m5WDq3JsF
yddsoVFgvfuMZ5oNe3/taY6wfbgMjHQCzSCTqnyODe7b7YHjHY8bXebuhTGLSoE37dWY2F0UZY9V
hiJ3mgJIEk0UGbw9+yD9aEVkuZkaKmbDdmOEXuIknlBpCq4il2q3QV0KPajDouU2x2SqoGf9z5Cl
C/ZeLWsKYVfTuSsYZJyAmPbrVx0vhXuaexjv0fWOXpeUZWrZQvnh3JPg/KIC5jqb48rEDZnV6Wwp
v8lOQZQbPRH/wnJw6mG8okgQa6xTQ0Y6nT2GpcDQEgmUhm5DO19sWwklkk+k/AW3iTCQWszAt7Sc
B13gy8hah7yFdHvIQ8ztJKyPSTh0v85hot1olA+wrmhE3T+doiHQV9ArlQDZBKDrsyaDum1mHtOh
2FYbrCma5MLso59Xpwpm+9NUE25JFPizIuM2C5gdFacc5RJnv62hdAIbVT+VQDfMxNSl7NRyONJP
hi4R8Uu0aKbGmb+rLnsmj00kl0/PMP71iA32puEiAoi5UPasNqwPzZaqwaZ+ByVEzWyNk+Mq/PqG
d5+vK3s7bBudOSUsJE39Cs1CsHztV3WeIj9kStmb+xqliEGV8+jKd+zNijXcRMQJjEHsr3knUW/3
HyxCA4I3LVYqLfI15ra0b87uU0c2/m3A94/2MsoJqd/G82C694vIydiO34teOm0+l9gPiXSIjrym
YelL3mafX0k3cmuGvM5vIxRTrhCRshif8O1AE9x2n1vGP6Vr5LtSczF7HJVag8ajFmtYVbtrk0ZQ
xNVnNsqatPSjZsa5O1uCXdNo61NzCQHIES2Wa+h/JitnJ7CAofAhzf4HfE5OxEB4E17aiUsxWo//
uMLvt1HgZ9kBWI+HX6q0zemNOtHQ6kVeSTbjVbKBzk9/Fw1tZZ99nPxCkqzzPckHkYmWALfBtC5j
HR74SjpbFqGhEno7EecgP6XFozpEXmfURZMKoshFGWFI6OXfM4vMjXcsKYO3ykMYNAaX4AlS2hPQ
eFFaOhX5j+4Ml8bhlNgOaJh1bTRLMO4msbtwVZV/fi0cjx+6ADX8Bhh1P57P/chWQrbLYgWs6sgS
6XspPnhl3b1VLxZ8n9lN51c5+/13eSEPAzXFnUoIbTbYUXeeVS5yFA+UQUtmf7imd6wQVXPDd321
dH67Gj9m/MMqsnFNLF4B44rH/Axyr6G5rjl4XfygRILJ47u3zpmWC6FlqnwyWdXi7hZdtTpbWHBQ
M/dX8QPlbuOkaAdAOp0YToaG5djnmHNYjSzKEgTRKUKEmnWu0ZtPyoBS4jtS/CVDW8a9G77+0zsi
rmIZKHxxg3tdBCnWeW0EkQCdZzy6lbtuXlmS/BmWtZVymyxoCAZ4/XbXixzQeNyjxINhXnUu70mt
TdKIr768jNCnuWk1drb5SDEKUmuX+ZtGKeTPvUZhfo9Yb9O3fpgBtmIvb0c0C6x/x/oagfGCYFV4
pb255+zev1dhJihBGNVejFmSbw1hJkKl1I1Q4qQASm2lBGiHsiq3vCDzBdLFhWrzB8mKVkkxrGc5
mePzkklQGmfQVjLIUc93zAhTSdZ+/zgfm7xDdMFVWVy1fONCSFMhBTioHamSLhcrDwmIemw5DZBU
4WbW/2epmeV2+osVRqgnxBxy2EGEa7WcyGYivleVlVO1gQc3HClPZ4ObOCtfAFKefSYc78nisU46
04JfeVD0ESlQqwSWIqUkYfsCTrTznSSG4WJm6xReMMAP4FFLWTVTRdOJwO7DRoTvH6eBS6Tl658b
+1L0h3207cNV8jnOz8Hy1HYDZpxzr677+htHf9vFbXNafC0tCoEiKfe12d3CW6QUBctJAKTuyzXj
CQPxrp7SzQDpTIjdza0jsT1Kuf+WLYfMUJsZq3nixaTCFDLVuL+ekZLEnQOYc+zFicJY8eqB6yxy
S8gVYb6EcIHHLIj7/vj4o+rtmyEtDdPcr21/JYcrUOLBIxYGzhVecMUB6hbca1AexhOHFBgqyc0H
cZtKED0wDAetgOGdCvlOVezdb3nFV32j0VCB2ArQR3l98u1qblWxR1HqIpHBb6n2Kvy3iP/xfFi2
g4uCsZhW4pUwGMSI43ys9rrsh5NWzp7D26ptGZVP9vSYkqTCPIA8hCzqKk2qPtLjslEKXd1/UzMI
LbfjBby0C+ScE+V9PmYm6AS4uvXmDwnSLrLjvkNXfT1pPeER0YiR+HfrZh+n1imlLeYNaQx4nKJT
eg4n4NBGN0yfl+73JYmf+s8NpOS3c/sVkQUGguN7xuuiVBu55zuXKydxjFAK9M8jvtoO99yK3Bgu
SvtBKffWhcTmQW3f6HcARQBHslWZcx4BgaMxql9gHU3vrsxuW614aNz3I0yyPfyK1mtJRcN/1ZlG
vgI0JEzLngbXc7avym1yeixmtfDX1Pvc4HBnr2JFbcuXl7VWoc5izxiEVoGbV+zI1brNtcA2gBl4
gTuWGlt0oyA3FcwYTfH4wFSi69O7Ri+NbWkueucpLy26MEV/9kf44QMqYXl/c/DD+dCNp57E+a22
IqYymBNPg4C9N971ilLGVchaugbAeLROYCL2HBPxs91XaynTg5OX6L392C9DRjDCsM/EnIxSH82t
ANclHyhd/n1GDy0FoLE7/hh6cdRAOFY+zN31HrlEbmWj6+Z7HpuEW/VJHm/GCDXltFnZQg3mqyCB
7iXKKzPKIpYk+Th4VvqoiqR0ZnJ91YkBbosypOWsQ51QJt7U5RzMAyQkEkkORjwDEhJLmvQNEBX6
ftGp+CJ/3WF+nJZgtRj5k0IesKRUdHXZTeFxPwJBzKK6/wndvsIhgF4+bUOq/EGh7mo769kiR71D
cO9crbV+icMfgmhpyX5SWXfRiBSezzzPhcLkXaDaPAdWx1R6IKZJ61XWlIyakJWr3QnCFgMq6S0k
1a+HzWkezYNel51ZLlYPps3Tdyeb7NJrdjoFB/mIa/2+ZH/FP24L2qOPKuOfGrMtIcAvXNIOEk15
uCIgVppMxGt2nCy8fmZ8g5nfsA2qIqSdJkT0NdQOU2wvhzvX156bAksyBECvPxTPkqMLXDy8z9Ka
Gvp4b2qVN6yTuW2fJsqEyx93+ZEwN8XGOxAtsxYjCQCgBrig1vCXuMBOW2M+cY2D3ivbzhGIjLhs
Lvy5i4+XflsCHBQK9Rmzg8ddU1iV9gPyJdZi2e+bSRjt2HT4YV96dBUHpAhRjItYm9cXgyn3tEvE
hRX+iG8OYoQ2bLErmhL9pTpU5tf9bWe0jsjCQHRiCVLMP1kk+/svzk97hnl65AzjKoL9DVzWLktY
O2ON5poSMN5fCs/KMaxNsOf4kjcTMXZTgolTHZa5fS4xdJOvAryMqwKQt1dZOcZkR0utRZb28O/9
e4x0gIhlxBDa8QoepCti7utmHRHY74FAoCuHAbfNDk1tEwt/b32KuMaRnymnPgKQpVttZ+6aWzq6
e17+ZuLdMywAQkotMzT4L3Svtp3UXMAVTHY0r/a44he3ebi99niaVcKgvKRTiAS5QY6r/VupyptC
jzzmCh24vbTfE1VlzNdseTaNfl4I1BeMrbxqc1+vCpi3H9F2wy7/SMQ8QYa9mDfT7HIFf50CsB2z
IucbQyykAMgv8un2VNetPZdKdU45i/WXnFvzjE6ElTfYAt2II72akIZ4JaggNrb88VjWftH2rlEp
oQ3CwXAMbNfYzCjAB+bZHLCte+zM7o28iyRzKWH90V+kzeOvK00NSbFnWPRHLYFYw+Zj5OcLHJ80
svMvsUbIVfJcuJJN9DaFNtmQibOIhQsjnBKP+6o8d0o76Cl0yDeg3rDS+hl+59jtvLiU6VICZRle
gIBWqaDiHt0b9XopSz/I9C8OVb1zdWFIMAnxkkztVorldQQxqD2PMESCI1yuyLD9iRJX/tlyKfAG
Z55JFAwQAGPMZT9wmJ6JJawWX76Pl6xW0sxlXUXK5eojFrWmDFIMyoTiEnm8IyLf/PobmCx+W3Qm
aI4C91GgwAiniNbHhhey0S5m+B0hub9ZgcsHwoH9N6Qok7QznnZQuD1d8FCNQyjjUnVoWmalrk7F
eu67hvIAIhJy/Akwy0wOaBkxdoIG58+gYVfPImVmfFPaYVriWeYMN/bz8QB9TX2d5LOftdbyDdLF
A0Xl9iTNTNi92XamWc6C5j+185onuEWwsB7TmNoWdERjfnwDqgnbax8GTuH8nGGok/pKSGLSJVaK
S/v1AbdXeJNcYS9pxlHtlunROgtjPE2m7NrzE7Uc53RhmLctM2oD+gyRAbnGmBFo1P8jkAIsam3q
U1hswgbkNcBJbCqZP+Co11fW9Cdx2yd8QwfyVjOQLIFEJeWGhWZuIZ6e2UJZenU8ayqKf9NMnJ1Z
xL3hCUuCdogRMmBHiA5zvN8BrzSvQ04KWrFOeDeZPyT3gNnTHE7a2vwIk6RvN5qi4akQ+42K+4xQ
uNgGOUnMxuoaD9kK4fVmJXjE8a5NXCPkhyFvbF4L1mXygZqMooHwm5/ZCDWQVk455qhnqdglaXVV
m+PdoiMqRJ9+Zv7m/rthc9veBGOoPeVgD/mPaqV6vBjGOqW7UN3a55OZnl/f8ALRj6RJNab/er4T
DhI5DYoNTjv1rYekjoWP4TBAxi1eLBQhpqXvYnUOIIEzF5R2JLIy+xH7K77PUyOu0LfEiDXP2f4s
HiOMFU/q5YWoAdEPRaloHQWvj3YNHqDJZfVOIZomVDqrwQSU3oRuL3K7sTDn+DdHLwhMj+ZUaCCy
hO8UlYT/bqRqLThM/HUAXngcGRK95klTC9kRmjcwxjbuzGNOs5I3cTaHOodlegDpsMdka9FRHN1a
EvBxKG6AC7hT8MCQEuyQ9uAGc6/ohgnaTCcuTiTfLmF282C+oq5MeSpCi/2f1tZJ506a9H6CN4Nf
KdGgwM+btSzFbgC1Q6lQo8z/kI1on2cq9ThTrF2LfeAB+Ay9GCEqEGSZlsGV9537o5nsVpnLA0J4
kEjjb5lFv4a7KOzenPsGqmJ7axOdM8jLxne4ZfMGz04MQBjwSF609v3UsrYES2LVpcEb0xA6qqQR
dL0vGLDXPZCQuZapUVJMlG2nx9d1q0r32+plgGKMLYbxdsVfwsVEtki9/NMXwH4hMifru9pToi5i
qLSM9QYBmZWzYksRcdGt1KBKjddeB++l2DISDOFYljXjTWfuGuqskPiuVqpAhF8Ih3sgs+T9NkTs
d8eKTw4DZXKaVD1/xkC/XV9pkTMVOdNmdBdCKTqDtGn14O7YIQt6i7tjmr90cAH7SpU7IgTS1TZt
bDcvvU7x+gw0nVFGXPVpxXhAbSsuV5+ccqd823OXictJGkRzSNIhmSe30rblOyFsB9Gbs7ODPT9c
yIf/7Gpf6qJurYtQ2n/mPMbw+qZERhP90u1/AGENAAFAjDitcY+3aytkJD1NOUubQcDHpnvU5/Kk
HL7XshezLEyDigx4SzZpkwIaJoTQrx65MGiOkR0sup8Ls7cUTC6w4RH1AZNNAtj8UbvXcHdxJ3Kj
JNGtW33W9lazTtpFUgTJeY/RrYbyQvkOdJEg52vkbo/K6sZxd2irTT/Vg6pOtfRKPHwBVSh9MrSa
7++12gz9+a/FCbuKUzIvszmzI739E8MFmwFerSbMnmb9hKbBDE5Ml5MU6Oo09Rpj4peRmhvqtHy5
6QZG41dgNn/wAyd72CpMMPKb8f/r5/yDQO3/myUCtkUfyJ3MnHSGre7mMrckKu+tsybZjXwxn+Rp
OKJmOWQAwDqFIohphn0gf++f3xfbWenL6LEo7KKp8BlVvr1e0feJko+gGROKChEsXlWJ1Gk3NzMj
sz/xetTrpDLn7R36i0NVIpC+wiLEAFp+9K0adGncfysjJKTqFIL/k8R3g6XJXFqidttJ9XFm6ioq
fF9V7M+c1bw4aBChhmhUmPbtJQ0v7EiPxzLmrqaZ/T965LZsEKhKO/1gX2f82wu/3D+p5gu3VHd2
NLJGRr5C1xRsBry433cEcjhSPJTfupBuGVpMuTQlgtsB+eOnipz2siMRzQIqLWqBw+/Ik3DotBRn
ybqUj3XFJGuwIluJSvrPYktQN2cirEug65eMtAYw0wVroSQ+AiQoPi5g4gkhGqC67g09BDAwxINW
QcB8iSa/FfN24MVjbx6rTQ/eh0DpS4MZ5lXesnj7OXIE9fYBQjzrfi0wNpNuW9sqhiuKXwYPDIkA
3gvhThr164+C2WI2lXEqtGVxBkFxTp8tP57f1YauNwntWiKNnpO+0re9O+gLx6XkzY6qDSNC14gy
yATTFw8VwKZTVg9rHHEnEvlm6+2ClawIBNgsSIwolEv2SFp8o7cEWKk8z+Ed8kclf1lA4XdsOYwK
A5PAvYxZbx52VMrPVRDo49jsw9iMJku6vLjmNwAiSt1V0xs8pAmpCtQjjm+wZ0LvmDhcgMFTZoUh
Kq3TO5niym50zYpv0ekwnaVNFuJNjruU4GFRt2rCmBuHz62Y38lwAObs2OW6p0Oz0RkGofq+99eF
L03FG9MT8TvEBfh7vVxQQzGEFAXSq8mGL+HoZ3eDMjfR0mMeGh9Q6W2SWs3HYHYa54Q1x9/r+6iW
jeslrnPZQiuNfLgQieUNsOwf6c31jRlE4Gthh270csWaRmivoLImn/XAdBrWyM69wA5nGROUc/lK
QSEm29wAeeWkZAulwec78P4H5akwuTucC3/ohr4iGhTEQSgYm4sT5hwCDsFwhw7ExSQowuCdaNdl
73fIb1mR6YiXCM8VTqs6c+1r2xwNgmR93OAEF2o/ZI2OfmnsWtuIv4z9Mz06UJ0VksaejBRqS/in
SwKkLFr3a1njrjhlaLaOOCZs0iZ+MgL5iljMZDU7n2PVXGfzFWkyVv67Lw9OskUsRVHXiBo6E7S0
RHlXEMeOWLTjh1tpqoqydGocU4+KvyNkwZ5s89P+z47AzkLu9+HPQmM2gb0x8KvXN4wLMSAGNpSV
0xdITEVERJQERNiprx4KIEa4NpxTKuTXXZdgtuyChg/ZZzYnlUeVeY3wxVHUyMxMXQMVJwLUwqBm
kXVHdOBQP5/d5YAwvQtkKkYJIBMVr3iTl5mcfhOvHA0o1ItFhdiNimq6x0bYLZez3HpXVVcCOMVG
rxCrZdVk97tVAxAKS159StHTVpdBai8RYxKduKMxp0BhIhxcePsoq3Vlzg4jTauomPJmBcuq09mq
w+HoYuW7Q/59yDJca76Fez8qOBKN6KBZA2h8hkQwHuSIAwA2KvD2fr9/iHxnAMySAN5ZmRIZkM2T
UDe9txATxtBcZCcrXkdJcTWzCYROiM++jv7qdJKP/MJoQ5H/z/+DIjQYVND7BiynsUbYQI9oV4Co
7gwk0L1AvwUKAtSvbLo57YUFchD280CMERbfo3MS23Y8/DHt8cWrtXtMrtCNVkofNGH8lPNYR/0q
A18TxjhP06GXrsNnrR3aLzHPv8xpQIa+A6a7+3HRy03UCF2JFvde2YRIWFd7CZ4w93sU5XPmbNlk
WoKEjPwKPKXNQSwr3mRYm1j6WHiC5cJ2W8XI0T7nK5045A5Ym2rT1nUg9zWuqqHSSdelXuRS5asI
iQPEd5Xo0vvVI3v/Vm+VczvjJEgRIOq4G8zcdcm+/7o36uJp7i+fDGXgaGkUSV0sDmHh+UiBjKYx
OFIizhTeNEiUWO2Ap9EMQ3vB7YS5xIA8r8lcMgAIc+z3jwoIWqRh8MkKGYCENzA3t7Ira2h97Nau
wT7nXWFr77K8dQc2Vm0wVe3oiOz5vr+PiHKFPQnuDmUjcLHgwVvCoo0Ts4IJmf85zwMzlC9G8wRO
3jdMr4UWio/0935XsAqu+pRLVqtsOsWki2YMD3ghOvpnS2q0YQEtBISFf5RhUoWg3lJm8b4LA31V
LXgMezTsnSO4jhkuoIOmXqZgbGMpmeHaZU+tiT23hB807rx0cXX8i9ZTsGLmD+7pvDTI8xphBzX0
LOIK7nuX6hDlDAs3gzhlm3A2YuTfThF4x4KkDv+aMdhA/ektaex9Qlutt7+TyNi4e3iPrc9Skuy8
RZiKHCQMa0x4WTPUWWHgioZecO1eRoGu3qOgxmSN5PxmWIicL18EF2LR0LCYnfCTUJ4HJskb6gQ8
uUr7lJ7jJhX6FZuqH1ymvGiWUBjoVacJ63PGyPZlgv5NfpgePKYOkLSeLEcVwaaLwExehPLwqJvt
0HFWZ2RQeY9sJVIsVQN79q+JPzNSFAxMlHpFCAfepy+aWMvrUDqkAtS409FZibIJABGnIjhw6II1
Kjtyn/Y1hADkqlBigyuuE/NlYDwEc/U1AdvOE6A49sTIv4WC2cOc9qM5ShAkhm4C2ZS86691u7rJ
2XWQa1JTGjrko7dkM7lQAf9mgUQly5NyN0A8ftAW23Mn8cA/sm3ohuyYulfVrbetUBSZ2ZTFzvFo
0CoHRMmqXMenHQP8vbHvNWifwzra0855HN4arwukL2DXP3ITGHr3SxrU1kUocZ6DglBRXvKIP08Y
DvXOQkpR1AdykcSVhU8dEMx8PqlXbPY+7Ur72h0yYJGDaaWuEjV6Ej2zSjIb9r4CtyTca8Wgp2G4
Vl4Rq/xQe+WemPZLRPklfhIdeTC8cwsekmmQcRH1B16usQlX/dP5Fn5j+feW+Nzz8w2brD54K5nT
LstZKPOloBniE0gvKN48YgdeNbeQtsHt03ewZZqpAlEg/qbHapruuSKcfT334HvRMxL+GxYU82JR
NbKlq2wyrrNQOYCjh+6hvlrITTklrq2oKLKpMSVKUBpueuyFVRlkR2A3tQgm5OHRYmea2nlT/H4p
MMo6ZmlF4tnd1V7riy8KAy0iCd05/+hmhWrlVZDOZQJyWFm4VLwpLF58EL0XP6/Q3F4WWN6nAUqo
wgHNw0tSQfJeIn6KTBm5y3rqq4PL64hcMiYd8MQa2PcbDrr0Gw9zX0ciCRODjvmeG4Y+zx1uM2M1
S85iYl3wm5uC/pp8rn8yN0Ie0vibw3VuQDB+UULm34JDGEdF9MrjifQD+vQJXMoX3FVCUPE2FEEi
8mEVHeebg70o3mzjctWTTj/Y8IlV9ZAN09A/4a7TDF+1dE/JeKgoiDm5C7eTFsT4VAMkt1h0v97/
CPRJRPjYH9y8bVySZ/N3rpe3hlrPSRE+Do0x+oRmNbVkiABXM664DxFmnC2erfQ/lT8tI/Ms+QQp
Z34em2AtnNGfUG6kK6Mq/qB+wj1kqkfdDxnhW78XpO6r7qZLIGpjIdxrdJ5aq+kjpzj8A5ADOful
c+Xt0mMbdjL+BHN1RQ93wY8b/OLVviUb0IVjCFJ2aGLB0mP+YrWTHclFaHUr64l8iSy0lDVcMwhl
eGfNXQfZLj8931/veY35A2BtiMWeuP3XnP+sP7ikuGITTB9OAMC3JEj1s3VjIo2sjCxVU51ToHC4
jLn0x0qVVzYB+P6FwTyVhknA6SDM97yKiAeNkfHyCK8P2JPPZyuAlidlT9fNz6Wf18hT9exCTr9K
c2vug7b465RpuB6DELJAxCBq4tNt0pal72K+gJCVDClHTQ2HAfQsc8tPn4Y/8k8eqUH9tj9+T8B+
2+lbssbHqyk6EvK2nqHQpvqocV7O2YQIjO6jQ1UlfMIUUb7NYcMFRo4e2t8kBxcO2YRRFfCoY0Tm
IeCg7x6qaiHasVpQyheXR0o//ZRZLHJ4CGbmpUeuecpm5WSkCeCQYKH+0uk0/zNaMM6cSWS1dK8i
jPVZ2q5BlF8+MvjgH38Ksm0Zkv7/ycC93kJTyPH+XfYSIFqVGsbwq9qeJk8QJJGYMi45G6wMxzZo
4gXVOUQqabdJxObePVoHf8EIywpaOdYHjRsRVN7+QmLIKl0U9hoF1IVUhLV0YUFc4l7+bTzy58wI
K1WhkFO4HuilZ0JRVyeo/j0eSBByqW3bCK924osYSl5S+LR89YxZ8LE7y/4xVv1JWfv5FdYtyG2k
Zvo7ZyTjZ7HCHVfTWVPhl0HmIjo7xiWZ56x6G+coD/h6izyCnTMcG6F1xHEzfM/VYk8tD5+9ZuSh
t0pBOhLPDR/xKbL8T4tShCA7GAefJ2bFYLZAtRiE+aMTF0v+sTgNg2s+/yXQmIXldKExl9k8fAJO
cjbtwdO+jPRwrWNXA4H8jKJePgwOtB4TPg9Y6tdFya9id2QRA61+oRiyDmrqq0lpYDH2dCflnKCi
mfNDqDNDCLO8OG7vECFTMlNHkGwV+s3uW2vd92PvSEfw47nG0nLJEafhxQC9O3a/TfcLEQKFHNvd
26AW1HWVquFEmwiysg34FvCuZbqYzKuWdjTrz8nIALwm73vm0WCAbSBN39N9Rz/3bW9beHmh7Hoi
J1RvUPN2ZXySlGgt+LX557y53fLF4ShECszqSieq8g6L76zuVGqDTEHMUShAwSrl4F35cB79cRXH
lWh9ZB3i6213vq70W4/Kkp9kZTOv9Zi8qDrFedDQv9eSr00uFxv1U2bjGIdYroDIZKhzk9v4zbFF
lvXOEgaE2Dlu7rM7T10fCwbIZCvXUa8z7O/zsZ/gj0SgXLtnlqng0t6BA1SpmKweRR5sgzJ505lY
6F2p1NTFJWwNfuYfbqC73Z+HmLEeEWVtteMqtRdztLIBiUFuv087fGMkfZbRHXmaYdl3FbZwMK4R
2e1jpwc32O3M2cDqihCkh5a/3juTRmCMKnJhSAct5rQcv3U0DazsAQzozUQcXITaUWv36fy9khlI
Wkbgs+By1LMbvQJF9hIgnSwf9Q1nfPJE+joLrh6Xq6MOk8dAwcYvIoqKzeSThxtzYjs+484KhUga
W7NSvV6rBv6SspuG5eKfRTwFUfmuwTpDm4KGgRZwpwMUe0TcsJMqPUEEokU6GICsrpz6qxcz85A2
EPW2rckPlxAkS0PiMggFMrh2FlGGSyqYNMyN6Y0N5U4ep9Y0SEcPUVRYnwMPzGRq9ch51CX1Fuec
Wki4oIo+DcXjuVeAZnNimqMsN7XKLQi/1LL28ZWXsRIM4r2a1ANJ3hP38CPP7EX8PuBDb2j0oiL4
xp/2Mi4eetf9WjucbW1sTLS44QpD9dJfUZU0Q0HSNjgaNe8967rzCnKo3yUqkzFksJchgH42MRdJ
9HSigE/xly1xfEv/bkl6efkNfWx/sfK3qRaP8rrC6aFjEIC023wJbzF1MQXfvWDlJXqcDD5x+s4R
5ENV6d0SKFeVfvy4ryeH//qw9VsiHHok6ylWDFSYR1RnqZUV6rSIIWWeHD9zGCpOoiO00wNFWIAS
yhD6RlJ8Gp+XJoP+vu4YlDER8I7z+xAUTBOZCoj7sHZ6WHM+vXz8rz1pCC6LWS6TyTiFFMvzG1yA
pPaAbgdf2Z1OYkhbZTleI5dW3JYoLxYmGP6FRhczIbDfjQQ2Toyb43BPEjbanc3qHR4mtQliBhz9
CC760uaDhzPPNBEv1C7XJpZw792tARKqcOLyDYpD8RIcHfzkuC5EP+IILpict3SGioSpJWU+Qe5b
xDCsmnTO6Ia9rRyj3NGW0h7mH8Hch33bUO3gTyE59WRHfa3ee3NvmyaCSQCwBS9nqEhpXqyODbYi
EV+DnD1RSQAeAVhrUL14oPcswEsfDhBg6bLgxPJH10BoZ4ZQdDHLiK/KxY36QigUVUJ2YqwVBPmA
g5DgbmqLpm12aG7ByT455SUR2hc0vEthv8X7CSyLa0O5BQSHiyhILwlJY87Gvb9EYT0MpjWR0xeT
weyTMyRtMv3scwPA4QA834LMLzk2WreM8wS/89I/M10UUB8DGUagxr8Nd1XXSVUADvE6WBsv5iLp
dPz9+DwsFH+fUldTJhTOLOQjNzpJLYmKVkAwEmaBPFoePTpQ0S//d8kkjJnajb4l+4bOMvJARKL9
hNxHT5JeMKhduRMjcDOhGog8mRDgQv+8IzDtroUjDSzQfA+HiBtjSGTW7BtltXqLIiDDi1U8DLhg
/iK9tH+Ama9iDx8tpeXC7WcY/Tkk6VPrU6HjYTxTaA4nye1u416IHov2JToC821ctW8yyp+dPmk1
pZYVz3f++WboY2/bJR3S038dFjIYuwF5Mo7xF2ekHnOs9gc1/REl+mN6KHcDX8jU9aagzeRcsKXC
I3wpgYIUtCUmpN6M7/+GJX+T2cParI4bqELouhIaZVHTO3H2uyB4u4EY5X7/ND7z46z0Gv41zaTJ
mNz2A2nM+H1U3SLjQDxRj20L6PrnRMBrKMY0nKQlDH4h6Cblax7g4D1Nm/DkAJO77de8MzIIkxqa
vK/i9X5ikM0jVvCSulyLXYwJwwSaNcOrHJ1UtGas4pcHu6gJVPaEQmZhxdfNMHJ7hj1f95LttoLZ
uh7FrVkXFlqfNLXJQZGP8rIuLobOl0CIghlwpp8/3N2Ga1UZUsPYvKbjbaRmONoUlXGI3hn0xf4J
OTbvQCPBM0pke6QaaN/u7nJTRAA6wxMLIPHr0Hxef/m8VbJgOyDajGZcvOU0nE9rnj5rzd+t/vwL
ZgqDKdysGEvbZEfynCKVpMIiiL5ndigkzHqQA/sNkpbQGkqaWK6NROGbpgypw6xJotqjYrItp1w6
cQLIxlUczHV6MLM2/tn9/ZAHLKnwnzNHxDJL2W5fc3RcXYcDgsJrDDBi46+lLGXkwHP9Zu+BCD5m
o3K4CjBGAB7Adc75il2JZi7Cv2lGDLqlwrz+d/pYbJyDGdcNL6y6kJnoy5Ntw6BFdgDHzUKQ/cum
2jaXBhyMAZw3lkBTQVRpnn9Jvdx7rbCM645jHuQc7URKjIDcE+xRkp4muRLvTowmjHTGNXmRY0Ty
fvW/DwhDirzgmp0RdfBVh/V3v4kd9Jf9JLH7qHyg9kd/671e/++RdpcUs/WPTbPRtW4Kr8V4CUnO
9s0kp8VGyFMIlbKLJ6iIp4sydOJEjGPQcuEy6s1QzXxMDoV7z8QSrdyVdClGEy8oyfTqngBO3z66
nvvMuL3Eh7xwJYDsDjgPMTSBAsSq9yQU7INSNXJ/q2LKEcMs5YHFEcCyEhcFdVLTQ17YI/k74UDL
otJimF+T7kONyVRakQcLkJ3OhoPFUOM6McGIDnbvn2hEEd4TvQq9VdIPhK031tlTLrGRwGwChP8p
xjp53Ckvfn1Bl1y/KzR8SBbK803GBAz4m8aEjU033Yk96JaVDAliD/TA8T03YtMbhh7we63vqTJY
f7EkL1sf1jmm0CnGcffXRCuLSEBKykPAGS/u7SQ2Gk3Ipdq/ZJiHsF76MA/7OpeAYDVq/2QZ09DL
/d/cELk7MdIWu+84RBvgE/Q7+k/1jZJWGLIYMcfJuA4D2yupbAO04wOprQPpiYNZakLduS5xBmdb
nY5kJ8fpUbGraY91ypsu3b1lDHmKEOjBlrw4YvqZ/KK9SSDa1VPRSkxueNmW6th+7WVBtMmFcUPR
ZNY0GeAWouulLuF6gkjOx73OdphzqDyXmkRgp/bnkNg1F93D0uWzf+fVd4Hu6LjmtqBhB0nG4fJA
uqx6m4I+uK+wm0/yIaib/Cv9oFu1SFsMDgTaa8j7pCP3Xy/bPfr/QZOImmRHD2XZ6T0nwCMrzeq8
C8WVLeku60QdtM2ANdWpC112j1nXVxLwSaPWbdVY2DpDb1KHRl8bZ1bH2fRlh9lAwIo1LVDQofwS
0kdhLXP4xoRQY2J5BKwH1mqUfbvuSI3ORYBpFlayvIjmQBDNgG3zxXeoIuC136uGlevaEtN+NwVi
NIw/W1QTvv/RRT7sYX6tepn2IKXW6QLOh3XFOh1Vmr9G6wZcP5OXXsCVysjMJgHH0FKsEMYyumkk
gqmgfCs8o7EHIsqLf5bxuLJjN4gZEkte30NG6Cz6zCif1Gl8jujTU6p7mlmuGP+sDxTjWKLgaTHn
2yH3tGj0D2FSW83F4p0juRiNV218CoHlELGLfBrj45JyFhlVE/gG/egOIACKqu5PjU5913FUqYJj
sBBqOADg3Qn0kMpwZEFXc3wnlF/yS9Z8TBr9UKleCMGCJwsoKgU/98pdZKsmwkxdr88AUYOFylIA
SDcwXoY6qx2hJ345flIM+kDbWLRIEr9VgXrJcUaJw6+zALWM2HpJWwNG4/lvMsG5M5yyRLY9hxJX
4XWDnvXY3uXSBR3HaLwIVmnHJz4hbnb2mJsZYvieBCy4xV++MX3enbYIwn3IgIEwhUObgXx0S8ht
RXDz/5cS2jDj7zSRAu6PFbPffo7CijbRu9KiIpH7JMEbAR3ak5C31O+Fd0roGGvgaE0x1kbGWBA+
ubT7aoWZaviBZqjoXe4iVqlA4cKJ7obf9dnOf5FCEbfxsXBEOfuTBO0qNeGDoDqMKF+/U/4xUuLs
3hfWyNrErezZ6Zprdw5f8zNqsb1RruL2Nr8+nE2dRk/kfxY0OmVj7FNp/MRNk+hPVc5wgYzUpaCl
sAt8yeQ4nVtzvHRQtqOi9NCSJvoMPX+CWE4dIV9OCRrQIVdTCknHb5WNGIIeqjp6VXcO7nLHZfpY
WqJjlscLeQaocEperTy4Q7JfFHr7o2lJWaBHp5WJJKYqXkoDLdG571geIFKPtK6y9Q9du5jW+CV1
pIKigF+0V1+Md5gKeT415cHIVD9+usOcY09PTJPhkwV8eCZfG2ZV/q1kxhWO9Ols3WHtmZ4VdQHe
66BDNSCHH3ZyQr6VKH3BioasdBjdPkf/djCCqjrRwMNXY8AqdUDl2T6NRTztYkld8aXXeuRXuhc7
+ikvJ2WgGeit8VfsiJ8FReD75kd9W3U5wJ+uc5j5WzNWn/REwMcbCv4UgdjHJE0rAkOv8K8L34aS
O+IFNHKU7OUOGE2vmN3XYzZMDu5EfoF031FdUi88azF6n2Ecpe/JDkrBiA4I6Sf7BlD9VEu1sddB
GmlPHwy0kIlGzjSz82PZ06lIXE6ZLzKErDsj6/SOBYYM24TvDtZKt0V3GfQup+L3RmVKx/1SRl38
7+vBae/AcelAT5P9Lv+iqUoTNOXjY4U8pGNTAYeYRzXAhWjpgDOndcFyfxBcTJxZsPI/h06Mxx+r
kHHxGNeEKApdmv9EDZZslzCR7j0eHBi90h66XEeofy2SgfNgYgfom4m5bRiw1efyHH2iWMF5o3gI
cTVCGVyVgE975Abri3E1wP9vxSx6Kk04C+8qDhNna8Z2bl2JRltaWZZwSqD1nwEO3c6KZ4FuNwRR
o4ZVZwJsgbmzvt5BM4fFywvtfrC6xjUO1k9pBgcHkuY4syWc0qr0VDZ43tVkNiQt/mliHdBnoPA0
gmsdo7dT58tMydEY5dwd7MzSRWyeH2wyvXiTtWKgW5pmDtofBVYO3pBsxkatM1PRoZMQ8HH2tgts
m+25/j1bq95xBrAq3lKjSUiFPwfWm8Xsf03V//i1+h1p+YBTXtyb5NQSRAXqMQX/3R4qX54SGKWJ
wPXOp7X9LgxVIGqOKlTeU2AJFol0o9esHOzhfUDam9a3xnbHg3/8GdweRhS5gCls8Rf5R4PX4Elz
I8AuhxFaRJwC8lBtXqgvOUQ/+GzpvcRJG/OH53GuBB59wh0dZ4rTaBWbQkLcOMeXLDHgmhi/FUqO
b0D2lhd12GnFBm5ewZV4M4fxc0+oJV1EiKcIhc2WcXk7jNGYt3UIo4/AGcf81Zg+JtZWpt0lLabc
UI+6UYHR16r+686yl3aJrgLdl5/RZX7btyUF/dXN1vXKzEwcjhRydoqVES9ymAWdbtHvSORk8o8H
cjS/BlG7xOsonjdAuEMSvDtcGUZ3qW4UT0L11w4P7B5Y+KeDFeKg4lmyqyhjW2qlbhMgkC2KW6vp
4bDLj4Z7P9moaXNgUD91wyWPyaqxpkXp3owWM2Zlf/O1vBrXz3QPY7SLe+bvsg4yWauvpL+De7uw
B6hxVNv8Exdcbe5ca4YZqdmmhi8VvUGcQqK5hT+NQK3pyClcqn5ZOf0TuSiUeHVRa8e3Pnr6wcyz
IoEMw4EsUDFIpWnW25C9g/lKdNfr5ZpiH9RKqbPYgBY/gkd7Sbmnq7ROqtkyphZwNaVIknrEWT9w
rTkKMDbv8nlX+RroASIxoLMEMAmx0m+K+b9GYYHt10Gg2Q56d+bDJK5gZtwlivMlvzkFZY9IKEaI
jYBbRYPzdTG+V0LF8f3+x/g9x9vSMHXY4iZzpPnYrxWWKKyVqmOdrS8ra5zloXM71J4jSlmmMkRH
hNrRhblYmX1/jFzgNpqYtK3DHCQcPW1LcAW8zWwXsv1sLdtUXm+PMsQ3Mg/4coSJJ7nSAP8yp6sk
BGGHxqs75vWZIsfAi7D//fezwlbEIhRA8Cxn8BbCowVN1j2em+GPxP74pqJQKeXms+WqHL/gvDSt
xg9ogRt6rtwN5HYpw6pnaDLTHd+xY5+G81CuAwHSf190Ld620eiN9jvUeJSpwjRg2lg2RZ7+py8g
qWaLUitA0PMoHi3TgigqLDQyle1ffTV0rEvTRhC923Pn7HA7I4HfUrbI93EPaWiH3mg1Kp50PG1R
bxhct0/8/V6Czeg41KgpdmRCUUBAMpkkUW2IHjzUmf7DLa3qsaZUa3ST7SqhpTskXzCT0QXrWXzp
bl2O0W8r/id8GNvFfCqWWXrJUBWYY3dWhrXb3O6Mg+fIcL0ORehdja2lpIDoi3L7PJeThXbiCoST
qMGo1cLUcWZhYo8QAEjTenrHVEXgLYKKulzghX3ro81kJxKNtLXldpz5GGI/ISnJJubjG+vXq9Mv
auE4y4zqiNJYHf7uxLG8cNOW7B/tY8P7/9Kapkepg4jYxA/BjFE7ZC8bpOQShzI+ME10tLukHK40
2iJKmFm6zxzag/XkUmuKYrul4xozESE1wOFsjGrZMRRFqKJtDZPfijOz9/t73Eulfhbh2VFuVi96
bGn/ssxr7BsoR7P8aWQ5ogKISORfxTsfe3VuAbgfM/9UErAYsOZdr40s4XL4JBUDCTzotKH9pIx2
EI/m1Bb0mhfP8UmGPt2awiBILuWWuH0SYAw2tHj/sxsjRkjy1Pkv/W7DWHLDBU0heUJaALmDNFxT
/kPo4J6KdsupL2wf89Zr0+tdpFv4w+gW5daJSxYac1e1ZCcxcXMEhK95m/JN9/xl+Q87ecpUsmER
rYngb1MrYOMOyENTej+Wk1T0Yf6S5BQ26CatYpP4qyRBjGrVXsqe09sDYI0WSLiDtaidc0do87Y7
PelDD5tJ5uR+dc1w5A/fpqFbsop5Sm4fekR2cxcZfZUkdvpkX67+pFRcmD1x+U9752k7EIlCWiUd
sUwvBgV+E9XBsgCnPamT4bS7d+DwZzHXqx2cUwIQ+53ZIQnG1+tYH3ReMYRkOmJchgPZtLz+F5f6
WQOnTzcD6hdYd3MBcesMdVOpuT6SqCgIKVWtUFS3gIUK6PrKOpL3F9m12a/P5tMCLSCFoltDjNul
m0zdK4GC1zN5VDRtQpOuqc3luS6VAdVWdQdpvTYV5GPOfK1crXvbsYUKR3hr7y3evKDxz8OrhrGa
diLFuF1STBjZbv0ZEZwI0RcbY/pHGmOXf64EB0deARZKhD3I+Rv8zCFBeUVM1wdlNH2mZnu7Cbzu
oHg5rpLO6jgJhDGHrt/vXn0OvcMu1+cGmqzPw15n78dXcyHg8GzeBIyiSf/YfYweuh6yb6yEM6kl
NROIv6KbVCKslMJSVU8CTkiVyiy8vHLBJIR1BLTZ4G5hL/4CthHSHGwBVHEiQ4US2gcX8r7K7+vg
Uw2VNlSBa14HwXm5bgaMyBopVRtij13pTMFSKXzNVaWwhZUbBi9xtr5YOnniutOchNCIzX2xpNbi
9lnpm3A6Vz4uX4/4i0o4JCOHwAIQf7dCJJjBXWN67DfE7VlUoEY1ZvRIhwINY4CKVpOfnLhiOgP9
rRUZrZ77++j5neIM3Y0Yei/WiGcvF2L7gdVs94SW2phhnUcq5vJE5Khtw41wowzxGLBBahaydrVx
X6F4Cs0yTD4I6iWuFa9aYTHzTyz7/oBxsscS9gf+muOICSAGzpR9IGBQdzcroqn0+ODVJmO2zZXx
CPbDZ+kl2vMepfkfX1o4Rnm9tePvnLoNsjBXKzVhZpbcTxvkLdDMDKAgc1RGOLOEcjWTjbM7aXYh
0EnsvMgtYEeMUmuSO4s3SwLEan+v16swwtI7GT8bIAAGsrk6hADwMUNTWSCUSeQzEb+NZdCsI9ZW
YVrydgveosXqtUUP0THhKX33mJUnTyyZXs9Duj6+b9DacrOsZXP9UUm/076ZPMKt68DEB4o/LWUN
yGOuhtf/OwQqw1I8hfWya3hgFQilkU2HAkRznnX1+tKkb3dezcmAhy4hbwTRHWD8j1RQP8ErE2DX
WpmF1Sy8qJL5fOwDHvtFkfLCa9QVQxt/1lUgJRYubx1fjKS7RsRPFUMMnn+FKDeoFrCY2IlOq3qj
k8yLXoemRvwmcx83mgPoDvfv47R5Efjz3DS0GQGdlVabGyUwFBfcYOyvQmFOnwu83/uk+WIaQl8P
iQdjw1BmYEvtAGTCdZYMBKeOa8cdl8CwxY//hK8tkaWJRW0ajMPfyED2XkxTln5iRq6PheOQrxQi
AzPWTWpL933+DiisimCb/gpjW45X/5U+YkXN+obVh+ZK2CDSiDjAXOFqSNGH+FRBt5fI9JkqOYJz
2u39Jr499ajbvegxTO4SOtLzXg6GE5+c9qB5bw191eUFckANziH+OM8m6AHTet+Cej/ewXOPafcR
akbq+hE9AbxhAF3zj6Ayr2kkuYzJLOCe9SnHtxvkw24V4ezTfF2IZnERBODq5xeP8+CovjQcOq9I
ZsUHo9jlCXbMGlKqDJlCIXjwhzWtFaTTqOLHFQhKhwanOYhUjk1D0u+1Ym3E0EO260EbDnJXDmgG
oQiEm2L0ckYwj5AqrEV7xB6U+qRe0jQjMhrE77b4eGMXTLQjgmMWFIi2+rA22yKi8IEkcihptuqo
G6Kcpf210zH0INtrpKzplbymvLZ8JD+uviWqLiD1X9PJg9J4ONjWsqxcSv1mQZuQ0o/aX9Lpg/xa
w0VG3YYql/fBCz06yk6AqzncSuHwyvoDj4sRjX6ST6rVkI7XAyRIibrc2PoOxHMrEfoqCmIEQojx
+QK1wHOI67yvTFWOjoiJ+iSQEyiHDfJOzCUZDfPCpg1rnv3TdNpFzUjNI78aURjJ95Bq5JPoURMV
/Rg0K2cdP30Td8dV8y748lO2x0vjlyh8ZmwHzjhd9043QLB/PDOZZJhqh4gRyn/3LSpjj41PITq1
VAe7dXUf9j58w0UGq38P+w01n7oSTC2zYyHxHQSrfQfEoaPnro5ar8uYGuZbPHheu7hQqUmjqVIE
ivDPl11UJ64+j8hlUw0suNLS3tq/y55oWaLGPDTpgdGjmhjSqWiPzb0VyRnX5ljoXri3WvpKBmQQ
E91t8drb3E0GA1/gi2u2VS/7utBMhM6Mfg9O++1P9dripJZd+qGEF8nrMci2be+tL+Wu54uufXcR
/e1vJa7BkXEKZ+FSzi2HKdCEkU5rNxhYWXMYbc5/4l6eAEFQ+Q5PqEqpNDZGGxj0OEbfAFq+KjVt
NODLl2t4Y0nQCupGHAssJ0vcM0oIt+S0B64MyDaqVbhBjDwnOL3HOoYcdY90snJ6HreZcykviGRe
29jN74sc7cayU/dzxhV2Sm4fleJnSZvt6VRrofHaZt6fHl1dVuZ8B+6OFUcxveN9sTHnOvfoePh8
voHFTjpUtjHyDrwgPff8QqNW7DwwKmquB6cfDOuXG5brbowIEtM+oUV0getztpiCOW3fKDHSLFTb
kJVce9bUWHNgwSFVrJ9pAxh/Hu7ZGcZdTkZ1BDvqBMQX9jKUGuX+kb+UZ+0OdLD37epJYsF0lcz6
SRXZVnoOqHxMLZX0ia25eGv/eNEJFaDlLnPRf9btI1fjFyQHfnr2pQrSqqwG1GCAcw3mJpy+ZZbW
vJRhocIJBCckVdfzomnl1/vgS7D2WOVbNwEngDP6mQegUPwR9HjtDLl9Ysn+FIGkJ5igm9nMU26w
ppCuZxDIsjJKAs6f8Zy6bX/is241DCyShm9U9fgBaum2Jdup10CBECgKleZu8O/mNSOwR87WsZ7U
MY6LHdjIL6EgoE0PCPoEtSSI+FRaSImdZBZhjtiOTamJmLh5Zx+2FvFnztcgV5ERPOiJ+iMh9e88
njy10MiqhaCtQ022S5ccuLFQ9fPpvaU3XJeT+2XD9DX21zWupxllYeSsWY9e+ZBtOi6GSv6gl5pq
H0DJZW1f73SzThaLkWWmqoH0wcmK2JnPnHa9QfB3efG5b91Z43aKP3CR8pjKUaK/HrftataqFvqJ
8C0fsP9Z+RG8/1dW79SpSjVF9gxLOth4YEBkdZTm6OP99YufXy5NscY/PXRyCbydMHvddY/aSAkF
PohbMmqtINn+QJ0RwPRoUfROfHp4YmmYqbf8VB9hlOY4xWNpzBKCyhhWHvuyt1ZqO6hKcAoKVAbd
ChT5NcH7VhrZssThmarWdC2ItpgtTW9IWe8yB5yBDO8esc9om50Y3Y5GH5a86iaoR2FQA2IwBGV4
/ZRzGnVEabRgvsDFcSxL7PdMsiwqrqZwzWlt6KrrBeDeZtMLgmRZ9Zfdc50i7JTuWfqDbxM9chun
rh/NbTCMIetn3Ael5b3lQDTKKH8VTMB47tlNpS/tUpPujJxE5/Sd99v/11MNAYn28QLaWtF++XG8
XDPoCNUn0twEYyxOnG+c/1ECkGDt17VyQhqgF1jkw3AsWTc5stkqNuLT4RoOHYAag0kRIFzqsQzN
4ehWhBklt1LbP2t7E3DCdIuuL8rhjVm73fltGWM4XTZeCvH61t2Kp0nSec16seU9/jWolRD3y1ct
exVNguB24T1Xv5r3LMrzadob/hm9ROWrKTn9EPptOQUXmVn5YD1mxILE9NP/Zr3jBRvjvaI8rWDV
dvbqsCZEgKwQxTh0sgNTnQuoQ4371Ren7MF6aUsWuxkrDoo6pEULtyUq2MA1zK+lX3yiVpmvH8Ou
OB6Yxn2EyE/ADs+kbVpuTcf8jzHzZ1YYuM1KojuIZI0y3gE8q5oRlz1DjB8aDhhu5EG5DyPaODyj
BTHDybCsugZOquoUbSxPNkbCt2+tXzMUDrpm+zWrZcQJ7IBH9q04Z8+JhnLY3lwH5DC3pD6eOeqB
saFJPhnMvuHUxyxmCUPU+2DVqeG/9zedjyMel4ZObeXRfbhZn4+kK1UgBL4HXr/ZFFitSQf7GAXL
p+j/o8cKNMb5fbsq66Q7loMAA4lZy+5b/jhipLudySJqz6YPd4mU5ZNlslfoe4CETStJhGWgxf2W
St2wrTcre3XgU99czsqVG3OvVFtqgFEzUiBrP3/ME+dLKR8SonBlQs4DkeBhzqC6dIkClvdFIor+
+dGAPAFUjjHwmxk8DntQNW6UA/s9C8jYMyD6NBgde30u6iI1XUL5Q3LYRnSXX+2kZFhvIFwUSTfW
RQFYT3BxfqplDfvr2GYLQVETKmaNpeO+YM61Nrs8Oe1I0Nf6mttATG1gVC/pGRoaEyvG+yepcTO+
P6GOVxMUyh30VZ4SanrCVK4JDqv1BEbmW+L3l75VDMk+6JH7xqHsQ9+9goPc5BUqheB1FwUU94lU
PviXT+0/Cww+Qh/l07yUVjIDpBjUn+qiUCYiO5SvlSsh+Ni/eOiRqPZE3BS6a0e1H1tDmleCg4/G
1kjr/zmH7KoqLvI4OgbPPxa27rS5s+CrVYO8A6JG+NHXNL5itXOScoDcpkzOFLiWrI0wbZfvXCMr
qKF7cH6zTymhh2QrOxKoXVANOYpO6OVhpuKM9xYMx69+xjAXd/qMJmJCcXd1Gg98i2t0Ar1ZnV3f
jzCK9WHYenpmZdRO2Nvrrr0ZM12eso66p3bXAEZGLPDXauWQLtPQq0TIYW/AN78x40I8ZoXg/kPd
VT7KlkXPHnRfIIvJkp30jGja586+yBrs79KhKmKs3CZyORtUzd0MzAD83riEX1XrqOtucKuXVRUS
BOvZUFVk8k3qimaRLM7XF9HLIbmbIagKlNW+uvRFM/ebOLq//svGxxnhzzIdJ3aYsMDLfQ9IsukA
UUir0kBjhdbge0wMiPkqJC8fmobwrW2dWK1gLIyHfFh41sEA8mroMJ5vMsMPlpP5b8Nb0fMFLoHm
L5U5zeTKLWEjwjBrZ3tkb+tG4ESV3Cwa3jEJfq59+ayaAlQUj8T0DbMKzoT5tF5voKKwtwDEt/MG
JoFJ2tyUu3USSVCkoO0sHTKBTtCfofkguRGy0LdN6zthZ+In1GTBZID9tPbVSOG8oJFvDjsi7uSq
OHNIpdxTb9hd2jpfG9olcklyO1s0EAO/20j8rGOYMlO27NMVCJIJSPy6UHpTzQbE+aNC7/1S3z6p
V+p0/jqVv1g6y1T0eDF6F6HpH5RFb5tXgZ9w4r3yNuZM0YNuSR+C2R2GsagTUAptV4tqjf/cmCKF
IP1lYeGYf1pu+tbkGbEuY/+wqh9FI36Y4Jzt8OXJjKeV+RF/s7VsEs3bf9rd7An4UaBD33YyKAdX
wjoeY15xLbT6eYk7mzcMiCC93g+Th/qcgbIVNLC8AhpCudxNcUo4FVsL5/fBdWubMoz+cw/5MX7B
Zrk/s5B3iBl3ScsjurdxDCAY57RIHWj0pqsVsWR86B1crZWc/lgmqbGwrx8F7QmPHkPjyjv/SO/E
+zngqhnf51abmbIPgP5Lhkmkn2oxO3s+zdBz5nZm5JjOQvEO9udQhEFGcqHow1Mt3yHxqgyjmhyh
t0fLY16mzMzRge6h0r+TLP+Am8NM26vg6DdVbq/eI/B5JUWI+qbgRopinlQxajsd8AA6zUVG5/YH
PPGo7K0EX7o3fEJy56ey1z8mHEWt1zkRIFzbH4eS3/EcUvd1jZHd9V9Om0M1Jos4zis45m9WSm4Y
tUdeTjJRS5SSj76u/G3y1XQY3YnAY3S4A3kghFPkiLIQz1n4gkCAXatPjKTHCXaQIz2cw/UyhGhb
+WGNy2gx7mcvCXtwQ3O7Y+w4fZHG6lz3Ic9W6/p0smAyOcSo/+//btxFcPxy2UQ2G9lNFYh10mxp
aD9oq+0GyWVL7DpxICe+2WQwIXItDreLzg2cToxaU+0nbiIwVuxvxqdsZggNaVbnzFLFH8CX+aWe
HfbjtQYE+NCTyLysqojbqAjnIC/P9KMe0pY56E5QUjok/hajc7FMIDc8T8gIx6sW5EV/G3d62VhM
AeEW/3ecj5tZdWMfZH7XFgxi2mV/MHCSgzRS6XTxCzZ7ktKQFP7g1ahoseDxaHwyGBb2ly9yPEVq
CxVlUE5GJ8YhlpYQxKgLjatiQxT6e3sRzUMjUQBRbtQFiFYDP+7mUlMou8RStABYPHyLR1xBesmF
wlQjY5q0GvOugh+yxAe+4hBNxigd4HhAo/mFUGsAuuYW9l6RL2yZKSQrCOiJ91hFuonXvpVy3MIH
JE7SygtKD3tRh6VFMI/ONRkjwFudQz62egK8DHGQAI+b52ift6rxTevYoAwXuQ0o5sNOSTVgwF7m
0meWJ2WDTjF/j/V1lyBPaj80U+1gPXETDjkhwdX7U7ye/QgAC9QQ3TdxSDpv/07bx7qA5fC7b+5G
hAnVFcMaaCh4rhOqACHJFbTwMmkqxQ5G1fxPhwKAstfEIv0VB3vyqNNloV+vKWO6s/Kv8vyQv9XH
9vCPSQqDCcc7+rolymiuYGV8i+jGjdiOmz42NNEsWz5oilBuM6cWwOEg7C6QnPhoQ0K/xnJ+aF9o
1MuNCvGqb9a2dYvh5GIMBRXhhmZAe24m8BxzJm3nQif6WZYioNBoRIGOyj9oE5DXG6hXost1a7Pu
637J0sD1L5S9pk6RTG5KSsmkhcqidf+mjcfBCaPBdK9NXXE92w/IfABmTirHJ24VM+jE5SQKklyh
iUue4ow1vfRc18f7M0nMr11HmpXRmZtjSX/ik9wn+mL+S2kq7NrXaApikPgTZi3OqkTz3X/opu4n
M7vQZIkbzAi9Op7cXnb0kMkuz/raplmdNnL/+XFR/k0g7ke/OS1dQgFR8EtcYnpIHtMvI11/mv1g
K7H7LAn7Wtk1E4ZIRZTb80Y0Lc7kHXX9uvNWBsYtyUI1WPAUKacXgIovB4G8wxsbMnDIGUSlagb9
3pVytHtkXKDEMhoo+/emQrya+o3zKoqr1vrn+WY+UchgmhwaWzTL16nzA42bOl9UoVfhrqcR6x1f
UHdHe1hLMBAUXbxgf0GbNECmdVBOCons0aXuRogWHTca21cWdtDB/da2Nps8lSxc2k/SyVGsKtgX
pUlLnA4Xx/ZydgnOwlsoMGYksmGLbqa5Ge56h8wQsnblxQ0Brx17BL7sRw2Jpd6Ds4Prb1mRzD3k
NPCqvzH8o71XOlDXzj3ZZtXpsz3So1RSM2OQoAnI6e90xmeMEENiivgqlrjor4VPiFk8MIZAgw5s
StlIIe86QlT3ghiKxjDx9mFo+maZKAUlBYuCHrlJQedzF8oj3+p4epf6ye1lvD8z/kodtKN+Pzre
Tyh+3zct874vfizVZrZO0qtfCmjLHWF/0+mwV1mtnrqYPLXXrqZqBB0HtNshESJHFNc2FiSx6E1i
xh1BqxBRGcygTdmVaWT93HTWCYZGbamR6t3bV3muLBtQeGXKA78+roShBignhDgJzBmLZ7rcvUlg
skJZZQouMFqVgVztexVBOa3h87NhsQhLKEyBEWESOJKqv3PGq8d4OqtC5bFgtplsWGVh3GRybM0J
lrVfJgZmOM4PEoZ/8mHt01dB2xgL97wbRxir/cOOrKpOlnS2gQX5REPZcT+8eMa58EmHI5cY8iGx
srpK8d3jYeOn/xQ6ULGwjwuRJGfco/Bfn0JgNzGGmmjZnTE6GKqorwIHDzpOpU34yIuolwftSDj7
+zNdERJtus6rHW8aw27/r6NSRLwcZtA4Staxaz8Avxvi5OWijq23TxYtG4QdFa3w1iItXBMMWKBO
e3pL6kVxy9fHIaotoefgzs/w6Hxu0bAEkWYmvsJDwc0TK6+b3Fwj2WtOi7M53pzze/fwV4alf9Sv
HU2igLKeF0IWNJEkFZKzuO4EOmkct/lu8LgPNyu2SwSxxvYigvmHgSk1mHyJXz8LXkdMKnFGdj9r
E/aW97IawsZMaYqJJDCHMMLFnphv3cciuO+oMJOxVMDSmhcddNSo6jhbqEV0Ek/t5wwhwKAylZ36
zFnKPFUS+nlryyK9h0H9v8N985yCS0Al/lz0VH93EYngdp6NLigqlULx5edfHPBy/8J/9m76z9rQ
KKMjp5LLcTKwAHPjCuyrntS56hDXZAgps9B5o3qMs6fC87uQct7CdgVsVaExqiqLBV4bl65yfCR+
N1DY7h7dA448caYal/sY8zbfcI6SDWXxeVox3cfCVeHQACMJQXEgGLS89tSf8lV/wsIzbPYdqopR
eQuJiWgCNHHiWP2fYd1FWWkftGMBTd+7oaefSlJ9BIvOL1OFFkGpWOft5C9yRE2hfLcjxdPkC/38
cvNM8/CCJU1X5TIAxA7VDidNyni1RmZwDRZimN5aMv8hVNk37J7tiq3QgQCC2PGPjum7yq+XbtNw
gvHFBYqZ7g9sNXVrf2Epmt4kUuDKDHCO/DQU8jc/sC8C4Uc9yS5bZf9MivdjyyDkgHun6CglswLD
b+LgoFggzbQO0Jx+ON26Fkb0wBZEqDKXw6N7te6wdJM9jyEr3Aa2I6Z9Ry3dpF5wHDupPTDak29e
odVeF5a5t5u5u7XNi6dPBOul8lkT8g4/tEYmLFeuxrZIeOIxDl5egpBGDjWxOxWlBmEudU/OaqP6
r/Pdq0Z+QtQ4dbrvD75Dd/2rcaKlMRig6Pexs/T3AmYNo1yCegNI4j9nHBXVkPnRa7EN71k9ppTU
T4qLiSG/3Bn31My9BQ2WVOLgAFojedItVjr6iYBf+RAINtB4dUI3DLO1qkXIKeVZsQvoMa1bSHxJ
8SDnnvxOkhD5U3EnNHYkg7eeA/gOhTobbe/0cSH4LytqBYNonAM35p50I1dlWghjN149xPmxqwsb
Xfbx6ife2VP6GJj2iQm/QS+NaXW1t3xLRd6c8zIXBND0EOvEcGMkg8jyrbhyLE+DaqHMKzAdbUMd
fecdRQCDnVZ7mNLbZ3uJkfhRYn5Jtd076nt2B6MT/jmreiEc/Z81hPohCFKn1+VKkqpzI0iguWct
ioWKppqrsE6Lm3LpcfENC1CZTbRpHanULwnKIZ+sgDmRYCcUprgajrz17t8A81gtS76IlxGfMRyO
Dt79QhWwTrIFbtW+19oYNlF2coVAZC0ZUf+BvQvTHH69ke/9kCVhaQGZIKMYYZuGLaPxnqSLrk8r
qf20e77HGlcB4GNV1Be4dNTKOt45ed59hiABlojXRZNgELbzaENBPFGimlNjj3HpkGixdgYzCXTN
l8o6/k95bBebBYZbOK3CyKG95c+/cjvUtnWSbQ7XaIczq/kYRgn7dVS67k/QQoi4iaiGa8gNkXw5
A2pc4ulKqoZv0r7wj+aZbayfgihHms0xafl/KgWjlbBoPnxIss5SJx2PqfEwTonlYPjxC2NinsfF
m5sog5S0w+jjndU1nDoi6Wb5ixk1OPrFOCOnfAJKkNyGS95pp6VvdtKDd3ZOgrFed5gMRC9RUx2s
gGyg0L1jniWfegcvC6BvY/3Qx3z0oaI9tUEhB8iBxdd2wt1/MKUQYWN48bQg6GD5iJHVtOJSaplg
tME8RpbLQXkLwYsBVO1B5TuN2114n0TxPLea46tD9gQ1r0TtNXuvjbjoTdL4ccLGFHFxrUq0H/7e
j45kBCs5fWbvkDiQgmV1wZ6VBDEKun7b7Wx0Lck9VG+dtWgSsACfmFC2smH0cXujt+KaV88b/4VM
+FdPPZFj3azKvadUlMqjdxmTlBwKwcSmYTF0FK09K7Sd3QJJi7nrSQ9/5YR3NNsoxHk+I/Me7F6k
528/tfzh0GsJXclRPIZqEjvuHN5m8SDgdr8kl95JQMQKbSZ2qpaYxWqQdWmxNYeE8/0J7iNneY0U
zPwD+rhRwNCSknfHx16/2Y2S5zIb2+6sQKZpSNL7eYTrSbluksoVtDUBnkJDbcLG0Elbp5haJbRY
1HoUaJ5NqQ7O6k3tQFy4JQ4TVQ31+tOBPV9oJsKHAJJmhQP8xmJrmP5P79xI227kb5O52fLmRNHt
iNcM8wzO3z6BYCu74LJE7QcvyElEjSPBU3CKc4OEdJ2mD+ar50RrD+YdyzG2RG8eV+S8q1C07dO+
5vxQjneYSFDBKk6k5eu7NlH22Ugv3gDoCoit2hKz/qLv/vCbVCugmLdt8EEzxGO7/UygdrQ781Ej
AWf4/E4j98/YKt3rH3U8vFqYL59Bu59nkfQT7He4ZarDJRioROXIGSl9NcV0y2IGoSm+n10fieJ/
nsUUGldgSEI9f+9znX95zfm2VXZwdloZq7Uy51kzdacFqHhIn79Gp5pXPsoBA8MoWCRgjzOsIixa
QkQOWhob5/jwLq1wRRMRxjbrEawIieJ2WC7P6ppty3H6grI09OBlIGGihALdTPIexUbmTQ3PWEFp
cJgfEwqfIm0+XsjqQMfIdJRxTdyDSOsU1yhZmN6mfrJwaS1aoa8QfEExPv+UuMrw4XNSbVkLghMr
oTos5NSKsoc8IZSfknkPkGQskI1cS5aNvL2lDE9axXTAP6IjFLE9gEA7arN1KBx61atxipj8/eex
DCytyjqndkObpEAUkJh9Lbq7xuBlWlwL63QrciYJMImjp3caF8Bs2VTiHH6gqpGFaSjQbS9v5+vo
72B3ZuwR6H0JAUbsPgWQYcCbqti1+CGi/N8m2+t4U7VC/uV85RU4ShvY2vVFKiW19Ld/DF5fGNdS
mQWFr0sEL2/GCU0nYjAGkq6pNFimANWMGTAKR1xazFMUE2QYGhyKYhHf9aynm09sp285RX1k7EAo
SGU6lfquB5Z2uZ4VOG56BbkyKEWkaF2sJ70Z5bcG444lVYZ+SjYb2lY920YGgHgj2WTkx/fuQ5rD
VO7FmFX8rskLVj+ApRkoGlbr+3i8Q1mxZoe1PhWE/e0ntca0P82Xhtwb2y5CWmnQu5vSVxcC8zZS
OOEshs5pOC6LPpdp4cr5Saf57FN3wNnfHZ32a71xXEhL0lqujfmLk58I0hmTDHnSadsJVZGyjnko
lqUD3ZYtg6tTmslYMdRn2lx8F3zST4BnP2XKfVb9Ytz+1A2Y+q9gVPwu+jwHFTdboYpJJWdjNWS1
sfIe09iNFAdLEXHrAsNZrjTchTtd+dMKiZZY28G3QXSEb2Xd+SZK7zaE1uzXWUG8OqA7nIFBZX3r
rynN1azxCYHYxYt0Sp1DhMOtxiVqF9FtgPlqu+Knu+OguqeTkK+UIFbWrVlloCdibI1f2x0P0CD8
f2E+xfhGMAA/QnVV3VQrk3SidVETjPghfk+5HXJSzSWJzv6dAY9RjN3lbUfnxVkElpgh7ecAaMo/
I0qDjeH6v5ZiqVoo3KCFYh+W9fsnPNIwBm515w+Frd39yAI6eyaEtCltYAZwQzju0S2ki+GTCghh
PYrl3DOte+pbpNebKyAkrPqGwrsllkDXRDyq6ApUCHF5QOfLZj7SDpdPN8+4YN2hKNfJarMEl/lV
ADQuYKFzO37Ji/Rvy99Z7OnB984cpELa3gHt6GHjDbwspz8KaW7OHXzixTrkt4AbrxMaITpLq2xj
OaNg2s0Y5FsD1if5p9RxY36QfHmoNcB+xskywPh5Rj45jxydm1ZFGJNVXGHQQeGfcxUkxzJM8Qzo
u9Wz7FIpNf/WTVCVCGDjcwhsfn4A5TzAuK26s6netpfM5K8dMS6cG5TUpBOnDOEzvG39bckl0xEx
5+4X/raV8SH7pmqb1WqXh/tAMdgtvi1gE9LFthiVqgyJ32uw+XB16SXhdGX+mICxNm/4jEz/0Xjc
3DTNfn2M1Da06zAVJ7lQ74QE8ApCWTauiVzev1yj94GWQUHC+CFNvHPd3YwJtxFgKRk9JmJyB+c/
UdNPmLvoKH5OqlM24gW8hEreu4aCAT5o+vfb6LQX7ePTdyFcDiVXsyvJlkaDPlpWqtcPOcvhG8Sc
wo3nzlTVZzN4YOVgMGQhq35O005DRHmp2cZ0rBnOo6e+cZa32qsX8fBAgvK/egVk5n443esunDGf
pMoRHrO4tT4E1oIMxHXm/NOA/HWoD46UIE9ROuNH5xorPUflYfUfoE9bZSXjvG6ldd8l890cs9hR
Um7ouDlAfvofU8I40alYRVfhgwRfIm4WBhi299Ecn9wzJHzzaKKHCSx7fXDaTSyZ5ZLlZSj3i+Va
Gc+SH1gD++6HTwuBo8dkMcsX9+PR9i5FPgRDnx70eyNoCdDEbOotIubfMkJFB+qm0FOYxhGj158S
wTnPl0lX5J+xJujqXHxOlmeQYHOekh+R3+rNoS6HtXy6oKmrOZxknhVZYO809Kv5EpboY2eRH1hT
YiyGjgKRqXW8aCip0Y+woEKpp6zvzz+17c8otrZztCdp0KZtK3o66wRPS5DaOtx2XU10/6e0MwIr
mZ2tBQR/nqHX2msuVxvKnct2tcz8pw411wZ0bquKziiYxTp5d+KFkyPFcxLkOeuFORo1BliRDB/c
P8Wkgt2iALkw8zPDBnXitegWJWtsmzGqEL1WVoQJfj0sorgb7UkEdN8fKsyLn+QnXeaQPNgZ0TKQ
3jppOgOwTJKWHxk/8tL/I1RJxYbmI0eTEK58LMV3rOtNEigKEw7088hw0Ro3+fncGGZ0fq+pZnVV
qWIVMNuN/o14UYANLdpSzjDdnN4k1Qx7cWKk0jhxGFV7jcriV4SoVsMJfMPM1gxG/C6UIKdGZ+sk
gPhxsRAB191lhWWI56zoaWXP7N1tF166vXg2iIHaSed2cdbnLKTQtc8SEN+GoNa5pU0+VhM+VDnS
AKmNVNSmGA1RBU5q7bDt5cfYJ3QJoEVcbcpPVCLDMCu9Gl/jfEYVdm1NdG4sQcXx799dw0Je1Cok
bvZX3ddMpfb8LGTJTfqneXHQcOt6Ztw6PO0BcZe0jMMIMHVlAVRi/VFTgGSEdRIyIttEJaMe8N5O
QEz3M8JFiCY/4rUaF1wm0yqpFGyFJ6niz38jo2LbF3fERioHeulf9yKOsYsA8NOMIhxap3K8wMAh
vLLHHRa7rn4yKM4E6tz7w4rqdz5mF8ob7YUDJL4Vo6zrRxcRjU2SgFyNa+tKiTb0zfJU/N7H1T8E
wvUC2YAY/vNbUul5PhGmCYCTnCAqrUH6U6O0vhqHDOfUZQL9wfmjlecSuCocGarlDP5nbeOOvXmX
CkZ8vupK1vCy3grSwH91FMjp0+Xwf8jRd/HX8kk5cHQr+ljd9m4aNLFcNbpjAX6SN3visK7K3knc
+q3QgdpKDdX8guyZb6HoD8QDBKJdAjcAPcMevjeDWCtaRCi0azyavqdsTQsNq1RJQvWx0o90Ry+L
CU3Jcqv1GfFekB5FVGFT0WGlclHcO3zYMjoE/Zn1qQtPnS3AUpbPi+ubO4B96FLN4h79bEQ7n/Gi
qiFuUfXDH7ydy6uKNTVHKcBq18EsCzj3TCm3KNx6rYwqhbCXPzG1jJ9q4mrB7eDA9ww5l59khptN
r03g2XNeWH540fg0JaGKLqE2oaGnKS9sjDophFlL7j7Ac1WsAYdgruMrw7utqVZynR3BJZscUBgE
mPooQSXb5IptNuQpnencrjiFBJEg/ceCCLXLw1QWsmrVnMJkBmHHdh9KYgQ7Mr3faa0RUNaqVGY6
z2Z0Y9OR2xummufwFfhViPqruwlmPsTYRjEVZ2WDDn54QmGVXZxiKbaE+G5+LLPqXNbE7Tt9R4eM
ap0fakRyF5TGmsyIBqme6dv8ti+6p4W49PCSRgPpC/n0GchBpzNAXF5q4YkU4UvQw+0pdQ/+tEu6
dDrSQC7DGfQy6AzR+ACFPAYV7Q/KTXc+VkmEjtFLaaGSgzM591MvH2zZICPYncqzp0ta9cRLTIjC
4dJUbR501Je0j/rF+VAu0Fz7cz6WCCMcngn0cKuXNFN6o1KEx6CJEP+zqhzjVUQBuAfdk08GtmDC
TX8Pixb5tC+kLm7LQh3qfUe8UU2iURVOgkHkhLvzQhcGL44oJtwrn0fe+CCtHJtCyNrYSF0bPxcK
amM7ErtQndgC7m1zhCavOpqqOCZN0nEAtRTk5R09HFgBl92MmUWue0glBoYt+rLUJkdG7Ydh8QPo
rVXsgE304VfJs/oWcMsWW8zqi3xI2naaLkzzbtqeQCkWsvFiYQbX/oKeyodvIirctrKgDTKI8brV
iOZyxAv4W/Tn8rdY2VEC2Z4MmFNN70lARejrn8cMTIucQ89ovCELpW9VnWa+pUscRqF8DfCi/D6W
/LcxtUFeYHOOp8W66VhuV5fRAxZywP3RL0lwAhycIC3rI1lP6o6F5n8lOozJXX3VUULM5eH/p7Wg
ZsLfviAUOa7ual6B6qQw1XPDOzBlkT8wHpTKobj7cZgIQRsq1pHKcz4XA1wEO5JerC7vvcigxnw6
r/lDqRzg8quV9Nc5oIYtNfjSKJrKbYyBN33inqvPpOvpl2ZI2xDuoLwJaIuzr+xdy6LodxTTul+2
1tw/R6rw9hoyPjJDfIYwpYGEzX4DGccuZXEDKK1mG/qPu05GzfX88eXNW2bMgRczoNnFoIl/+G4/
gjbHFna9nuYmJPrftolDGfum5jIh2GABM2RxGDmAJwW6TJJ4hk2CiunQ0KrVjftvlzkYiWFf3FSN
QGrfH9Ux979niL9kYD2wLCwz0AEWc9bRPgLULDE=
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hFTbaYNpkbRS4ev7bDuKMYo0UcvovzDCkbLR2eH0YsTOAIicZe0HXldEOVUV1GUlW9qFI/hHAQ1b
YZg1PPlfqJuikeM76T48ySUmVOEgUjCbauVqeb2vasUOeTgQ5lFlghaVfHxlO/JlM9BArkTcw4QC
XUhKBpzkPmPsf/BvSlFXdBhNidsl0c9Ye401zZTFSRbr/NCqOtlP48jxzjNp6u9vtovp4LR+jiCy
SU9NTZyNrKOxmiXYgf33AQlIAPUVZqpIgTpNAmLFIhmX/qgSgRSCsMjep8goGfrBbdAdBEbab/ko
W6dy1luVTpctHBg2H7vM33lym4srjZkU/AC5tQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 119056)
`protect data_block
V34oiGvTYeXLXhpgWDnUTcCXtrKJVaEvZIMqWH5RwAkunK0/XP9Rw/mG/MxWpKtYtVZh9uTI0TGq
dSjlxtV/F9rycaw7QvXSrrwmaBBByxJp/ztRbq/0cghHwdE06pzYpxoVghJMUwXhftdGEu/ekiMX
SPKr7kxxsLTxXM0av9Tz2ucjKt6btv78Na+uUdp4sRYWHfl/8pL5HwVmzkMou4i8wls8pspL+mRt
r3D+raa1hNwBaQjRnvJm8Hc/3VJMSuZUpfCy5L5uyiNy2EE9xWOfuSCyq3+WUOLx+Fl4GpdaVps8
T0lkdOyQZtZ6upJMuvMjjbhsZV2ko8hzPDJO3aYgsDJwF/ynewEdiLG2yNH5b4L9nZwNxGYu2j/Z
rzRWRcxmEEhPlegiCm5DvZcWzMcj/KTgCNLcK92jsV1u27pxUc5p0dCqql36u1O7DixXb4XClzRT
c8+8BYFHd/PxDP2wteazNAlwgsZUOyXtQo5D96YryGY2B2UWpoZbeEZsafycIP7m7n8DeypAEdih
7CnFEWkxEvJ/eVEWwremWf2j366gPqI3+l2M75/YXUHi+4UnsizN14cb9HFE1lDmo9WGWM/B+Boh
sMDXGfe506YvAX4H0hpqrnJhXc2L8mb6amDu9S8Ftl+jKnl5GjuzINRt0CgwpKx8aVXX96WZrAip
Ty5Fta4rbwG+Vmfzu09WNA1IMBn+ETBaCkME+gEV9dq9R5PWyIFMf8RewDPpyARy1mXUsGskPMpH
p+7LsRrX7kydsmpXVIu7x8juSkJjsOv/Euk8zicMuImvBoHaWThZDklON2ZnOMfPdefZABSeee1A
lZGZUUsnX/ydQPJe1EXAdMAXOlpwYWD8pMfYcv9oUFnIvOeUeq1vgCH5vKUVhzfS1tdYXGkOXSlG
1vNgIzVQVSHW/9ZpRi/TmOdT7xQNyY+yQVo84Y+1gaOJ5pHkREqHzNsaKMw2tz0d/aWPyLljR/Nw
etmWszQ4ALZWgJXIeQrbS0WPXMKqF+pT9Ibh+Wl3Q1k9RN3DTm+bQSPSQnUuoRQry78aH5POKJB7
7A1IExK+JNd0oXGxmEP2IjROlitkh7KmIWnAPMKHs1mEKlUR8EXwQMCCi+SmLDGYbI3CPMu0Ha1p
SwR0FEBvOsi7kCy43++DtycZswe/QDPin45xcNB6AojClX6bRGkn82ZRquemG858ub5/xX2py/21
M1dcLBl5ekukIu+/DSQeC2Jp/ucZa7zmvEOUaj8nWyVrqhIvTMCaiVMclJc8NIIq9468zF/qRUi1
XEgIQTRBeDArmAamznj1kEe+fuyZH1PT7ADw6029+EKj4mZbGfOS+TajOfjUSdcOUJok5uCnBPXh
HnXh/eI5DG5f8eBEF/NFTPZ9n3IAlZGFzWfGpUqTibH8cWQODAE6kGkl/TXq9lVlKBQvgZUzv5la
L9O5K5Ui74uKN6YYZbJNk74XVJlclX5wYmby98nZAr+QFvfcbe/svw71NjEKaeh1JVW2wY0LB4sH
M3fy0lwxcNApoD1rHurP3x3ghgjZDyeE+EED9t1yIN7wB2kpZNix4j4otZEQYBnEv9eC+nVgEk/Y
Zk0r9jlb9V3Y4PFaXIzn+jaxk3g3SFG7qHt+3ceA1Zh6WibrsF9OkH4axYpG+V6m9+LxaREmjmC0
5eZhDH+hUe69PFHXucO2OJwFPaRQQ2EclVPWFHAczwQav1u7R62OXUW7IGhVyxcMx3tMxoAnLiFb
wGR9HgzclSSJOGSeVN+utij1FDF3AMSTL3fCigtwNBq75TIN4XoTpUIpY/LzgcaZRr8dLZ/7axyn
TzmQsX1WPREr1q0h9JxEU3o+eIiiNH+KXeL3SWH00UGHs0T4Ne9oCTqGPwFFPVXQ9YIhcD6YP71k
ADTkrjFLrbeTYxlUBEzB+HPWhVCVyy8OKihkmhnh3XdIfc5Mv5O3ULjtTCDWylNewzkIljt9vXBN
AUJy1PIIfCOtfSb9TcrfUOdCXQs9BaY9EaYJS2A3V77E7mIEE+8OVILeI65unOAMQoxJaLrr19DX
J0dD3XxRjKFauEc13+rA09Oy6oFbHh9orfoefEgZaN5OKArH9azIZ4SIlfLjOMcFto5hKy4BR4YH
BkJnrIWga2lyly79dUbfxi1cLM9Yo7l7YZivti4oQ2tAY5DT87aOFRFfgyPjrOVQWTP2H9tKWRt7
4HNDmcL70oouNmocEZgQceMvf6JcPFxHuHUvM5OrzhAzDB2YSwQwY+/BsuGD10xgZFv1jMIiex0a
fSF/XBhhGNrg8l583FAR2OL/ZtEcNKuF7WsEwMxS58c7FtLtvUVYVxooLCPmT6lye08px42Cagaa
wR8WPYmA+GcHIa097fFzwMp/V+g4GPZMJltuYDJYtTnri9XFvUd116QMRnN+WmsPTou0aZiYayzs
650D3/WyVOGXeKmDGWondc3YkR5B1Yj6hgHdGUxmDgtF5YWElpd3J/Mzrjk7RU/DXGrV1v7bSUBN
OpWzfJVACAKW4ZnPl8E+F4ka8qInTtHyJ+QUQIKIapR+hwT958SXugICiT65ri9f27qmXjy4xhx7
9cBbI3fSqPwMBzXzt4sdVbdzPWxVTUYCdCCYWHglPVe8hLHC3SXz8l4dvlPav8Mr6JTDv32fBKY+
1Y3091rw+PUvsi6NyAUksiCaoTc3x870qztOg6WiBurGWPpFz9bDtv23r9RROCr1AS6vUkpOq+ih
vN5tdXnkrGQPhVP2uUOHcLHjtGWKPCLsSpQw+pb2IIbs7ZEKOiEEitVg+kbfpWiivnweLYkIuQIe
f/6HRw0EIhueA2QZTDLB9VaeayeO9iROcC6S582+BnLe1T04X7xohZ/Lhye/r9ypwwgfG6tgQqwr
CVkDX+5g42qf9mkvMF/kh9NdOpABw3YpuMQbOY0Gp4o+zPHozQxtG4tAfaXO0mMkmB2k4i2ftYPr
vfLW9Xqp6DVU828VnKZWHePsTyebvsLVQDazzlig7he6lNuOEJRUCN+Ox0nYxn1Pln+K8hEO1qL2
TwH+vd7H07YS9x1mEIWc5DE0it29zSLrFtjFIi2XROsUQSRU728C88y6H8807/VX/owe1Wm5yuLY
zGvvDo/EOsIBr6lQHAb6+ri0x4Cji3oZVl9NEi+29wkdy36pXJ0zp2dsonFsodLgi93YVAYg2ZEV
EEdDU5lbvu6Y5QaQTakUwRn9gQ4O71EWmnnpW841i+8XvxuRTPcyAVjsx+I3K0NSWGPlUwOQcwc7
CknuBo1Tpo1joDs8Of1kbc/MtyPv+QNaJ20+80K8jJvDTUllRDf9oOoerSRBjX7ibUrdQ16f0Gnv
57z7LjoSehOgWPgmqLqWljt9jkuDRfu8Dbhx8+Fb5rUwKSf3Dqb95bdIuFE+E/LBzIDz/zB96bdj
auA9OUEnIUaq2RO4Jdv+FSOx7BT4nayQdRauUu+qghy9lu1JdXIqnl2h2NjWYejNRawGrGDvFEOw
4fnoH74scEKbquPt3wyvBqX3oN87vRHwc0iZ6WM3t652vbCtNOHdvL9NY1AHsd0iqcoeDIM5Iv30
U8ja0ZhBzOQYB+Jaab8SVuMmdD1poOkY/m/2dyxfychtZQ6hrI9dqmota2T9e3Do1V7lKMYVA+dg
M8SAupL4ffgvyqzy4Tl4ZLJxicRR+rhR81Uy33yjNPKECBcUpsjCNLQowI9SWuwqCubS0aRs0mot
zUwhsmaJ4zqT/pTF/keBeeDwHjkIxV36QQIIv+suaaFfAQ+5pty6998jER/B3yrBAib3hFwQi/jG
0Pxwco5kxCap/mF+UAuG03VqYqf4HEt0A8zhe6FnXfbhTCCB5Jmbg7G/34PIPBub4WmF5jELuE9s
ukoYaR4NdydtI2/OvgAnPUrOOYF5WD+53xe4ePDdtDyPxeet/4Vat4zTV1s5iY5Q5svLg631gEQZ
KnWsVsAGDCF/aWWcNqeXVuPXlxjmE08P6WCJiUZC3wrnNbGc5xyAIdsU5o+OT+iipsWPaZunJKDm
vHcr/CoRkIFtCjFbAPQjNygjzzO69sMmrexKsdn51XYPlNFYY+UPvTZ+/hHCO2bi6vTNXXNGa+sK
GQ+3A0uAtGlHV9w0/ADULqaZY9bLdL26Wt4PRqwmdQ8c/uRZYIZvbfJnDwX87zScD/dskVefJ3R+
ko6aqRWpczEs076zIM/mCLXOghuLiDxqtrXQGyTDv5/wNZGQxGxHdlCzCb9ik4M2P4CcFWQwCzso
QYGBvzuJ1fF6Q0Fio9on0Q4XL9sby+KSVuBvDuxiwpSbIxyKj/4dIg5LXOz66WQ3w7OEpAVY2aeg
PaiMBdvieTGmrhGbdSba2heiSuU10SIkZmf3xxKoTkrAMpaJ9LHKjeWpQcUqHm/5VdII2cfj+u3w
gnykClAska9FpwVXsqP2pUjAyfvJcSzIMLWu0430AFsZRPelaNA02muIwGCoL3v/58KbsdgUkvQa
h1bx1QIqZJ8IYqm1pSAuEJkSwZMi8Y02p8X54MwJoj9jekQnngMhL/cgpi82H31CYcfo7Wi/RRdG
AD8yiZO2SOQUevjjzFvvaioMUHSi+E/VmJ+5s8SWfUxjKC6i3w0gbwappa8pn+Pc9ezMEXZ7NeGl
aOd3W4NKkwb/Ww5LPXzNVhEw/b4c3TxTe2vkLcqxAWJCSY4H9TUK+Ay/hkIxOVFKxxAhJH/z8xIJ
yd3lUa8JYGlyIuusZEyRnKEqfROly7d7kgJY+yNL/csibuHG+izbyNZb7w6T+fvuiwyixaQZejOV
qmPPrYw9biCwxxJ6tzC1ZW/Blpl1NTUziSSTElZNwRx9ywOaZbTxX2hMneD+eZedyHlqsKIjwgTh
D5DnvJesMpqaY7QfrdKHfqFIaAZGy4/eXv+5cBt6MMHUB8K56zMETMe6AN3lxC8HYYaRJHLWn4H+
4HOWt0eF2loMUQSt60o9R3DqlKEsBuMrWmayHBfajAtBVi9CbBJ7g1OWOHf79M6zaRlsxXiLrDcv
XcDQ5QrFiajKAUw8R8tjpvP8kuXcS8fbBw52eoTCgaVNKvrCeWfxF9Ze1Ants2M1FLBocGefW4N5
jjRbeD568yW73/+lc/g6oENInimp2lyXzWKtxcbo5J0CErT4XXyzCWQ1fwSLlsXyhPiGd1vYDIMg
9rD8C2cMu+lgh2HRFNDWJ2lyyzltb81KR40/0LoNxJXKwfMvP/vWxqHCxQO7HflL608pXGbszXRo
wbTDHVKGk4bVC6hErOiR2b76eRa3XWqslc1byt8kms8IoUfAjx5jE4ULqeTljmpk/z1loXdpoe+6
4gG3MG8QTPBb9vkeC9b5M+/6khqTy3neQ87lMeysdBu+kcPUDhcuHaX2k4sPMDaxFvB5NKOLhKJi
jxE5ztk0XHgFA2indY0EizLFe+MIDB6o16DSnB4gi3juJWF/j0jnFLv7SC2RbNsJ3Zs3uLSxTogJ
C/WjW5DKqHAVoDD5nUlnaVhmxZHXrlw+yyXBJwOZixCm4KEhON9cuIat30dMAeSK2SAxW0clvXT5
6/9mQSo2uj2wOEeLQSP2etwujpMvyZDrPZk1UX0a/ESnHydG8EqODXmAITCSesj0eEgsQV9QVmAx
OBseStAVQ36w7bb6dQcT6Z75W0zye3MNTVw61ZOPOTip8dF/zA3e6LPXZza7damxlJ3N+rlcURKw
6xtesPFdZ88hihvZkidvXpKITYWsLDM3TWQD5ZZeJJMPoWOQxTYB1CDaLEPRKZ4zCt8pEAMjaZaz
WvS+y6vgmaz79jpEM4kEc11EPvEgMgqR/MJM8auE0wCsl/4uR5LziI4Qo0vk0st4VZqxod5A62Qs
QzlC1W3OACzUhYkYVmma5o9ewwpBM9jQrIPxtScpiJinBQfWXDfKZWa10k1jwNeLHJrX6Cs6A5sy
FfMaA7aPA3WS/SWno5QaI3INIr5Y3864JTev7PT3VvIhE6YJyIzkQxdNK3fVZ4cC5djlggYWm85m
pUGEeui0RFaml8ob8rzK51Vboz+99Dde0V7nGmAvVU9A3J/3t3806+vAKSJ7kVEN8Geooj0H1Fes
b2+8PncSXsWoH8P9ev7LTsQDSaU1RuReeqquAZMBAb7esaBnVKBgQLJjtiRmoA1Z8tN8RS4jeOlE
gbWB6Gzwtc34EFjQrlz7quwoVSDeq2mVzooWU4cTjvOWbAkf3U5w6ILrMTy//Ka+E47tSwLGC4r4
Zusm6CWbWhmgm592Ic+vPGIfsfZwPrOCattO9j8w4emBSfBiGGJYu3CDXgllckelQ2JYNwKYGBI4
rwtDVldTpPQcWsyCtad6/1jdJoFNJgaNlIqkUi24080iYORzfRnpKCLbKr4JWoyunFFEjMNzMB8j
ZSVnUrhswP22sD/XIJuVuIYeNYC5XCugKDRFhdyYbnQy952ShVh65/gcaAj1zPQZV34o5Kild3lm
UDx1GQJzzdNx/k5bYS1HEtlUDVzL1NMGrqY01ufOOlDF+JHSZiNi5rT+XlIxdYsa5aLBx/fwodzS
nzL2CD7Z1pxkJ9VZNDbvkEOopj2OTDEfNwH+8zsRLnOGLVK49/WIrCNqZj8OUVsMLPyJAdpJsTE5
xPT0lOnIDcGjfRvMQlpLF5W8C9GO7vo2vdr4S5GMATbBS/B5oP0zFWBj+lbFnoZ60B05B7OGdrwy
fRHiDKmNhYd5kD7+vymvA9bUMR76JunbFfhsR/luPm/Yq8IlGWmqpcm7/mtljFwtaJAYRMeupcfX
IuaTi+1HNwd552Z2N1YvLARjBiMFztFBWdp4IrN1w26bydKDHjwnThKNPy3Jd8Z4ltBGOptfIqpP
ZGVPcX0Nabzaa2XxW6hUhA/GG/EwI/0rTnlrmCmRgXsW+/nYLUKz0h7vmATtT7A4wX2NoG6s9EHo
3k0uf5bd/gEg3bwKNx8Ih50zy74d6rH/BxKP3qLsR16ivpFn79zLzGsoGfUyMIYSJ2J1pyDkXDPd
TrJS57xFfjQ1lAAxbAtr2DZ4lYjrxPDqN3CBiNBrn5M2iF0vZw/1/E+nBzsNkDhl3zCBVWEbpz3t
AsCIAuOH74jvlsxVyQgWkweOiOEYSELTogkjVMSm5k7a0XFFdHYBNCtNBCj+nS9RLDQOANkxnOrG
V/+c2SofJqf0+NG7tpGwVrcGHXIkXAD3kfh9Ndb/dlb58Vbidtz9i82FK5W9C3PXV05yInBBP6Kh
mIuBvdTp3G7iSGFJw0fFLGczTHKmqelo/F4gmarW+yvtbtmN6wcSDlSJ2TGOKlMLeR+W8ZIXJnU7
SZzP6fyrOvveIme16R+NrApXAUUz8AmcFPIjtJ8+4Ed+G8T4v0+9jZ6/cJcnLVgoVym2wEkCJDe6
ka99cZP4TDv8/ms8Z6mD7/awVmZVQB5LLaVGrmNljhg5BrrDESNGeevulUzFrnIZRO2LwBEklpKO
Xskx/nDsqKcRWEKab3Py3capYs3r3/Ml0A4yIkB3o69gUR/Q9iVr/O1A1Qv/NX/ydqikB4KGq3Qz
ANjW4st4rv1uDbgu3bNiu6EfdK8jWdUHw9cJyzsJ/i0AzkvLzTQpOozhZVHLTXti1NJTwb+RYHPp
UrGgdlKobT9v2adlscJYCO1GhBOoGPY5c9Ghb1BAmLx5KEXvZgox6gmIncJUtKg9mf1Wt53kibIw
3CXTARCMzSgEUmL4NmuXQ+Di4b+rG9O9+Y/dH5E+ritTS9cUvmpt0NMIARQquOY8qop/Ri0R3g4+
L8q4l8Fs82uvUYOUWZR3kSzCLHFJgM7fGBhmdja0ErhKtJex1EeaXv27DImvTFIzBTGf/OVKDm8n
u/vrZRuQX2Ikr51OAlQ5ZpNIXTPSV6UNgLSUhjKxvYtnV7600hdR+QrQ9NwaCkq9i0yAi23gCa7m
9YcJf0AEKfAITMgJdO9DxCWdwVgVvIARAgx1F4KBhQhGywS9SMwpfQlrrMk2DVswL42nbhJTH+7L
sjp2pAn+WjTpho6hqBldX366PZTPhJPS6FtFWyLIiHtVHW/RX+WSUIGmb8UQbYmk3txTS25b+5DX
k92oOVPTR2Q3wIPayJQ8eXciaUcSnSmO411Pw1gM/ZOR0h0PIl4n04OFKpStH3bQRvQiGZo59TKl
MBYBtE790f0ueX6DK5lihwqmRfuT2kYkXFSvPzqjj6vXPFn58sMqFT8tpJgqbsYTLAc2dBBvPuim
CAAiHvahGMlyaSIPrOoJnwZl+MnKBovhOFR41No1moOfOTVcW2Ka5XQ5byMV1t4/fmBJW+/7hv4d
mid92+LYGMJybm7YcN+3TtdHdGONzjYSpCJpqZzJSwlU3RlXTM4szbqoVZaZpMxAX/Kpc7DL0E/U
2G/NKuPzFC4NcOootod9mK2K8Gcvpvhobj1BIuQkkTi/iCbzQ9FtBzVofpkRTMcbasDgb4XExthX
/vPj/rNz1qmqIi6x2wkDLja3IiVKNr8Enul2kn3d1N3X3VHu4Vnz2N8v+ZSH4Td9OMm5vjN2+K3Z
U3xkXS8OFr4Z0C5muSeJF2EL96mMEcv695U+vd3JceESBcDcsXaRDSGe25imr7Gy1TCD56wcPnai
9FuVbR0D/+fBvPUsoTft3+9+xp2XY+DyA+05YGiP+GjMbbSlZLvoHwTgLIpWq9LGpmqRHnmvne3p
wkvZGmCBWrdd7hQhHopCxuAGChoFGbNXAHI+4lvTel86+6PFvb8O3qXzNYKAmFnW1ymiz93MIYsx
dHi3b0Gsr12Sk6sQugYGsyli6hqXJeW7dpU+C4s2WKhVGLCGRqKBaCqyKqTjFXh3eNJ7KL3yGNFw
JyLeB8qdMsEtt19Z+d41Kz8+kTDSuZdxTK3Ujvp25gyZ4o0yUR4d4u4Anyd93P3gi9k1Vpdhd6FW
IAoEQCv6Kh6uq+pHDyDlCak15DlFVzXtN0eJgltFR5y2beDBvFjqQSlkMwk6rNSgdCkbRaL4VuqY
1ikTRU4A+M3dlVvm5oPhRRAaQSIUsduZ0aKyB9IJWwQTXEgRH5rM5khg1lvICEj6dj7vPq61yEaY
ci5GEJzOrxzkyz75ham53kcy5Bi+GduEYQMzyvG2mCzc7fRjpsomyLV5fwu8MMhJWXXCFQ5ZcGDG
ZvgWznToR0GqKl30Ze5LozUutbfAiVtKw5jsfElfcdoeO4wO55Yfkz/wlnLLGRkbVnsln+NUAhgn
JPL8S5BTYwLqDDNmRfqofz7aoX/bkgRkcvavYhfJH4GoHgKO5fi6uCeeeMtCjl5+U0K09qLJe0BE
Xj6kb7zaxtR9r9vAWRK4l/Kjsw38LlAZrSuRzfUqA9Vcy7rOkAmgN9+2ceijrYPdYrIBOenFowNv
g0nnkcSoqOSXGkZBBETzyy0Z959wgbSC1c0semgOEPzY/71HwRu6SWtIx7Cy2JRSAF8byQoUkK8r
9sOn+BemI+pa/CCnlAhrzM50z8FsqDYjWreHltb6AecxQsU2bPVs5ELdv/LZUlR71nXCHe4YXnPd
M1mSSpDDRvYjYAcEf+tKVoSR8LD+NP13jlLEr5ByxaM6+aG1yZvFtm7C84YQCewcAKOwtS8lo+tv
KO+m8IH75Xp8oovROPQ/i0r9QRTFS8kTQ5mRNVUDkv5LrE8OSx4kr6xEL0VefRPPIM4d9+LqIvyT
79bDRvEzH6vZp6k9OCd66KHORQqmxZP4qPE24tyu33RkYuRzJOZDq6YesJVA5/MrkTjTiMskQumz
TmlxQlfWI50C8AUoDty3t1eTmi83u0jYxTKW6xx0c4XFIJ/alFbyN+LviH4ReaU388W/MdjNalVE
D3rNs50gfo1iLRCeSV6HaIE74CDu5Y6lKd7NRiewkIQW3IshCnOVUgolaOxueYIGsvnNTGSyXEqP
HSRTgjsJxmegCqFpQVI+EtORI+0vVDsINoLKxe9k+Pt8y+r+Z5aBLkTRSomHXIbG+7jniunEbqO+
pf9ai4YK/EsV+OhhdCW3rKycB4sHlprIPkrGh+9xpQP2bfyA3Z3InDwq4M5gFQtwcwixVOjRRZ5X
GnISgpn0Znv6Pp/6WDko/a1vDpNZChgL/ERq6MrfIYRWzL837P7gGvduuk3fWG0jjcSVdZKXP/gX
udEDRRZWPIos4/Omh+0Yq8sbEZe8ful1enkScdOwUOI1adnczJIekOlI8DoSLQM+q0geAl5vMleP
x4NjvhWj/PaDK+cES8yBngaXOWxmFoHkt3isDK/RYyv+4mwJvk++ifNb5yWwkDNg8AFaeVjxJMD0
6vAiGxXBhaDXP6099QBugJ4HJIB0VIZOnW6YqpER3jAH9oW6+aDFcnbKpIk5fL0Z29vq/g08q110
pAKFc7FdofUwnyH9R/cp3xpQ3EXSFHRNq2zMzuHaQZXYGT1WboaYwgfw4Djuztu1j7Cg7Rc1jUAp
hzL+HQ4bo3c5MoqYonwZ0MazHI4s/iwI5Uke3vifz27NHneIhDTIAbapdtwzRCcJh1tw9fc36L/7
vtjBXRbUCuLruBfYLqwbCs0TaYH5N+VNo8baY5wanEYWV474sWnvxB48dLTZhlzFllTqzsSPx51I
5ENGoRhksq7eoq6c24TwP8sjfU4RgKkW7Cs98rl0Pw24PLjkMgFyCwbcbwkxfI6zpBOSlLyli1DX
5DA7nDVbKLfEufFYRm0x4DxZWYd8d4lduVVlWS3oMjAxrKvuq4/cJHJ1SsTKZ9bVcw44D1SkRNHG
6ucy2Py3f/lFvPOByzo2zPw5T/p0Nih+NXY3dOCI+zirdD00rdG3nP36NmJ/nfnRqBccBJkrzN6B
bBy5qCCrGr6IOxrXyzb0jHNZpAjJlD5OzEV90cfHRC6Q1HcLI6qmr4dWeMJQgdT5XR9+pNuXPUWo
liYd+pUHwlMSDX4I1Iv1kv3kl/sr2nI9cDjVNw6apJCVo79bifySNMOB1KA2+BoGfbTz/gjyPDef
LBZz3vDNziAMs9j28qXNa6jlQ+0X+iaU82FUCexFExJ9LfwqyZfPMxhgJUCEEqkiQhXZzxBdX8kM
GzK1/5wsdf0SwKwB9pe/vKvNm7r2e+8K/9BSbKjSSMEp5yivU4hsAAj46kPlJ6PidtpDAVQWMo/h
MVnDvE9s7t9B8f0nIp+2mHyKZm6d7jULfJE3UqvvqpBNkZ3F1rI3FoOuZSPDiOnzsgxUOIaxAuEO
F+cqtD/XYki9DFZ82PMIlDng2G9zxNAubefHHRjKMbtre6pBBjXKt52m35WI7qhHXYHClgCcWqyO
GPfaNX2/nLTs8nfdhQncyLWEiotAXSEi2MhwK2SWoCZD07Db0qlYfGofL0CXIpVyNTdnBxHcGfuE
kjV2iEsHQVt2sU2dZseKkwQ43x4PHw8J2OgK6uOeaIc84PLBvwXch7nvT4EE5MDBmQhM07uHgMvE
XLWyPEyMAWZAKPcI20Uoo2Q+1Y9NsjtuS64uEWkqbk78GAcYE42Gfvxr5adgcEvNfw3QpBVkLQcu
sAd7r90yRZtpYxaDEnieuIa5JgY/bjYhU4CaukfjMXRe4LgjgBylpATWcHg3yEywutC2YPxVBIXZ
2jQ7/f1+u++jU1BioV9qAuccBae6ThRpHZmlpjKHJpOR4JIrF6w8hxTzVXPwfVkKRWYI3ioR/GX4
z9mn/1bWuIXIrItyddjFiQ4T39+CLviZikOecynG4S6KQwpJOJf4rU5Q86C9aB2b3IlEScMxfMNp
nX7+gSTarE8WP7UudvjoE06r+L3RWrkunORoeDhDlDXSmGWh8w/mYEc1lZ7oN4LzlkMK98l/ev9P
uzN6Zbil2ruKCOzxWsHljhWZsBq4aTMUM0chLWJtEafYPBBVvveontEBqfwaYKLlEinE0LaDfLsg
fmB7IAMwalJes5nEecsSX1b4n99f4PUuuXmcgLPMI8zuVEnb9FIDvsAHLQBbniRbM5bRw5pT5UJ3
fxl4zmpGu1E9el3bCXKjuCFg0mASbojadq60y36KNP9yDjMFYD+lUhTTDT03RCHKAtsPx1DMGb2D
cb8E/g4dvmRiaQzX12LA9TtH5Xjv4D5Kq16MiNacjEVPjJd/1Fn9yRaiPMPkpQn6xNX23v2f8OcU
Tu17dKGpv0qes5Pkc9w79Up5sCeAqkB1cD5oSabYteZdfD3t2ZCZtX5DgQ7AP/G66755nBqT+3WC
ENBlm1IvCPo4qMSGKS4ZrcHOXJvWhYdS1B5o26PJ3FxmQUk+Jih7Fl7nyBqcvR5yt5hK4W2kS10o
5tfcwSXjS4Xx4YNTYmcBD1oQz57njFgEewBVVE7mX1Yeoi3DPUsNcZ9yD/mh1tpHzVqPG8+U5idk
k57O9jBAeNru52hE31cbdEkbJtrr/vLovbonPF9z0f3w0AAo7KC3201azXBUvrwE2pTP0fOI1rPz
kSdjF35Pk0ibPmREUylaaiiRXw1b9z+xUcrCnsb9N4FoM0ZwriM7ASKSDSY+h4LBfbMeeT0vB9P0
31WUMJL3skz1LgynfKU0LvCG/3ydgqJ9a+2uxlepk0HXrS4hMA4lpZZgtFZ/pdpCXD9qG97C8+oN
JSl7nKEfzl/cg54d86EDFUNMu0fSWsg2jLkpBBmgiqZEykTfEbqMEolq+obn2ktYb7FYlBBosl85
VrRz5YvuUGfniEEF2d63nysXjTfnX6IrlvPhGab885bIFjc6lFctQaDwWvD590B0LQNEoTH+Umgn
814Omq5z4DIt4Vxmx2RkyP8cifGL1MoFSJd55JITRRZ/mLqL0NRfuyBAvU0+QgUIIWiXXb8W8z/q
3awhCG4m6OGefE2dDMhQuMSbcK81nL3eTu9P/euUvurKbxzoDrDCqWKw+cJ0oVYWix1+0aZ+KQFB
7W4KpeoPC4X9aP8Uz799svDkiQxEiRwnbeJVK8KYiWw1YPiHFk9KKmg4f87wljJmRt4fC2A2U3ew
t+fxyur1q9PNzUwKQiAJXwGRgRb5T1QPZsv5N0WEm3IjVtJusM/nVvZhI94dL0iYXWvg6ZJ1xp3M
+/LJbjCRvpwQ6GrA8SzIp5X4zxvNNvZOcWC+qRvNOkhLeWsFpGiMpnPlxPCYaTtQHRnrtPdEGtuz
umvaFP+csqsx2VRcC8JTZcLYjVc4FNGUz1ICJTB8YXK9Djw6Vgk6eAxBFVrSsS39o8ZavcUr8CIj
cznkDgTuEPKNNLR9lR4yRF0DygyYZJZaa8YUHuOKhVjIm6/WrmivAjVO/Dwnidpag9PYuCIJ4G/K
20nsDvhJ5qKJWU0ZpywHuX+dYDYtp+SbeYoaK98eX0Zk2d5Ph0Lz9fsbnyukNLtSkTnd/7LXU92v
kd4yzCxmqmSzy2KQvrIDvvRZyat3ZyeLOZ+74vLtQHoPwLn9M1JWcBNheC0+3eiUfE0w4aXNt6En
/pRYfHUVMSymHcU8elmWVW7I3hHIX3vV+jJNx22CuSaRRd47K8N3I+lccwjMLl+IJAtbiInSgt+N
flaGDkwgnG2YwD4XSmxltrJBY54cnoM2KDlbUAZdqPUmp44YLnzmgg/ZO7QQn84SaxeKiUigC9ii
M5C6lXbXbvSOCgHOdedEuC4IpxkHwFWGJ8VLMP8AbgkqrPaWuHaXRDIft3nnb+DsgwoISweFZUl2
IDYLzuufoC4FY7mAMvu0yqSZJd8wPkINP8uCY3+HM4GQzUbnPAd2pzP+dE/p/tXdfUi/FnCJ8ESx
QFiQkVPd7XzKUt6kUORNavwX3lD5D5G4jXKgh7tkcIc+HgB/DNBPFPd4/Pj76/86b8D8T0qRZIZp
4eC0y5Ljit2MsgAGpp/gb/C/cDjt3B0W67/PuH477S0mQyfzdb8VGpv3VRbCwU/UFAn0FTvjmGvX
4caK2V3dFKgmU/ib6ZM2H/V2QwbvGC97dzUdGg2mM9UwToePb/Tr2fL5MonhAugsjjo1QkM2YbCW
XM2q1lTPrCpUDS4pMVbHPBbcNOHweqOVvkFbA+jZU8DMi019m7paXVMobKS1YEE7XLhL6s3zGvdo
d5amJ8a7+9y+iW1IHBWkKSwVfRVMVQvMQMDwYLlMCW91Eeg18kb27DIk26RUwW7AJQBEIF1k8xhK
4U2iZN+z5+Gjgy9rjQLtBosHy+/x+fgmV72OA1m0UG7rQ3i0c/maCwqX3q4rcXwWQFpjdcPd+pJx
kLHyo+9CNOtRpsKRxIEO4Jpu9msClBfGXt84V7Kn7p/tcKgo59LiDpM+zF/wEjexg03E10d0VzlE
Qi7+ynBQB/zI/jUHaGcxc4QN+KKeOcwfLaX4Mv4TgN3lFbpSBxfh2uXZq747eNTczkEgZLJ938k1
eKtAQ8uXYffk4tFKUsefUvA5iTIIyZxxuaOcoQTTr72HAoTA8bjwVDLS3lZJrNmi3Mk5wzDJuSWA
i277vVDZOE7csLnNqHTzYPqEQt+x60RlOwMLoGd6RxIwP5EmLc+yrLVqsCOm3JO9/yI9STJpZtqC
AtgAitc2qGytqnKTq2hHDPo5qHhYokw5IgXravpn96R5RRH4aKRb/BsHedV3SpBNrOHl6V+QI9/j
HBAtJ8KquyRkYZZNYw1xH7nGZ341Z744DZ2vcZiXXOVHJsLXWR5AEhR43SbMNZcPhiHOKUzq9hau
UndOEb8mSoV7bJdkN5Gf3uthh2PEC/+8h/bnz9l85HSVtyFXBF3J7A9l2VmcJBxxBY2P5AIhvDdd
aAB0VmEoXPKIFCCeOlAZgemfhZwCeMKXbX6gGRuJpSR1RWmRdbS8RMY7dV1YtmlreY/j5vcsb+1/
5u2eC+1EYH9DUC3l3/qQRJ7B6gklgk+Q0PZ4Kv7ZJNKFW+US+O+bGwfcPtdcs+IgLwvwWqFNLZ6+
F+DteoW5NtCNpOGhq5pzhYv36bEQ34GL369GE9ZTOGiz3GC1EIKYmvpPGUDcUYxYDNcEXBOSNLLW
bAD3PzNbYobmQawUUBxUeY7asNIJIEaN6lTL/gl2eUQqAZfreWMD3bUCzK7IFp56+hT14K2gvz5O
6yPSy72J9VPPdNP/NYU9ieZxFMzEqgTOD/YzqDiTMBCU9eAXSMMUD8f0qlP1Gfadc0+BR6dkvFXF
3BaLn7ZQyNICsrbXqq2oW+C23h44NDESVDTx9mGUswA/u1FgpxrA3jVjBw7UaJyeLOVKsyKvqkQg
Tw8kagDzosw0mnK8J+ADwUbx7MyemNcZUKKmEzBCHQSGF4oHTPcd/26QcWyPsZfa2WhvI+51yjX/
STAHPczAkqHewim9KGYEeQC/1rYgpn1A0dux7/NZibqyeIAwHbLV7WjrKCpRo1RUoy8NXdEeOmyQ
M04ew2TkywQhzoLHMpRxFLC/YThSWfVeOD2Xj9ltRpaJimjx/P1KiQTP243MEHGLb9t/7Hv0Bp3Y
Pm3bcmqCKFlhI2x0usMaD2oWHKt2ryZSuGLz6cDssxs3TkFeopEwQx2RX+I/FBD/Dark46vxyNBx
mZKN9eeOqfEOZsppEUZn6MEk2wp+IX4fDoEV5MFtUs+8XZdLdlT1tP2m9CHhYY2MEiX/V4JDT/oQ
8I53afs4Mcf+b6c+Lhj6qgR4rgQYRmAiEBmojWqHCLT2w7V8+Yl8ani8g44/mOYck5apdLvGse7V
xhhPuR4MB1dTI3ZNDCLUmWn5X6QLF0D7NZ1PNqw5779qErHFRTKbES5edhFRN6lp9ZlI/WO1qLkE
M4niWldYes7h3tgaHbTVHkJz4fLlfBelVsa0nYczIO6gTFFNb8ICRCkF2w/3Z0+hCV9XbvizSwI/
9djSNVdqT7BAFUIJPdfFOv54pC8kS7KDKTlJJtS/YtJ35MImjgXiMNfrkfvn+VibwwVfxyBISSiY
NIbm8lvbzv+n9pNueDAmgD12j6YBiM2jvClSxwUbm0I4qpaBSHx66W1P6iEG9XaG58KEmYUhUqAD
72JS3NuHyiA8B5uHdSTniO5X+12pT0dsAknuXPip+kjyxyQVnLup1vmTpvS3RY84oP3uxPvbyDim
oxsX2QwFTFExLA17hmZ6ABGmjTFSCq7h4fR4LdeUK2PbelJ+2WhwiJ1osqczMeSKclov1YHY4mf+
ZMWeabSBsGTB0MniWJPb7GDD1f7gE6GvAMFQNLDcfWay722tMl2D39QuFbhgTOwj+z3j7D1RyW/w
bvE1cjtGxNSNnWbuJHf5nf9I897P4vSHyy1zafFktLgQEJZJPAXiQZ57JPXTLQpuI2NDhrWaya7+
Iugox/lgwUIHIouIoyqdD8zG2JkHPKxmHLLgWhFwMEmDnTkNNZcpmJMgf3SfrwtBYveVoUpZeOze
IxtNhkucjTsxZEoprxGEKIrRhUAenBnojhvJL384ZnaWDqtrbWXWVyi21VQ3PZVgO0oEcAfCB61p
FQ1j1I8KBrg78ObTMQYveu0FYbg9ZvBAscI+9NXyG6BnnCM+IKoNAvYW/206gXMwsaEnO4r13Zwf
gyeyCz8ZzpGNDK0jASJrZwq5DzwT5/XIhBLmxbPf7D0ErhW6fMiqXNpmdq9Oaao6cFYdebtJBQla
VFuyrwnhfUnKKkgHLsujhYMv5ctwrsJ2LBVXJjQ5x12gkJhHN7faWR7Z96mJCKwoNJratOb4wjiW
C607lbQVcGR7os6bBxCx6sd/7ZpOOgZsWC7TmrYbvAkkBjtIWxmL4ei2qlCd2khDxrolQyf+9ftZ
VCcGDJu2/Dkk2Ex38UsqBaBJ3VAfo6lP9DaQBc2NcJf76nWoJ6TQl/yi1G+SB0dBn+/NjE3cIfXK
aLaSF2rbOUbR7VHKVP5ymrp6q/J6nj7gyWGgBD+ddJPPD9efbuwt8vyycUT89034Ay89G8AIk5Qm
kAUoFsIX5sBIN2H3dpfMpdQprXru7J8X/CfQMECqd6WvxJOZgkmK/IOK7CXMM2Tg4r7MVsYJjrW+
mSweDREBaiz2uFsimW+fRmkhzr9z1Aql7m7LYfLL3YMDTAeEZij6IIUUh5UHwhEBGZf9SZFM8fVL
quTciHB9WWywEuCZF2Z4kiCDjFgAA8KLOTWfzNd7PDvjklc2kwhr66EN0SF/4K+BwzCl8Yh2yUwB
nKUdqOidzB48nwI3CH/Nfgs4JKYuaSqhy00hYY7nxcwn5IGbeBjZQDEHjwEXZtTm5AKD1m9JxJf1
DPSrZno/QZUockDO2LwOPDXrdxAMz1RgjCtlAMUiJtLhZGKPI2T6N8rwRL+oX+JtTvLRVwXyC0EU
2yuf30gpYgXlvab0laaUNqt/laGhoFd0kq5IM+rv/ssR6LxTpPMiMRtLXC+0k1QyVae7TLVqzHMG
ZMPUqYO9WHWLg+OHwkQCGVzvk5+U2liWbLKrS04OzEFnW6k5GzVOFsX+q7KWyePl1YHQXsEibZ13
34j/+AKgoSkF8b3nvWEQvsx4Mso7jrpm1YPhxHJakYlmb5v+EOoQRlXLiE9JKP7BhYkHIe7u0ox2
E8v/rdY8W4PZc+vzZB2tw4q6+MlvwU9OoKeFQe1l56+kyRfeJTC6DK7WVYvU1Idl8ZqI+pejm7sE
DrJQ7tZ8tGpGKjD5uNp9viqJdI2Q9I0zhXyFSebhkFZdiyvU0cCv5h97gk519y8xyUqurMLv/y97
6GtmmBJYmKZpQHEDWfrxYR/0Ip7Wc/hmmD3lsNt90x6x5eiaQf8gz9t3Xb0Dc57BsKIbg63S/bJI
xbxk0BY49crsmjtEBGIFWrcftoSWWKtbb+MQp1PNEZO9pwJ3Ct6T4s4bmY6WDNwhKKEMkIsTIJhm
vFDN+50q4WdqARjbK510AkfzJywcq1GG+BhA//WsiQLsUi7FwPbZIKQ7NPWfqiTaKBa4gnAunomw
Oa7dZtT0iNt96sLgg8oP6gKYaF8mfqluDWQGwU7S0Kx1H4GDEoTmYyrTcxwscWygpuztZpwAiRcn
vn1hMmXvj1fcxTkEmnUzIB9QMXE1vzFwO1OtOauhRujBSMVsoksTtefJA7UQZwvkH064cCXWXdE4
wdD2dK+oUgdoYIUD/vs2zeGDIkHT2M36aJKg/KmdRFEPDKDQhyND9DTGTsv/BoRMkt+6VSQFuSsf
soXZ+as3eZqCPrXafseyv3F4iLhWjgm714txEsYZJNXpULFUbV8mD27ivU0K36VJLDYBUOBuUgv2
KtM4QkJUygJrVLMmfw4yDtKKcz3ypxZuZkI8FcXrCxM2gEYibzEPS9Ye0dnJUw5CRAnAVmBNbKGv
uhPNsyA/4tJI4o2SWp6tjHp2p+pMGrCagzK2NEKk5Tn9zZuZSNa+oXlUrjSrvI6g6Qv88Z5tah95
BJ7Li3K+JsWj5i8zBsn4RGAYtn+vGZ3I7gVuWpRXWL/P194BMpa/MoTOqNBiPSVkh4UiB5d5hk4R
5Hb8t6X7nSFBJbD5vXw3vidwXL9X945L+B4KdFPnpkl2CdfNWv1r/KH+Gy5coYDPD1wNFOaNe8JQ
jsAx0l29fxADWO9xoNmK8X5k7qxDstdez7yAvQgX4jNBlkoSvEkrY1D6HujL+Itly1KQyMkvUU34
ZDMdo2eUy11POlvtyKGyVeDQ+YAYWifAlVK0kRV735EeBDwHRz6749B6lumNmBpbzT/A0p5XrHH3
n0pRFeZwCBdumr/ycsCjafvMg4GWjGGVJVP0DQinB8GLBBpyeeydIBD0ndgZZf8wWNmgNR+beESb
kdHIBOqKr9K47pJSqcQAWTcHUnx9HVmKjG5atj/B6u97DQfVXc4JIRyxrW5kPqPpVmj5NULdJ3ro
szVmNOHn1+LnXjkWLVGv3fB4+9ucTgBeIRxWs2XIuyxIx8ekI5cae4kfVtQOnEEO3yTGvDJOdEpv
mXIvwn3Xqg45Nessb9/iFLZuvEDTjIE8jEiKPaZy3gSmNb/fOwki1qHkqkJqtPzGq7GrJUsrymfU
SPoLEZqFUWJMdCNNWX/ATwBrbX+U78anfpMhnU0r5AU/dGVPeWYRzDtsvqiRaeTZryiNZQVVNntM
zFitmEv6cg+VxwHC55UsP2UcFcbVX02kavT09BiMalZVh+AF17ecN+kTEzu0ZgSNlc8d9cfQF7cv
ZbFvT05vlSX+3sNeZvgdqlZzzxrt2IOIBa+8Gm36gHhFmAhSoTGz4zULzrFJExm5iU0Po7bssNod
77G7IXqfEMoJCc8SmGLykc3SA+due3NQYtg4cnKIvyTSOZJkB46ndOUusl5igW3ICP68Ygd/i2wH
f0CSdnEwF25EQkMoMapvqYeqRx/GTW5b5uCQ+SVaQJbilcQIj143UpXdyAaVqVFC2FUC5UC8NLfq
Y4ierD1cwbEmYFuZTpxaZcRjXUNswZbmpYTCD3zI6DtqJ6OpbAdAWg9YWQcgi7Od2qVo9tyXs1Om
FbcqcU+vhcTrg3kVfHnJzmVlXJX4i16Y1g/n5lqkE29lrl896now53o9euRJfflGgPMeH5nI6N+M
rU/r8/qmkNodr2sSDhTbRnWqlJGd8SejKW10GFoqxlVcKHrPMNSkqPTxNyuNKXEH+L4mPK06XnBV
0dnWrVjI7CAntMUnLjDTUgLFMkQCXLr+IY6lkaRyrF74zXGPVneLZ7DUHQ4+VjKL4Nx+uSrucAxt
qILPMZGHSA6IbBko4/xhi3RqwvzifiW7LYAM3ggE8t0P08XDKbmgHTJXS4ZGu5iWGrkBu/xpss6O
puKaEOYzuHl/mu74qZhWe4OWCukd/exuBRhC8nR5GYF8q+vifo8QrcB3cFVloaupgy6MLTURb68h
c4YN3gBtrwAuBWUrye75OmAM2B3Z+77eqWF/8ePSAJA/sXyPdZsNvnzkMtQe7+1c7eAMY5g27dPM
4exl5S2E7eRx/WF2OURD9f1+7YCoXoQDc9+5H+ORccfZ1mmPEfkyLPJgp2lh3hCsPm4mWyaFTo7m
ECrqcJoJ58/eS33cPBSTrKBzDPJ2AM2AobyK5GPP10BGFJwhD9ZSCUpERPqXmxEG4obHLu5QJR0i
LdgjtUAS6Zkgutuq3jdImLQCyHEJ06eNdCQEoM1uVzrq0by7+j78g6jBryO7QhtSzK9IehbSIFJ8
oX0CUCWneAh/1T6luHMEc7LpafivBacgA85KpIoN5y60mID607A2uzoKm7uMnZG+POosWhitHopq
OukFEOCMQG9lg/EiUVQRR82+0/3agcRNsiwrjALYAoYVwbcHn2ID4mnth4/iacZU07SHfaxP2UUU
+lqlYGxUYu3crCE8InHU4HGBVX4M1lzVhvQB9j3Qnmfk9/wJgCImLQ94wO8w2tJ20t4F5+fa96z2
aIMoHd1glCV/tJlyms300OZlgC6EchylBxSXmfa0ol8rLdtWaYZrFc+h2XNSoe0y2bpCpVRBbSXU
r/VykLq/jWZ+qL/wmK8lZxu8WJe/iUOlNlrFVZmpGCcONxxwS5uRJ+qE3lP5VTKmBflCesvgY7kJ
ttSbAtmN3Y5zwQuO7YnapnvHzuHoAWnbYyHVMEB1WVy0GdFYPEDh0wwkgLqPvmOMKegAWmDhUai6
G8vD38BNCe2bxXCpbJQPd2xCG7GVZLm5XNqgX2mwgn3TcHKWxMZ2Ui1MWZK/9u4bdq1Reqm9S5JF
oqZlFGX6FqXBS/PqWktBecWBFMOzuVOfgoUJgzIVKmaGhO38278L33obeKlixqBSmrgWs+n3AAF0
mus/xhQ4EZZV4wzY52jlL3Ziq+EBmEOevOOxkaKU1GYd0dV2WLqMfDki3A4fE4exkukRA4PJzcR4
UMYgZgyNHgkqB2us9ATn+cWzTvOBEC9P6GbItDejUVBqUq841vB0tRj4ouzzN2sM48WmX56Un6PV
rUbA26UA9N16fp/c1jHFEzGbqv25HuPJlTMajccHaWF38vWOly3T5SvTT2/6AIYnzlz1/ps/Z8w4
VIXZCEVHUFq1+3M6VT0T5jOZwJB21GzfP6GhdTZACiyCNR6KcQDqvIkW6ZOcERuXJPI1W3CPEsbC
1PDQS4CQCESV+PaSMndZe1kPbActMh4kVqSkCmeXEf/fBR0DVBd92I+vNsC5bT/0weXPYgHBG05T
JXY08AKJonYvBDCBn9zrdWvuz385MTnmoaftZDpiQMkgrePtRfrsf/V4QPusgkAweqs7nslGJfUY
DpOufTtHUA+hnGBRYYBWCvHsU0vHhra6Syl4GFef8RWyuIh8vedo6MsRmsSUp50h0acOIFOe37sc
4rJJeMYadWK4ttBcmUG551GJBEzUP5krTV58qwlgIds/zztLtU1vXjRRplnrfDJPfq+pFNHfg9S2
Uf4oc0wXZG7LWqQzMAeR6F7D/It2xOceJVBY7/ZVfnNHB+NRsh/xT4wAOWKR/k1Id2iPs2mi2/Rv
9trMkovWmtia3+oUxIX5bao18k4IV3SeIC4hfXHI7yLb0CMKKsboKo7kUcsnTUEk3T3WU0ZSo+Sr
FyVFP75WMSUWQTqPAPcaZiQepn22hEUJJ4IjsgXk9G1TEjn06nh3ldOY68pQKG97dHZ//RG/7Eei
5Z5h1PLl6FiJ+5sIUQ5hxQ2SmU/C2tFU1c+JMSG0lG0ycxwMzTQCUP6B2thEf0WM3AT87pySl756
Q4nwFSjSHiWcbQRwGGBhj9NgJGN2WEuy+9YkcB9ydjWbWB1+pxZTdABWPdLwrxZlSmHXV1jM0OBk
IiJ4JcyYDx2f3R6QnDt3LwzuYSNtccEnTWGQ+N5iypfnLKnQB33hLmfdLfHa7WN97KBwiuNOGkQf
x55073U0ee2zidBdItDL6Ew3johC1waeXZ1AkWqub6o2Usppby6BSQEQ8lA5uvT6lQFL2FQMvVsj
EEszP0bkRgoepRrr20+Imwxfj1v0a+zX19OXtYaPPxTyC2VHzJ0qb/jM4Zsre9ERndie0L3Ioj8o
LSaTzz8j+hg5G/uVyrfVnUzYo23lPN2WiwQtVijxkM0lcFxSTI06a9QyWHQ1vnnvFzJKG/Hh0Y4q
mrOwXiEZiRtZRFRS/H/CwYx1fHyR4fY1BtzPwTUiAyavbIKWagXWcL91lq9yFS6IeWEfKTfkWaXz
now1p1k9hwnmz+X1tcpGef9SaHHUfloUx6aImpCWUBSrt/c+gp55LnGFRlo6C8TZ9uMEdJA6ySYK
ac96bwIHcZVJqaIInzlVclgi6CtE4G2hTdGdipHnEx+0yOlhKTDpdD1Ej90MZ7/OFkgZV4kaUMof
K9xwrE4SVVDo1iAjJU7dPkaOKzvKP+Ez6utHU9Bp1rRo+kuwXvOaTe2EH+umhGY3B5VIl5giSw69
58oqePwp6hgznPqpGBYPf4g8p0gQzVb396r9Kp7zAJCvm6KezpEetetWrByXZ7h/vQI+XpOWex4B
0JoL+rM844SQWuSfYAXd1UothmMGQESBf4Y2z7TWd4qsOghGK76z5N7UYpqByCTEJI4u7L9nsVqj
8myCCqDr88GWUjfTPxVQ7arqSIG9bmRx4ZucYpeA2YG6sIbY79+eRNo2dIAB9t9UUVEgu2QiXL+f
mIGMU0H+dfYQVNNkmrBaPyvUko7xSBNKeYgRhAzdf8zUC/foY0AGoL4uczyX5s62p+C+7i3TSwOX
g1ef4S30+ujT1+YahXC/ZEcIUM5rEMXASgOE3EffeL0anpO1fuyS/28hBfVWrAahGjaF+CUDx1BM
FRM3KOeYvCGLc7bGNYFYlb/E5ajASVSdxb7nK+j9pds/LJzpoNf/FUChOhrVqI3BzqJUQwOOzCqc
rA3hbMxDBHoa/1x8hMmeZ0DilPfz054bkf+e4fcOUTrlH7PK8X5WaKRPnU9tXjiobdb16XaMubDe
JNcSSEgEOWolSXh4byFXCuLuup7u4wbgocadMbIbH/9YYRajYjqbq8Woa+eN00+Fxh7uhT7p6Es/
IqI7W+Hvi/j0Bps+fBUZQ2xU7Eud84CfsmipYIsGE8oQxgmE9cA3tjqKItJl36ycwrgOYR/bH6e7
27oUUodonPIAq/Kgns8e0MkpseYwojZlcBqjK9QGzQbhu5xSfZ7ksaNyPirlgoE8dT83+wEJ0Dxl
u2krnEJAdYM+Xi0su1rMUp5NsrUffuf2w8MOaWNvDqbVCm8+8JcA+Ar6ABwwOreW+UMbnZnnhWKa
De1h71SsVOWQqi0FoWBrcNcAypf5TYq7NKvYQ6bZGm64bYCVzQw47i6vmB0vrDjiif2eZ9E0aVKt
A2Dd63cVDZUv50QGZtNdK5VXwSdWnUPvfL7LoFVZtTpvSU9d9SVwxNh9gjGOor4AFCjcw8w2Jskj
H9M7bAysAg6wgFnc4MPkD9PF+ebdVyMc/NXqN54ncqOqmzIynF7Jv05LOkJ1wL1n7+C1W4lmscG3
jdLq6t9XiXpGqQA5BDSj/cNYJBm5x4Z2Nbu+MjgdNoGgE5AEhAVHPNKflOuPAXpONQGtjc7e2NFu
BmVjf+aPjyTc8uS8IYtlXRWRMWvow5bBjmoAy9py06F8c4ggDoCQCPm8S6gshCeCMx47kMOcGD4G
qJmGgldkYJE48vfXu7zOvLB216gvzxMxFNkd/zujOTrabxC5gzPrhM/gNfeWbCgBPIhWoIV2QmfE
cbC44i95HN8a8mbygiJDT3S/YNiuH79Q04w/K88uASZscwlPJV8SupP+ompZn3Ei2HdgkLDK2YYD
JnmQwHpmlwgxLaR42fMvyP/S2+TQWiLY8AUR9IjaHkAZo5v0cl3YuAoeguesngv4c85j9OO51RNP
lvxuRBvrRP91pGleXDMUFWHJQUQzLAU8Kh+chR5hW9i0cVYHaai42wU7pc3BI2l8c7u4FDmdPi0h
bt5/9T2kmOneMXWICm9rTPAs2tzz6gwxCiN5/wY501vfly3k7BIszKjqrU+r5LROmSwrmVQTjYgC
DevwAFztyQ2OGnWh3q52AYloK3LPVT9gzU2ZyCMU4wVclU3R44FtuwF0SyPo3Ixy1JwkIw0xpRb/
mavq13iveTCRg2y06+fLsDlw2OD5nSD3a6Ri0N+BK1gzA1zxPr0xH2oVLrqOdR5PWA2pjP2N1ANJ
5jdkzSm2NcxUq6xhaipGryFIrAEtWRB2s8GMrw9oKAPIwZFX56+0IWrqUIMw6iuZOTUP/MZ00qGK
yG6WG5+oFKtVH4Yc2TUXFp+W3vnbJWY6IKEZEna8rCiv5WkV0FqZN0sLIzJSUNUFv6HkhVLfK0RY
bBQxUFVHiu1oZE8LR/eX3/4h1PpTlmzXjnee6HU6yIHxbe0y6Up4xV9hjv6jGlEIkOvPWq9SVP84
KKLAPB8vP8mYWxlYhJvbBjN4jizAps9AjB9vVuRUIE/v07xBT5Q5kJmCO6ATdoZsdWElg9PROH5u
8b0ynPcQpQgCIZePyMQpXEi8DTpASnVben+JpAYBx41AoYh0/xUiOc7Ity2YYua7Z9l9aOdHC2M6
Bfcx1fuLi1QWoNez0EgxaXNWj+XuBQFNPLT9TMP1vQ94t38cX+KQZ4RLuY7P2Gmw0JzZCHuzi2HN
HBynb6yDKktDlGCfrMHXRvfQXUZ5RdEpS53L3GR66BbhUx6H2oZwVCkrmDCaMnQrcckdGpPHk0vQ
76wUSiP0W7p2dqG4+2WiujrF3eDFJl5K1f8Cax4XL9REXqcxBOAWYuwdby7VFLq5PurlJ0ITDhAE
ujzZReBpqfm9BkG0s6kEMCy9ZLpKSsCkStNh3wu9r4wyY52FyK9fQ5PllsJx3Kg9gWpt5N07iT6q
e9OJNUYQhBACzcoQuPrn5+BCWF65JQE0AroWFnLTFWuDf0M4D0E2Hfx0jBIHSI5bEWYZ+8da7UtV
Y7oYlVxfo1iPvwr/WERA3+N1GS47RhLM6cAotrE0xs5kpfFYHZDEmpp9dg4S0rwD4BiKAMdDu6WC
MBMu1JD7oEUve+k8jIvZgDZg88YlwZv4orDkr721lNohIdH4Zra86B8M6fWELhx5Twh7WSdT01ju
7HvlOFkCdN4PLDF3EBvMjVdkbjMy258nwUosV003hgGWWqQVn9zuBzGiGSFOwpDlP3OHrZhWn2Mi
PjygVt1adkQBtiIEc2tygp3EohhJxfBX+qNmLAu88HfhvYD3SPVRzR7SFGXIUgLe/irYMEFwSiJp
XXtJLNyh6jUqBXoD6Vzrc9VHUkjDKXAtoQMWL1KrZV3xe81i/aeTYo+rbVSZImmArKYdYL3iEEex
4FjVHF7t+9rnZGfd3lofTCMc+DjEOOHZDCXVLGYseXiL6+Q0n+GxLlGqYYcy5ytCKIbIDIlPLIgh
o7Xcbxh9Pr8pNug2RZtM2NJ3N8yI3UOoFYsFkYivUDfBNZ26tgx9Ke2j+8FwljCU6pbrtXHksWUu
zgOzIKzUfVQZREzofvmZHC/AMhFxRNAmgf4J9a3RxSFP2L/vu18PsNNhsNZ9oiRb817qRmiewkzM
wFnG5zbjTHPP2o4eoQtE5GGvSSwK3CeBoOd53aFrv1LzgP8VrnWAYBVYmkhGHFfhCHE5VD6NS6HD
6vF8Q3HcaM+SsMGrmHxWmgaG7tmT7LocWqsOhHdFZg2M5ReigutNSr16x//QThmgymj9ex2jn8Wg
urR9PWNaN/ImrzrZ+TaLwduumwbaiQWusZNpxrGAzoV0BvUNa4agkHKHhetT4ZAiEmMjTUKc3oZt
KmBxGWAsFrT3I/nW8X9YDju0Y4nXce+zAk7h7IGoWiLAq655C+I5LjBX/ZgOLo/U9z6Kyk5GOBts
C8PO4I7N808kWA5OJs8F8KPmgXkmVG8hWGfGJcC1pKz/5B4MzEfBRndLlfL3mDh/tYXr1YlkNdbH
j2fDOJ1R1pKaoSCkNawBz+5t7Cu+0yToWPXIncPIpqP4go/8YMvbF6zbAf6VSwFvihiVJ3hw5ZId
P5B3lkMQnX6POu2TwCAylY/kLAc3KnfAngWH/Vs1o4MIFe1Cf01//tHcwNNfGerzLV9IwLRg+PFv
tiJObzxeOsRJd5QYcfY6kP0fhJVY73lucVy54mj1tOcv9hFNxMCpm/bf+ft6chYNzVYRqRBjzNfy
dPY0ssnr0kU+lcF5koeZUwcD6A5KxJx7Ozh2zfyoG+HayuYQurvPgSy83ybc55WUGDClL++XihdL
grCiAqnLNrY1G9h0D/Htn4dFV5h2anZKiq/QFdfPPxAkY4CtiM37DJURJSkPjIgQJEFKcweOb44b
rm47IrlD6nLcGnvDuOmg0YDqR0jF6OHE6tbFBDERu4KtxR1+4K3e93fNBsfdheTi3eWnPLc6iHT9
IYuAUI9S7qabrQvn71diG5uzLAvDOhoNH+0ye9UsEhU+5NtduyIh6Z2he+ng/Y0ZCtNtzMuTQX30
a8gT2L+U/Fhoacvsnd66eQ3vbAm62QhE1A7Hz7i2rNeABj0CqSZaOozGUp/N0IriO+tWa1MHZvMK
6lPlZpWPmZIajcRUHrAIFPvGlL4RbGEanXihTiHeat4B3XD6JjPWqVt/VecydPb3GEBaXBuBJfzy
extmJrNW/W4PI4qNv3cVoca+hn07YLjfi5b2MO5Fx+vozJFpJPUL+UTF103zx9OXC/O0b92N2IUe
Jscr99uOTOqi5lC8F8+G97SFk/R2JvWb3LQtfLgNHKBzlQE/VbRYXSY+iX54++ml7VhlRTnoJa3u
soVnKBwM7KGLkmUIFvygJvZmP0Q1A+mLbFhumRXZ5Uk8qi14TE3IqNA2vrYDx9LnScCR6sQZkBHV
hb0abYHX5PYQ96bRdXXIp48OQGt9nOzT35KWJCSbCrNbtoBMxp1AvZWPKBmMkw2gun2xiSo4CimO
H6JpcA6zGoiFev1MuF8BA6JX5Ax85aO/W8UTHQPmRFrqwmYeHtc1KQe7Nx8RqxPq9GAzhSZm8k3w
4fI3yzDAE03Q+/h+3etek0YUR9VWiCsCyjkYwsJm3nDBGjLra9nCcUExWLRhzrPvD2ytQEnjpR6o
CdWgxJygQyElVp2PORv6EJJPdAl9QZOQdnGuNKi0dSpTxBKt3TBFUX3lVa3Nfph1CkRuswcRIlVU
+ZqolMMcLwxpRzdu0DNDHKMG04YEMTo31St88u1IfivOy97qCF6T+iUI7vkIMrOzE4tXzZ9tjo/8
Fj4IDPXeI6UUBdESfg5YdQ3WZmJflC6lqzmsIAHuTlx26KhYJF1Uhppddlq1c38iJwvJeogKjoKR
7dxwUyhCQuOfYX9VsWQ/PXIhgttz8fQRLS83+H5brrFE6Ob17d/Zl3hJkC0OlHEbVESTB10wpAHY
yRa4hoTqWzfBMoVsLO9mpitxqsLpknf/bQvnrQKboN4TnoFDQ27lFqCCmX6bygK/ssaEOoVnRWer
oOXh+IiUgh1wlevPllayDjrKlwboQejKCjcFVeTCFzc/JU82eIYUg3j+aRMQgY8qt+ETUchM+XOL
eJf65c6JSv4bIbm9KamBr25RaFSJPK30f5a4/FI3OkSKFtiwM7ZyIwWE1cAL9BkW2VpDXAqrq67C
uLYRNU4xj7nwFxZ7kpD+UGxJvuOYmyyKC9Vj0C+Zd7I0lDYHewXfgTansC3E+UeUzTZVoVyuUmjW
6aAhGGgvke2GPkwnm4eE3gTB3oWkarDDT9bJJM39PZDyOBXz23QNWqJ3cBJIdj11P55s5gDajnif
T3qYUxqQ+bN7JF1GyJuO0wikm3Tvkz/OytrTLf7MwJrKflEubZeBs6l11Tnf4I31jtBEQwuY15Qi
x7/gIVkJN6JHtG6t+MfdCnzxXVZ40acsMZmHX+56aecFik3vJA7A4o0l6NPS9nxgqwWOct+FLlDf
gCdeX80MAWQiXRN8RgwrcAOxMDwxn0+3cWr6ee8gdPbJeZi1Yo0G6RNIFr3K6C0CRNqHXmQmYNSf
+xygctrTVxc22GibVK4a6bJ5seLhRqfMR9XuNVFFS0p3fxQNI76tWPESFSCrMLR76Lpkvf3yvpMn
QSxhNP+58hbiEUXZsKzna09oa1IsRxlhPGE3wkVf0pCJSc/+fEVd/XT6TWJlldyaWeVn/F7YlcZp
HMH+siEi95fJ+hzi33EPhO0gPOqwAV3R6DfUl7CA48fILwFc0RaWdAnUqDs4kp0vTJWHbtvp+Swn
RFh6FvX7aj9RHE8dVHeVyX0C9JV7GAyq4SxNMbjIfEkOzYwRTwFboXXtZ8T/GxClESfphMfUVjUx
WjHeGJaD+57mcE+D0mRXzHcFzPR0nl5xu14chtUqRJZf3kVP5BQ83OZo0hTqY4xUuS4bJUD7AS20
3kKFSFK+iFIWlNPl4iinP/Y2T66PSxFjPaLvLYpjrLyT9JQqBBCtQpAtzst+IZ2i2EOTPNBWUpJ4
p5Vb/9nwXu3lsTr4yrJIt4LyK7uP0qVKJ8HMRWg+GnhocYX+Tk7SBy4BtAh6O8kaCrT7jcsUjo2b
N/e3wZE2avyO9MWC1V0FRbpa4+Iw9kbjTaJYKsRImp7nP/u3IMcmEfcg8226hz1Q7ZodQlgfCwkq
3iOfPmU8F5COyLSu+57wymimfjvX02COQvj6LCUeEr5jTYKInDuvbcdNNtqPjKGWuw3BOkIXCwil
F0lcQC5uv71j22M5C+0rbpr4pdTAcSWeLIkrjj96qykkks+f1CrOaIInJOQGJkObvl6znhKjlmFw
aC/Q1eTVdkKT5wVKLWfQlBk+vJG0dhyT1dndaEMzZrio3DXJ6H/zCH3wYxBbUfd0ijh7EDcm04dz
O16SdV3CysbwGKkVD49cFxXQOEDj4FoqSNz4NqgJE2qixHvT2AbVOGbASvJqf3lt1f9K03LF5Zf6
EFG2A5z6srPYx7iLVTGJQiFTng2HbzdRitIf36GCk+t1PtamCwBBnZyareHLTXcw6tjvNp024lD9
e/o1Jb6lwP4atgYR6opUyxMJEHJwcJeNn7aSHxWbD2EXXRHIu6RNsTpzAVRqkRJkVAUZXL1VwsIj
gpsLwfbyLF9N2/pY//9puu878W4DRqPP28O+rVTeoaBpCPfn1iiM2U1VGXtfoKaxij7v/Q2WpxVX
Cg9q2LYAztTDoBDfIY0u7FtqTSFSnZ2u+zCOMQiVeICIESwv9jQ3Eqaq16VdxE3qTrNp07nmT3Si
hNrKlwaZcINbCd+jWFbi6V8+sZ46kB7N3UDmbWVRAwDZTkcsUJ/juIBn9/jN+c22JmfPrqI4aMVx
APy6ZUpmTsX6tzXLd0alRyiTzcsbOKBO793QUYriqSEO4ROLzNRWgP41ui5Gr3xBRVMDVdtYkexv
TOfAuF0csCgy5bGjKUmaJcOUbHvX3M821ogNYAK/eOJjNuvxoWvB8w0nq4zpN6q8cXpSyYXG3dFA
lELRtl9SebtGs/5H0s/aLmPUU6KV7M3tsnhwqSBxeZXbfesHEDbT/FgxMblU/kQyZUC11r7GbaAP
wzBUcVz7WpVGY9ecQI23FPXiN6VHcyJfCYh1kz8H3rPDUkX7gtR4jZ5HHYsXCRFli/+hJM/I85WY
I10d9aO30KcqEdCmEcRMCr3g7rm3uDNYXVHPCm+/WGsh6pR1iFTvAFmedMSUCYS4BRU3sYHLqogA
cnbCR6zMEfDo08heGEhSZKf0s+mu2L4/5F3UZSR+QE7ZZ5DNMNRu9yGIg1fSLVT6D2D4G7NeQM2u
J5xZWUvd1ue6U9MFgLuqpECN5Z5MDfl2LBtxYqvivUMHdbvrG6DvkT+JqKBM3dtvUqoryC4OKAC9
ufIdmoCcStO/lFK7x4DWPHNylsnWdC8uX+9NvHRi1SUjUYEnwuqDpGju+ibe8jSxqjHGfumBubpG
6sljo/6WpA+FP5QLpdoqz/32K4/wbt+B2v/nUXtzcdCKQx67SJVIfY0efZ2yb200q3HwKm5U0v9w
Dwo2DJpZyuXEAcsxsOpK/kQv6ljlnkv6lbFKwtqD9cpqb98JLO3KrKsS2fYiuVFyaYNZGw7uAOWB
PLyjQ+dg9OGCpFTtVSRPWY5FrVlU5hn7WRJrfuRjjtoqgUknUZh/DiqXl/OSmdrY6Na+d5xvUKD0
hKoGuB7aljCoxgRPK0IdEPsBoo4ObUjY0GM0K7W+1rZ48UHBSmpyAiFPziXWtRQ3Ml4pySAhh9tk
XDTDQp4BBFz6EpmYSgNCq5mBoZC6b5LUuXct2KbOY6ZILqXo8SMXHCcnnotBMO/qi74EWP3iqWdk
5IxXtRFsuo2yCFoHzzr4EUeuTwx1ma5gVmoZG+UXd2BT1AKcdJ0H5YdtRWyIaLxzPGmF7HPx9gGQ
dlfT6x2yUNlXUOU894hBaRAiJ+0oDwavQ3Ytd+5JMfUxDzRBHqR5isP891D+1HuHDSSlxsP+ZxS2
8H8J2RbDylHubQP1oC+G3JfQ3VGYet3p7fvA3hSkkKp4/QPFANxZwz6C/97+cYjT6LdV7jiVIh9A
DR6pta2i0ZJgEJWpf9Rs9uLrQ6d+Z9azJPs4vRplImQbRNjVibXtgr00E5TC8Igmfko7HjGT1p1A
86DWfW1O+PCyr1stGidulasp/mRcNLPJsfSPuVcbQsrqhqJmMcWbrTAqJ4tVOfysOQPT71jlyeIb
E2UbhiBB4xWwjOwJL6eswAjV+T3hhjAKNOwTyWmEJ39TTmqtTG0Vd6LFtpvgiyzcVpEivJNeqoSG
jTwX/Ysaa1rAFi6G87KBhoLgDU6hafOzTzZ1LGvVyiPPMrQDfsBA/8+KpcjXxMA/GO1F+WxEavo/
pYDHKwD7OW9MzpFIShyT5AHC2Sg0I0uySphd7W7KTHH15a5ynxwNoV81f9xh+0YTR8r2DZPCp30t
oKLpcHsB3hS+SnnHE7b3iVRaO8ubmLaguyVYXh6+/Hp3VRDVzzgSzF00pddZsALl/20NYnBlUUS8
tJZTz0CObwD7cuI5JoP5BKFRNdDkWLRr6ZOC53sJo+jNgTXRxzd+KJOCJEgYh6zyv5loB+k5Q4fV
IBbbFc+2ylcY7zpwM35oQdD2BoXszvcyHsZE7nKLT4wWwCpIYCKiDTuBFeo6L9sivN2B36+Ie6yk
VuQSwpXBYOr1bS4WWVd9TF+9F5rl3XG7zvqMr8iItC8vzqkrkd7KrQk8VvtQkhWJOOBnL8kaUk0D
nGuPN0vAKBB0E3q7552LNL/8hWwNzOoUElRF/cRpy7b8zp+qgbeySohpm9R9f/vyob+xzuXKyVKB
nXHobNSHsK85CLHGqg7UU86WWl9mYWuIyLu2adWpXUd+L2jsD12zxgWYKPmr2z7XE0Oku7mj+x7k
agSTBU10wvDfRxfH/9zirIUw5Sz+v3RsIic+gCVgtRmRkL/RlAhuAcKLcv/JEWDuPfH/bC/DGVFD
OQxLzdUr69dXkuEPYM9M+yf4Tf4tm8cfVdTkLbWynU3Wv9NjOXOm+bxwZL0VcY9ysj8ySpkVcmOj
+FQs7yrSx9AR9lPdvTLayKBjlgjiS8FEHUNAndgHiuEV4iNKhI667vmo93t/+MqOPuM9R+vhi8kG
XcICdJEMCvqS1vB2hcE0aiena5AnCrNgllgqsD+wc35OHzEj0YA3fXjbXjsu6RxNl86hHhulXXLj
UxFZlnwPWSdKv8y7H4DF9nrRDdP8nvXP9QYUxmM6bvQEkKDU67mqYeeVmI19Jbdaymbd9cF8CxsZ
BXh9MC+ZgGfRTy/y+ux942jMjq5wYxL0kL01mNJM/kEhK0BRQW9zc5Y2EH+80OIUh0ZZUvKhBNE+
9LS5voKTIJXMN4KErLsufNb0x3YMR2Zvg1Ip7rpFD8zYNE63LHcwYLQqqtRrihU3ccvMa1ki94H5
EQs4IyQKijoEHixo80+34kDUd7E05s/jCCQUe2neK/9VfX8InedQmCZXb33SkYqYHI077SW0Iwl5
BSuulSfMzVYK8bbXxPntBDL61h4Hv9U/lyU4jsFdDET0VbpQFTp9RuTbk/Fn/9rEnM6Owg0tj70T
4lZhDwzqp9D4oYfI6u4ZPXLeLN0ZwioMZV668fgtnfLb7dVv9wRk21j2tsQJk814K5q5iVSp8run
OrDy0bU7YShcEgdAv3xdqtBkByEUbRbqMxrOEb3vX2rUx+q/djKYLz3C1+JQ7o3n+9eLRwI2h0bs
ny8Nlcy4IEiREGX6hhPr+4djDP2rEf+s9e4u5v/CbWy9a+b9l3X3fAOIuOlPhIL/5uxdohfR2rOL
Sd76LCPu8MutBopiRonpmHFGdWLviR9+tuV1SSiZ4i+Q7tvMzE4ntceFez0C4aIPxeg4ZBHkb2NX
9X5aBLG051WP/nNMqNK9NbZ+vcCKckLO0RIs3rlPajeJWfxnCr8WxQgRQ3N+xBNf13kcMWhe6jW0
+jUrpqUEIvIU5eVoqu7pucraxJ5DaQHjP/sXzUujEkAm2Pzwm9P2LqoX4FfgtaBffl4ZDvEqkjzb
pM3DDY+GjczbwiepCY+CKrfTAuxVE4hTsaSlUJyoZolFyR9+El11IaPYVbeVlwNLdS1I8Di4dWAz
m587fNtT3u6rEDRfWFVzYXbscVyZSlYSDKGxUzIKt1cG/wHzWH9UT8GT0XnIWplw9BUyUFBEtfIr
pN+ZbjAqAT1IWxW4G+/+rOwpGp6yjKRU5wQ2S0sitT6TOFix6WhbrSrNFUIdyeqcKt1y8VPp2Bfc
N496PHFoPHQLp12K0WTdW7lo0A36x2tDQrpy3G50Cy/bkkBkwMAR4mY3koRNw2zHETJebguajn+Z
cZd1feGneqbQ2mbdz7uHzocnEyYntI76l+AlufOSKrJGbFI9OJ9JM51/Jn0ZngzFIlZWMATzHbpF
/J1lLyOoRjF2lew19IsYUna0MgIaiwZvkWTdwOoxgVW5pvyToJDj8Q3Hj/0LFSYLm/s/D9qKcmAm
Knwi1p5iMqjN3iNo/gJu4PAWSZamBCuYloR2NJYXEpe9ozsh6TFiqlsQp+UWkWOlLp3Bs+2yOwSg
GWFm1wuOu7sLsfcfM4kflmT+cksHLbPucuHn7uQvjWrxcS0HzyRpwDLZhiDsh7/6tVJ2GV9ulHz1
AZKMnJcglCpYAyPEp+X7nJLMwObZVoV8SzFQx5feVypIi0zjOeLRMjxI+aoKi3jX0VDbDBghf3Z1
d+6mhZbX0jBANLL79tutm9es5NV2jWnij2Xd5HXx3MynOtwnvYI0rn6sy5TRfuXWRaGV8m1PzwId
86Elgxy6iw8iNveACXQLi1G7ZAw59gsixNd3Mh/KBzvNlyRnr0YTQbAmVRH0hyjS3NbmMxgG6OH9
cW0xPFaj1z15awILQBdcIQPvd5CF+HcSHHKeWfU2b7QgMs4HHVKAypBEIT3ytNaDlb7qBBTbxb5P
WOJVmZyeX0qPgWdUGOcSEJacOUn8fklvJKi7MxHxatpJheQW+CJfhlbhUli8baASL2edIq3g7Ucj
6a9y3CA1S2SDRkuNWYmdh9n0t1hVLyiXvDM6kYk7bRoaPOsfmZvj0r6YnSl0u1OXoHjtKZt24vvC
1kX7dEucWKVvP9tGJop5n/vvqfGv+buIRzI6WwVE1WBL3wzUzitZiKQHINVQdU6qdxv2iudLruvk
Mm422wycCqdphaCfe09SPin6lVCj52gsWuLsYWXrTlpSxfB3f2YENLX5V2dr2kQQ6fozVq51edT8
eapK7Y49BZfrnfTll1Ts6HIC5AI0wvy3Wc7cLRbBR/tj1SLQMlOCaf88nMVJ+S+VlJWSV3ztSPlQ
GIQpydM52TwgcSQvr1j0C+rG4PzEyGrN2rwJlQKFggmQUkPHtjAvkJYNI0IIPgrSHDT2bxzfedPv
8lnsqVKFo6WUxEp301Kbj2C4tXmwYhcrGZyZvcodwrYGwder9lBi0/oo/Z05xugrFc7LWysfnfQp
EtE8rIXWS1WeqmP24D5H45SaFvgD02tpUi2RAmLucFQixKjsUgQUHR27ENAAwWlZ6r3UCPQBS0l7
vIbwcm1WrLiVYryGHpoysXHojD5nRzgzCwi9I4GAIrQ6GKzivraX0KhxpwAcQRdweuVYhRH7GjZL
ur4uDq12DnwBkwMtFiOWPMj1Sic3qzIi4ooUsw4gOJ4uLmFmFwcNMXTSw5jzUyxk709/wAuL9ej2
6srJETo8xptyxZ3beUV8id/l56BkSdBqLCAH+lwidRmUJRdZA3Nt/ek6s9o8LdnphYZb4fud+Rjn
c3aCZMvbn0LLajlgxIrZsgVYcHWvPutf3c/On94IsuSYFtRWlt2hReSJvSVBfKubXx8mbd7WyRFN
M0wZkIBDkcrT2SPiQeluWIm0ghg8XfitW3ewI1byCxFrQBUnL5m0Khq/vAhod67meitR3APvpdsa
beXkBg/yWoO3G3JfhQmsUVE/jWY7PM/8hInGgkF6bcDhGWJyxEK+AVRrQtmzT4jEx/7lSw30CLYp
Br1x2y6/GIqVMT/2PH529ebJCHFAYtM2sNIyPQ61lftRQ59gRJei+6ldD4/lnoteMtIY2c0YlPFx
y5F3ZkXL5BDq0m5dS82gVUjWi1tVBQ2BzjsdHKOjvdytwqCXZEUrAh+EFiPGidxTDymOw2CSES/o
zkMuGvSRwnx2gcVWHPKsypn2iUcwDIGrwNlyQF8apsr/PqcnHxOAOuIvDL+yj1bjU0isLp0wrkpP
pox1kIP1zKsOnTU4WdK1fLA5yOi1cWFVAlSbaYi1vz5Tw+G9SLWNWe4bs+ucn3Sqf17RP3vwMJyV
KHDCcoW1NjkZ2jQamk5gMxuI/4t6UsjxT/AYmpq42OqmwZ5/ephizhQKTeBNptJmgl6CJJD9XSNg
56T32yJq+1zVx0opSIN7l+bjB/kurJ3+7bqYa4QCtMqlermwlZoeZMqpmnNAhF4gDXkY34UrTmYe
xX2ooF3SiXTjPOOQi32TlSNSszjSoBWeINjXBtfehV3vhxvlZj4CTiYhipZkm0pdik2x90POVbwr
6Y6f09PNd/KJq494Ek5qVKTvetGf9r/CdL5FZggU4Kbxs9/IlB9TmUPqPjrZWMDlJFcHphLGrhSA
dpcyTTl9IDKFnL+YQWaNXjkSGmXelyntnU1pvcFMNhJ1lYpE2zcs5y5P7KgeXGhrrOVnOFcMC6Mc
d9C6ibOjl0QCfT1Lllyio9FLaAkv/wMTEiOvjfD79ncNmvLXpjW+deJl4ytoIB2TywRLtRxPoDRN
rUeWik+ZKIC43HXm1ev3dQZsRomMR4ofBrNhgNnRGjEl2Gfn7vc5YsIfOR6DrO/UTBMhdFATJyGn
ZJjR6ds0IrC2tXQzQzr1hGdFQBjN0f/wwtRwkn/SkMSCsGBzbYdkvlHBdTe/Oq7W231GxE/Q+oVL
sp8MwY3YGmPhRQMf7/UQmKqzBNzWu/4GB/RMS2fb2xQaKust68n7DSz9eo0kZY+1S6AuossKbtrd
OmE3ylh8KJP4HXPOT2obYNqHnypw3EMhjdPPqdenvUtUbA1AOm9I8jTOyW1CUAXxtkT1GEcTA9Ne
s9U3Y7ZkLRFP2ke6BMtvafhNJnmD7xO2Xk99sAZWkv5w1f72OfqjOx0d4sdMXnd0MPWOxq8Y/TMa
un472q1U+KRt4hjWgGLDc+6qn1XbUaL54X6VVz2W1LC2R97GM442a+ElJisGoXAs0kDOemFxOVOt
2oFOnVJrPwG9Vkx7dAiay83XZdX0iVsfIN0cbpVxw5ZxOQIE053FbUME2EkteENjjdn7Har+MWuD
5120ercZxJKdGerL4TdQqGWm9w0zFL5y3ni62LkXX1jynYc/m6yUJJkV+DrU/UTkxnWROjK93N3K
pecdL9wQUv2zqJ+3uRlBARdGqdAU94Tong50A/IFIW9LOiuggHSgROxInlNjAgaJrfuUoRnTid8m
C0CrGg5KBFSxjj9w2W8IARKsqOpWmJ7xE/jZ23dj7l6tS4EC3bQHZ9Hmgz3ZMEVTaQHCkoYNWb1n
+IHOyFdIwDCAKgtYcbebdw7cqkiaSHLlLDieyQ+QzShc7Pcxg4KjWrzXpX2Ud+mop4HEGjt9nZiG
lLr537xVRVuOWKyR9uvIeTBCy99UZ7s6WRX6rWiTg1zd9DfPVbXiGJUD5/YOD6MBHjxT9SD1Gm15
esfJokVu866zairBzIjg2dRfqveY8Zs4dLWhX6ahxSWgf7fLUBDVRTBzHJtvKWwIkrEyXGsWN02R
UErDo+L59QzhIk78RLehu/XlacW44dCASr9l2Xh6PMDZkevoGOTF02w5ZJ4rYUL5VNZVn5bDnkmt
XZLhct9e++SO3Cnkl46gtF6irujRF9AqJaH539RB62gYHvW5golqrAM9RBJR6DirSl7odJNXFOMH
rjUKAEDS4W8KRs6SZLc8+0DynOay/KuNtMLHP6lpW42TUXKOI3Z/Ed/dlC/w/RFYGP93cn9zTEzm
Wwot45og3n2ND5HySt2VsNarinvapdRBCKLZcH1CUjlYyv9nfZ8lVxsb+3XxMDE5vVu2kUZIf+5V
tQgVfzR21j4wkfX98BWQ953oLkeqAsXWG7JB/7aPN/+wjkqHGAKv3/tlNdJ49tfeA9vQ0GGLqmIj
CzeGfS+Ol0ensa8g5yeCAw8wKjNnXqff5APTCqKzM4jKEtk1VNZh/L+DpCGsCPybdVAAlnaFmqCK
9fMLPJeZcXeQvcPOLBA2SCIXKzPXqQt15WfUJIE/1sQxWhzYI0rikWtVFpuNHDlBnFZDVMzGybj7
B8P/eSV1f6rI6UAuv8Y2x2vWz1Sig+0J1CDJ/BrDk9dzfDhdeBQPiSULaj2C+gfXy0tS+DuRQcE5
uJ4BuTtELO2jV/nU34rR0LA3dJzSx4kEqgDNMUCr52PIaBZDvw5odVYa+aSHiYkU8h34ITTDRssW
Ju72dn6Js2KfSZEncq2HsAU6GbeaB3OyHNEau9zHaG1vus0oDgzOdcNwYD0sxefnkuu8mc2T+T8q
eg4EPl7yfrJUQ6U0AdkA3/w5y5DgwgwQ72kERQJBw1ssV91GHnDJBKbmeSkMgezEVZGO5tSrij8u
vAC3w/aPSirln4BxziakP+vaRf+K6vY2KG6oWMHY5ll71rO7IP9Kq3OOgMlWhWvjeHulk8xOunB0
Q4W/ChyvImxHvGNZUmnA9SwZg52jyd+DZ1HLH2RVgWE4yT8+Qhdtis/Lx6RhxXzzov2fUgWSF/bg
HIDajAnBWhEKmqH3B9if6NoCJsrCkERVFy3Y0wpFds7TPmODevXJ3gRsYEz22zrun2MZTF1b3thn
mBhvBb3U/47SrKoYoUqOMxq8uTSgcoqLsC4COWWo72ECaZwLyAtrj/LaWY5QMqnocEdiGsjxwjbz
1vlzuEGB7LGVYl+p+KfyqfZw3QmpV4xuo1RlRIJKpF/G6Dv5ZapyfqsRU0BBVwdo66qrwahXknKZ
TkT7iPwo1uYwW0sU21J/PQut/IjCHk4ZWJaIt2JTRZ0NyjF5gCG4UgxxdrQqr+/os0Hz0dxffPys
yfmhmXK3nii3/Wr6EzQAHr0d/snwP7+QpJlsaTuEHEOuJ+4/VogdXkiEp2CgShu/UlA1kmvvyQAu
J67Ax418PTUZ6hLN+bEpbDMAD+bNvQ2R74CPjuxPifTqqSbztmE/chURFyMt92cs48t7CymkiiF2
19pJbCesqyoW6031Oga39rY4fhgDsej1nNaWq9Neq0hqKMUAaC5r8SesvopotAjtObDlvTMo2Fb9
81DNr1yZ/MSQNxeEfDI/5/m7HVLb5wNYib0n23VD0LdkP7gIwXZh2rLq7v/rFpHFd/0W+FbGPHmM
8/mayYKDLd97hRIf7XLRlHzOv7CeC3V+RigcYcQHKrenjfqvuJvtGmqKt2LMC/C8TGL0blreN0Kn
bc3BVp70wvn+/iap77CdqPMQE8Ke9ntcgW2tSihuBVu65PrBa9c1RDaftcv3L1KOhlIzZwaPMuxy
2bX1aChA4zzVc9AvyHBgpIm2PKaSiufCWqNWljIrJA5rlDgVc/MRASCuq37TeDmVmjURoo90/WOT
6WKuy+fPwQfmej7UiK7Z5+mWigxExfgAgS1DdyHDxobShm5/59lKZg0rfOW1CnYpml6vSU7lKrJF
fFXISHwDnrDSLdpzxtcVffi+STYwC0X9kR9JxBsX+wCvzvx/x/KRdL+kkTzRErCnGPWvQngRQ5nN
gc/s8kIJkQGNtk8+TOEcZdEe7X/DePAAJqdcJuZx/+Og1ui/A+zcMgRzlUg8ei42LEFoHPbQrozb
y/u706ZgYmlihx86NqNcJTwW+ZrOcyV6sisg3nM1IlanCOZFeCn0WQ344aQvCNiM6LE6QZUSEYAh
8dxFRXfTSpLLPjNa2YuPrXtqC5+ne2EwMmZdU86TWxXcaHrboaFQfBCLt4bJhhbBVUBJ1LhK/Vue
EXs5UlOi6ODmeH/xNfR/qFPBJcuB8BJ9+S8/+7Hfj3jTf+yzn5RWFGV0PN4lxMYB3BDQzEwoj6IK
XpL3fyWoiAzQCM24ED5xTgE/b4YgxXM1zJIV40+KjsyuRatt6IJrTlSM1PrSgYBWt+Hitlw1oE1R
6FqUXEHxidV3nCl9u19Gt2iMnd9Py9aE9c9j5aCNtZQVkHs1C8/8vb4oF40xYcSCAGxXp15uFbv3
g7j6IyJsviCIDBsG7tPCGu8i8OhQKmJ7WGNIMnIfSYuu2EGXJtg1rMj3np0Fb5s7lGnNiy3+zzFe
Z8fK0svc7Dd4/vnCp9+8ZEL9WD4XvS/gccIYFNKUw4HNo7c2fK9UlE8Gxd56Z8MEYQuyFFsTI7jt
RFMeckHZthzq9V9iA8ehFmBgj2UbJ8qL/z1W4Gy3Ma5b44dXpkk3gfdtBSFjA0zf6lGuozP/9GV8
KPOC4us89RDZMjrnGOGXL6ZAlYBjm46EFfnFATG0oD9VBot/z472etxzj6AdiTEbVpes5fIvv5dX
Mg2pCiV/tQVWmGofbUBpuEOvLO16yXBZK4QAGE7HFTT9gB4/Z8AwDbbUrU3ve8c2mfEU8QcyRcxn
lG9IxQ7hjCvdYxfxdEpL4oDOvB0d2t+U1qG80QtbTHxw6XLp9Nxb2ma1U0ABxkIGl+IxNQXkUeKP
iBSxUg7aNIA4H/ghcLk4NHkAc8pxEtKw+M2yM6cum2ym5CW3opBfpcQPY5foKzFkxaNExGD/mBgm
NWxBEMv4RgDPQ/zSF61ufrjjp7yXeXiIvPbFqAM+i7SCyLNINIjHe1kPGR9DOIy39x181DIgy4vR
MMiFX/JnXF7cZWtWSLwbSh2RYzJIm6u/7PlbrTFzyX8VHLfINHbEeV/MG+T/bAxRxQ0RsEBjPpfI
dxOSUC8YeMGmnrM+HgcslAtq7MVR7pKFsQgvOfZ9oEf73XH9+BW0AH2i1qTGRWDQSxUVg5V0xLtj
RuCw3xjM78MrEN5B5KJmMRmR0SYKLZjjxBQLJWvmWudjjHAJaWTOJc6tN6szWK5CdLWKw4syG039
fcMjfQjZF8b9UE2/TU4SERQXNYakN5Ru2iEQtsU4x6c8o19eElFd3DxS33kstXwc5R7BXVILLtYk
o6twVDaQQ8WN9jxAXWldd1bVQU0KyOAridsF2xWgpG2gIo75paz1DmUsSyiwiQJi86s+avvj2pys
f+fy7Z6LKrigySTlUS/vZC0EXjK77xHiWZvkpm5aE9eBP6glN+aDwxZiJ/SSOArabmdROE+nhn6K
5Nl5+hZ6K43Sy3B/Dh1Wi8ocNuw0FnrN7j0P6eXyiwytS4nKhk30S5HIF43kxagA4At0k4vt52YF
tpp6Mr94snGZJeJzlpYRaCjCeOrMYP5Qb50NCW4eJJqxGBh/jMjZph0OKro69UymWQLYbMc1A+8b
A44txIgZWQJGhql8FafJ1u5RL/+LhO86SqRLYSf1LE3icfjHU2OaKEb7nTuFq1GpECpeqx5STZCM
HKuVkTFjeLP0k5HBxPRsDxRgZfuXrXLeieWEWhCxhmG2Yw3phUiIDmJLUGSviHoo+SXKcclLE8mF
L/T6Xlu3zRfTRKtW2mvlcjm6lqvCyYzm0IhRtNrLbvJSCtjm7eWpvH9KwyAeEu+L0VPcGix06zAU
t0BeeM/Zlx+P3r0mY28Bp2yAqV3a4aX9nH4TocpeZFo0t1kyPn18gjKp/rrFOlO/sM50DtHRLNb2
BQ0UtWoCP7qRqsFlyIFKEkW4G0Af44TTKVOW5i921l81f0WrzFbFqOi+KhhC2DklfyKwDmDtW+ef
N1LoI3ytOv8U9JJKffKBj2Sup0WzLnBQZoypA49y6VJY4D00wCf1N4L+V5WXrebzhzZL+HnF+C7V
TySmVjMd96s3Yx7SrmgS45M9QGw/rB/Ljux5sC0PIubf5qvHpilFixozI5zk7YaMC+Y4JpQ768fy
aRlT4Es7ZhBoy+qnqOYxzs9OsuzznwpgL+7n+F9dyAxrTXZ9wzo85SeXmDdnErGFHGNqGVL09KBo
QEHlq9pQ9tveP+6p2WEbPJfnb8//yzlhbRSKW3HvVsS86Z0jrcN6bD+1xrYQsRNvLv0ez+hwjxPX
sGN3fBpNlVQjcq1OX9rrGclkvdukdjI8ofTbsetwqdHII5iKK06hsA+kxhoiUaLJMhRoMSFAeubd
NBT9q4gV6SZPBhGcJ0n6qESj/S0WglYvaHhIk0CExC52lAoINpCec3lLL8KtG1Mmgx0BVLIuj3aj
09mJnCySNweYQcypgW49AcqEQzdkNS/Cw3AmwtYh5FUPupW7zMwS3rwpFO7mftXKjOAYTe6k6ANk
jJuHdWYx6KjXdLt93bOpiWEtge1MK9JPEFOnJZO63IMXiXi5AiMdDn0pU8K2eRHwD189dRUJVSW5
DVJtLtjTXd5VHUFoiu58OxZbBYmJ2IUw2KIKTxwXu9U7umRVehrw7jvGOK7QIvaxuD3MfFMq4ehU
fdbxjzuFonihbmni/lhSoX6FZqjv8vs2kItKhXfSnbaL3ynpGbJQ4AgIg4g6F2WgPxphXPUR4USF
V4wCMGQt8KtiOl1O+lUoZpe8qOto60WPG3/LtO9QoVE2EytvAuf4jSvXjETTOU2fHI0H1opvW0KJ
F6BarorAh0FVI/7xeviArpe2Xzy3tvNon52BHIUY+byUUyDmfaDjpJCYmBXYcafTmZo89lA1bB77
As2l3h/06Ud8EJt9XPuej/QQJUZqfxeh0+tkSYIFKVmupmTtznxA8w0lQa9HV+beThtC/LUHSlk0
rfuHAYYMsVNMgqZ4nguMJf4L/dgYGHBUYrKt4hN+et7PIRsdYsQhC87RoZV95t8y9aR4As3Yr7gI
KBUq8JYqw9bqD2/RbH3N+1WGlKFSpeh2sX+1sx5qRSXAAA0JiWxMMjWDm5quYew4sCs++czN6iSJ
hQC12Q5nbdcX6QJtGLN5oVRYBRe9ABoAsrQQDRT26OlbusRJ5VnNkfaKaSoVUo2tyLg96Llc6C2l
O5+JNPlK7DvapSQBEIfiwTgUQJW9ZPQbhDCP5u2jgBGcaRiGJuoctLSdMZakxe4VjHWUyBBqJ+f/
m6F6LhXLBtzgdokx7tYdC8vKolWCdJug62tea+I4df/97M2zfTd1/RqZnNpJ1TaVUJ4uUbfgRFE6
YPrXqfjxfaYjsLqWjIHALrmtt2fz3y9guEhZAiFB9EppFFTAlOBYd395BmwLSC/yT+fB27C7+sBS
TIsMqAYNPVPe/pXop4Pe7t3w0gcQ8nruLJUQM2cBDwQG65wIRiqIsVyT75DEKupf9b8Uz54TRHu+
kFtYvvKXqCrsvhd9eyE7SBApdNMFADm/VKYmOwU5JRmQ/x1rkW8YROrsZCcFLHLRtVSjhVrMFdyO
GLaEs0SuDqvX+4vyFH13JYOMM0ae6XeIerf3Z0r+YEVVHbSrIaZ1+J2Y8PCgP999y0Ms1zVTgNDV
vraEqDp9dKjc/jppMj0r6wYVgfJxyNl5gArvjpELWQQ83TQskexscnKl+1FascG+aphAhzjFwMR+
qt0JMUEj0C2FF/dJSxz0nCp2PorqW114zn/nvc5FOKmCnk45KkdTpUp413Yikg+HMjEDRByA9FcE
lpyYtxlfSrHKxbKOp7XfzbAJZgrd8Nq/KrcWf0TxT/cYS+w76EO2CF1HN+Nm88J4BX2rOIe4eKKI
4zl4FH/M/CrFmmZeGrugtsHRPL1wB9CZCQQIAUmlrvrt6TtUchOLLbNzpuGnineEjqciQMtvg/aF
Cqq6Dug5MUkRMYLEM2vuVKWq3yCasGpgbcBdS9G7fVg81kNlspqhs+D/7YQ7ndazJZsxQ+gWSrT2
9c8spJKcga3rPP1ExpmotgUX3UX54b6mDdiWj9FY9ULtoCVB4fdwmT3LEtYjC/CY9pYKWmYRcOYl
G+79r1N+puhWmhp0I9ug0GwyXm6ApELDdDMbGQljTweiBUSZGnEHCnXD0Mb4M6xmKXWDCQrDZJ7d
044qS3w9hvmBu2asDS/6uaKpznISKJO2ipYNpHbEjfc2gYJDLXOBX87PdkF0/MUKhmU8BEBVZhBi
9LoOOU8Qk2yQ3uOOKZ7MoY+/Ae07ZupKLWFTrjD6DpMnBl1dTA9ec4jTtP8pmZSBnXTUricGVc3f
0pxsEjCiRf3jRcnLMtTDKc3uvD2g9+L2PiZPSyA4wJ0HRaEst2uRP7pnwC/lJRQ3EhXKmL7ddBOW
2k+Zab+MMCvKhWz42iYoJtHM1ltnUaKrV9FS9PepRAWw8AjxYTjmInz1hGKLpN0q6VtcqAmInibv
9lX5PM9/8MZNOumXX2WqUXPyaGpM2Q5UoWc/53rzASE8SFwhKVm78yb6Lma20h7AreVz7nUFWhpP
fvWzzWwlEluzc+dQeVuGz9GCJs5G3Q6Mpdiak3zB/8hPogQt3TBC4hPFelrphHmzRNi1ZJg3DzAd
PhGFs7y6Q3VvB9Gkzr8qDa/cO0ueIvLVzu5hscrIqQ+ZBYAoz5KRd/MDey66SI5Cape9LCG2CGhS
3oQK3Iy0YLZM3+/MpP4JvGDPow++Nze1DYOhEt0L4BqZ04QiIBgiZTcnCQkwsvx2xlMGWu2PiFWs
JmwBjP5jJNinR9tC9tqYId4V3sH0RFXDGr1WXBx1/NB9ymmab0d9U3Dpd0llRaHS8rOqlYOeHagA
Zl0Gl8uxJpwZepAj1LjtdFWg45gkewsSXOIqEW9nJ4QBWcAGlrGMDO/SE7mSg1PIuLgrpGA5AMiw
PeoUILIMKlgUhsVwFn7ye0j8I6DsApm1VCLamrL72c+zgNiHWoiV8D2Q8bIvWjs8/S0QmI1Tv6Jj
tUQ7jPN94qiu8PBU4/D+QmKFolwhQJCzqTGYqn/itjZsSH/2Wbhw6RDCDNALobM1vOwOlefvSUvM
Xx5HB5lXCeAbis5RCYBggPRZQKKRHlm7xDMICyuZ0ZWbFV638bRY7iljKnvhiiZWCuFu0cdwZ2I4
p1JmCk6nNsgTQOXBVJZLOgUtHbXeask05803eSMxakbO2vFFMv4PYkN+qIAErqEUqQ8SYRrv2znD
rec58ij8n8FlSi3+DGbYzwmiwk0178C0TRyqmJ0NvYnku0l+1TrYxYEVA2C9HtBtk2diK18U9wq2
SB3s9b3GbVMz258YutIOzXCJ42Zi3/b4/Pqgu5aa3w2DeIQc1bzox9OmAlX2fO22GMQ7mGHfgjTb
iTWC96IhWruvkwSE+9FH14zvs1ucKsBBTrFFeoPEJcXwJEdd9vpvknq5i66v0RhbaLMnPBfBJc+3
TKokrcC0RG5s97+QUT5bu7mPVumZDoezJCc5C5xA4onwoGZzd1UAeEkoLAFOQznuQxnaoWGmAlio
pMNLQI/0fn1W3H/8WBQEp6FJILSx43W+rAyX4I4sJDWY7UmApGVbYc8peeOKDxavpLty1nLXlRHX
IBf3THTiXRifcM1CjFSWKSfqhTZPNm1PhQ3SM5yKy8qPd2aB8Xfiq+3UYoPhW1vJdGu5ZoLNCnQQ
vSnKoEYb0mOUJeggzgO98Rurf7sJ99lKHrCbLLERRENJu+wrI0K3nSYeHng+R7nnDMgzbiIGpKuV
q4wUFv7M9K/4Np7Eb5CwhSJ9Cg1+ZF8bbxebQhAZQFcfOHfoVp4LWOVPYoHUBL6U3mDM/ivXgl8M
J57vWaxC/tqclsNZr9HWKqf30LGo2Wo3bJQSe91cZBdgrfOCvEvOvi3M4DHgigDnjYUc5a+PT8ON
iMj4ilrzyjJc4gcemFV2VI1dFRpUN+X+PWZEEvAzBxkjPHC7/qxh4vnxQJsP073CzmTHIBl8sO27
zvethF9/bQl5+5oUK/Aqz9jfCzvK1BvAyTKZ4vYhhRPIWx4DrFt2iG4VSIMUyqndHHB8e0kMotdN
0AnMfJg7jOi4ZVLw3AmmbMs0LLapF8ou6v5VbFhtRsd8R/HrhLsxqUw6f3o6FANqCP18BIXcOGuv
IntDg3TpYXsGP3ikBMCcKcfd1+zmXddxKHxOC4kWtYMIbtKbDC5oeKRz/H9hceIA8pu/rWMv54hY
TnyhU5k2PgzM73OKyZycd9hGEDnVTws45jJZJCZGgDCEZxHs2rmumRI4kCSxW4NtKA/mb5CZCK5W
PKIw9iPUyYV0FQYT/8MTieLBLZXCl2vGutwadvE1x3MUyJD8+v1p0oriKExdkNl9zELT4kDGo9JZ
PDEtpO/rE3tVaRT7i/vtVROatwNdkfokZPSEWytOq504gZwtbCsNZxMZnaFzxEysUxkc0IO4u3+W
ac8K67nzYP3LR5qZCEO/2w03SV0+2jCZUl67qSLo0yBrLh71bZic3cbrCLzeQdbQQUNO4/j7jAQb
9Ckz5bsSD3QLrYvAH6B/aCKksZ6BOETBVFdneXxi5Rzc9X37I9EXUR47STQduUAQ1q6n/5lBShrq
pwowyjmscmcYE+0142JiveFWsGIww/Vl0hXLXx0o6qza3El5Nvj0tvAughFz0KqbxUSi+OpFJwvR
WvwEJCP6tOdR2HlSpEv7fZscEgB7mmzucqMo6Kv3YV2KPw4VFDyuyW5fQQ3sP35jQ08dpOA8q7f3
TJEsw0RBOYHOgeJEM9x4nbwoMPVJYXBzvP+4hwbDw0dcN8yOunZYpyG4uHdjoOxa5zAMsZ22qSkm
dI0gprs5WSTnY1SlSwYQ1jWXMC+EA5VIQYwCrTNV4UeoVKIDVCUHeSbVY3Fj9csNK8gWSWCuapeg
zdEAbVTa7Hl50VOo4x949UxEn4XU/cBemwjX8xudiAIARFg9R5BRizAKB+mKA5r/BC67LCmNBub0
LsZQUbKqHZKZGf6HhQ/M+JEM8obG7TQq8mFiHKhLZx+/9eNg3vgUxhBpp30vXRAw7wTh4y2yGUSj
PcGUs60yh44nOWxfUE1LFYZ+yoLrkkfhpNAlV8eyl7K5PrhmOWfKZzR6lqoEAfdG/qbo79O0/7Ny
HxQqyzPJ8SAzwmbxwzf0uSo8KTJzWgt8f4ZYIRKGsfJ2Q49iEWA3ia/1bias5WinN4APuX2ewuFD
LAr+1hl3xceqj9OEmkKneis2z0cd6mcC96fPCemCKsuuxv4TbNfwCsddlZDLhCcxh42agacJU5v4
jorC/fdLYN5zyZX1HJ9iCON/2XoZnZAjbcx7ztSEH6xCqAOi0BBmMpZ67Uh8i4xiMkw/lag/iXyt
Uo1dRQ31UXqfun3ZCZ6p9VLvcHheGsBVcRX0P/zqRRngvhnhBpQc+PMpyj9DgYjqwuv/40awKSfE
wbS2Zt0wLCjlEW7m9FSGOa9JOMWVadBKxmXYL623VqBprHvf7XIJ6DGrn2t7TUlVhuArYswQPo3+
IGekFW2dsItYxWtqYvahdVQFnKuGVlcb0Ih0U3BGgcXw/CeV/JvEyLpG+75zV8AeCd+jNQ38hYip
iFDroeZYMfRW1plkhxrkyNhiu/RrrXvq34kciD+ndNnFMNK9leBQ5HWAl9tZ7fJHr/VfEBS3aiX/
+QCDhaYwc7kNkzofUHtSf9CUhjc+MfRkU04uFuxl7HUbeTqoCzQB6z5vuhfwAL+YNlQS4sVB6B6C
co4RQk8v/zEUoI1jVkNHZXJKQkscn1zqv4nGthBZ7870mdHAnYOHMacSfb+O7EzBO9C9DjNyc818
mZc593opdUOdsmYYFUueCS3P30ZmADFnlnnKbx+L2ygHxWjLAqT6iiHjilUptKoj/pwGogSRBEKA
HUdQSkrjP+TVrg5ajzFNf31ni2l8Le7PmrQ9Jn8oJRuJ/FY07X8vbzYHd5gKWrBNTPKud1U6FVHr
NshgvJY1cvAzjybuH/9RVStXIlamqQmrOCx1EL82t6J37W8E6SXShcGdUhbEhnlDwBveE4G78bXb
29sEa/ipUCEv+yM5cMAMYGjDf/LFV1xQTY7BSr7ZnDnInWEUse8YdsksYpEh5SMZhU2rHHFBJ2dF
/+xRATwotqUjjptu8Wp68TZqROcW/teHwsH29ijO8nYYgNQiWRn3/nhDa7i+fdwl9UM1BQekDA/v
pFCwZFKl5HyA//rMcZaSycoeUcMfW/3muuGmGCvifLs0bDTQTNEnI0hwOlRDaUOI1jwHmrG2lXXH
fDKZutxR030Nh8EG+dSlpNF+yO37HKSl0fDVI8R6WaG/Utng86J9PHD0gMGxLwKRjAdnVQ3kSwVZ
BSzLvHjJrSO0wbVcgTHTnsZIaHCBTKZkQv+R5/vz/A+g5YmmQaaVqqPsoR2Cl+N+dBZhtdx8XFpV
PR/pTyS3thPxygNMv2s11IsEKLWTeNGOF1UsVcg1XNKzOHqgsKjrOtV+nbRE+wefu12kV6M7sK05
R9cECGIJwWjaiBJseAI36e5gALjOvP9cPivW/Nk9woCzBNdSXwqYBblc/7WPMeWc+F3vy1E3KKrB
Ta9GmcYPZwnbtc/wL2IPciG4xielQSCtu037L/mU6TQ705I2uj6jhJ//0HnLCbIofxwbbXWwkqQH
WCak3/1z6PZnqf0h5cqT6x7zSewhA7mfWYj0KJ2eZqG8rUr/ak+kyKO+cDu8sW5V4VP53ou6PraF
ZlVxj5MHxJtPExJnZcrSHtBXkVIqUzKZ/TV8xHZnIUa43JWBZMh0nAMCbhs8Qfv9m0whZ7SBjhJX
znN7D/AklFmtwuUoCCmug0bag75300qor6Z6HASGpNEBG1s3DCzE+6XtrhD0L0+JjYfXM9d+5RqH
Hfzhq6+0gv712pyvtR2nI3FH6iAooWCzl+td3u18XXbQBu1onum0S8Xzk+Hke8g9vMhGjh0bpK//
OOzv257oe4eVXdIrN5Qctq6u24C7Yq+BZJVWd6MJnFhvkY9JqevOvcBNZFNyoOFgDhUGOO7xjioe
OQJOgEJdPrDitXw6/d/SCmK5PsXQ8UX4mWpKr+ADTTCootb9LiNDhzDQCEUYd6i14w8W5ORWfOBU
3347BakesB9ucp5gaLk/fEPt6G7/32vilYEz5P/ji/z3m6EF4qQ1o0V82bencaVXZ4A9QrC1hIf9
sRF8nXki4/sPGQKfc+q3ZfpBCq9T/ZtrpLndgAXvzH8KS715chbKp6muYbP6S4qnbdtbHCddNyjf
cw13wHrc7CCyjOqie+vYG+gOhpE0zxzI5dXGtIUSVhY1pbNxR4n9lzktvrbn79xQfLGhh1y9oLM/
DvG0XA2/sUJyc0BdMCwNvTQgOBfgQlPzxmz7vctZfbnVgMsPhA+/B/m6bRkfke+undhFO8qlI9JV
Ud5P1HeoQZNhc3emiXuBCpiuqenPeIMcARH0NqbXeKSZtCHT58Uv+EniwjD9bVey/i9x0gkveBP2
RTGnKPZQsX20TgBWpomdkIE7cFzr8UMVwi1BDzQyflsK37pjFSIBQis4Lsz9ccRbfo3EDULAccjM
68PhmMHL0qUf7gW1npPN3P9Pqi4DPSI4KtmWvg9zsLB0aSYr1vSHusFpTOcr5T0B4TRXLfRepokg
0KpGTjnDGfIyDlwyh9FHQdlHPlTa8b/e+tMC63eLvhugzUAGUH0Lg1CBGrlCFX7QrYmCSkQC+s3p
CraY0xI9Rb7tzZ/0676BThr3atp0gfFeN40tr6/kPce5VFMJqUHspLn4diyIyX3eVB++hTGNYPra
WLwiIXnA+mzz9R4GXQobKeLfzyMWWg/07B5kd1FT9hYrIWMIqg3UPYwez1hkCLc+anWkemzLS71v
odnRaceFiW+E74udQSo7iFwvbyIg2hrCPHa8t9zjfkuAF4dBhR/6bl7nNt0GKvvSoqCaIjEBCDsg
DIRo/J6q+XmYSpV5lCGIvHvVPQnehQYBq78RjYVw6FClymUJMdJsv9OqOsiLEx+Cp9tcsNrkNKO7
uXCQE3Lp2MlaWfBpxb3JPUCmXtO6U/jFaCo5UW9vFL0y1653e3fP93i5hZd5YSrKk/+iqgoSJvwJ
DupACXzutn7Wfg91WVmASZgsEz96qAXkJ71nXG7+bPcbCqYLzoM7zF9N7n960sKxRemR9UK1oQ4t
yFlfA/N4Yv1pH8tLsk1vzGRCQrMF2fXI6g8ZYLft7ATJ/PBTUq9cVHXa/qY05fNqcz6SKA+HvzsQ
OQj7neqhiZUQbvEnk40E7aqqr3ptjLUdX5WVY2VzOUEJ0eMTt0TDZysM2S2WxqL/o1dBJk7F64EB
WpPpdmV8VVT/vV8GZFTawm1WM22W2zAx90wccm5/hOM29uEchX6yCazwNfJP+4+TFcODIwrTyDJ4
kFQvW6cjSs2QrJJhy5E9KQ4KrLGOKVPDtWUua9neJ9HX10ifAd0Ai7F0M44AVyVkzS43WvPEZN1V
pYtqbyBC9NqW/m+D3PJs67Ww8J/6WY2ewQXDy8E26aT5vVmGPMN1DJ693Ri2XWqb9RHiWmbWTr7I
q2z6z2p/E+HXVOiQrHa8r0Y+kPMAbg+vlEl3KcKrX3DFWCK66nnV+Qo3eHYxNYc3KjPorkTd5qFT
hLzPJjgI1CD3T27LohtPLW8+hjUx9xm5gp0k4RN/hT40QUF2Gl2fPiWlpGlNWRcDA1KtHPbyOltX
QpUnyaoPiEruzYBMpT8VNXVa3N/tcqm6L11bzZ+6Ys2jzCQ8nzfN7ICyyyjZKKdeeyNMpuRkGl4M
OY//f9MWswXfSuDBE5nuvrCAMZeZpGsyXJucm6oYlKsru0tqRc3dKgiNniEixPUXThtscHUZiFPx
SUcNLmlIph2xtyLilPmSzVuFzkzqIbleDVBDy2jPug2OD9PvfIQUBRl77qAVyn8769skmmjAdydM
oT4pl2T84QUyaZctrZsXXC9qSHzYVF2Y+wRB4Hmxz8xQ9w3AUEtXSuSDSBUPn2fPlnTnjhkJyPVl
7fkeSGTKueAbLPQjqNj+2Y4IQeH7ptGNAw8prKogS1fSnxKlSzGDFY+B6kNqcnFNaxI2G7LB4r+2
abTmWfFIxs9JgqJaydHFq/m4/Us46U5E9Pnt77OAfqsZit+s/x9jxo7kKNYiaBgJoSkpXWVhCUHJ
yQlbnjTFdFMBf7gzBBQoMN2WXLF2CFYfWUUVy7UpQWv8UN/JtWS2AW69dynzv8AZi+ebBmOhPvKs
hG5b463AMaHUaydRKRuR8Iq8+3rlAazNEGkGIZQDoumZNBLH27t/TYd2en6twCLYPH8NawNH2b6h
GTJjt2SnP2f3oZ9PuVSbeejLdie0ZbOZL0iTH4SOxXN/elmy2Dca8DhJoYcrHJPRibF4LVhtRr1K
1uT6Fgrr/J3s3Hais/SATDn/tKn70iwdpBbk9KGzQOS5r8JtdhHkyoUafmJ+dg3vC1DHyq2Z6vrA
MjEKVlzRtg4nEdoy7lIO/8vLT+Z2ukrAa5nJXexaRK7eVFA9nZ/DSjmZFZfpy5B0rfEVFFOxrluh
Xp88GODg68BW+tK7qVYv3j1iD+s96rRZztlSv/K4AVlT4VTsLDNLi387gPb0vZrucamT7kyBk+6g
47SYzXDEvfpuz3gMsPsfvx95lVE0rwQ/o1Ih6bT0uJWBo7ztpyJ/s27+c/1E0UAeNWtmjPh1OYM9
qj5A5t6rqw+RKDEVxTjPUGF3mljA4epvQnNPM793GApa6eQHCk6pyol5t21tEv3A9b9epbav6gso
dw/dXM12j1lXky9ajs7KTTc8mGzuVakEpSaHMxFqNz2rwu5csPTz6K0ZD7EtGITtSzQGFsnhpElJ
8wU8MvGuS1r4yE3KqCqX/YP1KBR98bh3VX4zB5fzPbazGNX1WVKquKURb+4zFY6rGvQPUApyEJ1e
GVzc02VJ//t3yg/mdhMzq0BZNwcYBJsOJiB6XlTwDs4e7iAzJO+pQ9W89Bt6BdQYZIpG67LB0pWl
qh+9GsPiH6VwM3Y2+UmN7USpUkfisBHGFlzmPeqTNeMvbq1M2S8o8nhlEnYkzyv8iTfLeNYpDDRs
LpG1o3u7d73wz2dRG0BL1O4+y2DT4m9VG5990wiL+4S8LlJT33sOwWB/U7r8N8rOW0Hr8PDZb9Fi
IG3F5nnuxH2okdTjDB/Fh8rKk7r8JIVsQTQgvLk2zc5L+fqqNJ7MlWTIVjRxkxI4UsOjgw/nE22/
nK2UrzghLcEuUe7BoF29MX5y1hm5wptoWgwm7F7wWKJwtaGyFN46IRFI6gbbSphQlbrMJAmj6ko6
ozCW+ZN5OA5hwhpkiBFF+6C+KkR3NdbxIFnjUEz3q/3zDe6jqzBU3Cl4Z/xT1Z3NIkEo+UP9JNcF
SbaOsGP8RkqBxXUAli6IBoZtC53eqYlkwccms7pkBB49ce4j4+TWgnpA3noiM2BKoQ+baT/sQ8GX
uyHaWrCKZd+Bdtb9JBfmxG9V4jvWz9QyC5FB8rVhszj6IGh+m8WxT1mXMw2AyVWVJQFvoAAGrCxs
Gl7REXP83uR3nwjZ7Sq1jPCA40py2EKfATGz203LvclUWIhTA4nqfpsSqifQrdI1wfpeJjoPVkBK
U8Ioj/epr+brYoo0HU+q8mlITUDf8hNhqlhaQ3vPMVJZb7EIXkBZVVppcmsyDpJ3BJkAb1VWd8z+
3DmmS+t1E9i29IoAGIPWMkmIHwpCjH2s0lUH2dEq3EhfTWPdQSSENZ0b/zrZdIxsoTxvdrszNbgL
+U6QvrnUBmAr5cKWtEVodK3d91eByoLGFz+hQ+tyPPlD/HqVcdKOMI54+iZfGHJ+3mEK1+bgja8E
bIPumcugiHn2354bl+x5AqIEoEXAmj6poYRVLflFsJeiirUxWNOLKOC8MPX69p5Oe/enckWS32qV
HjrtvCKErwNPGFu7EtsQy0Zg39xxnP4L2RIQk7rrO2qCnuAmIG4cM8i70aDO2HF+Bb31Di/AL9PA
wNAlPs/tVLG5FWiJMmjo262zSf51LsOdSms6S51chwWPZLDIUw0qUR3QwKcIrK0DcRjTqndGufS1
gi+nmehfuUK09CetA4TvvzcUEC0UVxqMRsvRmkfFfA+D1rNNi4Ert+iYUh8PCxGTPdPnTWLet2ik
0y+G1Z9BZ91cheShMYkMWktIpXO6SNijvc0Oy1GhdKZ5jEtuua5FCqHAljPAGuKabRPZgDtwToSu
enI4a+oKUXJ7nf237n3qgAaXEtfz6hT2a+LhNqJoVho1OrqEbL22bxrLzy6pL4rNDzoFzKQDDHyt
sDuCm0CQKyWVXDltB0S7drdtkYNcmqjhxK9M/x+08EpjG3pzLrAa27Nq5lMNE0Zf6hJC+RdYUVOo
+nTCRTUnX0A/Mr0BrAgorxr0ScojW8PSlwMsewV6gUex8ftlG6789uIuY6zkd+ZT7fVBRsEnjzas
3HW8Es/KQIQugNLaVa3HVT1e3s3uaTyOV5xNDsEf+Wc4WN/gGG7CRXW+aSEVm16q68BkebTIzSQE
QDY52k31VCp2cya9jCJv6MW/xC/XlMJx6F0dciUsV1D0I8Sy95aS4dmOPiUSj122f1a59cXyMhRp
5vYdW/slzIkWWyMF3SPcbgs37Agrd9ZHU5qvGvVcGF4uaRu8w1XFP//0Kml+NWo+jBsw/asXNRcu
suA9HfdI15jms65TcPBfnXPXntsWeg+fC1rUUAYGQXHGnt9bjouFiX6ZNTcHe5iRe4O2SLVobCJM
0HmG+mmMtXWUGaa3U+eYI2WXGRDBTvbhFAM+MC2r5oR7r/Z3qSlb4eapFZKu9zTnuJi528QKm6l8
ZCviCDkOFs8FAGAMGCnU5mFv83/k8Dmx0RD8ym+Xibd7iGDHk/M5p9HDBG4cVDL7ZSmzzOQRHbuE
HCQ+eYQ/qNx1Cl/hYwx/Hsmhhb+C+ky4HQch5Mvh9lA1GNEbx8X3U0L96q9GWEc2i72X7dK9I9tB
i7bYOYkR/7aBUo5lO1T2EaaVVYl/35BlUKHLtHPJzIGCTTe45hNxkjOFXgoiXL9LbtWoSrVNDE7T
3peOIcAyQUNyTB8JWPKrf7IY7JjOS7wpXSLwfeYuRfK/GD+9+L3f3vwigOcVG1isUIaWEVvs1zHC
p4AR6/RbiDfGggq5C3ZpeuN+Lol4Yu+5gdTSFgtEZcLbqBIVrAGmExXOUpCSSuNM5R1MPK3SVg28
x/7KulIslf7U5MHj2F550x88pbyLvMWzzDcB6OKy/wHLc9QNS8SLKgVoi3RRDxzxJv5msebdBFfe
+c3HzEKy9Y38LLIyg22JtleTXeVLlGg2KB7I28oDlz6FD0n5ubR5EZhrSSc7ojzyoTgS2uncAROU
gD38mUYX56aJs+8XKUomyp0hs3OiG/EADPZkJJAUQShBMrD4QIyHR4ZkiTstXOregpvfWHwn1lGM
fDwFS3lldM1Udi3ZQi9qriP5X5Sr6mEBAiJPz3EiI4MPDnP917YVoync+4rm2AlK3z/VRmUmFFi9
TVSw0QK0pyTPi1EtUeXoMNGm3AP6RkWBw10P6C5ykHH+StEX0F84xjja+ffKMfFltnDakB0AKAzW
HpmPH90KvSYj5w/01neOfAv3S3vXmsEBMD59Oq3Eq3Lc6eII1O1eu48+CW+3/+ZMqSBMZErRs2GG
ghpXzaVz7akHQlKnY8UJSk+GViHWMPdbvvPmeeG2tkOhN+OfvENDf0LGFFItc+vgmdu9/A86c9Du
zRFT8irbwZyAHJ5GWpflOs6EqlD2YTvjjs8e0g8ETsfDoblHNNWzlDiXRK9Mc/885d+wwLwJ6lUa
DpY/sIE6S1NooreIFknq83oR84DYIl0NfUD9W2oG1Xc59aSr9EclOXgIt6AKVDWQxZ8nrwgoGEUA
mAYmWnvGWEGQCxCpwgK06h48hMPoxC4czqW4uoo0mF0Ni6iEDpU/LSrK8sS8bP6Qi5KBH55+UOYs
Tdd0YT5Wrbwl5zFVsvHqDtYukQw404YcAHPEv/JU5wIZzAgAbjlYE89M9G8ghlv9hzy9zfm4mWXQ
IUu3MrS/gZaoA3GGrKMRKrajCQ+mXNFGzsu4CXjEljbPp3qaZbYzfE2m66BHXH+R63YSJoLbFVWm
6rRoU2+dyx2rmNbi+QDPgReDLDEdgWbQUQHDlVwhX4EfRDlb8Uuh1h1e1J8lTpXvZmuyuag5gvfx
1Gczufm6mZgnCAPCk4holoJICMYUGr+14Oz47RwMf6FCNpoRWLGHhVJASqPAlr7GWMPmKeegJo92
Kk2tdkc2++lNel78lTUal6n9pG3E6H/PCLqd1hlOzRkw29p1rgOgK5fokEv9cnwU/N/EZftcTCl1
miQ2y/ycSmClhDsfyJ7bIss+zizYg/GBctaN55w4iC1e3i3d3kl9qqwlkxkC0rxwCOgVQ714HEHX
Z4juKhN7LFAYvlvR0Nf1VV6zAlMCCcN1IeVs7e2X3+cWsX293dN7swjF6sMjuxFQ0J3CeWjSf17V
ri7EF5KcYAZTnYip2y480UsYjrJW9jz+/2GCWNc6VGdeRASNy/lTswjQSrX5gDvHBP9EBuFZAqeR
rR26ixUNGhqGyjqc1tgbo63Yq5svA1yDKePKD2v5L4XqKXPVXxfliUJKn4ncqah+FCGFyQpIlMns
xw2m+oA5T7PX1I8J/1WmBAHoZx06BjSo/IAVBtP6y0cTtuYYnpMwOy98bW4v/Y+mvuvgCDR1Src3
Tpj1e38UsrJuadOv1H2smOAH72gBTFkEP/MeL9jS1MFFf0U+vpFPDmZOMn1P6Id3JfMaBkaER7xo
abxnZjbYJvlVvHMWWXEZpMwvnr71NuxKIt7LatSWMNugKQlusV0UxshZV2Z5Lr/7jo0t2NItYD35
EAO0rptmpDeLGhAkeEBQGi3pDWXa/I68FYM3fbw+ioyG+giKoaCj6TmRnLjkpztCr9ZXNADol6A+
bT1AkKIHwcE4JnWUc2IficBODa/vjrKSOkkc8RAMMzQfYE9wySgJuYur/oiusTgzLbrQj5pIdU4w
M2aGjG9fuf60tZtJUWDoG8tFmtDf6teVCF5DN/ONC4ESbmmssdGjVbDqvan3279yxL0U6KY+OfTc
jLAl+tuevhqFZVyIIko2y+bavgiwPnmN1elN96162wH6FrVD8n6YTnzxXC8AfpfqJ3fwLSR4Httj
Jg7d80zpvmKpRAWVZ+77asBbWP+TL6iZ0Y1LnFzOQCZy6zcQqusAvbqYkH+UHGcuD68tCjQHBrMJ
5MtYFsit9DhHA+Q4AS6H+EOSyxZzyXkbnKF6oat50aAif71J4CHuxqbxAceHI07Pyk1zhRUs/NYE
jXMWd9kiXpovTd/q3iEDne+Mg0eWJDnbQ6pBwhgMSfXTMia+r+SBP9sJG6Gax+tcJW6eIq7mM91Z
hjgSeUiY3wO9HqzFPtKMOlFd8jhbXJB/owVOfY+KvecFv6agono/Ia4aOL0m7akqV8wHAQ0sc+jX
XMlpiCVgvn7F4OBq7K6RNTQdtJf4Gjvr3dQZ5QYgdkxKE7BFfrNG+1tGPRNVPkE684yWBtXUQP0a
hRPloW58w4V4V2HwUHSwbcuXDKIYUa+AyaCS5by3pwTQxQvHOdJzp8HBKrHNLBsZq7VtrqoNw36t
33129hD8zoEu0r9IMdGBlW0bppg6bCWXNkixqP9kMNxP5tKMNq4cGY/ZKT+yRtZFVyUTdQ+PG/bz
8ldboQoMoeqUjzvDRKaTf++qsoANk038u3KbGS9SmRXQ0yROdxVhAMjEmfF88Qkg35kjg8Ts4RTF
E3U9tuH+OXU8RIGzgzWFTIj9IpEmKOwEahAyNn94TWO9awNqQJUTRgZjuDd6QESSFl4AFhQujU9O
xIs2/Huz35vZYDv8HrWcqfIfyugMPRPRGm50kg6h7z8WyLOISqOJai/p8JJG6VTozigVNuPlWaEU
pOVX5e/tZpBzsfaLtFpC//JU9+oPjfS0bo7LsXa0wHfCelwKnLyoDGkKgD5W4AjaTQE9FLt855pp
IwGXlhZTA+LOEgYrHdFQsJctyoF8fHbtbzSRY6oAFLL6UcGCRYMRC4bHFZZxpwi/oVwcwjGyX4w+
x8eKpPeJu5Iv5N0GPBNm6oCBsswreNiokJO+/6ksA9i/ktKV2/xLDP6UmXmRvXlpxG/gScWpsmQ3
1U0OU4jKW1Jw6cGypfJovVb8mN1GSIjlADLjbJ02yFGqG0SNPckarby5T6HyWeZO1jzQyJLxk+ao
n0HnEQjj9m0msAclivt4awXX9C7xEKTNG9L4E3TqKvd6v4jXbvUDKkyAGG8nY8h0LKv5/ujawfXu
LSTMRFPjagY7MLnbKw0bNQejTblQeGw2RyfV59Xdd6nVs0m4wPenDzKdbAtXk3P1YoMjHfSUQ58I
DWn/CDgu5GR0ZnMOkKKM9DJrhgilyWxouexMWZcGkFR5hQYpqLRV7au986Jh92EZ/D2AHVqsGJiB
wji1cjqALv1Hf99IPbD9RcSEIqHt37avSbmNLhUYG9C0OmcPevLGMceECFIn2EBm6HGQPWNvBC6k
q7j7Ap41u5eYn2PErbH/3tVHoIH1trqNA3j8YIG6iX/LVzqZcWuoFiKGwL5QI3sf+Yk0NlU5tjhn
6uhWr3oEL4A7DXHuZRfnuBedXNvXq2kMYoUtWBnArcWIV9uAGDBfoKaKMuS8S1Tvyro7v/Fz7jWk
drEKga+E5DRoH9wdmTYjc4QMu7a+irDR8+7lOK04SrLoCmUecDRtdy96G6ESOvLoeMyXfFqrRyKs
uBfD2P/Q6ehSPjSF8dNzYNQBza4Pfi/nmHY1U0AcmIAXVBSsu9obwPt/Iy8brap3jCJxbcJ2kzBv
kVmwMIvR4Kx9dfrqjts/vFrH1u6RZjjV/U10KijEkAzGLibGUk6xd3WgC9YufAwasKljROauqIjn
GSz6MHFqkoya0ceEJSHus+J2JT0zQVVEM7uPrIxvLYtGclTscQVti/riFL9oQubdCZaH0tvoOTnY
7J+5qt3Xu0Y3x8o+USc9tHrDMzwzJC6hV7OGN0EXJl9aFjaVc71ukE5lbEY02uC99tde1uWUulI6
LIjy8DnMGE0FaRNlpAb20YnUI+sO+vYIwYlI+/Gx9gw6NV+E66bNqlRkaXUCXV633w6Qipb8f4yE
zTynG3B/5XkPxYL4YnfefiyCuRcq1j3PyYHGrGvOUbSortmrvpMDl/bPkyoBL5KauIB3ydes1CE6
tgwuuYx2e5aVsmu6uX2KzUrgZr1PinKds0oZa7snxOydfh+OM1RCxpRLr++qAYTcwla0ScLjyAj/
D1wD4wdGBzXGJqAzqRanVrJVO1UztgLP1lfyhix+2tooc55J6mB96LqNXHntoNQP4pix7fpryrJ0
5rr1AAvisn9PuI3dV5mDsNSz81OV1lplxdVOPdO2iTTzIEBdy9r5ZdMiMZ9GiqwHxD0g6PWrwcUE
PkJYJnxQxhp7gUq2+rxI7qyaaYve3sQXV1QZpvXIlXxvZeAnKEiCdBctoyFDRGelp9JHGp1b3n0c
ie4OxZmqpuJf8ZVg1ifEO6nt2BQMvDNqOLnc6zJngh7IpfVwsYiW3B0MAY6lZz20cBCnMP3MIqxi
O/zI6Ku9uFNdWIlNaafU5WEo20Fl2pM8zpEFODfZIWBEl7Z8Vt8RWc9XVFGYAroMXPSQOGzV+oGm
HX30wJDRueSXbvOaGM2zuT76++C34VNGrEDohT/rfHbBqQLpkYa252CFZXDB7YzReBVRsRltJTvu
5XYBm3ta9H7/Mw+8n5+VFzAmFMMvZPO7sxFQZPp9VHBSuJ20IzyMVPNXTHxLS2mjo/7CV8hXd+OZ
GbS+2RYWWk0JsEIZe9pSNiyFkyxgKDcRAogDl/MQA8B7JwlcsQDpTBQT34LF1SxMucsZXWxsY6L8
eH3fqEiaru0iVmOw7OlH65ygF2S61Bp/pBQXd1ft6Nqvlhnh1yWXZv94rOclxncSYl9tY50dk5A8
veMND920bOntTnGa8wuZSJ0Ex/DqyIR7XcH7sd/045IIeXrY6jK8Az4vEuJPYD8uCD9kZyu6sha9
tzSiCVw+F0AsfaH/FlB1WdcJadUQQn8HaawH1qmeeClH7bhfDsiYn56ZFqnKMQuv1FJsWAGbipn6
lg2B90K4Qg+pwbVGkp939Eovig2IELb2pVgElBKM/Y8WI/5KYPnTlTDSETePTf99CnVP1WqqzLDS
eyS/irnODqAElAGI8KxJaat+BNakhlDE6yDjZXMamVNmTg8kfQwaJuLzuePivh2S4GOd6/78qX1W
jNe25w9j6SVq/HsRrtT5f8ud10nEjqZt0cZg09PPUdfPxfTW2kXo+h8GZc9yhX01sOUHj5jsGNb0
5EiSO9f8hCyI5YYew25SJmV//H7Davllbme8Vd0Tf0SWpMKSqrBAAPgENIcidvi9BsuTqC+XoR37
BakZu+leCgE4axquIY/j2XsVUEAG0Vq4i1xlbavsVDv03h33zPv1hVxGDQ/mfYink/9LvgcHgW29
8T5Thfyb7wHbaxbv2v1ns2033M41qibk0R9a5jwPtYzTjuwPvk59zhdrrlQM30SXzW99dro+53WQ
wNatDzHtsdM9w/+AkLaYTs6UsRx4FWuBZywwt0zw1kHyOYkBK7mRotNuTIYZNrg5kYzSe333vPNj
SjomzbEe9d7+yuh5UzTlmh7WKWtpdtObLmnwTR/A+qRzll0j3ut/Bfpvz4KKTBoy6w1xdtlz8wfs
LBPiVpOcqZjK7MYjS8xur/DvYZhn9FWg0ZKt+AFaFoabhGiOiOESaGe3lDsRNtIY/qzFpZt/l4kz
i8/zEOeJGOp6NYoBYZo4ZXo61I7lbPu4UfWFRCFbKyRgkWRC7N0bkuYnIhaLJxteJzVjwmpKT23h
xhvr53BUgfRewqS9512uJ6aydnjzLrQ3UeuTgz/CDCyZ5IX/lgJyLrW2ydRGkKCwl74mYM1MZZ4H
koVaGf2KYppImknRcI3Gx0ZfNHwOvhZtTgz0YXejYsYxrWpKR9jfHzstYbpZs7OrkMe5zdWRCGwo
8Ur2mnRquBfZsh4w5hanczt/C2vwU9z/1p5AoNA22B9+qeuJ5YgNsd3ULYdA0Yq8kKidKjAmO4wu
r9t4dmB7/Er/fz031NRHPkJkOxSB0uPPmNt9bgj59j7Q6lbRA+2nHhmHPLp7vAFZ7h5Q3rekAu39
3WN1KeO/Zqo8SiMoptQ3kEGIUAQxqyhhFhD+l8PYA26tKPK0tkyGQaLikXh7+XyzFzLg+/uvzpn1
zvrQ8/wbG8SFaG6QBYxUGC1aVw4Mz5qaaVVrMRgb4+75pw90I5d3S4xUhUAEV3Ao210lHYYn6b70
gM3VVM3To/YgjrRz63Px/R08pf/f3TCiccz+4swRVI45XQ1w6iv+42vATeRhhUqx+8L48XUQfnpW
JE3VEZPWlNwgeYyJHNg5GvNkH8UuY2LGC4sKl/a3wRHUufr4nerTPxoKZBhYa1KVtoUXTfo5Ya15
m6EK+3yDB02WuxTAtKASCpFRcAI9jz57AKPUt+f9IWA2yLzEhZL5piatopJR/Of7iQ4hDFD4TX4C
o1bmjoHMxjtI16SYokjS7woKybRxjgSzyI2b/fzeZGokkStSeG1uQj1lLk0BX+O3RSe5eBIcp6qd
VWbnKZdyu3by9euoUMan7QHHl8Fst/OETC/jiBsut9q9ohOlGgYg1wpN0go/bGC2Hz73T0r3LT/i
F9zHIMBW+Ng+//sP3UdzB9ooVVwYYxn55YuaRgNTcMvus1B6uBeDBsUX+sxsb2+kubStO9Tn3VDe
Xz7RKXMxBMvQFIf3BxT7VZOwrucROvM1NVvhfXZJq0PcICyFhbsVyD1R1MNXlJOSZ71TKCiRtyVO
Wg64ap770ChhH6MJPvKM4NEzDN5nEm0LQ0H6/WVlu7YwfSgiWK+0PW8hcR4jb9jh2IxzHL3H6E/F
BFAYseBmkX17gi+lsL8rb6kIJx0FS9HDR7jk/zuRI1sVvoeHrkwOp80WL7YZPNJ5DiR/8ltx9/RM
HBqGDqhhOgb96io3Su5CrBOFmUblRztEb1Gj2fqfspzOgMEySJsiIzV9LCk8LJAs4SijZDqBFfg/
TQNTVZEWxNyLH1WUNXqjxsL7XXGfPb2sZW6rDstffdgvNvM/DIAhs//9pGg+GpXxpJuOdKBSd5G8
6vNt8hs4//lVG9O+SMzx+wUVu2cm2+d1XNuOHIHysw1BWabPbmyApOyEOKy6aTh26CmRwF9Ezf0I
uKBHS7Mt+FAFeIhvdK6p5akD4j8VoytLUprP60VYb7FPoWCYnHUmxOvdCZsBPlMlnMFXPxc90li5
PzC9lU80wTfJRfS8XNHSXqTWv4h3DTjKOa3XUoNwh2j2/vw1ItvZ9/cR9K5tWZzsC+6LJ6B/Hv8g
e+6yn8gcSxZXsYSRF93hgX/rPkiLnUkD1+4QvNgCOZ9LQvQIgb6ziIax0MFMwhVtBmlDeBAJrLpu
yrJb2Jx62gA85R5RYf9a/B8QgxRh7mFHOYCefmFh+Xxg8fOtgEByCznNi2j1AH/PLYrb6o1KqRqP
7KIB7xnPZP5ezm8x7vm/R81oXsRpUUu1NKKY/vw9R3AsZq6PYPkLO93yZuC34PG3XaYigVbhvM8r
RQ9wyrb2zXpaGYxjuE/vegkB+0nxMxvrJPPs4AQb7TqkwNzOFFtp3iYT4x4mp/JbW3c5ueC66fNr
EM7rTCEGXkJbWcf83mxHoIyI+2sljns1w0PL2bXy0Y66x/nMgnHR6CENDkTozGuu/NfZlcRyEfOy
wqjtwAzs+CM0EejLPbCV4JxxMuwP0cDqfZU01VInMSGWCgsoiqpXPPQhaus6uJH49My9zNiyVNZG
l+zHzE2Z86FXWaJEoUy9abZMZOjPSjae0NRo7LsmS3RKKeYnwWr1ueLInYWUOUm8Qyhkm1QxdeHJ
f/7WaHu8TieynAlNZiWYUsOtXfFxhHMmfCZQMRWC1943IhgxbqaKJFXqZjH3x0za6wnJizpF8Lfn
tgtL+Q6yevzDdovKUDL2bv2ZS/3njJ3AgRrPdjl/cPeYFKM8WtMDSxmbZoKFeDRLiMlp/bLs2aaA
QjIuWJtZ6K/btIdRKxTbTC5deWJyYjQOudCeLfHNwIU2tVBfqPgeh8wYYmAoibAMjtN4JarseGnL
aWF6en20/Vnjer0f8il0RD+hoPesU8c8SvJw9LLaxXY6SdY9GtexWRSNP+/3lImwFw0DQZhNMzai
wSNrnsrlJg4TsgyhtuqMNqR0zKoPzZezE6+SxDF0d88NJPDhH6HBZD00HB0+qCkDWJt2VZCGRh+g
qG/aj+gyMrEDnc8xW9VRC3cnAhJwmFhwefZd4ADMZkxxvfaZfs2OwjZ/SItq92Fj+HmsQOO/cFfN
7RyrN0CSkQV2Nhz4U2J5UkAKmHm5yNXn74y1hYTzsaA+sZepH8smozfNi/CAfEUb5XUap3onMK5l
YVBreNUwTF8OQ3YoeWcDkezuFr1smRj6AWM1YE0z7SqK2uvKfljne7zVo+UDYB2kuGZjPDGUY38T
gUJwoUbFG+pq7jBH8vuK6dlyIgJWvnNEZE8uV7C9LgYp8cudKszlA1DQAblVZCC0ejCRc1AzEB0l
6bfI/TUVBIAipkLiZXPdsrCl566mBlaukEak9r1VJ3ccIrPMu6Ve4QeGQ402Msq8po8wnNfFcx18
GHEgBXLXKKv30I7FNRK+mFlUnYhNKSQlTJQcpb8R8F89AHChLCAVb1xHWLKDItJdZhJ6aJd2PwlV
1YH9svti86aevJDdZyKyc4EUjzcGrwdGWHILAipjoEBXDTdQ2N0mrj6HPHa4s3VN/UjRxm71zotk
HCiySOw4Pgv22Fv9rahWxmYWBwor94Zm8+Pn06qOnRmXjmJlcHVoS6BeA7jB0yECSq3NTJFvJILM
t0PdiwQszQqaD/cL1Cz4XdMBXG7hcnmwvP53WIaliLqKDRciEmSCw2GkJmEps1L+QvtZjnHr0doV
tzwOKW8T7TAYrDLzOv8p/gH0iYvOIZfMU8o+iFv/QDmSuo/SI6VPjVL5gxfXtEhB9SWqF8aUiuk9
HFtTKq5wCQm9hprTxjIbkicA3ZNKcOKjbUS8F+BWT1vDNRgUqtUdMQvb7Nin330KS5K7/5yNASaU
mjr7awsvRMrWHBc7VEOdrEBJWzTca2oey2YjplwlY57UEIAOmjsTxqfvuy3Ilr49Kk8YSC0v5jM7
M/GcmjzO83y/fF8FRqOh3Fdwz2jo17Y967C9fv4h7+CepbOxRqPHF9pHnWCMeIHE8x3jnYk5j/Vk
SelUuU+Q8Mp91mxRre43A06WzVr/zFUibPqzvIvEicUAwkkYLM2P0KeOyybjTSJKLPgPrKUS0yd+
+IP4WnOsyc1WWAAkX0x9cHu4jbaDLLjBIaUZbeqjQTIRkGZROsIsmQeghw4x5FsB3YJWneF3Fauv
QhxjmQWLG8py0dPpje1LZ3nC0sVjhsskjk9Q0HhEtcBqd0EwAbO10U+0dRoYDAkWgJjM/6CScYXD
AgpuBGeobrkwurcxMQadWHXWxPPZ/2YkNN/JlpgFTLBktDmmaT+CETsdsbf/i1B0DT07BXPjPVdh
uXJexkB11wjCF/neZTPc9r6HTnPillLDONuxTPBpe84GGBWhkXf77RXBknnXyBbUC/vtMFuh8jN6
fkTEucSFBpe3cB/uukFJZ8udH2brDl7QOCFyn6M/OrIFp8ekuoGo+f45muQKjoZp1DhUcftvlWR3
foWszKK+AXXvKp5EsdiYP39iI2LgH2kEg7tHqXTns/nXQrDFeuSNEmh/S7dXHK25i0Wz7dKt/Yss
uGnP33W6qxD3vf6Vn14qf0X/JLsQBm5Ed3AHnh3flNZZ0LO+f/mJlXZwtjtG7aS6r98ShimtDBXo
8EbT3Z6HWfg6t9PGVlllfNjKRKMovtuMexkVZL0uvHjooBE7U929siMHmoxEMwiENuoiZZi1mQnB
oOle+A9sNwQqvvhy7/0AIXktqPt7QdMY+iPzZTQMzqX/fYNYl6Gus2qOJOyNsVsaA3CvhkFLT1Bu
fIySexGdeVjv5FJd84756Ur4e0Yz6JdfKEc6DsY4TFWkyOHaIc/HpGD9juVNNLFrZoi/DhNebe8P
yKI2+Dm7HfB2QnU90sYxf2PkP6/P/keXAU09s62bEsmvt2Q/wY56bivDdbN6Rij5W8CpoqE2htVE
R8CnRAVHG3r7O6lr5jFh0+wmmAnmWLLxc9D3hnxaTNwsLfJbkZHE2sN4jCLqqoOxBBIC+1xQo6M4
UTQBTaluJrvduojAIJKOvH6GOAVNIrQkXl5GkStUvgqlF8G6Pr7TCvB7Z80+94gO8us1JExi/jpV
WGg/E6o1bPQXwWfqSnas1PnXWbnFR0Tl2vIjzCBQ7VHVYEgE13BMk5jZ7HqBS6c+wCLBxlmLiS04
O3kt4C40EQ5zQ7LDuowt9xBaC0c7LRlh+BlK4Z1ExjsBWQj5CuslxJsR/35RUCdNiSo5dM4oiEfF
KcjR+eKE77I69Dbc4H3AJlyKuS4vSRlPFhyhBJ4ayTvRKw5OX7nksaIyDhpusM2psdtOmtGpcWKE
J2Tu50vmL1QbonYyTvjkLJFinB6oBQJPwThPKJ/cWG4j3jyCQnJkzrGw59X2DCnqPzO2oQrPpkAK
0bBapMrqsWP+bBXAJ0GvXx+Q+P/xxBQgHr3KFB+ISH8G617BaMlXFuGrXaC33mI+8N1HZBftR3MU
2Lwl3aNO/vU2B9Bb7rfiN8iOXXlq1qmcHcqC7jtOkDccfsxDpqnnSe2yJSravMDomIqzeHb1cf4A
5fm1T/zXny0Htg61bOwq/YzMl4VAkb/BWsHPZo8hehWgvH3DmKS4lVZCEGMORs5HEE+KuWmvB2ev
HM8U17tQHGBaZv6z7P0NI9m6kWUmYMepYcvWoT5U7O+tAqbDEtG6k1FQ0EMKurEwfi1BPKm97E9B
kEhPaRD8wQnq5tuks0yt5fhfw2GrQk9im4ZFVcdSLuXbE2KcPEv8/ELmHGXJRQRH3G5UdVa6JPO1
pTKvxSdAkcROk89PfACB0aHWD9/mCu6B0pD4a2zZjOD9zF7Pta2nFwNdGLV/Dr6jeFIHisNQQ/5m
skjxQ8T5Wl5zk27dXnmwwQ8jnYMk+NCoW+yE+CfdI2p80u+1LMt5YZkV7LAs5l8pR/N+nC5IiPzd
eLpmctf73nqH0TAuLJBeyGOKilUDKUNez8StCUNxypuYyJjWrNHqjlyHvxkzWllaUAJqSdi9AQsE
0KMOVyimNwrsktwGrAr7CbO2uTSCZSWZJ1xyWykusxOmEStqzE+mYTdt1Zm0hyrvPmeeT3KZtNkb
wJGaULyivw1bff3ySjC+bOPnNIjXDe83je1jc1VfFdlvsk3IsaxY2h9EdxL4XGPn3DbMnAyEuqyV
WOkoJBjrbTjTmBjAxwxmHLAGpE+FnMD69DnEQfIc8hB14VQfoL6HJZLX8UuEzyhu4Czn5SZhUuMs
RSRRTnB4bQdbdhtTEiuuJEl9VMTTqZxX10fgFPT1TmTAMx+39hUvPJmka8StBIogTseg4EfT7TiT
H1qJGMZGUrzgRGdzsqw4im0UnzjL/8BkLUmvH/9N7K+9Sge+pQC+s5wBqqkPVDrWjSyksy4pgrRO
+e3aWz7D+zzuDZoBtkruRRwSOR6diWUvlFxoWkbyNSD/u0qsmKqxiqf7qi52xd17cnEojARO7hud
kG74TUGc7FHMUkQNy7XD+LbAw1kSprchAYLmrPqTPH0rVYvy/S5NsHxZJ8bARXYLAqIuDbkmaTLj
WwHpC/gOLDby8+GXe6ggH9HJXFIkAytyv67LMt8qM6HGqkDYv6zbb3GecMz4kambm50lxiIK4gCO
MQbQzqAgbQ9d5MVRAPvz3wq2cBZOtO//mT1dlup64ocq4LT4svrKfnp0iu2dsrcE3eGCh7N1Grtw
h0Oo67m0hOIW7spe/g32S1tyMgVftoe3B5C5ns9qa2hDYzJxx38ye9XGZQd2IRQQoCmxI/AzLEC1
KJ1stoJKAmADKMRSUWAEeX0Y+bHLs9HevMc3w3y27nkLktQjBpHQ71K5SrZFZrMu9hE4XR7nO2/F
iIa49b9asiWhVo/RR4fuakO+Kpiy5WSr1Pq/PVbbAjMwvkLQQNiGj210HfzARK8YFR3hLozVj5f2
nEm7GB1TYeWelFBQvp/arWn2oXuc3W2lnHVM3iy8x5F8MvpZJxGj5AlEBcv4VRsQefSsNOtNYfqg
2v1pwLjcEAOhA3VLwClCHc7EmDO8gKvjmca2Psu7qQviCW4FuhhMOWm1O6s/7BIHpKMiDFefWDlu
ss1uh226GCJ2Hu4epb8LZJ0WZnKS9etWybxs4XZYO3bsLiYTyIYzBFd+6z3V5fPv5c1sTlb6Hpgm
ta8p8sWhpfCcPXP148FND+GrCv1zUvqqQLFgIFVW1rIj7SZl9wwLZ8DWHydIRP+ATYLsZChcK86r
EUF/3eeU5bXlGrhfnRJuUu2pHdjGLQ6M8yf0R6gSh64cJlfEluXYLWT7EHkhZM2X7hd3yNF67cF/
cRnNkGLbTxRYsjWZ3nwKf+LOk+y92G5i3p9oqZQDId93vz+ex7JRCcRSVyaaBsfNxPNvNC2xTk7i
twb59ooMkFqO8u7qAWWNuLMTrZW8ld/QySuHEn7o6X8oaAObi+Ni5Z+Nr+UIdt4c8dv05J0uvI0s
krXaId4SpATyurnoZ/TZydgc7Y8t6ytXaQbd/WSVxbJk3NxWcehC0YhyHehYJE5uw21/KxpjJbjJ
HsxBS8+pDjnJ9sQ+dbHR2YlAOaG5E3q3tN1waV4d8W5d7R2jxZZY1gNjYAQE5oj7odGOP/iVPQ0z
eJkVSsQKKndm7p2CKrfZW1Z/s9HJ0sq1X73j3Ls2TYOVB6N97ouCQ3Wiokw+Du8C883WSqGjocgs
WKhjknd7Yz8aBnTemXHZgSXnbO7CpcJnYTWaCH/bw/9JqrMAtICkvpe6L9YLU1crRz0m5cvr/gPp
JUWxh+sN5v9LcCrvayK0j2J1Y3EtnEHXcpWbNrHVJ6k8VUSeAA1iqx75LjCOOYETsDcxZNePfDN8
lWzkswO7zt/rtS6b9PdZw1AcVuj6LsTDuH8kijnSJ9YhVSou4WoWcw8e4ezmnXwmfJ3iOvp/0nTc
FdCQV/se/mrWjgSugPuZa7k1tLZsuxYV/M2MJgs1UQ+Erz5K46ZUTO8oRpL0ycQ4ulnc4VV/lKzn
ZtscVOvAreouSzrF5Ub2uVzVoSxn2seuRj6K9b1lnRJDIDiU6iix4wmC9Eb4aL4Q4F2uAFoJrQlF
n2HyMxP8W+uzemredxEpYvEJ7cYH0gtd3qwFatm6+4VzaeriCObqhHzhioVLuNesVvMqilVwL5vk
sb9FtnK+cXtIITpGSR2e8sf70TfxsdgvMbu3Iu8FkFy1i4R3SI0PBEueAXXS8CPu+VTIAH+evCNv
jXrncpZKuzLHivyBR0FQNjepDUQ+/ik9o6J4SoGLvCCqrh1p8ONqm3EcFpix+Jt81nG4QavLtdrT
Jj6AIsmeyIbr5dDcfq7DhYPLXjeM3o5J5kFJbdeU+haUWf9aJ5ig7OR5GXetK/9kgHRmd89PGIDl
6AWq2ASYF1q+Y5jEWf/I+2Ec0qUNAK5LbPHT0hHcHm9KPthp1zOthxIqaF6j/Ma8I1yOIUctv266
IrwIi1PXWxjkUr11x9CAWmTvXY8U1Wb3wnmEmnUiJ5AIUbRhsqQkED9NwkuQqvzL5R8MRcSp3R1a
lk8zzXvCrhms06I5PiodNbBbc8PTVWuOtwwC4yU3XyCG6LALoCuwskmCNRwdRZfG1Q2wPTTSHBto
nP+gGS5zFk02wCdJCZ+qaurXdytLQ+b/aagOeBawVfEL2fxkbHTdVfBa1qM115reha2UC4fF8Lm5
v6kfxJUlkF0yUTGgiFHv1D2c9GvVM8rXslH8q39d08GTXOO7o+PqGFNvsJFI4c+pEGvM1Y5YwKXu
XHRoGhzyZKWGNWCn6Mg6mS44Yr6oRmfgAIA//5WZQlM117nAMw47SmckBUX0vHQBkPuGMMycFbqy
C9ikINQWNEsiw0sFnx78ikjSVMz9oKDK4PnwrVBfSgIRTYm5FNq9ZoGQwTFtHAX13xaljTMGB0nx
HXA5QmlJXcYeSVDy3qCO9fIrQpPG85Lnc0K/8Z6TLvY6I7DlswHNInElYVkjdzkgM39xpx7d4jPR
VEZGFTnHnLjHisyWQMcUNCvYV/otr/9GdAP/NbbmD7F8a2zNHAT4VOx3FiY1NivrUFgE8b5+ik+Y
0PoYtrkoCOyOPAPQZp5fPdFann3v5O7YjMwB4c63Xb0+tfXEyyJP6Cjh7/ZdJ7AyNRZLMnjUekcI
i2S7di66E/cJ77xqJEK2bBz7GAS8rQ6wmmau/51UH1Gz5CoazuGjv6hWA0kg4eYNqXeoBUVwOR3X
Ra9naC26TKwwV23VTjTg/8mnjPt8BTMq4kS6luKbVsYxGZwF7/PEQRs+QMXbL/6Gd0G/f2NUhqDd
oWt8YKS8BDC76Du94PgXVnggH2pnQ03K0/Nh0behlGfiSoMyuqCtFvBFWbixNA1MFMMZRdMnKggt
M1cHsYm4h94qpFP4ru9hNICcicqoQwkFf9F61vXatw0EYXl2ohvvL2gfbtBck4YUELuC15qK4/id
NySpUFS598IwyEPgT13Y056JJAMbFqBXWvqx5d+RmaNTSBpRb8xgXQcXIcpwwGa7YgE6KKl52g0F
jRPtjqKjeLB6yVhQoqPZ/vaIKFQTseGxDV4nZ4+SakKvQtf5rPyHr/P+oGihUF55pIT/c9mU7hYT
MB86w2hZZIfFLNiv154LokR7g6mHdNMe9393ARwm3OyIHtwEPp9Lq63JJ2kdPt1g9tQUNpQLDiwu
D3dvKusf3AXFgoIn3428iVPRVn9BmegzeVaUSSrk6MuoxOTOw8OPRBOjWgPX8/qOeLT4kXmvl3TA
qcGYrUeoauZ8Ix9j8ob9YvtSVThjFG/dv7m2APksTlEua0tk5kL5cVwkLlK+9q1UJe+ndD2ecWMG
wD4SbXxc6b+lsFnebhqB+tDnIK5gFrQBfB0yHxvwLb3+F094okGaao3bODWHSuNjIjf0TjcvTHuc
vhahDAw8z3/QmbKsbXI+awZbZuE4eBwkkX+KMdqtWSqeaLzz8dCkhzmbcZUUSA6k2+5fApYGI/Fi
+dnbTAfIZxG9x7bvrwHsK5PBuzj2jEpgBxvuJWTqyDoAqMm7fdJeDrJpWeqqyN8sLJNG+H4Xe1tH
MVy7PWk3/1oc860Xl4/sDFaUbbp/1+v5tZTmH57XH8DZHYTWqHs5aQz6Kd3kLuLG9DtKDzlMuVaH
JlLVh1lM7ktpY1U4wAbA4D4ke0qghy3e1c6egN6YHZ9NOOJVKoSL73Ry4DmqN7i9GhF+yRkoHBYa
VrTl0Jd4pcoDQcYUAgROOZ/O/w+Qkk+R6VyFDPRk28NfZZbKhipcLp4Gjbz4lL4Wd/RP28caHEZk
B+sJeWj5F93fas31FWNURoagALMGKLeACsQuuG8UmTMxAzcu8J4k+xpoeJv7diTav49s/BpQBx00
tu/YoKVX1yTFZFWDqm3WrvYiU1tLAv+Src5453hOOoPYpGV2UnOiSarrQsuoQ5Wu6NfbrNlEMe4C
xZoMiby8YcMVSHjs3wObzwjMTAPa5kk8L2Tf/BRmaOYT+vFcm+WiLbPQBmM0GjX2Yx3OMWZhYoyc
doWH9diKQ+RANh7tS58bNzYgHMCDfnbAWibvpye+OjUEY6Bx6+gY1K6tfDlHpe6uPDDahnoRb3GJ
6z8LfHE9LYCq6qWILR4UXAflJ3pbL91kLI77EvLSDH48x1fCKfzF4WF27GvJI00gU4f5csai0Y7a
Tmsny9ZfS+SaVwlJljLbASq69SNRoS+MAkSQFQkMl5By9xplT7O+GEJi2Z2Ge0FKk4T0wYAEu5zi
AZgTGWBEiVSKYOVg+EFfcK2KDNAM8SntuwxJEDsBXnfdOkLkAHQdvsCtzQUkx05X8cMjM+eF20Vf
UWTPgLimMNhu7fHz7MHXcNeM2PCaTr9k6mhoreaIK+Jm4WNyEcrUmff2uogqTur2VYpYtHgJfUMJ
EnGhY5AsOMSb1HVIa4JwPVrQQg2ubufsp7h+m/8TUN9jkIDeVhykUvM+inSJXpAP5A9EW0+Um9Ta
yguF8WldOih9ua8oSGN/79LKfKiP/Us8+NRoi8mr8vHpkh2yUof4FR6tx7NQ+AP8pjQofQA6bfZx
uCuxPGkddWQc1RYYvLMoEJKrHsRc4Q8DADccou5MBc5eIYKGebk2HVcIce1dTD7FBLJkNbi0Z9JK
cgDXIxgucxKwzaZfJN7RXRuBedVlRsc+yH5SP1Lrc3iokedWDTWyTarZ5GDrR4rYJr8Kk9beB28I
BxYaco+8op8WRkJKzrgquOw7NqVsmF34Wv2YzmTacrvttCv43oWCWz5fq/Ffus9wbQ7JhKoKjv+y
+QtefyF+Dy5BGo0Bx+9Z/BdTqKnEptRsc3yFUnSU7t8w2kPrHrOdHelePcy3l2GHw8vcWBetb1Pq
vXwoJxBSZwwegUUPTwRjGGcbJdlxWi9EkHf5uXjHegLvpDuuSdxIk7ehYaMAIs5xnFZf7CD9Ebrz
bRGBaTnDwNyuYDsx32wFqKbPh+Br9lrHTzx9AyhfyLjh43irrIfs1xsd0M87w3jVDv846/YSlhcO
opaYsrHoac1fb8y15ZxCqONF742mo/8y3NKcMJUoEtxKHN9HjXaDc+LuVdijhQiHBuDukkpuf5ge
fyAlORCWv6S58LD7IENoV5yPelnQBjWjDqoH5sC5Cc3wPicsHVsi4DH1fYLyVpcH/naemD2dcG/a
1VY7xgkizo9RNqdRV20HqpvFmRsyT66QLgNnxUTwSSLA91uYp6UifCTfWZLhxcC+oT23qFLzX5kQ
Iw7Zwqj3hBaLOg6XNgTzpT8wXn0ksWcbRxxGQduSnDFASDLN/eFfMUPBpAuTluv1jaBaw/p75lTG
qrscoK+AnkOpxMPPLY0j+ZcHQdGENTdnAAaxQikbQbDTjryjcla57cioGgdMVy+YmtQ9LliHjR/t
sDxcrNK9NS+7hN8KC66tuhpbmi9ErmjrZsaeU6zTI1zH3eM2/UwoLAzK3Qzz26z+yjfGIXCya+yh
FcCzvDcZO3TAs0Sy260ooP9ArUt5l/1KgKVMQCUV/yHihCnzlYpI/AH4Cc3uoEL9NT0QdoTETjGM
n4cWFkO8GE95VYW6ybW2jsH0sBxYiTDJM3EDkP3KCdcW4Dtw7SjANjzTM0zt89+JSx2ULlScq3dD
Vki7mTXJQ4zKMjbHN23ZiUcUCsSuLLkN+MN8O/1p08/W36uR3suGlgUIUYBsie1siHcczvUQZr5C
Q2G0qvxR+qv/59uglFwr5qQhQMiH5euOJiww3Rf5knDue/HxPAJx2gjCL6rseubBHkC9abjwdlKp
4WEaV0Xsdf0qWTiB/XDBKrDqq9lGK4hFf9Nt24Ucju8qxeU9s6qhsem8jP2szLcONt5nNVs/VNY6
gXmCgfY3XEWZWIoZ7HX3mtfrQsHjFQDksewSzs2lhpnHyAxYSRpx1+V23tqgUBJxv7XAc04zCfhg
yZp3hfo+Ynz7GJpddOBLA+/7mFHrn2u8CutY7CvsPnLQ/CvHVqfgxPsJ3wT6kA2BEfoF9kkSNP+s
rEgiecXBHKk5ukvFyqPRLG7RQSEJpsgHvPkKakHm+6VZjV6wz+3g542nue696uEfzejovshalZFA
fNyZkmaAj89+cLWkH2k5+un+dfWyDjs8OPnT0XcuYzYEn7a0TegHsUnwgQ//83m5maiHujsXjb0p
k2edc7Fvlrj4WahfDB4NtHP4brgEqSJASQ4GTH7vUSvfzQP0qJfTE0u4OOu2fbAdVlxhbbMHhy+v
EE45+t69DkYLB/eR6Ti1JS7LlZyNhFc23bdhzIE4Hspa+y/owwwng3+bTGGlWiZUYSFJeE7q7I9K
p4rdBoBounUFRNZZ5irESdcdymD4Oe1hdZXvuOnaxYfSB53sA9RzGNTvayz/6SiJtXXTy+6kf2n3
oNIjHc3XE74QceOaRwIaRcKj5I6s3Rrdu+Qhs9o+41AXILdMlOcuNzFywCjSevrTPQ/CFZirgv/H
DPmnb9GOEamLCSCBeo+RCVC79jWJftYOb4tkStDoAhnTYytZ1mUYTdOwPlQesUfc6HXuV1fCJZzw
WZkMtRwniuAXAd1dFmLpKtXB+PeI0ixAfDEDk43N4YcBFdPU35HqMQvTUqa4qaszBumpscm0Rsjm
65gccykAz2BuNuBDKTxx2wfV93ALzmx1VLqE6yGYh8DkBngOJ9iiZZhMmtBu0OWKbQ8a04KCo2tY
jPgrR9KI3dUqWcEB6la4ofM2UWZLRQFSUE7eZACs2R0Mcb8zMs+UGmmloGZ58Q5sgzCLeOc7Nt86
yi2KLTa51cx5iCxwTviSxSt9RE9EDcmCt0arQsLnl8F7aX6ol4I2s/HfH225jkn8NCEDw2XCZvcm
JiOJ5tkDSjkzKzIQcxjwt3tZ0cpgJMjvPwIalPobHLNLy/rlcL5RckNAS5wVy86nr+Pf3bqICywV
yig3yY7HtTEjwXfQFqC5I1vMO4KOaNhNJL6je8P+BY+v3CL83n2yI/MOa9BV5GBxFClXGKoVv/nT
nAs46tRlTtOH3YIvwd42cgXnKh6YGAH0tDyKy5sJaeY3XhZolApybJq3112TfhfCu6+upYBcWvbK
WA7YrBB5IQgleTT6TNcRrxgaOKRQyaGkVzoS94c0r3yMo39FO4sQc6J2EpKKWmwBJ44DFkCXek9n
Y8d5QDBBECTMFhqie0PUHRh+wYwpFVrrxwbOuN0YD27K3zWHd/QG6Ghcqf/UtqgjUsvflIXtdasY
YERrFFFzFbkXGOGy6C3cD+o8v4+Gr+W/iJZ6Zl+gbc5Dwl9wCBKyxRL6kgekkBj87sYbwFyU6cOp
1/ckg2KcefIMhlZCg3AdCjxeJ/CLwKJ92r6lkaEKMFi36UnfVq1G/xvrS19rH8eevvT/VUp0JPdY
33npKuVNWruw5CSll4I5PpY24HQhHldlUuMkD7h6gg+RFg3PjHZpwBI2Kp17ULaD943VCssZhzuL
9n7hZfMO/GXFfqYm7zEG45s6C2tPFF1ZrYY+4ySYv8z+9n+JGY8s9Pdmumu2svKmFtl5p03lkAfq
wyoZt1f117PAqiKDEH+/1FmoXKNV9Yo6usxpt0IMSMOtbIQHVJtO5XMuakBP6XYFg5ccA5jd39Vt
aup17gzvPuRBQrxYtzhAyaLCcVS+EDS3N5OxWSrponrMkqYJhLFn5WFgHOA/MRYrNwwppPicxUzu
/0FIqbFpfXN6/jB5x5HP4/HkSFJBeTx4d4HterneHLQmygyV2sfHZP9OB9bT1AY1ofeuD5S7oUdk
B7LyJaSfb34MEJXD5eMT6Z90U2J/w9kGs8zC4qrEHpLR+qlza0mk0VltdoS9CK6FKss4XKGb+g/s
bJFvIKPPyGO+z9soWBJbrjKbY+IF2Ptj1PRt6VCVGWBVZKZkcnZd5uRpXhHyDxYvYf6S9e/O+BQJ
MB1bEh59+OZoKwHuy1UKzYT1PFzxxPUS+5jt4jdQC8C/W62aNp8fs729Rh9Bo9WaEM6mdWHNNkwz
bm2mQChnzdHiGvEfHB9ITIkqfveUE0M7r5LuvJBD3mhKC16MCZrqTreXF4tU+CSHy/CneufS4+5I
eDVUGZh6J3Fx9iNkNRhZbQ+dxRe+ye3tQBAxdyGzuWgPR7OJRHTbMY6KEzuD4A845SBVChJTpGPd
fPwJ6afLY56CYIwRNJPaCc7Iw3wHRnEGTsbuKfFdc7hZbvWD3iVtb5/dOrwa8UL7aas81mZdRlps
5RdMeOhb43RFhczReswfh/+TvZTfrg+FrHWcLYtHI0HDJMj9FQxnx6/ECO4UezdvnjK/kza+IhJ6
Mw5IAzq//+9oph9G0YllBm0pli06DBi5hcouiRbZeC3bhrAw16zFYPUkvv1araS1YMY66Mz5VzrE
D8a15P7sixz4wUpELpCXBd9iVAd5JnOGxPrCk2WYOaZc3GiiXq+PZwOvVNUqS7h/1H//XYKT6BBl
KxNlKAS9zkNDL8UrsHLJM1iSQnDHF+QohfJLNCJlp7bzhi5RZ6Gu55+2khiYil9rP7PtUit/E61E
vX/+svdZNM8jTP/bJ7IPuuMSsyWvYVMawI+fZ97tR2wqYhzo0fyrcNQC60WtXX72nd/3jmtSH2Ku
/L49+Y0/YAXfMDbIxcFHy4eKxn7MukXZz/CneeBOsfHZamADxB+XyT2rho6EU2AtYq6rkldweOEF
fyWs65vSmOGfw+t59LIpOhq8ez86nGmOvmyhHYsbKpXkINfhli0d6SaX8VLD4rUf/J8gVzsT9gyx
8WhSCkNu66o9QMrVqua4OyrqtaKhfUxXlRwawHzT730NT+FpXY9S+GWwye0LDeKMvFL4oS78IGRU
+wohIFMjOKbrhoaCCS32oVV/70/VKaR2L8u1xn70mmZOx0XRVpUJfCsv9jEozXTYwlmknwSispHI
xfVO6o2bTAf6FCbdunLtT5KzC4n976wTae/k0RWP4RJXa0yNe421jHhBdaMme6AjStoqAGUKe8Jj
NT0VZfKkw7VRqMarM9IZngbbxeeCcnnVvrZzwbHhFusu61gs1QKOQtros+g3nUXNpI7LDjz1KG3h
72GBD9evUegOAVoWQg/ViNyHFb6TgOixtZ3EIa11injNUX0dnw+AJDWrLz1jgG8L/6ozwMpXXLy7
G1lFU+xJt4SD5a1BWTdaDhE3hNlaKRP+xpu3M20UU4LAdp6OJ932mUy/KplhKLTy7FgZFTnaIpYa
t0UWxbWCUWn3Nj2u7Fu1JxksKja11AXKATneXJUm8yiwd3S9a9Hal/t8FmNqG2VjZqkDgK4LgVBK
Aj+9W1wr/xDTQn2cK7nhZh/kApAzGHvA7AJEugufcirMDOEpgyleiaZ1haw9+RGIGiUleksON2Vr
BbnPeD6kSI7rV6HMQAM/p08o5vE0+W5EhLWFn1JWDZIvYhnmDOMKXlgSF2Xj8fOK2oNYqOol8tpK
3gPy9p4MQKKHtBXT0VTHDsT/pwYuleUgLg+gbG/VFG75rXVydzCMEsfndI/pvpY0JstI8zGp9pmt
hm3pTU31i+IekTFiUq8+hkmf7+0E4HiOdwk3zO7jqpOhrq8twgHkDuUZkVARbKhSEJzyTp9EKxqz
uOUuWPvWHWctTfXR1Jqu29DLN6QgIvl4vcbRRwMzSGQtuEt8ccaz/NCLLOzfQWgrKsu9dGialyBS
IkNm/UN+jYMhIY3WALmyzAdaWUxJhIbpCBSE70Cs3I/rSaG7kRF4xbBNmqDkpq9iNBdc+5AE5reQ
kXZ7qTvO0t+yMPVvi6L0aNr+OmESXtNNdGw8tlzMdPOijTc9m6tE8IbA38GrLPjz8hRkgIy+0nUw
lnmzS8YIBe2HJRzri8CZzMUFcqW0hyflJUNd5QMlDln+1lNK05HEzaXmt0i7Q7U948lsYm6TzmGA
bhqXNwLIwvLJfB/9nOZRGiiMM9fYXKDs67YPYN4+36ZfLoIXEmJl0fO3lBqrkFgAnzvOCx12lDaB
EGEyh1FK8AydbrWBwmznsKme7HBKRKwZOiF7VMTJeEvb1AVYUJ0qPSt+skrbqEhh2VrBu/mxWHRL
5J0J4Qcnsr09VN/7FKTmE+IOP2WIXpRSwpU6Gk5v6ZOpjcP5kHk3N9pFUqzwhfJ1ckIre79PgmoB
gfDPr23+7jEswR6dKwP+dZDWVUd2WviOmr8vUx5FxFUMYqYBow9WcqvtPnQzcC1kROnWzfl3Z/bk
MV8UrHbI+OL7wtf7tBc6eB8S1JMeAsNEkKgKk+VsenuAQ2Xrms2jW/sJsU0T4hFi5eO9D+ZwXmEr
k0S+gDFSvfW8Rb0XjWXEg22ssetaj7nEK81Ct9Vr/ferNyHrma5dsjPnd+Iy55lPFrgQVgjLgPcg
BhB+xUgIXU/jXshbN3Q7KAR/fhS7s0XP4IJyGMYfCmKS63HLGL+Iy1zgpsCrvMd+SkzPVg0naDx6
hF5gknfjrh+hqv2nIm+RCNtC5YLukCdjMVXHFhzmcbs/75yf3rT3bA4i2qo8ViHJjdaoyDsK+uWF
P/UOO4tT4+ZB8knC79TLe6gOj28EE6YauBWlMc8HKDM5n6Ae9kymcuzH2Wf0nBncXtM2Ws5k4McI
yBpZah87zSRVIuAebz3VtZHLaCuN63jZuTed63y6cwG0EmV/dG28HYz9bz/M0JBkq9B/M5CDi6b4
rHvlKwWmQjlQ23v+7csF7BnWZZpHmyUOEoNDXi3n5iJcir9KAefnIwSNLkvwZa0hQqZyI3xz+MTw
qCYmkeHjb1xQjo7pSAsTJhAhoR7rEyKwhUDPm8rlNs9G1fxJjA0k3Al16mTQQY7/vblIdKRHboqC
xtxNG7qO6OKlnIYeFkT6U5j95SsLbLrXrwVuq39FvJ/bOMcYf0HRvUEnMbTY4rEQLCRmTt90inoV
iy91lx8kkVR+pN8j9e7oDBfoA1md6afGG5j9w0vr6L6eS9uHvQaHbrQ7XOu1XqKPHChv3Fjbqo/k
kzwwZH9ASOcOEdLR/CpfI7aORxQwpZO1JXb0cFAsncaYbF7IXgo4e9IR3E+CS98PG+dz/ep2jP8S
AcXDPj1DvNrTUZlOBu2bwBr1ltaUxIvCjPO+wzAD9k1RPemGULAgeHuQsgRSSHMAjJMDHIm/nz45
hIEwbB4a0Z6JjoXvv/zHg180Xi/ZQ/MY4vG1fOC/JcMi8lxrETZ+w3INKShjS/0B0EwKkls+oNCK
RW15TBtfuY0+xjb6yP1dqgCFoQ61wYNtj20KCTWPW6mJ96VIQHsTVEps09HiHU0RzMELAN7pCpb0
EsT7JBTZVWGt+3vyPVzci+yzvVci/mGBk+IHtt3HXMs0/w0ypB49Bh11CQUgcdz4yPk+OfY8P1Sh
sOWryvIP4ZZPHkTR7K3bn2YzCef/8dQkGkN9EtpiCPfV6ZXtnvQAHQgwK8V9eS9L1Fidwr26H3nX
6+Z6zSU0hl08uQz7jpxoWdq4fy2EJQknqXpit74WQnNmh+yptn7Moq/g2y0mF4J+yfj6R0aeoZZW
oVig86wcOotdGKEDsPWYXEueIvP4eIckKb6/JSQrpcZ7fiYimX9QMO/6v7huNgCEt/17wnwvnEMy
G26gD8iWff+2CXUIwCCeiflIUQDNy6d/1vzLcZBYFM00RmSj6MGxMwyFa2ulPm5gNWWHiQojzzC+
U9DXJe8mDNSGJQNXH3KSTm718ZLcVUbZL9Wpq3YhXxjdgmqvqxwlTEVcfxzDAb2/YhPGxKVxvtNP
ctusB5uq+k2C5GlziolY8fVdFLqfgD77JmFObm5J12/X4AxfZYT5Cj2qwzyGzJcsmK/dLXGgpOcR
oFalF3a6IfkMmqhb96+CpmrHkWG4LnZWcZMrKfudstre/Ds3KS695zb6AYTraXtplhlz8/me6+MC
grRYpnW994IcrIAiQL+SueIMTIakjsEwOW2Wu+S//1sV5kfWCVToIyAQ6bPH62Te5kXEPDBmhhgb
0UNFA/GLHXfgRyjGx1Ttb28Q8TUiHA2Fll/1FDLZQKC+lVC/PzJujsqdaGySoucjbH4ra8nyr6kn
F3cQZbIB1+TAGP3jmHaVCVxUis82zDmmTc7CK+Odk5axQtrOE4KWxctrc8PgSJBMlZOIj+5fY9pi
aYgrTTWE3oCPnZGksrQF63Ik91xD7Y47ojFp9DMjMwNow5LueKisF12Bw5oS5c1i03Rc5p+AZVIk
lm4zMeklcIQOuSRueiWgpIoHoMVdnCDWLSV27vZ8DWkr+c8L9StvXq702SEonzmAgYgIIop+22NO
lhkYlq2qxXd3mBk09n4hfI8DpiEC1yHeTbhk0H6/AVVIREcR11PVgixNRAgOzLaImVyJoWbM1PDK
tQ17AOmMEAv/DVh6Uo9dSQoIrFrRc64/XZRXI79H24XpEHWUocQUm7dHGRcOkxyniweyV0t1fCML
cH147J/Dnv9qpFfS+56nAIYluHM7+lJJyE7FDAOfUo4P48Vhpd8nMqCldqfmDI/dDo5De6H7mxYm
YoW11UoIAPKvkj01ExwVzso3uzFOn5xJPy6+6DaBhj87y2v27QpflJqkV+9+nUSaWLDJvVJqfhZG
yigmepGNlNFsaKXdhCHUJfJ6Yrd0xTCJQXQJA3W35kzjgZXE1wLAH+TG3+ppLqxlHKqHcSZUUjo8
bfUjE4aAFGfT8DcmR9eIgRpzwTdjzH7rIJGusRAhYRecvvb4qI7cqoTCRREe/1NbJwou2B2DOIJq
gmPeVuwKzsqOzm4/83Y+WY6WDqRLQZxJ7IyDZFqGbN5M/G/HTnzMuime4WAgIUi9GMvkUGkLpMpD
C58yVyh7fpJg1QWuGRsrE592sf1+I4zzGN2id3VPjv8yrVruW8cmqTfIy76VDheQ3xaaavT3Lw3/
uCCejUJQr6VAjxYZMXVOm9MihYKWyPl9azzB7B0Xn3WzZ/2GKuJJYTVuMOpNBWLwC6RPgPUXNayt
hOcp2mTZDgyYDqkEBuFVrm/sRdyFSyKFBBk9wDOSrJ9rwDz5PTo70YK4R8F+cFpXAkOiQl2gkkZo
jzJhw6Gzp/i9UVkHt/CjyUseKNkNZyFkyO3U4zRU5iFkIUL/lT5kAOJrYcdpzZoa7Aw+92hFx0ti
QwyiD8CU7ZYIJF6ao+Z6oGBcI/3Ku67G4uqpJCxxtuUJKiHBsRutqVVlniUpX9B8e59/xTLsvIg1
bN6TqXVHIWpx0NwSAYJA1EM9Z4OyYDb80YmYhP4HrGipzadfveJCd65NFNfRs9ije+yEWFJsK9gH
iSQCWIjdzXpwLMT1F7SyROP8CKIa293vw0pv4JZy0vZgsFcDp//aX060teeShc20UiByNtDKaD5J
b9aseRNLVCpPZiqeq+dUaBDmL0+f2bregZ1M63/GjwUFlJFtiPq0bGCTDdYnuHtxveIEPO9twjDs
B8AVP0hkzFMODCE+bP9vq5tiLA7DettyoRndJevBmiJni7+rz5GLx4dVAZDkH4Ij6wdj/iP5EM6N
EjsTjuSc7Fv+3bTSU7K9T4MJEZjy15Ym1ilsnkEIF6GHhR5cbB9G4zEeRxLR5DxejhItZ443mCrM
JFdiWWb31UB4s2iO1oC59kvXwe2vWI74onzgD2GT1/kWs3kO9eMeiwrUkzcLyGH+8p/TQrQ4saFs
eMa+MZkRkpjDMqakpjlHObuxq6PqPRUVWuIGKA8LHfV4MMs76ZnzsKTdtlTgy/n1FJAahLwRN/E2
OagLw8Yb1y/jRMwckHQ2l0NMGfMExO+THell2F6HJoNWGVtQYNYTmxpAgXuphOkHozJEhbRmOn06
XGqO0WuKpyqFLmKRqxSOeTSRX7dsBxjx1Co/fTxXhwz1hZpBIfM3kKFLmwuW0HXzWbMSXlxhRKLy
KaUR0JAjUZiL/oQxi+P2+t7XNi4MSHMSgQUTIhhBJ5tnmsyKix6Rjzk+1OaJbNbFW/1P5vlp86MV
dpyVKOXGOmoEsnznP+sVTuIJ+YIyNMd6XkBPZf+7sjtXtfIGQQPg9U7fIDpm5qTHHI47rJupr0KQ
p80osPRRcNWB7DIGdWge3bX4c0lVKA+3vvSeCmQQXgSwzJ53EQf9om9I6Kr8JMn5/cRHJyzLt4Fb
/w5V4zDpVSh8xi9kAzkRMNaLMlNqj34yNN+mlRsFMSSApCFp3ZD1YqT54FUnfjgYgK+QB4YoPiez
ni9HassYTgBdrOY6J1bKxkjLgAdGPgtDcX4Q5wVXQTuxJsT+rPhjd9WWhYxBJVZ1tAJCWyxtoSO1
TN35L3M0JLdpa8ylyYXC9PjvVmw7lmRH/5Cb67q9HLlB1x0pNFhfkP6ggUV4G8SdFl8hLTa0eSfF
CA7oTKA6/fLbSDF6gouTOa8SKCV1Bt1049IaslVLsWHolDZ4aXMpWnK7Wink3rOPTMOfzsysohxI
jkkG9h1u80TrmlALrVjrl+JA12Tm4yuBRqTNtj0n0SAKoW4FvwOTHvFhwo5lUnas85o4jdgVePBR
DLOyBuIJQgBc5XoCo/zewM2oVxjLHrGhqQ9YEdyLE7Petq04B4hiKueHrAJiex7H/51caha6YR4q
cniIumLDigfNhU9heiWeMR2hT7TYEXglXkLrBsKZe3gLA3chMoKo7RwrFiCvx7Ds12GnKWjhJmea
jR50cYd+9e1WzRR89nWjWrb8ZR7oqpNidV8HGWOILRfcEnz3fYcTY/x/tcNA6uMJEMVc5wtiLFwC
wFFxVr7q4GGXDPHYU0JurMEWtNU5FnNoMU9sXgijpEKnZ4dhKk6G9uzgGksLI8DWThJRalwvuZKp
ebZbPM2zlDfHa9XFCkjEJBQiEQDx3DE3/GXkDEkRRndTjhHtBogxTYGjOu37D5Ke7Mz0hyS/J2q7
WfaKPPcUE6ksOaCNFz8mlo3eqJAe8/xbQn3M8XyIZcZbAUmFjb/qz6FQb/bXje5xod6YsOI4B8sk
maHyX+QSuXz1gUxbc2nbKbKclr/0Su+egS6LcGL7X1IFr3I3fr+pgqPb9x5Zyr7bBtf+G0Zls0hD
tT3n3iDDFMJueNocZNMN/RD9xHSdtAhzdHYcAfFOTZd+pwPjPeox05EurGHSYbra5Yry6T6QYytt
n2nXg10Blj/Tf6lkCsZoRukWPiLSCCzCqglOBeh1os73pSL5FrTUu0Hbp0L0Ng4S8/OcpRF/jVMo
iWwGosfCeO5dxntJF1Liow/LzfpLwAptpssPlA8LgwsLIXkJalbw1UGXN2s9R80EBZx74igqii9t
wDHPttSp1P/ETRoQYJ0AwosTyNhk8ODwlcLxBo5805T/iFKy/354M5Xbjb/uBtr3/L7joiP+U2IW
Vh4D68H+WrjxjbgLh/KWSW2w9l/8i1dXjHXSFPxS1lco+FmoDeLTZuX7+4jTOPQfJt2y7GSmL8np
ItEX5xHr8QETuXx6T/fboY9oZ9ZALyn9TxV/pXIkyP/XJjNZvDwAxEP+YxpCifZDTzXTzGWNYACm
4A+PhzL5EGBEfjsDFwhcZBq0kyZZTnPfOXObCfjS4sGDlC20FlNvAEqMTdSkQfCbypbXJNyNkhcd
KmhtpWIIKp1Qiz8le3zh1dPdZZREd2AyRT139Sbv695drQ7agmjFkDOApq8xCbKZSZKSssjUZ0ly
aqci7wYTyDWd370lwAkGf+Bo8oXO6ytWmCzbPFTzUBM0MRmMPtaD1Xe/iGX0eNAl3c+5+I+TLTOr
Oy0wHdEOy7WPpe8Bq9hFnKFZbQywq/MxCvPbuOqjYlzl2kGCJj9N0oE5AcasXGEFIpZ7OvN5Jepa
wkJbfQn/oG8Lds6Rwf1ihg+0hmBgByEz7fp4UkPwbHvqSWl2Bbsset6IkwmtUVa3FDdDyAIV8L97
DLT3Y4iJQGLRxFhPZ2FhcPdmckFUHM3nMNhRrgaE0IEMH5znv2sdQnRNKwVXsokloyUiaNeOlzzH
CdfVLmAlKNlVKxALTaaWUpDipP7JMgUPaycrfZsrVSLFMrlt1aLGvG0mJP18BDasG5E5uiHtJkvr
j1jsXBTekqSeHoG/YBHlqG3lXAMDj8uzm0pf5Ko8D2zmt3bH+81RJpU9ACTKtzaGQWEboh5MtoMN
RaaCSeCSda/hvuXttgWoh1vIwbBTHxV8qyzrJM9gqF5RBDbImgB81P9NbgUE+lLm86fAjxfJd561
YtWujRCVpJ7THpaxbtraPKc59KnUuF54dx6GOuPvgPBRa9iNykkOaK2vTyAe8ioxx4qVKPrjX2OL
TI2WvqCdDaXUwSKWODMZ5fRdFbQdGby7vEuq9xvkF9VMAQSU9zIeo3y6s6nJPPiqIJkGckAQuhQk
QUC7DYS9178N+P7dPCvJqyAY0s/HnGmAQjqBdLSsgbNzoKgEsy5RwcMcRmnFruHVxmmuLXMm1I7H
QR2KBnbCQ5ZeUXG7NBDDe1cICUdjRGEOi4Q4LIyzetF4LmKQ+hj1pnRDS/Ip9bLBVi6YG1MltJ2m
H/YMhUsKRh6XOgvok6R3cV455Ai3Ou9780APfCNvfki3hEUN0O2PEApU6iN6OaqO9HKPfJCf+olv
waAFJtAhJ0CDlcksK88lpDNFYXYFRUmPQ4sy1HN+Wk/4xmrYA5F8XUXtSkpndS2s1ACp6haHGiSQ
e5hAJbPITmHxQSF2bj3HKGsLx1GldsgxkJ7/QB+Nnt44J8N18DxZnytc0PXqlfJyyNiXsWOLUoyM
3PECaePQoVBpltLMi1czSnLCG3r/WnVwPASLbWwIKloIk3BFAb9kjO10uTI4rtVaozWojYtbEEFW
ZnIqtH1uQax4HuIQ1h8oRBj6PlZEBLbXVQSNNISiHjfep63+3i0Esmgi7b0gmEXYsOzQen+mT+Sl
Rxbmq8+lp8aNvFkO/TuAJGFVRdm0Ybr542J64pc982LkupNPP86/PWKIxPcA8kIgvMqnHO55JAdB
HuywNB+xUvLEa4MATRxVDiXoilCsp0+UInwV2iBQBv7dJgWyz8AmBcXkF1E+VVr1fi87Uq0bfJMM
HR2GsqTa9LifkgEZ4P92eGZ/N3nNN42isirStp3XSfcV/bvGTAfr+QNh/7EesTHMC+0MJZVCSl2e
Gz55BPP+l1tCOYf3/HzY4C0iPPNtC0hdHkvv/7Mu7VJN4Awgp3duasaNopE+SoG7XdKTUzoPSNan
PHGB8LxKd8l2Al4XFa8Rg9bk/V8nMfZEJyJWrA9cKzTWO7r+gZP2mWVRaEMIb9rj6XjE/veGIS/k
jhIpL40nw7TVC4C/mjmYav7OFOgN2zs54A0+pwsTGywrZB1fjxyupDmnKtWIDqDvSEIG4kHk29JD
MxyInULKsVWch1VksEsY98hnQ/9ONFbyx3mZfIUMYGR9nLN1FSXYfX2G6GCgz7aSaZXSfEtGH0mr
Ab5hPs/qbX7HXw/Qwc/1csYv8+fHPbrV2uzIxgfCXZ96kNgoOVn32wYXCzaw31eJ4NRH9s/oDN92
3lu+JRxeunjX0rOT9WKa0rtvt+r4UVlHqWHZPP2Ro0vXgIPm5tHAZkk3hRcuIBFdkoexLJ6ClIym
mxoZNj7ElD26mR0qbt/zGrU+aZ7iW3KaQeo1wta1P5morwofC+QIARik9RfNTrGTiJr93/bu4KDa
mpWvycq96j3a20XhVzjztA3LaUtroNQ4zqf6RSyTvqQ1R7uW5ule3R/L0Oz0V1eVktAFxAgmztVA
QQMx0ssatwIjT4ycLC5WJ3vXqZ08kQ/c2ayq2GuYFQp9yGv1c/pt36vHL81v18oHC1eQjXxR8JIi
AkW0WQI++c9bQa+oMolISkiaPRUXzEQ054Xk/+G+Zw8C5ICMdjAVqc0hBdUiQB1NG9uMd3iYu9ze
D1qlorQUWNMVifG6ayfhVKh2IrTCoy99fcmhbM2RujOYdnrJSJEfc9GAVHrkRgxQ3hRKLivGU9RX
VPoYqnzUUQS5W28dcvkQ/RF0+UGTeINTcNunWLmME04Lr3tz9Xs3/obEqRMyb++vm4yn7M47Rv+7
S/q3LXhv1sDeLq1itxIu/GCdEsJu2vX0RhowrcJIaQJfGmK7LOcLs/YzBoXVTo+EoroCkjBq4eWu
pi8pSVwcqW2cGpPxOrG116Sq3JhejlAPbpEywWdW89VDUkCDRYP+gndKBfDG6WkMdTLBgd0u558Y
XZg2p82SDevnflBrTVmbHaBb57a7PGZQl+uvbgsB55coy8a9ogYgk0jRVsthHDuopOppmePdHtUQ
BZ3MekUpR1yMVq4qwJOnSEtHqCLOttPaq6KhRsAmM0817IOPrikTs775CxS1KfYPt1rSeiV02FYj
QyfNeVcIOCpZIeOgpAYAeXyfTyZV8HCGEDw/lJWlm7J0GveuPizwv2LYJ2aSAbzzQErOwz8rrZgQ
InmS1Kfbx+qrnqH0SYE6y/4njjd7s09Gqfk7cgGSaz04ujWhP3BxwLZotgqL9QSWflyHjL/YNn6L
Dv85Lbz1oP7ITYqXRAmNXh6gOR+8LWoSOBpZPEtj+2JvgzR9HjDgKHs6N8/QRsfQ5R4JJkBSTxt1
XLJEMTF05BTdZQlWZOiXaBPxnTST4lGO1uSv4ePVHpopbhNdUkpnLvq6+9/iWKQUuxtsp4IlGqGV
di7ZtMQBMB8FLhKE4PQFjjlwQkGHF+oGF6iA4NupUmcwTl5MEGpyGIMQOChPj1C4lpdF5bPq65Eo
eJjb5t6CwR7MjF/34lMiKii9JtXzLH9a9YZa1b5g6UJlbUVw0lvz9GXcSJ57HBS2iZTi8bcWoCIK
uxuQjf1rqQNKQQjRDqAIdE44xK1/kyEIGcVXkgwrR3Qs+Fs6JPYfEgSb2Tf4mvaHsZLw6gzaiNUt
FrjvXeFGCTRKxwELiPvlZ/QKXEwX9EAnLAWgncyqdc3vi3PiISwGrZWxWh2Wz9dbCywAccHF1NMo
i/n4FujCPPH9xJKBvmOZ/FKWIvaCAdt559BWyF4P4ht7RCGj0Z9NGhN38l5tp4hNGShG58E8t7pa
effQ5u4Zk99oKWa5LvWkXF1hwVtnO0j5LV1LHtVCCXJQoJqO+Za5pCQOjuIUe6Q3PxRFxNxdOLjn
gvmx6mPjB36Zdn7F+E467wwfluX1vrVax9iW3z+V23E30UwId6+uYjRcx7+PDDMuH2/AuPBpHN1e
NspCus4EtAbtbq+VV+8jGZSYTlS7sRm9Z7iTourFfYofuwt8XEo55WCNuFOotFtGYjmyqMEY4/qZ
Fv+99IHqDGXeayYpHeVcjdIeE2k7/nzj8xI1QXMv0YXSgXd/h8iBrAPuLmmxUfKheR3XuYdRANr5
Ke/YlXGb9rB6U0yxiupSfD9yNMC3qys5b6IFMCG549lenX5GQ50Ck8rBwFIMt58XLWesow99TmV+
n75SafNTmy+/h2CIecUwxbiRCJr+TxrfbDfUwOgg+E4im/0GRhLK05rpJNqJ/pjZ2M4Sr0syrsao
Dlr40nWO60LNgbYsf0fMQkfzgtSsI/qCw1YErlQtF9Pnec2HYumyw2vVN7TPqbP/g61hMseno5UN
jIW8WU296L3Ac3qQ5XR4K/MUSzpeU2TOCpFewPJinufDZifxjvVgJrjpk0vS9g9/Bew/BkuF7pj6
Le+iseQ8vD8E06cYZN5JBfZIT9gQ+1PzxOzYs9kuHGeljaS9P0muMKNjqDRk0+sfvJx8+1js6lHR
9As1suI+k0tU0606DJS2UN5Z1Dbaxb/C30o3I/lRQNmVSdSJAEKF+nTFeC0PhF0TguVYCPDYz3+/
hnghlTq+eFIWfDhndsMNl0Cs9d4Z9tInlYGGVqNj8U/ETUd6DE5mTvYOVTmDi2woylxyQIHu/0EP
g7hEkkE56L8/W9NA4/oVLUcmHLHqIKHU4PtK7FKXjZ//LlLpWdPn8apxD5cztiGdFT2WR8+mZ5+0
KRSGp4pXaIZW7CHFh/gf7y2AHWF+2BjHNrDjuFGrEDAX9661Zqftn5gMNevIjNiVeJ2H6CgVS5iE
SPSTasTHcRh4eLzHL+lCZBgMFGJPF9W5r+5gZQ9Gvs803FVv67r3TSoIYs5VtcB1N+6xdZHJu/Nf
9EpHm7l6H83TQnc9v2Hyv1W8crOcd8U/L/zoywRT4YjnByoby+wzoRW6hRyqYsvwk5kj/9a4zPrS
vGSDcfVvSRUgSXtWJaG+gOLxHSo3mMIRpANuIizPaf6ah+w5wRheIf9AqajPgLxUAiWz8Acvc8Ww
Rmk/6gY5R0Oot5qbd3wFNrNEI5N245zFNz2aYomC8LfHntKBcfU4wgsmQ8qOks8k6p0h4L8VYvvL
gp2/0G/hDLTN1bf+SWaMnxtL2m4raN0iusPNXAradlxtMe2rtfKlsMsycqDfVU3CKG0RojptOKQn
viuVz+v8/x7dSmyKeY3DThVUVSYPoga+OdllBgiksmG1PG80YBDP66+B3NK0z8yFqhV5Y5IJX4h/
L3TZyYKujPRGDBcJqpyJujGD+e3wf0kMuJkgOVzxkUAIPT/4dA3GXIA+W2qyRYQ2vwWf7Q8egoKz
ZpE08lk+pWIV5v/OgC4pKTh+PdEV9JXI3+jwOQ0qk8zxXaCn0m7jO4Uc/3XVvFTC1m15VORHOeIP
Ssn1GOXziJmF3efLt2fAtnaOAOqDlVRbEuIErW0zrO7frVQ3C2iRGSuH07kckq1UFsUXJLSolwP0
W9W6pfurfB93hiHVsWS98MKMQmg1InSmBz8VmvBlzEVReYfKUL5+5Iz/THmarOkmSFl6qhaWRREw
F+ejfmKqD+PyCRkZB8EZrTugBgozHHun07slYbaFA9Id907UzRNbmj50X+PJrQMZXZzo9gMHOUQr
SS0bhJOe0Yx0SPGnO4gY/ezXHFV6OyP/dK8G+N9if6MTKakWEaBDqK3GnbWWGzLxLrfKDT99mRWr
KDsHNOTmgy35yA/xsOQfZumTzg0c8jzCUcw9koFLIS68rkIcc72kToUT6fr0zqzYgbksLJ+ik3FV
uQdjZVS7VkE11PAOg03aFq48+8QS4SiVnRzL/lFRXUtgj6Wnfi7b7T/J652Ve+/bE89mlu2q3Ikh
Q1L/MMnvrEhxWIIBg8IXlTGufx69kBHee0Ngi0cq5UDsFhs74Dhhmnh48H8sQabpfm66BPEg+sL4
n9WOERgLxeqkd7feLbrhZeeRVz+1Ra74TtU5exHVYnnmjuxIViBlxB9kABIQYiJHp/e5v8O2A+9I
CNQZlXnVoOhETdZdS620/pRRBW75P75jLJLWn+eOm/dnvN88nx01je1ybtJQd5i5ysQ+OKwJHv+r
gftiBD9BeQ/XQBcbvieI7/UglgwZd2NyzcaqLfkCrWN5ro7Qrzv+1JMT9Kn7I+F8YMPVWzIooIGG
bvmxfwwbxen0BisULdFRK4f0z4Yd0w5jS6JM8VGFu8MEB75jmboFF1xakutyPLWshVzYo+FHe+Mj
1siCyVlPCJez/VMve4ScI1T26Zj1/NYtR/en9Yrk5Taamo27C8/rb6KDJjSNus7o0pYt37psI192
covmudvRkD1C/L/shIYJaHV9RIjr+Uiqy2dDFXu3kGnpYj0ILbMisSJtwA12rUA7JnbRm1ECPYNW
8YSnsuWcH0JKsQ25QJnRrbViCt7NVJZe80HyjzB0f7lvuiuXzC2d1PJM6K7RxD6CzvoQ1N0WqykS
ZeW0e3qjB2Bryq90nC3wK6PyPqIeV7J6s6NxY+SYeDtw78mtxw+Gr5j3u7Xj9XKYKl9J4Id3+8Zd
wgiks58kos4jtLQPbgIw4Ao/FAgNZkHeWOUeEd2ySzyHvj4/V8PysbKyPFWh39lfazz1J16WBGKE
T4lqq94/GNlqWvY7Pzu1bwQVd7Sd+c4g/J2KZaVDNLyWAKQez97JiKofQSiLc30XpOgwXIcbSaet
6+sPIfhNBVwHNTlXAEqIdw0/p8BgtfeDTvhFFiz3BL6fZhzktMcXlOP7jVpzW9LTvhRnM2lj7/zX
7Fk8xbNSt4Yh1FSR7zLqChZl69TEtJA/kSAjhzvwMI/MQpmsFRP0+uUQ54DELvpFtmFQUDNsnmSc
ZqpzM7yaKvJDKhNrd3GOnrLbNcoyVy71H+E0qhCB3sJdvyw9rRWmM61F316L6m730LF9ehtnPFoO
BYSF/IWCRzxYp5e0Oh+3T+n8yn9a0E2+NJ/JmQlegzAJqvOEAx/5GrZTLlH5AF0pWB9vluDdpLzH
JoL5bGm1OGI5TxCEURjl4yUsmE7wXLNamqbd8KRUuh+LVQ20DiWv3yUQ0RBwqGb7f2cQewITrHK7
/Pb15qBK1oiHyr9hD3ChKhfCQwLuIiQbd12sWfbrP0NLxIL6jo2pJKyWFu5kggIRHM6q9cNML27N
VsJLcfyFS7etoKK+eFRf1jkA6+TZS1362LTfsX58jtrQEUaM/MFh3Zlp2ALrWj0xUfYd29O1FCui
s1IArxiDAATwSLsjp5D2m5RpPzuR5Ptt8nnhD+AUZnbYT8gKE0Qf5WY96QpIbIxNV9RN8Z0DOFE6
6fMPrOFgDe3b+/w0FobtukGlf+hWmnT2tTVTGwAgnE2nxtNTAV75tqZMGU/AEu1sfSBH7YCUvQSQ
yF/u1U969Ut/SMeCJN+7/ZOHPJoHQH1Pnx8tzbEGfsbH9oqRC7YN7ZytEItyGvmRT/vuY6+bM4Up
GbBtiGe8na5V3NKxTbZKDiAzwjPQ4znM8E+mraOQj0oOxNAkrxHto7nSa7TzMP2b/PncusCVg5Fg
b5rsWuLIIkzD5YZ4XZ1n8ARYLEL1NeuJihXewm4/MSOvLh1NXmJRSWc5ItnogQ97jLv3qbws6lxZ
b72kHrquloavd32oWT/fsc8N0ibh8RJZUoKXn8IsczmMtc2P5jTPIbNAIWts1jWseNw8UBXZ6TjO
jfB2xlw6Xl0gCURbc5/xK0LaCENpwvSJQ/UxgX9SOcOxG46k2VrNZoLLL+uv0czzpD+XQ/plKNea
w16udsF7+YKUPLw913J6ryx/3y+qV/Z1aNpE22vmoqatyP6pr+TtaPgj42NohXum3CCvgO46mkZ2
zeCQG806nKitotys3tnvh/LZ7sRbRU8y9M5EQM06rEPLHrm+Lbneh6aUdYusjbwMbZCzfXcsrf23
T2KHywPJ8UGnfihozWEIZymG76ZHpF1K30DA9NwZZYvMuWGfRIf1Zr98ZcpJTrsWjUhRyWbExMpg
ivA4HP22Y/Eek5p+O4xQTIJpdrjhwc63a56C5po2fGCn276Tu9FXKK7Jo5/aySnRvbMgCmX+AlI7
CefgM60ZtdQCuan9ThOawZn2QjrYS/q0nYHSIHmF/8U1LOwa6dImwqCUwYFoOBgXrrFSQr/T5KU4
p+MgjUf95Y9ZLjKKa6+LSHW8nMugih63vNMTqZgmiuGQFX5rVftJubaLtfCMZgqRB14wQcASpUEh
TBOIxPCIO4crGOgCR/RnQpxMfulqRJ+8tjhrPfMN8hid6TaI7mqS1NNJ+1rqA2r152qW1mRZV2bg
ACQRaRVAb71Yv2CJPJxMGEZCBSNxAYRgKZaQqVchLGyZl+ppusW/xKLsDcCQ2mQEJsFjvgFkJaEe
8x3ADz/og/qwxmK9mLbbLl9TVrCM6kGmOofJIfqROrPOgTIbC2VrrxxTlp5u0fvkjuBQ9UURrUPX
0Jll20byHvXUYTDyFT2w88Rd3WQ/lvwVzwADRCVumWGX3CbO/fzTRtYwPWhRosQBHeuqrVAatUVD
/B9Bwih9chXP6OlNP3nawVmzYrvVJDO3OSiDTdPk6tgZefTy8rqURklAUUWtYsW69CEnD1MuxfKz
Tjs/ve5HdmFSRX4q/vB7qh5OxxtxE2NdsTRI+QpwNUWxs5UJauGfNyc4OAZ1GcUx4DhTLPGLmKS9
318MrZnA2jQNVNF5aAOvjpxFfyw9fkEiOsb84RBVCzBR07Hh2yRliFKWu2TTnAM10sBSd4HsMpVz
dOOH9vRBzQbyHZTlaHMozSotrGipPr1BMYMPjFORqpM7KhOiar1ndyByXdUtDHM9m4i2FeloGBpK
KejT++K4LXT1ZxytKvmhaJHUq4RVxKvDnB5ciThbXV60kOl6Z/ubTAcALDtM3gBGy2W7H9aHvypD
2ZqD6FgHfVtSRvE7Wqr8xUjpM7BaYzs/CDtmMYaTQoqKWFCkZljMcqH1pv2Vj7jIZBtuGXwcYUc5
W+ECJ3NJdUV9i21D7wfr7rsX0Swm5g1Ae2gimLvSjGu3QbwHS7HnuzferdhWpqAfcNym7iEv9Qcy
DzYLXsB30YVU9MxZuOdYH/241RQMPefwDMhuNFjPbkZNACOwNIyE7DCOT3wwdO//dGmgxgFQL/0C
qHeKChcvEmt4Un79t+VVn8zuIcrF2C01bqI8SKU4ZEAmJZZcN40/6rRNFDq0GNrXp9hdHEbzZ8ut
JQmrgz6yKy5IIdXzVxkLtNP90Y6NSglE6Mms1B2k/nCN6K+sgfEZH4s9AAHy1+QP9vGr9a08hQBo
TeFH1vOrB1chDQMWAXDoLrv+9dwdi17kibGvQR8Nv9//RRviONtc/OKH6x+7LgSFXpTzd3QYbNVc
+khlQAthkhoHvSU6aptn+GEtudZe0QUMijYKbgXP2TFKSHg/FEQRRK2GsPx5tyC+/aDVFy0ZYjiD
ImilYxkAASvEHHK/zvavO6vfu+Tni4f79j+AyrNhRtzzJscBIJaXKA3wWipbvES1VaxQ6HU8tgvo
M5NeU3LlofaMs5qA1f7aEP1gIFChuTIqJNl6Fgcf9dunzkS7QhuWXdgmyI8yEaP7v//JyrD5gQxI
d7TMR0HBCt/apyGOgFFoad7Klynx1/UAYogpyBaUYGEpGOiZ87mV3Af/hh2B6FAe5WcLBID7wF1z
2P0DI414D1cEfwY4Gp4U1h9GqfBDnLEpM9U+b/1M3rNogX2VGqMdsxxTVHW9MBmkNDKZHmqJAy8b
lx+7kPf9qtd6L3Yq6uueo0NMMdNAVgPNXhqwoVvG3SpJFaBk25v0+8GzntVeBS1TBRxdvuoIbWf7
AIY7+DGM+3BUJYWW+ccCC6p7UICV4vPBpUuaOXY86fDeqFICyL3Q0k/m8DMaVSLtps4Omi7rOqI0
OTZqOPRxpBbnK6BmyoMiGTpqNyj+jsFswI/8TvAvZ/ulNSAHh5Aai49gL0+hsQcopqQsKHmckWOL
SsjWYiLndb4bZzkwp+ywE2uJ1h3Qjj8BdyjsLNIsdG+V26ao9z+5b2wwU0YUOG6tDhjivrJqwMSQ
OzqmCT/kfS5s8K46fgbFKcZ9ypFbFBPqgjkNhSsKXRxYilJzUXcqzjHtZXL03bE8LAafgWqGPerK
7owCJW3sDH6qZX6yrQyLUb4fHH+ch0oA+NU2FpUzoMKCp+iGw5CF4vfsUpd22EN/I8Dc1dWUmM93
F5onCZ9nY5A8GyN7Q40HpjjVJ1ZXsca5BVjq3Zzk0hVq9UC0XilZ7WuYVbEFLyVhcQWSSfVrvHwg
kiegJOknISonlhKfOdz4xxvaiMj1OjxfQzVcCwXGUaTO6AkN5Ew5gYfxNwrO+MvBKKXWAAT09fqX
954BtZtEhNKvuxWfN8ZQsmFliRH49w6tekdwvuN9ptfZLovWhvxou9TTbxIEqG9HAEbCNqWBLNzQ
1TvV0q2AKKRnfD6Cd9chjZBzQ5jiYUClXidWHHtHtg8Oze15714VvNpRWJxsbY7Sf/oSjyBzQCXX
n35lQAlZelwY5xKh+NwyvmgX8PjcjCWc8Vo0k69qaYpoe+Mm4qBWrk/u4ocLVgrBNhaYVDIXoOF8
4J/z3DnHAAC7XF1/zXH56fQxVlFt1Mg+E136BsEot2NgL7+dIgH1QORx5ouP2Zq9R+qfc2F1jdUZ
rdiVunfAe5fFjawLubyX6yxz1NSSilH/txBqQIFfmDBD811SryvWsoUgaxsjTDaMRTzJfZKbOp2J
PrCLIZgPpE0AHXTFreu0UgEiEL48SSI7Qbizotd3KJYAJmwdfd6nJae7ba59hTgq2mX2hxdEamxZ
bbjBuGyDaPP6XTL/9pSulJpILJFN/H7d08R1SOlInKTZj2VN3yW4fLxNO4dUc4bdA/YzQNylxQMj
vDZAZfH7BUG8vnECmupUh7IizgpyYMYTWw3sW4SKkdZLtJsodfCU+6qWxKt0cd/eHUvlNGN7Eqag
ArdRGcG3D0GVZRQYT0mcp2Yb8zo7pv9TMolGYUUbAszdd+ixgckY8mBMsKX2H4EoYDFP4Vv2PTS3
75bkcVJ1u/vKUQR1HN8NTgd9nvOyhJX/JvV34K/Jcx1Z6kLONkdG5Xeqy81aii0SpInBYAlCiVQI
CTebjCeps2wczMA/ksGu+7kmGcm/SYpgyaFqBMlCSlWXd410RhuBbFiJxuP/jAfFXmNZ/x59k2nC
snA7kB4GrQsCmn4nLk+yZA8DeFSfljGWgDk+GpPzdy8Hu43GKDAJK8+LPsbSNpky3FWw0VcGgOz/
PQWX0Oiud8NscjwGmVlskOzWe83rpRgwsRncOjBCoUlR78rQMN0NzZiSg1TCNgC6x+Mg1xEEY4yq
Cpw9kEX5clF4El51AO0nCg9d2TB/n7u5COHxXhMetYw4ZZEHHZMXmFSOOWStQv56IaKWKuHCgLED
kRW/zbEygvkVZRl+hMMjHkHJsTAu+MIGWXEucHUr4ZZ40OFVm+3AnULJnbUj8ic5a/5duEJoOs5v
mmONBq8b8Xc1S8+MCRmRuNl+H7RnPmNsLgonLfA2lxHVQtDg3Bw6dCQD9eFasS5usjZ4MECagBDD
qrT4vCrBYhYr3nlmAxr42fqZ9wUuxPqsGzk0czb43yXW6T15jhXrgfpe5yCdNROKpuX61NMf9X2j
V3JiteV/kuGWOnM5E/uPO0q84ETQyzGR6vDUqWsEJycviytKn8J+4vpcFVKqY2vcLdRORiaUnVNu
VMjRVh2LhsioaGPl9n5pPC/ptwhavqBXp2IhER0iL3TAyZ0OKZQtNSmVtQPFdR53adYB72jmpsNo
M/AQCnqmAPvimBaxhJ6FurgcnQuk9vy3cWC9SIpaZ7QWYRmqw6TLsRCY0AD/5L+YethG22OHWhxP
MsbFgrA2qsOkgsy98jglGhXDGbU/0D+7WcUSk4Cj5CgFqwVr6E5V+n+nfFYQtc6r5qWAdBAEHoif
FX6AkvjzbTZL5qheCpzJpjbN8W0v10NoTjV5CrCVqBuDRFG4HsFiqbS13hboxUQ/SUo3UJCcd7g8
yBQ3fy09CuxB5lmWJphMtXAI6nQZ0IGPCA0iVkxTeDwu940SWIBE7kA22UXmzi5Vi8OkVJ5hVoIB
AV1zKlxg87MIYJSJoa6gEr9tODBaPHmuV7moPKqVS+UGI6iZoZvLuBXnUG/znARH+DRWkXZD9KlN
C+EPSf9iY8lDlz986bQpj9BBNY+qaYLAHmaTmjoKLaWEVFk7QGxFGznFf06x+PIa1dAHAq1BmBbF
4xi5EJvy4SsU17ZZhlpNrMykcYr7F3Z7jMMc6wGHOa66AkIEYnaL42AEC9fcE+88xppnr7oHGZqj
sMZkUWcR19ECJO4rlVn5DgCLHTBy1N2U/pDWSow63Afq4SxwgRTW4JSBP7J5scdZq0klEhQN2NGv
DPq1uNCY69vgyx6USm0z9tvutxaMQPNTlY/My+fe8pV4tc8V71ZBP45bKOysBP7AxeyZWA008Ako
gqkaPQKq8sOJv1YX9sqwfZ4AnhDMXg30NvCl7QEwkUAUCbmQwJnqTxsFG7/e/ezs4C/7K9kzlzoS
LNzfUgFkuNH4EDycYXdi+XeuYTC9oqBaqcTBJDku5KwajE4uUUsIGAex98/TSKS+uq9HORDR8J9Z
lZ7ZO/KssNcioyzYaaboIvVDZ4C0Ij07sUWBlj53KECFPx7whIC/pSP19V36n0Jg6JgwQcrh2E9U
s4ZBhXWMJrc/BiganSiwmKa1gsIY6tNTDP9+o4SE+Ua2HzzvXhBPJ/gGHLMWMI1af9E2/7/pRb/C
7wYAyLbbkp1koW4+a3zCIopC33Vq94VWzlU+5zDY37pI1nshOi4pkV6zNP8rJzTBE+EnoEgzugON
EC3lx2PEWEOEEhRc/NJf5LMgngsBNPKTLofDo+RPir/gno4eC2XJs4oxWlDkZC8m991b4RidQfBS
fATyWVLCJORDELb33xgE30obeCFxkQkCub9loXqvdO2AqDl1Ok41fSLKnak6Fi1lN3faj1GMm37z
Ntq4rv2EonFOXit/GGgKEhqycgNdENEb/00XVVTJU/wA9xOI9PrBphWEroc6ueY8UFJ5x45ht6C9
rEw3NI3Y4BEG73mm8Y9Lid+U7W01Ifxcft9c4zqrlTN0JD52dqVR04shNjnK6IdDbMb2dGPjtOvO
W/3dFVXEFqNfNuwV/bXfgDIDOLHKeHFJ7hbggl+boZmXZN3Rz+cvfsFOtaygNhgkOWnMCP96OtKl
zYbJec+QgzM5HqtOR49emVi4E9wRdt3dih897H+l/PBgWVmngS/9JwUSlm1nHAVhv6Roi2YMfm3y
SALBVX7mBqxQszHMdqRje2Jsdq0PUdWkWQWOcU9iPbXeWOSODCKq8XtwP0yN8deDDDNvz6ldEgiJ
sNOb5wLEVQUY+nqrEfsgsvWVvKCF1d1YMq7OrSEeXaCHIJO/G597UfFLtG/SeCx3XF2mH/PBW1cp
RND16tR2jNzoyqtYbIMP4sq3K2P3EKIxfAmTeb9Yk30HB8056wWmKR61piR4vFcwaq8IosPBrs7W
RaS/cXUzQYqanO1cd+Dbcr/DXTBoa1eXOM2lJdxQxk2UXaujSaYZSt/1DStuz2nLe6n1hh0DluYK
oOXKIGrpyJtXuFKKNnVegkqW7bm6gysf1g38jhYeKjLHV9aDQMszXHXYo6mhjj/yPC2mRGANP+UE
3b7+ahP6HD9kTtXEW6TT5dAiXVmtrGP2dEtkB4nXfxdsKSNws19zCpTkaj2PpF0AZacLvxscEKrG
wWQG2yzs0lzAkP0VjBhT9Gs6TcuUi+nWv108sOaiOBy2qUToBTniWbxebZd8gIo6xCAsx+1Exv9i
+YlEekB0OveJZaX02LimqmEdKu1QtxzS3MVqX6Kd1YmCTIHgQ4zzpmx++rsxHcyuYD/HENJ/uEer
+8yIjMWVXnQfWPI/KSNVBiKDYcMK5QcTyi0eLQV/1yJ0zZv3SV057/RrvSqkT5Fp7svL1AWmOty8
uGpj8jhJ5okK/aeJNt5iGNbxvMHEO0yUDQhbNgKVLHD4/GHCpmYYjKKPssIAIzGyRA1hqwHFRnSC
5A3wIB8oNBkZlwIV41wADKLnEc58AOX2IPMtbdfcHHNn16bpiHoTb353tHBMehecC2loGVJQY3dC
72ILQEEn9VjObM2hIoNbfc/xwQiPADBjw4AAI+GH9YjXwCfqJc0tcVt4vmN6kOhNnX0sL9dhXSH2
PgQURvj4pl9dmm/9Xvcheogk+xpSuEnd9LVGQQ5EYOHeom1ZPB1Y0gyN3aoiG5mShElG/SXCmxns
NP6OS7r/MJBegMvOdX4m194PtkxtnyQ6/3vhgVRP01jXw4IX+ukkSXGWwHyS6MEXmoUAHYWpXzWy
6S21MHYjKU2l2AZLfX86LkRrMA9SzRGakHhHosRPM6YtSJzD22jlvPSpTdZHzyVQwnPQN1u4nUhn
MEzyb03iE9dWbVgl8x3s/xRlEngErlGJQtD8aw++lZLFcwHTRK/aTeXnWazVrEoj0x54aWva8ASe
vlPcNYgz0tzXPj+t0IwGxC2qlJD7xBB4skFNeJbBRfM+mt114iik5qAj9H/EzUDOENBiUwQt8n1G
Yct0L0YvKTt91C+qVP/LAqUJjciePnH+8RT3JYbtobd5dzd8pFfN/jD6xAO/jDc+cnZ6X5Fi6el4
L7vZtAbccMEmR93uk1ZOoSUvuE0Te1aWNMRtp2VEi2iWUHTMW1PYJQiFDOWi/N6vAxTX/fkcwR0E
LZOf/1eRXmsCpunY3wDIIRSGe1RiD5ETGgv4EmotHHu6wSzZ3VKquvKiiqwpvjvDmEfuUFZJCIDQ
F2w4sf+XZBSYgeml13eMjBKmlikVrtfLz3tIXEEAPl/VNammdbdb0wQOv9BRNvOsppoCkEaHhCNT
x3v6IVkYT7Y7aCEQT1gVQtBkvJVaBwEWTAoooJJjIBOcq9yp4BvwQYUWSlY0yb+KHNl5lQf1pY9Q
lmEy0nMV0Bqdmg4jUpHrFpK6utWUkiahcpcGvHa1gwW32YeWjq/GxquMAW7zTs2O+wkj+NtGQlQE
xN8BgKyIg9SU0tCIxgAUhXLMevKQlhQzbihTMtt4+wI0ynh6sBL3F0ZepSVettP/TJMQxb6y40dK
IShi+ugNzJXAqhB6pra2EZtvKf8fy85oqvKBPoKndY7cy3Yc7JsL4WtZrbSlzjr09HsF6rdSBU+Y
BSX0fQCWWZUIh1zZVYqvRVeDQcRbEbIozgM9VhCN3BwwA8Ns9vbn5M0TFCl18ZyO89oi+tgXMsWt
OKt3LcxGwyPByAfvp3BNzkWNme8rt/dwbRuTXZ9orZCWnUBmLfGOM1Bsnivf7HMWfnx3q4AQyVCQ
DPOXV++URrtneHU6H7voKPw7aOY+HdJqrYwPCe4qyXlNR+AWynq8Jnk66PVBMGNUQxd851dHnotg
h49s00xxZZ+kF791P2Al0rP5V/Z26L+w76oLY6po0NZP/OOKi7ZgqCt1/VGFj+XK7mXfuyaJdFSP
guEhmTxU/zveS5ibQ3FqMrn0/CCXX69rg6jepgpB/4fODDirCXSYfuzy+B4JKmq8quN9ZKcCLxf8
NxifU+P92PfO8uljWJOumLPzNyQ9N5/wJXv8L+EzkSSw5bMvN67+cv4ZdEBDs+72ivO4dENI243c
DXLbxQibjUbXoc4ynpvA4hRkNxndG8Vb4EGZJgHZ4iZGRpU4PEqbMpEAaKLR8Md9AMGpo+iZpirv
L+YuocDDfjylBbDIwYxgPL41ZuLBS4CHPjETgyYvXhA9aG2pR6LkjP7crWT/3ydjysZLTZKiRXjx
3674ya9gwYAJ1FJdtk+VQz6nFlDGVCBYpcispu3B81d2HajyCj5sWjCdJEYAbfObW7v3FOXExVrb
cAY/yKOfxdQQiuc31R1Xz86LGV2UEU+PxTMWHGJuQVC4jodxNyB5OzyRLMvIRYTh63+C7aZPWeQk
c9qk9jwWYXlxwLPyWJ7CB98brqBnp4POcUKlEHprhoahrmFyHsoK5IUJ02JIfZ6pJmt62kExkvni
yQVBdRGArhoGZzE3j98BkfI3G2lsZjzW7KNrSfKz4ycE9jxQ+VVC0l9La54ZjkJMiTCU+yMPAn6q
diTZEasmnP4+6lOOYdZCTsGr8nYRKj9tMyXKn8mi+2mDn2n5dVQa133nseKzlbaimw3NrMZJ44kX
4+SJAFwlAddBQw/jNSvvfO3QQnG8ZSYYZN/vTf1v0rPXynlCsTjDmHKR782scSQ3hfGaq7Jwhs45
G0ihPoT+euXMT1CNf2w4MnENTOGnJ9DNsUXFMCy1YhP5nXbZHujQ2rRRfSLMqRiCxGtizQb5xzlL
ne05pu4AooDIpmrj65pGmsNSOzBD1geSRckRyWZYFK7/aap5Ljdd8Smgqsvu5G4xQMZAGcsiSWAG
hz04oLpbkgdCgn4gfVIUhFGYKXALanXLBiOn4Xzo5x8NpxMuCEMeahRS+pwS9NTJDW6Je3dgjqrp
o1eXEFoo4QVYWNXWZy+gtLvkTECQ25LBzdwzgUmqaIU+HDvoycQwp2YiXly0uHDUdK/G7AvND1S2
294i8hOqyoExP+Pc9hFryf3XCNvDbU9JwMjIWy9bkmy2kHJDnRFzm+JCWO27Otpn+tLmxjxcukg0
4zbfRFhYmDS9WM8kND9MLorexk45Vc9prfEvo4xaohHli9vYyk6S3HHFqXyHWH4ZF+rbMFCBGOjd
z5u1k30QnZRplQBHcBniWHEZ/O3KyEaPzt8BNNe+iBMviHilzUIBEZo0YA0nABa9LRXMlISL60wE
4Vc09WAfKD6rcbAN1+hR7qPkxhfJvKGqXLnD3OJyGak4w8UGvpq8T+gzjqm5+qPb2lOK4zOwWA/S
arQ1QwJKxxSuU8VwQGnjnJ1m6rhYSpORmZr6xQ4AcuZ0weV4MysGTFq1xFXskKcAP0zUGm5QO0ty
rPbkjuBQcJCB6oeA3OJ7DqJcT1twoZ/qmnTwXC69IeGi7IKgVVXtOhjveKBVojXFYXJbhdLzoARW
u8iwoMn9rbem2T9liruEh5A0E+gATRg7TpVhi+BE5nGD6XI8c0nG91NtiqOPRIR46vy0YHiXR8/O
7GwfRYLyWEL9QYZIR/uPlPqrK6Zey9mYWk7ADL6khxALks+FpOh0CBPxdng/Rrg/WxHnAcxsrzMl
W/gcS/Y6q1e8xbtMLQz8DL07LiUo3MVrCT3zj42rEcGelakgnFRr8l6hckeFoOxp7GoSXsmCY9dd
k6N7A6eJbyfiLUa1RSJ6TvVzSmExMyXYJxX5YdiA0gRkH8VVuLm9wXnniWxhIDgBcjYkT8U4kxre
R6HQpQO5ZTPlc1ToQvbd/LwKtinucokzwPW+mVN5HVLygQGkNuNr0POb34ELaFgxPoZP9hTk9GVh
Knixl8ephcOvPIbiewokXwyfwzFzF/Zj6p7Cdnb2zPbWOiar255rP43cHu497bSUFwpglK9XYj5Z
p8fjQkfsCBcRtpbYgTRekBjLqgP6he9ujPcbaSF1rIAA1S/ZAcyrKg/oBhdlU7duQiIO/6TMBpcD
kRj7dBxXTJq34pVuODb3Sn4m8S8vELBeCmJQ0M3mRKvd+cgo3G2ujgLpA1xVL3fL4qHGvYC5ALpF
TFs6VX1vnUyFgvsqs2azFKKKpi5d8dsKDcNLx8tkaTYX5D6gLRJELdFm2p+B83BnHCaF2L4t4JP6
tGlrX/obNBW3bQbcdxk4P+pYkuuo+ZwaIUIDDOHIPnx2GLkQfQQT9juSyNX9qdQQLfFrI819A9PU
VfwBbmKBjZo034n4LOi6NVseNNMW7aQzlYwfAZXYFkuZv69u0hWukR1175as0RA0bsfym10Svlf3
jA9p+aCSkEBBidkOmTgPCR4sEIH0hosYBH9iid4c26CBu3/7tEequS4OVd59KsQczqWp5PAmEZnx
LoQ0EPMN4Mt1c9xwP3TWIaUcYXtk+bwSYOelTwt0OkHBPR7WP1Lo55ISrmqfERGqI/xvIP+yOi03
+w3OmjMHsu1oyLUh35T5ZYdgQx61IR29NDBhQ4045WEWe1AJnhAWQJ8Gg9H4va3y/3+w2a8ISKoM
FP+ojjiebHt5NYvJ0HkyrBES/VWNvFPvACl4IRUcZ7C9dSeTJD5lT4i3Vd1COkx+vE26O+wCL9gC
JHyOV59s+M4py8ljilxQjag9SGa2RKB2kBx2PJGb3Mxh//xrv3apt+/TftUfcIv6Wpe2pRKrUrvB
IqO7j7HUyeKLjVBIYAPUENxwd6I9gynSwG4tseVCh0tmxl4r9CJtRvXVP6CZMsR59VT0YN2jyXsX
f2eb9andqDsqFLDglqnYlUS/O+xktfr/9/jHpoIg46zwrcpQd0V305F+0pSBbDdkUD2ZoEsr6Id1
bdsv8ubiSw+qv/lPaEsKyg1km4VjBLzqZJlXXJYaN+cGEK3xHyZLX43evhP2ZqmqPYaydcQqVyA2
1y5dRUa81Z9agIG2GUqRaeccwVh+j6RBVCSMrhVN6vR9YjPIqdVCs4809vp7+gs2Isix87d7199f
HsXZkfFDsOnUiglOCl0CWt86S7k/9wtoz4ifZ6fRk/TGZI5kDtwPYjXncOamhGXOwrpwyAA/yNee
XB6nylaNMlRli/wkgKZOGUBaSDLH60ze5LDLXdlzMJwJFSsn1t0bqrY2byQFX7RrOSj4iGriJpHW
o7uJCFfeaHyyLsIkY3SF9z7lCNuf+Etk6umbYEqZXwo7e8XfcILeUE78WZr+GngEjjDyX2phjotP
bNJjBADI96QhYJdpIYfqWxc8mwvp+OU85vluTvGKy0jFphVKcG99MVrEaHH/abOzaTHic7MC/tCY
8z0xwunnR4jdzLMYPs0GWb6y4ncURon+u9VyATKoyWHZo2yeZQA2s5lW92XLwwfm3U/XAAJCxwC3
MZkxVmc0HbXWoklvmxq2A6y6s+JDhUq4CE1IWOLG3LH+rOnWrFbBIRzsX2Q3cSwOGflEFES3JBBs
mxZQ8+aU9InTG/stqGFPbzLZQ2GjNkI2oPaQkS8IVCROYGLVZryJV4PrkocicSdmR9fBsmHzZXiS
MRfKyf74PfTKs77t2GYWOugr/9ARGCE52ANnymzNX02rYAVMRJLelPG8kukYCZZALLlUO/q/JhCA
myQTJ4/mpzfag88pnoKbd0V7VtV44+xIVw+6z0pH/KGHs1QXXSnjoG1E1gJQ7Xrs0j5MrENqxt6F
cSCiXMDhL69XlKB38q5ExWPMF4pIGOq9hRgI/1kWkMbjlorrXR70ztyEMIU3YpGKo8SXb0ZSO7VP
rp0X3FDaGUfkEHRbrnpPBQHTVdY5LnWLKGZYw59cL+Qz1nDdcfO72XHgcN5+ipO0D2xKgTA5PUen
djHWbuvQYSY/iCO7fUkFXSjyf5UvFSesX8eqpLos/yVT+4t28m2aoH9nK/JTxwLz9hdx4akD6w8J
L9jwMOIOWoVHWoq4w5DSJrh8Zm7VvLn1u11JuyQoVj6s9C5fwP7x0vXrsqwCJZQbCFy9x5T14+vU
6Hb3s/fkN3rQfdT9jQbM/M0GNSmX5LW6JFFgaE6C1HDPPiuNV+BB+0KB9SEKVe5rFJHBwicdjvYo
KfVx+e0aVZNkA3HhJMqnx+d9hQ0R7amsQW7KmCoJuCei3uymbyqKz6Cxk0N7+jvh86xnzKcwluPf
jHLrEIPDtGddhjwWtbgNzQsFPWKstqspuZPPj9r2efByRzsDAT0ymaEfgDYVlFEr6Ev+BEbnnBRV
lQIA0qdVewuWAgZKiaRrn6xS1YnsioeHxp5svs6JJqWIYO3lHhmuFyQgvPdErsURBixsoWILgotE
2jrcP1YxN9qn+MKSAgopldueIKH7vtP1XkL0vMRKNHjUHG1xPbQn0IufqgadQJvFr2g75+eb/s2/
FFyg48yj29guu1MvFxReZdobi2bm7iA5ewFOQV+jOheUQFSxxpjQE5+rzt41bQXAaWTCl6ojOXjZ
fxYhibIjTUqrQY9j0NPSvchMnr9lKKU+uGowOA+m3HbxSr943oTPf2t7cLFQeAA1wYKyHhauOSri
1fsJsn1ykABYyLb8c4MMH8MQ7EDz4Hm7PfvbnWda26iTAmcUMLNQ8BdMzsXH9pJH90h94zU5sMCK
GUmCKgnFXFgugJr5FpAoDAEIZ7ygAa0Rr8nBxKb9zO2g52ocBWNZRBdw8If00Ti9CjqcOInhUjyB
vxjFyaLqqq5AZcYeOiDH3ocM8uBTXd9fG39Eb96Rvz1o090WKlq4R+aViCVpyUkmquj50dTU0vSQ
/VAONZaD5VtA7FM9NkXguNlRO45sL28ZdKCf1t8Cozn4VVSGGLuOwtkETPxbd5bpVKa6g4pGcruy
KKkuxciTsoKjHlTGlcwJ2LH0JfIuFryq9Q6YDP3Oe1Qhv99vR+h9Z0DEy1RUXS0OEkGVmYCdFfzz
deaw/VmsziQFULEPiv91ZoZOOxfhS0L1XvE70diOx8M4TOXDDwNiLVR5DIlBuxHLuJ76XvfSK3i+
zLnM80QiwQajSwDGdBqhYh0k42hFQKMykqNmZdpQaGWiFHJp0QRvI2Tf1u89jl/4jro+9ZMxQHSa
INJ1t3Lr2WvXvXMWhdsatFdI7eaIvINgrEJJ0VNy3xrZ5CG79eLvN3t7bj0MdTmkRyDoJLWeoh4+
xs60H+7Y2t5u47eUBY9DBo5ouxWTHyVqQDSBsynnl19LVPg8MINIoo35Fah3DtwK8JcsNY4Bot2y
XHa13wgcTPSEWHTZjhEinm8hyI9dK3aE+0okE+6rhOuSiP2hLUt6rQU8CmRKzk9lrjjzZe8UizRc
8AE2EZw+V0ieG4oGkzsRmUJH4RHr8K4EAqmwcEoEp4VUQPQC87Pg4VLAe6O8mBWkPRDTZdB+pH2q
oZwBagE0rEB2/WkHpeF8yV6T3QM621fgLe0iV71Ohr0vp6gMxzwdzi95T7q30m/1KWVEotJYhgPy
x29GxkAhFMlpcgTPpxJ7tM9j4yYwPaLuvlTW5GU7oexIAQKpoCv2sdjFKLwB2m0Fuzvc1HRA4m8B
j7V1vsBYdkBjrEiO9otLdRCKsaudbAcpP6r2w7kwFTj04sLUmSPxEp7L8xv3oSsROOluULnXaO5A
eP7B5XnyjDatTp+UQy8C58Uw2JinSzKiNjJ8OWFPKpp+8CyKIvjhiyPNh95kAkHlAOfM9HxXvHUV
Dd5YVm0k3p/qruLq8eJY4TsGHY1Y8iqsUPFZgZkAU0TvkX4tvq4eBySqDPtvs8L2yV8GHTCmtnJB
KlJa+SYcOQ7X7khhVL9SfEoyUUmuKk7eetIj81Rt35oc5py2rHFofo874w0Zi5kFreZLnil2ySxG
okVXMqXqvg+mp3Qj+XaIoCP1mQh3kfdLfX0Jo14OPG/bc3eA2GuzmQE6mmIqQrijJYiEMR9nIOHi
qKnK9OwraQB25ndsB882Bz0Z5/eWxouA1+Tr7WxVFhYrJjMAXTfXg+kT8chk2jhhewosWR4BF01R
F+Dq4N7hbqRnTxAVxwf0aN3tzZ6gjyuR48e27ee4y4JaeaUFsSd9Jh4juTVqlM4J1OKp+DnkRsKL
oWEdi03wPfZiqZ3CGlI+Cc3qJCObDWXE/Ke5rGDIsQjKyvCIcf9IuC3TkRFQS635bJba4dFH+oUg
rsoB2xew3us/QITj8eQpvzBrRy4XDqmQ0OGvsXlg0omw4YRLqCkOkiQwVcw6kPh+0RdPxuUTDmN2
xvuX7Z3x2feYTonWKurVCurptA7WQ/Hu/V8fHt9+Oe9DYhO1mJMnk34EvgtYBC3LW3VkrRinVZCG
F6T4UvR0LkMcJyPqsDsb3hOlmSsNOGslsC2jCRcXD/n55FCvSFWWxcslZiHGVABN03WzFN7uvvHO
UW66mnbNtltIm3zf0zmbIgFa/6CvMvriR5IlpunX12MsDK0bnr0iDt5m1OJ8KTvuQve+EBzIYUAO
abJb0Ak+t3XeSqT8Qrr6tsGUkKXa/KKCTySTid3+t3sui6Sjl/RuLtk0T3S9ChmF9QupIlSgsojy
UquNeSg56v+YoWnMe/qPopf/FFarkeyeev9aFn+swnYt7S/Cx+xGYGU5++KIfBnuXdQvz1p/3a3q
3ZSHMoxd8X8n9PtvrLjwKSt6FR0Vq1Mgk6KufkXoIYGu0kdlmqJAuP2Bw/90XNt3iFIvoMaJArJK
YAJ8gyhHXYa/w6vgR9NFOOy+Q0c2ygNRjvS3X4CSlxNK7dj1lCJvEXeauML31v6DDr+Y2T8lJeGq
RDUT9DesD0K5BiRFEydPUKG6CJ1aZEhPd6Gi2CDv0C3t0zYXYxdAkIk4iV9gRZfISOkO9wygs0PL
wFah19LgtNi2x2YC6zsPLD6pk9Wkg8tEH6xG6WgEe0qCavKO5JV+HBaZuCG7yZ2wLZL2wQ3CZeav
It1NMC3ahmIHJvrgce8rlb9aECLd/NQ0naYAkjEAbblYf5Y+oVA6TNNirhhfm4g4gaMA4ObwR34U
e3eICEZavVsksRl07a1zX4M33wF7QzvWj2+ldu4mddQVHsqgt/CLSvyDMhqRPeM4sLE/V3hvnouS
jCteHIRGeY3vow0VO+PEleycGUKRQfprOnW1pzHBZ81dGa1yPpxmvmusINBLIdlx9RH+RhzTeq/k
DbFpVfhYl73iMvYTavskkFzCOD1k6R0MyjENtVodDEVHqxd5eRExvwrb0tk4vN3UEeACdReXHC0a
4179f/lQd35SQ77VUTZnencit6sJdwmWtY9Nq4BUdhCDBiTqPBTyGcc2r7pJ5fkuTMAiDZMw9k4j
HrzPyYGLg29XFB0fLmgjwFOa1P8wyHQSI7rRkfQ1SKhsMTuYOjvjzW3kXsJua4pGdi/OxiSv1HFO
gPRVyW/j58/zAw0x+fh8x0sk7edFPItssZama+PIIh+Hbmur/gn56TB2LYUDz+961FEdEpIpoNlB
dYCXzuo8UQKO7+CI9t4NfxH970nmmnd03lrcIlWRRD3ebb1KSuQPn5DtaNIx+V5vOf8O9DcOBeJz
3gLJSGiF5EnnEjux5XdPrlsMVY0DmLnxKkqAOSROF4HUkwxARsSSYBVzDgbms9pIKdGZSnwnids6
UO3A8wu4BrsFTS4wn+8kv5GYiQZrniKGtLqDPPAqekwQ4NykuX5FnziwmlvwB96yKsNWN1rlskwr
jOAVkzWUmx/Jz8+3g+9DmeVIQxZVRTcrEJA21ECabZU5lYQcxVeBEI9sjwKhU6+FXWx6Xo5Hrsay
VLDCFqN4kHLSQBZb6UGH0q3A6MPJ7K516+E0IHWxBGmvVxjyjBX0vBMYZx1KsyZx2glcnXG7o9uq
1GiEFXJlpPToZjJA3BPMzQ07kKfGhblpTnl+G50UJrju3pua/02KgT2nrjjJLbBoUEzdg6uR722D
fIoBK1Uj2AU0mTN6cPxFae+L3e9tCc58X8si163OWYsOxHEJZDiWuY+TIUXreMf7mMvuQyvnlsk2
NH0E5iccIZT1Ex/khaw4ACF9NUXEWX9TXA4kRemMCpPTDQq5VEL3reMtZ0iWEnMHrdnZY+c+Qaxv
N3c6EqrUEpYg/sPX70uU9uiqAPHnRI5ESQmqQa6RsmB0wIqm9oup/yYkUsKY9AOZfMQ2eKcse4Vx
IqQM1MwbMaaTelUJgyczXLH8lTi8NPJ8pJ93HX4wP4yEV7Fr2bj5aL9KoGWixHLFBsDvyQnJPOeM
nIv/BG/1DnfBOE6R2ULHrsJQvh2YnKcUaTB1pr6qX8uAaj2Hw++tlHIuGe3D6O2Po44s7OWVgfs1
ujTHrYHmrxnb7Rwn21sxfsnCztl6JfTeRlCRrq2zkVHiyDsSNfdfPHogyHCe0BgUShiOZFEFvD/6
Ifuo6nt/d1O6EBw8ftjuR3Ct7hKNrZ7BgQboaTBL7RNROB8vo1LPCQnOeyWHl59yeMAX+FdbCDd/
lgaI02Rjf1mtG1wXjurVPGFIVQTIfSvO3GC0RPvoKKHzWttbOwJ8d0OnP72EfUUSjgFTMYPIVJS7
KdMGLhtFoPIy21U1eW1KNN+R1nD6gC7RuWHaF41vxFCFn7rdTaSbTbHggU4pN9JEh23KnVgLFgkG
aVVU6hxue01hQ9aMOfZvTCKgZP8dEcFQ8RcvmtMsy7QQuG19bC0AgHzU4QgrbvmADyOo08dbj+UX
u/0WCzlkXp+mz3KyfpFyE6dv1nti03+7ZmeqYSInwL97mGNZUqRGQsBxsOPjFjE3Y57kZYDOMkM8
9s6z1VK9DkQgcunb/MJGMbxkn4kUyZeI3T71RUsyJKV22fWwhZE9T+aAww0YQ0hPWnxo5Y1xIXrM
OMVwzfscEKDNLHZcVDTBW4QVX4pXAMActY5jincRxP+gianWafdCpTjPdE3MQIEzIWsE4jFap9Fp
7QaUI8mAFxpNmnJTorYNMM3A3G4D7KfoVqbBq503Zz6FvnaFtm5ho4qab5FSyCVSyuoPLtyrk87p
b6l1pE9Xc8t8smaq2lAtLi35Qft/k7s1Al9WSyMJx+zVrw1gX2K5V5Bv9irsfOCmenME9BYb6J1W
lkTFi4WZtxbqZUAyFFLv9aTla5aUh3YBv09dTgJFCug0ZojFdQHo7Q0mvhgw3pmuMdljH235rIcw
3gW9OqZvN1R0dshAXbd9/3FvbV2V/9wqzuk9fdUgpI5cSkrEp/Jznq1fa2I8wFwpxzbA32u+x7+Q
2TzENW5Oqyf1h2Dmi3iFeA9Uwifuw7coh7HxvRhAPWrcajYYkR9c/rlpW6Zx8eXK2Kiv+BYaD2W8
hhPz134YxKL7fpPgwwGvI3tmfFRFVgRI6H9Vb0cNfdsF2/LndsK8vrDWkhV08/JbxshPSA6RpQNh
pSmBt9TsiYb89WT/FPuFJL89MhyjWnmrVle9cSEZfsExN+TmUuV6yN52keIGe1HxB2YXqSwvytPu
UVCHqNvylRN6zYVgCj5QUbJFHTe/xrakm8/Tz4SIw104CaPBmDhQJ6RpM3dLnjlzJgoyQM6klClv
QhghDkVloqE9hbCwtDaipYDvfQxwJtYl6cpWrvnH4/G+obdy9HQ5KNcZ5MrmqK+UaqOMc07U51IH
25YtOdU4K+GvO+SKt2LHyvg5Gb8c8jVXnxyEkyr/5Ek+sOmGNeUH5mhkEUNTUyCsGekSJnAGYjnx
sqB/QGcncAqI/5uvWfEgX4Vx9VKCv/+1XqBVmFuI7T4O+E/aKsIlVCFU+m4CKuMGaf+PVmEqWIoh
faZ3SP71nJper2LQfqN31a38L6ASCsuyOizWs4SLYaGbGBSD3cbV8bsjCQpwe567ksy1in6QZ56e
wstgJkAgeiPU736EjfL7gIOSSrVsgdsQ/9GJRCZDijmK5+bXkRR0SDBeZZ36eJAoV5lN76qFUs6u
9ETwdSFMUHfyvr6EcU/xEHbimayex9qSo05oKXw0/rhe2nxCyKrsMGxn9jTL4aSagDvoG4IWqMlr
gcCEcTIJVKQ8qeErUZ1S+tnM1/cwI7ka9Rqhg+FYDRLeVlTRV1UbwRawS+wLN39L42DEz0GZKGuw
t1zUPUKCFSoRBTMIBEmkqvyOJQoT4/tN1vFS5Yv4QxhDzVTGlXunDcGK7QXsaVnaHIneIlvlwjeA
KAk6A0YgFV7ne/yAvMtcf4fxwcAU9GGLxxmeugNzl50LmzWkoie7pNYwNNyE59qPl3VPMxUDk/P6
FpMOaLx7DAPOCRVjLx3ZnRElt6rRemGBbgkkewd5aKr+uEzQm68HFg2njfrfKcS9i2dQf8HxZDTZ
YzmLFg4cFisPfr1TelTPBpF/86F6pfXgFA7hNNxcQvPxv/ESZx1Hvb9NBbQZ8/cR1y+IUq1dPdKN
6/fZwy/Mv17Q+QfWGOLDZqlTiIBhUeIAwB3r4cym3hx6bNxBOtptfhS1X/yPuXUo3hfrO2maPyR+
AKg242CA6O7Kt+cSRr2VTop/vfeTjnkhnsiMFSQmzUR8lGr52KkpZPvI4A8Kwocau5X/KFT+JG1m
239k0J9oBifqZx4GXxpzhVEz0Q/gyZcwks2co1chYJYWiztD8ynw92OZSdCbvv5h+pglNsHWHoAB
ekli7ByWSUODk/FbXyQ6y1hkbicPPfqyUq0O/ahcJPzf4osMaGYJX/w7MJwb135HfW97T8RPOqnb
P5sNiTvU43fzAAD35pvq8+y0yWE86r0EuZovWYUzPQaYJ8+f0L44cruTdFt5SftnMiHoNZGF1hR+
vKhN1zscgzgaq605XwdlYbVIDjFyHpuQFv8nWPQFD+CEB6KThhInpzLMY8/y8ZYtiOq1vckjDsH9
uKiWJg3wgXIv6l4Bo7+tG6O9IQNJdhMGycr/VimPjwYD+U0H0ElnqtS3kqRjYwoRE6UIuuZBsphi
a50EKtUCVtZHqO0RSzPKacXnxu8fyZRFA0xZaLz+2CniRXao0DmmyN9xAS+NWwTUrQ/0ZElHtp+t
ru0CuAApDN+FUIhaVs2/dc4VTmcEDdLX2EoCgYww2TKO7ZYxWADtCTKYNNGNRiUDIzhw1fvr98tS
ml/ObSrGvW9E8eYUNoDEkW7ODcX4a/gAHnjTgqyXVDDWgXYoKTVYuGw8WEKRakiVX6SSUTqSZ2EV
L9Fmm9l+H8nbzR8EYuDTB4WPjLA0UNFwC4jBsG4EqWjHg8naPPOcQfwO5L3fXiR8UBLEivECU9fA
cBgIux5foTqWD9K9HFM2zQkF6bg6PILiKQ9GfW9hpAt3QYXixNx0Wzu+rtOtqg1jtOr3K8Nt0ez/
q/qfv2TdfIdGUyXoUMQRrZ6whlOYULHCY+SzUy43nJc74KTIU/GPEYjPk3yieupcZDsep3cpMdvp
SBBdcqHDWWu0I2Y6Lceo8CIFTZbdqx336I+a1ypL7FwMUncAfM+nunquMXzFxpopbrdHtI1O+Ren
L9s0IFBchdleugxk5qI0p9FmNr+soRxB6FwfW2CNndvAAWdej7y7hMQ6iA50iiIonRZyBFo+juBf
u4Qf1gn52xtDk2ViR9bwJpFmTx/7u8NcczuoaQpq0rBweWzfcemxLSfxXWGdGXUgaF7mskkdrsHG
Mi9vSzmzSgmf0t4BPpNdg/gv5zPABLK19ftBircUY7KTMZGivBXusDwwb6BoehmraoPFGmQW7BvP
qzS9aHkuKOOHMkq46gEYThs5A+J3it9clvkA32aaPpYYPPWXoqFm5/6PQht1GKhuYD1rVEjKckSj
CDu39Xu6l8E5MD2i5D8hUFHA9IH75PpNvYDbrzIc0bWGXzhk7wLhWCKrVfp8lnFyu2QJ5ECtw/CX
VEs96uClFhgXf485qPcMw28ebj2G/4T4G06XXuf22MAHVDawmu7ZfQAwhltXlVPJrPtCpPHaWQ45
Nt/7hvQbIAfsc8S0wNCRFLjBloDzo60B/xdQ4I+3E9PE7g0agrTT+8e/MqQorYK2HjJMMxm3sw2O
jEDaxDbxFczZ1t0HB/dkM5DiAWI3qLVvhdQ5kTpPKYyrref7V6UFElXm22B4aX9U85GLaA4jxq/n
8UuVs9Na00P2KzZURBbDtT90inKvqwjqPzIVgfzAWP0I8Z9Y3o9IbCNBxCeuaE2yAWTBUPMnym7d
vpTKQOelZ7Bv7A5H4LC80HFZ7aZH7cDeQAfPKqZRhOL1MNbVX8yFOMZouwdTIt0W8ggUaZiP894G
XwG/YfqoiNQb9fGCCnp8bK99sD8CEbc5vtyKMMyqe6zpaah+/9IMiwKtS1iREbXaeVX0c1Biloz9
Fs91q1hbswpe9MVBdd7p4J8VzfqJbywZYBemwJ4PSWV5eHuOz0xK3zHGvzYYVY7yT3IDqY8nX/03
bqOjjAeUl9GIPQ5GYObsEEnwHq98RdEqVZKPP7NWf7csKzjjUaixszevfUob8xzYIkSiZcd1c40k
gVlXmBg1IJ6XvDTvECroX6BNW49Xn7DTn4xAr8WAmjkfwzxwaV39AR9P99yXGrAYF6DCl0xyhajO
CeuoIq2vIyKxldURKS/aTTaJb/amqo/PjsTsyC4t8LO51sjGdu3ns5zdt9pq9cZQET4GYXCqAgFB
4a+D1K9GMQR43oboB1mNm+DxjrtbH1OBhSblZddMcYXIRzNYN1EU1buLx5wyEkaGg9lJ3+SEToiA
kjxhHu7psBmF9g/Zr2I3JPTczQCBYXJJS2TxGld9mvbIa/V88cmsBq+hcUO2TC92hBzU08/Vz0Dd
/xtO/3ksZKjaUek6edvQcmsyCl3XHF9IO6y6TYPQpC4p0wcgkMKyXkzxgbSEIYhr5CsT5tCjfVNH
nrfjnN2pnvR5pDaD3ZqzeI7olakSJ76eE4YESfcKEj9nUo3icEKoxbCQINWqIj7uBmLBhlplkOhx
iqvwF1IUNh5apdKf9cGJKJE86nZuwNPbzbqpYltcRjyl673fwq/KgiMid3jFv875KGMhFtbodYnU
BA7xbU2mbtBQzbbFj8XTkO9S8DdIh5hAoc/k6RuIW8DnMp82PQw0p+50dbyJtp5xlPhoZiwm+7Q1
Ol7/NohPaT7KiS9IhsjTiLRR5ST95yGqMncTer1y0KIxSJ7sTsAHbfblh7RWV6VDG7F+yUSTa1/F
BRXYm8LXZb81M9gRJg8yQS3DjJMKdB2O1hVH+oZTd9wiHwvxjtznbY3mYA7Cs/ISmik5GfB/DiSf
PN9KL9+2nWIkEiw/+ddegjtWUUXknJnWJ9x+VNosyjRL2UKfojvJw30HwcakoDdG79gfk1nyAjr3
Dp7ku4qoptYoV1hjEwNPKT1jhAMCm1LpjK63IAeborTtT1rmNZ0jIfGG49ISPJaVC0/qqBCow98n
6mcvn19bXK4wzLURl57EUnu37K4nmsxwIAvZOV+KeLPrRE3yRvA71leyjkADTXfIjrkCvJryrsXf
MaIS4y6T4d7ZDTv1NGpZV4FR8SjccAovbWJnfrm6kuhBd2nWENNHJRjGxxp7hibDIZlbUp3pAjuv
voWgJiUD7ZGFCXExi2uRMgITiTdh1IlzCl+GpqR7H4APbu9zxykzbj8mRhAmXljSVFb4rcVdbWuA
K9RRaIqs9pGzMuUSyLXfKVPtaOvICFtUcnHaZynZ8OSPBIMC89MM93LC7H036GOc/3cwArocbs2U
Bk0LN7ruVTFUXCGyJQYT6IHB6bBnH3XU6hNluZTkpI7UpC93pVNuBhWQeFHmBCPgWIaYI3uI9u6A
mVAiYsICsVu2WV2ZMwUed8Dcr+bHglpUR8S7v+/7/eWV0ylZR4shjyAmDOi1EbOMZjBKlcUmg20s
mPuTZXJNEpPs+iGTfxVhtxDf0yl2O2HLt8uIZVWcBG7OX5I0UJwG4ADuEcqO2O9+jUSv/mpwrvAo
9KQ5U27IKB9JJ5jA8ta3jY4CTCRzocZD+CT53FB9+7HnIlhGYx/29uNRcuTePjQOj/+eUsc1JjZj
xF/e1RscrgBSzky8Lp/nkIXk6mcJdmkKyl1Gjp2FgaJnMWh8/lNlYRH+eNvsg1PX4j7/rK97UcHI
kxI3gwJ8y2FHy4MuY3YIGBtAEaWEI1XONIZRyhuPHDNxoPAec60URMOyjUARJSLtDU864KGUyF0N
d9LtA2yA3sEfxwaLdwchmsHyI185WlgD0UOEqx3c4YceYumpoJNWAi19lEPR4qJQvqMq/b+BkBjl
U/RmMMg2t5rqwPUYe0B7TnYnB8IE9yuQ8MoZpvDOtWd3zEzTzUB9PBQysqSJ1CirBfmi4m09YdU9
iWRnaLOIYe2RudiWoPx7Bw2PSOa1PtxYjVncbMU2SXeOHA0Gpe97tG1MK0t5fp5aHy2oIs1wlO9B
SiPOy2oFcVGFiSFeensX991nrWF6AE6lRHbsZFgfjnIJ4tXFfKPPdCgy42y0xSuq0ZzeiCSoWVDN
d8b+Hubhg9gRYOK8fx+5jezaw7F1yKa9vS//d1ca2YulI74fGZThI52c8xjcqMVdQeylA3NNqRaQ
+pG1zBW037dBOHbfwbnANTS8zSFEtUeGxhYun0ALjD6JG+nCukdWHvUwmZnM+DFq6myQTDXtxsa7
Y5VbbYo9YZLOOFIFhQBzk4hhKZ7UxIAXMiWjMqwaO3fi5ilKJ0OAsUI1VBkoMZaNHibKqZuihC4i
nZHZxmqPjvEOHlZwL7plbv+XpV/z725s7nOa4V9ems0gCz6jsM/ybi2t2XEF3svLwM5b8wRTFolr
rH/W7WCTL9M39phhDx7TS/bTnKVJQKSm1ywdmud1mxdHw4DDdBKMuhRQVTjwhv2dLBSwI15Vv4+z
oFzLBMJqNKWc7QkKeX7jwnYqs3VL7xYxNRkHSi6uX9YBGEY07q/XYIMAMRKnSpjlIZkyIVsqqKup
crhYbK8rkS7pL9CCbBj5TFL0Xi5il3g4dDpophyIxuRFVIqZRyEkVdDTJFrVEkpZiACkLeeRQJyK
qvjvsIE4t6hXOLI26GFtqOuCFG1kf8lr0o04tFrkdbSwVKmNV6rwSucLmYK2p87NePPPEbf2/MNb
akPfpVOxn/+u7VYSqYptxyP/vtHvNnp1e7UJj9iOG77Uhu+ayIzlWdIgT166gzsrtuDoYdvowVlf
vraBaKd0H1xMzBRmJVv3L6FLzDzWkV7QKYEU8HTLszqb4sLSWDsZ+lGQccbxpuX3+uxst8JK2dof
Q1/tduHXNVQmOOpzUuT1gUlc0Mm8q3ecpwQKOKyKz8LKs+ELifpWYg4fO8N6e7cfiJIkWY8TmeEH
CS1LcBI5HGoLJkruZ3WZ07Sl5A5VMf1eBYslLYQm/hEi9u1mUA72tRLeYlY6ef+tW+79ywcgf8bO
RkeCx21D8nslZPMUm59pbseURnamdcmZQU6RgVql0RgA9Zz3RMqwmaq1AUgV+cwNNa19WD+shU+v
+aIH7XdiDLTW9AgkQv+pH7p+QQ7fNznpPOrsAE7kdAP3iby8Pdgs2byETF6dG+0pdr1Yr7uNHRwk
uxTJJ3fGtM8BWC3wKwaTe+vJwV3hw2VZleNeUJWZqE4Dhu32HtPK/8zHjqlamjzdX5DS0XAcLsbe
RVQBkXvSGKPJgCbJQTKvRN7OXJs8OPcctanxgiT0KkknabaxFeRqtsBvKNy25HCz31mm5tqa9ZW5
xeNjsABulKPUxLrt0NTE8MLHb+FfOk/Xr34QSUYR/jH2c9YjrlISIFEBLEH/kLSUhRUEg4Nph8MQ
vaU0iQZR+UF+a9v1jkjG/cUsHWUB56OQZVdxfM6bq9fI489SaHj9Pldug4eHYC75J8O9SZK+FkSB
ZlITLCmC2PFe7t0G8f7tjSNLs/p3IZWpXLN1qklRQpF5AAi4L0QNeb47diHddR9latA1n6ky6an9
Pp0W0aJuJuM7iwiL3bVqTJGGV4LI/1yyFmJbrcnsWgEjiXko5Ajho5GhTQLeWKXmDC315Dw1Rlpe
MpKWy8bw65YBw3yyZ5uP3DKeVzdnbwGLPjE4j31F5/rQu8TjHfPDWfn3SyeUKbVWLgyj873aD3j6
mJ77Wl54fDIXl7QqLYs0Xm1QY0ObMWY4DLe+h8e1r1yLZ2XIOMkST2lFLTtZhohBtLc8exKeILp0
1UsMPi1R9L61zMjbH9mSMGj91CJE4Dp4Fzw109XvHmx36ha+rlKbjEM2g0fkgGaq82GFSwa80uip
22GC/BQiKFgier4CAtfOrvOpkIwhobJJtXbvIgzmxHffQ7Xm1evmLqMRQehvrLRLIFMU6ry/hUQK
LdnqKowyvHY01KzpfhQvlP8lG+FwOl1C6GgLfAPLoWqKnqEeut04Km50vUjAuhn7rxdsKIUGc4Yd
qeL5kWK7kQWU0tqcrd7dT01vwUcKrWoj7Ezac58kcEosbnplYYwhlFjrDWm/5sWT+B9ymnaLfdOU
wYjJgZAytVVZ24WSmvSvv2m4ol2fN9EA/l212IZcuXrFTZ9yVteahkJ+SAKXz7ly+Ta/lSucwQsh
dWxl+DZTZhQG/HcuHXIn8jHRi3a8mOXbh0nvECQj81Gapw89v8wUfDedL/kMy0a8L/EA/CDR2Fth
7uSXVSlQtHDck/m2+eQjaeTzOYCGO3aY4FP4fswN6f2mIySRuMqPxaYYbrk6H28Uzfz2Rem92ahK
oUz+HKEUl/gka4t5Ej4ubLk/GbmOQnwxgQ1IQ8kWGdfe7/cmUNIiBgS5ojp7Ri6brrUvo6SoYYwN
jHb8IRKvJrzffqj2+5ZTjT9/H02AtpQkaPxedM08vekkdwIv7eo/97mDYp4Vy6aUKMdvv50MvSIe
hoojWxWnPGfilYgfKFomuhByKEYF2A3yZgJCmt8w4qf1K9Qm1KBNJL/F8fFmV9Wd9yrS/5JeGEpk
TXkCu31pPQoCAR64vw5xjgimeCjN5Gu7AOjWC2BDwAE2rY2wff9uGK3eUeX/DzhbIirLOe8yrmf0
YArJjLmiPKH48ciItg4jUY50Zk7L5P6cdOHtkZG21vjZgVdEh2gBWp5XjLFIFy+t9/btqnZvMeV9
6iIze7klGcvbW1C/4CwyQ8FTROLT91cR/0iLGsfKU8rvHFs3pA8eKtafOg3jdbZCrnuQ/Zgag1dE
qBtXGlhgEzbKX6U1KvJ11kdTAHKvUCCPWLVI5+LVVlmHjQ3ks6daeiQf6mNI5LavNtts+wRttN0h
ouODsv2031ND5Cy8gxV/0lmsOxVUW/SgflvTZqxowq6U3htuRUQYolnUZDVauw2epZO+KjiVjvZl
jFvOO+Xlxa/bCOtRT4nTu2Ht5/00d+oyVmGadWCYwfzt9CHgRGOkqF8Xe9eXTcx1q42k5XtfVCZ9
xAQ/6f/opLG5JVh7MluH4NKRhDmnOHoazc25XM0t5YolGb73UZSZ+WTQ9toH6ekbaajzCW8yXSgl
hebw131o0Bo9Zvgvnl7blHYS3xc/TubttODQnidJFsfcQMJbdUpeScoJt4FAkLqCTPSxLPxSUx1J
L+QvBuVrK/DVYuja538v/9RnTKK3WKLKm5UgZ25exQPQh59AfldDl8K6C/KbrHr1IYKJG9oTJGz+
ykZeCu2dnQcEDOs3zXxzwBoQGikWR2XMdpVC8AFfg8LndNFJkEFo9kqa+YJOZhR8ioYCex5VwVzn
RnDoPcDhpbgto2yyqh9jUiIV/cRc8dCpe2tmtlOgxhssadVlBbwQxqzQgB94vfLHBAxpS9fajR6x
zbbD5WfKFZB8GiPFqAi8tSKuWk15QUpEm5isdmUcGAgfBcS2SXUy1HHnycY2tUBM4qMthp72s47T
v0F4yWwEXWFGxR3INaiGjCFBaq9nKeWsXM8uvCnNTLk4VavDxNnLeiHpgPuXf5cIbebS/NDIK+tb
gC9ZMuchRQgOZq2NDpDbULVvroofGQ0qOTdMJ9Ig0sMNEd6ueRZAA+fxvgresUeLtB4qMEvn1uQy
N9+EhlowV5I5MoWFxGvFERuGogrur8wWhz7wFMyPKBJOZXRsVxs/yQ5BJvGEepAU+vw7dZMWFo04
4r9e+K2PVfCC9ffrn92P28MFH0SuER4B/pa3HS3ByYDlx2cVFS65oDnmNDWWm4aM4z5ulWmnLinr
l3nTEzyCVjWIjSZofSQDdNzjRFubbMVgOzLi5XG4egIO/tEiqq1nyNNFlp3M0smq+o4GNIf5kwO0
l40OSnwS7rhCzafSdu9/LWq9riMciKl6/1yp8Lvf3X2WN1rUay4X54p7HhnD+sPwobVBWPersyfK
RBKXQjCoU/WOufoOAB90Os5jXUjz4V+SRCuoXSnhWMmYBQtAQZxNIzfyI9WfjNxTbQs6BYzglawf
KP5wSNJo/Pyw0BKMrrbwTTvrEPcq6jp0x4pld/L1X69qHe1AGCrk8nLKGzGsqfrzQ1RpNNrRZKBS
q8akbRS3ud2Kod5qBMAiZ3iyr3Hd52j0FzoEbGRiRpmF1vqnxlABaSN5liJfael56Ck/8EIiF/Ox
e5o+9i1FaKJqi19dnianZs2TmJy62owJ+c8jJcmK4mxqyZv8Fji1iPPkPPVhZhgd6KE/X4Xa/ZVh
U+b3n1tfgxHR/ZzY4hl0eQOJsjJ075m+xYFib+VibS/yx83nO/7IOEXwba3JJO2yB/7t1R/yI3sF
NM6216HRqLSO95kB5qHedqu5oX2TeYnLafkG6XTP1q9kYk89lZrwh5ajUhwxUq3eQ5Hgb6qJhpuq
ou067YQ+t2CpCJv+wjK5W17uTXopccmEvayxsYO8W0Ky/R4h+Fn840ZxHa2yX1b4I42yJNRV+gUB
Ay2aew0Vs5tdOmSSjpm8KdnU0EGlaD4xL3B5TepHiVO48EwHVWEveiowLYp9JniE1qkFKy09LPed
wHzEoPUPyneEmBgo5dSCnrwjtoGNuIvyr6fyywmc6w2hCgWnKMEBO7q/T30aWmY5SNI8YQ+Kljj8
9qZCeUAyeZBoT97T85gLAY+nD9Svl92P7YKkWb4/m8MntlstcUOrt+JyBJ6BOHOObiSuOL0qw/wH
O+F+HFZn78xDelH1l6XC1CzYEkApFMUo52YJV8rmel0UHKBC/YUXQr9tR/qpAmWqK1IG/E5yog4Y
BHGJ0ZrIpJUjfb2A82jZrH1cCrpukaoy8DKfdhBLExhjyCEWvpcbsxbAweJ6K5prycz224opS+CV
YPiL43yLgE63q9yp9TT5v5E55ERykg7Wj/UbCv6sFw9LgsneheviN7rFz76rlCUCZUhunv77DArc
hzndbJ4QyYk7dhYWIyY4tORjgHmGeeEQLyhoqpdUUAuY/+Lwz7kuSlzc6PVQlr0fceSsHKP1b9ga
M/3BYg3+xghIuwWmztOl6fuJdyWQvbEf/GRgo3UjAfkz73YhrLB5RtWXN+t1VaePBo8l+9gOnR0Y
3D9CUz43ZLztIMYcQ+itHaWob4Ccb45OJ+jhMOmQN1bFdKgwyBXcX398dBvSS72YA+spNe7/tbpy
GjfcPsHbK71kH6Lv8tOntFx8660R+BtWpDteWpxz67NFfdUuO8XYjT17jNmzgSEhDFggJcijzUJP
4LyVOf88feA6wE5wGITW42reb57uQNmgdjg2A/Cn87mS1YeEwpx/n9kiJdeZiVwEHdWFTEKFbmic
5r/tP2HxJ7nU57Ph/k9QELcDgT3TZlidZbnhCmXsmoG9ZQVr+0qwxWda/cjQJ/PYeJM4WAtTYD66
mha7TTXDhf/pOzuiRlSHGn6WKY8yKt/bZOXTZySi3IrMK+3b82naV3fj3IY2ib08DmOvk+0CpaaK
qsXYhPhgJBg6bV3+IrrpMUzVu7VnEV4fVmbFja1/DGFfich9r/Zjlh3lgDTS2fWvL6spZYeBgyqx
IDBTfiZ5fB5IwhineHWmMVPUioB0Ixai8K1uUOfOpTtb1H4aewoGfyNlhsM4zPvFrrfQMH+9CiiJ
71Dua5BRkSAP32mtEFmFnkC3hQOanTcR9QuLhV/PqZ4GT3q7Ya/cJkwAK3R2+Gsw0IkVcVUJw1NR
2R4v02fLhpNY0+FomWoL6O96+xi9Z9IuXBiNjx0LdFfsbUxLW9js51aRBke+vnfOVgCf0fk3NBLH
k3S18SIZh6eVoRFqTt4O5rhAp+uF5KcYFUQXBnc0JkI00PdzveCZbxLTiYydTyacXffFv5De5Jsj
dEDasYxtbdSnePIY/rDuIXYce2T0OQjKxQ7dEJJMNq6Vg8Px56LjWNAjyiiP/TbssALcXQLWOjYj
92Boe0o1GaLV3jTB+Bg/tdnz9G0BNPseiKcbMkVQqNM6NVv4jfME4EYbiFnlJTe4566ZboPE8zJ/
7fGDNVG/McJsOyo10mIqn+H7HjFWLDGoE4RC0TD1wIQ72ZsbS1VF/pg/lks2d/dcAtoZWUwqYwcw
hf88blHC2BaigmB/8DwCX/IKNs8hfHNN8PgZjCIx/7s/G0EbQdjTURg5iLRY6mYDmtuDgrrUkY4f
aTASQ1T7jVFcjsIK+UZ08nEiu4b6gCPOMlwI2qyf7o/0tYUCPjMuuwBbGj2orroi2znnvwFJcCJo
MmJ8hUjdxQQFVgt1jNsxQbSgcioAGs6Ke/fdUOstokfEg/3XV1A8p91vvDj3KxYHa1d/ghpM3O7R
zV57A7suk74g87TDvC8uJFPZzbhWyiIQDiNjsHLxAXVAodwutG/dkq0GTQ7YBQ05H1YVsMSZK45u
rrNbADAgY3vF0gXkxnuGqOjMZoOAg5+Gno78HL9w/lhJ39Yn1GHZLlYcoRh5SjLfoqwBzRRAGLGj
pqwjc0Y2shT+AA1NWqi7uvxcyP4Rl1F/u29kIPzvc7Qv9j6tU8K91EzFRtVUpG99vEdqJMI2Xo7x
BU0FLP1okZs6oZmxcEWyqe9N7UNhS74JMWI0AaPMba8O/SxWGK16bS51R2CTGGmVsuaIXRum2/QH
uaKloOAkwtn7iA7a0/s5HKmWazBbJtyXZzwKpDoTdRyUP9YA4EM+KpocsVdVbslIPoD7eTdwy/ZK
mRtGA7sPtNpZgnhYTtPNMSDpGKNFfoi4WX4wm8vbI6CDYnyEBUPACnUQLJe2Juq9L9IN8CbfTggA
H2upcHHcvsTkoX1ru5P25bbotsAl/KBn5f4lfkGO2aW5lYaPWqDnhx7jT+X5NFCg/nd4Aw/Oni9t
jm4tILTudt+5PoQCcLB+ScktBp28DCeTOkCVTvwmD+r+4A8W1afxEa12a+SbuLZyg/y/qjLVWYtY
HE79c7JsK4k+04Sq+HHm27wISs7LyS9LtRa5E8wFiFODo58MftsWMN+hqIW5NlQqhTa3GcoomZma
+GXitXbd6m+ALVWuBgABGUygaVFnVWdrQmLjgtAOW0Qy6P13jZFuqx54DljzVpFjZPdVYvopa2iI
ygAiLUx0cF74W01f5T3FOpJwv52uoJCkfdoG4Ze1mqNNIlfRC1aftj52SqsqQUC93Klul2b1eBGm
CEUluf1qDtL8lNw9ACpIabKGPAxT5Jk2TM+ecGSZ0nnyhXsUwB3OoVHBoinN5GqrX4Tmj5r0qR1x
XyrQb85DeFJ3Yp51C+ZPnFQv8MtKwG+CgUuPQUdSug+etFYRy/eamJaIjEsiHbX/OotCl0qJZa+3
+APjWUGOpTakl2Lw6xTnpf1fr3GJH8Fpc0i2S7aOQneXjqeKiXY3dMhqetbuBTat9OfrENZAKVDE
yOLsyGNPfOrQQRNgQeMxzIBrsEeqejfKKy5u8bQmdde3Cxr0oIKYCwB8Ov4FUREuz1IXI20hh2c2
vIg8eedxXBqxm/yOkmWSzs4RqAnjwPgUj8zgiRrSttoVByaanjUlBBV3KQ3SD60jdncBqjoTlAQ6
EzFdMzoImb/gCyyiIzkSHXrUOi6TPKZkNiJzVRngeWaQPpg+cAMxTisJTRfx6NEFtcaIOFDQ9ufz
RrYYdbl1JiVdKFQdg3ydDcN/sv8mnxu8bK2ho1YK42y52tOFMQgMynYLG0eTKatPRk8WQi6GH9v8
VgfJvVPY9i6Sjy2xE4lmfcztlC8e9iCvq13ODBWmMkL9lrBFySSEAn+llcaTsVvj2HpmpCNT2Stw
a0JriDtvGZ2xwVsQhigRTdtCEU+K9b8N3v4baVdT8XQ3gFy5ZW+UeT3eV0G7zA7zCf4Ztt++3nij
I2pSb2N5xx0WFH3EhZ+kYSjWa6twFwflEzY24CfGMh7s6pO8lnVd4PzdckjMFWfgKzgmpUS9kpT1
e2cL21gc+G4i089h3qxNuO8E87CUd7IBWX+vOgXURyhqMgneoGCe2X2mC1sDBBnUV3sHcl4eS+Bz
5FWjGcnDvXlX+skkK+mud8wPyYixw6ckR1/jKQvAAdpBAptjGT1oFtFgp677S4dzPe16FDwYlx7u
YaebKUg3yA+eXXgk8dSdnKJBm+wADHtTUqOtVMsVv5lff6ukfco1OkoF/2cxiOJmCGemA3SDLGrC
3ePUf2mZbk9Lp0knimmCgPs2jRUOyCpMtvS5yQqQCCS+Gfr++56WB91QtLOAZZrcUSiIgS7rjxF7
GDoR7jZI8L0MDKoZVcAhk5Raz5iNdeJFoVWk6gU2F5MAS3ydJ793BVGLDX9G3hTgrdOH4bMSF68z
SBO714k5Eb2GjnIxZcrHBB6ejYFGa9JwuBKkzX5Or/Hfuix0OV1MEZ0zhUreGvfGEM9UXNH2kN+p
fNuHrnKB47gQIS/9MYCZ6qzvLlFLQ70PUZEQQI23jUe9p6hibyuyTXTG54TsbO+h5xB7wFFxOHlO
giRuaBpmlC7I0VjI9jHGKoFG3QYutlajZqSVbTzRN/veqCjACJO1M9GY8FoCanAeXaiZF1Mtg6VR
sNR50LRLyFTtjtrCeLqNomnMzJfiaZA7iwIiZAmf6eu/QmVNM8Q0HP1sOcuC29u1i6gX+7q98INc
nsZsD78+5Vedkjsr3Tup6KcuXAWFHGpOMWmo1uWZYNisNmTX9cj5b3cSPIO60os4qlsi+OE4y386
uDj/xdYmbVHiVsVZgAftn6GYuVlcQyvDy979c+bQwUDkdM59nIc0YQiD5UBLa1zP9zny4Zgz1ITQ
SlyOJ/ntPzkyccjqdWApVB3lyuUpfolA/PriTAR/APEz+0qwvQHcCEFntJ7TsnzW80cvuXclp+Dl
XHo359qWcQBSbWlxOpWRZy12S5HuNrXfO2WMp7Jm5fcHh274I8QL5I5Z2YV72htigAEYc5KG+vKu
/2F0/+6nqj43hunXHQIb8o05C6roQUq295w4PqWIvO66w8yw/ZNX50aQfQ1JcwDQQP8rvr18T5yG
twgdpC5VIi82qHdvKmULYqtvhJXfkHzxbYYgw2wjL9D1TzXbWCKBWQJqnUC22t+zaB57sVgdvXX/
NyXNd9m0ztS38QrjN6DTIUdQxgriB3M+ZQPKKO01zUqegUqkbZnGDZdKQy/i4iAO5NnJRsxsIO5D
t7V+wEB+mazQrE+a98VFMoFzuROWrLZxjoRsh5+U8Vi/8E+Cb+D0wA/jeQAci+fbX+L4WBYdpYTx
fLiFYBtaV3szjIeDY8jR3LXjNb9bo/fCj5WgaxEepl9800Okv7aiDHX6sSF+ZRwRgDA8VO5T+Bmj
0apIyq4MHeyHQ7ZAMyBA3/6m8LQx4BcoON3ZLI0KvSSeKBlVzUKecNIihTlvQ5vNjUHwrI8G5WfU
sMLowBKs0CbgyDDWw+7q7+fIlJEgZLkkvja0T0/6zIWsczjZPi4nOeHLdQ/x88k1k3MZaqmCFh3z
ve/9dBPvLzXeSsdaSv1mF2BGy1Xp1dfMsuXGNkRQtaPwfDWpkiZpzW+xpzjfEFw0VJzm+6nLZWT0
o46JCabM8BSQNpbL92j8KsIPX+3ShnjmFJh35SjFne9jjzz94rPQgmCYLfglB4RutHQd19FEHR54
0e6sloJ/pSN5vcuDJH9aoNR1yEnB7RjUwD9B5gr4McGoTkYUC7NmLgEid7FaofGDpjhF6K9wYGBh
6Ql5k21V5Mw6w5c7u885TqPgk6sa7TlmtG9/9mSUpxPp/dL7oaFfylfoLr1rz7gkuUchKjXOvpMm
wdZ/2kJdcH4Ovj8+1L4OmtGw1/PS85DvWi6pm95zLmKVkKJc75uiRL4vGBf1xxNV8i+DSUaZd+Hn
yTW7/k3z68aO4ybydS3irEDDJE9hvlLWZtPR8/0aEMk6rkFgXYe7rEtpNezS8pnOgV34LACZd3g/
TayRUrTfOy4BU4Fh46/uGtIYSIv3h8+ZWYcLAila1uS47jQwPSrrJEiUfv7HvwtJg8R8Z7e6X4yX
amPgj2tsN+RK6rNARepbSjqFdCdV/KypAVb94udTS/IVKpHKwbT/iIV+jBWLJocS06LqYUAdA890
2I6U1z5Sy/QbX7/MOe6sO9uLAk52sRDLu/pwJMFFQ8XxXN05gFn0qOoYm/+Pmbk/nYjoKAYeBgqN
tIyd5Q/w7Euk6HNoygxFHxWfUgyp/UfiQej+0QlUvmkvUDHcMyVZgihojbDiGFRjswqMEphUyv/H
1ZNzpjmQomUB/ni6itQ/Fzih+8lhC/WHJSWVgE7R6fUFm7w+H/En5FizhL/Qr8zJ6WG5itpqEzB2
kEyEOegdITdX5TSY3ihMEjUbUOLfEb+noj8Wb/qoyFtTkp5uPFfn4aT+HvgB2WfnDeQjINsg1LRp
norRe/U5+QzHf4HJAw5pgR+oiK5qYpuP1flpnA+woHWVfu26OvF5nlRB0guYzRjGA7SeUZJK/qxB
MKPEtVxnbZn2WvdK9dkUuGRrGghOf1VXKKQgTW33bC5bhusQMn2LaZw5Pr236SclRpsD6SM9vZS4
gPfNjel0KnRVLQzTiJnsSxrjNMIjCiaqkkkng2F2yP1dOXF8uU7hYXUD5+HSt4Q6x1Mz/2iePhvZ
zjtHOW+pXYRrZlSePKRUoPBB0Rm3ZrvNntxJSKhA6/2jflllpPsQMEsWrEXW/FxJBnqINHZmCbWY
S1uiI53hK9iunw89AI3PKqOY5VLsaDbKHlBhTgcrwEgG7eQOZ+EW0Akz4GaCDSdngNJymRfWESD2
nXyJbTVGl3m8hfq2A9Kifd1XMgPFeq649aAg9L2V6hLXP8fwg8e5BNCko7K5FyTcDkQQHgyKUf8i
TueC+UlupT8xcsofB2zzs8BX87ixprNseQs8RN037Dn74Ow1gLcXNWmRRCSXRDOalkPv7cy7eeLT
7cGb4mb3Mqg52wQeYNCKeLLyANrGXv/cwTCOGCx6kMShxbOlHBQZD0j8kTIIZq7GUHkOu+bFEu0g
N/MzkOdnD8lIDiV0SEOOYKlMxFfs1h7VntWVRcN+KROreBAhUx+Uo3k58XyMIHMnmSO9hTnmbVFK
OMEoCHcpV9jOhPKEuxSKQLNj3KWiV2VsaipqG1lM0ahnXFf8iSerV+stL31d5qlNJv2r2FvEmgsq
XSwgiUh/a+Zg0aLjyTFqpGxvP2lybgXYR7mJY2YcmZQ/reG+P3siPIoWxjy48HgnDyOkn8AW5yHc
RSIvW79J6mSAwP7pMIyEMMOuqGkZa63tiCyxOyyRYUHHK+2gyA8V6uy1y/mUv4K2uwtxA1aqFOjm
Ng+yY2AqNMmj+/Yjs0m2U69GTZtPgW3wgs2OzwOlRWDF81bx9j4MjVZgQJTOSK9B1/+xPnTAcHD/
2vYkca/EDMUwXOx+eGTrMzbx7HX7CnWPerMABLu5yvdYADxtXEBb56eubsASqB9RXJSXJmniOpcs
JHLO+12PrV1TXq6ArScuxUyH8f5OeCjM6AUUXdBg9u0SShkcr62SawxDdPGxkkDcR/17lMdSn7/c
b8XsxduokzNz6n2Mxw8vTHBK0Vgo6i2ZnZ5NBgPGicBSSzGiLMb0nVtSAF74oRNQUtJ/OzEAiwXs
YhNnMEttP98wrBTWeseOP5ISf14xGHzDiuoduI9ZbcS2iJDVtJn82ldGbWUPFUCLIfFdIlD239Ia
Mm63Kdyf+wNZmXHvap+bosC9+WNKxLsE9HZ8fT66fQ6ToIPWt4c7M7AZzOSqVf7RdPlTsZMw4sEX
GX79JlQmkPPHHfJz9Zk8h0MUgChYVHzmRZGDC+zjyQX/w1SdO1QZKIDAiQlTK2gIbfLXrIUl1OEL
9fyyRdevAlhm5cL/4qcZYk4qLwo7iq3v5nK3Lc+VrHm2GX+cNjJwADZI3L4rXVd5TV0s4y+zZpRv
ePzjqqrj/8hrXyMezrVdBDnKsFe0riUzR1PkHn/M0Af/c3n0qBzC+67PHxTQb9tpe1cROfuEdvwF
32d1Mxp+RTqZOswVeJpeKGRZ+/1XLd8I3nUqKfvfOmvA8Q4IhBlzEsxDzWyb1drMrppfYpcSuNIG
SW0GxatTxrvUWfpXDMOMG1QenIbRTFGQKIRagPT1VwDFMvCL37O7NE7AtePgUd32ZV83WcLKLOw1
uegIu7YKgZ+JXQNR5WX7cqoqKtYXdyBop75fvL7zqfD2TPflPx3CUfyj1YNhfbWJ8OivINfTu2ih
Wa/qFiBoYqLcNzcKPh9Jm/aypnotUfLGsC2QuQkE1PMSNM6SSNgmpgv7iEhof3uX3+UV4tdiVqRB
4oeZMKmepZ6xBY8XE/9XDcqgd179T39zL/ucwz1jVD82zqQ9jAfOcQFhIw6KnvTFozWXpVLPcFyD
o/kZnyABVgEFM6wr9VjVP7yLMb834EUi59xP35xOHvSxJir30oQd0amGasjtrcivRm3C6hsJtIOe
98p3n5nN5JuqI30EylGzHqcmmrMetNhdQYjcPBayGM5rDrOnOYE2M67mMgouYewgydzU03G5eZav
+J1nzFmjWeIcHj+qTHNhV/5fvAAWJpXjaxQVkTblfy7BGc6ZLZIo69NF5kVcIAI8R/D+RGUfP2tx
W0Bn8jJUmTY3N7xUrj/LG8ve0lT1DYSsFzaMxB6+MjP7C4bT/T/NFm4mU/atMN8fcB8b+RLt7Ka4
htOilJPXploUn2Z8M772HWe10CAfrp3f8k0xJ01me64ZqCbbC0Sfci9no47LO5bsecmbmIk+7rDv
1kvMu+zeZsKTuy9UOlSTSosZXdEm4BHyRBsGJaklQ3kWT0+/2FEcfylgtFimx+ITuwqy+shXLMQO
R4EkLbs1KxzI9ZJiddHLfG4r2/kCJct4uIVQPy2Xg6MJP3B8pcGieTxZOuW6xCDN2YPpDqnpj+HU
SYCqEnQ7N91wJwoAKw9pGPN32a5K9cg+RmWz6Vg+Zmrzaarlh4xmizRgmZ25r8LpOZmL+SsVZ9Ii
gVYfYkPtZe6KOjh8Frpd1o3RyL9PEC9AUOsvaPARW/IYwLID/kTpv50Vo/v0ONFwxL94Bq7eJ9Gx
KQ4hLuNLGoBEUW80Q62IH9KPSI2l/ptWwu4kvmyWyW61xQ4ugjPNWrltNMFsL91afbkCaRsqKs49
HyJbsT9ZTD1n7/eROOqwdMozc3xx+3DHOAGiu5pPL5u75WZJXi9XBNrzFPQNWBHFRfNaCCPdOnoi
1p9Yvv1v+5Ja8VH8DK3s8tks71RjRQ2A/JZtg/4LTGd3hvz7LD/XEQVLPxPtx5LcEoN8yqAce7nQ
Uw2GSgwwLdTsHupDK4ZoPY2fI+STPRhnsDZ512CbE3+pHVXilnlq7EInqtTpaAnLZNHm/uJSlv3v
P5SpTwci6DUjYuxmbbmwRL6e/YSOGdB9gXnRPfLm7weoi8+ScPR2wVWgKbF9Itd2ZktOQP4mQU/J
ge97ssgvlTZcEZPpmxThb579/lgaAqq5iJVP1dOBNrlaRsmxl0uTWLftghe1BoOk3L7N0nCNygqa
OIrLYv5tbxBGPpJzpzWQslGXCT/mDKmddSuTBrMynI5jUj5WOwdxrJE/drf5oZHnhJKbfIWCCuLV
ITmobO7EWlwMHZ19WltIMjBFNOVSkcf2Gat4uZzooYfTObKbIjQyyqH8ryN2s3pKMDAqcz8bWxy+
Mb1bxJDH/MJFfnkk7582f+/8MXbq6QMDbhbMcg29J7XcUyPKBsYYC4Z8yOVdxwPqXb6BG5YuXnfA
wc5ScB7eIabtvNYMLsIhfyZdkX613zjwu1oNLeZjmmw8seM9cn5LOEE2jlPtrGKj509d7ixsgKK7
CXRqubteMon7Mv4tbvbO4ID8p3GyoM/Lot3yVuYUuPLIbZehRcorFJoZahWbdF5BneguyVYWGsJJ
GIlcDSvi6Q6jU4DfQGhgl9mSpJsJEAaT9rIcHyGt1KluDgrh0tO33IDS+Z9lo8YXOEGUvUWtvg7d
geuBMLi6YIurkfIBBRBdx0TJk28qkuOSJuC4Y+9NyqeuyKLvv2Sa+SDX7k9gAGzuhvxbNjrlBZIB
da1hcGKJAcfVPrT8/EONn7i5H4TS2JFVqLXJDYHMVEukPZhvJzGNrU9rZJTyGbODNih3XkCsMvvO
08N54DiWqvYVMYxeqLxK8Os2LRjsftaLaLfCDqbsCWAv/5K/juiYplolJ75vEqO3NRfVx+rRJEwx
TLBRRPq2takXDP1OxGKzz+XDgzOAe8fYqmv+xuQiBqEv6wOyeUa0yzkktX6CCCbvJQWOZcDBoEC2
sE2Fxqk1UPyLYZ7AX4Yfk+LsPW/0oQ5/Gpvq3qd6xvCvA6PYsojAcJw/Jzpr8TfRM97N+P0RhYzR
K8wgQKhI+7QlHBJ2fFv59Y70GLVS724FDzukiF/zmLCtmOGnbidpfHEOEEkeBd3JRX1qVxvDh7er
pFeAJANpsvjZi9+bB4kCvZ6eO/z6zQTG+RCjtGj+igCituYzPfXngs/OZ2gMoJjD5tmISU6mtk80
JK5aUmY2djSA1pMNPYx8Ou/PC/skwkd+scvtfkqN4bR1z/ZF7VN52ZD9+1u6ykkz3ynq/neKEU5m
dxA1BifivUWSNPVJurJRidRRw0zXRg51X/sdItaC9hhaOk3LLV9MW5qkmNWttpTYVeOCz388Q/dl
URaF7zcB08/NS5LMhiPEwuJy4udTq2zrWentl55x4yfhXvOg1S8KUuLOs/moW43KpUEUSIR4YCId
IaZaUlxanDpmXWOUeCo/i2UluOZkzQXztm+E5o5S6ZQADnDQ+x/CNx4FgfOrZk/rEuQg9MVkCzCs
lHvEEyQpj46zbmt3lNrha5OsQNeFRNv6DmezOprv15KB8awk2Jw3r8wRvU3PO1hvhhHjFjgigShw
7Uy+Iu9+Ly3V/qwiMRLh0U6fUkOnX8OE7zs/j3kcMRlMqv31bc5z0Ii0e3RBad/ZALoOOf762LPh
sNRdazoRWVhx7nXw42JQJm5sXaJTiTOwmz3iQjuRkxUO/Pt6eYySRYGvPkHTbOflJVvOoWVKepcs
HNzRHMW3gbLbdAY8XtEvprOcElNopqgWHXJWAqWVB83G9URJnsOBccLRmQnuTISR1+Ry7gMamlvk
7Oc/x5G9BxJxB95trhmq5b2g9q40mF3XnAcqMw0VDlsCTjlEQmmDlyv1C4q39clzEVrkLOO6qwNC
go9Nw5PUJMjYYdNONPADe2SM5UTWHIPRALU6bwqKWKz4SlLRfhctWjv+G/R9Nmshz3yEOtAZv/0N
6DomD+ewNkszKcwtl3JaBxMrU6naQ9ImdcLG18bNO1ln7OXNg4jFcBXQCNdCFIKIBl+hpQMUmFsV
r6AvutkQwJG4txluTsT+gU0sgvN69fFcG7p4MDZ8P3y8rioasVzU2lp6rM3i0gf1ZceI2s2r6Eui
Z4bHXiPpBnYETy2f0B2fhLV+tBZVUb7QbU5kgoQA9SZPj4WbdYZjE860KIC5GSLnMG9uYYoPzF1J
PVv/mb4KTRyDbSt+YAoe12qA8pb0qptgcPQ8ypW2kS/l7c9u4hlX8sUeyCMmOIQwx0TAHhHNXhXJ
rb+m2cVPmy9KfNEZ2UBoMmCI/0trzygxSUbQ+AWA87NNi3G0l2ASZpIgDvMthEi0pgcS+U9MVbou
9/cghW8K3yg03H5wXxWVWQRd78ivvPe5LVwJK/u84z7+jvErG07bKv3PUMsrXutPl+nUc632Ihyh
JkxNYcX4125MQ0RVfgsGxnixu9fbLQhkCaA28qtTlUAm43zq2FzfEUom9QcVPidG4Iht5xRkVdcY
Fp4leUmSU96ALzfymwFdR3vtxJMdpNKc5tmswRtowDJqUcCJeXE7ElMHcCHU+v74O5n/urO75tE7
ubm3Ixekt3j+hFaaylB1tq1NR7EG5LiC+5oz1sFp2LFD5uQ34qk3ifIl1hrE3Ayu1/Xeo/YQXSIo
SHDbuelKs6WFzsMiyixxs4BnT20SHG4pezDVw8LFtjiTws6m+K6BpgEhPFK9M1cw46TOCuptItrS
KR3H/Lmqf9VjTE4Z9cycVY5jjq9D0QZRGZgsy/TzBrtsvmT03H9jYWvFmokUlTvn3TuJ4ECQp9dX
lEfEUigDxp2/lz27cH63TPDkq33LmTTyWxYvvfRJVl43RYoTR5QLfGmDi1h8ZLJs7TBEe1gr+U4b
aaTqby1sLocREgKUBqvSQIpgYh/wWW7Vh1nulthdFY2y4DiENx6kdL4CAjz6py503xbGAIpDoKWb
M7vXQT/Mpf3nLgvnhgIw5DkV4H210o9Toxo4VTjQj+cpl/6wZhH2yow6haMfEsfnFdOEXTeET01s
UMgMyN7/wv6xf9NWhyoP8UVjNFrkJMczu5ckEpIUV0GHhI6T02y1OnxxvkXARRhmDwimdHXeUOfZ
6CPyQFt0dPIqogt8fGWsZ4Huvstwz31H0YJ5k8Fmuu9jI9c53+AeqR4dEpfLPai+O/tvSKNXfSF2
NzBFc8ywSDH/iDipL9Sj2UdxRUwzhd+eXBA8Haivsr9UzKZiXKYbbOoDiKIkNOHPy4CdctzUvey3
jgKBbsnKteZrOy+NMd/KdoJrfR+Ws2LAAXl4xfm04r/gjWbnSzGDHOZf+QYaVeoJYI0NA7flAyE3
5prClPi1Z5LwVccSLs0WluOkTwNK4SatlKjcwazd9x9O7VQ3mwIB371dqlo1wgNA4aJz68qa/4Vt
8msUnr309Ja/ZkVYs8KsKyDa8HXTznzA4gp/RafcDNQX2Sli0dpsToFREETQUp7OsG2tPRcyJvXu
Vgync6RnyMpNcI8Hp9u1nHI3RmBdkUGrjY74Fj3x2Tch1yYjU19gydNPSTKXNSyclXfZbhUxUXx0
H9H4VEVZQX/Bf9eDu3LGPrRnBdVHGCTkeGLKqIcP24fVjzoRFprlwZA7hYJj9KO/QhIRsZbCgu1U
kVLSBDHa/v8QLNF23zSXGs70NmYwsHpIz2g/1MwuglnpWZMnhpLSDZH/FgDIIGJEDGaRH3syYD58
tIIWa6yyZGxyLul212SlwvaZQBsy+eJtxAdJRxm24NwWtGr5unHFftkHRWRFqXjXHiwFsyStDZig
+dWCNLdzu8UTfh2x5+kEV85IUE3q1R2011rzc0rqpMBn+tM4F8PzPrmDWmqTTI9EnbN0y+1zZ8pp
qYdSiOx8lIk81KBys9wECIaQioABDv2+Y8E7IAjRgCxQ1joHyzJJWWuAbUQIlaPi/i3RlEyEk7mA
CYl9uV7M6q6C9VYHqhrw4JcgAcn9pQM91YSUSWO7pnfo6obg9Lf54r2P2vOd5taLi5uZnITJjBGR
GEi6js4Eo3FsT+/MWP841UHsr1GVijh5Bmag2MKrQmN3MvS28QGterY68CxOGMohvnIc11F4fyXw
qLPbV9Qm/4mA8DBDveTWHXHJ+6/X/xeDnJKxZzoYN56fbheXeMRo+tNq/rQNHl3yv6TSYSRV87ju
jB7IHsdjeQDvexlq1/DdLrUV6bA0RSFnyPP+giTOpqMb/+YZgLdN5OaouoGCM73bJiyyKM+tDEkV
EfXwg2jNzJDHlzGzPmvysEAYrJz/3b9CPTNShcCJtJcpsEfDcV8MFSSw7PalaBNOHgbSKOMvuZSc
AkW8FIO+oziNU7DL1he2NA/c/AVkZ7ho1+NbKJ6yJ1mQBf3PJoSBaJ8OS2OevU7WGGYOqdgdJgJX
oO0H5OGiNHb3PRfzQ1tzCEwxSp5W/JLK0cZ923Iu2z5ETsyap5oddM4Sy2Go8QIfYFCD2IDjkoec
DYDDznQpeF7k34mD0/UoWx+xMgJyuTj9LZ6wFHDXoy+iqeEMzvX0uWH3fpIqfYhVCu0av2BRgcFK
4HZYMpxfdDezXqEYx+0KSXVSALFX1IfSNzqwsqxBPNulQg4nXTmF5NgU3vrxAhIw7nE2gsCl/0O0
elfceYQDK1GgXARSgS4JxJ2cE0akxjE5eBH6lyqxApEpDnkajibQU5Oz6C3j6Re/jVscjZEZBwKo
NFcT2JArbbqoqY9syVGn7BJotnQX4xR4FgznJ+hF2ISYA2n6x4wuldmrwDi7bnOLgGFE07A+41Lk
Ym4bqT8ZzhqSoTWuLktr+Mt0u/jlgpXqGdu1zUFzy3RMDY4SoQS/jlOgoMv4LzZnfZArKpoKVMy8
w90H5J6UZWzEu0AhmSXapslXLlufSBkbaRyoCxt0UnxSp2D86Fvb1xqIp4HIXsWIU3VQ9iJp8YaQ
xVs2HxigaQFuIjTyYnBny4b02btrSLv2MaxYn/thPhBWIWvH7nPKvqEg9BTcbCASXmsqYXl/pOne
ZW90+74+lQ98e/xqvCkZeqoGVdq9fyRUrX0B+EgO/JU61nPscMj9JyERjLE28rQcg+dkGWEbF6Uz
lD3vJlaK6wVe2Px+pTzqUkGMbtIkWEu89flvNvVCyxmsnNYu+S2bkhcWgMCZF91+aYOVBK/FFSxZ
RTCZ/8ZjrPOqJnOlYbI/yPc5XHReq3bWJmgVxzSbR0Sfk01YbdaEND4HDMLKONBGHvQjA/z8Uvtr
xq6DxTzCivak3wGB+7B1sLPWCCLp3RJcvKpdjVJSTlsJfVtizgKVYm7acy5VdF0d5jZ6fB2mi6VG
VZHTghWi13UjPRUhFvBIew3VKUMm9Id7CJW8eB6aTjIAGKZPHkOb3IBP0m4ftFF4pzScq2qnf5U/
V9PQ2r6Ia+8qmgtfLP6qADcitpWVZKC58t/QYkMfRhIsyvTNGjvnhzXXqBXC44X+qBMfH+TYrQQ7
0pokCK1GQc23xbpS7kAltKsJTU1uFGoZIYIdh5xjbQthkxEyyOJfxfdpuaVt6tvNtLR7SRToVdv8
f/+7W8ZrKLu7QclQr9FCxSHv01C/gvgIa5kItem5kgaj6hW0id4AQwNIVpIWY/IN4uq4tncUtBh4
g2lyp9NnHPe+rUO/fMHEBJsCdgMsy3xaASYrBubpcHGJzpHjc/1/ptM0IdZDr5s4Wg+BiWFUOmMi
57/RjFGJeF8FLeYzW2pcHan636aNKvUckcYT9JVazY/6NUmLBXen9USGqXtInAaSG1NgOxLIHf40
YpA9d7RIzi65jQ6a+V7viFuwzNFCr1XgI0BCNKnEjO16VfJNir+v0KxcOwRagORpCBn2/Y01A1lB
/q1KmMkC/oMh7puq5q3rZUb/CRezWyPME7n5yN6JfsywQRiDqqVr4QwQzw2FCq47fAQPJYKXTxtA
zD1MeonltOTODWAGPg6lYYO1IBpYkQQf/7Aj4PsfdyB+WAhg1r8BP+Hq+Gpm9DF1lJPQORkzwJF0
yDp+aXSNan35my76GlbbKv2xJaETkrPDS73Hf68E/eaygXU/JhRhVuSLClY9y+KpRdiLd0PMDZwk
/paAIPFrKoH71eLGrNqPA8cBUm2EHzwJf72We6g0w0r10iwbYYPeJa5xxaHNjdu7hub89+nyI0rZ
eFnACbZn0lwQCd/hEBmZFBG+t9/sk5fdcpAKgrR9/cjnisu9iSA+GbMwNzLNkHErzvFceqRFa5cq
okahcD6VMS/JOnro8j/Z7PNAQk7mN9hZX46q0oPRNrgYcMh0DFj2vW2pcBnKUjIT8646m7Mzjtsy
+DTvymGq743cJFPjH4SDfGzlwIiPk7U/9sQdf/an2GHgioaC5Dv61z1Gv6AZS5FYmFgiYFqgk1hq
s0GrClGMT1np4Xx2A9Jvo7HPy8Fv+Hg+XlCvJHHWKvixMs5owT+HwjYSI9Rn1eLPGaOu3kyrtDUi
f6aPUcUIn1y2XwQaSd/Wxb18jgVJzEozDUdREsjh6FR73SWC4OpJChPqFsK5oCtvavRLN6LL2jTM
LbPD+rc9y9nZXNB4cv4lgBkZp4SGZA3efD9vY1NOwwDMkBr4c2+O6WzDPSBlWqIBRoUEKARPTys/
PUs21O2InUm0Q6Db+xCgHeDK8Hq2ns69xiLnoVFoSRpa4Bu2L5GYzcxIWtNIZBPH6YpbbuZUEPbg
onXhquaYyElp0LSeU1X2W8kOLHQDjl0WAN8VgLbTUDFKY+30BVAjuuomu3IyfBvgorzfDvfZtW40
A6LbfGYsiBHKYY0kCyd5wMLxv2zdGCrsUm9eYQrXl2iA7rsze1j3ruNqdT0I8ARXmUJS773qoCqH
UwHhpR08BWGfKx1we+FHEC4Fi3pozh9ykKyC1rQixlINuEOVqHb04kCtdy/u2V6R1qe6cZtxpS+4
rxZgWiTXY250m6M83FsmDlXBFRjRaLtvSYs5YVc0Xz+ecahVKijoI0Nk9nkYVVQckJm12nrZsr0V
5cjBGyv2q04Q9KSwyU9e4qRqAuIj/3c4M03ET1+/kBxi/r50aHxR7hI0r/LmkooY3ZTkcKTFQFw7
xXmrr2hugqGVKJ7LqflpozMdPXdj/Zw4Ucd9nQE5jUksD+kCrTUcPFg4a5BWuGdlKnde9qCQDIQy
55NiVPgDr5A2jfPc9j7+wYjiqbbeUqiXSE0m+F6H3mGmLbJ+BJtUQP3uVmUaiZWaE8qUYsf1Z1Ov
qHdOtbJk7AdxqVT6SJWgl1Qm+CCBRuhVgZ6uqWg8kdu/P8nTSPScyLurwl3KfNmR/ndpQvNZoLiy
AKQDY7ySXK1O2wcuQIjTkQnPZ6IJB0ahWZ33dHBEKi9C+Pdy0IDZCceocvGVOQxQj5pUX+iDlrEq
XKNX1PSp7djIEbcOTftY8eraZ6+sljrtg3G9TP+qvh/mwhZQ71vnc9o24j0ZvN4xtJ7pwoUchGpd
4IUMCmZ8mlIJNbRKnyFoqzcNaVNbGw2gGDhhu1PonigNV7Uy2MbDu4Wb1Iiaem2tbDje2n7Oz649
Wc3ZtP++pgbOvJDe7YouhFAVhexYIhwPlSCKccWPyYb8rP2wbk+LxR9wtHM2zDWJmDaAxFSdu5RL
q9PSoCaNRIzrHt+DT2TDBCrBJgeodLCPHZehrh/Qf4mqkCHeb+7AFCd7r9W8MgsVJQ0dmVOJDfXZ
j2kIVi0bVUm0OMw0D+0tmSkgugovVvWW0ZW+dpVaWE5y++p53ElPjBhjg38ICBSSfDjMtFyocQ6f
ooES6ufh+g4IXZGL1tCbprCE/ZA6fbNaX08PKXTKZoY4K/xzIQsgvWYSC3aUnWt3kyn5YeuPLyIL
z7pvl9y5289sSbz4kSBIDlUf4+jK1mA1FAMBrf/GNyF7TvSurCeaoFlfXfBMuuFvZHDKwR3NZmZ9
yPz5Q+oQ/GQelzjAonCjbIotjwoa7wa1cUTMxf4C8lBX/XmPKQRlo2y02PAhfwAgoMcYlaBrXgzA
EevR0xOo2u5l4HrZe+1REnt0pcI+DaDqjdNZVgsCTej5HyGvSj0hn3iLKEfN0tv5lWsCORP7SbF+
mOSdkURoaPXWCfNd45qh0R1ZLkW1o4LJNtdu0Zq7SiSH00r/JcheUgcqpaMv9R7eF2jkR/r+rvHj
AGFlRCF3dOOd8ZfU2GlrpGMrPd/F417y1Bm9m0sAbD+eJoZKrUw23h0r3TfzpmyrGrvIYWeWPIMh
wjISjgS5FEpsKLdQAvh+fdK1QcId5x3fUIKqC9Ssss8TXRLeoaWlT3OxKKHbVb/Px5LJ/JnE//6D
up+B7xpxwRcjl3bpQ4nk5VmW+dOz/ANKJHF0kbo9LePauiJRVBLemqqZOr7CKvqFFZyIJu+elwH2
Oxnn6aJoOnDdU942M+xLS03ddu7pF6FoHDNlEE3iI08GRlLW0NuBguE1oHJq5oxVQL1a5t6P3r7T
s7GGO1EmRv5rDfiOd1y55dmjWXogMntTW0Dv3IyMkSoq6yjSFuB8OsXz+ZUkdTzb9DfSHdTT+Oo1
mhwHeeUqDOMj6xeke7WwVcCHfMTYx6T5cfFcQ3EwpRtfhJXnNy6Wl6YrXqocoaKOWiWtcumjSueF
wS4weKhZosV7mSdfd3E4jjXLXsiMJ80LHU6dvdwbiopNQ3Z8nGt490/1wkveaZnN6t6XyWRzcadW
En6neMf4lzKxP+bmeSUpRK38tVJCpkaAoAhK69AH8ckfQ5pa4+EDPtFbdTBarzDuV89BZV2C2vVQ
Xxm/S2n509W0sXxE7eLfEQ79zZM0HQxhOtK+T6D3yeMtwMwPpcbDMhBsn4S4/qrAX7VG9kJQPvT1
uLmCDb2aw6Y7bsyT3T23KqV3YB0ePjEBTaDkUmqCr2yE1LSKPYs/Lk+onvGCHIw019HxlDo5xcHV
f9rORg9tQ25FX9w4wVgPAzd9V8Wg2Z20WKNqZFSFijtYzKKtKYTqutLQNQw771y0T20ucbWOn/8+
lzcKb8139sJ+LQ/7xLX70X1uNtqCKgYAjXn44XyLkJgsipSoP80X3Bh881aqaH0E69fLNDxk4dUv
BmJMfWOotu21Qa2svrkcl8ItKN0w/C+pl/C1U+Veu2vYfX31a/BaMggm7JVgdhIJL/04Kj9ToH6r
vSxizIUmtC4prDUcT3wWXd+lEr89HkPu3VF7QUqjV5trlTq3pEuAiZRTPo4ntcnq7ssXvoTfD5Fc
HNYDVfuYgKEDzTA3VANl+wRW7hPragKYGq1OCqb59T2uk52hjbnNfDXACS3ZDhnhIRPUi6BF8tS6
7L/6HpozAOw9NV8XCLhY5WJwlfNrlMSzAfrnYCbUnE+XHPTApW0EYJMFeO6jKpFYeSC3x09GB7VK
GRFX6aL12K8/nhj7WUYusGy+MTFJsPbIjEytmkbcNB9G2Kt/FG8o62qfKcq22Mk51sXfnSCzYbZe
1COX4sK15sRrgxRC1QAjXidg3Oq5UTuyxtEIxcUYd4oyXOt7/l/yyHGo0GXsBKBmmvXhoIM3ZRnk
4XE5zsyfjaQWSxY1cnuZRXMWHoXSMgrwwtRECCbrHTMYBL2dvmCa5tRMLUFjmngrVgRRv+zmM1qt
kErNYLWhG6NTik1Jr+sAf0xyzMnYzqxN2dD8dQsCqeQs6RYY0whxKIGKIm1POW+cCHygyJyQ2OTv
k8ZMJ+HBc3wKYBSaJpmsOSfXfXrUd6oG9uagGcMjVM/UcSzyl5BUCDpmOLNHGkCO7/LSzp3K/sJ8
qUaoagjfsWL49j0mmzUMMkIWwbUWIQuYHdtdqVBQ1PKMIwSNTyI3P3Izay+WHUhzoE3UFItJJZx7
7IrWrlQzR0v8e81d0X/+eTidYwqrNLDc9WZbYwXjpvEC3HR+zAoKVhhjL7EJtW3/3UoDN3hHxpwB
neSyeTM8fSYNUGyHskPPZV8ARgV/XQYEHDryl9+2SelJNrX6AtXrV7jHAbGuMWBjPlsSFAPbOgp2
ThGJMgxrn/s0fjXj+mVV9ISTLgvv40wOdypEeIb1hQXm0b77wM3zlNsrhIDlo5KxjTx2c9qQqAv9
mzE4cH5ayd5GmavBHrbHA7zcp9LIPqVLy/wf3dzmO8ZzYwXFMnp0pgz/fjlGSF6MSWhPwxkDW4ah
Q1h+gazMaNzQF/tPdUy+2iyIMpA0BZRVO+p+NKQUsVde3QGDGejXeyZ1wcV5C/k7T2xBc9YhDeVM
8jzL1mqs72wvV+0kOxowEwNNaoh5fWgWZu7Tx9p2HLJ2kmsGVkU079EGX13BAlhNfRvuxH8GkJxb
rUlr2vWYNrKrARZoRjrsspvCIsQuANycC4pFm7GdFRPQPwOuYv9jTOeKAGQ+Wb3G2+v6ibMpLBkk
edXKDMgwP6ExHNJEb3qWv3EfLVTSH1h1cJaChU7BK/bi5aq4PrVjaDV1XjZR3FtyLdOgmJiHIa5N
3ioswS74JnDEaDuV3EMIrqAQSaQYzviLzg2UwY7gx2I07ND3Nww3qumDSyYcuaTrnlaNI6HQKCNg
cZKFzZEK6etBRtmrjfCpAuQgPmzqs09joI050hngeolWvMVQ7eK4PsXWAwSQwHbNQR8WSHtYCw/7
B/BJEGN7S2j1S81dC//miWH1XfDmDbHNkkwjgmbTr2it/6kNUojM/OaKZuFZq5v3sZiTdm42LNu2
kdzUuRzT8G2KYjObfl8OvtsqPDNL5Mp2bTsHUn7mRswE058gUZHvtkiL96CctpZGmuZgfLIlS3c9
IgJNklundr1D/IM57+3H3mGvABY44RFNQrzDXMmBvJwAlv49sgzLPKqaXyC6QAgK+VX7YntV3W6G
g7xOji8pSy6NRMHL+E42DnXhQ+qZi31ps5baoSfZGaxoFs2s9pTfwMc0J8PeOrp+c16tZHZ2eFfB
5ClapHkQERt1IcLb5hE7ovvkgUogfWuNBrzy4DNW4q5p5Bu2F4wrCMfT/NkP8pSjQgEFMjYr0izJ
Jk4vFouzP4cxi3sd/G/RSpYKa6HMg7zHydKboHyG01db0vpeiG+3YsWvP1oGD/KPzXL5+l9Cn9Nm
WpqYoMQue0164uD8thlc4YP5+582QUSoK0Jl5Vh3PweVKv+Hts7oE6Fv2YchBRgHdTityVXczVff
LE1lnrptw8Y6Cz/5aK95sPE2kxcQNGKrOFITKnrOrktWKKIur6eS/DHeR0A9e4S/f+AbzO4Fi4ZL
iCuEfi0ZLmZqta4HHpMwy1tKPcxZhd5qAFvizy/LTZ/deEnCiJ3c6VAB725RDwOhTud0K9DQM34k
ceQmqDqiVFUwC1k19BIcQ4ASHRgEbWl24QNMQpOX1WMt6m2f879AQl3D5Tdmxry5zGvhFpRHrd5L
9mef2jIeyHF+CJXn3jJ/W8WH3enKL5zJB28Kqw9imf1Eyau3IvCYWDTJVlv6SO0JToM83vRQUzpD
oW/m02n7yEMdXw+9ZzHsz5268pyqZJoA4CWTnVoTnvLpD1VwSW0YtNvmH57eurfgD5klgtJ4ePdS
jbKMcIu70yI/jnmQiXKYhJha+nUCrR5SNWR+FOupjJxGEXI+D652LD4zQKWpPwvuAPvrkrXJmoDB
MP8Ro1SClMH1QQDjRVPcgEx8L2jknjVR+agukcaQYxFpC2Py6ZK/QuXIMTHo/H5GfbYiqKP2x4xG
3UUmVVhlLruJvkWRaL6oK0aA3gyAfuNi28q6p5oSaxDqMK0cxrfdvcbbhMGs8ciJSWciT2XV2boq
XfPS6kPr1ItsddPFHWlqHq03iZG5LRfTcdpyfmBtoInOkBkty/XPz9rl8D7zMe+14qCsCvq0rF8M
pCT+jLLRjboyKgRUqau8n1nDGlVcfhOzs2qGCPz1BtC7SqHOVQ8Mwsqto+G7GnAa88zNHUCtX45h
IG7JItVQyowy5kpfGOi2LGscv/Cbvw2p/idPXInOoJcPzXEUk3r4sXwZ6UbnCRKnVHqFvXZdXjqG
4W9EgG0a3DNEsenqXDN+PhcUe3l7hmHydFKrM+Y3+MVrzq3yehhg04r8XTkBrygK6C+YazftvCpW
+tZhLm7JMvP+p6n+9X4CmtAJVI8FIB/K4DLKezbA/bmBEfenEQJlJ2clyyi4LGwNtbgZYzFCCmGv
1w3aZW28aTFIx3MbUzzgsVM9ZBZDx+sNwRzaVepz3Uf8xKakb5Xix8DRfMtYVlmciyX2o6vU4umy
74EIoeJX3pCHSrDINkjv5lPS8nFSrlrm/r8U7RoiO9K19xBOMjYVZSfXKrM2+//HWlyNbOtJHshY
TconeE7Q2M05HF96Ybef0Wa78fcA8O5yZiipUbqN5X4p6nWv2iwPWHFk0yQfWGmYc+Efz9+twEgF
cvMccISO9FSEn6N0+8TsLB0nLaxCtP56BTyrXH7tQNu9sp3fjwv2HK6BbKq2jQOlyWh7EOZmZwf2
JFMIoUlUmw4kNc7tc0NHW20NEFUDJCznFeSKgSkCbHE+NTH0vzpPOfylquCBfhC42WvuPmpu6GUc
VEHJzgaikpVeGCGC4d0h7FIhxCTeDkUUxe1tJ4u/zq6jCl9qw309aueh/71jz3C2ya9Lrr+yZi60
VbmXRnfmjTOqbMahTHmaFf/hHOVm0lY0FcdbG5O2oepUS64fcLneg0qhYuzx5f3nJziCKg2B9dsB
NPSKrY4cA6hqR/BVp5+y8Lds9ZBV8n/Kels45f8ye1hUQSMeJSp4IVDES1jWO5guVu99GoogOzYW
EenWDWjBwC7CqN+e6cdnjM8O7RYL6WaPaqXFhjGAgIScmdojM68uWsiPrxgPtoKusQSAH7xKBuaB
3oUyz3WA0mbUX1WP9bPQpvelbUWdmlsWY7IyxK0R+QoVFEjP5Mkq/td12+KmgrusU+Z1bosbHqGE
peBaXICquHiYjZAybQB9iyJ2c6wdnoVpcb60ot+WMULtfbEtbKdJNLsv21GQOgRnGs0x+mEBU/TQ
tgjbDJMZoNCDZ/+HVe8oHip4t8KE22vPfWLIUJn/Z48V/Hba3jyOHk4VzGOWiH8qOOcNHJtyyprq
v33jXnaPkL0yiv86JUq3joEgS6ctT6McfH7fdomc2SI+l+JjvL3zS96f8YL1Go7F2NIgb4uPEvI1
hUkmujyl6r4pwenPLNGqGqELzv+4OqPnl5U7/wucM1qdNuv0YpytBAh5NZnmCKK2elzsc03cfYGG
fkWWp9r4WDY55/fqHduDy2GZIvTaPGePnXhWnuQ6mr57/fH066Q6l8iQsnhSjG+1EvNIkamS7G35
ekoYE5K82HGiNtBXdl7MafwCuPFlp/57yVar0FdHSl4a35ot8wsCDtEFF3droRrDTK98uK65G1fg
C+n1AZ/mrZx/9wAREX0HaoQl4r+lEu8fm3C/u4J0NSOinzjSEligp85nRzTbICSPLABUVrxG7CNp
0vaAZV56EGuJnDgk/c7bMd51unR5oVn9K6FVNDveryJWpXAIQCzoAryzP/c0FUpfwqFa3OSMLeeK
3C8QCvHqscXzEjWadG6fwmJZ6LySp0zZq3eTvSUTQ92bYMfi+pVr5nd97Astv82HTJg0VUy+eB4c
pXebjQEsyAYLurY2lo3X5UO1ODhXY2cxvv8Skvgtimy9/5KSOgopIsvrtNSpOyu9Kte0DHqEcjLC
OIUgzs8n9rN7SaGTvCzh5Ap6hDK3WHFuPW+uDs3z3r0FYxTq4hkBf/djyLkFeFc/CpFyuLWoazus
SHZL/ZMNarzaVjDcqBVJ2U2sRM3hDrUhYid83BeurPIShGdFpslfZ8Yao0TjqM0Da00panUYUhhe
/nKF4a7vqXj8F4tlY3ou9PvuEfGX8/4NMXJvd8GCReGiY4GR16D3A17BDnGjzZEA5v8u9xKoGRaX
wAzhwHpBQEFvxLrxrpn0pweeIlAf/ObHl+RweCrfiWSb76L1fN27j3cgI56JS8komZNMl5W+mi32
2uqAW05M7YHlr7JiYrJBn0ajvHYFNDB1MYF0IuGSKnz6PqScxvB54nEtoquKmoW2CW9mDE/HHqkQ
ljbqllEqCUJz1KZn162russU5frzUnIBEPJo70BNnfcrZkzJqcTCL83wtwgPPGwihJGreaqz2AAa
iHuZBbdOU6eETJrnBWYssQTFwHnwF1yoBuut3YPd6MNOCLLSXu83R6juPXA5mnQoTJr+LCep9qWp
2/w+pWj8X6j7j+1VExLS0O7txcqfZ6Ysr9edRzFMtMjkzRqzyGGucUYLSUUvjgMYLVYMEeBnpUnt
+NBZrs/psTTHrXVjuNN1CDHH1I10/V9wJlJ+hDKAFpoR9wkfhmX/tST9fO+FwErOVcdtVb3oD3rS
SqvwkxIG69ghbSBRyOLx44Z4jLyVeBrTqjBWOJMqQQ8bhXZbY0F7oJVs7O4gFIXd2bZabGz9OYbA
oN6Zi1ieLO/bZwhWygi4pEhqqxh0CEkl37VAjZNS/P5f9a00ZaoPtioy58sjULxET6WZ0h5X+19I
sY8IG1FEeKGj8wXmJBWuCf8N5VSaWVZciF6nBevJ2qcCEOK3PakwfKqzIG+QmTBCt3+SjfbWKFS7
OapN9MBCY5ZhRBNjXPKN0S5cc7Yxgpfh8BFyDxDtZxKSm2i/Q1ilAZrXGazPRy94v2xfkPoQBwZT
IY76ZxKFZC1YJiSobkorzgXZi6ovzL4QMoT3HE7zhipQSJseR/JqtY+p1T0pbDCbHhE5ikPXV72t
iSfuRmQPKOQEOY7Kx92jTxxEWieoayrt7lfx3t9qtLOZ6vpQd/fzUQ6MnjFUeo/2L0L+Yj46HkZJ
BiPWdV55whdcosiy0g0SS6WWnKjwvjYiOPVoCjElDWje2VJCkXezJcdRwAJGSXRaIspsLYPsXys6
i0CxKlhU63HeWzpovIDo5iKHNlotCg4+1RzyNijclQKAVjFPU8QAmlOeegpJqRSC24XlG7xBWYJc
KOpA/R0+5UlAlfvQsMbXSGy7S3S1HEjRRqYmIe7y0+XRixGwNltAgzXbmb7LFZG/8oGSmQsSqYcY
PG2AgulPviLF61UEq+GTxtJ4jCYgvbN8NHIRVgROVjY3O7/M3fQcgnNGWwyRWXaJFdeB8K6uuSx6
iCliBN8tP0tWaXpZZ6C1R6/W3vNfveKCAIlsrCVeAZx9Tcl2IlrVQGq+7Mdr0PP2+R1yt3w4RbJ7
j4LrkEQPAHgrRv3SEhN+ZntVOCACXHmr60R412/1vm+fBdsywP4u2fC43yNyUV4JAF/d7dmkoZQp
fRnM9hz0jR/VbAt65AaHCt0u9mBwoYnyd20ItK2TkyatBxTcWE2eiPSDbgbq3QMSh3FszxqzTEfI
THjdIB++XFGgTjEWe6Hz0nvpdVyjVCLMwAEc3Fa/hNnhCRWOlPjTsRREyNlaIWa+4KESUQSoDQlr
7NbmKnMrRlp+xgIeDQwUnkYl8F290vgNVsApeNNBlH10qGuGTrqXK6PYlOYVBZVwWTI4/q1IOEui
wm3oB8fTv1aehFcgw4YJzW/jIB1msq3+uSmQN6zUGyrECMlJIA2nrQDzMcBVrTQ9sMRRFUwC7F13
zJHjxkdcfUwpfogBEzBJfJtqoLI+y7b7f16+TBhtUteCd9ho0GIgdc6PIeqZNkavRXecsLSY1MLV
X2XuJewKwhWbgBPQ+Geoj5qfPv08dQH8/1u1maB4BWeJI/+Sju+8/svLHXXKxexsdDhTSh7WTlIl
2XphrJvEjXPkw91SopBwmK5vOtIa8zH4IGZmUN3VaLOHtM0MzTfeivR4P2VZOpKsHSztbpnH9iBy
ABS6I9sMTx3I4M1zl3LbpKRXhl/CkZxuGCPJBNpC14av4XlBeiUfl+G+ukIahyMVx8yzUXx7KrGF
T1SLq6ZRHD0y52MCI9pS5wSdrVIsO0XcZKFv5ciE4KjJFrX/4wKVh+PvA9GnrwFXOjPWTwl+T1Ai
7aXdUlSJkdwnJj9iOAW5S3B4ZKCMza2bAASWqfqvCh6uhV+XxiO3cjiQQzfui2AmPxoLY+LF+pTy
WTP4HYOjleI62zMXGJrtij9SindGw3OIhvv55eowiqV7Dbo9JVnNqQ+IYDZDoA7viv3jHh2hQ1yA
dNMyHY6vE1dfcHXU8zijsks6+14V5tWyd66tBF294/PNo7yAJz6Q7wKqir+O2dPD84iSv/kVXuUH
VPahu0ANawal8lEVEikvt9ExMXRzMCi/aQSvn0S6pmZXifY2WdqHQuWXrnLH51+QkJ/80//vuM2q
4IbmLSDGqp6oQDpZfD7oLiLV9CSF4rlIZnbWVNhDUs1zGabPt6PJs/Ggi3F5XuiCgcERyje+wjJb
xPBik80J6RmPDap/yy9jdmOVZMlV96EvpAwIu44n4h2EuAbNxnpxSpJr8B8VIpbwwaHhNsxRqDmO
YyJ+sKCwpt7xuy86uifumlxl5E3JBP/TlG5UUaWqD14XlpdJJ254/I4LzQTYHL+TYsc2ne3A4+vL
fmNaIsh3l/Z7Y45xFJNyFm3Vb0OSl+sGV238TO72AHyyhuWm3v+VyZ+lw/wUZ/lQteC8vIQiUeyN
b42JxpeYhdWa8aJJPOH+kdjxbI1LziINproswA/yPUOmFtgM7RpONRfnY2ktmXz0Y5T6nUBC1J4B
KTtqn6VXOSPaZSolMGGp4kQTZYK2qKuo16dQ7Bq3uR+cOA4EQ8/J17KJHDY/mdcV/7JBKkLZDWAO
U51taDbwjJYiozFp7Nxs2ca3S59U5teRRJN6fkZOgMylFszzDMwf1/dNFeuoo3mw9T47qyKPpOQQ
XHZcIktu0+T8V0AW6NdgJGULZnYIgCaCEGNohIpesSWJ1MXWlcsGl2eFh2niB2lvF5PgTHp6IV+5
oSctpMV4uEomsxNpg+aolnJxUGg0LL6mnOF+6C36Ew5SPsZQbnRXk8rbZArFhyvJ5BfFFuSqsfYi
P3rWXT7UdOM/vhBPVFFBYIUYObMhQvLRqMxzPvhF1ZW9onUoJv5s4eGWm7VYPlO6B9IbFw/PZGzh
e7IgNRZgwhrRZkDvrYbRX8zmcAH0xqRJxzxILnK2DaMb4imOI62B4oanqTc9vMwNsyPi4hHfSW4r
MNHTzpfGDc9/5TPwV0EzpgE/cToMGFrgKPQ3lbDpkZULLLe9W48rw2Yt/reVpgmhs5gMRrHdt0GK
gOad1JOoBQru2h+6jUKkOBExxsKKD2FCJU6SPjfo/Y5mK2uxLOQrUDQ5TUER6mpyDNFCvTJcqryw
yvO+LcNPxPTymwxn+UIAqyolb/4OMi10jR6xi+qjdJ/6t5/now3LWT0ESticEolopzQZ3/aBa/zQ
/6ltbhOY+hIlR/hXzGlLDlRfDKQHlNHuxMQBzC1hTbQPumOJGpzp08lgFO7kpqYj3vBZhYWH+Jvz
8zlFj7sZAahEHkURZbsvrtOCtitIGPZQIfMU4fyWtgTCSjBXRD2QOGTlxTl81Ho4eCJ/9Avnmku+
eCfqemxA6hxlzWNC+e60YnnHefbolEK9gvVg/tkqoLkAH2L/zLG1pXhaY4LfmIQHLzgoHTSlkxZY
DigqfL4S9owLWU3VeDt4FhDjEo8wlPsjyn4ksSfjSh5wMFZ0MDZ8mi/4tMA10YGEVZAtqTFxh2/1
UwnCL0RXQbRZomjMFlVRV/HKRfWOmKPMpStolaBMCuyl/WSZGhmoL/EzHfc6966Z+avwD1vxpube
NBMkFmEbPquvWWax5MapDOGS+ljN5KhemAnJbg+XB2H6c5mVYSgyCvcDKoq+0/TJ2RVS7SD5bXi+
v6N320h/aS5ESckNr2o6gjvoSImIaIUNPlgguSNzEPHeK5mndOpvcOor2P1DdrDT6SNSwh+QOq9i
f1WU3EfmltCaPsW69zKZMn84g8g3/KLlWbOj43TM1uCjG20UjHJZ7LbN2Jnjq1mNE1rS31LfWRFW
ElPUAMYeQm/8Chg/yyORk3k6da/a/4pdVaagM7Fnxur0b8qf8oDizzdP6HI/mmhEYtgwCg8Dp3OD
5IUw101hcQ56xd9XuCXx7T2vjuqLi7C0Y1wLFYMNQyrbchOTE5nw7zWJeJZyLRfXxi8HxSsaa99e
oI+T3b6S3InhXDqNepHZcFXRsroB5C5tgmaCibviuLx03xV2cqnSspM2qxus0VqK8N0MFRFdkK0Z
ly9w1BYRSrOnnEhDtEr2g3B6zlt+sgdBTgt+l45VulW1IOrGGeKg4T+beyVSkKi6dvX6lbs/0KUG
0lQVCtsanK5DyzQ+/epWPz1mtr+r4PCy9M3GCumBVPspKoDbVIhiYsbO03BgZRzwncrRDvs6sDMR
rCRk2ySoh9MSWbCAJQwTcRCXYc61Xk0/L703yemsUIaky2qdLkGEtyVZOd3MKMs5QIfCFgPRcs3k
RfmAthNPKCbrFMyYgGkrBdFZVuqfHUSJG4EaI5qrKt9E/gGuG3+RHqACkAVuy3gO60tPHWPtpFio
9+5Fd4JRDRG9k4cMmAt/kh2G2W8b0MTQ2rhJTGMUVV5sO/lPjKn2PN9h3fhf7mokFWL1tiJe57rA
Es2AUwkzW/UoI0jB4mDe9PL0/6NASp9BJYPQvYSDssrDxew1xEWLdmmVPaIfRjlAL6prnQ7jQtNO
uIhUsKzdfFdc/XRExd7RsgGRn15+wHNXcmvBMvTPwhOUY8vdfYQxFhbJj61IC4ZiB3GvFHazXP/Z
bum+5q2clTga4ijCOYY24GLZK0Z7EGDdpgTPZau01lScqLVJ0bYy0kB7c/KGx7wvTNxgDQ5KnrZ1
TU+OJy/P73Y5yPftByLoxwOF8AlhF0LlOtt20MQyJT9BQgvFvyLkJE4gPyD1KjBoDIjpSJHLHYKP
mvBHnAKChxqFcMJxAGJZ2CBK23ozVpa0IN156GYpLeaZMwudeWMMQXs/tpIE063kryJVi8QuOFsp
z9zqzecBgHqO2S7yWdcCbwnW4czsS9c0jMqxClEIQpibdCNPKGLdpRBlHn/KIqG8KwaTidyS54RQ
m+Opd/g74fw1Pd3A2C+WPIopAJu8cwAKQIoMeW6Y0lSBEmJp158Ma9QZiPwMg6sFDLBwiuMbHmlw
fkjPJFEI6iz38CxpDsd60wDis93E3MbrEiZoHm3StB2OYnH01guzYXek8rjuhJhM6oisj6MAL99s
uW2GCh35B4owFOtJq7uTMGHUGgkokI9HK0QsdAQYbtNkmmkRWcPIudze0+ysK76yMSXxiV23GbCS
ns1cBSVKtQDVe7D49IdM+hAWbL8JgDeK7GtetjRkqFRl9udz2n4GFA58xSLiH442tnXKFIa9pAyV
qhwYjl0o+CsUPVnRZgmA/VJxJ2F61vb+gBgWRZ5RySMt8TE+oncXEWRZ0sArm3ICUOwWFY7y3ih2
xW5+6aIVwIn+YqGmqjkqiYajG3e0fk4Wag+sUQaPM/u0G7GSLjm7NajcyyPFI89qZ8oFxQr9jNRH
CgOCInyYyQUhsf62PCee4CIyJKhphNsPUbggK//cfL7bLC/3gikLp6J0LfUnzAWzei9xbiQigDXC
BcwuhZrbMQXshDSsDXZuYXDuwE44uHE2elq2TiQd5VY846aOiDKyOs/6/jzj6/8pSAM5pOGBvnvA
fRbV3njFwHUq3X3STzgoHZnD2S73NdojaPDKVLVA+7cxR9LKWEuVOGiOqxfgaVYX9e52yCwcaxC0
7dqbJ8q+Jr8XwKZt8FysSz2MKsPRWQk9tWTJxPYQZxq+q9oFPc+d1AwQXbGh0sxFrYo+Hdi5AfGB
HBhtVxWQpWKV5D2ZFijhZb8XJdtqdeAMnIWv09wqJtpd8kGKG98k9q/Z5ojm8Y+rjt/niTnWowi6
weeI9NebVNL3OJW78P08cR7l7BNU+ez0W/iKWilPW1rCnH4HsgoTnJTAkT9e/Mbskq1oF1pVPNsn
73QNzj89IKjFoXBRgPwomB3QbY+QxQCj9f+Vnxw5aAblSrWVYjffLfS77I5xQLw6adi617QwnVho
cJAwjLN6hhGuBPS1dFHt83/4DA8O0ENCf8/bibZGcePgrwFD/vqcOMU3E9XV0/DhNVIw4r4JEB/t
5rafUf92X547YZ2t63MBIXacsikKGg3lLFnX5U+iLeMA/YOAHpxZBB7GbVDwoarKo2M6/ZrTwpEh
/Page5kBiqk8ggcovVNrczzmTTu02fnf7C5AhqJCFNcrLO/EdoIyjwJGKCTcP+u32ZhbF5CdWXZm
rneQbP7/EUuZuaWSkfoUd1AwiWL2hn/UznBVrK4mZVQyGsXj3aXsc5BqMPgGC/Hi5LyaFoZ5aa+3
l3+M7/nY6onWlt1ngl6n95Rc8Mg1n7OtmIa+67TPk7h9XQRo2mi/+CKycdsVP+zn/p3zq1wzuDTI
/D2MfaFQFVG+WnwoVpGfy6Jh0x/UbrnmJ3c1b1A3vcwvDtfcubVM/psdxYdD9q/sLz3fq3/oNVRo
VwwxZKV82rgnyGVDynriuHUOKaS3X4EYcBHJaWlpHQYvqeh9f20vza0uJg9rIvCTqs8Xq/Bi5Sxy
OIzQWvg/or33LByrPlU2U9dtdZSVWvWoHP7pv7xi2N4DVuSQiPKSzxNdgTvCN7O6yQZunCLuwWSa
WeLH5Xt2fMCX/9Mhx6IADFd05a71A1Q2JOskl01FCW7SRLvKODkg/tV9JPCzIKMNds5D1YYqn7Ws
1RQmmx4BFNG+3NYW1kf0EpwEO9DaVstegDFGVUIfKtHYqzcYhhcoZTfOM2IsNF6AmFEpumcqlOqa
gi+2hVsxL5t/aLjwd32YoIElJXo4mWH57tRWqLkiF0pVwOuqAqr3GNzDbgFM0B0o1EnJltJE9use
6SHsXcPuJypXQnT8MFws4wAhQ63Kr+7IRWdCKt97+5+mELXj3AJdoGysXuua7O0d+YwFa5Q10JD7
hqY5NOjrLfOYjkXa6fb3r0kAgLt5QvJ5Dcg4deq6i+gaUtFxbItPODu5HcGHQWiCdCHSFyZTRfQf
zBTZAe7M0S67EsdaxfECHajSmQUuTMecjDqbmTefBc0PU+zIsOJegaahRtNGBFCZxIUaG5EVDK1h
pDVQheuPmeVdUuVlZ7qdbwWIzBEk2vtlK9DZY1RQvgkjbYVdmMxdjgMFtcVuz82zrhaTMWx0MdtP
fmGg0GDSKJeCAO9xVfUHZVpNdlffqMGlc5bwBdYo6M9aMEOq5hs8tTM5pBBkCY4F/JqxHTJj+aW1
kVE+pK/WPzMmWPBJfZxU0dXz7sK6F1qbEyp5tysXS7VPRSjsprBbcgQH0eTN2BwsLDJRxEImHs7Y
ga+dqkp+5B8AoH4A2rRoRj+SnOMgcyOwteuegT34VBSvMN9PQ5CusL7oIG8ZTuiKVyXL6fI7/HXA
M1/pw5XXKb5FgxqSTILQY9EEBnS/bpCOXhk4OwfQ08ByXC0JSmH12KWTz6YN9ZqiM63ugLMoeYqP
woBv8qLiQB3fGYLHgUL9fWikxMAc5IGz+EW5OZUalgEwOWBgq3neaobm8yVc+ZOSw2Kac2yeFS8t
RjXk+JaVS1Q35BFCjNeXRtvgdVs0v+8+5/WIgD3dzyiRbf22x0aSH5BKRV1ZroDjgw5+uNStXfCU
XI7bvCiWIGHXZvZviHMNRriVdevZEBLmTaMtwF4hOuB3op85tUZYnJJafqKdgOJ2oRXCIo2Q4rSL
wwzR/zj6OkEOM/Joo5sbVXt0sf1AqFOSZpOyAAGWOppgcGuATVVpZT8Ns13HGHJhlipUrkfCrOa/
4lRWCztCd5uJSfhESlYheMP5NXoAmSIoxXrIpj9rU/nYwCB1PUFoC1D5q1E8HSXP1d01p7tidIAk
xPy0UgVASMG+iZYXaHR7iS8rO5AGdDQP4JgPILdXcIwuVHGj7BSk4yXenPUWfdm+8yHRx0T0o9NE
7gEwyETZwKxdMe+6nN/y8t8tCyjj/4W/AejFf6X2FJyOsHetVZG13rG79TFIx+WHYaZVxPlfCYM8
OJQkQWWBjMLUzG1GgZF3Rk3vgPGb8S18yHHzgF+rHwYH8LmIEpTBlVT9GCMrDOLNP6zxGMtddbIm
SrqTKMLfPdIs5h+OL/zwLvLHTl/BVvCPtyS0FjcaOmXbN/96XaEO9iCkE+tCgxrzR/itRyqATrjI
na/fMoWsaTs1bnLyEvL/7SgKU2Ipn6LChfSVsHQPO2VWReNtoaEQuffFSchROD8/L3+f4+brpHCj
9pEZ7SWL6lXRYlrAmUK8fSkzjSiajigUvtmWGpLIpo0GZ5VO/soCkxVa8aFTQQBM+7F1sX7I/OF+
SFyECgGMHXRFXs3+EcxRJCYdtMLN2nQL8vyL3jnpqu+vBEFaX8vx2P5yLmRJQo9uMcpTDi+LvXiv
BnnhBESqk2BSajE6XTfrg0Gl495H1s4PpLIk6d+EvYTVF99/zNHG4Di2qG6kGaGD4Sy1QjMtM/tm
LV7N7qFonUcELSWwDFQyFQMcqBSqmqEjiHc/avdruRlhswrWpArdqzU6jvkNeEi4EP3tPBQVu4wC
6hPjU6g0y8X+qD3erzgHQzH20/gGVZcRNDlKxUFoaCzMw+iojrczrMo697HJe4m5HLl0WIbCsWEL
u+troZoCypxt3hm6WBGRMW1giBNq12OeKhfEz35uw23I8napXN78NXTjKEneueVMbIiUpULtOOef
mPXhNhXRC71niB7WHg9B9MEj1oBDs2YL3p3PMgGOpe3421LHmNNElPR0vg9XB46ZBzC4S0EdeLmQ
xEQh5o/x259v4PqAmpuC56PXyVMOgS2relZ2Cp4pWCSNVfTqLJNnDD9inz3kPrAHUjYNazG4is/4
XPwB6xyCC8Tl775jhNVrnXL1tTEMHf0TPVl4gcrKsro63eh0GyPrFEMZYtsrCEBYXzURMYufovaf
nHhXug5ZtZXQFSdllEBbHcVI15KuJJxz3SvHOUze7XyIRQdRQq6dpF+Q95bpceQZevciRUQRa9j8
pjW4E5sAixXwRCLfn7X+CmYpy6HhAHBGRaPm8VnuAEvaQTWqu9tqsmOdDb0gEbG7FlDAl93JTXfH
WJA6MqTyi/2IhDe6fIo5b+YSBut1E4B90S+0Ve33qnxkmh9N9fwDdW55u9MzLWAXk8VtKkvQtQD9
pRctDOAyUtN3EWbV0aWMZw+yvIMGplBpwNC/A5K/OZTSFvfRj15QX1aN9iBtCtZxtPNBOvaH6v7E
cm/OvDyikoQCQDCcwM3hZ43kzhLmIBfvtLjpD6Uqt9o1bFB9s5p2kjpD8QECIBvK+Z9Pu/d+qhPL
hlTvr5O6PloedRFFnGiwKvGvrWvqutMYzPvevS/Ni5J0zWWDVmdyiZYVS3TKtvLlvALPyHEA9YUU
THGceJ7C3yT4KIe3dZJOxGTjjhDNkQevS4O1HIBaiTluerIGqFQiN2eXViddlSo522mTTs1lBtXY
NNTpkfA4O60idFImjNQUg94oy/Qd53cKrMvCQUI/Zan/ke1sBO7a75cbachZbpuTX/HhdpxW+OPH
2jadIPlZ/is70yk67JJYuHNEfObXlBzRMj2iE3WLxNl4ipNyHmTrxwRGwO7wSsNbvH2ZSRsag0zW
zxtGBPXDrQtV2W/qw0bLRhDi48gWv92VEBwuG3UUY5zHjdC86F3Qx1TU7zVQYXiFX1Bi6rTZ/4rx
9la65a7cqiwTEKq0fXo29vyViLZ5CZSwOk3ic8TVVUfaq9RGvRpVE5Kp748C7F0yXZ6OhQl9bEaI
BmcCbT6z5msA4qeFlKZCQaXg3ZCTWAth34kp3L6lycaX44uCpCoaxvLnNToODBkjJiECCzuNMuU4
2KaAdBuQDNuN1MPxu4Mqsbh26M3zGpQuaLiRWSWmYPTlx5RU3bsGXe1w337fwqWnhe/r5uKJ2IP2
gnLzsFVAk39+Xlw71M2PqECtwClhJ9vlSy4jNF3JYwNXl/6QAkXaoq2NUhO0uJFe3W9IBd9E7YoW
zwBRKYvj0ERCbSiH/gYiBb5s5Ar8Z/8geQRClNL5DBvs61sM3lSG4WbpOXr2KUVilctsDe413hiS
EI39UbWrGzky4No9nzvsDfjB5ij1UCqjezcCKfzW0RplzIv/o5wO8V2fp33kn8+a0iuV0PtrCwek
+PHvLvjoGyHLVO6x8xhwzC7yyvbJKM1EJrV77At+EyNbG7su5ReR9IZZP70y7Avn9sVNnDIZuFsk
Y53XWK+1FlmdEwV+YCHmek9OdRMoLEmJw1bF1DyzT6g6ipxfqjROQj80grPZuQjkqWkObh30Yov/
GFXuyMFJ1H8yJkQZXgEmsU9Yik3i4BoTeoDc1v62anNh3z357Kx3b+N/OIQEDDBlhH0S8qTasq8H
LQPgW4cRXM3jv3APAkv4HAa5B3B3qk3jmIqKIwdhR2auSx9c8PN14amQLZgU7d8WRk+rW05CfNhj
pU21Z/rdVPOPVUefMkMx0fTaNux4kOTTfiPO/xza/kWOvrcaB9HCmFyWnRem9XVv0kA6bAbnUCLy
AnHtu3mREdGqVRMnAwWrRzIxVhhcDbSImYM6EQN+8xArEPxw0y6HaJel06++qi23IEalODQmiwX2
2Xtf6UAUYDBP3aOBGslJxjnZUzkzTf+wYcrjEZPFC/YS77fZ773m4vPcyHkUR0pNeJGN3rqCDvH9
vpHRDQTnoR7/tCM8MGOKahmwyJB068DVU21MjUek34b9Dbcq7FZFev6HQI0dCMdTZ6E7/MsWBZqq
RJKvWo5dUFg99sSKAB+Vsva7gpO2WqUKGkeCD4sjr2R6zz9A6pG1NSzUmRi+B5G7ze++Tk8gkUq4
D0LfkJY39G5ZkCVBqzHE3sS9Dh4a+valiaDZkwLx1QNTopAENSuWwoSiy75kmMc2cxOGjzZAXY2f
KviUvQiDsSaNlpCKXadZQCnQPwgHnWenIfx1iGbFOsDOwGaoaaSxHfUXcDc6v68unnanEBgIwled
oA78eKlwXdZKNcCLuxoEFyLsDgrquTtNqWDa7Ih4CpXNkERWq30PD7E3XAwgSQPSbA7zbeFaOVXE
o4rckMfNbf/5f18WXaYM/51X+XqfIKBSTO2itbO7hCoFTkMIExWh9tqHGRgIVft4FeVODfVSlhpt
gom9f5HYSJzZjRgGKQBuaTM+1gK8evgaH5pFleUfnpdlI8mkoL4mIUuZxmDQOcIRW5hAD+cioeE8
yPpzc4CpiRuiCqDTbwb3UDmt4MhWyf6JK2BgQ+7Gk0uptj/euwHSvDvKCZOYc9zx3rsKbVMkvCtm
99+BjjeCLrnDZQqZIM1t59xEK+n5cigpIgEVAUDd3ib6KYOagZNQXJ6P+pk2WnlZB5fZpsQ6U9vV
04exOPEgFEkIhYLxhFLdDqNfXyOC9cvqooBah6c7kCwfTUljeXzSPDZhLsTcR71IX4ur+Mmpo79j
IGov4FnAch6c/NhnX9L8p9P6UnuBL5818ax+T3relEdN4T6WoAKsCt1yZ/wk01VwSjYGsqN2LcAf
iTfzxbs3M313u4y44k7KYR30n4NHzQMXlFid6WSJbWBoP3rzxgRIHmkg1A4rUcQXbv4sSJwACsMn
2G/tglMsA4368tfnmWmKHeE4kLRH4vmkonTBkw9l0PAWAmvVuXNawyNo20XXcS0VOlmBq+HOAbZt
xO7TrOOcsS4WRU7m+yX9oHSK4Cux9Hr0GZNdBYvremoydXEpMTlsBqPF263X7KNX//6RRih5msls
BSG71KGgHN2aO/EpS67SCGPpiirIaCp/SsDJGALGm+9ZsiAPGcjqgDBnYQ1Xt3pVTllrL6KkeRgp
fiDVrCSAaiNOZ8JQjyA6jjkQpF8ZEv6YXo/YsOiSK1R/SxFu1Qna8DbCjm+n9ZBDW8VP4K1hrBUu
lU+lo1NinAyuY0jkZTr2KSfbfVUVT2opFoptCNqxrq8lYtAC7Od+4JdryEiFIAU0X5s132Qhvwll
jIOEuLB/z6yWhPcZ6M7PtPRQxrD6xy+LT4vMYTD6rbm7JRhhu5s9u6CtUibiHVCmIZwrL/hsTPfe
JQsE+pKoEWMFdFYSi6qkJpJHC4Y171qk/QX9cQ5e0ocDrl+WdtRpu5cZ2br6QjRaCxFSgYxxACX6
kPxk+iCZpYKruPQD8or6mi3pNCj3ffRkTrus1mLRXMfy0KquGQwCn2pWmUc1uGPLjBLJzq4RAZZQ
8qpY/Z3hw+78jZLROBTtbJISPfFa+pikAzXP37D9VSG8uK/HNCIT+Sbt62j0qMyM7aZMOexq5tfl
OUKmUOMYeO+hh+q3vPIRDKmv/e8Z3FW4XC0A59D8MzFeR8BDy7R688shq24Tt71rzfmr8UEOGCNG
4wcPSf3b/Vc+03nr0bupOWoSx7baBnngz+R5dnY1NdfC45i91IuRV8lvBnQ6MB6B+NjefkwLxtMf
n8bNgmCdzI1Z+WvT9lOOFNjoG8IefBFQAGswy/uLzRs0WT1h9nB40ghADzoeu1dwsR5ZQ55Om18x
uTYQtlh576Y/QlHWD95aMPcEyOofuZMD+VyIf6sxvNYUxLwfFjP1rftEOJpAiTvokxrLNi0t2Sxg
wzfuuV5LsQR/6FWcdT7PgPUNMk+op0tPXsIjWKyGEnLN4QRBApvbIkzCf7Ep11zofeTc1nRRZMGS
s01lOIkC4oYpEMqS6mmB6mvAE+71VthQGJE5lqjzfLMTNpzFofH4wZ9xQ1BKnQAyEQfNvEr8How2
4x55vX87ZFMPwwrQ1UvNRnVQ1UKNwHTfK9ux7D+4hJU2hNnaT4nU9CaAOZJtRQawWv/rG1IDzRkN
RcxfTDIDH5TabvGPdODcujDXgorso6zI5FtEcMNubQgh1X/9MtImM1f5oP9Gd1ayQrt0zYXKJwV0
PP1FM4oJR92eUtJ3ksCJLOTWgUCQTTy+brCiYqqWGT8XcM1DfNm4X44Xwtk3AcsqqsQCZYQbMaBy
HxCWJPACq6mxck8iEX4b7fcCuzBD59pvaib0H2jTcnxrffPQtacp/4i/NiWtc/TJUX+/g60grUFa
6PjIA9WaNdK5JVMGqsMBxDi61jFyYUJO0V6lTHxIujjFlXr7KQiVicx6KzK5fWs6ei+9swCcfryF
eEDIxlcdIqgx09s9eqf+B0M2i47N8isBPxSs2t4JAyWt2i2LoT7qEB9cSlbaT4sAxWd5A5ho3jeP
m/jcEbZNsQetlztQ7blK64sP6wJnqijRkIOqClHP6xBa8bJUAALgYVbdr/FjUC5KRcygFtRZQW3i
lHpQAhyutmDLDflQ8iH4MWu3tFWLiOAmx0AFzmDYvfkM8ki/4Dg2w5zOMWZgFhSMpi5TKxmAcaE+
KYMlYwk4DHN3/oURCLFBNLzZRQQ6+LugnTTo0XZYDz5whO8+fCf978KujqaOQncC5MzYzvChaoby
YwGmHKUAh0jvuGtfbW/dhfFqRjbAs186EQnvOPUfzjVM+OYLTxCxvLpYy0iSAHLv6MQZK1QIrnYF
H0GDHFzEuN7L1Jlob1F1sTiHaAFo5u/dcvWHFnZzl1H/Ni9bYEsBfYhhhh7bfx2eBDfYMgJ3gua6
1922MNNAwkBZ5I2hBOcCYG76vS/IUEWkvCvUtxRlZrLKUW0xZTOGmmshQS+jTfiWlVXu4sHKqhTs
aTlIL3rdRcL6LwAjMM2TATE3h7g0vRzEEXw3mpNr47cUAogIgPEo+M2mpCwfxaU/TFW9P3NqHz1E
oJ1e2D0ycl/x94occ2+3yLn8sOKZtOk6vdcqkldr2ZFSIkFujwFMSVdpVfKkI3/iFdAgxhCwlQ97
f6drrH4+mEy5RxQgtbpE0CoGLsWL7/8YRVEAYhuog5j3QMl9TBLILjMl8dOwCbOle43uqNg/AVYR
T56B87gsn5f3tzDlRuA4sHwQ3DXoI3zcCrIrA2PCuB64FJyZEfGnU+RzkMQE1IG16L7C1DCXFOWE
E36oo9QGaHAuS6MUHLpvVTJkHcjVd8v6DpQmrP5ZvUolasv1h9WTPKoo8pTBruzKJf34h7x50SNc
9O12Bn8Zpq7lLu94eceVeghJlRiQxjriXBjRgYsaN+3VHcKoobx6NVVDFONpWiN1oYQFjiv1CqSt
pDZFhOiSZvf6st/1M+Qeiuymw2w5/rtUddJHwukQoQfmgZNY3v0p3E5b8xu/5gU2ikeKJbojvSzV
4QYBKGqVW88renp6517YRDWyZhbYT5S0L2ZZQ4gV8Fe+xJ0BSGs+dPsCGbR6Eh/eF7ujkW/6/Uex
9yjVN5RhdoXDAsPQfineuiWkVkfvDRXQauWmkdDPS4Bslc4Wli0FRBFke7GIEnLk67rph1tXx5nG
91gKxTQzKh23cmKSXhJRrD8K1aI4QyVz7g12xTqcPRd2dt/hYJsKwc+qxMdmUVGQM1hJB9zb6Cn9
Z60HWtVs5prO8yGpgsAwGTkgg3lA1fSE8NMXXTQtFIBr9M3rNh/AHRt5q+ZNhnaHQ/l9NziH2AKR
J9KoEOFemTAU3HaTooSC2menrSDsrm23fPOLu337Nv0pTqcSwJ+6u/RpJiOPKu4iONwlj5XVi1JD
hxmw5JVpZcYOHEmEPAGp6wSOqWPK8XtYZNC65NNjVRyca7mub8D88u2eQbIjxeXrNcPmcvSs99UJ
s8Gvr488mQhnCrhmtGr0x7dhqV9+wpBtyyhFvM6WXF4F/WpzrJ8GWVHIAJz6qeIAvUI3lXi8PyjJ
CiJCLaY1NA6SikkDymytd35cbLgzqOxAlN+ZwWDURTueFJmnJ5YejGBBi3UsBEnjOCTPAI7/K/Kz
ytdSfh1JQkflgzXm0h25+9jNeotMCM93THJnrqmGugQzEqqjcD+pwRDEhkH5p3qayD6pF8wMqlJu
AHMlN7RFyr/9lj+be8eJ8fnW/gYiWTCE5tjC2v+ffaUbKoaDzNmN5TdUNCzOfaU6YoUoFqMZeFek
XirogO5OwUCLvaAQbL6axh0wpapoKM3rm0lw6pPKuGdD9bsPEquXsdtsGS7wZaW6FOKZArARBoB3
pEkQ3D1xzmFcFdzbpa4i6GOoIR093hXGM+3eFolKvi5Gy2Ne1v3owUiX29mtnDB99oovu9n97+0K
ESQQq/qiolPJML+j83XJa/eDT5OfXyYMJOjbRxt7oigOreY4PXE8nYVFyQQdoKzZ6oNsSYEmBMjK
7bKLWAMpeGQSG4qEfuetFkVuBSmXj5BDPAHdFGuNy3P63aHsjcefPnO1sWWaELF1DjZ1Fwz3KZRE
wASLSvM49a3HxGNQnZlHP1PmoP9h2PMeiqrF1wr+2hRtMCrEywUhrqmcSJ9AT1K2RTYCcoTmN8A1
uoVtchhmXhtzadsMuOPfAu6O0w8j+T0jYHfbdAu5A8XcYTVLjH1r7l9jj1hwrolFt91PfinLMzhO
dKWcbG/onM8TzMyLwPcJDN6hyK8NfL32gCPFvz/04ni/4aFtU8AZPu5A1iT7Jgjdch7W9dRp3Z+6
vpAn9bKy5x4OSSMGlupBYrABZ0h4sbFlBfIwlFhby/UbPfp/2BuNJPVWSmTSTuJzbA+43iEzUA4s
LS4nBNLfEl3IciHg5r1NAbS5+gHKusGBL0QpMJ5LHagPRfkFEOXF7GsWqXrScXE/OFcVkRE658zZ
ge+/bj+DrzXfuwLN039Lpn5zbyBz+f5qU1J5QhN80+bw138ssVV2ICxQB4EfK+eEH3Hj456Uf+VF
zKHbY7YYNxO3v14+V1SmS27SMER68UjPHaN2M3GBsu6mjttWkv0xDaJZ2f6M/XY8zJemrGHKlOCo
nM7sv3tdqm0fIBHihbvyo44t2pYsbLQEHY6vbhiKHDuPqFC45MpYkJ4RIW/kyoq9kn32DG1UTqq+
a6PHDy8wQBe+SLAjQj4WoSYEmdPuf5Ld+EoTD9vaK9FsuK47OaYJJ8pODwR15ceWjhXdGDFQAPVt
ivLUzkReIs9NyFBB673rn1pmTOXO11tThT6sCtRFvnumBLwr0fHxO2GlbBFV4nszEkCRLTRodhdQ
wHsTHDn9P4Wj3aCT1eT8/Ej4JdxlTeC+uH+1Yg+qugW+crD15sNIDVyQXLv607G7fQzhfYv/7/eA
QcE2BiKETAVjVk4vJbMCFiSmcfdBZrxMb2VMcfDrOPvPhsTln77TtdyOfGtRjy8LYhtexCACSvpt
9tHVsjOFZ/BzWSXL9exLnNwM1HkceI8n2pp4XIdRscMkBld4/hbjJ7tLWCHgVkCIsSrlgOlYVwKT
yl/QvuFYREKwaxFqSg7Im1aVmNsCKaXWK2NVRH5kT2iTN9tKNswSTZAAzJrFxXlP2SFwmRSv9PTj
Wquuv17UPQWNwc9ObbDGS+skEYPlUwutLfVGHGwuLQ67JvQ9ZE++7aBlu68TKaM3bMrsJ+YO5Y5k
BsFTu4vm5HmjtEThPKm2nNnwCWZ8fuvKRQrRqnL1AYCgOiGr0iG7XLMWhWPf1Phwc6Wiey7m2eTJ
Dq+fEXtDFPh9DVwYeYTV3R/RW8v0QEVJ0O3bWR6SzTi8w7HsJJigQErY0ZhB5VcNAUNH0UTG7yuD
p6PJi92TfbDMQ4FdsV61gnbyiCJeS2A1riE641liy6RxFA9EtVRXHYipAyk2JcSQmNVU86DhRWh4
uXqfQeapklbhWuT9/iMyy3EmTsMO+X2IHJqhCU69NjcWEFd9S6e5qIDo5YLZb+Onvr/TBiEyRfnC
S0nxW8zzGcnNGM89VEs3BDeWy2iACv3hbtEquw2VLtX+u2pwn6ZeKueQaZ82V413m953uMl3BAN5
Pe3ZisXXVFsxmg0zcbk+ICW5Rpobrguxi8mbYba64EHjoTmdC1SiW2wCklvtr7eMNv5zLQPD8Hty
EUgo51lU6eCQPbSBg5/oIJ+sIEoMPrey48qCWNXhpEUJc2bt8cyFkkGckkjKuY2kGmVZGio6hN+r
99Lq7/wB5lq2dlv+EVLNq5VJuJBFutWFz7yK2EcI8YIWX6c5ZsNMQ9YS0V1QmuQsvvpEQPHS+p3p
FQE777vq1MSnq9FgEIFOspaxUuqLd1VG6BALVuqy/sAGr5a5lgRdpsy4vvTlnimeNzWFbeT9Yl88
uptfLvCWUdlRXC5aYatlCoC8v0ufM1vBI1n16zB7CCyq3iSbtE6kKkq13sFpbyn5awYNiHG4xHYE
XX/A/lbXd3mkU9iLjhgCv0y87EFGq/c9xa7xfy0yfZ4e96UZ/FRdjyLT8mYWYu7LtGtWQOUqBFj0
6Zy2ZQAIuEz6wMAzTAg6OPNL3XJr/Kkr8Ccu/l3YxgDugZzqzBfChbZoB9jn2F6a/Nh9CjFPDkl0
gtcmLQHi9bfmQaNFANIqSi2acvhJazj78VR2Ws1cyUPjRqDgYRQk5XMhmvZQLu4ZBSGhLmBqQ/1N
ec+Q8bRt3Hp9H3Lhg4C7mhvfrwuhQW/luyzezADo9VIlYi5rIiL3MTP/JR+YQDEFgp8QQFkYNI09
LV+ax/+jwgPh4R30wK1gxClaBShTL2A33Tt1cE3hEwlD04blE/pA7UbKOk40uBh+y/J85F8c2PZg
YX/FLeKs8tUFTfJCjAKFxMM7mEcr6FFvAJ7S6YOB2bz6dCvaQ/WDBmnPbodzxhbtfFDrBkZtrnJL
R/9actbCtnSJhCxKEYvhJ0VP3t+EoFpOpSKA2drmNXWI8RZMQtwZMbW/mUvfB78dmLDNxOb1fJKA
e07KS6Lv+pa7dNJYmcILuymKNd2cnNUGpOgoiTsMuUsqtHJmtd1Lj1lkaqj0FVb1TUEAA8DKiVte
jGcg86Ke+T0+sEqjNgscgyScgn4fVGm/g5fH4BEfk645jmIjM7ciauFjW4fH7IuBvyA6bYK3bTVQ
/RTriMBBMhuXiFvFIFe+xMj1x+BeykuT75C0XSao1RFC6h1C2eFvGGJd1zlbIUPaPRGGL7ysHWax
ax+VNHaSLBJNKViv9XcSu1lV1AUfHxfQ+GOvxgeS/fl4fFYkJMhpNp9mLbbZXEbmLQQZ+pc9hmIg
/j6TVN7GVLNoMRmGMMKpBNT08sOvgBAYIE1T1o3aYgQaLCk9m5CSRndGFq+ESo0KrWW/odpHyLtn
lMjxi+kM5/UMlZWx2c3/VtcGaehy1Yky7T1UwL+2+ORrk/K+U/OALb5/AivGy8KLJBuYI2qoBs3J
BRa6ioBPNvQNj0pZGIYxuA7OTeUC5XVAYqtajX5u9WPKzMF89i5rIPy8l+EWPba74+qclAKjgz1r
3VI9eqHBlrC9xHGEBMWZ4bdt7JphhYBJylEmV+3L4MjhpA0eXPmSlaQ8GMLsQY2FG4zyfhD80wja
CwzOmOF/2OXwzoRR6HVox7AhgypJSA2m0a7Aywllx60EB6UvY7MF4oAbTUT8hzWk39035+mMm/rP
5MP7fyKyN+ycUlVDCoBjc5V2n0C+KvB6nq4eqTYMVdf1ApFPL1LZxXZMpsnVp8ni+rX7+2SMcP6w
BWY7j26CaBMb6Oegcu2zBeihCgjjBrsdzKNGEwrh0whoafSli/4Z6fWKUq27h/fjyGtsSyMVv72l
yJ7PKXkwmRVhIcIiW47MSD1j1LD8CnraxBQxprBZ2kxm9LCsL7NcT7WqiEzDzcuSc2yO5LrkyeYt
Qpp9/LSp06sQGvG+Rb05kHLZwABJzhIWBKFeRyWkn7HtgK/rVY5nTC6aArE3eBuh8LfBwgDaoQgo
7vvip9K8H51K3O68LtaU+0GGWRFgt5+d8KsGpZ+e9mk18ON2Df6WvFp9fCSV/1QMh/TikqOGqqjb
um3L3//D/KzJifeVS3UO41Q85QHFGpwqN/ZHDeFLh2bQG+BCL3k8ll0YlsL9sVpqK9G9EyKHc5vi
1Mk72hCMTcZKCk1dVXtCJQHMBiMgkVIqTODTnadX9SpHWhjFz7NmnYmJprhuDaT29ctuNXUhnr69
xf+woGWeFumiPiIHronUKJY/OCJMJwrhuyp74t/eqj+pHTsebMmVpvMxqEdIXYKJ8pbPM3kc+5XV
KgL0qnZ5ZNmTgI8eowH7DjDeqNrDVfRcdmhIOYqEAu7rM7ekaiePh0tr3eevG0c9kGHbJWtx0nR4
53M3613N0vkj0B4Nfrx1EBJqZsli2bk9dVBsRrP/3NZ54nRzO04HtCp1feBL8BrC9E2hIq63OnQU
jG4R2L6qN4VDSEppNSjUAZUy6fe6q4jsyvU0FQQfUdfFK4MuCghkNKPwKhduB7+RpiEHPZMBMQtT
3gIkB/lpwsn7nslyPokdKjZ65pBDYKPr6qH3VLHEtV0jM0IOPOIHxpBqTuUQVyOGsVXFm/UC4mRm
vbN3FieD3czjm9Ict0ZY4DJd2JOdOaJQtpPuAdeGcHjxo6B08HcjP9X3W7nUCK5M0qNJZyCg5aTj
TE0Yg6a/RAbt+Tu4jc7kBM2jthw/L6C3B6KRb4pZR7I+ojtdhuK2S6+u83K7/GClsr4MPTd6s+Yg
4DjyheTKLbL8URKd/GXEf+sr0jxz5+XXG7M06kPo4knRenjI8ecZsUKy3ae2pn6kXV6JlMESXQCL
eg4tj03o46xPWA5VsQGcokd4CSQ1V2bTgnhkig8Av34Eld5Z9Bl7eMEMq2eFvhjmG2efALpBVkld
MsO6dDblFOiKIw25T3tSZigsNhJ8Yp3/kvTh77q20H2gs936IVe8rML4Le3lz7GyWYnGjzmSB8uV
bQdf6USeUb4k3CWW8a9DyWGZeyIflySkzY410w342cPCnSnkyOf2+FeVeTWR1fJbwXpkggCRj1Ck
/507gOnKXuhJ3uqltAGau1Rc1EPmWPT+WYiUE1WwDz5TywYtzm92+2U9khfzF83HqdfempcmGNHP
uzMdqzCSk77nE3h40r7hvXTKO3gg0zTyHmieTHa6Tb3U1D4ygVs3TBx5ouBrYGvseEO4BmzXQ21q
TkLc53acRmbm7rqnTCPvwKqWM7PJUOK08nThGHh2LHcnGQwAPOy559VH3wC8CPGlk5PgbFMOz8ci
ezc/SICqohc++Ibo6MPRqfVHH7Pxs1nUwPAMNlBBcGuuyMrtgRsUOnTfasJndpWro5EN47x1KBcq
wyvamqqFfF6Kj4bUtdSfXEKLaqznOLmZVVoSFwuhqTUWL4JAInATO8LqIk8lA2P4Nv7UzJbBU8q0
9BbzcdgrQ8W3l7RiYyZztiK+2b1hbubPJnzFgutF4c/ZX2OAnx3yIGbHZasTLBFvyhzi/+CP13Ug
8pmZ3k8fXLg6/ApNmyU2gaK9SSMFSC9qMjxjI67v+qjZQmJrbT1Who7Yp5ou/I0XkIZdhLNFrOVI
3lyUqJ2+FVDVOcB38v6UZGK7YpvE6WR9/JbI2ere/9Aj1IT3busBx431ht1USyUK/BoBGy7yTR+l
PiFALEXvbryi/GzyyvtJd8onM7kYQ+LCda2a+uBFzqQkD6+Ivtt9QDaIJJGqxTotNpLXr1ydTov+
nGFz6PPNB9A90Itqz6quqFxdQTHLumykDIvvPgGAI7DMDIhTe7KzRt4ZoGXHuRnrK0ly4RwIw5WP
b0rmCGFEtYOUPcZX2ZmKvz54B9a4eR/6PHQEbRLMSftB4XL14QgnWp335ucIdzneJwweRW71b222
FaWjw3MXYLDFA267lr2Zhf2Kk2vql+CVh6/qyyrQ8wYAcEGn0wlAL4YdLYPzzROW6/IVnBKZL/GF
vQvhdw9yNLuOV7zkEnthAYiP0L8XHoudyQBJ0MiUqaxer/fckK5wNrG7mfDzhNWmZvpG80MhHYZP
CfQnHqOFaS6ZiZyjK8+I/foFCQUzOl9ToUrqDGqnZFcNXkI7xrNiTM3tBppj8Pn/FhO+IPuBbkLx
NYFOQFcLJQVu07DW2rhspeA2yzUC1zsR9ymAjSGTLiVAfQl3Arl17g1yiYkqgF2n95IMhvVDvJXO
FoLXuaXYEPZz5bj+mdaxWL0qxR7wOkjsy1AC1oQnTwyzF9xJafO+nduISrozZurCzaa20SYOQEUe
xlPI7Ax+WMJYiCvKFLbBhVyjq9CFX+KBOnF5QEjXQtcLiWQP8FZugvJszJxLwBqqGKDLUksRBPq+
H500lCKKrzJVJDqDc7YF5ujUmBJNLI6wHXeUCPbSW/kRrZ+F8nBXBefDiADggcWDz2wz/eGn/GX2
eZoT5nqr82TDFTnA2moC0XZZ7v4LVPVHX/uR6Q/FELgu0fx8e+5oZAvv4Z0sRVtIhEu6Iu1xDFhl
skc340984zMCVOAFwLQd0T2A/VILCJF0g0Xo7WXh1D1gbCNm4ykuNGvZ6g4ecjFG9vLtDLrMwd1G
uXzdHHe9DhVfaWqOpzUVMncSpAGy1EvZ1kLDy7h02IxxJUH0cs7l/1G4APFfk3DPS33NryUexFEB
yl1fdrOV4fAadx8XJChE3EkbaEeyRB9U/KOzaqhDK0sXEetkgPL+isVsuZTHatHEIicqKZ02OoNN
hduVF2FmTg0CqAZvUbiP+3cwp6KS8HMxcos3Sl9VCPB0Pd3KF+zrbfGpx0Qyeg74hylzR2w6GPBQ
A2dQo65mFH24WS+8sFD7Y5f8tC6cSH9z5p9mfnj7lcrTRW2rHOgEaknXRz78hbrggSS/PuzDRTgT
VvwkzbUI3YoU3bHMQ2e/1UOqBiHx8zJQcgWEAKXKyElECCbgQx+GnWAuMuzNun5ypkL2jfykY/57
y5NaNnAmuPshlbHxPuPGwSgoWmgTbXyQU+1vVA+fs6Nxo0jTCytCKNxrdriv2w81IieQbevLmTD5
0f0uu+P/39DfEMa+WPyxtXSqCuHwr39lV6KTfAAyOviZ+FSpAl0ltENHopRCmgDX6ms4JQG9w1Z/
lvFtXooJyKXbEiO/Ts8s+jSoRtubuWnYJiRnHSfTu1/WBa2JQPbjPblH6HVz5lL/dOMnUkwYEtnP
4n5GKLkHjqRMbFUV4ppt0IPcREfoUABNpBN+N6kS3ycg2ZwGEvkqndeU26YNhroUgicH87tXobdn
tGfxZaas1WTpN5qrV1FwVwQoTvYXvh/IDUKnTVtxVYHOidOufJR/mVLVk/hBG3ndQxZY+Q592Ok7
8ok1m1sXn7ywyEp9cVsrsQ1M6eiTf+uD7b7xHxntPgYkf/AJDogkV3ft2aKpHf4M3s+xOLQgMntn
+Keo2FWFhorpw6A45BRzePLxyi5jYXR/K27t43qXcf53YZMCSV/Eak/S1iT7brLllD17CR7plTuD
GPBv3uY2++jSKjhAP/soPU8Wqxotx7FmYxq9FJRuZIVZy6C1u1V+g1bGWcURIpmRrK26p/SWY0Im
zV5EeCTdZoKMAxEvnej1D3fz3ndMxA/WY9ieH9TfmSQzR4P7jw0I2eZDi4D5keWevzhRmoe6ViOC
0Eot1FYMqvaseKMS8YBl1hGCXjdPqH37bVeVY77sNFTyVAC4fIUSCxLcbgp2bkSZ3uTj+NewSFRN
3iVxfAcrj/Qe/7KSim8XnCWt43JWemhIxlV5faFbzs5/LoqAGE2/rnAvYAWi6QJWfMxLCU1805Kw
w7zSf0HjxyKaV+phm70v+AVW4qC5wrLKgV8wmE2E81dXJEYW0rtwUeOry8xYDhPnFPMASUHBhxX8
1Kjdn1bMo3M116800eZNlC1k/xoNSXt8I5ihU6eN8taa8kDwZadWcfrYvPOmCgBVb1aEUvSrrBg1
1OYAwFqw3B/50oMcXFcNKjJtqTB9jdFB7SrYYKSRyKHbZ2GmWYaL9Ugfkxyx5/nHL16PUazD3yZ7
WKoK3p7zviHBu+exYC8dKm0winZRIXHYWHP+SLSs4UVdkg5JHK+jt5pKcYl+eQHszc6QvWRJrC+i
uLvTmikGCdevxNIsRq1ra8LT3NCpK+p+mhOrjjQJYwEDMSLaWujfad1qxANdFP/Ft7y5Corqy1M5
Dq21YQYmLeKoFoMhKU53L2nFobD8JQh/snYSGmkGnk0NbxZ5DVImHll1ryeJOcP01pdjNfmOufxg
DpiU/JZcFN36dKIgRvJh+nflMZkAQAKnD7j4Hmn1Tu7PlVqtLPYvDk5xVw8YMhQTqEL1IZpoxg+f
clMqGSEzvfvOohRP3r93zAxXF1QfhMCAUS0S4Bzh/KEg3zytpYSmMQ==
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sps6dkA5WHyXDlApvW9Lm/xYIvZkKe0hBYo79frzLpKZJno/J6u885bT+1l3VS9kbVKBz70g4gvA
R/yrycGhm+a4Pcu4b9zbm15M0Gp7I+BB6HNtWdL3osnieMjwDSc5zs+J4AKACdAGob9ZusyBhP+0
N1otttRWJKG5wfoPxx3jsxORRG/da1sTH12GmDT+rV0udhfFtOzhKYFtPN6KmoEGkACCYUDtU483
7i3+wHrqNyCE8OWOfuxbKVAbezEl0VS+pI2E3hs+99QqFAWx2/xEyDabLe0vxCgVrhEteAOvoFkN
V7UbnvwLHXNNYK0lS7oWhUJppr5XZHTd2acMLw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 53376)
`protect data_block
jMw6MfVOXv2tgloUIOswPHdhYIi0eOAe5QdnC8wRVGhkCqocGTSjtkU25DCBxZD0gWbPd3It1mEM
tN3E9EtV01yoP/SrVkHsCqZ8PLhuGcvLIFPetjPMijRIlOC+LxETZNZ+7abO9/R7G0p3jE6wLtQf
ksJ9SDVftjTV7o2Umh+5+jI9+KsCUa9GAOqzGuJeIi8x+1gkVSjjUYterK1JzqRyZ6Gz/bsFyOmN
BDRL36VAJj5smhfyARuql3/9QnjGJ95UnW732Cpu80noyeTnLyWe4gDZo6cOjfH+e8b5FSGTxhuT
iKtDn2OrTiABP70kUMZiJaV93+1rRiE/0GblaP/OaV7/5BGSynAxG6lxybjaxEfQjoNboIdGAmGW
87wUH2j76yEC/KeKaWkR5NI8AW6+UA6QqJG4Q0XLPQ0fIgscwLoav0N4JQl/GwjUeowI9TUIzodW
IDcayg90V639Om7p/2gf/XzKeYD2s/x2IOAPZLL+D3SF7wiC8h8TYkFUtCBxbSGO7V+cstxJBRJo
P74+g06QPxJ5FOjGXRDfuebyR9gFCy5q+TqiFbH2vo/M97tI0R31WybtxLzIUE/3mP50iQGhmfe8
0RnWowOi4Su7mGH5GI2jg471ts4g6HYgKtfZlWaGceJqjovY6LxdMJpRMn0fiu+IVXRJZyZVmR86
0fMXMpRh2VTEmxVlEiU8BKN9aABeUDqaRKMbX8qmBIqNWJD6qtT91zWsbfdRcJ/ZVg2K7BYldX68
GHsFOtcQYrEWPlRWlm3qnK8LXCwtjOshOeWDOMXZtf4nc/TmHK1ULX5jG5vWdogtMAErDYjOwLgu
OP819Z/LrIAAxh9QMuGf3Ao0PkdEWmDgsC8K9wTmRuaJJN7IR9CMkZmYEFWtGGrj1rV3n6IyPE+0
ukTHYemp5B8/6HksqRI70znUlgVXDi/Cv8pNR56KZw3MQs9IwJt+MCeGUxLpQR6SkoutFvxud2vH
fCOgj7/o93K9RTigHyrBbFnxXZe+89WzK5g+9HcxsMiAz4vLaw3C/wZQpCgbrKdE2mNZPpUcTndU
upShZbd3MK2xY4eUZNNMy36XwtlqHnyV+Fxt6QvnQ1hg6yD1jtIfYwhLBEEDm0BjU9usdD5bQ8cG
yqCZhlJNpOctsVtac/gJXXl6jbEWkBND4CuwEzvbTfMgNiNIwCXitHJpMsZCAlFAUsmPXhaJ87bs
nz/MYoww33EgUNUWLPW14P2UGln/xvF/ayO1x/uAGrFqZEVSN5vTkJprNbzCiReYWtVqjPNh9ggr
R3tHt4r0sj+/QTXprtdVnib5OYxA5bHUSAlF0mymoFO3C8AKm8kN6Joh4dLlEdFKXVYB7EDZnY1N
HL/2XGtB9yZzVTZ1tn9nWosYqABnz/areaQlVCwEzlUvVCFHjq8+6K0GnDAwBHbbiS8sCkj8v5m/
KFZV/WrxoFMxUil5Q8+TLDg5TGhx3UDn/TFCj+4AudxoR13dLEvFEmRf0Y0LrPeSvtvPBJ4WLAUY
rBX2tztH6d0uU0FahEnWZmjz30WWFmxWzTb64lyCGl4Ka4anXPknNyPQSjdIjCSvxamEjcSit0I8
yaCbMkpiO3sctq6zisrvymr29wvvIa8ZkiOsrTdyawaAhkhEEfmeWxFUlCmaaoZ5I/Mprze5kleZ
a4gFYP+krTEt8dMtoEqWA3rQU+PLUwI8+jYoxXxXoYp/j/htYBfL9beB5OOGvBkQRQso+s8xQ8XD
S89+hL09uPo1NiHwbNcnUaiyu+OTa1U8jQchpUVZk5+2RcmYv7zuOv8EIz0I29E0OvtlpdYWFgJW
+9fyD3TrFRyUWDzwgfW+In0DC8ALNgqNGymcu3yissWv2sLsz2NKiMNbFDGK5Cy/f/XWupJVB9YB
AQX8T9BKyRwl6FsmN6z7laVnqXcesw23FWSztwAfl4ZnquI4Y3SX2qnZuXk8zvWiqRjyo3MG5pjL
ewNkPMVNk/PAs1OVzF84LtuMI3qf/0KYzxd2phsxshvA6F+3KtgabT0R2RHlngeR8KgXnXEGjC5y
TgM0hYGBDZ6BkU1XibvAc97pcU+WI2ABQE4+Ml1LR6Q81QLFmavBLLv0ArWKbBa4ab48boy+Fkkj
tZyG45x3I8J3mwpyESE+btj2JVWtszXw+dDjcLqjXNjvkv5g9ULZkDjPbdG3KDSHTZnXqdHioSEE
EY03j+djAWDyE6lC7KuHbOlAOrgtZ2Ch50StmvlEVY2xMCV2mvhsE/JGGo0P8YKr4WJZVZp/XDCU
SSwxkHpbsphJIb/WvjZUP6nswGDGZTYAZqyJsVy61mRzq57rYBgVBBEv4N6kMvDJgFt/Mgn00I4d
pra8nmlxOr6Jj07jNzOH1oU9xZy9IMpZ1lbr9ykkJPmCMUR8+ISX/yZEPBwIlRza33YUTQEFtmQl
SYl6UWYDnQ83Mutv6zBNei2ytayXPu1I7T9Z6ah57VpTjvTQTeIa1foe1W06tjrvzvgjfsoB9hqf
nyzvmOgIshUPWyfdsuN8kNk5FzmODBrAFLbtQFUxyt7a5lJlpvSONbuSXLz7AyjrmCGyGXhHxUvJ
k0jRRzc18/xyV4DC9nym4/yrLJtlh+V9MzGuqQ3yYinpxBhdM5PbS41Kf77A0MKODbZ0ONB6GAcS
vs7W71dL5ciL+dEevOXMOXLrtodNYEZkGQ5ZD7s3QExxPv90jwn0o3tDFvgl9Z0BhfGDMcdEEwqO
wQVv4r6sPqd9ckAsLWW5HcO/BTozZFD20V3I/oVpJL0ztBxO5TZTC8r0pSKa48OMeRsl25KDpQkQ
9hKEsqzDccdLREDBZiZvijHAuxMPMrXxRERlOpClgskxVCdae5wy5T7zMfAJo6khsaD9Z67Up5Zb
fN+KkJIAtj7HxZq0seYVyekMJA+8PpCtfylMOPCUyO3KW+lmMXZYqhPpVufB9ZosxQT21fHIKNhk
jva/Co/wNCod9S+ZXXUM4fhQnBpdzzvYiMlKJeTlKH5aNHDz66Zj7VbfcxxZk8behuZuA+3US4/a
kx7u53+1BegyBLjssvCqiGvvjgY6waFleu9ayHwdac0itQTjW+y95L2yfGxurkqJGTijTewkj4QU
50H99/WswjZz4gcMUWPIu0eavaNrLJpEFarU97t7yF5wP1zByMWY0sVGr+iUWHrA+blE+ldMhiS6
7O6VHf7Mqg8ekxx73Rz94+brPi5twwPB6jBwwLjxmbgwFu+MWgfvgyveHr/JwBVhw36STyITykDr
5REdx0Qnwq1zxgV4DvBFfXxOl48TrM6Ujxh0BtnKE0W3IheoDsdcuDYs4VOxCR7xwuE6Vztb6FdX
JiI58EXNXZg1EtMQdSGdCAPQzb1xegfxBDj7LEM8wGUNZjeEoCqHcxYDsOrREbfX127d02Chlfk3
idCxc4uzl7kSM/+JeLKGLTBfarAewbgT3E+sjGF4aUsGYWO0y9AE5jiKAwhLj51EDfkT1Ixnevg4
0LDY/h4AS/VAMp/7qYxRv9zkHKO6JErC5gPZKzfvuWcRSZT7sXexdLYfFc4MveLLw7qO9n51O+Ij
/7Byktnv0O8Vyw0kWej3iz0UYt+JRRCWjQIg1lSZJz5FuWazlsbVoeZLH3S4jWG8vySqYJHkTvtO
Z5ORIPBV+8IjLd6WqvY16Nj9QnQcIyuNrSuZpW2xmOl0roGpnpxFjLA7eFhzUgxfTen1aAbGOH+n
YwmnuO/jNqRHbTgVO57ccERLUE+HKtgnZmM14BvB6vfSPlhiei1LYq4VVqqCgA6PSs4fwopX+HxT
HDL86BzvkJV9ggb+tTnidmXu+6He8ygDenBR7/0jG4PnDd72/PDw1niQAD5Z+wGBuoHtzVGJe6eK
vkhND2tylhOKRSuTrTrIkJaEbblfAYi4CPyKwLxw+qstUmrUlxekYyYgZs30Dt92GRLrHENx2Qcw
9JLEWBlX3YIE+Zc5/dbye09DY2DFJ6W/F8QApZlc4VarmYxnuVJBlCr3F6uPaRh33P5SOd9y2el4
br32diySKGNvkMWWKhrBCn1CqeajqLbMeE6GxRZvJ7j1eCaKGI1/Yj8a2DZIxu3z/5EcEHuJISpz
30VC4/aEBU8JXaX15fYAfMNKKwK6FGFwfUU85N7XOQb8g7PR+XYYgBlWipobLyzxns10aFiqmYAv
LD80NgWtN0yrso3XzU47JE2a0VeVF9od37bVSAmNdgrikJdoRTMwQlvjgKAkdK+CVjMk/jrRtGgR
XNkhOiVkhyUx+tBbd5nznM2mRnEROGonIU/etvS0XU6THwwMqDZZY8jt7Wa9ekfcUO7y1fnsLk6z
2HhbzgqKj0l5vLo36M+arVk7YYOxbSsu8RWWPJIco8bc0VH0qBluSnz0+AP5vRpuuYAdVvWfGfJv
kWDph1faTivOzjj8/WZzfPJxm57lGULvpQUtEhqm9AP/Shk4asYFy1dr/bvJMRqLJSkW6tRicccC
RJ3g/QhDnD9GMZyw9UdqH5xbIrWFKVkR22SghH89s8QqtqEH9Y71+ZTA1JL83/7jhUFnHSPdElCZ
fqiJeiFT7zjE9bUHUToAuuL3HZuxX9cOAPJHoelV7dCA+ZJaknbP2+Zv2lwI0g2VoiIlsjXc5s4m
iJkNQlKZgeIkob0Rmdb1YH5V+XdeaUTV7yHaW2pov8r/NJdi3wv5EQ3/8bdJnek33axGsELFO4jH
cNj+D30oLK5KchTI2mjR4RRuWwunADRE26iW1ENMe/hpKt7hWW4jU8cKvVBATpPWgqWxguqhw3K9
oxX8ifLhqf+Ph6nETwem7THYdRl2t8Daw4EEIYCAMnb9gfYxNdIaLvZc0eJax3zAsp/ZVG1cFxxs
L8Sqppl5KVIY67u05ihvIZ0nPVhHLOXZVNBX/5SFegsYrlrT4mdgKtauma7P3XYdQ85kK5LLp/QF
O+2GanXCedn7UsSD7VO9ZDtG1ViDOrfu2gp3FgXtfy6CKd1iHunejhZafu0m86qRz2JpjLe6SKMO
lDFmwuVcPV5C7Kvk+xrTkr+aJkMP+NSU3g53a7Zw2ZykZFr/6CLzNN0SZTHBV675sVdquHjlgKw8
2ozz+eGk2lqBxQabSwmYVeBbFm6JQYphJNULZwYbqr3hWGy+I46Wsd1NvDpONvU5Mgz5MmtY5kd/
59qiaUf9Jy1KKZiPNOv01USiH+rMulhRw9VNPvP7aTgAIgN4OdVKCMoMzP8m5gqBNpzL12jyfE4z
89oGLBIMm1LNcbRPqgwi5C1d8nhJDFvQSg2CIHLT/07j1V/d99Lpe6k7bwn9UOIdcEQqslJ8lr4L
kIFRQthcOQGkHP5ERdbPKJ6yi8cJinsB1naDjMLijwNl2t7MtadttWFA68cv2pz5TXOusnLVnipf
+GKxLyBm6WlmB2B+F1+oeBrB5THcPx5s9r98x7E43HJMdHkcVK335JFWE7u6kEs0jhqZVt7jXb4E
Mc5lLvj46dxzcdfss7aEDUw1T16ZRfxZzNwhcdrR6+6W/AZ15Qhvk4a7ooqq8bCHbZktTKe5tNDe
VwE6psKpTl1GSrXGWdt+dnW/kkr9NvxpwdnfF6rOvXHFQb2fOvNJrQPfJLWkVPMJMbaDVBbSIE71
p9fkITbKtinW6JR9QgBr8KaMCRweBTOI6/7Up7hNalw/qvS208z0kM/7JCoJksON13v8v2WUtAwB
VfqnKzRx3OuwN56EUBBHhtzwRoOvE403tyalZ/t4MkTb/k7MEQSRp/N0Sw9m23XlWCVnvQKpHLbr
PV81Blm/9MryZv18W8FDOKgPad2fvYz9ZWUnvCG0aJnhDHra3666gng4jtEHBwrIX/UsJKnIXLQd
4Np7bZ/LAahrW+l8xPdE02mlhlbV81eeFGQpJfk2iJNnLxxnXT6bpcWA7+CX8RQOpmgCOOmgSIgn
Y80s95VYuYsQWlWD54TvrpE28YD965IBCYJW0SygsrMjTUJYX0uxSchpeALMdh8TXlD/BZnc/UZN
PdZuF5lMVsBR/xxdxO/zXZE7eUHeJhOtHF6Up8Wkf4fK+6oUMBnsaSQQbRQO0+Ak+RxAgM4dubM3
/8oS+pk+sx4H3fJsJqekqilInzz3Nf7oESHrvAKZvT+xcjXUfzyfphTKcz4PapQrIFAJNADf4jbH
FLHqkBkwlq0bOSJv3LJZxDWQKnoDPOpg/PY9lZ0aZY8uUKktsIyan8RKbVHJI4TGKvMaqiwVlsnL
BvJ0xgs/fRz+8VmDPuwtZX4JaMWwP9UOinEspZagD4Mjk8INY9uqcUIlyt5g0pWYpur42JKWs5p+
RgPag+biP0LoVE5QQcLp4UR5nrAqJJ1+oxNs1e3r+aKqKuv2jZ119ph+LBGZV/0Ly9COsboAqJJA
QDs07U9uoAazZX8XJlcV026LV42T/k2nEt6BCQ2NNgLc1IxCrVS6MXqD2q7uT9lit/u0AMTK6KHQ
J8+sN/hPv5O+IgkWNazJMj+CSXQxKV+BK/OR16bRUg5V8pNzR0eMTX820vlSyqm/G3c3PR5S9j3K
fL1wpHTgwvjBQBw7prJuxwROmvI0nYWzTGqjKq041b0Nw9inBuhIVlwFWUmEnhJTHwgGjzIzmMCa
MHECRiW5UhP59BBUz1qBxGcIrVMvUrc8sdsnizAnXa4pL+BBjyHNI7Q/CL9jOjexKI4jRBoaL8jh
l3xbdJpGt5HzN8CiGaUxoj5ojaFqtvyaODIk8q8Gnu3GkXL9DzhriiWWCK0kh8Hpp4Jn5SVD/U1F
uZRVRJAI+Y9BQWoh9qmzobV0oK0t/Or2klWBIfz5N0K2UthUA0pHVHsJ9r1QjXkaN2pqxMIopYdd
qVFszHyLdPg97D57FNSXv78l39HFr+1eJpsN4eM7lCeIRCokIPl2bs682CNRJiOgzyJFCK0UUElK
hLyPiR90jxzpeu7iIEEk5i7bgyTPndKNZ+6CrNHx5rRe+FDW4kHI3oQB5hh+JWZW0UPF5mnqFu3O
Zgmq5cYLfYGVqN7J/Aij28DxDqLjDUaTodVuITMN+dalLw+8Bl2YqGXOL8l3rU6l/yUYgwxi7miy
bZ0mIBSHqBMX6rgkvY4PbpmJdBHqC3yWpqGzJXnwJZyQz+fwYZQGTG+4X+PfLB3RvXqfCUSCeGZs
PLC1gRyZLwyxdFaDGvNpfjP6wwQhcd62AuLEqmgCbn98XbyJmfrkiHdQBk90+1z2KAJRub8Ne8dd
g3XCYF9FN/mH6LGf1wEPb9+AhsqMYA6Ovqlnhidhx2YPiuEE5jS6YcS2tTg4ZiTtZgzpuBV4RSZo
xqCjkEIqyhg7AWk50byMU8Wzv8FP87SKP6t4q16baemM5uXi4smpUc+heISaaXZzr7ElbL+6bFRu
T/T8StUn5ytk0havG1nDBVhTAXir+okdGubaTkDxtnBjrYK1kpC70ixpoE1DBUvKS8Gy8veqqsEA
oX6L+5+CiRsOHLOmWg/4do8+x1UZOm4fUzJgIg6W5I0lr2NgAfPeClbv4ex23fh06J6CrakNMpsG
K22TsdWSQnXHBd8T9j1Rgtbn1a5UJ4E7awDWHtTXRGS/zme0BXnKU9o0GwcNIowNqa5+5VRhC9nE
xhPl57nBvNcSxz9IV1FQMA/4bNob6Uy08rq57Bh7a+YnvtTIvINmj0xdXy2fHVNHw0bBPvFeXg22
l1AWtWbzjnhSNyuKKriMhTLtMxz/QJxAI0j1aodAly9i65yAypS7BKG7KSOax5j2bF6t7gGIX4od
q4fHG1l+UefrciSLxn2Qm2jc9aOVe+E0Boya+AoxpIjwi/zBMK0lobyMb9F1HCldraEtUfXeHQsB
4YzTctWRJH0IQIRmX6c4NMzoiFqpsYBEdywh6zNMC+hoad4u1TmRHfd6h/G9qICVcbQdn1U/K4me
ZYPOA03N+qecojGHBeFeqKCfbyyExQMriBGL5OAMRALUCgIUnOzQ882Z2zB+Bgvz61UNz9RJMkp3
hRGmXkcYDBqmQp5y4deldNdy8U2g1T4jd/CufhT4DUZWO/J9WNip/HpUSC2JDvQ2Aaa0z1F3X17K
oYXy5lBq2IwyGbUhodWdDBzlPKIi+M6P7ax/LtZy8wGOeZb01AwBRi7XlHOqYoxO5hNsTQE3oxik
fwAq0S6x4nmj7+RG0WoMYnpFDZpxVwrQXwYwB+342dtUWCG1oY7UHh0nkiUjAdHk0ey/EJpplzNL
eSdNC/zn6pJ/D04T4CgkRor+8vaQ9ke/ZAWDqibs1euOrIpfR329UCY5lG6YOVWFxGml8LSR9/VH
JcIanrfNI5297i15FCB11jwMqyyuyASUGcR3BKqbTBoAkuPkvWTW+0PIz4rJPLdqYvE1tUZTUthe
bcjDp2VOHFvCT5nEbcMQP9PgBuSdOrSIbb2minE/i7ZxPsCA0QJ0ACIu+R2fhzZuxVzGCGKw8JbC
IWHC4E25DQ+nOB5LzvggbjQihIkdq53jUYIGhzOukmNnvB9mK0qYqbqeSyp9j86zfoUbBdZRtUrk
t9XiQIvjEIokq+iZpBrD2y8+Rm1y3/yEMzvSUx47qHXYMuKwTo15tbx29Xnl5dYw5xwfRg/I3u5b
TxE0mHD/8j735oYxcvFWlQzYO8I5OCC4VrF+ZzRffYHVaOrikYNb7rK8EGRJ2i2qsuA1s109w+t6
t0dddsjEpf+mIGU0heXdJxQf/WzVsx/ZiGPw575UqwXgFIEM855FPfOuaGCqZjLSfcMTFHOUM+D9
RHZK8LSUNLybIhjt4WMQE+rZAjzW99GMD1RlS7A0xcCnQY1nBU1ByFLtN680J0MqFyD7I6hZvATU
2zEdtVfLxM6f2hK2Xfj/P1XNETcXtuICMCas01ClL3gOskwDQqjVcNvqekp7+qwb+OyjqY32cAqt
+20lIP65IBOyCJriylubq5KpGTJ690fiXAwaEDTbqUReiLfkWdEQmw3z0p83jyQH9AKEWHUpNCCc
SdHN3en82teals33ZbvI6J/7L9fg6b65LHbwVrBgnl4i0X4JMgxcRHETzYjXa4dq1bGtz/N2snTF
l9Jj2Rhu2kZJuEohCUl1/q5LVbVM0XFHpyuzKwxKwSk57bJFnpFnnK1lZVkPC6qBacdyvkp4hGSW
AjcohFcdSadrLv9Yp3sjcV73y+7NlA0JtTkNPrHgjBdnzoLIwlvUFlassF9NBJiH+o6UdiB64hQL
+ynfGbcJxIQ0sY8iZJc04/2Rlc9aXelyrpAZA5MifrFIUIdCSHIoCYg3jpCedS9DgzmH4J220shd
6aPB+LEG31dJ7TXwKknXEbUDS4Px+tQhqMm6GIO0kIU42rj3Qkm+vLUMQrXmca5egbza+W9mckuB
ng5IQ0nY4w0QIlz8KS/Pm98OerNVPtNo8W0PgVhAl4lX25lVI715vye/CmdV/ad0VFWooGFoknUG
MoGGO9yilp+fFU3tBifnycjLH0TO4bYcgtb97jdiVfoEzEQKPkmFs7hO68KnYiMgyX1ohUX4Slzl
OSVYeDsF8QPVftNrPnuXupKSArqLzHiRSXBqf3dbD6SMWd+sRVj5VUuJ8LjRWh1pJZKgR12NKsGw
Lof2nJz8aFWhKk80uMLtMI7F/ppp6TJ7z2KweBv50PP/7OTeIy/jecNNMkjHCSWtv5hXN3F4pypP
auyur3q2TpL6lkkkFndW13rPVbnHlO3+qA8fG2JU7+CXSs5GHWuLutTL/m+ii2yOMDXaa0+krtai
ZaiZ7xpLqpCf2lYtDUiy4P8rMWZnrGBQW4zaQUToJ/4mOGvwJPVNJM/qJ1xzOcLhnOJUdeSuvPhl
TnBrC2VdEKMv+FV7hfgi32ZrdNPHP1BmSG6jJli90CuLueVR2xgJLKfTjJ4m1nNDZ7nloLDkMWbp
JunRETw9cxmQVgUHGKaw2Aasj6fRh3VRgXZmqvQtyBiCAfF2f5krDoLfxNmUphsDREZuZPqps21U
LcrUd3e9m4msvtpLhW7w0jYhRj1sGEXTOW7NQDFsUfz1GlPywNeMzOmVOnIHMP1vyNmkd4Th2fo1
W8Pehjguh52tlnQ6unhSPloqcYdB0iO2lpPulhDeyIozqjTFIrFN3Iwr+fS2cq8enrRF62gNfWXO
JGfb8CyoX0r+59XKJAEDw4LZ9C5och7OFWLNGjPxfq4jP5VwbNUSoz8BW0ncULGp2k0srayU3xq5
zxHjPv7ETUugMXvCGotsya58F6n0YnvX9GITCdHtXEkUt0Q5MDSb7mfhLubwJOqNVckcg3DeplL9
8VTHyqFhZsRlkeicojD7ZJGDbdnu7R8y29r+HHQ9hybn4e/RE/53z+X4GdT+MQwtaVfUmoq+zVm2
j6icGlur07JrFMhnfONc6DMPUcTDczPmcoKzERBOgRwXr4ojta6KhcvlZ9JvSuKZIaMt94f+mjLc
bIu1lPGjeHZTm3nIa0LzAnH7o5w2l4KfW+8u1mL+V+oDwLXfD3jCnPcKlTdPu2GjJPLPvXjRi9rc
R7IqwRuhhPZdRQb69HkOFJM4mdEYWGx0QJWRahwoYpHZNgQGV4yP/iTljawqPLTSC6HU2PrwJBXC
Q8s0bB2YW2YdPoCKNFxsMtuJhfT71cqEXlmfWxFgiKIkicCacRxrCfd6H/pd6qX35RRDKOM08v8M
/1e00MxdyfUngBKDx93gnw+1GBtQsLrZAcj8KGRHlGm8Bp33JXsCOJU57VSURYx/AEw5cFcVgOJK
Sj+x8EmnJPjJIZlwsmcFD1JxFNw4rcb0BmjknYPO7bLpF6SSp7hxzbwFNT0HqO+jRZDqsb2F8mYk
RPCR8+3Gkp6JL1dCV2QIRcpM0Ic9Z/W+iShjIRbUxHURev0Hzgj/T7udlpKUcas/QzFP5TUckg7P
/eW2sjrezWJGZHXx+nlujdDXqbrWSnJYSBYo+/eoDyMbmK01IrETy0dyky1b7U0DbUE+W7urZ3vp
LyB1B9SnA9Euw48ovOWTxGbsXACG+STHzFiDjpC2UuiK8toxT78pm6l20jGs5uwKOyqbrDoN24tw
ENHkhNjZ6WtiRHR9WKm7o3D0SysTyAowpdzst+avFsPjL81ktIhjw9EKOCBslq5l0fqWHvh96lwn
76Hsx9P9FwnhoLjEds3CXee2NFI5BddzyxuamVNW+o4CE+5fdm4H+r5R6jc2qtYhOjkZRKgZGU6C
T9k7t1cmCti9gxsDLZxhosUjczIT4mNgGFcZ03+Dt1jb5Kt8S4RkMhnI/baQ+5z+rdsxGBZKCXJ3
AEovpZf1qshnjN6IxdmT1NNDhw5o3tXcD+X8CAR5peUhclevpmT4ijcAWQ2TmBLjXg24CjzapHjZ
tm7Xv2lNVy9MfHbYswfRUFZblhwiDzZMkqZB4x6ibINGm6JnndcZ8QybPBlRAYULlPaoh4AOIF0i
mkHn0S7F9U2I9Lfj59Y8KswURGPpg6oK/V2TLMQLmXsmDWqspEHAkfbylUbpnO+PcpilJYKdYonC
tHOaBPmf6rFrTVFPMda4z15qukph9iKDCvYlwkSw80BWT8/c4OGAPgMnBHrEyuG9rOqO6qhBPQup
4u8OQM1UabMTNXW6au8vxrVFa+1kQLuCJQXqulwoTL2CeiRneBHIE4+gCPOWox3LwpAqUMLZONeP
aFuWSjnYvk2hdvWhfmR1lFdHjEpOi1hvJMkL7GY//E8VRWled0GgMdjSVjJhDFh2U4FDsRupPby9
3O0vrxHBYMjq6xTG31T5mBIO9A4YFklfPpK+dIk6QxCFuhVEYz/HNfjQ9LuxWuujgtvRy+UHQEyj
M5Vh+ZzN3bJUbO5w7h1PgUWWvkH/tPSfpMzXLefGYyW4ECP6q+XZIN7Dume9ibrEixDMzgAg2EBG
EVjVhpsqxpF2Rv+sNlE8KGQ1van2J06xaVb87q5F1xYsnSk/vceK9FjqT6colVjlEQQKko0ekHKN
UfOjfl/0rOrhhAS9Se9OsESyh+6o6o7El21OEGSVRiXCAsixiyP9JzkAHBqFwRNzmmjdP3QLHzWE
68auIZj/6XsG/P/k1QGnhANvjj8CYFlHMn7sHrW6SEyH+N9WSzhS31XjaurFgpt4QM2jfyIEmKWR
PyaAp8KmDQ8RUL5UMTiMhtVSFUT25S8GyNPPYgmLKdp+XCtgd0fHR4FFP1uwKhRBvvleq/+loJ1k
+mQrNc6ZnARDtgQVnL9iOz5V67SQWIRQx1ZMIT7neN3nMpjDhDgWy3KMMbNygogavhpzxrYOHD1W
jXgc5zpvxrf9vSVPL0pWyC5zzKc/gFiIiTnJgQzjubV7cdu5hzI+dZbzzdq9gLIyUWKPuBAvMmLx
krdoFrF08m/T08cbpx4BmTUFBQcLERi5BX+D2opeN0Gsh8M5E+GMbAJjLb8LSzH2n22CL0/eoSF9
IUva4ImfZ5Wz5YY3z0xocdQPPCTV68V3FM5QwyFhXClRNoN4Ug2OyocB3hoPj5YaK78mDxa/N86r
BaCuVAuxCAJVCK2Tz925r+gHIf5Tw8USnw6j39FrPD/jXypjbNVjY9O9d9yNLOM12adQsgLwg5HT
Z/0F2zc1P36eIq/9uJSU2nOVSXl2B3Y6COqV3kfZZ+cdhqQfKd2NkFEabMYPuAJMTU9Nqa1dca0p
RA2YOEv+9nRgDiJSmFeQG6ALfTADceNcGpjDuA0kGbFjVSc5Qgb23xL2t2OGXq8Fs4E78kOEn+AX
Peg3AUIrujpBEO0wX0z/DcvBKWTkBH4T+eb7u49jgMOLcXgy2Wx4x1utEAp04U0lK1377MPW5tHV
77xOM6cMouJNfIJJUDxlYvawOi5CnrHcj9BhNDh3oVmacMBg5rvD3RpCfVBaAcjgGWv2sZTC1Scj
yRAHtDnpeHwdmjhv8xaibTwan0Hh/Lxhrl6PZWF8uIFFrm8Eeu+BdM8LVpFeKFr2spV2RX2RnTiU
ooNmR/Ini8F3H0UZiIJH3zu9rXMbX7ZslP1iPsxeMQp9pI4vAfdfRCxlh6uK2B7W9uI4h88jDvwJ
C7vO9JYUWCsTUcLtLNnBpZkfVewqW0zuGJ+sLqCelRW+TKvzi+/dAj/Tg21U3FPCMRBugo2/zOOA
vBVtPxRfClWrSLQ59ORLBD3tzKoiMU8YisV3xdYKt0HaBrXZ3UBYcBF6mepA2iF3oABE+OfB7WfF
nzaKg+cJpoor/aXWhDfZMToO0+ZcIohokn7Fj1Ms4vg/vFS05ZlkEn6Kr7Ed0ZSdTvfEPOC/+raf
2sd2f6gB+qWigbdX/vZWs8HOhgKVZshHMxR5/zEp4Mv2ULHkGH1vazrl2oKLAkgxB2AKzBoqIoVE
VVp7mv2mDCo0O7ZQ8yeyHSnan4o7arcL0zqukyb6LHGwwfLxx16WpVE6kd6YvsSYmC5CaEC1cCub
eIYkTNfkip7ej3A1VC7K3FkkT+nB5BxUXoDAsA4X9V2NFwbhdxPIYvoiBMjb2hbmMv2bPDfkf8gD
yUvDdLlo59runXN067fu3hWQDGQGJOc5osncudjaCvAQRmtWgWX4ELp+U5X+7UnDbneLGuNiQd3B
9Vn1wgMG7bcwXXYxDrARvEF+s1RMw2JwTJOU7mIABy6JluwuD7qnJdDvAC6r594CrvJy9bdQxOS2
LrOQT5Na/jTakf+qpvGFQFYIzS0YK/YemncuDOYcgq4X0olhS6nSvhMxm47RPNlWDbjwtJ0Er4Yt
L3XGVbnfb5qttfhIBFM3k0ec0XDC0aVKSJR14G8HWjf04gqds9nHYDzgSsjgLOYYI662TPgg9UGJ
U3E43dealVTO4aQ9pgWFThfHQ9+Q5JGIkmhotZ0gdDGW2IW2L76w4YH1e7hh75829FjJSBywAYbf
kZA3H/2+SRNZuxbCQaCMB8yLhhtC1nJt9alyLDB/gxJtvRAEmE/bGgISoTx90tBs9ZEhQ+qkzTI0
VHJ/ccQKuQqk/8Sn6MHvmTuA366IbBSGi1H8ZScl3n/yMte4pky86Tzk3UHmXerD84vTE5Jyhdl1
p8s9UDDFUtCo/gx2hy9wTYOV9MJi59PCn8Wko5WVkSwQWYubFhbGCM82Q0G7WiIovbTer5HOCtz9
FqUVHxmhl8enLwK2z0bTXgEBVAmREwi6j3SkxpzadKb7XUpvXDxLdd26TbM92BRRqDe5lrezaq4p
Rp8tgoozSErlu46pUPpaGuSmWyvXe9L3OEnZZEPpupeBXDvmyOTMr4IJheHA70OUJYcnv6IWyQwN
GRmX8AKS9L7ZfSNuRhsq65z/madNYwmRRNMv76IKztZjwLQhYWDoNWxUAzljY4QLdD1i8QnJ48lP
MB50ZBQy6ZXlJ0BAiAgr9OUNK0xXRR2wMmTsFAqajnVotP1Xqep4eKtNXSMceJOjNrdqKAYohqF+
ISabE7LYzBsOd+6kfcHOx8Ceyl4eToe08exLg0unxrLE6NwnlfR6dp4+603w35qKqlVKRXmBgidf
HN0EGz+ULIiGTv8zNPTChxe6Ipm4Ze4e3+PDBXBzsYgbXueQlWp/F7hbdo95Xfjq6NPHKSr3hvIB
lh4+HXQY726ijfZ+m/sms1N6W2oXyiQ3cCEuygWO3ya/SnR9RMXj/s6/iv13S+IOCANZKlCR1qtS
1lUeEiHyIJHoD7mPYTo0UrYSyF1/w0YMy1Dlic0xdxAevo7G22TtiXWmu4AyoNIe9Jh7i0T07Xoc
VXqzwlgKYH4TyPP0wnB+8zqmwpKziEASXrZnLWkFhR7kqZ/D+arrMYQONWlktgr9UgNnqHaQWgeG
1ovatG9ozgbCyhXxzZU/qwwsR0OUK66euUVXaM5BoANjL8NB5H2vANvDgElaUTjNFak1/H++PY9q
ilBIQ71SEMhydp3YN8uVVH3eupgHrLQJqp0d2fX02XvA1peal1vUiDrpTecMtcGYQsykFtnmTb7W
506q6fpfulYV+G3qoJOKN8uraQ5MsnTAnORldcDCKPNdJtxFPBXc5eUriUbcLuTU/E9OdUwU6U/D
dhl/xDWLb6hFmvwmhZ6HJE4jxQXzRvwwP1e8WUbGL8a2gVS/cRiroCWsW/EfAXMGGOibu1pZ+d2z
+G8JlATGhPLcvtg8TxSLZgzTwLHw1ujlSZkMmsEflUZnsOoFoD1XFvO4gfwfcpGV6AAqk/00aq4D
OGYezmRmOw43iaG3AmQnv/lkXhuYJ4vvEiyV4L8t4rBZ8aWgnNva+W1VyQVX8cCavB5P9jPo3Kaz
FGYM/g3hbA1NVoPRLLg4Y+gAvY5lRpGIfu8qvFuc678vUKEoaNWG9R9gIvlZCi/EqVDgQLBd4gFN
OnsPHr30XKfLALDbVvw6cA+YUdpinxwunlCOTF0zFW89e7RrzGfWAqQAOoczl2QZSEdT7ugQ+F6g
oV8M614hjn4c7cjrklWATl9s2QTuwGR7akgZ1j57+R+tfM5khHp80dUDtHwCpT5rXhttNv3h4BR3
zN1ZAw07BK3rb1dAPrPGLud0JlisjMwt3ggT/8p6R4qtvp/FE3NAE1X5tS2Gh1mVPgm1RUOIBbzY
W0czDXqfDLAM2qhiY9fUjuY5hB3OphKL/1kGI5rEZvLO27k5ftAAGaUi3CiRhJ+6H8J8re8m4me/
j5RUbyoF7RLjPryPzkQFNOfIqt+HJhXzA90BTJopwO+YB0AHEtz7qj5PKvZ0hWVsW18rSrRFQra7
TfuxfrnJDYl9sXbjfidotDCKVWida3TNlSUrsgP9Y1IiPWy0lINQNAIja5eAL40TpSc2nOmLcIyL
niLN0CJXLJlImNciFCmh3UxDoOoVlfwE4OWL2Kbingu0XAOuhei/Io95TraneDDR42Vu9MWRpzJv
L8o7XHS+35hyCYOrDnGlYn5Yw8BA1hNDuAv8ci5i7BVQY5jvDjeI7sR0J9OLkuS+q2eXi+yzhdhe
x0l2/Lv2NU+IkkCIAKwNYL3mweptUJXEXojf6rg5G2pY+Hu/3CL6S/lXWJt7+sjGODgrMAsWGfbA
sghJTHESWZtm2AtxkVDzO51b3I05j7Jm6fYAfJiNrKQtxQR7Z24Cp3xCP6jDwygTLpSXNcdhL5Wj
TeJvA1LAZToxaLtBdqBCxjkmZLFZzkUNn1KSJIX3+0pRVu+TAdchxoJCF+CoGPavoNM8VkyDthl9
JXUm0StrBgUVbUHFFu/EiKH0wtzLWRaZEVa27UTDjt+mdubpy30lx825Dr3xrhHiRBfM5Ri2tWQA
D/vonSdM/rVmqk0Nk74UG3aB3pqQ7KOFhHdLhNdAdbk4GhKexISVwUvvDgDxdZpZFULc1iBjkVo+
ZwRuKQa9rjt9Ru6QtWdtcq9sdE1eYhclZ099hyT9M9BDOHqM9Hc1F1NK2G/2ob8IGXngTfliOWts
d9xcCkkn25+b7q3+QAg04mbd3JZzFmMd6ObZLSdyzBo71CkC7sDx1GzyOs2/VsufFSPhqfjOW8eJ
uF/p1Evy7Uzz+7AisSjoQ2SZJqR/RoqAi/nf3+mKm4etMsD6moX6Xg8AdQsKfI+8jAUqvGT9/SP8
wtIXrctX37lNRQ/hGus0BSWa5+3TBzhZ2P6CDFagIzOUx3pHx8HA/FFQg4iHLhnGbbU2Ou8aHG2/
FC/kF/iNe0TE10AOQThyIehsrSZ83zXKFOAIG/yGeiYluQg9WBrWsRryKtExRhSg5JaP+A5tvoiN
OFmQq/P271DF6N2W2sG7gfWdfX5aKYzl1P5DOf6zL+U0qjWF0I1E8bqNz8/Rnejwb+OG/rEiZm0F
Rm3rq4mdOiBkwhVIMaFhjMA7QLWOPUleWWaKqh8tiCTewOJ309U/J+10XWt38vqXwzK/+yt3/d0t
nIikcB7WGzzWeMyoaQ3AFTmXlW20nOPbeDnZOoJARnQrI8JZOK49u2THzzw3YOBISTvLhIWXq0z5
rqyLif9dI6W+wsive2o9Xrjvz8Gdta7T67ayyk4bVCs61Ytow3o2v0kX2QHIlXHo6AOcECq1VmF6
aNgVidKLsb/fYmRhcPVY8rhyJHFWofPyyajslWNhyflhSO4c7LDStwt9LwuMKXvMysVY17MzbIkO
Zu8Vd/joBj08qS7jNzSVqGGfYk/Ox0iD7GwatUrbR4GQfs/HYS3DXQZFjipLqNauop/r4gHBL6ds
0IlUsjxhLgmZznOAD61BW1unUJ5e7+Ir/Z6PNJuCo2bcdlTbUDWfz7uKKT9aUZDHemI+KTf6QQIp
Ng5IrRFrFfTui1MY1vElXDo0XkcRj07Myt/Y4plXUdk3KRaNs6Gu6okiwc5Sf4nrQ5pcEITTZYrb
hK9Mo5mBCpY3PlaXA0uAmn4vAPEm7Fh9X/ZkbHMsKz3cSCAnk8sKUohpaSTzTbRI8AUWAxfjvAeI
/Lfts4ozQsCI8hEZ15ZatusiBFhQBRCok+TQz7lY3mWgujdEujwaewBHjk5QDMAbksMGNn6PEG+9
Xevg38fWsxk77tQ3vzUoHdfrtFFIytlOyM+8394p6Xez6R1lBj6kEWFE6KXrzpMIiJ++CJxLw36T
0+UtLgQkwqzd7wzKsj/6v12fob5jDsBRO2lMmXNxgnzRoyBgbsXnnbdvRcCaXdR7Imyup/QFkjn/
YyhylGrvhBHIj4lt5Ax379uGKT2GW6B5xhUyyCw+y/YcCvEg4US4YWwiYHxzmgtthkaV3rYHGJN1
bP4xYWNkWQgYLSSQhdpkUXzrKaIWgqulechSsrHsOAu2Wj1Ej+k+L6zMFjsdTrZ3LDqC5TssEkOr
YDcScptohm1cFa+w9jiYQ7aAYWW3xzY945CwwZkG9V6VphHRmdo0G0n26Llah5h9BO/sN98/y5Rz
aizW6dAvLStXAep+EXeKWJlX6LUWsceMjV1NR6jMEkdT70o7WWd6tDAe4RTa2Kq5w4McS8+IGDLx
oSWISc9Er6dQ+XO4yTG3wcTNaIvzZsLHIB8QOPEqBiA42jq2qddJAuwXqwZhDc42R3UatJP4TmEX
jfgmrm3lg+eeYuu443gFKPwG3q4vyKQniiDga7ajyCccvnXgoZfipzXf6UAa3RK/J9CnaowYVuV1
zPAYkPhIBpeUEoi6yJ+ckNlTX/hTr821ucSkLaVVB1T3AFc0HpMyd+QhjK9uJAawsJSQWy3FMMpR
fV96sud0JR9khOHtzRH7ANUm+nxuheQ7gTaSWkUAeJv0X+x4GTlDPtR0uAOsIYuiVANvYMnmmQLO
AvTSnbltJt8Q/CfPHmsBE0FTM1QOsbvJ6urj+vx07d8fJGV8yaZpH7zHScpMLgVq2o05rGYkhKr8
dcPTWCJ82RwzfBlnd0lblVJxsIsm1ZpeaynBxullRsnagplVEZsbZhM+I09ktGxyB8cleI2py1k+
oNQ603wKkLJRU/zEA2p2M5HYviMUb+F4Mqy4urMVvXyT6vxv5qz1YMeN9JbIvBtAi4fxGymjzSEJ
6f6h6Uj3J6f+mCiTz7zL3WSEQkB525hMhbfBB7bEUcKgcmOEkIyhilUSYHSKPfIROJ+x1NBDu/og
9XUPdRwBy3tWQW76ddItFrhBmBBWSJg0INeEcUyPUOHZ5ipNOEVojD+YMjTkcvVKOYOjMAOSKYRK
nMPBMTAA50cl2xtzmp2C3lCIXfqF4GVkWOWkxmCC78p0S+W0XcPNN6IA52nUruTMetThRJtCOM3R
0nTq5w5FewUTrNf+WL14ILtqGfh/18BYmIGhxHSVwR9hdHbBjHMwOTmPbWJYi9NH5Gk8EJfkLq5N
TUcubfvbPCuNEpalb+tJ1YXuO5UJY8Y0+w+JXn31OpcUXkr0TfW+00UCX0nPTF4uK+bBZhiqbeiD
npEJ6sY0DG8bH8zxlZuCEPOWIQmtBhEL2g1SxmspHj0q/7zb/08SNlI1dVvnPDFM7JOUMTtmKwTL
TYKLStRoOSxIaJDL8SwQbIi4PyJ+YNd5S6rMG25HB8oOpZz0DVlDZ/5duHzBCQc3NyhL9COpoBdb
KaaphweY0Jp4Dy2qbZb5F4P8RcPznf8HCHevhY5kQrpPz6N6REvmYSZtJlpevxRLRykarvInh9Dk
l4PzvBP4Hsc20XYrAAea40pkUIbPF16j58ohDSyFF7tkbUN4xcz4NQvcZDGzMhLa6wtVb5sFQJ8m
nyNbSgPU8z/eBy2lgBIUjIFs3Xca5IYDemY7JNNFb4BLOAGydS1D4tgmUI7FNFa89fiF++skLT1Q
OMKa8wgme1nyQ6hXqueZcFMwNGF0DPK3Jq55ueq8yG7x83Byf6RKOUu8T+4OzWloU0VGcRuTgFum
6QcG4kXGUcc4OJWfNWSGvqh74sKhKu+YbHlnyfOe+SH8wiNYrvM7FeeJ8abaDcBR5cBmZ4Zr4WOh
OsT2jubdPnZP4O8sxyn76YvojFeP0kwNw0Rb3+iaE1CQAjMLa1xdVnyCiU19tAUke/KGgbkxnXmk
xO4IcRTgn6ZjP4+4Y4Hor+ewZRDaQ0E8J0HA02oxlONM+wriVvRpWgd5AhYWAyHuu9yWEbNc4C4w
7f9jECCrxgF61YcYxog9beaj5B7cZqxDrnhgrBxhD4fvuh0g3QxiGmcQ//pg3X71wysdoAJPy+15
2raVdJFiw86TUhxmmCO6ULRchX9lsMHrHTSdB3kMbalXIKlhDBBybZAw+TJ4sO89D4dGmRKqEd3n
DUNqQP08nBhHerGUBFmNzPIV8Mvs4P+sQ5ip7AMzPfke0QmjBqkAAvrtZthZlBLeCPHNP7mCdmqy
ujeSqhzOfBnzv60+ul6XkbTOPJeZ3smRVQW/r3ESKNNV3CFte86GLuBuVoHjSVgCD4LS61UoTIiz
z8kQSjY9OlyqOFApKw1sIQoAc9Lm5bduOoNJ9gYojF3Kk3TuJxmx0GAFHL45AdUkxoJhOybh3Vy+
cthLU12LfqatpGMXy3qfgzO0/EZN++yvcPFnk3yP1Fmvwj5UUAZ8sHidUDnTpKdD181vVgNv5vOu
PDDD9X41wBi7rICwtBg4sTWedEq59r3ZnK90he08FnMIJcDYYcIy2h/C4cb/DfSrc1mk/0Nq4T/w
rED+4ixsZhGr9r178rprxht90pHMUBIfIFv9l3jVcGyMnwnN7ZRmZoFd6XXmPrYWgIPRfJc986EG
tC/Bw3ZGwKO5uyBNQdSGtVIQ2cCul8hE8c8v6QolahhPY5Sf0fAo3++L5tvDvVnx+LCBvit+jQ/D
neturC3Cmsm0vri2BKNVT2GUnEiELvmG9OiYTu4WF9BaghC3ZIzaXKXY973mE1V5KyfEQErT30ep
ao4XuITdFsnJrxtFSBf9gdzLu9xqyXceA4rxKL9csWzMUezx4YpMH5RNOnJ3yrvDkmf44o31Bol5
//JXccjdO7sArl5g+Lv2cctGhkeKLUYdnrywK9sS3ELEJa7wVUwFSVzXvxctaD9sziKpxawIsgAt
YeCt1ldMSYa0aKPkzKW/NxTvRo/vypSW3sPC58JFLba8K/jG/BfhQ09n9/ria5K55yV3WxFY3mdT
Ct9+kqoVCB+m1gz7ytocK5xpahQVcCKeVJEx64mry/ei5tc1aZCF44gsb+hbkGsDEhD9j41VS6/S
LwIjiVRgteJx3SO9Ket4DnUsozP9LJ2MhEqIPHk1oLjhN7WSjo3TGX3x+gEnmVMmxvODCUH77t5J
iIKUwYsk3hDtkcLuNxYLzY4t94jh8PaZBdbv76zvde4kyJOKmcV6vFyAPf6K64Cai6zqNTz7ZJFT
7KhAhvWDO2p8XTAwtrS7Yj2xZ70GsAM9yIojZBkw6nvkpr/wgFRj7/MyO4vVgsB/pkrs1v9A74k/
i6YYKqBNa2aUOzReg0KAPo7aZ5JGccdWGJCXqrU66klucp4cVTwGxhkxAOhwlTv6bDkR1oI8bpez
uS/y0X4Vsyko5y2gqDX6yYotCSfGr4xahKh77czZDWEDOQ4GfHhBKPTag1rZ7AJJYn0YdUmUzlkj
seAiYWeqghnMdPb4t1WM2JKZi+POB5cQI9mbGyNEaA/RY2m8aIdPyD5yLg3QiC2wbZ/JnMbfWT0Q
m3q7jL6TnzkzYjLrdiZWHvmZxiHG6+5fE4oy7g5fFvhxxHyTKb91GwO4kuJ9PlbZguTZnV7Hs2G9
8XjYkjShj98QI1R7nBIqMVbOcVTsQGXo9RgciCUSVBT5VfFrfa+zVyy008no+jL+luqoATBCLfju
MywjATcdfmGi6v3XJgNEYZG3fjh7RirD1hDk/dxGQB7n0zYpC+tZx4SvMHh69vaAidOHwH3nXUx2
XWpnWWkCt4pwE06xvGoKUnCVT6tpuigU34+NvrfwkbwK64Lb+ZtEprcPqEDgHILshP+z7dgj/b9U
zwEiWKJdPrdB0lAtH0bCSmTmgt5LOUPPGwIsDt/NQbuJRoCl0rOr6QjKaj/EFnanAObJB1ikzxVL
m7FZCRygbif0wq1EoahUQNStXSUNq/HjeGHT5Ci+iy+cNpoWu6nURSMurgfW4S9uEyIvtNDY6npA
lAQI/9rhz4Fbz6li2TuNsPIku9SBQEKSpBU2G0c2ShS7JO2brHzCXcqHjWUH9QPjT5Q2ox1V1b09
x0a7V7hHJS/xzwfOzojjRCyhVwDEwpIbGF5hGKpDUAeFRKb3R39fqyvZmoWWz8g6hej4BbkEfWkj
N6AkEDA+MX09PDjAY4V3X3hIqFWb1BySt2La4YCPBInnqL0mZCMLhBeAveKWufy3BKKRaMJdBxXb
Pd6XVBpsgJJMemkp0GD7dDOlPl58pLPiqXEw605xESOUc7BamVCDVyi55i++HuCBSLju1xkRIjnH
MBE3PMmYVceK0+NX/5dG6M/4LJiyz9QRIjgdp5S12XK/VMkd2AyldVSkTnhJ960jfnYN/apo+fdW
kWm9IHy1/XtGvaF+9EckHqSTudMsyofNdaGOpMl4vFpgMnqW6ziK+ezudeiA7/QSXo7sJDpGMuEE
EGkSAXJDHQ6nzWQm0yQC0oo994kW858Ul+lJOjBrU0jcvK/s9zIz35ujak+jwG7QpEO6jRO89p42
g4wv62jHlmZ3qIY7STxpobg4n27Pdfm7EsHyZgMxH/gRdKFjf0Nr1V4lkdLvm/kmq6TJYn4kJR6F
hhsM6EgkHlNvC9v+lubkmWX6BGYpHMSMH41QrF9WRCyVeSoAuB/WxbN8BFfeW2RMQ7ratFMnrYLe
xLo5gswQgqee/25s3DJ/Rl1Pd3MW2t+zh9fG7ap1b7r+vvRVz7hu+xEEbZ7GjvywQUs3J6RHJk0P
w6WY9kmilEiNNIhT6mE8T5l7RphVENZCAPdGAT2kyt6cPlfUMXSHs+CieVJo9544pt3uhXh0x2tu
wBFecYB9mZLKOc+VY1TsOqSn76G8R02crdWxb3uph7o15+skjKJLVPnQcuvHhOdLojAWyeFZ9Gfn
zY4/23ap0G8Jj6cn9w+yH7TZytdeL069t0INVyoARwh/i/wGmvJ8+hPC9uXEoAZfSWxNlLjZaYW7
qS6O6PVVaYcGRX2y6N7iHNAAZWd3pr7VmUTbmDAg9OOJyHA8yPG2AyKlr4tUve/6kgNQ9Fd22Bki
1Ljj8zHa7SF33MKRHays9eC7ynJeotqj7+XGdRlbPsVWQ+uo8D09NEKrNI22kuaF0aj0do1+gvVj
9byRUMGoVjGhuUiIJX9RZtRZg/rx1sEdTXvsB7csiS3HwDKpBV5pm9JJpNY5Av073xQOenzA56Yl
QLb+pXTzAaDsXgHYn5eZCqT90qpBtzMnQdpfHhLLuIKPNqD7hct2DSebLzRt5dHfpSwvQ0uTqfDh
MMFMIn/CRuZaxVTSf9eurq2XDJ+sopvjzRWkkLQlU37+ZHfAM4SVPk1KugdlW3UHBwfbbwyQzPoA
ITIMPraAUMSWFkDErEJEYHTaJjeGUQKL8gUq6QB+yORsquBuHqoNQDuZaZ0UxFWAGhfkbH5Q9tYQ
rzQvaZmRTOe8G2kFGCRJdZAwOHtXi+KTzf7LkrsxFrqsFzKtKRlomRuKCvGdYE02nAn4K0sf82be
RmPm3EmxvBbCn71SSSZzvtohWLfQbuDCcHudnfCHpBvOlprOKgO5i8rL33lNO4rL8mV3IQCGngNv
edV7VwySnfKClgy6MtGjoV3UZOHDjX864hHhVJ5goBLuFmnDMH5r49PcAi3+3kZWt8B3ycAU3ab2
lEvTfnmZO7BgBL0JJHrN7NOTw0Q23gv8vacUN71QLTgs8jl2OYXf/e07uqR9MDUJu/8jfPioP5PU
5ewsfA81RPonZyGrG+lCoVDpkIkjzsXwbKiKpRPok5QZ+d/mBFgVTXbytmagiOA0N5QXM0+o3Q2E
lZgKjSH26G3p2XOFlB+aSwu5xbuzk9lWhqg61ZtdoNlArC/BngsP6MAxfBkAKncY/E7wcvaew3M0
xdD/LpeUg25MSIxufnld2Nn00TElWp3Jcq6KY5Eq/ZvQiXkq9wzRQ+xv9w1osKz7Vv5mJ2nHuKJG
jI3FVyJGddxq8fxnKlEAhyxFI5CvSt+TOfDY3tnU+YCDsYZTDWDhH4h4d6lPQqfnW+J0FbcYxfQF
PuUgKmgeslx9GftZycnf3pYvZjG6A04xAiPH8X2as+igba1wcQLPjRUJi//trKQ3eESy6WpRE5PH
G5gVyRfsQwMrnnzwbFSU1NWfWP/aEAARJmi2A1upzqwY2N1gXqdzTNPXdMLFGqtGaqs/462OXZqf
rUYkC0EEiyvAXdLHxLGt/q9CIobitC+Mv18zPum24qVKe2XoIyeeIGaKH/86y4n1ZNKPXU1FBgMq
XA0d6Dq9CUeFegzUT/J1nLt/ux0dc5I6/Eryd3SW4/fRFuvfVHsIJh8NWaNQdAL9GQT+/PdP3lc4
frAlF7J9IU9KXLRcK3YkgqymhaGKctW2fOf2eGzhNAyZfh7frM7013wPC0l5WE0JjHmwXbj4OjRu
z0UcyHfmzTpE7G27sZBCx/hJqMxixeho+9LyukQK6Te8ihwyEC6Q2L+MnLs/uBmLWIvpft03weoj
JyfVsv91Vzq4TOS70zRr8EWdxUe0Ny22XtAMEm3nMGR6tujZR+rr5JWeHG118EpEt2wKGHKEfKkj
wii/1EaOopVwGFMhNnbwzurJ4+nNDXSZG0vJHTjqeTJW0mho2SDpmTV/M3KPl34icoTB0YtQjCqE
J0I6SaH23d7vd7xtIZePLBOzuLfxv9xeN30XPYPerSeGT4F9W1TjtZmOph+7g3hcM0dTj6LUDfd7
JsThtoC/dt3C0SGV/pc5iCUgvSmgQmWClNcoejWKiSpXNAbgvM58vC+1Z4Nz0tTbP2xv7PzKNKDk
L6mmSxJwcgUsFQ8TAhgeOPJe+CRY7oKk0UxavRH/jDtLkDk5L54GC61oBeggemmzh8GW2H745HYG
PxO4JaKWPI4HtgYHEDG0UqWpEVXvCfDG7PExZtjgw5OH1qX1jJsx7gCaoBP0wqVZTKq/Gr/Nxj8R
d/26H4dZgI8gRtoPHXdYqDJg8xkKqlGvJyE9d0ax1yE3+D6/pX7ZhSO79yMb+6EAR9e2rTPCAyw7
cZ2Z2uTDSbDXhoTXtm8h7JwwmeOaksW1fkGKNwFeWlaaaDLM2BS6CwsljYya3HGsyePXejzUZzdL
YFvtolgc7RqOZR5aGULbnTtufyKwT5oIYmdIA2xocwnLIsJAWroWJ8BpJ8runC9nxUKmNYda92LE
kyx5YdIkh/0cUc8Cr8fvsvUHYvFOfExDScP7bQ43KrhM1sfIi+cOGIr70EVpUsRSmkyaQn8A3yiL
Ar5tZ/QYc4G+ktz3C1PVVR/ZlBjDiSFTSTPG3y80OlVZ1X5jrQJyoOZC/ZmW2wnAe7QqgjVOYsGR
6gwyN1UTxy1WJ/CjXCtYM4t33qHV+wczZomqe5gV0Pp6Onm2aVUDVTvxXGf5WJ2gEb91P1nGyp7g
CTtdTCLaPZ+61IWgLpWJqU9nckMmwS3EPiBSafp3AGHIH3UEsmgU4/rYFyCYCQO1E9L1an/Ux0hv
9cmedzfN0s6HVU8p0tsXC+FBqe7H4rcQ5peK7N4LJl8uCs4RHmU7Wu25iLTCI7jj3iKDx1dO0v3x
51ee3uxhCKj7fB+o9wSrl38VXNKlAmV+A5MnsIfucdvaSqvB8SkPIPTM0sKQI83ibbyzsc6K1Nz6
D7SfJkgpiI2vGQxrZryBO6EFpfFEE1VLRkNBZCsTS4hv2WLkY0BZlDUK2s8R48aC+KKjNTP+DUbC
EjwYx3CcaclQuVvlKBFjPtv7K1uFY92cqpJY7cVquPR2OEd/OeyxEx/0bfjZ1fdSjp6dlKtOWwWf
EumfhAnsqDDM/cjwmfVscr7wDiZbtZD8ysUttta3fOsPPxxU0lOlpuKmkhvXzrGT9hA3wC30D+Rc
f+JTCi1qxzA2AhoSyXS5ZXBlLBt7PK0vjA2ORNHwjm7NGWZNw2/AZTBFKj2/YsknsMYVjxfPtMtl
bhoQGaKbQo7HrSxtD2pB35VBxjke+PpsMTJei2x7/p//mWP/cCqUfJHBd9LPymGa3mXq+p44cYGR
KifkG8MKcBzRQpc5pHreLC5neuG1O7bYV+AmGW+IUGM+DXW/jEptdCbv/F22MOQ8ov3Bf0NGHMGj
fvHfNIOiPd35ZPlZe+6p+HtTwZe0ouGZGw3DTkzCO1SUmOlKEhaOLM5inNzUzZr7KsvkrVeYPuqa
d54zGbwT3XRj+IpXV5Yr3usCmLHWhz4WvPleQhZUT++PLC1CjcNswcLiixo1jLl5D4W0XFHRVLha
6Ms9ZOa5Uheco2Sv80LK14eB4hTt6M1Lia7iru0BgRyTmsZugWfBuXhRqbMQJGSCdrSJGhu2B3Rx
Lxrgmd5hO1s8IiscEvn3xCLheKR2p9X9/egnI8zr1qGyJOYcsmN06kVU1/VKe9UHofhmuHRF9elN
RNIQHR8MepF2wgBoeyj5dkwgO8rzVboPvufbkxs62wjbMcqxwjSmVtPUGGpcViZ1joMrae64W8fH
RtN50g15Lh6DvKr0Yq3Pb0dAQ8Gld6jJnjeYNKID21d9ElgGH8lKoqUj7K6qvPLaQO5F+YSk4I1G
cNPoVsjHZRqEcAkpoNIktzwLAxWa1MyAsFGEQVITSmOmtu4kocog2sYyyqH1E3Dj6eiDfvCjuv92
kBQ5LkzVLkyjfYXB6Bf98YkwxxtIDNC9xpGi5u7451umcjZsmChb4ioB3/wFJCf5xhjJuRv+ByZ/
10iwpf6UjnHpjqma//ik9tCH+Cstz3INHTXtVWaU9T3Nly36hN0BTawuHOEnFiRmrYSsBGzx69vQ
V7Kd/QQ8jLh189BlGEFyIBRROBFZy6UoguJ003Dg2yEQduFXQ5V764IJN+u1rPUspC4weeguin8w
glbAnygTjGInBBPt5p4C/0pKweJNfn7JfbpNNU0AD7XYDbjBkulyg+L50ZVdufZUSaLmP0Lt/M4X
35+6ekhG2Xr43mkt0y0D82WkRBvV7I5uWgVyh5TWotEdsyiOFAkgdWZTVGDvjFT3/tiKNO6r7wfV
DuDMT4CKVUfqkgnbPi2wxAJ0x6J/9jsfsL7KAYbIr9Au/HK2D7yX2DGvlgdwrFBR8uKjLIRsIC93
Ihq1LfH2uh6evY6lpgPkYsR/k+YyYoXG+1LAKDFSOzvdvW8+jqFaAcGUSOXODaDEM9Oh0Hsbx7du
szRqX7AGORqfvdMetXQ+ww13PisVRORdgDKyZxDKLlZUCUjtM1jGiASxLd/13a9zj5/GedBl5EvF
qS/FNqYXMyNQUGSztaOeM1WV9pPHgLS/BokiU0AJfCHytOHM83G2q6ch5GpqT15NGf3Epx4zLAlR
7ZOlcIvyO6daXcQoxjcBYhqm2I6pCiQ2uvHEfOSxF1NmXBFC7xXmap/3O2drUftgRTD1gh3LKIkB
iOdsi5nAH7+Goo6nmntyiO6olF+EQMk2QpWSWrQKu8QMd7Zwtv+HfJ6jMDPjN5U1RQwWHVq5OCnB
xXYcFFu3MWCWkh1EkQdAFpgRmyd4Hi4BQLYoSR3ci+cx3qgCE5FBV3g78GUAIChkRsuCM2CbfMEc
+8Bx1uP/9NDp+X8og8z1RgNaepYawnCVFF4r3LKuYLzlqp1KbFJN5A0j7F2wa4LHcAyv1TpDjXaD
SKYmii8RCBmXNB0HyhijUjepMdIOpJXqFks9PbqRY7JJ+TphjP/jkP8bSdtNG5gNGn1IlDfR8fpP
u/MbH2wyM0M8O1crekqfA2Rd31vBvJNdQWMTjWQS8mmRFwsXFln0ajapXkEfOgJYOyH6MSkGUPNG
PelpTtx5MaPcmfzASQLocHqu1kDQn8MxwqDgMQvymhci02e3tTdbHzeMTjt5+jScRUofKpsWuAaN
BUlL2uoEAFK850+v+Z1EXfn12wnwzwDRPrx8aTSkomn2GWbgbXiPvXAM2MF/49123dxgY1TEdKr2
gFP/eBhBWaqbFdE62Y7sePxUbFhWVT5NNbuIYaYen4CdE0Czrh5QpFtgSyECfoSiN/MCuUT4QCj2
Ht2ElG02X/BFRgUQoGdHl2aBVF9hhu1drsHd/24CWOyGoXHIetbVo7xD7g0/zp7H9waGI8zYTPyW
im0NMiWFF9xKhPl3WQxTi4X7aWfF/mJ5a0P2WVcjrIFcmrZSXDgeaNe9EhmsPNam08cOwGM2NT8A
VjOFESXUEiQ24VtaY+QpjFOwpLWUmKRSrvbO6Edl2HOUzP2skWFMIY/Bk+W7yfxIeG1cjZdFZk1k
3AOBnaYEDu1AVPWC5NsjdmRbauieS5HMS4UlSSvEZHIkuawA+pJ2DKDvf/cb3OvxAI+PLfn4A2fv
9NcTM3WSYHx7yFNlNK7IvwEc0HhovRffl3fNU+64lJO0YGCzT/9SwNcp7QcQw/2T0hnk+BCxeqPJ
0UBZoRtS/bCOhKEfYe7AaQWTZuM+RT/pf64aIC8nf4HHPrI2N3p8KAhqGPM1pg1/m+hiJzYrapke
paJJj2Sg3J0Y9SMT6M9NqguLpoCOfP6Wt+VXxDP4Ar/RGETb9egLIlAC80eXAmHgU4TYWfz71Lb6
tvKFX8lyrw1sLkiFTi4BUmifD3sB3ApGAw94BtctstzLpmLe4E8PTjA05pN/TUiOKaBqlet1qQGR
dduKqbN8HPEehCfNFYVBJ4um5CeEIRMO1ZNGTFp/c/sKDd8JXG4IAlDNVWsqu2+vh8P2feYlCetM
ug+1iw87F0XVkuFVPggRywvBUHPwcFU5ujgSG5IbQaHlIzn3sl7zS/tkE9hk/A0IZqHU0pOYWrY3
Vdg+2nZYXl8zT8RGM6OyVjSgOMwgWXrw255sTjcC3MrIF6k+8UffswYsse/CkP46ylp0S2sT2PHm
T6uOfR21m+Ao2VTqHuxjbAeSH0Ss7JkbqdPTw/bj2OezbJRPe/DMHW0bBdlClUi/b1u/xVfYOdBs
Qhl+C/IAlPtDu/KTf4q29hnPwEOBu7Tv8N39EOTVcCwA0m/SwiK1eA+dOxcGT1InExywGTv09Cja
5HLm3Kk0YsZqVAeJahqeBJeqcn56wdZEBhzjrvNf4iXzbB7HTz/0XnwLMcEtt3Q0Sh5JZ3MGNdY9
o18UVBQ96f7sD8tkySc9QDlu3oOPtVXkB8fMkec6aUA64btB3xhSI8gsFGbvlYkJiPIPF3cjeAt9
M71kClGUiJGaz6/3RRLlhTVl/cCle95Uz/rnma+WBaGnjpiyeW7LxRo1OzF7DYluNrrAFRziXjrK
KC3ThZASelXn5TjWLly4WNjiWLw9WEoeHZdLUGfEuq2EBVxQ1wOZllu5+FKkqn12i3KuYhReUio3
3c4iF8/08VAW6BXqBapfGsWqU87ToaSntoyGg6/LDY7er4+X6yGzw7H1jNWSiWToZtUWgkExtFrd
eChNYCzBC49B5NTiavlJQhH7PhldwKILtpa24dIsk/F+TK325tugQDZAXEDqc5e4QTS+Hk3xCqW/
T8088N/LT1FtQyqp6/A51tN5Axck2D3LAYM90blahhyjkcrbuOJ6eRDR0nQub6Iiz5ZP8HepXkk5
ppNsa5HezGoRAEEIBNDW0L94ObbhrXVKcF7b/NM/nMXESMV95GRU/nD8glnPle9b8LohB4c8O9cD
Wt2pKbB9Kj4k2OVfg75Q0JyPsKgtJ+cu38pI6xKaT2bZRVr5D+3ttNqNalesFpXD0syGsU6CeBwL
VupASv1nG3Qb2Ga8lojtsnTFQVduDrNelbfxYTP7RTUVau3bJD3KrXPYH0/b95OLpVbr8WR7ODOg
hnqr22c8gu6JO1+C5OujRXlDPoqmQWtrQqqdHRQ8jFOu5KjCDoxhMDAnFM9pKC2cceT+jMPqgiWB
C6g7KAGmZh+ILaUR6J2ceMYaNYZQks6RUgaktScm6497VgX+3Kk1U6mVinzRaflPRozLHE+YqlqY
S1JGvJqZ4p3znPRg2W591JL283YzMKqxir0d58/UvlyDGKDM0A+6UX2yNnyLdnM4S0WouPE4pLez
jazbtEDfzAgsyJgM/Te7BdeQLUUmILlEXsNwjA2nhuZdJZG9mkBvwC3hGXgcCCB0ucCZaqCDwQUX
FO7gICsCjP1Y9LSAifFkeJB67toiD2/EWFl0I0lUenB2aPGRYk4Rdp4IvnxQ2nraosYB3S5kZ+dJ
b7ziRq+ThOCMn/1QgoeVrUAhJUQTm8FpxqNENm8VPZuLvbPsTruyuuY6AGg4jrFCsoS7p3pJcGPK
PZ9WR1WJQD+/sz5MvI+1D5+K9inD9UVd5nqmNKCNLQOo4OmkoVZANvD1G/pyQ16bvdc0o/1voCSu
HpZNA86ZcNKVW6+omuYpygzgsn/Va5KRz94b4434GacUCVX9tiG3o/MBu92qHHzj/N3GS78clmBO
IOG4LKQIia6WSWn5/+q0RjMp9ve2yAR6CPZbMHMXdqvalxunqwY9aCuiUCTICPqwJpczaCldQ9rv
zeaxt0NAKCLR5egSLxO8lMKvgksD9wW9vIgy1Ir4JgNk/rGk7KD+fzubpC1j+BBPftWCyrKWlYvz
QIxxHDoKXSaFsM4pIiYSgoJR+Pr4FGce46P+9bBDWCkTQ4ASY2SdMMQ4mR+XvO79CTT8h8YMiYHj
6/5C5zMSFIKpolu24J2elJ+N/FFwjpz8KKC917i5fNqSDWwQ0JXbwTo64Y2y1X152hT81vVvOG3D
Ps92d6D3TbVxCwCFo6j0XAufvdXistS2QUUcExtbcSKoumCUzlAq757yt2HfFMOvvK8awjMsl5F3
SEc0HPMCYPC1ikJKyg30iIcezRN9p+wEvUJ7thCBHrvsxd7S6GMe+G3cnHW5dMPvtq32PgXS8UWy
40+FDrReh5/+6HNMTILZPv4njq3pCTHY3OtS3VMXqc5qP/jbVJZ+RjH13VYmfKffYJTh3Ip+mRHA
gaYZajEF3PwiaqCm42blntyueUxQUr51UKYKnYBoDF3F4T8GHOGb8GXhVYm+VVC2EaF1I0+hvdW8
N5GALBgOgjg2FXGXIPx9j2G46AQ7x8YkWjKre+7i00h5dr8mVBOcilXbDaTsDtbj0ahkIvTxLbUP
12hbX1n8BiXoP8/7ymgOe9izReuFOEe5PAdJXFlbh4pEFnQ3dRqtcTYTLz3t0A9shnMQDqxqBY7n
ojiexfaQPfSHLZPsSzbiT331IxGiYEIcuPaBmiBHIOQFPOFVLUZavQzmPayDpiAJFCO9x4K2L1u/
0wuj97u/gTDihziZlpSiKmtWgCbIT/Sdfwg56COzSrMYVQVmv4i5hLy+bdLs+FTi75rNtTgJA/RH
HT9r46lyb3kSP2Jq2xfk2h0b/sMt4nayai1qprLzYXCZ6FTwe0YhShepY1fCTTTxOQCexR2nbEiz
VIgTf0kjWOQdjrVbR9E/kqs76qrTMEGGZfVcbAanQRexe4XLhtCiTnKcI3QhWoBPL2hauaWh1hP4
0Cza6iLMPc86QbFPgSn4mlL17utPX7T0FrDSllFwZf1MGoZJ99jRCHPK7wC6SSD+XmPzLe3ki4Mv
edBNKSRb0fALpR0+XMdUYEdiH+aoRE+0OL5Eq2HN4cmlr/k165Q1wEcdz/mxbOvDg+wH25NtnpSn
cHRJv6vPwNm1vGJFpIDqUqtNmkCCQ5zVLp0im3DRSxVCN0FdXMzVw1vLBhL7cpNLBOINNHhVaG1S
Pr+/a6KWqF640PYmUPqAde+yr4rOwH6tmnSn1tvMpRYCuGNk3pj5Nx3R0XB2XymZIqVIMCg135Iy
QnjpY28euIlP7vAPuURk09gcJwFab7fMAD40GCj9jrB2Of+Lqd38ioShutvy2G91yIpDvujMmpu8
uilEBCvltsEzYvDpQNZtD4wAKlrK6W2U8sjsDK20y+I4lW9mSaolQhGZsVvxmIgAf/ODx2UT6otE
RmW95taZY0ppVjlLEFnmhsMEn15gPdof1a6dRil/MLZiqj3yCB4Y05Zvyjblzv4UojsNF+4LNDnm
ldDSQz3VO8UaxJj0d6hbpZFYikENyDvL4f7nRDLjNHCdN7XVwly8k3hPp57teLmZcKggUjpmj4hB
Wajv8WHggMcQOcIhgRJqPVHUWSJj33qFY/+Byc+Z+aOb1dUnXy37diXVMkuQ8J3dDdvWwqxmO9et
SgcF1o11gMl3OPI20QmuQlJiQdzyOeiXzibVwXl1HnLTRN859JSMCf0CCa/sy729l/qeFEXrPXu2
HP73FMb8j/m6SirxsmpxCkPjKyuupGQ0qnF5rJHo83hmTumbJiEDm+tZUQ88pdAOGNEGqPzjIoiU
D2PPmcq1dzMysjeFgCoxAuZWYam9dqs+AlFlZobk6PXCveQ1SF5ZtAmmmmgeJp30jypvXCbVPks3
A24u62XhhHP5R7tXqHACeTefIznfKJAIDA/2NCZYPrhk2+PPVH3k3IQ4Ui77LWhkbK7UF0rC+TXM
CFRqL6B4Qv6FIML7DZDTZ4PvNvs0tKb3yA4UDXplTutztxozbFzoYHgMN4Q3xGTL60pQxDOE0uiG
+bHc0BfcpuUYkv/FcSi8iWGLGEWDGWdSyV3/1b+WdINFVEV33wLb7nIZofBr5ZTjG5ddGWKarKHE
M3KXErxdtBuA+xlS20sZscbX1LKS8M+pEKMdYce8YwiVwHYr9dGg2xbPovrxncwMW8PnIc0Nxyho
Eqi3AeuUy/AdHTSypq/h3H4wLH0YFoOiyOAWLj9y0IQFIiTrnd0lIbujKYU/6IRFI4/35Khr/upO
tNIqFd9woDYIfM4LKlhnopMkCXMduaksdlDW6/n5SC3Xing5ka1n6wug1DynDn8zuc9/udWLe3HU
92Fg/GemwEJDbrcl+pyRXKKzLEmD58hAzvh96x9ok4c9nwj9Ace3e/dNhe+tuoZi8JaHCuaRIOPP
XRftrTSPq061Y0xjUusmrpbU7/jYQpUS24eZQZ9rA1ML4s2updm9HtGkhDoecfsVifBfo5MPYYFh
sMsG6YC7yPH5lR4dRpVFhG8kd4jOy2quryBpyAP1JJo3btHKD7MGjDdMCM/VGwEVEimgxRSXr93r
Z4VUMZvWWhNsOiTE9JgPAyYji+kDEmsK9h6V4XG8gXVZT6CS5T93nFniO0OIWsNd+eohLLuXNNUR
niy2QskyVajplBEjSRmGdjS6jlpgI9zy55PHFenJTTUcb+u/ME+ooB27VD5MzclSxumvl+KLrw1X
Obb1srOC6uqKDNKaXbRYMlyUoRK8FBs+wHcJy0VhMn85GWs8EpmjYnuU+BjJKus1Ri+Nm9GIpI36
/nF5KFkLW8eFHVrsiznceOoHkG4BJ6osoAWHjPgYOSL3FP06yHmWj0cLTrcwbHvmd3qo7WV3SlnN
eWVEtjofikFLacAMFi9xjhWWnX7ZGtahs84kXOihcOdTjxc4cVbF28eQMIsM3GBrnygCE8g/egGY
21Td8YHSbf9Z4CrlYED9jSPSgbq4ffmE1jHn6zXVKWbItuiNwE1pgO9lfQLtWDGje4uYD9h+Hmrp
lECrZ0SZkZSTQ0dme2bcGRVCYo7pYS6wkdt4Vr+YrmGXSxSM5WQ8dAYQoglXLxoufoDpdREv/fFG
K87i1kmVMMbTvcTd/c1W0vfUwT0w442XUf5Dw5qgwhUfKcrV4511ScT3r5687WVLI3XFYppnY6XV
gKb8NmLzkCcwhYar3DaXWCb1Y+rG2Xzjy0mAlQUktgwGK+x6cgQGig+QmFG7whUIjHHAYbxXomeW
f7zIWY2v3C6LRmel/sF44hx4+ZlRnd3Wz4R0XSxMLmXaU7RIlnAq52/9Q4k5aMbNsByoUKl3V+1t
4YbWqKbeBKMTHvyiG5PZdTVB8fnz/8uBGt25Yw7dHNbLHhIYyIl+vpZVmORCuFVxIpFyO3s6c1wy
ZH+jqB9LNWGdCM4bFX7GRPtr1SbD/XQTrUBODsyiOHjPZBwvXB93CThOtEIOZPMttlNm8MAADXJm
DV9mQwa+RdYMFeBYB2MOchODB7o/KF9reb1gyiwTeYgbfVq93k1gYOc+Km6++hJrWqf4ew2eeGJw
U/2n8H7lbgmb8Qdqi+EOTej1WKBThU0VH3MEULmeTO7B0g/L4oCJfHkMvqtZ8IEoqnwnfbzMlM+5
VMIkd+8VIdcLQgXDS3l652w+gHCWsGWolNllXVYWe6/R6tRZ2kzhHti4K52Y6+tV6TOUwDzxOPct
aocygAGsp06FXtUmzcEZwu9I9XzoeVheWYmNUnMcDP+k3wPi9Q1TSAIvYmuyyPuk4G4j0vHd5tgf
UB1RaKblCpt1vE3S4C1rGg/8cab/sswdeddhF+23Cx1O//pw3fcZNIpCguDs3ORT7k6BT7y4K+Mp
YN79BngWc7AwIKM+8D47/k4ypZLidTQ6r/WwqU3GB2sAw9BNT2a9y8OtUJe86UwGlYnS3/fm1zTf
h/8bTpTO+mERE/i+O2Sv/GtlyYw0LgYirTwAjo4kwC+PnW4e+YthRNY5+Ep9hkoKNR5g0MgyEB+U
5/RhHBkBhVdf9TEr4MnnAY445M/FV4sMzf0P6rygMkqk9rHCLGylfOCIm15blVyai2cjUM44kD+n
PyI5KJd73ym7UR9C1k95H/vd4hjl5L+WCfMDfOSK4m6sUwil7xdC3nNtFq9pY4Pfj1LTMiohEMli
GtGjH1g03a1cqKdI4rlRxRGZ/h646zXTDYcV/1n/Itcm7VyeD/A0yOV8K/FJYU/GhSDV9UAsRoWB
Tg9OvSJsOzaKXJarYdYWqbyZsikR2syQK3KRyLtyFKQRUzqvaEfRYTqTyyJxTxvCEMcnky4cbxgU
XflwtW3qAyGfi0MdiosN/h+2+AK9kX4LLKgK8xFBhY5oVnmlQV/jZorxOH+2y4yUAX3U3QsF7DGu
3AhJK1K/PLpF3kg1LOZTfkVzKplOP6VGf3zWyaignA94UyLvzLKHYGNA62aECb62oBWp99QHdl92
03rgGo9Mm29GJX+9+chCLwRhDOQY1LBzrlaJaANIdkxqwzh4WZZnsv0IPUohEwZKqqOAH+F/nrBE
/NhocOrZ/jC91NnftRJN5KKsmUb43bObHjodRmlwmNjND9J4TGzdN1SlIjG3WZ/j/yKAN5VEWLe4
6ozufAhbmnIZCHC6V9WMNp7uJWGVEXjAUyD0BYYPB93X9gHoX/MTiZ/dvB10kPQ8nlacMlzKSMLz
51EO4NLOGsk5NcfIRevP8puVDUJ/OLkhZDDuHQi2TWysGDlQkPhRKTQB5eB1looTK9jVtH/zj6rp
mhi2FSXOIAiNZRXQQYO+4v7nbcpLi1ogjVna5PWv6suMsVy7LcREolBk91ITghLto+6nLVGjHjEb
dUqCPG6Lb7uSVnAPqgNABbKh3PjVGXgkgHIigIhCzOOqHTNDzne9K/tbZhbdp2mLdAxt5YS9IJ+r
ou0iuEIWe2nIHmM45s+vk7BmrVVDEC3g3s+FcwC/v/I/bIx6n4xeb7xHLS7nB2GdYJhLHFNUq9gb
UM94yHrsRwHaqL3YcEzwNpE0YvNp9eI0dDzoK584HfWJ8VeS0XDJqFjaY3nEgs8Djgwhr6A8MBgy
a3HUFAAwMGbXZHCxThpQnnqCKcIww9ZKjdJfly5QqHAmi23FKbeScKFob1aeQJmJW5ApGIkg1OO3
Ma2UObu3U6JWqegsrYp5KugHWevT2zpMqF3EBXL3avBQ4rB6Z+gu+A9wLTV2k2QtQXRbDgQTBxgE
GHLFOyBz4rVCaUE2yWf54eeq+fXofN4ZacUyJAR91yqrE6sC7aVSVEoqlTWhQyCYfm3taXmIeUVU
MyMVChaV4dL9eGf3C4IlVvzo3ndC0EOInXo6Linmrpgpu7AmnfPCqdj63Ws+Fx9RYMZM+PxC66Cu
U5Xl1VNL1i0iZEPvIz8ivylMWeqjqWIiagIc5MY8sbCSQfnj1gUTuVMhNdkNXm+XbwRzEJXX6Fvu
KUwOdkXch8YsIBNTn0J8t0uJbPTIZ6tnFgGQIeLKqxc7+XVZ37nuGb0oCrkaDmb6Q5wRgDCJLiWp
Gx6hzqmSTR6cn3Cw4mS7AFhShlIlX3Lzfp8DIyhTTqMMKuScglIc30rzBobCWjMaQSrMZ0Gy7VBI
gs9l8k5k0ePWvyjwggQ8J0G4L1ppmYY8iLzWPgXWelAC/1XrpVKnztlBJezg98O3+z0P9jYV+XqW
xYhhRRv8UlOY2/3LH1Sq0GIthQVcGhccFnbZyFMdA9leRz84KAD/Oa1O5kpgWCABve6sMmWKh9nK
wQ7iGTDAAuL0ieDzXxiQw1dCgC41+OxwF2F0kML7c6Yrfzj6axb9M3uz8y6FW2N3PjpMcCeXJDXp
oXASw0Zh+A5RnHPRQiDrAQoUJ2h93qUmbYmAhMAFdr1+lgXzU63R7yhpn5twhYaFrJiqzOjMB0BG
ZDQ0pHtpHxHZMUtY/T2wc/t3ZaB8VvN7SFnDYbWicxugPqXEAxaViTKYcPhTwFfpos8ZyIoueZDb
omyGX4CXWMLDf32pUH40ZNyqemMec8MFmKVhVKeVtHN1f//kkSeCV/GQkgfxQOehHMvsaPN/o7vl
LztuteBmgLGRvk7YC5ipDkljahm+RuHfEjapv6iEj3keTs9/VQYQ2QzjGlsNTIOXutlYTKbLfoI0
zmKBkvJwFProNifg5RYgagKV9cts0TUBlO6IJuo/PurLblOgTnHf8waze+nPUk2VVyC/pZ8lx9yt
UscQ2bHQclWVKwr0nduhHUUyqPncPa7khmf/vww1zodxnJPrU3xvTaoO0wDQhghk9jEru7v3hjdB
M/XL3vt6GQ51C0F8MPm1UTMqRHdgtfl3hMz3V7vAhtyOqEQGIwBa2f4F891E2/sG7eWank8kThDO
4r33cuE6sygrxjZl4uQz5ILgKOjIU4GPfnRXaXMM+oxgQhVkNUObc5tgNrkGDoyY/nuyd16ImpV7
w7vD+uDGpxG3+SNTMWOI5Jhqy/TaKGhjOqvNgMNvkH11xJqgJaRXebcyVUXTVj68OfDjVJTrDxkv
z9A7BtB06/gGk5chvYqg69/z4PF5uPfQgQMAHsw6PpJlnWHiI+z7SgIzmHeN+xi8l4Z3FRL0BxwD
uTlPbXkm+X5JCtevfX8Yyf3Q4vvCaYsREEYCKTUgFsgu6PdMSqSElCtNaL0XgQDZ0sE+k+dkAUhp
/ptxKpZImx44iD3XeBPnKGn+IZfdWCLt6wNZG3IuXr0dhIDXyK1CPWPH5L13CNpZ8eweUAcaugbR
RDiEA9OmnOYdscEPUKaQ34x6zimvwSsZ85vSZiXl0YW/jxdyalYKSCf9SDCjc1aHa1oDtSAhIbOz
xvp7QAfWEddjJR0gKSY9q5ZjXcUjmKQDK5TwtZQiwkr/HzM6Zdixh+BR8d7zqBRh5dsEviZQYPV8
iSr17SUSk8+CICxo0jN7PKSYL8lHxGHzYy31dO/bKxD7APznVnIfoqEFaPMWLgyFX5vIidzuFHJQ
ZoPi+07T7Aoy9TZJRni+ZbrxHu3c09LalTy6VByf7YDW0NZ9+f2yOuFNgzpsuLAarogKGD1VDKaL
bTuKO4xBzhLV4TOnKFlm2sISrDW9nwAF0NgYKEeftT5juXLHTO2bDY4ocIZz5gtvUntpStM0lxAC
/QXc8liXaU5ZUeidIN28asBwCZD/W+kx6eaW/fcLc81EcF8ChagwRSAB1WZQA62w573y7mM7RhVj
SaV9c58R6d3g4ye1Sw2hFnkgia7/7kI6jSUg5pFCJRWd/8jEzV7m0IjZp8s+YQFGafVIqQwQN9q2
a+1ZcOGmU0XL5gDNs0dyvzZQhTn8AHwYVMrwqjE2cWTtWs2VpMzTB/QDwabNilS2gmVkcgC/Unag
CJkC/5ezvqiWuXLLCp5mquwk1bzo+Y4YmPJcqOF6VGBtIapkPvo/h3CUMplvc/BVd5oSg0E7CPsO
lxDHxLMimXClK/hgXLvYBmhiv4jGXa7OSTukwU376vOVzDD/SWUi24M4uiz7+aUto4DAgCtOVUSY
4i7m5c8YxMpdlk/A6AgAKvNpLjhnDtEoq6dpfn0y3ftYUO9f0O3mc4xsxFSK0inqjNOGVKRVh/4Q
7ZxyQ3vHmYSRJmSwDBBNzAnIguUQag1cInsvMfWnPvJsTk9VXk/Dekd2XXxTxOPVLrUYac8JhaPH
uZJKkqtzy/rJih2IJsQXWQdz1QN5y4inDBJkdtBTHjhwQbQJs+XrLNBzqeOVQXXVOYlDEsUoux7D
XfLv8FyKKATk4zOTZcYU5P5q+1DjQbRY+0+wVG2T98C1Ef7xlQ5zVlZ5Z28eUlI/9h+XbG1YfpIy
EFYGYWcUlwzVtYD1AmlHNEs2sHILE8CoD9mrY/9XhRDPfiVE25XHglUF0edgmddEsTUCWQXoxxhk
BpZYJGId3za+KY+lFSQEni0wi8hKloBnA9wReZgx2c5nNSdp1t7wbrG8vPmew+XJSfpwrzxQb6IT
UnCJJmAQYnp3kjWPTK6VdgcNsmgt5pU/aiPNWveOkyyro9Xzs2pxi1BOipdXwbbfPnOAQBNdb4q7
3p6nGRyav7CJjLOKhrvBH9uuYFbZ/OJD+/quNMz1tzyQ17tyd1ZWPuQp1ZKzI5NMmcjIBtgFKCGS
4GLLFHjT5/TeKp3df7i99LICv/z50/zI0ynU4rQNaen67tb8CIq7SLg6vXWRsuJ2/oznCUAxQfv7
bf+fEOYIsw3KZE0SUVUb1dYo0l+XILVZmo8I32dHCgkxD5mczdqvkKTu9iCSnd8D7dGTXJYfTWvX
a0p/3P9D2IZhyK10oDN7r0I2MyjU3b2iDn7GalOPQlYIO9QUGnhC/eUtE4qDXklx6upPIP4nvMe1
HxEaXrWxstR8/H9zgIrWj42/m3ZSq0hfk7fuMw6fJgwW10JVNBD9z9U8/KrQyXGVssQp5I2iU0CP
0gvi9UBPjjBVVjfbq8+CReyZ1LLx3qz2DR2geMJYLrbkAJNJWKxC1HYz2xcW+yAm4wcJ+6LTiACh
/EXR41YfP5mfguJW8sPmxl4HSjMpXHqLvtPBiKhRtAkA7+nKP7q70DJ9Ffy7q374e+h2PdZroyhA
4aAkMavXUo+LfGRDTTIOIjPvDXW+0Tq8SbDdLi9V4yHklfk0hJDFAFClDxWLufDYCIwTuQqPrNSv
EBo1b4nuEvRvfbSNDbwp8PRU02NIG1It+0Neg9Wlw2HQVGiLQ4hTsGUsNU1FfpW56sIjTVEVWyGf
eRrWCwDVPMIL2qOxohjsM21x0cmqio191kbwJr8jisQ7w3d9uQL/UzCI1adDhwSQBm7XNN77pIvU
AuMSyHZ0WwQdH1eYpdPuiZHEyMhPcIf095Io981sTvy27KR1xSDkh4YGCK4rOa/0L+d4EBPIk555
pr3T/ilCurQAzVJTjO1WgZbIE1w3MdF6P65fGobIFXvTGc29Pd/pDmNqn8geysCgvZCRHZZkZzFw
EWoMbTowsvRpEF8rJsMDqmMTSF1/MoG0hHo2uYYfG5thFpzkq1LmN4oZXPHpQnMEKY0vjZRUvgRz
A1oIuOddneqrZHLYC34+ED/Ffjloi7zPdTp/mUP5/ucC+PaDU14Ok2ywVv/V/8yopahulVb8YbzC
uGFNC5HTJbiz8SjgcEYvugjUC8XqL91dyN2uAEj1L8Xqnp4nYJ/E4eThArF0aRm3LyXozwoJmgCS
r7655tpcqzYch27jQLhFULAFAlLhIBfGtjBjYMntplt1siwYvFFtsafu5niV/hCk3Ob4h1HWUQZL
FjEPyJ8WWzQXwhXxoRTMVUUCqIn5/8eMGzw9GFtgQ2rmaAY6b5Sm0Aqw4FZzc06zV9jhYHJuWqM8
ugZDcb2TYtdySKq55Iem4IzX4fp9HY5sswwhZPKAkMbxuxuxvpIiemmhZPe/DOUPUsmL/tGL0/1x
vgIArhHgJwECop5JHDUta2dci77ypEA8BgUTMCGTbpGedlx+Jj6dxzF75tKbkY4/XxflrJ6jolGq
7t0yJkewLABUTXD/ARXqEpd/jyBAuB9n9iO2050JCPEdrpZDfaWKeyyrxsT+pmcyeluTEizXsY3S
Rnz0eQFrS46kbawyUpz6W4GGX+CKkxtoLyoKMUaJA8++EQJ6NClg/MHEwn6b9Jr42K/FWk6NHLWi
hSMPz4DANtXYatfwoaE/1xQ68keem+IfDcsnv5299jXttiw3/MaxJJ5Y6XpCtU/sZ39OtVGyzGRY
UWY1maWITxqLAGfVhWacjuwqFqR/z6OR/eND1G4hAnIPA/nGH5YPpb/dVRBLE80edK7PgElHEvWB
1APwksLgrXvG5g+dw87gPj9d4j79JpqPYAlt37VjnCoDTjcGymmnFg2r16b+KjD2iqdTtIlNcpx/
bfRoWUGXuWZO6vZtbneUaHlKkAooEgOpCM5Pn95B3ckoAhQek0SqEnaPgV6qfyoScyZMqjR3DgTs
zcWgYPAFmqInEFfgsqpXzqAtUcCN76YICnjJJfsoHgGVwVOdCf1UnS4BoBld3ObdsYzmvPT5OxV9
kLmwASIUcxRqy2LO4Wt7Z01tZ4L05rsD8UyExRMMSO11ti9oSNa7LkAD3pFe2y2/QoJcCsFMT9zd
XoEEw0/K8xEJ5z8Wl5ieXSVtCLon1NYfkJgnfBXMpe4KBGch3aoALCiHJ/vWLNwKxQpdCLKH3NZL
OcNvyroTQfUgY8+5r4hmbmck++6weaENeH+7VSk9x84NMxKBBQX9UYtHmwCZSpfuYq02HmdfaQkP
ZlvEhuGWXa+OYFiJAWK0zjQUt/tM/PD07Y47fDegJ348gIWP0NZUc9TFlRP51cvu1K5DORPg1q8A
zpyWUnzbHYvtvO5QLn1HAKxb0exZRTgv5FrFDqeHYyl91W9z1Lgl255QDSmLBw1J3qbtibYh0Ovq
mUALvrWG0S9sHCEdbBeWRtJL5pRYN9DDT9MRf+R4gxy8dLCXwSh50SdXURCFEMHMCYIGutaFQfxU
94L8LyvkXbHqCVuo1AgZ0vLYUiUgD9I708TPfbugLauj/8zqRc8hkD8YRhLWV7kREyyq2G+QVJv6
nXyF93qiY17Xmyjtxg35uRNRCbz1jbPsFvGlZj61F8fn6pMKkoOlq+Xc5sCI5J8enpvN8WKI2G6u
Lf2hd+3ip3u+nERALHp6e970mW+tUaGBck+vC2NTtlkUeSRrx2myTGUTiL7K5dru21VN02KUc9dZ
BQSTsuzvQNsvBQhQiD4ishn6hSpt3C9apS/wO9GQg6YXsVQPJmHwKXzN6OF4hGxr9n58clinUwAN
D4rFk8dyZ5Mzdv8+iMNSrV8+rLt3fOKTNgJt4BDdR8x/TVhZ+FGDLGjWGuGHuD1tsMgT/eJQoO1i
CTNl60zHLVPKm6TYNA8jTDjFZrx4qtwfia6mkd01Aojvy4l0SHoh3darkN7ub9A9+0eSY0XaHsv/
CJ8FcyXCohx7FhbxRrMHQC872Zc2KbGT7MYipZVrxGoi7vZJdhIL9SmC1W5IMybJxveteg3mNzIu
28Tbqs0FlmkHyXYn2UWsoyUlfrR1m7RqVWB/Yixc0YfxEBuUL0ucIXlAqa2XjSPODIe8jaxRxk12
KJYWATyO1+VDW/loMqFbjKla49wq3so03nLnF63b2ZG6laM1iE9wzvu+gHs93FC9seukiXWL/PgZ
MI4dgxnRSIrUwHZt7qiRTtfCr9MW0t24xSzZNNOwVVV8dGVdfFfyALKiD8m1Z4VdI9zZrLC4aeWl
8iPUue6zFlZ00kGMl0Se/yBj0NKJ/FM4hwPuyrUzUJFowXDy4lr3c9MUsD8Io3PssdsH8BUkPsF3
Bgb7Nrj5dHS808kO48vEQXJ1wpDoPaBrspGOjyppOTerjk/HzDIaj8S3Jp8HsBn1/2VnlNH8MkQH
6cCG1KgB6e7GYCPiipDgx+XTfYbgQZKApjdW+x3ZHqGhM1WxaTOYK9HAYOgJoMnponeEBcAlOYqK
IH6lbQIq/8AocPNG0gRoDgckXJa+DrGuaCbv8HKrFj9hReRMCNd5m22mqVANydb7i0HxXJjqiXnP
BhrE3wd66dL/zAEPXo3EeAmM/5pQmIybKfRHJZdoi92Ek6NKlMW9hfuBwAD9lD6x4v42KwmsoOOA
2Y3VcS+Yu8iE8hz9LqyG2f99cvIxH96EQOrAxx0Scp1qzwK3QZbwfANdf1boD0/3VIRFbh+pRLFK
h62WIgC+n6U7Ixhh1Qjv8OKmpBeKD/MPq3URyyqvcTRmLiO/U1nleQBW6WKgVCEoA5B/AFgOpsA3
5FZTWi/ImGpsI0y4m5VIcY3KGWeBKqOrMyG+8tiAaKDD9AXz+tBL9LCiu5I5k/vo9D76US887guO
i5SP+EzsO9MDAZ4547TeG0ZI4o/4/pk8xKS/3LLe36za63Y9w9goGQC7a+Blblm4zfG3X33LuDGH
TL8hbUA2/DhEp1B8cgyvwbZfN1KqOOPE4OZiQkWPds+b4b7I+vXrXeAxhfWzZxUVYFlH4OVgW+V4
7nrIqsXRDfQ3WSd6p0hIQAUhdWMmnPScY5Rvmkd6Y/uVgBr7T6TwHDDFDe3ufQD/z8HjM6vd7EOy
6KpOL/FxEDW8GS0QECXEvUX1O75lCb3KMcn4rq1kk1/I3AZBT56vqoZY8feCOMKDboHoEu+chI+E
0DtU6Pg2VRtrvxvNpz3KEgzzjsKgHouHZ8/vjp3L7tdfEono57wO9uSdOG0UWR9X8JWkdA9bobx8
Iyb46W9/BWNTqwl1kg/SRKeTnIHurwo9nJeO5TxBclVVYasux+jv1UMx45ZeBLvm/8JutYUWHOE1
kgqmek0C1Xw11uc09bK/wG1u1W6qrpI2vdoMz70Kl2DW7SjUaEHnNANInapa0coPnfBjWcLKDwm7
e6dmNmGDE6ijGRdhQdVNb8xLSsJR20uYU7hCP8y8qtVcTDB77EsD90az//9XkXGePiAS05QanOyo
yHiVuJiRzBSSdU6CgR4IL3C9ciC1V/clysLL3RTGU7b+tCCUxy3kg/NYdP1k9LjxDJPkiK0C/cjq
QPXmDAZHzh77dlUimNPnWL6X2XS1vLLotCVbdpoRWp8JSI8068RWwV6E/OMRM0Ekmw4mXJFuh9oY
tOYQlp1qRLB0bDREqlIqPlBjFscDbwM+/SGap5grK+HdLlDWUMkc9gyy/uDbZsNGtNm8HkMDFAS6
BIZO2Va3SLMPdFqWX3l57n7Alm20v61b5YOETx+TYo77W1mce8Z5kheGBi/Ld4g97YuFBlx5kMNz
Z86O12KcxP582fa8S0XwF7OT2tHC4ctw5CfZAbq7crUjr5dc2R07luQHXo8UQdDeoAJqnuZ5ULPJ
tOIxLOXe5rnPXZ4i+isu0/UE2/IYtFaLWtcJ0Dp0YbcDYF8Mz1kbGszPGnAYQ2fehoR63pHicE0o
jURYsQa41JCTfZbmeJ/jIx1rinjxOOZA2jPJxR1vi1hYIIAhXQo6r/gQBJtFQfbMgCQWmVf+LrDR
xL0AiGXXvttDIlUpgxsm1+KScBaqhAFbYkX7P1mhVl44Ljq823u/H54dygvQrmOsQUbdUxWAHy7Q
Ry6cDsr6T5GTYpT06XV22g6XSYDHghTK6dr1k/tQ87gE9Gxsw78QJo6Dfn88dmDBEs4kGrQJ9Il2
5io4r+duetdezeCgxiIuKXMeSFgQ6d8dEQuYB9M7+n8GMoMkJtMW1DSupYQ4STu3hz5gehsnBmyO
cqzQpFn5z8Y/tjqhHEUuNRohzjygVxykDsL9ACXHloRZSm7yELGX35fCWG8j/7dZ9f2KZVKLGpT2
8pGC/kFXT2trFL/MqfbO/09kXW/kQuDMI2XIN8U52lLftmkmGMzmJZ0HwVhA50Vno/bse7nU5cbe
e8QXw7oz4ILHehVxSBVpaWDpM1gSKTpyU68kU1DWTzobgR3mgF7jmMKuDvBn5tZJwepE/A0BDyKA
dHrrFUzS+DBWOfcggTvF1o5pKH8RHuC/yOAX0TUg9plzyEF+hmbV+keiPQSBUlvdVEGMEuzP0uXY
ZjgPb9VVcBMog2eHR6ZJ1tK1v7FyXL6ApNayqoqy6JTzQMsQlMnYk+f55hhcNZSiV3C2GwqSHvTf
TpcmXgnynenNhTVsR7SCr8HMneuPN9RGhy4z+jldcXCX+cIi+zVEmK83yi68SjfiPkxl4iyxlMpH
uCHEGUP5NYVeiJeY4dgwoPuMpeQGDSW4qtq35zBcjXCs8uqC3MBd9ZNjaTPnqwZRzCrajQj7/WYO
SLVAII2BdrLMqUolQrNKrGVhsG3ex9J88OONHm1P9iPa4hEsECiGrPIxV0ntd7mSjpHd5O8+jr8O
k7qaxngG6hu4wqsu33aRyrauhyNEUe695Uyxg0/g4it1OQsS0aXJIAuFZ99Y68U5OnqtAf2QkVum
S46SosZgrQwScmgE5dE9FaYhLJ3lEEH9fdvwMX/MLVXMl4Btr4jsUADtWq+v/NQyuUwxZS1BCq3L
f+B1fzGXV+hMg5JVhkA0anTkxOdTgbXdP8F2q2KfLwMEDzsou8hWxC9cst2Ns9bQS8psOEJ3dNV8
Lrr337uaG0NFTnZYMHsmGr0GNSp2q3UISm0jmk7GKh3/LWjn2dOWbtVXMIgKFZpu1wTeXm8/eY9X
HDjcYcnxqXjigZZDgKGbFkK8Lo1DYEOWn1+uD8GlCCUImuua8emoS5APadFvJ50J5ngq9vLBrZXc
F2+RCa70xKSj7i7kB/nbuBQBJCV6NZcjpfhtqjEEu49SV0hQoWIHEZZ210MxVbLNrZPmvPikesH7
SAUcc/OyWw7w1aHd2oIMQLzAr7SPI9JT/K2VoZx2bz2vA8AyYKMpQQgNe/Syh2A6jjlblInxAH8k
mLIferiba0OhDGhgoWD0CkqjqLGSzWdg6tfP1k1wSsXbESpYVGoNzaZx3m07yvArfzJjZ52voJWT
I7unJsgaD9LDEagBlbuA4Zi2Ju6pgl/QOqGEJCS4y/92Uf5hb6h5kmUysRh/4kNCmQ21u8llOjjC
wBPLZ1MsHGtCBXiG+bO+EwWI0QZiplQNGXSqSMxdKkBDByCVOQxHVA8m2zoJJmMfiXFpt7zhJD/F
vtMwVws4ZS+qpnoZDPQQH8InIqXngxVvnsfC9qCtWOznxgP31Sad34d8iPtyJBsqMVXZxVG1tlNL
E7bZqOHd2pQWwV6lsz0Ns1C+fgXCxTeL7LEPsdtCK7WDcTyNSVBPnbUbyQ/gFPvyfsaFQ/2lIFL/
dg0I/43d+spze0PtsxK+IGi4yzttfqnack6mQ8I9l18nKS2Mz6e1hqzbhUsLojF6GLEF7gtlkdVV
WTZxusdy44fdOC7lBz0rdHRWom8vESAl6jp/CWsbuBnGQYQdijP9P5On+MMq5pltk4Jle8n6bjB/
fW2YpcglXrmGccpsiCG8q0NGT0drtvDcdoFf08w2sE1XKGtG8umnHPWfzPZUFyybp+FquY+3kOFG
hyp9haKsOr1g82Epok/1TeX7U1FaZpHRXi9XGgMFaYi6HblP4nt3PU589dMzcRzjfLzLFrxMlvv+
CYHE479KiYNbHv2zUWhfw8ZvZIO2mkU9inQE6ohW3Z6fJhNaTb0MzTSqRL1nOqIVv1NpbmVxjZzH
mAUHqTbXmIRx8/xoeh8mKQSfGflD79XNjH4KZC6mz+S5XEsPjXkHwWDBkrUwnKS7m05RI76T+hwV
ynWf639ET0Zz6+TwKeNfbInH4WO1UQpccUNarkol9PSH6Mahg1w11FnD8MvWLgjaiYedTDC6LhMQ
OPuJgUy1R1Ly4cZVdmKcasUDy3ijyDHqMVcX6wqr5YQhlntz65wB28mF1xYA0m/B3O+AMj12E9t+
0y4QTpiFzwA+helVPLWksMcP23Sh63TNTWhmQYTKV3E3mYhNk4kkqRnlwF46+nOWit/jggAgqwqb
jLx31Q9FWqa2MjC011n5Btry+S8L5nMyxFjX389fKnzJFVeeJCwW+go58lSrJN343abbUojf17k5
78yV6xO68EyO1bTSv3cyHLVrYB/bLx9SWVj3/uCe4OTM/ChkikzaXfS2XMU1qmjkldthhzmuncxT
qhL/CQV/Ejm+zAq49GlKHYcyoEpb6v89RgXhbh5H6wZnKtRRqMl2hd1G5cRC65BqCh1zTh/dzJRy
zt9mP8dTymEeWgcNIpFN9HRL1OtKUPBaHOGZpfzcMkk4Fy7MMVAviZO6yKRulHuNw4K/kujLOJQU
MqPka79WN7zChfRS1BMe1byHZ73fEUKYrCpYG6Ox++BXK3g7RMg0C4/FjrHC8jerNKwG5Zjlk3//
DYHhblLuLpkMkdRFTfS0zUzWXFBe6MebFJGPywqKHcVlass+14/hgr/aV1U+4XBKYN8Uq0zjpeQj
A7tq5R5bHgb5XcGeftAtzbNfLJVS9V838NJOA4Lh4BttaW7EVt3Xw6P5DPQdkUldgO+PQkA6EbUb
j/PMrRv5nE2noBgXq5KWKhG7fDWxjNthnlvbVQd//pPOBApin5QY/w9lWP6us6MKWmoMs4bTqCty
Milxvtj7ACruzLel/9ZtdOEDztEGMCN56JbJR++EZy9QYCaSqciZOuraEU7Qw8MStrKNtHB6n1Ze
RvUOiW6uKm0EiaDfkZRm6Xvhe57BFVKtXWwHJbrKE1XmF68xwTzi+Ir9Mkagqc1TRrAPtlXWgSES
PUBgDDziCkuRbEJn7qnVAxDtnsFLMUWWRay6PPQmlOQiqV0QwhMN9gIPNK7MF3OtCLI89GmqL74A
fUPbnAoOAgBaYiVynZtKmzFDNRpJ4UrkPFuv+E6X4gNfxjdNB2xGXHqaGMgE2/BKIERA4YRvnnnX
/YLvbCzr4zAhouQc0dYf867XihOI68T97z4AMIJ4KaJEoIz5hC272g2LGN5BEh8hb0yrhvCV8JWs
oJFRX//apRUFFONTDRxCvFqrBzWMd88xIuwWrucIgJNm1Cf4dHeHvvq1nc5VfAXZClQoRt240eud
beZS9q9CRIjmd79+27OOj/Y2ZSs2FH0O96S9oTdmhFqk63cIZ5GSCnnk9zujUq53SRq2+2dx2LYl
eewYsf26QajPGsq8Q5XG3pkhEPhcqHwt9AtQYomDj3Kh43JEENANH3XWHs4LqpULwOu2prZB5wb8
e//yNLEvnHgzoMUl6jz53pbsJtQ//PrBBUt2tutPDveD0r1x80K0LwPoYPEegqqq5Dh/enfss1aX
qRugEaAjK+HGQdHW9XWGG3buyRVzKjYbnLn/xqMzkbWML90/vyJ3LzGNxeozQNMrydr6j3iwgCIV
cqL/i2KyucwrfOic2Rs8YcyHedyVRhpAaN/Rg3nzi6lEcewB6pYZ5q+qkwHZyUxCUxm/Cg3FFIf/
Nrl7iYlPrbIq1bEHeqblmri+VXayFKdl/U2oUV0+nvQ86rFLi3xmShKJjUgH6KWn9HCPMnuTtB5x
De0ybmphK3tLICg7x4nlMlJf122UXsq1ydWa4Ib8o3kFjG6cl/SPZN1nCHEbLOw7qIf5SIXf6qRF
xjHAh4X2irJYS5RNj7dF/UCkSkX9u3jm4eXLTMFkkejn8mJ3xiNbaOQTyOZrcv1WDzGd0gqri+hZ
trMlW0IjBN1MJ0FomFgF+54h2rwX62MOmHnL1Gg3ItY6Qfwd818TKhLXlQ1fyC9+c48SAExgKgfJ
s+uhhi1YvpACCWARxfNEdjk4yVs4d5gKTK8dsboSf+fHvOPl8RRV2Fw5VFRMc0MZHE7JALqrGmDH
AOdMkP3ScB0W6X/T5nc9jA/ECPSMV29IlC/MjqRDUeAvflrRsxn5ZfGFwi3+ixM3MJ1Worg4bM3v
vZ7CIr/oqnDRwc8PiCx2j7YvmDipqWC0XDOk+8sZ7zcDqr7eXC1uNJX9TMnL5X0L6loEFo0Y5p8q
upe/lDdn6JLapcVdGnjE8el+P2RKFqEIFGA3BeasFztkRZov4Id83uUYtmjIaw+R81zue6V06jb+
YaGiNBuYgkC/uFVZMvc3y5hJirg1SLBXZOrl0XHJF+jNm1bancbJ0/PqNtzb02Tenp2EAZS0CsH7
ri4E8lopl7bhJD1Gz+whzgMk+C9fX51Bi4CJq35OdsCbFwfsOh8fUKJsZF9TXpk+hvuFr0aH0OQM
IgfWc7pnGR0YWxK2Kyc80SA58hMMYNyb3/AWc2N4OQJOVFGAbkfXi2eSwDE76U0snWHd0+bu5A42
ndrFrIEZyNpNJPXM8UsieyUxhPIWRzaHHBZ3/GZkxTmpi6I7x5zLA8kuZ6rQgiE9/pOvUClOSyIW
BB9rA7/rcld/UVF6OkWhRVA+HudyCqq4kzZrpHEewa4SALp+n/m1UyN9hBPBWflbV4WSRU6EUyzR
Eys9BXyIgE693Jyj8x8tgNIe9nfwYNAWCKjpeY8vWTOuGi0SFV1rJc6kZn7OalDEImvtr4i4PYGQ
Ksue2pl1mvd10//kdQHaj9566ZqdxNphOoy9dmGJ/3VeNaFAGi+105yq1v+YMC2K+vuB25WsPSyH
oSTwno/wPIiunztWIxP01nfjQcILYhOiL+D4tjNPBZOcpJGFjcnhu0xN8TALGKoUVIazRkpeIWlc
Ht2WOyvhjoioRYf5lrrfjVXQ/USWeNLJA0u8veT2ELz4AauQgGvs9RYb68fyx8hSCHPOgQ7PqJxU
pxnQZ5ePAZNmmj4SBbijhH81ohAomIyJ9OT+S/gJQPs/PBFk4EI/MTgbAJlaA8t5QYLKCn6Z+oUg
doDbOCEhSk2FcH7/WbQozcTLMoTdYVSEPH6HSNlwcqfAy6g4EPbCRJu7hnIz4m+zf0bkJ1S7o/ct
9xSdopqQRj2ONAri9G84EssvigezGQChBDmehMydOHcGmJjYmEG+FI95+W3rA6eqgE8LVhiBYapk
vQThe/3pTaPeM1LYIq6Z3HTIXgWy3PnJ6Nof8TNscPC2cWqjtZpEUMUrCIf7tSyvGoT/e6G1luKN
Mg69I1UtTPTncFVy4fNJ4pmoFnf8oy5STgkwEb/TzzHT6NhK6tpovmbTn1IiGxu/hyruBiVpuRMr
q3ZmcCtbAedvekIRSwowWBleV3X2CeUsw24TmCqzEzpxh10p0cT5TrFqnnQdBoCqdom5WBwvHall
qb8p2xJm/TE2n/nbsE1u5SZaH5O4EcH5HetKY4o8ks0q/zCFqsjZCKzKziWtDTiOqEqZGHv5CBJg
fWDmZcWCKr8VKskyY/h/bu7PbL+K7tPCckma47tMvriOlOfuyBOPBXvWVt4JTFHoiMfCntJe48p7
DzzK7G8q8BLCu67BNQcuY5pQ7ZIZq8lCkZjc6QJpBDQJF1mtzVEgX+cllZmgjZ1whemmpj7hdiAO
DbfPaujMdoSSoonKx+cVpcf1LxPUSPcT5o/FA43Z7PuXD3Gans4ppn4YpM2kELx3/KV9cy7lcNqK
Cm7tk7yYAM7lEFMtkaWkNCEBOB7OWQDI38KMSFCtLhuBIgZ6nt6aybX2dwlJxFhbz4TvuaSw6uZD
E8ycl35wE/PGTmx+m0c+43oRnM+eRVYinotH/j+KSPtk+FMMOTUxAvVss5ZDM9pFjTtCZ0tp90h/
ZL1RQQWpJywLyAlOWDlW6vt/7PvRqvhjrjUN28+bhWmeSCeD0YnIwGfcs1RyYBNhnfTBPVK1nApO
9U3m67L0Y7YKgnKtrvBUjOf5DMCcto1bhyzHd88Fr+k/TSH/oiopypygI8RMtj8qH+crLD4ijpk+
k8aPWGYffGP9ysSfQhD6mPpO0CxMCCbuqY4RRhkJq6d2bUB5evwLS6I0qqliyL5IfYVmQZYkcA+g
9FQ5TUVt5EMdMw/yWxYPWsTwapnMX9GScB2QfLOAeWRkCpHjarpiCl55yVcvDgYMMmnAA8sFfhSI
yMniBTZaFs6fphc4l6hFUMtittyqlUdgqWkSjhIj5/yGrfnCCzU/tUFXfk9zVJVBvWD1Owp9DDYa
nWnNCtD+b4AM1/z/218zCXq6o6aTcDbpQuDWLUNk6ULF7QFYB09AWMV+8uq2l/8kxGBga/63IQE6
BEFYNWLK/djakGZ0BB47vI8DLqgccAzEyS/JKAYEWIe+Vl7oywSkJNwmhuTBBHcveEQluwDE6KPS
T/yT+/yFoTu6gVCvhsSGza4tfueioUDS5YLkKw1R9QQNLh8Bf/Uq8kvojiDMVe6XjI3qBThMFfpz
JTchM7tKngbMude0h8aG5RItVQdYaKlzVn3Hg4hf9CPLhLA8TRJWUj3RT8D9Yhtj2HZp2RE/kS82
Sayt2BlfX8KxWiXna2jtraAmtSGlpKmd+hg3rG3ilKvJiz8AYkZhSyU6dUZwASMaJkvaBBjV5kXy
fxo3oDSQm9v43z1Kf+e+4O91CAqDW2XT/PR5R8qUPQ56SWW7aKEN4MyKEFarS92E96WCdlHyxHCT
gcDvplmtDWkoPKN95VbRAhxwVjUo2P/ZQuAC4aC6nlMNdxwpbnpZSmCHjf+ojAqUbo+0PGg6AMUs
DRiq6pHYORWuUdGULaktRBDOcjwNsfrUh3/+DxSJP1bXPxjfMHMlW+uRorZj4bqemQ0IYdYCcl6B
MiQxIUoNrINgs8jp+ipXbtDUF9YfkjxIZAeB/bEBvn6XpxzIGmvezSugEyEKB2UZzhy+w1rU4jUc
/RCdeyQ51DzMjVvKg4LEeLogZiN94luboCZl4+qcQGbQ0z46Swnq11eSIF9DDNXkjZtxmQv4bvIh
HRiscx04UDesoCG8egvlwju+ywGaDFpXwN+/ovNBuebj9nfzcKbx1gUFEO9EFkh/fcQ/E46wIxyw
IhnFwGFkVilbuNAUecFFTvRY9PKD+KCXywZf2Dn0lE/3ziqASAmlc+PPpjiJNQ/8T4mkiudeo4T0
QgS7sp6AFKsgckMyTZ6DFpNO8WKVnBQd6ioLpUEN4Ttd8bCTmb4ufGHwYkddwvrEM0chSmwvP5FT
OTPAHMKN5yQy6DI6XgXhl/o2+aiyWJHhgvtr1fymMQ9W2DI22zhGRBu3DUIKF+9garPRqEaC4x/2
+RcS1qsGGiMicYw7yvarff4NCWWCnplCLBVaeJiIPkOmNhv6G9sY46reqeENNB2QRHSibz4NVmsy
NLT7Cab8UrXkefISbr3YisTctgSrfnsRvQClVFCk/tX5mbmTVkBfIefalkg9l34cmh/L+YVMJbXc
9V2dMk2Aqur6bnzlaDTnxmGj93i3iGugLVRHnitHvb5C99fE7BhMCkRrvUvzH+rE3dxkSKjG/eeU
kW25K15gTmcaaGIqKTYw6CT3wlu4W4vXmjM1Rr/JcfN6lhHE+sHVJ6KUWRK1wpjPiDAvEORJvivE
1LBaPBX0dNbT0QfU9hlDkkMyRP1OsT8S4iLmHnCs+7+jM1sIBjqOl9WiZp0tW8T2OMmSjYKC2or5
mds+gguiATj6iBtTlZxyX6COZMMVHfh2hRupGYXNLbfYTrP7OGaF5NL+xz+9zF386Ow4hzLZsJGi
TblvehZrZb7s6nKKSN/KmX+HuQTpXpO7K/hPRI+k9Uk+jZQUgm1hpnyWtROTrxjOnKJIxkmIWxeb
UeB4OlGugcBgmFljrexwcqrcy5TubRFZMXpQPF5+CWZ/eXCCZTkJSRSWWqmFVdvXku9ZQN3o0Tok
Tqx16F20RNpz5XSHplYiZbzX/G5JFK41YUxOQqeXbDRSAKy4mkiJuU7SMW4QhcCYUw6v8vIj58f3
RIfMu2i48vzZMnCqOcdBqja6eqYVE2d7Qq0gMRpfH3duM6+YKyJdwjTp1PBZuUJ/N6z6vOPTFY2f
N6AXfJL3m9CuI3Ll0RuAZu1q95AFi0hoU3YbaAYCyBf3PUDvEmX2kmqbzEGRYxFzVfddNfYqxWd1
EvjExx3pGVlCqblzst+xGQ7KALtdxKf5cgBsC9njsHG2yrg80pReqANt94Pzuw/bc6GO1dKALBy3
VcdzzlFCH4zcIrosaefHqHOcm3mDI5aalxyJLw3cql5qhobFJEd6rveB44OTGcZbGpw3e/f57m2X
+sYqJjQL8zkywwOKyHavVtCsEticewI5Vfvh7UOit3z6gdq9s6WTXCv/n+rH1GNzMZaQAGMXI7z1
DmgpPM+TBhFIH9PQW2mdwT2IUINjX/XGcz76z5m6ndlpEvNHCGvJ7G9TAXari5k0Zc2CiXwjL12Q
1lbXbn4NsTBeOpGE5jwYj+dT7u6gHTAQdy5dIp660DTDBaPCY2Qn01+REWgTGblyUEqddq/iMKmQ
ERD/Bdc3urIOVqZ8Qc8qX5XL5RjBLOPwwn11u0Y7inNnj0Yq+4UCsHsFHBKiY9PIzhJuOYiY/q7z
/DMaoWOIMHLlYG0syemNR0AS1deporcZOepxmWOfy5hRjr/L8EJf38HAThSr3aqjAXY3uiQOU8yS
pDPHmhkG5sx2k20NFYJo6i/ISYDnf3MVf8CTfs9RwvBfgvowx834pORah7/SW7q6+JoQMn4a5TwC
PT3rSC/7MLsyBZp6Ec6jqpU1t7VFvgbOsuH8e/zsvbhts5UJJ51pM5zxwutQq6j07cBIeoPv50kC
Pbntj8KwK2pt8OG0Wj2+32HGTtniKlm3i+9SUKV2nBR7yB6WTfzbwJVzr2qswFN5lSHinUXeCi8m
Mz7GmVjBuoCDXOdKR3fF7wQC7QAF3yVotRUXtMoguRbMPlh7YJ5acNejSAqUMcOhZTPMwnUQ5GGI
tTYJYkgru/HcNLLXxKNzhtMO6Cyx/SfDvCAWZrDAa0hXnt1LNDyrAfxRFEzdIqounTGYwnhBk8rg
3oiiMloUsA9vlMBaYejgYCRKduu3zacWAFdrkHI9jJQhl2REPHYkGf7EP5FOG/jdmCxeRj92r35/
d0EKaJAEZok/LvIx27z6hwH82Mi4up+2CO2bzKtb5B+mYXSNlPmJ9tkc2fE8k5rybYwGRaTCR7I5
IRBckvm2DMUBqwXpclxYVG1d4gITYYCe1vOyM9ELDMSVg09jYpcy+ysooYLICi/J3AI7VxDaS/pC
PQ540UxSTP1PE4RGcEbwY3ePRVuZ7pJ+aLZ9t9MSq4ad0nuFjTsqDjyTi1yC83diOBysT0KaDlMR
VNLKO9AS+/WvD5RbVfOhYeCw7wRc8W3W6WRY3dJob0SLMETQPqUx1Q4UZ2lHnMCvI4qAKeNQlgz8
SZWr4Lr9hK6RKqbEVgU39ZZxbZVwPD0RWgWcp3hyCbkSyA4s4WHCTnZLVEM8VBc2jU1gLRfrWSrC
iY6NcCdZvGvuxJD460EW5d9CIcxRNmPgPS3mjaar3IwvfRnEIJucctpYr6fDwM/iwP5deyrz5jLT
GaC5JTSBOc40h3PMGLD/zRNApb9jx/WRsdVxHwusCJ2dN/VTlNYbpIc3x47XgD0wx0NvB9g5Lf4k
DBSPlv22gBD4ZmruVXWtw7Z5jCMkGmfRYifkkuc0CNcXw7+3jATSRulk6gdycFy3e9vFQrxqXZ2c
Z1OSkbj8jdTTNAxv+jKkL6H0V8+wWse1wQ0upvFixBuS3QfgX3aD3/LTbeoON8MZZytFU7bHRTn5
VOiWzQB8eHK6RLaefGplodNcniRfqtVauFEIydKKQdlHAytgv1HRT2deK+pSi72RLbfr+019rI6v
UQHdQQ9HhgmmAoMXrWDaGF8wRMIcasjL6Mb4ei6CGUHTml+ynYMV9CWc0QrjFXeLZXCPUELQ2dpw
7qrn9V4tlw5JeqbgYFOkP3l0uLhQfyAkDZGl+ivRM+JYo22m/0VX/chbjUeWuwMm2rF5x95ntgBH
wyUoG9AdPz1iytS0+jZdN0zQiRyjxynu3YMsfsjUxE1pnaS9dO0Dt3TsthxgDyOk9353eViE3jne
Xu0XyAv2DghJGw+MqHMLTucjlcfpdDCkFi8tZQxGFeCL6xOwpwixA+64SbBNprpMrHM3ulB0YZNt
5uoq+ljNTKyFaMUFf7aJ2tjuKd8xJoo6EiQK3/krvXGrIvtzJ5CR8hdeKXvsMrjQsWD97iV26h1p
1CbV1BH0SHZl1r4TKSF0cknhPL4lc7kZrdnvvwo2zdnx+FXyD6QceR1wBsf9SyS87TggzUSj/MlK
MT9LGHRchfED8N78fMyCJTvt2dyKTVwmdDdzAp4v45enRRQxTHIQVk6tJBTJLCx5EXeh15zqArJj
A4yYI0rN/Elz757nvQUgE1iA4x20gVkR5Ehxi+v+TEI7RmiEcWSnqp5/GRl+bB47MAzfBVqrcHQI
obfH4NNmOmoKb1xOLsaliu5YMangE6YDPj/KegDqupX757itRGkO68RKpmoXzRccdwK0d8iAVGh5
+OPcyX4Q5wcrmtTy8U5vmQuHhGisPxAouN3CRd6mxFaXHSMh8YTOHx/bcNCj6UnjlREqMEUxt//g
vZvOZNAufvKLN4kHo27WjP9KQShmOn0vBf7gkl17JomFVt1dXgK8e/aR1JGN0ABxH9AQg5NSvK+o
Q9qD8u8GcO3RJHxcFRimUHyaxqZFOveG34eSI8ZaUWvYoyAwk/PJSMwrmtGTcmHnJbiF7kQcjNSE
RuzBdZYJ0dHwkAEf8fFli3OHuyIKuL7gATwsah6MkoVOmCb8ehYojX0r53/Mkvr+QQU/q2CzvtFi
0ytInIj0tbTRpR6uyHrm7n0+nnvlHPC0Te/msrH4eYIIJNv8gqRE0lXYLf6e1PXcN3qxfsXI9fQf
PIbleR6QGpYUeyCiiAJQGyoqgqyfk9HAZm874CvEU/r2Mom75lQ29ob8RotDvMH7JSHBiMwKfwNL
c2128dzSt9GSiU0b6Zg/MX+cT5RahTUxSZ492mGACjuThgC5PwQpd+c+CO6ktnqPWQIL9LfGEEOB
eZju8bcFcqviwSgrjmc8EEpwQJRj8KiEj5hoHFG0X+DCCfa++VSe/ojqkhnAFZi4+yesYMOg+UPt
9jBVagtxgJBxtY7tCJ4ecMFVNhZP5YPM3xL2nu7P9YpBvgUhuAC+jRIhzpx9l+UHm/RtMjdgbFUT
8MWev1Annjw5IyKw0zWyt5W3daLPGNm6hln35pUMzyhp7SL8QQ12Y7y5Gf4CrsVecTNHUpxwGFBO
cJ9uGVT1cnMpOlTnxH5+DDEkGufaRvD9XtmunSgabsrhwuc7UWeE/i2HrRtfV/7VExVJ4EnP5yF3
6HB05CNGidoKZ1qARSKZ++ueEqecf/5OEtu7PWJU0asFhtaanIXO4HY95kcI+hnktJqsEiQkFiGC
BFOArOTDigbrqSk1Q0MM4Sfe+zVRk5qXWWvj4VHi7Q5MiWqvolHc7Jn9RiDxyLZF/l+fv2dx0yXu
cpXWk69pqV2Ebh2M4K2pX+3b3OwYhOUkoKeAa1Gfw/nr5n0HEGmVtOBsXVvQquZ01njbKgnr4UT6
vW0c6iRFqKG9dgGHXdwdeKGN65MzsELZzg83wECsOhkGRTommeINNMJT2Lp86+QrTjIKEktHzZow
nSSuZ+EVzXQTMwBd3MhHF1l51hylf/zGUcnzf3TIs4S2EGjJZmE0NuxZBziTnyqQxYLxaQS5AkNl
wbZc4mftaTBgv5EHLEXhpi567Hxf8ZVwhnJSyiUbndz/MAjrnm1jiPNHoAo6cDRsmW2LXt6OULCo
qjMYG1CWvBiWfyqMrISaPyE9csSThaxxkFKjvgUS7GuUxaA++OwSr88BA1JpbbdpjJY91l3ot/Ym
4U+XTsxYzWRAAUuSc60I5pa5cxQSsit9rolEI1JpE/EhqLvexW494OV32M7XiXKxEnQos6YJguKH
zMa4aRSonajM7YsDdZJFSDHd8gqU4cuFIf94LbFjK8MZuqBRFlorNwBIzuib/wiKQ0UHvUooa1wI
HJZvdgVq+08wofTcUfWTjGKzFoY2oJAnhBBCm3kbmNWQpHQp4mboxWNmuv2E1/QVG70Kf1wfcQmV
m/TvQUEdomkiO3tboMTmJ350vmDljydPxPidAMsJ2WOq95gq2XrA9NXXCmE12BDA1LWIScFtAaFx
crM2BPchkrfwkUe1FT9V7og22jFFQOBSaF4x5G1ZALrvQk7VR9+XgbmMmpAGk9v6ibTYmwHz3lAi
mKrEURj2a7bVIT3QJ+UbNoae4l3Q8eF8xlGhjznWtSFnM8Y5hVz8jsobDQRzBo53pxOxXeZhJXHQ
dJSDMRDOIiMwl/BAMqdwI1ViLjCPZBIsI6LLw32fUrRA3WkyS7aQheHU52Gx0Z120QoLsNzZ/1eQ
u4/jcjaWMqfXgTlksKbSRaMf/dsAads4FiS4CueCwih88ResuyK/kpboy6eHnLa0zUPb5SD/Z3L7
f2UnWLf5g6prV0Mz9zjoa6sTRJe1koQtlQ3wPwd3Ny+W54T7WKhJSKM4WiqUpHdAJCVWPWJwqPob
aee/RONoLxdoxKq2zucfFPjtMaJ8bkvLbkfl00b45DmUTGYDXI9dSvDSIKNnbYb/Ro3IPuNNPqqf
VFzXoTH665RZjyuN3aobBStPm9yTn511acd5Z2jp2pcCzCaaeoD8IzcGHU+kc2HgNdPqVr8dcJIt
7ZGmgN+tMh9uyrKa07BrQSyeqFX7kTB3rcI31qsDs0LbyDcBrUMDgGvfwgaQpvFENQ3XnJeHU4Gj
5MLjOnNEH53+8p93qTUjhrCkNEWxl23NIpIAGUYnNvLJ6fca1rZvNOpYi8WfV/i/UXa1S4kLbQE6
gWIECyYXeuQ6CmhHe86UOan35W8BemCV/28uHHHKMxjovLxUDgli4aKb82dXfVS5Bc0qP4vnARk8
KwaZp5gaSlGBvrpjd3vF5xjN853QYkgjOveAbDrUBO4OwtSbKqJhf7UJSSa+3JE9eomB20supKRC
wHTItlDfgexI3qvqeFwZNPs31VfI39v4AXXgDsYTW+X699VCjT9Nr4u/qibWOPxHtn6hS6vvlVg1
Wz6N0x5YB/GJViOlfJoYBQIOAa7qH15rsMR1yBK3GTFQOpPUyY0/H7c4ywBDLBHQoo8EfbuuhuZX
sdkUSB61JUHZA7NXHSTpvKJnWWJka7NfIDrdim3rMpRUBMBkfLfc6mmH2HidnZGR+hSEpoALwt7v
TqDGXKWuZrR1yMpbpVmWMDDWv6eFthCxL9cH8W0W7tgwy59hXf1Hi7xt+x117kdYxRkccSCTuOcO
XiyGtIz7YboXpmK5LcVNxQYWWqvj2EfthOEUGaK7HXnmEhvwqm/r3RlTriHKefrtFhBNaLIjjO3e
oJlgb60mHhyZKxJrclfD1Ot2Cv3KpJcmOgWjlJZjKyLbLUDQvn6qSphp2ZpsiRBN2V6W6pfG9jiC
d2fgaKLsUQ5+KFJJTph8Mbdej8+fZu6BbM6AXkolEHbHFUAEJhITpdF3UwvxSu4CgHMKo54Zkbw8
YXMBVomdj2RfQK+a61wpgedwvCokVdNkWiunIQGzKykv/giDnCksW72n1BAkuS16pRXfL7LfyVr0
bgE8Iiq/4OF6zGfG3v3D2IA95X3YuiRXWnQ3WBVSIT0kQaAZUg/FYW9nnuDbzDSs9edekMK3z8C/
hTaXs5jZtIcmlc4zToCTm9hI3Bcn2KpIJGyXvuOZCZ9NsmlEICKQp7BTA3gPjpotOzogIr4aHjKR
V4jafGjzGj+i7CJ2KWqU+CskPdXe/an4EAmY75wYsBGvnM25hIhCqL1zGQt811BEeyAJnSptoiFz
iKAMhrr/lgFDJ8GhyHO16T5NHr9zPgLxPQJp4Nf7r170sdRcAwp3LBCRxmuxHiy17TQoZmyNJAHy
9F3r6b4p40yydotPrjWHJuEZilWPs60jHCvI7HEfgZrId3aiqYsjYzcR+dbS1wR26KPUnUtf94tY
15nAn9EntGPZ8rgDTmDJ8Yt5Fr2a+yBttOgqDHjdYJ+eYxq9BiF/OtqplzMPTMyoaGVEGbDcl+YZ
etp7zhl3VR8i9mRFx2EHtz0Bc/zWN1nodkBlCnojrA3v11/69/rfbnBDK+R4rwm+ZqClqwyXwXlQ
DizOa+/ZBC0+t3BE7mg0BQ4LwuN7dA8UKb+p05NfE11jSXrlZ/bOIJejq1AcNDvhb4DsfKs5ss41
f2riE1PN9lmIo5QJrLc25mQLDqnYHKDLB89YfZ3VRIZRKwg27CfSMpYZFl5ZXJxcImIcHb/JvHUU
fzujBPuuYpRgvO3g3faSesOvdX1fHIr1cGjGejv2JFKp6fm9b9joqLkJlMsc3gM/JX/0sKlwIqze
S3UC5x51/kL/y0ngT5Az5xjVifjch5wnnOloFa2ixi4am2bmF7ru4/l1FE5iFCbRG4HCJ7v9s5Oc
mRvz9GXUwYZ0lzkexHw1BaxzUNXso5KTTAAmgsYS/IeDHzWQyrwprPPyOdBxYZcoX3GekcEjNR6V
1xUwQW4J5iOqc3O5hqotcRJHS1NYb67C3TM/KqszA8y9eg/vbCSudjimQYOts3NvuERcFIlvXB88
PokxCzM3ahiJ+D0/VQRK43xJYDUfIwo6rt4K+c/0O6oWS+km2fBqIUB0MKmlNYJKJwvqA8TOlHww
rLrpvnCYnfD/eo9blH11hhd5mqHU0ySdxrSaNdiRtfcYI7e3j/2GnSnFWGgUT9PXZaXVrFxKmEJ5
rabZCfkWxCmUAIkgXG3oWhrfohZd1bVzHCqsM91Qoa7tOsUqLtZQFuqHLkBEXi0y5+sMmENpQ5t8
zHMvRkKhC/mFag3H2iqey1m8AkuWlmklUKZ7eUieKwCA6Vk7fP81VZz4N1L/R6LEFyK8OMdJsfyL
6yGRyHCcMTLET2bVd7upa4KbWp5eaPpTfxNNUlWgz+zoCwhqnBrDJDkF0Ce6KkXh1aP7Se+grKtv
uNqxBxPWTByeRTUZBl4rc3cuKgNAZAtfvzeOCZzOXkAXlujkYQQrXMHRoAHxUGVCQhKLDdEUGYCX
O8HH/rinAH8aGZ0F/TiTykO3YlK5pHoM9aoETpLyAQcRknzsyX0g2dErQSKGna2NmSZeSij6K6Bg
X+IlpVeYil+vcrrZ0tLcPAydnQ+nrpb+HYQbQlO4CgUqW+AuqLJBgJCJ3I1NEBbfHJOZV7eI33Db
VKe4U7Fj37KHyyBORPJxQ1F/Vng22/BTgi25hu7tGH3qAXFkFFNFUqpyaodHmJrKW1ndznQLD9p1
N80mgfBZbddgXdr6BpVHAf/zwDd36eY1PF2k0luGmr3RZ5vf+RVng+zIkSJDRd85bj4MVobx/GOY
M2/z490sqpyn8/4dLJhC0X4ZiefmYWmWum4SzrFMP7qzLzrR98KJt27rJRzW86b6O7g1IypwIdsZ
u5XMvzF37QTqXBPg6FKj4JvW9Py3k8GNRzzqzhHHZ2toU2YEEX4CzKoMstSCHuhQ5v1NSVSEejgP
57kAUaraBrNO9pAGk4rCjO4/r6PfG3c+I3yybwTfHD7fHL+5kBbNMQJnTCygYaF8l1HXQeT7m/6M
D22gwOj5Bf9q3TifRpfGIO/5yJFjNHXmL7JAcKjpak+wfZFrtVsRwPOnjylTaFlWCFhqZaml/hb5
fW8Ap/gA4DE9djPIGOwxMLvRC/be9Q9bjqqKMEN9tIiQGoY9+mP67o3+25KObRKGXzixHYbgUK5O
jhtwDbuNHozbeM7EfArxopprL7bvOUGlZ+j9Dft1Oq7lCjZYG1p9qy+xhWnPzQ+Ed6gQzo7AKAH3
xIEFbpkiK1w1mTc0FNobVIjNHGQvXqBhcXlwmu5W98EqxSH8Ma+LHLOEF++lzLWlgPsIqmO7/uYD
b6WpS1tcuNWUriq6MPb6i23OQM5+uRgyo2eS8wufqRDc9OSYcf12q8z+6XDOk5HdkjECJCI51wul
YeWQjYI9ZEBFh+7SdYIFbDrsiI1q+TmELM4vMFV1u0Wgj8UUUwYDqJHzNP9qtnXf7CooNtHjxC3I
G/lUZSX+Di+AIQaY5sf7FiqKgPd1d2v+P9jd1GrrZ0hSLf6IhB4DuuMPYEx0Nm9wMks6HddImK7g
7Xr51pSiOuvRK2ZWS65TYAgZZ2klatCFHjVtsE5awu3R23Piv0n2bSq4tJBnR+UzaZJWZdJTflLm
SqXrQuMpUwOFLQbM1bU9ZDwuUDO5/MH2EP9YfWD8vICtEJCh14P8dZWkb1xk8hDWAYpDo0BnavXq
sAG68dJj5E/2bT/VeGeBlZV4P7nkC3eg/z7Bpw3lCINf0yrjBfUZ2zFzgkXKZ6l+7JpIikegjQoN
VhxrdDpZ41062IGijDwx9lsg1dObSwgVIN5n5K9wSEQZknZtU4zVN0iarsv+yTRK/qRqzXq7A1qp
rw2TXN+oXWTl8ZCGmu4QAn0xX4m/4Qj0jx+Q+E3glX+6insIz6c3xxuj1xfkE/bG+IaLuFn+O50/
T6Qtm3F203XJNWE07a6JZ1Ur+RnGtbcX0SBL2x65nbeZzmObIfC6ZGvfMFDIgPVuSuJumpYD7MIw
4bvevhW2jB8fSTmWr6nx+JrXXTsYHawuKbxPRBQKzj7W5d5k2Iy0Ix/ygsXVuYl466Qr8FaCt9Yi
lRSMHX5YfrHN8VpvUauAaOOyYt8KXdzGFinhfBjog/e/h2US3pwbOFurYB7gZQWVK5M6nOTU9d3H
Q7fe4l5c/rbdUQ4RjEb6r5COE25VFHt0wMOIhC+HUsucKjp5WbXDpgeD/My4VCpz9LUgHQe+f8nF
L+MAXiIzJA9otttxeEqzijvaLxal/nJkRJLYLfj3apmrsV6bVxIPGoiG11sDcXmwf8yqDQ6t6xq6
t8PgFjn4tzi3rzWZOzxa+ISMXb/JyqN7ShTyEdqFxqJz8ZUApgxqJymnPtDajZTqvUIds8bNy5iF
8iYMAIZrK+QyQyrN4Lya9kvDYIVTE9X7yZwnJea0wB9fYIkiVks4oMmYJFahJaPnXd683Txp6455
N3VmQhLUn/pqWfOza8XK4PBj9mkqy1/uRCxFNiPy65LHioqwsCxxXmkhz/n8lngr/n0Kkx9qklvu
Ha6z0lNz0ysuXSSIkMrp1InDAp7HeGKNhOe67A7QwSu/ErjqpXQZh2jZIY0xENRLS0PLPFO9V3KW
S1tlI7o9pvPdrRGi0hdvcPFfhwhthODLdQtp3QUddNs7H54tfoq7x267J7RbujcqPl2DI39iYw+0
qhuEFze2gaVPjxRf6nC3goI4TVZb7lMvCvFkkUHf3sQaQQ0c6IpYH0yebVDphxEZNa2/MuCE0kGJ
Kfdm+3QzwP0DvWkSlpeOdxTCrmmjQiD3OkZSd8AnFU0RCfeSin8hYo+24H3wAuEgvObT+6BTH1JB
51fqNYmss7WZsidGHZbFgf6zB3H/p19WiBwK1rQbcY734KKMMj+IReHaW5LdW85m1u6aYmQuERpu
EJ2lybeNenkNYiFXYLVkaqjicvlxku8JtFfJ+ZCPMzkVxHOEa3CPYDwbNg5Qj3rW5Mxfp/uImQqP
7psQ3YGSohsfQ5e1u28u1UBDvRq/gIwYyLyRE/xOkbD+TrVpxNAhlWL3WEbgnUg5ggCQm1H8RWxd
Cdm8arJWFh3iLmBDnioMp+x6FEBSeOrjacRuEfWKItLMlQJjXZzaQVR9FCA/L2NN6N+fqIhT9akN
fHOrjd87mqbXpeJ/BegT8IHpJrtNeg9cuSkHvvE2HdOG1H4seP+3duwdVm2tcCwjVuW+ECBrydwc
CkI22StjIwx7mTZ5BN/gqajjj8Trm5zJEUG4vG1hWLQJOBQaIsrA4hcDg1/ndUIXF99m7R6K5j2/
ViqARpPCyBxJoPKPMUwY1zs6aRDnp9ODBCkjRUiZPr84Wez400wtlF/4WvirnY+ky5hy4MI2gv8c
qFzR8p/yvxASeycrLuapNofIVFkPpupWMIQ2chO0Eu2BjnQ8ZKhgLNl9IKHSDbgTj7hYeDZXrY5R
z3ymis0U3wlTF6dlOALmfXzERln00L01tMt6fWoDjXT1UNEq85XCZdphUjyOOpwLAyWC2U3qpmIs
IlFCvjGYxlao8faW+yzFEgsLIECr+xxxL6dgJ62Lupp9Yorn7wLdV+spfXm5BKqiIqsBTye7OY7Z
YfkKrQlxijzpfyUjwr7Z5unSWr1nV+VSeFuTHZQ2EFCCi7OGHK1GplYK0UFxF9IyIWXbyXAEhuoK
V1UTfqjpLr61DCpW1PVVuK7o+ls7R8IZUG/02J7rHb8F+GUMEsKp6igFWj06gkF5D6fMeyl4Kyvf
AffH8/GCdjcaSsjtFSwD5ozO5/62ublisrX8/kIq1or2oWCAZlTLjD1Mr41z1k2cXl0etmItemn5
mP/WORUl0BzGhqFJBQDM2aU2NOaqmyryNAqqtL59s+2MLE+Tzw9ZHsRAIFRtg4xu8M6s2t358wz3
RSi9yJYv+n4xNXDjqirOj6dZ/TCmibCpMqJA54wL7zZvCgVl6zWr74ZNtBg88QP8yeTygOWOsF3b
/Xih4j3OyQC3ZN97fXxzg/XDKJag5QEU1DWGbplQR7Se0ap1PNs10daPbLvbddNodEW0D5VvgMMC
dKRJv1FtozkhPhdtYjYQfyV2UUEpGhaWtIW1tR3ILP8Q/b+Y5e2G0dhnHoVXUvYIf1Mh51MYXwtx
WzVwta/DiETBFqNoeeALk4u1c9yIGdm2kyZYkNOA/FdDGm7ISuGr2q6QJnSMIea+TkSzZud+Pr8M
Gct9w6EL8UQFvFLqu/yvv9wQlv4Hv/2lleL9t7pE7MM/u0YJWS1w/L9dS3ABMhbZeyO+L5MIdePs
Zwr975dG4yAuu/i/7z3xZGBTA2yAz1netXNiP76V2cg62gZMpNwEs6JHMmlAy2cICsQDY1rIz9vB
mednLtTCByDXO6jfeLBFHioPkYcPKHpikOLEVxPsyHg8XltyA2wd5c3lkwy2abLBpLGAU/EXyWOh
OxUYNu6uMTr2qIvXyTt77RmQfwzd2m/lRxSZiNjvxAvMKgRB5pHtxBAVd+kQ3y7l2TOEPBxbO6Ea
fKHy/T6NmFtNzVZxfTGbRP8maM9y347/Da3IW9mG72ST2TwBcevSngba+cyh1+o3ahGALavLZYr8
gyApSYtRCuvkQL5MAuePqgSKWk4eRAj15iF/7uRDSYI9ieoYLT0RsaRlF45yBl6uq3KHKFZ1N1pS
rUg6Ig+E5sMjSylQu1GfOObBLu/kaMExMOZkAShKOtodrLnjGeuYCZbgENWjRSiK/7JpK3fJW8Go
Qk6Jm9AIM9/GL1SDL8xMcw2fd2HBKWfweoDpv+74ndrQujvITRvGdFuhIsTcY6GPFdlGpkLzOSLH
qE5h1X/K6d0DD5KWNklz3tgALvU7md1hIhJK+COQWUfNylgW3Vg5EvPo/UllegzM/khc3yCWqS8B
yM16zGO/ql3f+3ZKwQSFqeLk8WBa+KfDVsNaHgMhWbKjw/oVk6mCMe9PQjQAu0cjYN4jgNQ+2hZp
WaE9OHrNwCN2WZ/7zskGwokeEfmuuvKHCl876RqAOe4pJNzvAEMZOB8gd/iruiGPg5lmpzc4QdN/
q2aRUUQbkSVd6KC4TD4zDijRMHuA/N1kdCi8YvTmiisWKZtlb2B9T1jqqVm7ZtE88CTObqAeUsvB
OY9e1MK1WTOUWQfU3fMOsoIZDri1ycjs8ohRczwiN8UWIlH70+wKJUyCimnTEVsmGK997jZ7kPKs
DoEN1/jltvpSeVtClTsr9lXBqHblOGeQw1lHYpQhjR5+90bFJF37En++sHI93AytmEPfkN6yCVNb
sfvRs67CCfcY2uU7GTAv5ba0KoOeI4xe9kta7xuXnaYeTNcbbd8cMgYqQEc/7jNhwo0XV29jsY1Q
chUOKkkG4mCHGkxV2uuJKxGHAfdHTcmy6tPFxV6XEmSgWWC4TUjywBXP2Q9/cePdodUPvkH7eacr
svwpuZjRH0tN7ulIyfdPfy3VoJTdB11DSVJtlx7UmF8ICn8A6LVYiqoV28rkkBm2JqqCt/o/LGxm
yg0euhYN5hO6oorEj9FK98iVok7vr5ukMyN2O3TTD+Da0eR9vktn7mi7bsIaVBF3GvLOd8okheGF
OC1VvNdoqivtwy5dC1cWATe6pShB9EO6r1omRMjZVhiHqwlvSMCnSY7G8PbrH62y58L2tmvkdmgV
8HEyf1DtmAD9hufnzRKwMfxkoRPoNetKjHvLftzNy1XvyRx0mNv5Pzf9P30D+N+mdwI2UfvqSqjd
6D2XeA/Q1XQQO+ynbPKdQKMATHouNceQp5xLY5Af88ssP537fqetBoGfDCq40AIah5gEbtfYhwW9
t1sQCsg2gsggqyRk9NPmXOrxO0OBBvvm3eBhSahnMCJE7yuIBa/IQEaGWP8W1XQoHsPnCgiqnLrg
GpS831SNY/GXOZELfLuhMEPhsIRMAuRmUi24rIerNj43qXMhZfXvTMzDaLm+eYKZXum5n7uvGWBZ
eP7fW3ItbZj3/ZIu3ank3PunL6YQZ+lSR3Do6nc/H6oFoNUMvJ38HS5XAAQ3XnuFf0mJ5UzRq8Q1
CsaOf6om56pwz/7y4KreM7B4V6cSo7vVbFXGN/SkyhoMe/Z22kHtz1zg3BAmjgTOUpzKlV2Eih6X
1dY++0yd0tY70bMtJRVae1QtSjw+kMcwo13A7UqDxnJcAlZRArUEy+dKyOky7OL05aCLN0OSA8Xr
OGc+E4BdBS5Geq43UZLTcHh4J70MF5rSAaZ7ZbcUj4j27yaf0a8Y3qcuISScN+YIqV+olL+wt9jC
ObBkas522qhCcV+YYIi/+/91H/xBG/CW5M5QQ4CsRxY0ZlIJ8Hr2GAkOeocESCGexemhlPTU6R3r
Yqky33xVjOcWsEyhIac8aRO6DvsE9uBxUXDack/BqH5ykqawHGTrtnwcIGm1Yflvq7qC8D/yyGVt
FktJLZRzvuT2R8enZ5ulnXp82/3z0HSyjP54z6H3uD26Q/p9Jcq/5x6sT1dKMaqJx9nW5ULd1uXD
ylzPUSXer0y1EAMmX/aQCB1xs2lionSY7ICbqR5nhbK5CggnZTLev05qm/Pr4GtuPZ+DHqjkYxaU
fbYjvzPqFtEFbTB39nX/EwVr19kK7uM2z+4/1wPEZYv+RtCkPenaX4Tc/xNm/EtkfvShuXweRXd8
LQPIWlojOAc5TPPDc1TNa/N7cbE+RccGwbN0HIYxgG9p1Up7GoSZde/r70YlLv1G6GXTg7aCHBpI
M3LE303ZY89LCVJ/95QGqPJlXMWBiBie05GRClV7Pwu1GItEly6FjZNJ3rPtWZRt6KxjarVFt98T
f3B2wOyaeofitfp0HKBybP88OCWJfhsgv0vbPvvr6cMwP8NQZTSsQvaaAs79zHrcHCbRTZygivR+
pG40DKPMNrSaEHIOCPLtmmEfoae8dYBFbhD4Pld5/CZNukpCmoSilIdxBBhzNAh9E8g3AcNtU5nA
srMvEpxE72eH2OPlZer0pe1FaUY/kdS6yfKEDdhUfHVrD23MrpSNmt9S0a/RtHBRzLIifytQB6ZT
cj4MEgsYiivApnOiW7TmCZGztKjM0Y7DWJesM6rQj5lev20W02LIiI8tmo+QB7pocTaBT4otgwBI
TJh1Qgd4ym8ol+rHWNLHWcaS/EBekVUvKp0arbwvwpad9N2EEZSq2Ul7SeWS/pj8QYCMjPMfJ6SB
/oOshRIrvCn0BKGXKSPKB31Y4tC06DtmKMMiiM31eKQtGM0zO8NasNDEy/bXb/85He315GOAXZUV
DWPgTFKdh6aqlM9NLY36cXKLVwwGlKiErKWnzyQqgFc4Cm5kJpYhxq7ahy6Wnta3D8+zECzmK58H
Mgof6BeziVtWRVYEkm0VFfogU7HLO7unuD2SA9Q2ahFQ5Pmx5iXcbyM4qBy3/b/1lLRkgyt2U+At
7FVU2+y8HLCDnFbwJ/iKo3TGBU+ifyZWjjzz/ot4VPwOtAippLcjTNxm1C0xISoXaPh+QWJtTWKZ
6zcwzvaE+2D+cheCbDQ0VsyPBJ9PIWPlaf/2Ry9aG1ba2aD4/V01RzLRDdREtQezvr6iG8Un5YBM
zqpUbJIIyHKwyQTRHMriuavldvaJmRDRmaq+B7TTGO1TFI7/jjwj/FCYUJJUuoUzixlOhwTQ6gNU
R6uO7rMi+HVeMfVz2diSftc0hK0Mp47L01rmvGV355Ev/JQMlP9n1gWaEqdCRttRLUwF75Y7wARr
kmr7emR04B2LqOi88cdHrzQ1kBXFg2pXLcixB5oHAREJG831jPaqk61H42sTzDZStPmI0bpcezcA
PiALXimvkoesBS20CKy0Y1kW9y0QDLvzVbPKDMY+6qvmJZZPjzjyvUrt2dvevy0fPZyRb+utdW0z
11At9NAJdpo42MxXbYRaunup8Aufd8XEHDQGTmjZVtaw2SKvNvaJxGc6rK/EleF9+aZRvl7E4iKY
vHjAJAv5yCs2mjEYsuyRTRWGcPdNn/nhVkVx+n+fhGw313Eu7GNfPP1rzrtgvUdftZYAatOHVQ6p
A5WoNhM5v34dVKUKvkyGPE8B8xEn0Sg9nUMkytxaEnlKlplLdRxqKUJ/opkDnPp1zTco5JR5qsd0
UbUO/Ks56HmussvbOm8zgz8n+KduzZ2xhwWlZMG+aZNVCH7K8a2392yGozAP3XyqQcvwn6MSE+6g
xNRVP9W86wLZ1xXlAHg+Z01bZC1yfPygSI/v3zAvvYh1jSYYEE1NdOMMoOtS+kvIhiS37Kj2PFH1
QIAOEwWXsnvE7OBL/mzs3Yw1rK8VFjr6NDKNkq7Gfl+yZA+e1BYKvQVb3MEoIlfO5YdS3ztoYcKq
Ojb6Rs/hmnAN6pimqvpfLcavM55EukppiEItI+iKe0jshAm8XG004kbYfp/LoPJEfyoioFdLOxNZ
nkaDqAZvNWtPPMQudeN6FJry2s2jtyUc4ZHOo1SbYxgxTKTyuZiuq2aIJRFhGM1lkHpO48GyvwzJ
sjf+Skw9SkOTdU3HlLLakrAtQUrmA4Tv8MBOS4IFDScLadECsygWepMFNzx7IRvp1eBPpGKjF4sI
kiUegnr86hCMvmo21lNpiZt+Uh5Gzt9C37qp2Ysv5nXxQiL/TYnZUVU9LhKd7ruJGz7jC0CoWEfY
CuLtitODsSPG+pLOsoz4YuZoo+vAy0wnQ9Hpd1so/ZDk4p1uAMjPn9CULE9/eu+AnZDoGYsapPBP
6FsFQ96WkceIlGVehePbXZErhqGqFlMF9eGsP5HceqQJq+A05b9VSHVgSFn/73IaorbAAOEvH1C4
KfpD8wIdd5YZribQu453Y/hMMXkPZSpWmhC37Kz6iX/N4ppdsficlg1+pOYzDA1sBYWXplRm7SJE
VqUmdu8CfvidiYvXIc6n4Em0GwqT3f5sr5eMlsde6mrAX/vzigOUyKn9lBZRuxTtC1acjPEF/ald
S7HiuqzTVF/2uj8rPcHp368FHL5gk0Myuzi4WAToHtLuIvCafNOZSwIsNCcVYAjXvdLEoOoIdrj1
oRKCugohzbSQpjcvFdM8fVtqx3RrBrCcafRQtmkKcojZWz85uR52lQGDcLplANHXrqhtxuOwCiHO
D1JIr88P3794wdwMRjLUoRf1bxrAAVJeFJRrnZtbCZB5/5gPOdPHCQfd1n+X7XjBIJvwmr+83M51
59SAecAslmxna6Qtp+OPCoJPofGpfG+ysUZSIdCQI4Hat61Ue7gMuclPNqlDf7wd7qX7Qj/Pmjab
pQ07HzTKvzzPe601tIMntTfmll82nG0X3lkA2Of0Jn/38d7/tUPwwsryUbtJ2MgdWzsDnIao8cEg
PqCo7ChcHSoaJtln1j81U5eV4qAVRce4W2beFPkipzZu+1Qh4ikaDMV123Tn58UvrQGWfsRLV6/o
RirqwvMza9VJQBRRTe2ssgHPoPrL0n1EHAgSmtR05NpWvJvAKqevhZvKIjtZ3GxPfCi/0EaBtgRQ
fzwJrpM0fRQqF4/ZViGF1J/X87V+Mx1PnI/EsQlrc1j72YL+JqkoqzDoMuO2AaUfiz6G58l6jFZ1
rKJYU8VMTYJ29dNZhdakz9rPlqIfgpXT5jhcCsRRbigaJc6lEVrMmU2hrIynnNFrmiCDEXbdw4Ih
LpSZV4jrmMFisU3t3l3YNhGi6wum9KnbcpRfNTKEec1QKEuqEEzlh8WqN9k2ZWBAb8XkKuLaCT0H
/lolkdQau0WF/gXFaA9ys+iWIxxJwGl9W5PSwYMWTrfjmQJv3dPRzxtugJ3zZY2bAAFbwzVhJNws
dFA+W/dTzXbZ5/j4M+EMZRyvbH8i9Dp7l8KdHJnw0uZYwCAciZ8LW3V7BGytVsR7SkOKT8b4tt8T
EPtJPli5ilxgoYsBpWT7zQrZyBKudP1C7gv7Cr2+9jPxXgnVr4Wf+6xShhyyID7SEcweQPqzLSv2
PKM6d/nLrC2Q68mPuUYPZ6wubM3SWHIjkiAeVs0m7qkyfPaEHQHSi5xud1twJgt+toJNcyU7d3E+
QWjHJScyszogEHuepmMDKc2czugOVuUtTaZb1ByQOUEVaZTqGlycnyLJI/FSiJg3pDKfGIA4+9a/
1+xqb3DP0MeD9y1FhvOnDt/j09wa1sGTNpeSXRuYDXZdvG5SKpXXZW1erSCduKyeszWRnFYOWgAC
yYBi+1evxzqrY7X+2AysooWGCbgsyKCl2uqdF73WICX45Txkm3MqCRjXgN61HoSqNeHUZ796lIPi
Bl6/Mi3qGlgbVt750HKcyuBh1kWdymGpZh8CkGLUvOB4OgklLP6Ge5dsUHFpl7uZsa+xNj9iJtiw
Qln0jXWxkMhAZDt8qVDwOfaaOfdbQXNm6HTbGxdKAE/X3RvGQQEyDxnQkgfpiwDncsoXIBonkdwP
hlas7gcw7X+LYDtNkoKjT9JLki4UnBMjxHrTyocZ/W2bvLz/JcFNU8p3d5ddXshpoUF2nYbPUj/w
WCYvOUeGvEC9C5wyMyVJZZYzhMRyAmJVSjl1E/woJR/6LdrlwOe3BV3XBDKvG5iVJRL8sS8ABa7U
Oakd7eOmLiBWSZXoAc+NJ2pj86/qHOplhqx7zQsFwSwBkELNQts5xzdqQTPTiu4VOJu71oyWzPIH
ShhjNSQPtXEt485sCereQHOQcF6PsYHBRE5kV35TYesgQkYL9I2K7UxySirS/D0GyMslNykALVux
OFLDpDQ/c9P4MNz9G6kX7eFAjFSEbDwpyVWGHzx69QK2itCUNXqVSiTI1195uTMaZmbk+yFPYxop
zbF2DXx7mIOJ336XhHXQpGDelgGV60R10lX1fD/KK48te3gG93rYPB9aU/az2aKcVJDsQl1M1b65
LxdcjYrBNbkfU12njfcMfZvO3uEnu5LWyyuoFp/Uhgl2pw+H/t8oYJc0nL/TsKkTYKnUA85JKpJ5
iVraEUzLz5v4Nx0N9GckPdZ3hHg6LYwMBvSxVnWp8Gh5AAKQnEsXU6nDvr2OmDv0AMB6Q2ke6TBp
GFQNydnVWpKiHTbIBrOcA3CPC3FAyyjEmF5gjIb2U/O4B9Xp6lnMHIpbDFxK7nhqE1qlClc5C/Zb
QeG/UYh29yy7JtoyPfjr+N5F+J+4+JT5wQh7Q+yt3Ibi4M67Eg5iPeHG9La+m2YqVsDFAm0vBMqS
EB98RXlWQq6NPzp/Uj/0cUjX1d1A+8J3YL/MWcZcfxf5/5ZsEgc+F2/oSRATQx2A71nNCoErGoK/
oVxxxJn9lsnfn7oSxeobefCGE7+vbEBFJPTD4quo5KvNZMDCiRgCb0NR3x7CvRZWZklEFqg67geU
CF61P6Pc6IcvYinRjSvwaIH8boFCyWOYB34spRwf72E2sr2GlwBA70pWgwtX4VQko/iVMaxAfFgo
oKJ9MMv2idMxTLKqWeqjkBb8OgyVRDR6wbnMhAKUIRpgghZ7g0yxZ5E0roXs29FKjgUkECIcDMGd
4Gr1lHQn/EUb65xbYBbUskD1LFMnugPhyZztpgEhEEfA6jiT7g2i3Prc71c7HG6cRHzS29WVC9Hk
PAVbpNTM88Biu3RitgmCk1AcPi3i/mKEq3xUsVVzhoVZQivw2NV+bRbyLBYwCa+qFhBZrgX0mScw
Qxo1IG6NGNHxKOsiRx/C1j2NhezumwormMcOsVH1GOexrpDTHmnS7OGfABO3Xk0jibYXv8YkTlzh
wTMly0gFOg8cnGOwupVEEB/u42BxY2tHZX66MJq5e1kZNdDKDoXwbFhi3ibVpfU/tfDztEpinIMc
Eozt+NequgBtls9U/BEM/t5CeNKXVpJ9RpNJtUD9Umk/Ji4SpBi/F6AxvLD5bRwAa8ygno4ndVh/
4dIxOABGEcIoRPPKFFBtLC7x9jL+daaXyk1TqxvjXZMlcZG1wKdXsIr9GMDweS+CpCtuIuj8O+WP
oAd/PYXOxNV2XrkAKFz0H+SDJhqMamvdtVbp8/PdpfuvK2WmSAyvoOzJDusizoZwHhMIhoxRXGnG
GIT3mKHxa7jXaI33r1yVcUg31umYqihZjkGqpY9tSTh7GE5lXXp1SprM75AaKk+EEa/IRGhLGqu5
Y5lT+W7dPT0MapuN/bdMQV7Aq/IizcG/ODtbX8rGH7mf1BjaiqL4XhYVnpN9pmYx1Q6gZMtJolzG
a5dSG8geGVZc7Ckg92b/WxkIyPSwXnzNdNl297HTPTGMU+wVwrwvWlNREg4gCbjZLgEkjiBGT8kq
T0QYGJClfKeXIee/WUyJmgjXNosK+NlqCxYQg14ga7f4QhtMu4fTY/ibd4xn10EK8RxxVQOoPZ0G
cCr4ufrEJ34dMKRqaUppKCwMqjboszqxw80TRDU7jQ1tXGC8ERiEEwozSf641Z7YOOY8zwpRTF3w
lbz+8WXOkLEaYQSh/OL0XlprTxlLaa8RLqOYR8FC9FTGLCrvDhCA+OZF1hlL3muPnNHQSXdeNOm3
BhFDRRJsQZzDLU2Q9KTmKVIeH2vUlMObJjvwHf0FJ/5fqO0oilENAPSztN8C6aIFio7gKD3xt89z
zttjayyiS0a1zEGqF8BKJ2NSdkBBGJNAM+1O2LyCtyJZT0DJ11GSdBRG7LFkWtXS1SqyrxODE5Br
XZ+bqmWDW0NeiQrnGjXmPvE08XvmpStTTfM8xgYXiRylVoYjqaMJScw4VbseZpI+8/VrI1fuwvs1
ydKjhUfDpGncEnF4xA+hXQlncQbML3jcSQFCaVkNcdvUOkb5PmQY30SSddtbe92tUTkTy2IrrzTI
Be1zXG4T0AF+U1PAlcro7On8ijxWxBHbTdJ4EkRd2HKwRQcbSNvWoG0Y0KKForye7lfcVPx0ndzH
0odpT05yU0D8yeR+ja9xErTq9WGE+LickDQpVhx7F0XlmxVvQzV4cX+6UIU6mJpkaeYR2+p0swXX
wNim0uxZpR5AsI3wkbz7PInZhFIT8ptZg4ukyYiHK4eE4tZtIy6pb/+LSGgZkkfF3gISEuUwaslB
K6Ib1MGMJtbHBsnzZvz4/IjEEKXcqQHyC2IHU6/8RJDIcUAgBnh5F13ijDT1LVtOM6c0pIDSYboc
Yyjei66L/uPp07xdgXTbKBCETLraFiWu0jc5AIDTRlNbrZ5uJXd9vjKTa0ZN7gr8Z9evM99tbIxV
m94AaLrPx5AMeds3bI56nFbeFFmdDyQ4VRUFpoNNMUSBjhupFjhi+iCVyEqTRBkDXu0z9UTC6D8t
+r8pRfzJ9kBYtRd/4GTWXjy9eMYnAYSNUuea4wANuzA79v7+LE8y6VxHe1YB4ra6wvfeJo28rGPh
AM69TX4TLWAHM/FKo5o7E44BU+e/2cRo5AZObAVesc2fEDaNmgUpIHqdGtvvffzDnWSLI8stUjvJ
mNXqazO26wvZvXy9Pa3FIMaYG3By1BTgaSUfQS5DaEfFc0U67V2ohwyj6Y8dHiWSbwXcpiY3NVIX
rGT68zUSctkcvIgFzEl/Bz+wT10yFE0j
`protect end_protected

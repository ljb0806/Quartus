-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GS36v9jA6SFFXjO5m/QaADPTUbOqt/YJQFaVF7ASwAJ/ybG5nm9F6XUijHUSbu/FHjmAGmEQ1yCa
wZH2S2i94sMvnLw4mX3n2Ejrm9yyqdSxoCu7j2H0Cf6WPnwPZmXx1RqOcziW3GAW3Q3wf/lwd3WJ
IQlixAV98T0TCQmZ7TcerJTovomWG6+Epe8wVbag9Q57NwTCRkZjGeeTDQKeZBVkqXUm93Uiw3pK
4c9xt9VzQmrQjNAYc7nVnNIj2Mxv2eZcesZujKKYzFfDfW1x5cqkLLfnCGqd67GPxBLG54nRZxKH
1bK7ZmnNCrdEqpSSVn5HPswjD49jXx3+cMRuuw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18160)
`protect data_block
YxBmBF9dni2P5afmA9/xR4HmbUTN0sG+Y5VhUnEQyd0X398JzX6trgDACy0UzajbCOgBMcuLwt4O
eTqFLpSdcLWnYWFohMBr+Fk8he/ciz/uwW+LOmQAI6q7qJeIg7JjnNX8URVoSUGRMgyzGMKAaTHY
BsR8oDlE4GMv4iscdIS2GhJr0Ools2EjvNkcxMUOA3o7GoXUmlfb8JzupSVtzHRLNZ/7z5pgUqj1
1LClrE8JgRyYp77kc3cPvZaczuec8vHQCgPYaHLJQgeBeQ4TqxCqTuRHg0S5l0LbBBl4aCJ1LH4V
26JHt+21kS0wECdIqmUFsBAivC2vyh9UUcf2RknpjOZ7VTUvDqCtnYgIcAaYSCMoJaH6QJP0pPwx
Wefk2Iq1XNPfnlU2yi9UCb/eh3cVL9XKMdICdEcrF+YTAwCiYOuX9SQmGYSUsXjgKNDGWEeca+Jl
xSc22j5fBTUhm57r8phsAQ0f7xt8+s/98dMyVeN2KLNf5hH9D5MGJw3YnZnsQSwD8PIY5i5CCiTm
VuGmQ+2GlpfIaezLx9ArE+l81pER6C7AHuVHz7hFsAKbmrkviwcQNMG+fAjWpyzk+OW5V7no3GP7
sJLl7m+xvlkj3AL8e/Wg35DGtSsy1LoWSlhRoRx8bx36txkGNQDRycsgT3LrgFo7Ll64UIMvJei8
1dSSyw7itGY670w9/aUGWT73obHNOCGsphUlnxsRxzLktd2R4X34k0IIPmjmuTDmxM2QHg8/BjNo
diF7u3Dq4Fqak4jW7w6lplhxcqmpUeZMMWO0Eqy29k+LIQdv5mqqUf3rdoGmJv3SGVIGiNtjNN5i
vpcXF4XJ20cye/nuGVAsGX/ZVGwunOLsOXTTouYbGlWMWcPaWhOvkyrvkUHULgggvjCLZ6J0rPpb
6db7NcJhvaCJ9FA1kMAAbPVTku7p1yMxC6hI7ZEtT5noBrBbq8w1ywtwkhQJgYnxDoMZoWAsb2mj
9ypbu+/mlMbomu/fqTbPGpfObA7u9xOQ+F/rNp0As/z4OKCAdadGXshZFHUEUAC3oJbffADKNG12
iCXBblM0qec8smL3XUYzufqpdYyH/OhgVYwnpycH4ZC8AQNjAUSbDuuh2QogV9BTyUw/rNbSpkc4
Ok4Pkai95DPPHTCOOpM6xi2Qv8F4CawFGgwdZ0AJVlSOT345vqmqT9+ct6G5AR7OI0j56fAWFmrs
/7w4dMKdEnZGfRXd8Ug8iuvyT8j5V+cZr1wLa4UH8y1LYhWqWUKfgBzkPnqdRHr/0dPKJyIF51g0
8qHUwjfZOKWkFV3328zs8yvffOhieDsYKC6P7m2cIXNSQvFet6jOnYkNSWDQqFEtxAz1eAGHp+ka
kUKWpkYcUTZFDK5WsC8R2v0iYgjDlXg7enYb20u9WQwJdlroxLlNTLF6Wt3LOgntTTfjk8qtD13C
YiMB34//4c6OGdUsNBn5m7Xa4NYGT9dj4EKkS5+84qEPr2BqBTUydYTLdhfAVxK+WCkkmGPeFqka
2z1eQuNwkFuRExwhWtEDyC/qoUIAdXE8wNOmxZsnlHVm86SvzDiRsTTXsIZPXZ9sy+pKcN2lfxTd
xBxrlsecNKPeGQqS7P72+r+sQ0KCVmZ0O0j0GO1LRbSgB+R+1wHH/s3EEwxQmF6mu5vNmuDzbD80
Ir7GsHyDKnvob7jpPMgyIiarFCCzHV9sTARIsjdQW6KF9TjQrYRVXf66IsxwG3ivImow9uf416Op
hJTvxdtPAVtSwEbnEoO0l30mtNrI3FbjhlzaE2dhfS3z7KksJPwW4vkR8wlJJZ2QTQoFWRrHyyUy
/2cIC/zQ02bsxNunjCnF2b6Cfn819TbXTfH2D6KjbGCWCDG6RDec5bDwYrDgMIR7nseWNOXbDbUS
S3YZUi1k2WzzqgzpkXK+h8y/78IQdO4VThjdPmVLAHAGYUTpigeLLoCQY3sjJhdun/yrusq70IE1
O7ksrKUWxJrl9evQGgleDh2Fyd5QgoVckeUC9luYsmG7/XRorapQYse46/N+C9gpPXTHFxmD5oDQ
8I9kn+yZ05lfSU2gNsz3QyE2AZRIBa1WCVzYCRpVZnlV4e2PoXKzP/xBolOp8+nn6DeW9Epw68XK
AjWxv8impu+1ZIFpmeGpDkQKoPPaniceERxrsMjJ7DPPB+UGE5ZCT4FIHHvE+G01qlixmeTbCovt
OS8UiwoD//WRDhznK8awzhSrJb0E5jyHqyOjyAM+a8cvx6gyX3KhkEqzaOLkwIm989AUTrmdE8aj
F2D/vh8xGaDh+ZH3RKVPadfUCxJT5MJ3zKUaoVv5++ZjhGAx+sG2+PuA63DYmp33y3eKz+XDjzN7
XPfh/KzL6S2OkfRBikNwD7cwJGqyXqTIh2yPNyKGJ6zwZEpGjTZkSKILGjOjXualgPZpfEFul5n3
O+6O+hwyIYkvZ8saByPb8+x1G5seJXMIFfJfRuMcZTP9aUY3N2zJkITg0GyLcAHsFc1+PMJ0mmAB
3SXGCMnzFXB9apFw/+vcS5ourt7Pk/E9KngMDPM6cc9bEDLfkEaKObHTjhN7wGu2XC2jYoXLcWsV
T7OeiHzu2EZw+gU2524T8yh4o7YPgbCvU3vdOZE25Whi+sh8ENl+IxXZP2F0MRGMl8r+C8PTh6ZP
8UpKxZmsTRnIrSxecaS/dwP8TFI9ADrOTDm973YGp+FvwQ4IIR1y+3HufHSdp7cBMy5rr3W1xYwZ
NJ5KFROrlkPW9sSeY8PlvuFGX2pMxbKuCFnUzZd+GnoXrVlpWclMvttEqPB1T5qPLImq7aBHjxV/
SJ7Ccb3z6hYSDRD5cBZ0GRsIJNvz2Ainz6ZflUDjLVzMwHh043Y7gkAr7h9x9qHuXWl2U7VOJm0q
T5ZD6rCTWVDTDofCdxkLbsYUsrvrQbDrXYgf7yLmvSitWthO3hxbzZhBFdmvefAln9AoHQgKeDAF
jyY84Y9UIjbABwkirusIcogqorrJLkyy/2ZDAfUuzOpGTrbVTohcleJYCQPfi20RhOkBItlayXh1
a6fDHBBSQOvF/TRcWq/+E9hG1t45pBWBYJSVN2N4YOB+VlbGGv90r7auAOhif4zFrCq3A85YizkF
gVkzXi9MhqJZ9cfgfbnmfXU4AisVDKfkSiFLnb/CQp1jML11sw94BDJQdVNGM2j7C1nSRccytSTs
Z77h+llvXM9J/bAys4oEE4+jMX0FM0JISJsmkEBxu9RDhEhkgPuV3O09OXJP+Y86AMpbTW4izQ31
3+C3N8P3tCAgCV0B1TPeN8gAoYGBgDJzfNwIEwdCzzq2eIkFqx7zqKpdimqNr0IaVO292FExd+I7
kAfFKgKs4UJgyP4FbkCWyAFQvBsGzAy26CKMX5VEjjTO3dZHD+DRiYG6g+XdIf59C5ZnpDt7gIXf
csJfGLCtkFmkDZUmeYo+WIxbaTQW475AWhr9TUFOaFdxFuov051Qyd2ypYGg53PXG4vZQf2Vj6A4
NYvZKaykmM3nbq+0J3V0kFq2je01G7faZ9VeSgYQ1DzWJfDzyXa0vx94QabAVmfKjG4myBejTLA5
4+Zs5cIWAm2p/z0FLqWYStJbxcXLUZDMUc6huLebmnKmZJwNjUkYbt8DSUmET20gCalMQ9Uz9dUX
tMdcanhXJtNFZBSQsj3VSwzDleQfPsXbn07H4YTbbNtLq5cocoUNOHaEuxe4hlciqyd5WFPIdd51
jMawag0OdkQ9szBwKsN6bjABTUGcoJu5EWOLL91+o+OAHAaMnbN6u3ofx64MXqQpN+mQiPTTxTMK
PBM2rsh2r8cOTDNE7b+OAm7kqW2Q0JdCFtTYy5dN0IM5Q2QLuLIi7wV61B9fZx/fkvenWunI480o
jamJwo2a2cnDQKfv7QcySwddU53/AlNhtjuhZbabyDHkVAOIZO9Exk4xAn3xJdzM2Bkd7ziXar/T
iUxh5sNyr6u7WTUmkbtzepNBsKnwK7K97fYf5yss5grjh2kPBpTdDIY3GJ4pJnaSd4ejHM2bAoBC
mRGIn54sBvwoyXQo8jNC16mfHu3gNShQS+vFlP4JonNoZlOSTrrL4U4LumS2cBPdFYsRXZFiGv5X
P84+gCU0/+vRCkE+4HrPILQrlhH4Eci+9e3lyLkBu/huY0m2MU94gsJ3zOQC/brlPMSh/IB2FzuL
cLFnCkXFdw1NFmUYs0ElnZbUholHJ28cgy+RIYu2abQwhtQgsAtgCKgplW8km5Nb8+bZkGgHHUnK
CPKWz3iqyu3BhCI/x9uPR1POub8iKSUCtTAIenDw6AoTt34i06bJbYJF82zsTRrDScsIppGHotZW
5O7DGPFkCzZfywFGBBRnUs5+OvxDmXOw50xMtTLuPBRh0zf0UhKPrYKNrKHm7LVbp1V2DFkWEjR4
RgZX17mFCiSg76MBTdEnTjmH8s0lK7URr6gKMdDwwAaYoi/GtF0psfYPl7OnT7Sc+R7ZYj2Aa2lg
1J1p3uh9JbDwc00hbX1828xgnTfs2HGG73F+qhpCiywPWxc6CO2bAZgE2XkMwih3tIoIjxSbgMf+
Fjdu4hkLpIfEZkNTM2pMBZ3zQB+2BZ/xisfuZa+0bqZ12OdmZXwnNvXgIJ3wkM7nIl3skbUUFGaI
StxHrJFRqs9+p/55d0WIkC45kQtnGk89uQIhmX/o0RtTtddqGp7fkgJS+Qltnyn5JZ2x0g+T6uPX
5zIBzKQlwyXVfAWraID7O6NXn4ss+fRkf4Y9popW90BaCjWsCv0TRFMzJkboiSirVD/n1UhVqZOB
AFI1S18X9q0uQ6RGa7Q5rbCqCpYQlgj1YaHB40SiHNSEsulCysekrVkzAnKO9Pca4FStUx2hvMFu
rZOw66cXeE3OPhce8dI3/aehftpMTSu7kxMUX0Upfq7s3I2tszPKd7HanjjTdX9LG2d3kSc1d6pW
eD/ISOUH5tHFBsXmp1qIUZPnYpOgwEkD23IltQm3+sGf3Bwp6M3bYz4qjovhpw4SBkY44uciMgGU
j+p/SSfICUgWP46zamP1tQd8paxCuvr50bGEOBH3iLWnh5M1eTm7xfGetF66GXPh02O14zfdTf14
vzNpvhLFP+iz6k58MvFwD8/6w71JxRUF22fLJnKz8vZp1iLIIyLVPcGn+VvLdg3gEYHJ7hj5MO3q
vYkwvfcH6Luo9Iw4Mgnu1QaeGDGGOAitK9rg9SwcZgmnqFI2508Mlkx8LljNeEelkg3/U8uoCOjd
ubCaVn9miPFS1A0xPTbrMhMWnFjKr63qpVMEcs6kRHF3EkQ6rCueS61ypMf080YwBmN3gjXRv6l2
gH39Qx8UBRpoKmaD8YnkbazP6GKklKMfQZlxw16Zg4utH1/EelN+Lx7JSx1/SJxr6NLgsqP3uVtL
kx3l/6Nm4aD6EE+P3ZJj/YVoSN/Spmgsy8lnpKoivfT6Z6apDZ8sfGh2s9CJQIk/35Fxvayq7VSK
q74snJC9sXTdt5xPk+TwZyFvjmvizQtx6j9C06gKSc4oBGr8Y0KrsFWBBS+3s24nGDdZ5MMFy9uL
0T5gG8GTn5VPJEc5J8FQSkW07ac9hOFSfYRb2ZcJXVoCQe2v1713of/0g65cxM/MiGFI1phX0dr9
V338uimQRVf3eT7FP0mS6wciyRmR3dPvKFvc0aB42+0jK34+JnG7G2VVuRHCks1cqzW/4OOxX/MM
R1148cMT+JdKXMW0W/7p1rfXwYgJ2S9QgU2PwyVq9CWeHdY3X/nQm5rYsG6n3gnzUqxYmVz3swRl
4led9u+5bTn2fwEPbH3BTmCSrf1Tfjpf8JW35gjGVJb8EpD3noytEFTuq4eauLRtJ22ivupZI/Ug
niMgRtUjpavv2r2dv6OQhaQEtwPqnn6tqHFscTcZUnOQQ1mLXwHiI3IfMZsoGNGqGg6PSfn1gqR8
R2A6hCySKcjuPbjTm34i+NLJ8gNxYuqPfr64pA96rFAHjghKs749qYRhG0nvlIPXW3BXGdjAFUgQ
5l+OpVwe2tT2qHyq7wp3yzofS/5eaF7t3F1B2lzQDEOCd7tAyQOIkXtmnPZyOQeVueUlq7DumJ/a
i7xA4pPhER1WBZhfu1LG91CRP4GYpBWp78mBHKVoUV/ePYIyn2AOh9f0/PgcP/0fcb3xFLRDjFOg
5rFNBLl32EhgMfvX4M5znhuV512mZvPTCZDY/lz9JenF5Yg4OLaOR2vuHXwmPVq0dYNr2NxaCagL
/yHZ4MiJRpvyV27QjP9WhGEkyr3DRVjIdDGk1tz9P18VcQIBmMjEmrCXKr/3jVO/mBNTi6d6ZF/M
/u7Vwx0t/RI91cCOvIixfxDSBIUfCVfmOg4fY5K3K3KlGfg+KwOR3tw23FBKQicqu47204uvA7/e
6zNhYfPGHabJJY5gK4+CNQB4j3LG+qd+DB5jia+1Q4L8PeHEtr47NwDS3gQNDLzaFor1+vBqns1Y
9XPSsKAopZrlRuStQCXk5+1fGnx/XjzPYkHZMzORZ/BuEN5YQhkJ79cZKy6J1Qmck2gjJqPWfixQ
KvC9ATI/oaeKUOOi7ca2DeCosyI5Gp/kxrtQc+D8WOXpfwQkc/cUXaXq2dPK/EheOtDaOHqg5FZU
GprrykR4n4L8Zl4xL0oBguyyHC3RnAtUdSavK1eagHz8HDaUz1N7a/L+DiSCxe6+8lQr01UCoBve
e291yplaN/oG4E7qUKC1AM3DbC24ZOYNbTG7GVua9maHeIvVC07oUnzJyERpSRwRQJVc+FoPvLdu
obbzhvsGg9U+5OUZJrphO+zW2C29TQybAKsO/tPlfhTcN5F1YCMq4dPrBtFU1e3P9DpOnqx7CnnH
eN6j7PLNfdKYCoth9YknRrCy9Zej/fAB1lJ8cRQLUEf8Luygwn7/PL8uYMLcAHnGzLUUmM0qltu4
++0Q5K3gaH4x/Ivs1SQxl9YpcbjLJmbdwzAouP1fjvIrAxj6gbmzeDUdWJgUvpQxabTPgDjKMUPG
BmMnXIfMpTt4odphy/EXGKggDbsmt/eZxbajN0SFulB6GHHnTl2//n8egSAbSkNP2hJVJiI3cBL8
X2JhAbYLC0eZe0xOQcWv+8yYk98ZtoFWvTjkwquzgGSwg/iZzCyJYJs22WOpY8FVcu6IO+7lPV+r
qEHmr1SriyBdtSmNd+63fRndytI3S012cmYZhYLyhjwIc0wJaj53IUCYPFIFhDJMOvw1/C4++nYN
W048hjUGu3HbxcgOG1/UGwAzoHxegql1+tJi5z+asvrbYZvGgubPcftjMLmD34XarVA/CvUQdvP6
B6MXNJ6+W3xYAFVWx6IdgjxD8qkGvwUl2UlCrndsbDOKztKVwVjOGei0eoL79aVsP56wG1tlnj/y
yMlf6bX0NGESEwPkcyY/1PdjNYb8OV9YK5t9Y5NTRN0Z8aY3wingLp+7DvQC1mh//KHkByxN6aEP
fNU60NI5wiJRuSfyJH9RK3Q0rSL0ihFK39W8IqSBNjtWLDFVLWyvFcAXiX16NfWLq0AhuQQd0r1O
7pSTQi1aefBsL/GsGxbKYQ7DtfB7veuLDyviay+emCz8OsYS8kR27esXZYtZ0B0wHQ20R2+yrybe
yaiPe3lWWMlp1t1X/g+E+VsFXSd24tFEC8ISBQ+tyAlGNf2Q/6+f3EEttp9nIwBysS40BX1aZlO+
qRoBmUkJgmL7SkNF3RhxLj/0itIvm6O0f0Kkv30PnNGKcAS+ngEvqfxlXwNL23xZKRNOZzPlTsvu
9meUszL29h7OSY7JCLjFqHQ52XfGPur30TJetYIJAbRNvnLbDsY/K9prIHzwSsHg1r15ZfdKOP9m
nMSgxWY9PSaIwCxju9sOW+kipfv9opYheOTy0+HiAqG3BuvoaB9QntwMg6DTAuus0dEW+kgNW+jl
MHdVW2jtnMICQoRFtINoyvPVVY0M03W9TCbdLBwHTa34X+yFHdLxirYt1ZR/u1S5sU6iFWssd8Ix
crtxbv3xnDSq7FA8w4P3NfkzbQ4iIpJI8U33R2VFbWqgv8qGWeLggWVjXvJINYW73W8oIDgajIta
x6ukv1tecdciDT7PRXmy87wUKjvHa/M3qzyaZex4Sai02BtP5WvUrHvcBG4pAqIV3VOFiVGe3yQg
slTkA8OM+8NrXJW1bC+HYdy45hkd5T04JgSUMZFWlI+f2jy7gG/bKh+cHEwDMKwO6UDDeWR7l3Qs
XnMmJSK3pLpFN1KJxmEp0JeAETkU3HpIouPS9d5TjzgiOP0QEJdkz0KjmW2qLoSoqfpUS/ddfKRk
HSgT/pfU5qRrQvXF5+Fom+bmtXV8k1IbLit0iF9rX5puJ01OTkTl63uxZNA7Y29tJIwsO7wgoorC
mGjfz9UAHRDvBP18/g33pYT+gVrX8o2mnl3fIdT9qWkmyQ5Ujw9Xwn5cf8czjDDlA0WGUn3zHuoV
+vdqvnpKeBZn8yta1meKEHCh7wE35uhhQRT71E0eXem7sFdHG7tm/gwUdgfjnoro4yJB9hqH+zvS
G+oKEVYEjMszIlz6ucBSMcXweRynWqxigySudpDEHh/ydpb5wrt9RPZuqXH65g0XcwuYWwIzKvVl
6HtjoEov+g9gkNB/C6wtR+UrxQKzPNnhDtcHSV36JRldJvKVj62q+UsXoNZXNXh0Uvik82vSoobA
CwAVNs84A+EMWXknuYBfJ2sDiurtB8y2ZsQjbFR594NxmNzPH0wSp8uwWJz462lSSn1xckmOo5Tn
LUD9yFYRHntmCipDwHG2Ph6N9A0Kzr6ECobqexPTcAs+siAo9eJC40rXg1LK2W2wKiy2+H5icsJ8
2nF0E7S7TJJR3V3R9xGBbO4kP+DA0UWsJ7+T5HLmVpBs17VSiJ7g/rbI8Sp6iUDe1IrBxPbdmmMs
qxmFUXyxO2otr6xRt85Vr9ePyAik952RPQDAEP5EENFl6JSNsYvJML9mHR7MxWsH+6E1VHBkbAYP
UQXxEnvzzG370Ai6vA9rT0z2noSUjreB8HazINSoREvXyZprgp2G5ioC4oLOYjDbyf70ES2qb/yM
kPyQbDpD0A3DtOf61KwZRnjJN2BFVvY6AtoibFP6lWU+WrrktLIwkNiovU/iaidC4Soo1GDZQ+eI
pfuWYJ2h+z/2K+u/PqviDu2oM2qEnjqnNwmrYiagEZ4qetv+7eVkdweBkBOaXl9TQKB2EHlNWj4t
2a6IZu79vvVNXLRqoo66oZxmOhAY7UGakOYUfCnb77MgMSZVq3BudHMJLuPBwINkfxQZn3tNaG3T
aEsngHxX3MJ/MfnwsTp0N169433STEmdiSEiCbp8PQns95N8ioJG4iNra7aDncwRELXLvD1DshJ9
mjc5JNDmOkkc/U8N47PjPVasJteAJYVZ9kqRuD57b3AP9apH/C0vMgvkaqCj0iYr3rRAhpKFbLLC
BUaRgPWqdLNmSJ3zuOSmFnvTr/FlYt/2wwi00lmRYZQxwpQCL/f2kA+IG8PFbRZFEqcFe91D6IMx
dRcL7ifLKh8QjVbtMEF0loDFlGSNYUwP75a7NbyS+Ev6XUDgN0kLPSxbzpTHr5vi5Cgk6slfR0XY
WFY1MiiISVL0obFDSez6CZQ9waUCRovxcfMwwowLrwDGbXHhj7eY2hMCfHpDcY2hwICI3RR63Tye
iJxEKC004lL7Rmjo6rkryicq/WpcM2XXTr5KFp0rV/qdHbyQdf+14Z7eSnmBEkPUctBLcPEZYZNr
G1wIquan3EIqdlPXR8MiA4CQTxTXaC53UXghZEeeQvQP0TG/Z2PhwBg7WyLIv+tSlSx2Ru85MyP3
JbnG6aLXX5mlDvSZ4rW7q6lk56yYFtmBoZ/fFW2CBsN7gcLiQ/gcArkK4sBx52xprS6SK/RaqqNx
6JQcf0HUKQ2Is8xOqJ8fgQDsUlJoFxzUPeVJlYAAOHRTf6hNlWpU3W/yWFc5V/9a+9yPf5A4Hx6z
6qiDTNAarEz4VS1Bclf9tpmmhM6UFIgX9nros2kV6HC3fTJZdqNSrVD6pzhMvR4kSv+swJn+84SD
sDtE6RIjmFf+WBkK6mf+RoYjvEfT3OG6XgD7DPGH1DR4JOJYJYu9qfuBRat45zDdy7zj6InhwQb/
69hD58hhXxbXELhNIjMix6J5caj+liFGt1fCIommfryizfNHWKGfUU6AF4+j3O4P6Qtq/89Zn24j
Kutzpz5IRJdc3UrzJVTt8HWfrUlJ+xYmoU/FfemqvqS+sYsoWIGoP6tLR+Er4uQiFyRhMIY9SNOR
8wBo+lyMflHunUo3ztKOEc0SrHDRo233QES7VLHML/SYiQn77yQQOSaMwDlVg+0sVM9XBq6uodIy
7vKE+OzeUacXqH2xqW0vmzkALTJO6fpKqGfnmLZr8+EyqeDT1GIbZ46o3C5FDuGYVfommcv9LIb1
kXOdQ6q5ac39vOPv39JLz8HT5GwzYGjlSPzhl1W7AnYcOSorDxoTjE4YwEFFWU6c7KJ95BmLa8OZ
WNzLYWPX/jO71h3L4Snfs5muuia9nwNn65W+t8SPu+dg77xZfDPq0jJ0zuUjh9y1o01irnrmHbcR
TqYEE+O2c7ve8Ij/+XZN9XNX0lSmSnkTugf5vMP1Punul2+HMCvDa9oTrQnvL4FnLNcF+kUyrYvk
ldfwg/hfeBx+oicOnoTEl8dO0YfOiTgTVyfY2VtEfL8x2Xo1YSt+wAIuPTJIrjif304W8O7Wp045
j6m+yQaInzNxh0sDbD7AmEDSvvXIaI6/yThMWAyhR23aAYyRY2yegvVu01WEBuN/V3yDfh0J6Tr4
LXCpzUZeE8wnwGXJ5mCfHL+GDvkYUrfNGLnhtg3cDvOIMCuUnCtaFjdMY3Kh+k9UxYyvoW29Ik9Q
Gnvt1iZDmFmgueUDx5aJsK4GIvtqVEQmA01dy7u4IE+o8NZWmDYptcWBtNQQARPOitRA+sAW/U5r
bEgKTZPwvqruH4xx6ZaIr6Ha6kIeSX63iayWwBo14eZTPo1h1OTkOrcaaBLuQefIBEOvNQs6khhF
5EwZh/P46eguwGhoKOncwixDY0W6RIw//qRL2bH6OFVXn984HA/nfq9MRffun32Rie1FyiUL4/oZ
DsTpgGqYIdQSJfL5YgalV+yHYylqcfRayCbDOeTbW6Wn7crbu4bFvMReLroMd+VRBJsWJzTt0DHC
Sw96TQFlu3VPvgpc+QQ2grlSo8LQWgeAzUUI3ri9kCDguHh9EaQcDzFobZzIAxjUeZum108DsG9w
dCZSWzC25cCSMHkh8v70Qns0PazJEhkDwUUIL5F72kHUG2S1nrXdzBauEcHCmruT6elAiktmTf6d
bgaYGheuGeTg9x3sFazE1uUpj2MsqXZgaBst8MriYq+m8KL2DcpxaExUpVrSq03J8kXbdHAy3taR
x/mtymcvp0geBiQDg7mBnlOctjvhTG+eKul4Q3GvzACjurTAnzBkMR0tFGzjKeldsjp11IiLHznY
8sISHRflo8PZeBX4rUC7MYVV+XqwLpwT5z3K2CJBkDSUzmst6/ZnDZB34nEYqHdVRLw65UMBR3En
oKozvAPw38iCDiTbe/8ujzvdEYzj4Z3B1qNrXkrRjhDU+CBY5N2vOrE2dPtEBchW5w6JjuuuoNUI
4dnyPsYURvMsOxid5uUYsAoZzFw/kEkdT2tFWooHfzpCuaCHJnkZsDB2BXpvfsqwHWRjdFsfG4L6
rkj04bePHLb+Yt+na7tgODbuHloKvAerMx/w74W5orVNlzHcRYBji58o1yz9VSJqetd3C2vH5u8J
UV87CrmMplXHfdLHpUwqlQ6VKqtefiI0rbqPLUtcffSTt/LnEt2JW2CyFDA1Qkq5IIMZQuQQwnVj
JE4hT/fTwAsWCVPKRvgui4vz3BpcMpnqSCigmW/O1TQpIwwlCjwcS/VsE9374Rw5bFVI2pPMPlbL
/icimHPv6EgOnq9IcHiBYV4meUv3j/zRvSmVrM0Zg0em5lYGMGM30HkMYlHsVoUFjf2ASllb4xfu
1k6FRUcJbVNZV2xmNifpVAefgsAnSE8TeQjThHcYuepZ1g6Vy5XeJkaJi47km0NptRGy88xRJUNM
WFCDJ+E0fzZeCHGxzI0wALNHv3dnDrkWI04K42gZF80wY7opJKgT13FRaWgqxuBF54W9cEm/MdkM
C5j5dZu68K3ZLP0yCjjSBRYPLvKSIYz80ezq/DywVcfV6DayvCmyjKfpCQ/zzh1FGO4zfSttmQXY
WQzJ3+S5fuok+MLAxt3v93DnGm3SKg9lULGIS6qX96r55JPFFuc6xavJrwd3Y3Y9B4gzEgypQ71U
Iqp0UxY5lbKBj/viiiEMLbvE9iga75ph3RpFxsS0DpgiIEod8gE3nmTEi+skELO1vQblFS3YvYY3
8LsH/Cp+H8suZwHLTLUo5vsZGxVCMrL9yEIfKxl6RHcfU/IY3xGWs76PqI7dCSsYiYA+PGL5nyLm
43y/GBGpsoIeyFY57g6QHUpmkLE6u2EMN84u/cSuK8bKPyUG5TUPpNRhsp98IfCRC1y8cmvNJC3x
eBnYJ24kPJNJZ2NAa+cZMZgnzc5foh2yPH5AYpvSyk1rE3x0XRy4QaZuZVATOnIZq/BWxnUXnw7g
FflLWkvX7KqcIG687Cswk8Ze0qFMmKRKMThfwTOQD3pQsUT9xXnCjHTKDrt6dsNr3xVmasq1+AG/
89A46FGu96HXuGeio49AdP5LuzaxG/ToPWkx7REc8akFn8CFnopet0e6NECgXCzHwXaT8TSvHE5M
dlSA7hNGmU3VcFWJkn5unWvJ48PNPhrpSIngPbaQ6mag7Ydu9qUvkqwg5q/U4pH8GAT5fonZGhZy
+ipdoyHe8cnv0i8cdio9bi10XL8cYWVs6SsdJPz1F1MieP2nRvVCgOPOfRuF4HrNHWkSXZQhAtl0
t014Wp5aiEkMlA7aeiaOAjopR8aYISOVLXfS4Qq/Vy6OlFUalqy9gmtypeQgeEsMbBSgbwy7dxaU
DTyCkjiLx5W3vU/EldG6uKIBEkezymWAQY0eQRex7YOwSjygUPMuHwdT14mE7bP8QfDiWkNN1r4F
uEU4LIba3lifZ4dDdMAd/rKpaFL6CXRi6yPPDy7MNtMpN31KufG4GdoDNFHQQLraOSgmY72Iq7EP
FasQGNtSvySllQwkKD2PpeYK2B91+bHjpYAS43xXyhjB/5cScZzwoTcD5MJ6cx/pV5fhZIqnMaq+
/kjZ9nJinV5mSYowTRcRX1/7QAWCP1/vuOImEA4B2DehIan8ZMQJN/oo6UH9eeEPqyIIfyIrRk8D
ocf7efTdCStt/54Cjo0HJf/aTmX6eeoJOw5CTAK9Y37il9ZnWEFIHmXQBk4XvLLV4QGi0tY5bqmp
ovtxaUqYv5z8YBZP8xwVYz8CbBhSRji2H/TQiQLL5+i9acYmkrBshPNLlVohayMdIgQLPzvGNJwm
rYY2bptCSEAO0/xYX/dr2/VG7FdQAX0vTeK++6CO/dDdjQfgBV28pz4nJinGtafcJXfVdMhO4xSN
z5wYlji1HkriqJmKllQMKFicIAt/p/u6m0PCAP7T6hDzcFqsTfZ3r5/iGu8dJ1K/J7PP7q8FnAsX
XQBwVftXnswsUzfGecUUMAISmDyby2WYMlgT5LUSyYiFmiLLDg2var6+7rJrFT2Bb/i7xfRlbKES
QPXtNTKXWQ4CYsWKKJ8HRGQk2lLf62qutNoo4JOtGm7GzfxNTP38T+W/S5vL+CilYK9zyaCiLclI
DxhZYa8B9NgAC6HJDavu8bDppteQIBXkuD5vkZoqoy8oc4KkvrGoanRV3WTvcvhiPtaKAgec0Ctb
+eXRqm52/ubQG4hrtPi6RlEjcu5nF8ydrIFLv48quLiaIcbshDADPNFSyhMQBxdNh4CCPj4AeUct
Bjfoa1LC45iOOWqjaHytz/Wuo3zdiVbZUvRYNHjivmdQadbxdw9JIOBSF6Dc439YYZB/LdOePqwr
cD5kBMAWACD5TUqSvCbjjBxEckENSbzkE+MCbSoXK1p+yvOgru7tHuNe55CkEPEdIqUEvqYf5z+w
lyqsxCMryjWL1+EkPy6vc580UM/XRToIAzqsAlSCBU6GO4eMI56Wz37PhtMLtSFzRyrF5TAPJxrv
74DTb/i97pt/6WJCjswbDuHr9USKbPH1W3Kp9cLJj8sYn77YRlbVn1sSqDdEejdKZM3nJkRYki+a
iN9QfCq/KRZM2R8grY3uEuUkS3wqFB0RXDHncWYcmTQ9SXqupf4OMkzkjaGvOAimkBpUZG+bhM2b
RW932iI0ClrvNU/CuGLSWgGT1ESOwQHA3MqsxfrfSxiZeTp//A5prfAbImdIXnb/zJv1Im/21Apv
WZL7hb2AC6c0P884/4OzX/tSaibEZbVyqvNv3GzDFxARzl9G7EpOFalGDaSOTliPW8o5/3MfXY+W
3cEdZOqPc4VkyR36JF06lxomMN21kScQlmyn6R0q3ipD2Hemmljfv37dVSLs0GQ1J5hdpmaoLzOJ
Ux0tr21AvYlJ+FFhkLP1goR75vnAZIfhOLNnihZxdsCfJkb/RCQTAV+Sd+9RJJZUGZ/Cy4w8pY/U
Pp388Kl8PsWwpqYEvhHpEuBk7R31ve/8W+ww28xMEgMVgLYgv0yQdmkEgl6XuYS8QEgvGLoNFLUM
WUW4LnWPa2OMq/sCXv0IFO+0G6rCcFXTTUdRhUD4DyAZFKV2SYnSb13CiVPupb5L9s2mfwF/mH/Y
LUitLcaUrn8/AyI1dGuiUWUKH6CsGnQJ0695Syf9S9e21xAVpu+7KFPzkt+Xf/1eyX4nKeUTIH9F
0MEPdabZewd8j148/bYzEZLDBI4d5PMTYq2NbGRah5PoYT4n3Tq8RJocbKeyqvCjffHAuTQZJkUe
RkevBLDBnckc10sh9Rz9Q65EtgykPi3WCC8xfxWX/GTzclCNWz72oJtbNoXpTzii0GaSS6V8KE9M
BvO1QGeKL4rCFB+f+9UQ1E7vIDGIgN8oUq3DVS3DqLRzlTqH8uXt1wPoED3t63JfARJqJ443p1Y7
kR8DaQSEZndnk0DSTHfqGmYV86Z4Jd7xNrpkPUGcnTHPV9sD6MZddYssW0u7M7fhluhpBSnkDIWF
d4h4qD7Jg013Ex15ikIF9ZeyNb6ePeay4ennZ01do6JVZvq/LPBik/N6MbwAw8oGcArf1vkSpFV7
owvfLCOnqSQpl2KqfNSuIu8FDlc37LueXKhbqi30Z5SjXwDd4ausmfYV021M3dbABx8z947++lg0
q825HO7pSrem5y3r66Kjtedr3x8IlngvfqhYwypUqjuMbt2ovXO1LevgNtKT3Od7Kr17G8aletz/
Y/pMfYFOZrlfikPXH9RkocvrRSA5YWGjeU7oZTAgv5Q00nAr5a0XWEodqf2XRDHbZ35XPEPpmgu7
xuL7POcRb80NdlRGVMVoCz7dQ1TeMQKfKWj1Dv2G9fGoFSB6xf2tlxgMNV6cZgQJhGUsfXXPmpGV
X8mLSLr/soe0lK0JdBnphS+7KHmF/kf1+1tkb41yzGe1J+PB5/C1XDy9g1kefbOPqyKjE/iA+FCl
Zw5zuRyEtwWP3zuYgFNJw+KKWa/7NxcfdztyCbBUvlh1BM40tCbVHfr5Cab7tNexDbotykLo+UMa
b6O8AbwjyiCmaUdCC5Lamjxt+q937H1hFDsaJQGG9bD7/0AM8RiP9myZG7lu0DL1hkaWoiAdwDgr
s04zeLfIH3++DZ/QmxEovcIsMfb2wVF/OhlXBMIB51RrfpIYI66N+1dO/bG0fmn1c1hWA47S2GYQ
OEpChc9MCY+CDeh3QGgqq7LEFWXz3NJmf9M7eMHBtrDJ+/c3+1TxTKNpn0NJoMR5zDwVjOi/NUnm
kQ865YvcikGlTVSf+78Mii/g1VZVFhs6qvE7SrNsl0lFzcmWJ8USysWemEaxGaelQng9cEZqGOLQ
LYAeD89gJIh1IuVANitfox5UBZe/vQeLjiCaaL27rVVbcdz5GTiqfpYa4rAkbhUK3ZcZ6UOMXmj4
seeSY6a97/D8a6OSRKCvXJFqV+KYwV8IhslJxRct+wLzS20nHRkKNr1tTtBq/jtzmTODO7p7lk0y
Sc2uPSBhrZQ34jjMoWS9tLAlbn1z2/cKkh4Oe7Idu4eIByC0GSqs7lXYctFZeflAN7JE9pG3aMot
AxU0simfaP2ESKMX/RciZ2pxBPceVUOLMQMihIOTg2OII4AtNeimlhSgDpCoDsMF6wmuCJeL2PkG
usVXvfuslw98J0JwjQ4VweHo+z9AxdwkDfqTNhRDpej4nDZimFL4MHuiPeqcT7BdUaGbAzU5lkEN
CHGPqc7sfUSKYSOj5Q6rwhmZ8roKvqpOR/ifu/9f7wJ623Mh+KqDlEBaMsg2lv9Ubf3kZEiohAtS
kwf9fy4FYARrmwMcReQDEj8mLdb8vli0uvll8v6UeziqA5xjfgfIW5TlmHOGL+V+rNoIr60zH0Nl
NANd8NEFqyRx7kzq+TetoBBT0rXPspSidJ7J9imoT8q0tVqPAohYCmcgAMWzYG7Dh0aVWM5A6ON2
3LihUwgGAw3GL2b+Sd1MQ9NAXOo2FHY9KkCO5q7+a1ybM2YfUL9JkqaH9GjkUZ6pIY6AJJ5uLQmF
EYxO0MOWixjlsvwzJksEKvOu1Tgs3qiYEtUZcx1VWwODf2VH2KFCU4VJB7+lrzwKG8eFyTD0z3Xx
uQr75QQxww981WHdrgxGjLse+cuyMUMc4j+6z7/HXZE4M4h7tw599dvDjFQuH1iReiUaMzOK94It
l+DBFZ78AUWHgWABE7Z7hiPMhJoS6dhqNynYrELol+c7F1tbfa/KboR4FJHpTtovXCeBV3yPLDK9
kVzLKxBbCy7ayqHd1B8IqWG5BdOlMIaH8LKYzxaZFNQdCZq4N2blCYq+FBRsfIl57BMtPhwMlkO4
lVtJvt18OSlZwqQyDtE4StWnGn74GNCSQv5BzEPXEMC7ea0ux8gDW/KMo1mgPm3CcDK6BbYs+EX6
aruXmn8jGei51Ed1I0GCD1+plntDXnwlk9mZBBVno5ii/MpKUyxe0ICSsNKEmAgb1EskZr87E0rW
/9NKiWOKXb6N0Oo3fvLMnCLLTiAZLIFwmIQPkA6L/56q/haoyfjkRkndFAgmW+WlRbTbEih39XzB
KkG42VlXWAPXYfVTo9sbYfh5jFK4iB24lv/zE8CP1tRHXZqiTnJu+qGamqVJsHvn/xh5TzVc6cfp
SeYTnsj27fHiPbLV9s2HHx8Jx9e7QoYAaZ4Yb1XKls69VzaK3GxhMeZCGGkpHd7g58urNmK5Y8iI
L/sajtsmYyezjf7CHaeEifveNS4Vqo46uEuVVsULDwA1ACffpJiJFWZX+2Cy/qEihyfdK67Fus0L
agfNsHAqizi34Stlwtu9vjjmzBYLA45Jwem7/AhqcTrpgjNvKs/oNDqETY2hD8Sv3S2ymPU6C1Nk
4L9LrWjz+WgtGjwj1vl9EdW1ng2ZFrztVhapSdn95WUoaRruQJ39JZyIv22IxM3P1SJE3mPVd4A6
GEmTJ3KNlub8mdaYzcHOCofSgDK+Eg2aBz90jS1uvKLqzT27a5z7jzAXqo01Hms2iRY+BM1I9XMD
/PUIji+k18mCFNMfKJ1aQX9FB9l1FdyURAwjMgYBHeHbFdt5FolO7YgEeUhXsMrR3HXobFLazsLi
myxEA8tYa4J3jfY5JwoNNc0TP8UUx8rdXUcRgFrncUISCpyYDT6/C3dBAB6cQZ+oynBgqkS/PN+W
8ekw2E9BA/h4VNrwVpyrGcysqWPD7nwzgCEctCHHfAbO7+FUKJiMnRuyg+AugmdS0giWGdJQWmSG
VpQIdSZwMrX6kIGMFdn+gPRLMVFdOY1YhtlQCibs6BB6A8dXJe1xZve/EIyyZ/7cQs3zFf8CL+pN
nTobAQKyPeDdrRLFES+s9gAIPiVDIqcyxMCQDHBHpAt72RI0Na+GEbhbWR53PK9QZ7CSA45DTtg5
VTmbhR7MjZQDGp/lvXaOQrwB011hSQ20hFvipMYdc+3IL0cCRwqUlczq5VWAvUIOrFMKM0J15i1H
xBJYiM3V6pz4NflAz2LoLEZZSCZI198ibB/LEaMJme97+1o5Wsjmf89lp8AhTlr7PQDOwAuN3JwA
OSHW9TdJVJfOI+vQa74xCGtfGSP/B4+HL+8Qtqddyji6YFhepw/r3Ai18kSZ4irlQQJ0ZttKCsA5
fpfKuJoh36VNwRkg88z/9oIlafRPfuj4ynUftlGnG7tw6ziPi5HP3gbs+j64cWzkZSCYJ9PCA6h8
nSCfuoI+xcMql/B7vvMDr9GYzlHTJcEGDlbpE1AJZZyb5g3NEfHwoPx1mIho9mhQBuMqZfWM1JJf
rha1F+/1BPRyd1Ly1jOHaJvlXj3laeMKEPuLaI1Yuv/JtpBLzXjgig2VJ+SHq9KUyFARRPG3pCAT
0l+s3WNrIu9sNiC580YeVFad8u5EGAgGRqav0zdBG2qMtB+iXQK/MVpktw4aSPJhJ275ho9s9l39
iWSNUtm+85g26vOP1ZN/7+2hiYL+BAXXYicV+9cJSp4cEdyvCkPsDcBhsWNEZMQcMwjqCQPH6P6o
UiV43V65u9CdCCp1YaMi3chKuFFzMVsOlXSCaevTuQBxvPMFQs+yRgbvYoNU76ZHpQCU/e7d2k2o
LfaI94nzj4G7m6hgVcd41PAOHJng81aN2RqN7vm4X/+f9wSqmaGMVktIEJM7pyeCUWtkjW1l2iIV
3BiaKABvbPiDr6LgE4gpJvd6OtCLA1b+V8/s9rajOlBJwmNBuQ48mT2fgF9DiS4VL8XWwVy4xsC6
tL3WezPnUvO9jQyjkh5qzSr6+NWv3o5oOyPkahfpraJMsbTi2qqJkGjZefaxPTfLceaWO//5QL64
w3nxyzw+Zv5LQCYc1li2ZQ0JV3wJUBDzYKlfeSlyBkvNQMGdHinmJGN9UsIcfPWgWVwxQ32BMPx3
lRCYKcKMlNCWKsvtAyLFs/UysV+BhuO4ufO1QCQpgk7w/hiRTTrvqOALlkYa7t4GNge6PnFcubjA
emoTyVw4XvlPRfWPAH0Crm6ikGAEj3xp6fq7kNYU70QMSqRCYOx6mMcKy5mcl5cmdaalyg75M2my
78gDb1e+Kw+6yiEAqiPdAjnrUBp8Uj6Pobz58sPVYRwd9NvM6yhjLjL+6GPMlVG9hNoaW1r69Fxa
ntlz5DJRm52fIiInMy5IkAoocf7xVTbBXByvi2/7q2qXbHTHiQ7KPDtaVnPmjoSb1Sh9bC7W36Hd
GcjADN9ks4RAYUiYeDw9hST8yffxIlbSDRvToKBPDGiywdyNTVlHhpUA40wq7pgE/UaXYW2rtw0L
dZwDmqWIRzdXZqzl8oB0iKfBBk35oLXhPWWQ/oFYFI0NJZkrusVjkeqyZ1KX5wWQg6PrDO1ssMfW
csdl+Qnt3A4WT71DMov/qVEjxzzHGu3mc/0yr4Iixmu4fD7k1Ku43oqfv/ZdNZAOebAnQvudflGL
VnY8w6liXOamrKqU/gNwUY/SR0NqBm02oZVGVEigMzPpoB9MUI5mT7wclWct+uWkgAJ05T9rOYd1
hNIcu4Ua+1BGY9y7tzowFsKXk0E+NlJFA9j2y4XhDMhK5tV3xhoESkdsrF2moeV0Du3+jdExSM30
B39uraJXEUaFTC+KGheYpT5e435cNkFzcDcUclVt41YIjmQVpdMzwLSrRGyI2QzzfImN3ECrgrfb
PIpaZ3bU7qEibBwQ9ZRjpHDLja8Mz4Trnd2jh8e80TbkYycpQz8Nd//E09r2aXBz3x+4jOTY9Mca
oVakf1lOqzCgmdKsBx1VXcKbN/MZOFyztg4m/NSUfIuYqcksuigpgHEKpbBrf3xvitp+esAhpMKF
wkTo4iHCbsZMJVFW+XNVp5XZToDqfyZyQYdOYddBtyplPbeG5X7vo6tXRfVDnyB5uhHOviNEAh4O
0odaJ+XryGpjFQGXYuZhpWcVVofe3+D8Q75mrIh/Rdnc8aW5raUJRYXdG8X2yXKP19JIyRauwnd1
c7lT4/F1nEW6gL7lnNx2uc18iirif8zd/9qq3kAxwaXp+z4obpkVTIs7Yn3DJUricTO3XztEvIkI
y85tYDKuMjDnXqHsRrGDw9FzmaXcotT97mEqrpfZks6YbQHDavYN0y2P4vJ5a1lRdkYbSZPyZQId
4EGj3a2Hbx21r7yMijoOY3uuVVrx2a1IfNFu3P604Q6u1pgiAxU+p1yOiOV1B+T91z1IUL/O0oBA
008Zj1yv5wzlElVwTM5QwXwgEzGYBpCKJ/TPxNsTVpc4Wjh46RVyDEsy27oMlRsSWeHt+5YVn3rU
vgWTTSFEZdz47f/QW/XdP1FSFQyEmrO3UHubYX058mqrz5rskkKxRADuWGiLrgUMv7qK3FX7LgQX
sWpbR3tkifIj/y8A36e5Djau9oKL4fIuExUgmf0aba+ZljPuDNpxY4vj6OD3Xy9sNQdTqDIbj6lt
qUHJvEFhnPZ6t74i7KrifoRwYVLn7Lz1rl9dFOJK+AmF4EXWm1wJN8Eh86SURq80AVs5nziNXWcG
Ol/UmLrKJFTiZITOQqyH6/oziXeRASk1glfUSFmeHe8jII1z64zN8Y9MEN7E7xlcKfL8oqDVfs1M
gyhP/mDsrFnxc1Ne3Ue3v8gRbrP/Duvdk8fZ8XFD59w4IYMhlkxhgeN227roa2V8Ii5pXDTXTfmU
C1qXeDSOL9UGr/BRFaq6unf33/qS9gdFhOimcQSCVsCfovNp6o8ylwRrzZl+StbLaNfURyJt1aFV
6RLamQ/sYikzYhbWK03woglQWWBRYXv5z/j67/f0l3ps8baKfk4lmqU51aC4cyReXXO8lNu9/NJI
DC7xhTtmnNreSC0HwjLgyaf91QFse8mU3Heq00CZl6lJ6fm0X1t5MSgY08TK0hS4f3tWDA694DOd
CSfv5SR8NLXTFEczvCEAkKNyNsnjY+dVyugGM1h+ljEBs3lq/FT6C8TMtcWiazfmIxwCS1gyIXZn
xyM1Ewqe9zGFRex6zG9JvP4zJla/G4E2MwGYPn0M+DrmawCKeADyTRwEVkdPDcQg4eXCkqRn0vru
3sfnXT+psCW3nfqqNG9+7tq7K/U3ubGx4UcLoSUeUJQhIGNxN2DP+jYgYixCSN4Gmesk8zHpYf5m
iGmtmSK1zB/o2G+vwL2y9R7O6l/Fx3qxgXqnqcKudopJ8+VDN4w/uaWW7sHTxBsCRQRzbxAtqR/V
Sf2uqBvmnVJDy70k57KnG/tkWPyqlYlBwmewtAuP/veB/dMTZBLzjKXVle5KClFqmd5U0HgYzEQ1
8WPT6B0q0kQZZi7VfC70uKFN9sV2NuyfT1nBfD2LqiRAf2LuWiJ/hF97JrKt5QCwvHenEQSaiUU0
boCQcJJBx3Ga1yQOaMFUtHBmbD/XxeqA6n0EsQc6wBaXvOs20fDjXU0t0wzB9plTv/iE68ddjcZo
J5GprdBYH3CReWWk6OKxZvCTcsy2O9lj85tfTLoFVfPr8S6mfqW+49k2OG5ej5l7YC9+gXzSvpeU
aMmOZFNSJpVhW1jwbgTGPh1Q+9wZpryv6T7lQeZEaUigeL2zyV5qBJ1SVHYtGtw4RNVvMXe0ybt9
E6SisIjO19nLEPL9jgMpeQZD1jNDa/prhBCPJOt0worhflqPYwbY4Gs6FFYVmZHN7K4cEBX69sjg
BOwfuH/FAwocrHRrOspEUoz5F8+CUT3HPZZtC/Nv7hXrJxnXTk1O5UTMOQDLaLD5kkVLbCbUimWX
Pj76TcHEQ1UeCw/KGvpEL0TCrnNCaDvSOkG1S4Cz1xzph95jvlLRlGvCcK8f+BNmjWDUM8pbJEK5
HrlZvnB2Fu+3kgNDB2bFIOT0KfUvJDR9thB4PLOLpq+yaS7732Pn9DrC2Dpk8Hmp5pm9M2U/MfOb
Jy0tuUEZFmCK6AxpNlNhuJFyuSuvyr7Zi2bgTwr/b0KPEzAFGGEinBR1MVYAWMWp2Fsw0+g1Dyyk
WMZn+Muu4iGSP3nQjcRjeDmmu8Fzl5CjFdgRYOxIN5zXZWrMEmo3e+QyvtbXmwTZv2d2oCOOINrc
6NhvKdvdQ4lDXWD+6/n1EQ9q/VB5avqCtDTIMTZljhfIfuA/Ku1jZuZ2tHxvXPmsernxCwSUWJq4
x8jgoQYOL0enCAERnR/YM4sfo/Uen9Z7Fw6BdcelrK3pTTHbpLaIZ+aoAiCepOrVNpcUgvzxLklI
sr3MHdkWXhSON+5TnyI6eP129jBUKK8w+Wrl+zgekZrrBGugqZUbIkZwR1RGfEfv/iyTlfcv187N
JRPfaUqZmEgzNZs6Ss092h4e9cuPxwjLkIePkqp/8fQy3dUdIb2pW2VMKMHyKo1hCQ8nYMs0kJOQ
3eEPp5+BI8Oq/2XQUKnMOdghgPRSOXfbxQbhw+7+yeqx7iX+/fP/05VHMsBplvAMsIfTEJsZLRJw
gloIQJLmbtpW+MfArmgLMRWaeJgyH9UK6xsqFCRkjJ///esEhhpKSXtNGCtG8GSupJ5tgIXRk8y3
uPkXMgGUTP6nQK0Wp7JQJ234XHv5Qr2iPgdYCBTmY+ZdI0Kl53gJTIYW5QgdV3jJ7/aW9gebNgBb
LTumCoVC8bLkzaU3L8Azt+VMYevcjMMC5B7Zdn2n/73gqYQNPxxDaaoSjz4FbJLYHp9U3faKw48S
aqOvBMaoPMgNGgTSK1VzukjQvZMR0cIJxhowvPJbpKH2hBAw64k36R5GLtd8plEeUkmWf/m9z3pb
vw0UiVUNt2elrG4ddBwXqvjUcP3A6Z89+YvlNZ8Abax2yc6hf9UtdeuwSmlNsUiiZEuJiumBVvGA
aT+zHMcMFDdrJ/KpGk8TtmW2gyyGY/aa1DpghoFMcryIKBX2/jGpx6XPHy72f4uojRLbrEmOYabF
GxGipvV1tnthbWdRU+B3i6JlXWNO7HEhwraN1stZEYO2H5/RsWNuoYq8arGegKJXCWmq+u0lebLA
DJpKHTRL4S4TazvEsubH8UUyJn67U1fIadk+3wy3pDfOJzLhSApRhmM/id0WmHjq4HpltyY7iomU
9imch6Kegk4xuDh8RF4rsY8JubjbqBEroxXsI4W8802vgqMYAEn8JzI/NF4KeVoMk3WFvDxeU3u9
Mj8VPuRc4EvGjcwfljDPAhUeQmJ8KZk3tzRtviimlk3q42udNlmJD0QV7hLkHyp2d5EfLsWg1Wbe
dGYSjPx3Qd6JkHOC7JzhvFokLESHGqOdtz97ldn/aRF+MaVcbGjSCmjjbFxBevr5xitrOY6rBm/D
Uq+J3OGdxeFBWlWT5fZslt6aqY8p4hQwmGeLTS/MyavDnvRc9tgSL7AeYaBNV2yuGJmW61jqDHJS
mqOIFjUoOrLWROLJ+oTgeg6oWxct0JGaVq+UaUSZNLJO2c6MM4Sgjy/6bEqQzd/aekHklv1DVVOx
0OmskRToyacopk/KRZcovJesWHgK1aPnIF7lBRUB701WD7DhwcCDwqVFWoNCN2DiWrAp9Jy6jwHy
nvtUs6O8/JDsso/dFvAQ6++wBi6SSwKwmu9HpRXltO7g0kGzDHczAnzCcZuSnGqnfGtQMoQrKbFL
/c9tqLzi+rsimmjeKMXUvWjNWqFyqcJjM8lZhC48ml78HwLXuULpSenc9AggZa42JH2iOjVRxovj
DIfYETzLlJI5V3ZiSZJWmBpIKyWEkWlO2hcEZjjh6xZWkk8VN1+xD1kLFYv0pB+EKFj8EMEpjNBE
jx98+txDQQkwSO+ZzHd0upPKgIGM/ipJmuMItNsww0vGvjcwhVqDSuuOHSW7IpjS1D3voHWWc0dN
im48jL8X9u9NO5smEip6g7eZ54wqfHsANN9Bpbop5mnbAltUE24vnvpp+xMKcGG3aPmyFIsZH1b1
8VUSIcqw3z+iXT1T8FUKbZ+KLt6mmz2W4NnthfWOh07PxritBKebcbwJeetE+9+9rWahxTtHxglc
2aO0880Zx/MzcjGMOW35j8TDwoLmbGl1kZJoBV5wWLFuWKQfDFJnY7v65Cmpq0CNy5uVF8nCDsro
xoBPR1lCKEZr72ydhPoyBJ+lMKovNCOjCYJ8/RYmxzpSTUvAXuWn6t9cF4++pseAtjvkcRJMwEOc
NKyz6s80OnK6TWBQzQ+YqoYIoIttb4mGHBaYMKq3ewZBqQ==
`protect end_protected

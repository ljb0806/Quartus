��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��I9*�33�%B�t�A���n�ݐ,�9��ѬNR4L)"<��-��ZW#N�{
y�v �i��l�KG.o���?GD���:��v�
��)O��?}����v�J�$��X��2 uc�Y5�,��3azT��ݏ��G�J�7�Y����F0DOu��"m�H�����AHm�m9a��^˽����F���lǯ�o��'�
 �5�d�s�}�F�ɏc4%�!J�*�y���n�܌��p���<{ך�,�~\��e|��X�^�[��g&�?�@�p�:�`����߇ԣI�5N������e7��L���)R�͏4�_�.���/��vk��0ʺ�-6�H��=M�,h&yud�FVМ�E��	�����j�c\� �Du�"���܄j�[��4�#���(�W�ToQj�ݐ���T�`MF�n�vÃ���<�VB�������s��k�ɘ����z�GM$��#7��z��L��7 ��m�n��)�����8Tj`�Q?P�[zq��I���!5�ñ�`�?��{�8��u���Wb
e��"�y'�R���t����핑i�t�c��P�l�%��J�Bδ`�Q��U�@HR�AD-��u��萍�׈v�+;B�	o6�x��m?�.X���,a� <�AM��򳣾Wk*�p��O�;�>K���Mx=R����. �D����՛ʬS� ������������\� �g�=A�'���?O�(ڞL{/�:��/| /j�ug������M��Ӌ��v�&fS����\�HoE1x�>r�ʑI��#G��#�r.I�^�/@]�{��Qc�h�Sk�wC�ǝ}�	Q�F��l�W/�k�n���0�D��	4�ثv�hk���z��l�]��sGϟ�ʿ#i�|�7f+�_qE�?%�ܡ��Gq�vz���`.-�o@��<��q�#�F�Y�d<��PԔkX�l$\�p%:.m,��F�{ޜ�;�)��H�S}�`}�0�<��C��zw���J@��2�Y�M�;&�D�@��1��zw�WQ�z8l>V럌���m*Z����~��;��9�s>�w����G�q���Ii"�5eV�e���86�Θo��P\�y����n����v�i
v�(�9�Y�I�ǵ�O��V?�F����	���C��|;ͤ���DXM��n��P��Fk|C�i��K=�t��g@�~���N�`���G�]���)"�e�N�A���e���\�Wi���\��C��U�����]�|S�.9���:�&iJ�C =#��%mvv<�ӑ�U��K�wE��(�zH���ap���-�FW�F�m[ql����x��ߛ�\�������J�a��n�..�c]2�Y�>cV�Q��p�A����G�&:��q� �?����K9+��J+Z��fz�}�Ŭ���US顅���|�+���O`�3�o$(��,�Ac@��![NZl0_+��E�Oc`Is�.ē�3��t@(�������/D���oC�����]ތO�mƝA�E��3�]���($g(z���k�v]-<PJ�V�J��ү�!��;K��e�Z�4�$�k������`?=�p6��T�,���4"�Xy�_��5U'���k�Q�m�8-giH֩ y��.����͝�5��o�����m�Xw�pU�6����-����x�G� \����gY��&�)S}��U누�C�ٍ|�
z�^�1r��*B�"l�?^��߬��T3�z!���N@h$S����z݌hU_�G��Υ��^I	rzkډj���V�>�D�#�V?�x�u��ϰ���I���u��ƺk���B�&~���d�L�Ds���3?�8�����Y�$h��-�=S�6��[~3
7bH��j*4g��!�$�h�S[V�a���CKW���{׾1`��,�)c��{��+g֕�4�ֈ}�v���`�^uY����k�	p�+nH)�1v���6E�8���k��#���g\�+~�(4(6��k�z����t��?��kP/����ݸk����-�k�}>��L���Lkm����#V4�dm�idq�t�A�Er�*�k����ip���-Z7{���FH��J��g/�bC�w*�Y$_�/�4��p4!��Μ�D�d��?�f�3x^��4��w��t�w��"A�kh�sE�ҡ�8�!wjMc�_��+Ї��/�⿡K�"\�~�Sۄ��Z����U������ņ��`�ݦ��ڋWlf�*"fIۏ�`�hB-�r�	Tү	������ԑ}bRե��Pr��՜�!�ۢ=�,���̂��\A�9h5W��I��7���2yWY�4��O��(�s�����
=ny;ʶ��l�c���.K4�s��bAj�L�\Ai����!<�+<s|�
��Y5�`�Up��N����,���n	
ʜ�9e���*�1�S)��#��%22LV���wN= <;��ݟ�ci�8W�9�Q3��q�=�PY���y�~�1��X�=4)��a;'��-� @?K��c��͈�|�;���� �u}O��?��q�?ࡿp�XLU.�fu_�sN2�Ga�!���^��|32�h�*Qn
Hk~>i~hWY���<������4��T�o�!v4�\,�id�n>n/E�*p���\����&����c��^;�s=xъ�h,�W�X��-z9�&��w�s#�x)O���닩�1[H �'��O��F�"x����>�y�A�}kh3�
=#efm����$����� ?�IA�?[��X^�E��>���q,�ln7��C|��ܕ$.j5>�M����0�s-��Ί�!K��7U��b0B�J���C�.?�dz�+��3	\�(�yQ��L�#�hwy�8'�~Uȿj�Ѡ+��N�Yd��/��k��t�9���r�iUu/��)Kd���h��ލ���a�14���r�s��k��b���C��uа���"�����zD$f�"��"�P l�*c�J�1@��뾡�3�hD�4&}��k�ο��3b ��`� ������#�(�	�����MQG������3@6\M	��mŞRd��M��WUQ
T(6�9G3��\��g�`uN���*�V?|>�פz�����J�}�9�礎T3�o�_�2s��������w:c��*Z��e	�ő�z'	E$���I8��ѩ�<67*u��z��WL+��r<�
�]]W0��:��3�x�c�P��Y4�~����C�޼,�E�欰�?�q#dO<��;//�"�,@�ԋ���	����.7z��<}	N1n�:�0�u�H?PT�΃�x_8:.%�B�ERH �D.cQ�ض����LQ�;�5�H���¹Xˣ�?���~SpE5�I},��tַKN|�c�!�R�� WD�����Of:RbG�ˆ%18�R�ϗ�/��޷#Kض�me=#�v��8X~�\�) �rAOGo[Zx��D��:J���L�U��Ш����)eָQ���v��jh%�Y�]��M��Dd>nE�ؠ!�W����DCK��fpN��
ş�������B���`���Z���h�|4Y䬹�����3Xc�"Wj��gj7ˇ��Z���#��.��pǆ�S%MM���a9M�`��a�~�Od�k?�S���iI�����=7-p�p�6˯L�h�5i�����jJ:.����m�w>,�7���N��6ӵo��a������25�U��$�%H�k�a�}�J�%B�x�"�4�����e��dB�<Q, �T]��мXq����m��W���T�*�i����}�{�UK�ݚqSк��Z��|j� �����n\���L��sr�_ 㓤�j�����7���N^��W��E��WY�a��k�҈Yjh���zt4C�;�4lL�a�k�#3���q\���� B��Υ0 XB�gZ��}�
%/Nt�כ�r�Ԙy��B5��g)bo������o��\�wY<�k�e+;ϋ��b��&�WW�.XQ��Rl��w�̔�M��_=!��toGJ�pMɀ�z#��)�3�
���0)�Ī���_ �A~8�~ ]A�Mo}�Zq`Id���`'�"�ϳ�x6Q:<��7�-¯�·%"�w�8�F��+!��V �����Û�1E�O��br�\k�)AM�:�	��g,���<��+a\�@K�-g��1x�6 �x�d`�F<<.;�+��^��PB�x���{�Q��A��ɱ����oeT�tz�-]���Bb�Ʀs�'/�A��)k(?�>�6lc[�J��y�i
w��g��޼�Al��/L�
���II��O�j�A���1-�/6꧐��ޤ-���ӂ�?%в�Đ`F85n^�v�1[%�oY���Zߘ�1�m=�\�Ny!u��B�0�������k��WZD��}D���v�9����M���ôQzF��=;B�T-�L�QoY቟~�>�9��;�ix�-w_2;-~�ٕ����Z�5o�����fA���x�scN�$wK���[_9T,�l_)7�wm�#��K����RT�70����}gY:�Z�Y�!�)4CR��'0�.���r1C�(-N	��J��:���v剿��ˇ���n���xW�AJJ��gXUTy⃸!���r�m-��*�����t����w�9M�ʋ�@�k�=����Y{�:T]e��hz�c��&2۞�mԢ�l-[kw�:'~��i��O�"�������$��?;�lA�)�u��8!8X|\>W�쁍(�x����cP�*�fʶnq܂m ��!d�b������rr1��3Μp�}?G�OR��ߤ�bT;A�g/���WB��8�0�f� |��賵Um�3?JK�M���]bBv�SQS��9n3��z �����f�I�X��Y�_�l	HRQ[ޜ�3���P����F��$�2�C"����NV�IMGX�u;��7wn�(dV��*�V��%�$7o3@��h��B�k�$�-��P��T�>�����?I����hH�4y�JMz�8}�oؒ������ܼ�ņt�ެ�81��~Uj$ ��-�`��c��~���Ԫ�a��[����)¡R/����V5���Y9�	y{|2������P�:{���qݗ�������j�TzD:k�BKd^3���̚���A�|袞W�\18�ʙ�T尼)B��m}ю}Rm�.�*ʭ��k7_�)�m�mZ���6��{Q��CSq�6�����v�b���<�{	��2�UZ�U�F+X�ׇ��c�Z��s魬h!v$Kx �'���ԲƟ�͏~!�@Q6��`��աCo�ʜ�y�a�
Y�=e<�����c,��U-C�o���\���{Kc�s��G^��{u�p�O�T��F�ǃz��Qa��7��������B�'u��j���F���D��[R��D(��w���8�#d�4��"��D�CxtV3*� S[��$�A[�C�՞�Ǌ��C��a�����k�I��'� �-~ѧK�C��E��w�ձ'�/����0^����2���
D�syN�@�B�%��$�(Ӯ�sY*y���=�|p��e��a�*�kD��Q�mAl$�D�,��6�?���e4@��Tf��O^�ְ�g��7��<Ѭ�JOa�����n
(��8
��Y���j�'�6t+$�g�Q�T�F�4���QN�̾`���;�j:�ϔ��ֿ"��t���g����z�H����fG�1~�f�
�+�0.;��e:r��R�v�ҳH�凗��ڴL��RX����}!f�;����E��εn��.�����΄�|Bb��NƄ����z&��.���|b%��'�F��Y�B�� ,%���;�mV�����|�s�޸"`�!z��݇�ղ�]����(�>���bw��e_��f]~ϥ�,$K���і�kC�C{eY<=����X�"�~qfr7%�SE���>��S~$�ʊG�[�E$�9T�g.~B�g��$q�/����F?%CW���b��5�8~�e����"+���A�#v�)�c�.LP�[�f]�q^�T�GP��:-T�	!]�z>�_�;�*~��f��i��G/�(�0B~$��⺲�pvvP����ڥ������
���E�K���P�_�B�A��g�KW�Z9Q�;�3��}�W�.ad�"�@f�����j�䣫�6�qU�5G Ws"X�S�3E�?5K��!�$l����7�k0+l~�*p�ԟ�h�~����/�����נ�5�8TK��Zp�v��\�b��0GCg�������}&�z���X�rCnI.t�����(�K%���wd�E�V�	)>
z!S��q�szT�>�e{�w�{�����At���Y4�\��6�Xc��-'r+��A�
����;�i�;�_�{oj���}��T�u_��	�T	�,����%�q� ��%�ͷ���G��t�t��q�o�� �Yz%��H�ŕ�T�S��|7�<AV ��nqX��g�����,�m=��J+��Ӛ�e������P�,�]6�5j�c��[�H�t�0Rs3���p�2��H�v��c[�/T >c�[Me�;�C�?D8[�S+�����g���h��������,V���o�N3�5�n�TS[&P��۬�"7܆�ݘ����/%E��hW�$ް�Ol�:Z�Bn�q|���E�*'˷)L_�氳F���^̥bb�q�J�w�5��~w�#��`;DK��'ki�!M�?��s��Ò�p*�imD�.e?v�'I���!���b˓����H�C�d��ʃ.i5�X���'��v�s���7���׼���l/ѻ�,TGaJ�Q�:�͗����$�lb�f+��B���$UT�yS��d1��@_]X�m��
�HT���ǻ�!�4d�+jx�煖M)�i�WF������Vm��o>!ط�l|@�
a[���Q���U�f3��L��2I�@�c���� Z�O�Fc��n�B�[�1���L���4�*2K<hE�_����;A�3��4��-�]��>�C�:���5h������A+aQ��Q<f�lT�!du��q��_R������]�4�Qw.�����d(��}c���Q���^�S�u�X�i*��i�mJ� �ش�=s�}&��L���b��� �o�XF	}�u�X��du<Y.:2�@��ټ q�R ;�����\+)�=��R��ȧƞ�4�TKJ�C�D��M~
�{���O ��?5�f���`ҭ�L���Km��s�Y�cI��4��{L�,�6�#z�����l��,��O٘C��lɋK��u5�Ѯ[���CG��$��?��pc��3K�M���ty���w|S�����[7�G�R9�������5>�J.�`Tϐ���_P���4l��YK	\,h��z�lw�w�K���%���ް�{�(����y���&@h��H��X,H.5�?9���=��\�b�W\�q���\ �$�_c�.y���8	�)�5����������%m�1��G�����'e����>�l��)�$vS5�/lme wMu^F��-�:��.�\D{kz&�N�8<�>Xr�o�q�ua(�$@0��\�ҏ�A87X%������a�zy!�z�s��CY�\��Lk_P,r^�9's��I�]3�<�����M�+)?��M��|�"l$���|��Tnɱ������Y�o�H��g[
�����;�#���(�n)�C>ZL|�$���ts,� ���m4�W��/����ǟK׮���\e�����2.�~��ۙd�w�-�\���5��C,�a�As�¡SWm������l5�!.�q��ʙ1��Jݰ!�,��=����%
�=��c����@D��M.-s�����W�Ò^Wأ�}g�46�M�2���~ޠ�m��tz0j��B�m�vS�cO�p�Zn,&ɲa�Wv�W+g�S�!��w�O�5P�x���`��%�L0�.����9r��Kc�%�=����Ѷ_������KL�������FeK�#V�H�q�C�@���g.���W�I] cj���������F`t��p`SKS5nϘ}�u�
��8!���4�ހ�����ַС0$���f����V�U�r����ĩ"��'7��� xP��U� ��,�X�/.����]�x໲
56D���9����ȶ<��.�>�ȣz��Dӗj �z�N���4ؼ���c7ʕ���+#�ͩ���އ��ʛJ�Ӎ�?�:���-U����@]�o�qd��ǳi����e{kdF�>�&��qg;-8�yԄ��S]g1�x�ٸ.i��64�t�9iBg� ����}�ck\Fˢ�`A�r�w��	)�6=B���y�ss�g&c~�~�+�s�"�5|֢�K���|ɵ����#z�.���m��|Y�Tud��0뫐�XI~-5�$O��Myv�#��ҤsR�"�qnt^��X����p?ZAGբBkU��_�(	��V� ��q���qX���d��
�?,��=����b�*�q���r�q�>>�><9���������b8`�g��e�!��Hry<*�׌�B�S5Y�+�8���-�Ʀ-l}U�<2�E�B�M�sw\+/� � �� ��0H��z�)����g�WK���%��~��l��+�Y���XEn�e��f��<�XR������g�p�7`N8�֠�e���WF�n��T�y��/I�Y�ɲ%5[2?p�"�лERV�]0�+�eD��S?I���$U�wT�״k-��`�[�,������C��2t�C����{�|�1ě�~�\%�* �����Œ�ɿ�����"��;6̆��2�l�j�#U��E�SRZӑ�Nlu�k���YÄ|Sw\'�F`�
�o�F�`!��lY�eV����y�ʂB��gׁb�9_��S(�,[�� ���\��c��L�I1cl�rW[~�=d������|c��VvBu���*�l�$�&֭�&,��/>/�Կ�\Ď[_�sb��R�L��d��jF~��#�֧A#1���dv��	��/��rV��*�(A�]i<�
V���>]\�Fj�k.����T;���
���},�����zv/N���3[�A3B�is�-��>[��a�Ʉ��腖<u7���8��Q��w�fo�T�l\���Q~� �E�12Iw=?I#��؛l\����@�'$��{����J3���O�������u���k�$VL�Q����WQ�b=��B�t=��I���o��!���xI�~����������<?葰�$�����Σ�CE���+�ϣ������c��DA�A=���L�������r���H�^��n~ac� ���0+v!B�o�;�.=a��>�\tͤ�k�,���ZpN�����~���%��m�c��z(Ѐ0W]�1�wӨ�2�d�%�e�w7c��W�Ň�=^�X����#����,��v�Vx;�!�vd��߈�N0��h	ȏ'��6ZY���-<u��b�SQ2|&Y4H�M35�BŒ�����+�G'��U4�I<�! �)�ۗ�&(��E���t��H~�c�H{��;�cI��%�M �;�4�B��t�C{��.�Ռ-p�\�)6>�o��SU�m�������j� �c1�u7�AM@�φ��o�?:E��ɧ�Y��y����3I�U�c]i�(d93�!I]���8�G^���1,�X�����(�,h�gE�ͮ��ΎMD�f�����n�Z5}{/n��۲#?(F&4h�?k�y�XC��?Z�lX�q�TW�7�j��G,��_�p��A��!:�!��%S����ukD�5n����{����A�8����~�<�RL����M�ў#��L�δ*�)g��:����T=Ƿ�CWh� qPϏb�S#�ڢ�� ��3�IE>i;qs�$�S��̥�pVX�@QK��<Bz[�2v��6�L>��U}��m�����a�C'��L��\72	��<��Zd�N�q�����K��uL[p��Ȇ���!ew��a�l�^��Gj��vu�ڱa(]���$���t
��S9G���|U�G��>p���1��D#�ҝ�n��u<oނ��8�T}�1��R�Rߓx���� ��'|��6��j��T�,J�$���\�x�p[��y�A+����)�YܭY��8��;�-M� k�����;����J�z�~��d7��CB�p�(L�h�B��ُ�q��\�����`a6,EK@�j	�-��$VyZd�a�eny
u&��a��.���k�!�4��<��+��߫etᘯ˗��|}�ѵ�o��BѮ�޾[x��Kr�ܤ��ftP]*���� �5���f�zQ��̯�5����v�]�tyA�6U��h^��w�Xb���%F-i��m�K<mlZ���|z]?n�	�0�cS��{�舵U��U��0��r������<��o3&��e���	wnس/��te�:�tR��aUJ�ݘ�V��:�Ġ�ml}��f������Q���7T9w�^|�K����P)��G��DRQ����<�3��6:�ʹrhV�ԗ���	���p�[�nÂ�i��.�T�:W�'Z	����U��,�v��9������e��0���?1���;l5�5N�Ҩ��\��P�2`��doS8Ʒ�ε��imo3��V�9�#�qdi吺����M�aP���h:B��撽0dU�*��'� _���~nLVx��+k��� �ۑ���T�LX�\0�� �*������!������'wKX}�����v��64���<����f����Ÿ�Fk�]�����8ʞvi��v-_�"h�@ξ���s��^w�Qxo��J;{W�%QBh��.k��8��}�q�(��%��\ 2B;?�c`���}k�7vV�,�0�����`1nܭX� ��I@���[�{eO�h#q�/�Ȍ扖>^K��a� �BX�����ɰI��{�`P�)�L�Ʊ�)�&v�l��aQb���ԉ�{��27'��u�pS����z>drƜ�_	����+��Bd�W���\�L<�ENô'l���f�l����T�TY9jӿ���.��,�9%8��(��c�?9�yB&z;w�Y�ÿs_!�1dLK4l?�v!�w����.���5��j5�~�Q�oD��/�E�:�+��;$V�gO�9�i����&��;��s%��� �tg0�m�.%efB�*��уwk]��Wk��[��4��U�D$�����%�Y���ǒ��Q���Fq�W~�f�D�b���R��]�_�*�
��DThzŠвfUz�"�ofm쩺�)E��`g5��)����G�Ty�]b��$�1엻��7���Ә�/!��c��?�ӑ�� \	�/����3\)
#�eK`1�ٿ`�\rπ�&�Ш,ι�cV�'t����l&F���P"(3:��'2���O,����B��e��[���?�O�n.��!�l# ÐʠI��_�^���YŮ�b:��g�{�
M���j�8�r��{���t�|,D���	�z��%̦9����sa��p�YŰ��f�牖���[�e�fcdZe����ҡ�6
F��؝/�Vi��,�'��%+b�Ԥ\�At�1�R�\��(YsH,�yx�2AQטy��3������VSr����奤;�=����D@0��c�d�۟O����|����;5�O~��r��2�C�����0/P���	�ZH��}J=����q"-�P�0a�\��ў3Q���%��;�X+�ة�XOa�@yl�ҺG�'l��Zuh�~O���{�sN~/kqac��wڰTӌ}���s��>�Wq�H�#��<aaը�kN�c�HH��Qs@��*� ��<�;�.,C�2I]��D�J�T�H���Ќ�礙��kbU�:�8�ȑ0?�:y���r���Ff���4K����P;���0�R���)���)�%O�rz�.���z|��=OJTw1�r�p��2�"ia�Z��N}V�t��5�B��*����u�/^�.`��Q�ߞ�5�1�ڷlB�<�n�N^&�JH��ut�}о�v&*+?��?"`>��:	�4<��~�C�O��Rk�/~���a�jx��UF쳃Ǘ�yk���ϐ�A�Kb���(h�gw��6y�\�2,^Z	�0`8yGwp)�C�b����ĵ�����ůF�m��l��p!"��d^�Q.)Yc����N���AG�B0C�}��X>��94c�l�����I�#�K'�Lݦ�t�s� �O��u��,�qM4��H���`;[��H�3b���\<WYgI�������"v�Y@p)y��ت�V�e�&��i�j{�,�3���q�Gb�Ia��iA2Qoȶ㤌�cצ�x;giϚN����]��0{��Z�2đ7��3��N��s0v>�Ԉ��&L�2y��tu�9���I�k�Llն���D�\�C�5�G��þ��](O����>
{P%�uzb2VD������q��h�|�=j�eV��Vs�ƨ�����
#.�&�Sҙx��7m�O�_X���n*8�xġ%4��%زW����C����"F��>$�1#���1�1=�8� �����<V��C��J� ���))$eS�1���PJ�˧a����d<���3t�1��[iY����fT<�I��:����z�Bg�܇����uf����lg�o���?��
(�$��$;9rm���d�r�\ύѹ_\�䏅)s�)���{�$��s�������a.:lD�-�윅cr*?��ٖ��J�(���L��%�}H@I;b�xB:�ɰ�|P�Q/u?Z��=����~����dK��D�P���S�ީ�j,�ݯ�d�R�*����dG�o7���k^"��29[�k�)L��G6cR�l��7��\F Ѝ�L�)dZO�E�[�����K�މ)am֛�ß��м�m�5�:����׹�����J�r~��[dEvs[���N�
x^EШ����_������Y�H��QS	ڳ�ׁ푊�H2�Y15��q��۩�s�������	.ԭC������3��V���y�|�^[U�j�%��C$�: ~#�����S�X�X��Vz�Fp�;&�w{N�hr�z�3�W�<�)�*B}�$i��A(D{+��)ߖ����pu<-��~���"�Y�������kn�*H����w*k\����0�G���kW��d�f��4�OL5��_u?���s�w:�#SN��S^]1��qU�pb�g�P4��M15p�����DlU�{���۵�EZ/��Qx!EGگ���0'�1�/�*L�Z6�f2̴V�}�{o�f�� r��nZEkF��������![��%�q�t:�4��K/��I/�^b�nߧf�o33���V������[Xhc�c���Z?�b��̷$cD�r�	��0�+��(Bޕ&��5�JՇ��t
7#�rPP��D!�6i�sU���+�z�����;�0����6�Cx��Y�J���֣��e���r�+`;|�u�Y���>��/A k�`�#��*�07[ݳ�N9�7^n�Gm�
�R'��^H��Z����*٪�,��bu�Y�ʦ�z@{)H"�S+D�h�4l�5<��Ӟ"k�^RUA]���n�^Gnc�|2+OI������r �� vtK��в�ƶf�~e��?Z���դ��%[9�X�Ꜽ��'4���g�H�6J4/-�;I�˂�OQ�W��3�&�"���H���+���
�>�p	di�����hэ�f�Qy�Rl��i��E;e�j�?�����rϯ��� |p~ƚ���1�թ`�0{����.�R�8odⅾ����a�t��ߝr�)Y��9{���z��T������]�EG+M;H����[�jvu�⿀�ax�^y���[���~L���Nh�$N��c�R��T`�<su�0�B0R�nͲ],GO��O�b�i�W���T,"�<��j����
�铉��#���I�����#o�2zI6���L%�f��2fW��n�/43�1Q�N3��nV���*�
�����`�O ����Km
�^[���w&��ZΦ�q0M/����K�\>��~�)T4-�zxv��6JI�aM�1��}"'��7Z��R�M�CD0uu�F�(;e����B˾�[�\�m�5=u6 E��Oo��%�#�{Dh�mV�^�=�o�2�p�'*xX���r�~L=cP2Lѷ��ʤ\)"��q�}���J�ӗ�$¢�c�#��3�� ������}A*f�2���k�\��-ٷbm'qRt�������ϜM\�Y�5�β�,�0�g*���FU���[�ϐ�)/:�ܑs��c�����	�i�&ֹr x3h�"�m_wAh&B���,AA+�����,L���,�Y5��Z���bde=��)V�wU{*Mh7nZ&�t0��N-��0���b����B�D��[�$OĂ4,w,K��>�����j���;����<ug����2 #�~�>����n����d�^�CЁ���什3�b�=�=czX���RCLV�Ͳ9N[�[J��}�(>-�L���v ��=���*�E�F0B��0I,�#�#z��F�
A��[K��͔P�s�țc�5+�0�3���I�U6ش=�¨��/�\K�?��~ �J�����|��y=�Ҭ�R ���Ya�)GY{��F�:&�S���j弩e�Ș
���eY���߯�&������Y�E�93��inLa�E�$�E�f=����t��Z��q~cv���Y�����n�8�ڌ�a�Ez�	�8+ I3p�q�����gp�����a^e��q�dsW51�QոQNߞ Yr��4�r�-G�2{(İQ�ڣ�A�֢�Q�¯])vz���6��jH<J?1s�8n`j#�h/"g�$�� B|Ӽ�2����%����ت�N��ʂ#�i�
�w�	c]��v�� $t��eP!ʤ��5,#�-#؉R��ۤ9��V����	��%#�F�"(�����a���IX,f�����n>�����H�r�+k	���%���_�������I�`g�2�#!�t���9e~z#��.䁟��)FA��"�<�H*���'��w�ը��Y�CΌ/:�&:�~J����2�-�Z�F�<ȅt&��0+���A�ֆ\�,r���Z�ʐf����v1�9@�y����y�~�`NÒ�p��͖��[� �m�ƻKWѳ;P/���7�:IS��Q��6�p+����l����G�`�k�PJ� ���
暸�C�­]?k��9{�y	�Q���z�)��l��j�dl�����ۭ_z^���s3!-���t����n$4�+3G0��C�u*��$E�����$M�~V���`�4�&n��i�����㩐�l. �QԎ�NtG����{$ݏ�#[��p���S�ӕ�T��%|O��P�rFh����+ĩ�R��랿9$�7�ܷ�.��r����3��@)T���K2v�Ϭ�5����:Ov�͝:#nP]�U��@�'�(Ҳa�g��.~������e�'�8Џ�vi�wvx��~��U��{��������qa�A�q����0�� ��o�
d(Y�KbgY�bJ�~�v�l-ܮ1����&����t�z�!E@C�ah��\Hl����=��!��U��.�R�\{���Z�KdլL+T]c�>�I������緃ҋ�u����.�b�T�<oZ�
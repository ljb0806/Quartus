��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��$��~n��4��P�뛥J���h�c������j��-	3ǭ=����0��YF�4����1���� ژ��8�*棹�N>�,X�O�!-���iH��e�	2�7й�^�/����1*���}�|D�ʼ�&$��ѿ�DӒ,���Xҡ<���kr71 >5@���,�p����ˀr
е�����|B�[F�(b>�ęHuO����a�`�y:1��}|�9��I���p��*��)�;��T�j�D��uv|b��@�}s��_ˋL��e{�)��Nt�:?s�>�-"�Θ���k^ �Mm���~e�t{%y����p/����fIP���M�Z�4��b�%/��v�Ex	b�
��b�����<��V��KdD�'c�3��W��'Ƭ����Aχ���"aA��SO�r�f�D��iH�$��3�N�d�۞ ?N\�%?��b9�UX��Z�3��R4S�2;q��@�ci��x�P��b���~+-(�c�˷��� �8�K&"��G!�fSc���i`�F�f�M��gK��Pxyvҏ��'��2lCy�݌l[)M��#����=K!��"���o��K�[Z����1j[�'�Bt��6��c�,R�Cqj��*�l���F��,��S�=�������N�F��t��sΘ�_�!���4n�&��R:����l�����b�?H�d%�����ض&��\sl�0��"��A���Pp3{�bYD��IoڅM!_�5o�ˋ�`�|.G��hD��j��>\��҆�T���aW�Nyʥ��.at"� ���wՖ�^d�؀ǚ���Oq�Ck��DU�r��=�����N�7q��/z�%��u�Mq'�!��Qu��,�y���:�.Z|��ì�F���_�r����rt�/��Z��)�q1�_#��k(N։����^�̮i�.S?u��B�3]q'����'A�ʛk<��M4�r�ȱ�h�a����8�U�
������nr{ RǐiRV���
�;��"]
�l
�iL� ����&'r�F��W��>^��@{x<U��ada���S���D�*�=;|�f+Z��{)d�u$W<�fRI$*9&�jÔ)��+���6�rC�=ށ���"G�^������%ıd�b��A�Q}C�-��C7����N����U%N?���nQ���'�ܵ��EE�����0���w�t���2��2-Uy���y�+�h��"̩�U�և�<!@^����f�7m�SQ�a",�V��
�D�ҊE΅z�O�1��'�g:!w���#�K&�����?`;�C��='��тOA���H�MD�ts�
�Z��(�0qXyHlШ�x�e��!�XU�Lt/�A�M����� ͟�xg/�O�:�@H4���4�9�?w!x搅�	��;�����p������#oN&H�|�*�?"�d��$�?$(L��)�?�)k�g�?�"���*nV�s?̈���t��R�!�Ԩ7H�t������ɏE���a�����4�!�32i]m1 *��#��~�5@�:��6E��K�El�w<��E|[�`a�ɪlʑ7��/����]���EU\��AN�'���x9�"�(����@_+��4�*����hx���{	N����OW
�����9��A]��M&U�~��QD����C�� �v��u�!��N&Ɋ���ą;�I3��=��£������
�u�By0�?�8��A�Ͷ��ƂG-�ѦgH�a�v�AG���Y���HN��Q#'����v�_�Xu�F�D��,�0^aX�(�W`0���ߊ/U;��a��ܣ]J���e\\�
WP�2ϖHb��FC�?oa���C�'�ha=Ǣ;J��9�5O(�I�W������͝��t6M�(��*&�)�eRIP�;36�?_iLO��:���zٟ�A��V�n�>0���2���v�{�?Aq�
	��pލ+���d2���ʃ�T�_K���>gs�t䞺�`��E�5��cC���t�o Xum�'�?�'�%|� 3�^�l^�g�ˀ��aAf��?�t`��Լ���'�g���0���	y�6���<��?�#��	@v�rT:�էm��A�s���M)$h���1��(��-Ok(��c�
�@�P�)��?���U�۔���PO(��9w�=EH����#A8N,�P�<ei"���\?��$��W��Nc�VD��gT�]���S����Fl�?�m��C�c�7ER�f@�/ �T#>��Z#4����_�&џ���rW��we��R����G�]1o9)ڥ�0��׃&?LM�g="~1�������]�jV�2:�||��c*��o��9}6����oe�2�P1`���A���z�l4)�f�<,���&�'�=Ҟ?,�t��fٜSafH!���	n��%v�b�J �Ϗ(��n�Ŭp��O���+�©ң�����ޖ?���[��`9x����8��o�Ů@��^���>���1e#_�� � "��ڝ�O��i$m���� X47n�'�H��A�w���^^1y:"�"�Ɓ<c>��/���Q\애邱��,C"��U ���̋ߡ�Wsj��y�m	��E���C9�J���U��O�ҏ9/{f��~cHpy����X�baQ�!='��=�NZ��lT0e+��p2�XS3��	v牒��F���>|7-6��p�K��� +x�J��E�?$����4t߃P�oū�5�Vb�n��j��8�qU�8����/`AZ�w�!�����O7�'�?��s�����3�'�ó��Jʃ�3�0��@�k���,�/	�!�� ��Md�j�$|�VU��P~}��]b�fN�K�:϶����@YB�D��Zh����S��Ms��ITL�"bw�^n��]�w��1i��_�!�Ω�*�.D)ʶA`�䝬 �J���@W�@�'��f��$�rz =������ e�n�ڎC� �2F��q/�����f
��ܱ\�]�|.�e�����m�|�@�¾z��Ɖ�En�����n7���M�-(J��CLC$��E�����c-�����=�L�t2-{"#�jKH�qR�2�~݂�xX�$<t(��Y!�f��V:j��ق��B+���� P�LZ6��jq+�={5.������p�I�
̝Æ-��G��I�kPv�T�YX>B����ŗ~{�F>�jw���K����n�o�>�	Qv�]?�D�#;
d������c��	P!
xH;�aL�hb��=A��PĖ&���"r�N5�
�!Q
Ly@șQ�ld��
����5���i��rH�kE@V�L�l�%|=�E�#M�c�s)qm_�� �42�.�Q���)���i���.C�%���~��ܮֿ���?Y�O�x�L��0��ZR�4^�Y��|GÅ�E��	���}�<)s�_=^ګ{q�k�,{���5�з���tMO�)Q@d�jq�SY��Y�-�����1��N*<ngf���rn�(��A��𸘇<9�c�vpO�u��G�駚���|Јw~��M\Ah� �ad�oG3N��Ͼ�4�!���]�s���r����L��%���f��Tju�!�v#�j�؇G�'�IC�H�?���ϯ"����T�"�UYd���o?E�A�j��]����v	���j�R�-�&�z��,�)Ƞ�~27�O����=>�"�so*�'�a>ᥳ#�
=A �߬wv�tQ@#��S�k����?еT~nd%$��O��fT�&*+f&��k&��!�_�a� ��
��y��5S�\zyhALE{��B\�cX�ę���(�W�ʚ�)�[ 8xS]�ٙ��hw���9�f]re����N�wGZ޾C��v�Ks�(�q�捨�a�1k��|�z��bK��q��'�)^���5�O]%D�s#�=��	
0�[O��5	޼��D�z������W?�{�zc5���2�D9�]��LH��R�K�.��	ў��3�o�m���r���3a��F�ۿ__�V�~fBe�yQ�X?g������	�)r�C�j����#"+z6v�8�ͻ�<1Π]Lp�����Z,h���x"l���`V y_V�~1]#�_�Ҫ���.�L�!�w�ի6* z/�~w��[I���\U>F�K�A��h�xI�$�Yr"��\u��U�N5���1C�l�3����6��/2)�d�2��c�?U�u L��#���ȘY0�K��� a���:�qP|��}R����ܭ�Y��A��n�70ʬ�g�鱓ޔ�����{�nQ�����^�^�J�b�ۥ*���;*�cM�C���kˠ~-�����La�*(S�M>^�E�o�+���?���JFRs@�vӎ��gu�N�߫P��k�	��d�{����ᬬXH�|(��.m���n5����ړ�8��SclU�⻳��,�+�]�
%�.YQ������e�[Y�c�i
�@�"2��i�g~�1��z:�3i� B'�LWǔ8����5g��դ��s�l���GR�-�!���v�i��$�:j����?���Q�;��Y�<�ǥH�0�3�H�!|��
Up��`i`HqV��r5z�lp-|��@�4�Z�y���c�[�o(G}K-��W���-uV�+�
/[a���\��-�{�H��ڈ���5��N����m����PqYZ�^q=��:�
�N��wAQ�m�{�GJd�XP�����=�?C����}79!5Fy���@�:�����L�����%;.5@quR����_������F��Mn�����;<�$��㱲/V�C.�h�,4��c�$�x�� �o����D1�ޠ�x�g�W$}i&iBCW>�3�>Ph{7��Z��� :x��u`�ݬ������]���>�t�~�w�sU�h�6������BFȹ�s�Ɠ��V�����f�߆�׻i�c���)0t���XV� 4��靈�`�[,�p���V!f����︜����}Җ\�E�%����w���Y|�
��f���^���X���q˭����
��u5�����fR���$�F#��"�N����	�Vy�J������:U�l���H���Fwe�ǰ2%gVځ��_����Ӌx��('qLt,���P_�"h��ȭ�^�,}����������l*m�K���J�\����I%{f��X;�8u�^���{�ɚ���H� �}��LCz��d��`� su��mvC_T&�p/�pvL�#�G�tǬ g��hI���2:�� r\|�Em���W)3R4��J_�=�������hۍ�Zx��_�C%������	�����18Q]��������a�0��!��t���zO�k����~v&$g�X=��{���b쑵랏�R�����Q (AHX���6k���զ�(����2E`��B���c˒t.�ac@)��rzC,�Q�j��k�]/H��9Z��2���
q{X�iJ�L��]���艶v�#�i�逓l%1j�pyb�9[xR)�������`�Q�ebf
���ڷ������N��S�>~��W�?�[r�(};�lm�0�����W�KVA�m)��ؽ��yR:)�4�0���E�'�&t��2׃2J�P��%CHa��B8-��#d��#��Km�<��o���K���`VsRb�U��)��)-�"Zk�s�j('K�ؕQ���h�P�*�H��x� 8���ae�fv����=�3\�I�5����ħZ$��J	�Fh+�6/������SX�'�˙�J(�U�j��;��Y����ԗ+D껻�l��sj+�Ԗ!]�{P2�J$����w������$T����U�'N�J��e\]�����3#B]��3� ������$)!����`3��yk���[���s�=^Ūꮘ�:�#�dG��ƍ�/0㘠�!��%<���Z�������)�Bd�~���7(���t����L�EW!��|��OBL���J�-]�D;:��o#D���	u�%�y5�K���?{-�>�-m�(��O�F|�	ڴ
�#D^��w��-�Y^C�e�!��� 1Ì�͖�IU6��̘�H��S_,��'�YO���t�m�����c11&&��{�����\�48�\T<ٍ0ǈV�}I봱(��U���A��'/	��
�0���j�W������t���m�X���}�k�o����sN5�3���
�4[�o�W�e^<&�dl���5�3C�XY��}E��b�F����v�=��_��v���u�n���u����iBR���`�EF��%��g�S��לR�\�@oz�%�>R?�"����A`tV��Eo��@���Ge��﵅?2�y�g��i�@_8K�n\�z��TnH"{��@Q��oP<#J��>�����m(�R�4H|�A���N�ܜ�3WY���d��.4>�C���t��>���'�7Fڍ-.��H��"s�j5�� �\}Q�L3�H���!�K��	@1)���H�]��-�9�ه>��s�ox���Y)ˏ�u.����O1��Z�3�?ֵ��r��� ^�/w��S�;@�TL���H�� �D��u�M��g^H"ܥD�<4�B����4����j�=�}�J76��nћ����
M�1xe.K�0����ǲ���;�q#�c��l(;�Uڐ*#N76 i�ժ��_��y<J��= �z��0
T
$�}�*���v�Z���&�O�{1��F�vw��o����������Q��\2Q�F�����z���7��Ɩ�a&�7��^�̐�apfb�FZ������Q��p����Um������Ż.�}5�mj1�/�9E%Y梢����f[�����Ǒ�
�&���bW1�y�C;"���g�A�'��=�:y�V��R��Χ��AW��g|q�c�e�F�K��-*-n���-
}Z���`Yh�P\:�@ҐCH��@~\P���%����M�1�H���vMM����{�,� t��ާ�ɣ�E��M5�<P�������O�l�Z+����*ǐ����� �.����<��C��d>�g	9l�"Ce2��䖁L#yC�!��k<����0%E����+���!'5�߁d���� ���Iǁgp��w˸���}�&�D���,թ���[�L�������������`�b7Ԁ��
�% �V�<�{u�5!z�%p���M�p눆	ۄjH�Q-FO���x��V���},�ͻ�'n��!�
!��q���**;`�b�R.���o�5���.����k_$��+���V�;���La�ڐ�%wԧ�TR�ف���Q�����x����K�:
y^rw*��������Җ�(�}�F}xV�����ĕ�g3�\	dN�|�g9j>��ߗ���.0Ԣs��>��������M�C�%��9/|}&���*�Q�p;ڌ��V&��u�M�[���#���$���x�4���/m眡g�g?i/��2����ڊ��a�r�D[a��3�/��:�ӎ�N�T��=G�^ZUKZ�_e\���������~��?cG�Oh�x(n���r��VNI�`����塀��Y��T0]b�l�o�)�fJ��s�l[�G�V�P�ȱc�}뱺���>5U2m�_N�Өh_g��j�����U@s��~0��N�<LS�8�t�#�r�4��@�d�g�þ�Z�9�@ʔ����8����Sy�A���h���oy��_P*��F�U����������I�J���8�@4ą���^�)o+w���j��<�!�Ze@�s8���-��!x5ݳOg��n�seR(�u�B�d{/�/���O �+*����C-�Cb�yJ+Ƞ&��5�9bTm��ЫF�_�����)�4���~GJ�t�?$��Qrw{h�Ve>��~�ذ��t\?���N��8�
�a+~�	1:)_���1\�J��k�������SHG<��`x�0���.�Te�f�x��{}�Q	�"��<��Pj]e��P	�I2Ee G�8*!�����Τ8SA�L����utEݹD}JO��v�TSɴ�i#�O�n�g�6/6�ŭ�s�����`����Xw׮���' X�^���W[î��؉k��Ns1XG�lPP�\�DI�o�J�-c6�O���X���z��D�3*���}p0}���zaս �o���#n犫���N�KCmn�l(���E�a�t��`�в��!Ϩs�iG�� <�����ucȔ+`�x9�ވ��b��4 �E��`�����s�~p�*q�-	�3`W�*P�3��:v,%��"��X��j�d-� ە$��X5�V:�
8&�am�x�[]�NgY� �h��oM���)��s���ݓ������G���3��t��EU\e�(Fd�O�qڀ۵?�?-H77�f��F	s��<�B( y��$Rd��vL��
R����%���C��6~��xB9���'joo��Y�d��v�J��*�n��q�\�'�d� ���e�l!�!�qk�h�L�	����}���π�����%jƩ�Yd�ο��\G�������%@���h� ��6QE㡟�b�>E%\Z��'��K,s����Ϛ�0��L� \��x���E(���3F��N�=2arq�	�˃F���'�ֲ��|�9�nl��=7]2t� ��P��#$L�~$�>
�L�ɬ�$&����Vrm"QZ����M�^p�]�Dl�)PR��Y.K4�FN����=���5�.�wiq�Z�J���8�ׇ�|�˭O7�=t���G�BF�1�`�9cXN��ٯ-eT��o�C��w��z*��ς+e�i�w)I$�$�(��l~4�9��Kk�G�0)���e��ʱz̖����,E����*�fC���-̌_z�.`�9���p�VrT9�0dÅ佞���Nt��)���h��d� �O������i�ڂ���,�����+��z�i���|�[r�32_I8K��~�}�SX�^����{�_�W,�3_��v��=}��bx�����~��hy�����Y68V�E�J+vSc��b{hv�{���ե��M�_,L_�Dǰ�V�ڭi���ݔ��c�j�o�`�n��5#8���zY�e�R�]��p��4�n	d��c�M��(�0�h+��y�@;^s�5�[cJ�S~�r�PY+W����Nn/�D�@��P,Dt.�ڹ�0BM�rdR�:c�
�E��A9j��
��P!�.����?.vؔ�&/�2�J��7sfЛT8�����N\�)$bW�:a����c�T>��rC��i˭h0Π�5yU�c/��h��tBIA�敡���;��p�*NF����h��|k�p).>��th�kFvݠ�3� �6ڀ�������W��ƣS(O�y�-���	���"y��W�ӄ-�Mp�L��RX{�e7i�nP7�)�;o��A��D�!�U�o�y�ת��J�ev��w��C��bS���x(�$�E9�������6͒է�b^0�1�l7%¹vܺ��~��L,�'��M��)W������y_���y2Ogɻ�&8k����CS�ɭO1���	I}�9(	>��BV���g����1�I�A5#,�	�}��Bd��h�Jf⶜t�Ch�6��=��M˴FGs���F�(���<�:S��l-H7�&���|������|�W/⽺��ַr�ݯ��j���#I���^�
����?W�l8KT +���{5k������0��{������i���~�ї~3�P� �����XfqT~+U��϶��lP]},��s��9�������t����8�T��[-V��Ɏ2���m&ݴ1�ӧ���s�d��#�ȵ,�ÓYXk�����<d�7�9��h�gOYec�= �ʛ��elN[��!�~�2�~!<��h�1��Nj����t�0I��@R<	*P�����QΘ�8�Tc�O��T
[��.��E�Z��)��Rs�j컱�*e4<���F؝C�\��L�?g���p9�cp��� �,�=�\����o����$��ҵh�=��V>�;X���Z랹��x�> �l~�.����gZ�E��tD������|EO�� ڢɶr��o���p���S�h?=��U1�>��քz�
Z�0O����������c_,F�fh��*3>r+��7U�3�_偞�5����Yv��.���*��LUq5���-S(?�r|�+�/]>-(=]��W�$������B��q6^q�xm������'<����'c'�����"��O2R�C#��`���{\#�-v��}��ұ_�[G
$�v�f�T��]�@������g�P���܀�g;�Snm.\P�[�6ɮ�ZK�u�����%`}	�3�"fqi&�{פi��W6���J4(�i�:���#�����T�V�|�n���Df�墚m�^%���џ��W(u~~[�"�Dٷ��e7��mm���[����ӽ"~�
���dXſjq07p1�Ic�o�<��R�7��:u��&��x{�.�X�<J������J}.�]��S|���"�"���F�-h��
KԆ9��P�&�/A��޶������#���k�����zY?4D�š����JG�vt2����'/a�LT X��ֻ�7�a4Ltw@���C�M_d[Y�r�Oԛ$Lo�{u�Y5?ȤZ����f}�����IVYQ)�8��E���9��)[��Kmn+�_eJ���k��q���id�|9�/��^uhw�-qk\�E�M;S���ja�;@F〨�/�d؅���˦�	"����d8��Jnޘ06d�*��8:Ê`9,uO���5o�`�q6�fs.F�ȹ��F�J��\�]��g�3
�|���f*��_J��hTbU���;L��qmS2���o�(��s	%8O�P�U0�
�y�G3M�̳����E?l��e��0���+�^b~�G�%*r}�jK�o�QO͹I��#�Ƅ���ѿ����̈1�O�=�+~	�'>/F8���^���8&l���� �嵯*;�w7U�;�3bj͇4�BlX�'j#�,��bںI[P~+]P����T��ȫ�S�n���(�,Ҧ���2�9W�h��N�*7�g�䐓�bj��E"���\ ˄q`3���6n�K���c�0A�;P���&�L��c^��)�{�D���J��фj5�E:`��P4��b����3���lɷdav�M+�/ՊΙ�p5�x��K�� ��]!Zf�b���q�:�>7�c�](����Ҷ�v�����U��R��ï1���U�&����ɿg똍������0�Ykn2��o��~T��^�\����~�T;Z,01&���ɗ�i����.��Id_2�2��\�t�����ٷ��l4PLN���rR�d Z��s|�h�+C8_� ǵ���	a���񔾖4���d$y\��-� ���Wlm�<YB��t���|��݇��ʦ]�T�����b�~&.r��*�{\�(y���N��pm��G��	����D�)��{a�
��#2�Ї�+���m-��\�w��حÖ��[+��ږ�f�,�*� ���Dv��@)��ׯ�|���Ԉ� �S�����s��-�L9�G�cb5����j���jrfs���7@�v5BWmQ���ؕ]��5kƷ�m��tq�ԜOV�Cx��S�>�X]`F�g0㛦��9ߣ����ƌ��>~Y�|~���7����X�p���gVRa�S~��U��b��na��~� fm9��i$��u2����ѣz色�-D׀�F�hE�|��|T��zBy��E�x��ׂjs8�1�����h�|�Y��%:Qڳ�~��-k���t�o��/	��*��{����-��j[�Fb�g;��[;����"�xe;��{����5	��Pr\8[��*��T��1�u�\0z.�ݘ𱪲�����&J�0'��d��.~lE��)�=����G�����&����hH��z_�x䒌o�� ���~�O�����J�����*�۸��p����7�)u���Ax��{���-�-D��
l��z���+מ���66��ֺ]���
e�?@p%��k*}� ����ʴ�o�`L{���X�Z�ĉʱ>R���5��Y�.a�mĞ������%�ns0,} �  ��8��j����w��bOT�b9�J�R[J_��������w�垉��z�`�9��5���]�8�c�N��]V��dgZ�ǲvL����҃,U∔I���#a��N��Y���\�������ɮO�X!Y��=P{�c����WI4A�3��]Ќk*-�W�Ҩ��oW`9�*������׽#©:X�閺=B����W���xY�>J('�B�
:%dN|�s�F�(dC5*L<Z^U�����'�炮�޵T�õ��Fҡq��]�H�>���V�D�	�'S���O����ܧ��}����#5i�aD<��[$��*�l�;M!w�?L{�{</:jjs�����+��@���TF�p9��G@���f�9C�H��@͓��2��'ʿJ��oͦ.��8�y�_D Z0�b�|��뽟	dn>I[X=����7b4o�@t�>�C��� �t4qq��a�W��?����v�'|<��x�cl�Mݵx�-J�F�-�A��|}�$�{8k=yh1�l[��}F�7��&5^�D���n���|����sgts)���y�F$"�Il�"1H	rε�Faԯ�#� �z#����[}%�o�C�Y�;;��|g��� 	/��9����7&�Ү�kA�	0��q+6�#%A�!��(���b��� s���Ȏ٩iO5I�R�|��F�zn�5�dF]���t�Ω3t��~��T��"5C�L��G�~��$9��U.U���+�赀���c�rsH�}����6�96��ZN�#��?�s�i�`?.�w����̌��r�뇥��t!
1�?�6�p�N9�VXp�?*O�݅F�sx�������3ܙ�E�� �QGQ�B+�tpR�`g���-8ݿ��r���wo(8g6a����YAC���D~2�R�q�AC%���{"Σ�{�,-��xx�?�UL�AՙN� ~P��=]��b$%q�$��F��Er;G�����h"�����?Wu�z~��W8uUe�7\	}_��A�M#���Uw��o�e�>y����r�Pm&��!u)%������VX?[���G�n�Ud����9w��H'��\'.b�ӛҪA(D��vL���w v,,< �p���ba���T�6���8na�3	��N0o�A��d��m��D�)S�	�/͠Z�7H�d����`ն7�D-�a[���)_��@; X��"��`8H[h!�����Z:ӈi^�GBrr�~rnh^/�FN���Sʾ�誠8���{�D��gՇ���۷�7��F�P��c�fV�5>������;���E6w���v����py�uӭ�O���MM%ӌ�d+{Pd�2�|t4!��Jsg_+��N!�,X����_]V�Qj�*�\����
�)�;��\�
����1_j�j�#%�a������m�}�09��:�X������y��0,8r!�عHȅ�eeh�F�3Mp��C𠓰ʍ�ܑ�����d����"�'� n2�>�/��J�/Ѹ�be����ɴ�ż�㗭���_.Qta�ҵ����hNc-~V}���x�<��H9*P�5�R�k��r��9��w�6�6�;&!f��k�}�D(t���d�@��0�㲽��(6���XU$���C���k2U�����Ȧ����m�%
�s��Ͽ��AI�m��8U���@m4��lhM�E��_���ґj,���'8��?,�8d�j�Z?:^�i���$�eؠ!E"9I[�pi�oE����'�=-܀7�Λ�M��� �:���h@i]h�"͑�Z�������	��B��1\]���`�s��Ih! B�a5�s�� �}�"�<��9=�����Cat�́�!CS~�=��5c(p�u=P��
�
��0Y�t'�&a	'){�w�2N��K���60�\v�`�� ��Ӷ�~�%VV2�B�����I�(�~���g;.U�X�T��,��>K��X����˥�t��E���6��<�fn�=��+~ �@U%g���X��"Į>�-����dbP:$�d�1�]�L]Yk�+���I�+{��9����3�~WB1�i��aKX�Y ���qa�#��u��9~<�=kN��4������.��}lE�m�����!��9�DJ&����tvs��Pe����=��q�%lT\}C�E3_���y�\��X�(���4��3%`_e�C����Ya��BQ��Qt�x�ԭ�行�߭�r�����'���mhD�>j�aB���1�'#�1;3��668$��x�QrE\&��e����xE��l���_d�_p��;&1}��xvl���/�HB�;��ED$�%(���b�+T!D`��ld�&�ܒ"��¢�@B�s�u\[����8��d����-90A��bQf�|���qì������{G�\����B�O����iTo|�%r�B�����S�e͉�-���Uֈ�V��ƶ(����
RW���>-u��=,���l��E:i�8MpON��_~�CV�v���~G����`0���c};�-�I��ֆ���V�y����>b�N�;�+�9��\#�m��4�����R�éc�~��4\��2-�5� �����>�f\���s��m�}!���u�D�}(B{�Ī�o�Rgv�2פ5�Fu�:�M�=,Ũȯ�_�uU;Բ�G���%�����*�����S���D�,���Ɓ˳��h�:�Y���(����?Gc�t��a����՟�<}�^Y�Q��}���!Մ|�x�]633���EAA���R=���x2r�����t��Z����fM�ڂS/�T����&僿�Ŷ���ʞ?V��jh�'���#��;�0P��G�鉯N�V���⦂F���}��'VZ��(�E��^��'�JB~k�=��'��ߖ�i��2�0QNF���c��vL��L�aTM���Np����%"��D|1vØ?�M�ً�YO �,3�K�<�l�x�!ܠFF��^��!�;_�T����Pds���;��S=S��{�N(rq�S���ڟ8�j> ��mu�lӳX�Q��7�d�J�ӻ�Nrw�D�`@����#�蘌>\�=����#����*U��/|����?Ԏ�[����	�r8��4;�ֶ���� /�M���9���J* ���c;���W�l��Ȧ��� �;�@��<��2
x���L��|��=�ueP2�P<�|v�%���z>\�!�\Š�v��[�Ѱ�E ���ħhu����f=�+H�T�wYR�O3S@x^7�O̸8Lٰ��pKEw4�K���E�k4���q�^(^�5U�l�L��~���5���3�HNe�ƪ�j:n` J���J�Oň�k�~��/�B��Ԇ#jl�S��� �^���A�����5B�MO�`�/V�#ie)�C @(X�6%F6E�}m�Ikv���jZ��❒�l��{�"��-l�r<�>~��o������_�b�w+�Z3b+���SNsBL9��N:Q|�	|�04��5�R���4���s'x?�KD��Q`	=�
e�(�v����]���
�쬬����N��#�^
DM]�?���h���Bg8Wt@ t h�u�
a��g>Kk����'����-N'����ߗ���˳��v�3;Z��-:
L�u@h?+�7:�,8@ZtA�v�0d��%#��ط�{�*�5��R�m4ҝ����5��A[/� �\��!�D�A��`w�s�mF�,�ZKt�UɎ9�Y��60��k'���D�XP�|��x��̥��2��R�7Y�}	_�ȍ?ϷJ�Zc
�e�Z�Z��*l}�#�G��RO�#�hV�����]�j��d6Y_ v)��~�p��1�xfi�w�?���1��N��	���H@�t�x �����"Nq̿�se��j��	��n��$�@e�Y���0��O58\�ҭ�Je��שcF��q�M�D-�C��;[~�-�
r��;@ø*�&�?��K�$V�f���&U���C6/��;��*$�D����p+ �4�?�|�iT�	���,R�.l�>ؼ�<�G�@�r,d��������*������,���`���iN�-�]�y)R�^�cQ~��5픆�ȹz����u4��w��`�Rt��!��{����42 �ߩ���o@.��N�I�щUoBe�N't�?�rt�bС�(4w�b�D���	o�М���kOZV�'��93}�5=�Mե��g�D�+s�Z_B	��oxeE$p�n�Rm=�hE��u��do�Ư��w�����roS�hQ XG��{��8��������P�L�Ջ�.y,i�-���	�f��@�v8�v���6E���3������ �����~uIs���.I�R|�.k�s0Ĉ4@�7r?�ȷ�B+�!p�b9��F:���ɱ3R�_���q��A������*��.a�"�H۝LT>����03��i~D@[�Lm���\.$�!���	��4Id��`K��4�p���,���.}!���x��ƤL���͆A��Q5�Gb�h��F��=P�b�����~�� -;g^�n���*L�!�	���Ӌ���;�!��yH��_Y}�f�ۯ�%*�)�'᪌T˸���r���H1���nC?h�ج�ꁇ!��߹zeWUҩpl�װ:z�8G�(fc��[TLø$i�T�#�!�+�.K�H�β����wDT�=AZg�M�EI���m�.7�-�߸�!����9�e�pG#���/X�&��ț#X;7����&}��k=.��N�����0���=� �9VAE��3]�Pq�p([#u�Š��N.~�U�5����u�f���+�ޅθ��T�.��;C߳��Cj>�U}�([�hdA\��=T������sQ�Q{=_��Rh9|6P%̤��N��a�S ,�q��P&pkaj����}9��]�K+Z�lH��a&ۓ_�!���O, ��7�@jy�9�z�p��5�J~�����iK b˷�3s�{{�圊ݵ��0� ۑ�l73S��wD�S�Y���0��iJ�v��[^7��V��gVy�)�P�l)�(��BgU���PN=� ��/o�b\���=��[�Z>��G���l�7��lsۅ��b?VZD) "�1������j᮱�ޱ���m�p��[گ�f�|c��� 	A߭�jS�Ԯ+X:���-l��:��44�[6p�#��ǚ���Er]���U���-z�忋��*U��8q���6I�4���[�>��р
l��k&�P�/:�j"e�ß>��Uz�G��7��`D���p�P'���G��41�g�"�7���y��~J^O;��v�.� 喚 �{�|	�����!�r��X��oZ���0*�*O���W�S���DV�;�o��g�B��-gJ|W�ZU��o
4�\�7>*5�U��:DU�[�l�dд��~Euc�Y����n�	xuD�����4�$�m>��T6:(���,�6�e����I
<�������t����P���~�B�c������0�]�f/�`�ow)�G"}��MUJԲ:�.6����5GO�����l�{���{=XG��S��s��J���/�4t�n_�],���ZT���7E��t�eĪ�1v�H8�x��8Ţv�+�$���d�do�4!��&�vM&�z�����Y+�t�����n}=�[�螡 ��Ԏ"��	\}%T[��e�����5�j�Cw�)㞒/����XO�	�����,��툧ͥu�b�;z��騻-�*�	�%_����@q'-vB0�i�.�Mr�x�tx�<�� A�j|G��܏M3M5�����Ue�,{F?�f�k�ex��OON�TrS`ŶE�P��8]f	��g�pc����`��#�M��ѕ�K�{��~� $�L�t��q#S��c&dv�|U}䱢EE�BY+ք�(!��l.�a�]k�<�r9���0e�I����4_�к)�}ģNpT���rE1J˝C&cOt���1T4��"!�ި;��1q������C�v�R=�6�F�2��n�hdeF�r��t؉ZiS���ފ��ҧ�Qr�3:aA	��OMȣ{���XO�%�su��a3�o����}�bV�ߙӘX��dgύb�{y�M����oa?`z�����_��>�M�H\�桍  +�n���L���M�}&�G�fb6�H<*�g�:j��4���P� ��Z���ا�rHt�D�m.�%Uh���u���Ru��9CFc��{�sS���Dך�z�F��ˉ��w|̃M�C�ܠ��q� q�_d;�P�J�}�#����z���l�[�?(}�C�&йD�Y23��{�@;F?�vsx���͊~��';�
�e{!����B !����׋��Wp}�1J��h���:/��	{}�W>ȹ^ d�����pc���@ڷ ���R�*/&�r-���p"��'�A�|(������_�|�i@"_q���\&��b��py��=8��HQ�Yu�������?�i¹j
���3?�rgj���v���~$����"�0�\[���Zu�G�t�Ci�|��7���0�N��)��0��7�;U�^��T���W1�2�nAP�׊B2��ב��c��3����4�/m��F�!�`}ye�_9W7�¥dP\����M����7��Lm���+&�P�`~���#z��z�8Y:M���/���&/����yꝫjj�D�������110���(!�!~���VҮj��L������E�ΦX�	qPF�ݙ��b�h`#��>�3q�N����슐>�������K]�����Q����Iн.�Z;Z�r�>.��v?��\1Cq4	G
1�i��,��SuַS�@�/��\�Fu�#s��cU�[���˓P�=���8�� *Y����$h�r�	|�k����ã쏲�����F�Q�m�)2�Pn�{#��E�E���K�@�Ј�9����v�N��s��Q�e������|9Z��Q�,H�4���+l_h��ϡ/gS9��ݾ�_��k��J)N�f0����YʏH�g�2�Ġm����m��0�݋/Iv��}��	m�ڠ��L�mn�Q0��w<���M>��x0���T	����t�]B=�流8�9�ab�Z�;�֡Ou�VI����Q���(�B��
j�s�m��@�yja�$2Om� ࢮ
�7e��	��S�g��K�TkP�'vpU�ڸT��kvyɎ96�ɋ[���mA*/�0���<fĤ���{��R�j�຺���1�Ct���#��<B&�ʀv����֧��_�	m��3�D\���ta��yX�3��3�o�89Ue��^��&�d.6�q-����(v~�@�U5?٦�E+����nR���X3I���H���FVr2"=�����k�\+�j]$��v:�'XV�R�~q$�-���k~ݙ�����4Т�d�W&x�?`\�j��)��5��g���3y�"���Ab����������h�G!$�^�B�qKNz�aZF�ٺ�Al*�L����{��a�B�_�ˑ�/g�·�W���5^�G�N{�����E��e~2ϋ�V�.i�(N?
�XY�rt���}$�a��'L�|-����Hˊ�J}s'<������k��0�f�CL8e	@�*�nj��*d��:9_?�ժ���>-R~���X�8��0��~*��܋R1;R�˄<��bȋ�����$i ��Ԩ-����<��x��T�ǵ����������_#ħ� �9V��7f���
/�2|�31�L5���{�.'I��5@�����=�1�d�O��Q(�@!kǳ�gS�_��z�v���\�g����!�5b���]=¢�c	 �����o{��mgW���C���7���䲶�ɏ�p��㗖]��.�����3��=��l��/�|U�����,O�`dj��:�b'((j}m{�o�G�f:xf��t�ƫjU���^�H"?���2�y9�C�Kt����jO��^г��cK�羟�R�H�%�������V�"� �ya>|�0��}���8B���0йg��0��׌`AM���׭��Ǎ�.�	��Z�����#|> �N){�9���ہ�BtY�)d���r}]|J��0��W���(��^!����Rn͋�V��F�wɚu�҆ zO̜��S������D���-0��J��X�n��[o�5_u�A��F��'�C�X��~���)��ɾa�h�ϛ�~��^��Έ��<��V��TR3�Y���ۢ� ���r�N;f�i��|AN��Z<V��$/c��u8�%�i�#x��C�= �=�
O�m0��hA3?��a)�n���#�ĩ��~,�S�(���;Ԁ�W�î{aH��`�T�wه�!��c`����e��T%��R$,�4�:�8sK�Z�����s�z'�����RT��J������'���~�l�v=n)S��
����s��� ǿ��Q��iv�G�̉4�}m��Ng�������%	�qܵ��g�m�q*���0���7��\G�II��e���U0��}b4��b�H)�W��!��85>s)���Z���l��|���m��H�}`g�&�9V�W1�����q�&�zZ񄠥�  �Z�֙�T[����h�jkQ��0yϩp��y����uP:'~��$�����sZ��.�< �aɡ�����y�i϶��ԓv�r�uAtT~r��s���6Z�����/¨��v�{`�6�R��G2f�;x� ��p��ƥ2�|:�с49�A��X�g���f��"A~�	�L�,����� k\%	�P����VuVZhL�D�C�s[-߭����b�~���3SZVE׷~�q:�ڢya�u��/�t0�����E(����1��ƞ�疥JL��
��Eb��F�2Mm�����Aׄ_��;Ĵőxy�Q�=4�4��kbn\�{�A���u���2���M��'�D9������G���\�P�g��������L���b>��B&����)f��$qމ#m
qm�O%>��J08u�Ct>y��o��t���R%X��cT�������
�ޭv[l!�b8w:~�v\+(����<O)]�ӷE�մ烸X����sX�h/���Q+z�$^HJ�A��B��B̛��b�u�zQ(�u�.��ѱ��'��k�OM~����M��fi�0����CK�Q�6[&m��b|�S+Y�V�`&�1�B�b���θ >m�?cX`$@�u=(X:�?*�e�2��H}ߏ�2�M� h���.���}L�_J�zfS�x�@��w�^�������%8UIDp�R'3��C��mǌyq�ز��u���RTi���5�D�(�lE���|��D0��	(i�Lۍ�fQ��w������t�O�e�0�|�_V{����kl��Jj�8�lZ�'���vW�Ql�4�P��Rˑ�/�*�%�a���$���о�CX<����N¹��z��^�-��EE�%;i4Z	�"�v���vͤ�iv��=T�O�������wIPۿ ��GK���a��3=(��eG���J�6IS��4;���.��Y����`�VyuW��͈l~���^�[#���� ��&W:ɩ~S�	\�,�8#v�G�fL1w�dE`�]�Ԃ�r(��ꡲP6��q���ƾ+Eh��r�M��,��;� �r5f��0�{���¬Y��Ԉ#��u.l�����	&�f�������Q\��0W&f�����s�����E�����k�%�k�ʁ�D�R�C�:	���������탎hc(Z5��D,V����h��&�6�
��x��I��j��pJ�U���e���pW!P���e��t��n������1��F�T%r������^ź����������|>�5&Fk;������*8�V�ܖ��]��3�	��j�\� ����ܰ���AD���q��IL����[����]�>L#�pB�Fq�1Z�K.Z�����R�$:Z���}B�f�<�ń��'EW�c"�ᰬ0��q*��}� �oZ��$���ۍHR�c?�	sAŷJ�#��1� _oK;�@L�anH�{bȩ�*�B��}��:������'?����@�o�jS���)�k��u�Շ�Z�q��i+><�2%'��*�V�SNH��C�%/|Ɍe��Q?Ox\=�������4V:a�:i|sj-�ə��פB1el�W�'�1��L���ڃa�-Z�X #��r<�RCy``��z�t1��s�pWֈ�Ӈ���>ХV�=�	����7��y�ec��N�>��n��*�'I�Y8`5�����d��-%4
�g��z�槱+���wx�\�5Y�lA�=Um�p�l�y�
��݄�#�u�f�*@�\��)�k�� �Y+��"�wg�$���T�K�HM�X�5tk-'.���M����m�Ť*@σ���c�t�X�j�Vy��}�<��}�.N6,��D���^�lW՜ʏE��{�B���i�u�7��i>�𚆫2��8�g��S�*��|�k܌b�Î��_`𹽄lH�ʞG�mo��bt��9��7%u����A -,�$�{����X*�l���DHy�j��i����������)�[�^�MT��M��T�Ң_
���F~���B��=�ւ�9�<ps�n��㞶8��߬JK�2�[��5H�xO��:h1�W9	kw�(|��%���#�6������`Ѷ?+�#�θ�Q�y#
Ѡ�4�Z��/�Vy����n���9�D���8�vs>�f�9��0�߀�Ap��-��훜���@�4AAY��'�爹{5���5���R���&��k��,s�D��v#�d3��kB'&����W{"&W�0T��5x���pȓҭn\u��ȉ����ߊ�i�3)z�B�fϡ�OE�w�kٍ�"���yA{f�Hi�->��Mt`|	f)Gk���a����b��v��O�Ηhˢy��YZA�S[��ɯ��Y˖��E����x��E:c^�v�۹�V#�P���O�����-��p��u�'�f�LS� l^�Øw�ٰ	}zO�0����ￌVQ�cv�/��Nv5N��=Q��J:�9����j�8�][T��i�r�V"'�RL��pE&k�7D���[q$�9�5N̛@��C�5�L"g�\b�7,Λ62*��lMt���w�a����oB��5�֫a�F��J[��9���*�����C��j+¡��*�
�q�p_�������)����~�?�	�tmd��M��p7'.�S��.��I�¢O���BD��~���� قj���⃬7���j�cC:9؊:6�,1W�al}��Jy��� �#�(�T^ƍXP�3kn�}�o�!�GQ�3q׆	��0�2W�j��h�+m��[�Dr���7a��V�'���t8�I�
X��b��԰��L�]��5�n���`U��-�mƊ�<���E�%��g�����x��e�B"�Y��.�3��ےr��ǫ,&�8�rH���Ǐ�e�sU�Y���;�����B�z�ᣗE6c�<��tu�=����:CYGG�B�F�6L*
\�JU�0Y�������X�&tx�M���'��VR�����`O|����C31���-~<H�س�0�`�d�]��#�	������1˰�y�4�Oя<�g6ъ�0���>ڒΧ$����Ki�SИo;'�t,DU�+��7�����4��\�@M�a.�Bv沊�+����T���ri0�ק��(�YK�]��]	�V�a��=�n�xm��U���đYRP�Q�W��� �D6P�E��#����9Q��h�Y�ˠӚ����Z�V��2i��='�X��OgQeUC�x��?��ws�$�~��ڈD{�!��"���x�Uq�^�̍:6U{n>���r���>X����9�Qqu�C�=��� )�z���V]�<�YCW�BP�f:d��P흌����R�^�gqO}X�sk����NL�P���[٠$J!R5M�+D��~�!��]\��:J9��@֩0���b������k�����(4I0�r�{���ϐ4H8�Sa��tmN�hcb��\�d���.V�j:ڜ��HR�i��l/Fy]+WG��W���qK�w,h����gʰ��,IoU�a|�M�fϺG��vDS��P#��h���n���� ������:��|w�o^�	�W�{s�}���^��{�SO.F��Rb���!�mʋ.-+���wܡXҌ�͚S�~�zNA��&r/��;�f{daw>BZ-E�ݏ��f����9�%�Y�?ܘ�J8�'A2���h�2[4xJ}���/�n'&A�a��Qa<�׈�ը��cz	��0����+��(T+��<�/"�y�v�rߧ�5�Zҭ(��LP��b�t�/u�Z1sח '�1f��<�ϖ�.�M��j����!��|�z�}_�:�dK��7/�����=�Ef��[
.[�$�`z�i.\uD����*]�}�F�����W�a��RT�]K	����������(���M�{��~6Ƹ����p]�.,�%���.��+��*#`Xyһ�͟�۞�yJ\�wt�*�0d���x�S�)(�0)`} ��i��R���`q뫵�^Y`���O )W��p����v<��%��Zv��ɭ��� �e�換�4��r���PW��C�Z+0�p��ĢqU�.O_s��h�D ��OץRV�,w�����_�ug�c< ��w�i픠���{��$�g��!$F�r��.l|���̔�F�亃7@*��U
�����ux�l8�"cM���;�T�ք�a� �ʜ�Xi�6�^�l-���ʩ�OVƴ�8(�110sh�x"�wi�����b�{X�tS�p'X���ȅ���K.����F[zCH�T�����0o�qhɴqR6n6x\i��LE=�.� \��g H-b9VI��
.�Y�u��:�cJ�0G=��g@��-(C~�4\7)�H񼔫���$�L�f�M���#�SJ���,�����Hj��>��+��mKY����ա���6������4w`�*�OM����z�.�N����b��'�yPQ��M%������1���'�]���G�Dޡ������h��l͔�*���&��K6R{�xuc\Me�LH�\�G�'.�rY-q��u�~+�+垻�D��I��I�Q�j����@=�j=��8��p4��O\��ܟ���Y ��+Rz�5�O���ii�ʿ:5p84���篝: 5����dvW[��DK�C�<�����e���"9v��K�:�Īmu�}��'`
l���#}�NlB�_Ku���v��0K��?&����d��ƄW�����!+,��XAHL�l6=�<?Ns7��;���BO�w����t˭^�?���h?���[������e!���e���v 
�:K2�_� �!_w7�U������tn��~h�G���b��h w��t��
�4K�X�J��T*Q ��6�M}^��P��[�nْ�T��``eFO�(,KB8��1�+��j�g��Ar�yw �� ?ަ �u�D�-5��R����[-%hŁ���k,;�c�yH�U��|�Dk��Qtb-����k��T��d��ɗ�|�`ˢ�&$Ĩ"�P
�AZ������.lRk�Q�,9ug�kHLGQ���Iq(�]_��g��t�'������������$��� r	㱱�#\�Y�*z���B'�k�RN"j@.5��[S�,f5�>PQۘH{B��E{���v���$�U�
"��.��|i�gV�o$�O��8�ps2�c龔�[;��x��_?K���L�JS/8����,�҄��:�� �����דmrCKU�,��=8��$4P6Ĭ0���D��.[�1�����`i�C�0�~d�RvaȈ����"�b/��^�5&(����`;���}�
�;�}=��<΃+���|WWO���CJ$1�=/�v�@���ܕ�{�Hļ%�3����.�5�p�oAikT����#�$�82ǘq�Y��⌄+�H$���<�2�	mV�j뱷��P���[M�i�(��Zk K��U#�`h�&�)�Cb��/�++�<~Y�DƱ�A�V�庘��uU�Fk�i!����A���w9�^��i1xH�J���
S-���7FGȝcWg�]g��D3΂?ڇ�"8W[�R)�:���=�N�k�v��1������,YrY�����[��p�}�w�Z�RJ�P_3�بm�t|�F9�`c���<���Pa��/�:.�_IT��8��V������r�eQ<�������Q�ѣ�;��I�|	���2������sh�pep�q��7��l�����'��YB��B�+,3�m� ӷ#S���{[!�ǀ5�	dD~�׽�ύET��|���0t��O�)��_wOj���fnF�\�N�0��Oŕgy�q��<	�5K����:C��	��!�~{�kGg��ɴ\��MZ�oeżg�&s��cgG:Y]�J���9_��	����A�Ϛ��~^$+���!It�1�L���9�/��aL�����Ԗ<&J$��:kb��=�|�?�����vυg�j�st&���[ C(b�����U�ig�e���q��u�/��c��dJH��.�)]Q��ojb�
�Ƃ��	Tݥ��������P����~nɈnQ��S�v1��E�baԍ�F�g���oy���l�-�������D+N�^F-7�b��B�hr�ش����j11B�5��,B�Nh���~�4"z]�Y)�f0$NVAp0љ�w��&<l�d���$��Ww���V���$�?�+9<��{�S����io��i���T��/ǡ�{/1�Pr*J�����#Q��vO�����Θ�2`�"J�%�rsk���/��Xl����#������r��,GIfَL&?���z��ޟK���t��=+�,&/G�WT�Xzɚ�����P�#�2?ҙ��H�s�+�e0q������}x�B���}.�fKk&R|�H���^-�PU �a7��	����	T��c �j�,�뱅�X�ϩ��=c���8�ZX���5�r6Lzc���ܕ,����d�t�>]G!z��a_5�ɋO�EN#G��R�Tʫ>>�~�� �n*�Y5�-�Jp�ޢu$d�m����+�v��//�P�f�H�����:��� �����i���XW�x�)���������P߶�?�����(!	=)�CQ ���<6�l>9?��7n�}k��t�����p�&�����Kr�C��$~-{��0���#��v�BWm�
9x��\-�}��d����+�o��б�`lX��Jpp	Fn�����Ϲ�J�8Z������h��?���#Laqڽ����WRPP�BÔ�L,�f�:�N��C�?�e�����Dog
y-��pQ�oR�&���g��΄w��F$lu(�w�|>P𑌴���(g�I8T&�
N0�AxB�r�E�0�3���!����7�k?��D̿d�A�h���`���snx�ļv��B�2�'��)��?߯��QMV�����ّg��5NN��é�g=0�IGU�'GÆn(�ӯ���-"�d��P[Q;���8�/�n��W
t'��ߦ�^\K���D-�����RnYW�e��O���(J�ީd�4
���mƕG�x�J�~"t;+�����0Qy�i�n�V�"�]ķ䏤	6͋2h�������<،*���b�E�e?x��g�a�g���v4*D��P�&~5Է�p�������ys�7KAr<�hOHO@#$i�.nx�l\�{J�Z������O���vX���.�,�f�Q�%65�b���s�
U,/.�<k��zAO0�;~�#U��)�E�ys3t����r�����w^R���l����g&�4�J�f�-^� �k"h�QV��1{�Qk�W���;�I��r�V�'��ߟ�1��ވw�=�6̦ђ}F�1X3&�歾�l^��FD�-�3���UԲ���9&�`+����ì���,�|�p��pm�{w����||�K���Nذ�3İ��xFT�i���!�A$��
����ٝ�8VS�*��V��%�{)�嚉2�)�蒯9Z�\�t���wdf��.`�@%��}��#�]a�n��q��g�Su�I%i�R.NR��ӆ^ ߊO!�(��c��Bۈ[����f��v��Xo�و��g)�BO�����n�pu�u�j��Uc�'�GP˟I���Uq6i:��O���?ve`r*��4�v����dPG���~^�76�w0��QuwS����-P%��*�����F����*Ӂc;*e������d4H�}�A�m��o�R�
0y�z����$ [�)��p=N�U����R�O ��z ��x���Y���]���X�M��ed����~�I\���իj|�;뿊=�"���Gʊؼ���ط��<���?��]��lڐxi��:�m�A��>>��h�3�N}��zY��4S�5{�k��
 �%Oy��A�h  ���4OO�����&�c��ςz��y0>O8�7�J�Ѳ��/���A՘�[e�O�=L�θ[S���;�R�����^Q#��Ϫm8�9��λ��~���w���sܿ ޷�<�B��߹@�����S���QS��,�I���H�X��s��` �Ӎ
0���a�8)
j+}1�{o�H�/�M��&�J9"���� �]��6��x�x: Lt��C��?D��z�FM(�(��yҗ󒔓R��{�Ǚ�����ׁ�NM*K�C[Bw��]�R� �4ŀ��P���%qH@�v��C�.:<� f��K|�кu��tMU2	q�@���g�&+~�G���-]BV�����p�_��{n�$+�A���i���H@f�ͩ�~g��,���l�u��/��]8$֨���K�U������v�q.�$��q�-@@���M��.�<s]�G��Du5������ɺ��^E7 %�֜+T'�q�toW6bw��@V��b��U���2���7D��ۑG���7o�b������D�P�ۊ�C�\2�dKy���_�w��R��ʋ½�J$�imk�˸PYP�'8�4`��8d��f��n�L�R� �������1���Ӧ}��d��i��y=d�K�)/����d�*>0@R��s�(<v�|y
�mV�Gf�As����:��<��xZ21�s�LD�;�y��|�,'9_P����U&<	_�t��O�Iy$P��\�����T�ާ��p}�{������]Ui��m���y��"�w�k©�4��������&�ȿ�;��m:�X���KGo��z�qB9��*=w��;UU���,�k3$��u@��H��]/"ƤM����߫�=ŕ�z$j𶱚=���Y�1p5���%#�F�
�|�r}�^H�l��=��������I%_�O^ǔ���i= q��2a���Hd��p��(��A:w&��RL,(���Z�%%/� OA6&M���9SR$w���͐�L=��7�A��oV�e͊ƪ˚~Xdx)�ۇo���2�F�J��F��- ��T��F�!j]d�&L^3��-bG� �ZT!�k]ѹ��5̅;�WK�J��;-���]���G�χ��r'��x��D���r��!�Y�,��M��N���=+L���Iw*���ؕ(ɓ�ܚB�kIx��]�.~a����c�{(�MeK�*7F�8�R�Ě���D�MfC/��@��
�L���q��R{��ȵ陴��>w�=z#R7�E< J�\��!���,�w]����Q��N�p�v+|$��B�
�{�H�����ֹ��i��5�P���'�#f�y�Ȕ�&{$��[q���@}5�[�?��Nk�d�rA.)�<�X�ѹ����\��r�k��ݠa�\�72����H�;M�!ax���H�ؑ� ���I���K���W����:��Њc�uN3�?5X���	��旹�墑�p2�9��c*D���
�Hi��E��Ɠc�}U�*M2�K����
f)^�w"���N�xU�Y�zm|��^mu����qba(�Z�L��{6{~�Lψv���}
+��U�}%�>ɖ�M������V�DЊ���Υ$�t�Wd~�S������ ^�ٰ7j��B{�r�g[;W�9�굌�U���WڛǸ�k�@�r9�������:��ZO_�w2pJ�8�v�6�
@b������5e+�%F~�n�φɯ��ǿ=�L��xu^����,�-Б���4�*�9T�Z�}��?TWwN]U���SI(����n��*��%)�?DL�dv<��	~�;r4�ζ"+������/��7�<w0�ќP��X��ԐO,�gt0\A��7Z��< �m��G�E�	3ƥ�w�sE|�?������E�Y�F���[��y:u�n"(��
�5�H,���vѮ[�_��,~�V7��·��1i��i�SU����e.ۢ��#So��(u�<sV�K��2�X �6L�N�`��,��a�hT�����JA��[���fx�� �����\M�>�O�ǚ��
�GZ縯�'��mu׸�:�R֤�d%��daA�f���]DV����Q֑�U�%5l���"��]+��C��D��~ȏ���P��-�&��8�q��c_�?�#���6$���Bwt��"�fZ4��\�i�Sz���RU�{��TL˔�/�(2�+2�j�ױ�R,���č�d�".U�]�ћEDTP�UԱ>�縷���>teS��H�Jj���KH��J�FC�k�H��J��\<Vq}r6?V>����V�mwoM��Hő�Ϡ�Ĝ�K���>�>{a���4��� ^$\�X}1����]�Ct���A�)�r�G���7��Z˷���ׁ�,�#���>�Ysā�}��Q�:7�R�J:����
��T�v�dJ�:����]1y@�!�L����MO��vu&V���g��k��^��1.0��|�m���@���;�X��/�?�E��`�FAxr�}������p�E<H�5 �*9T��#�y�1n�����4��1^e���s=��>�v��
��K[x&IÌu� �@�]�]{�<���.�����w������6��B@ ����9���RZ3O�Ɇ�_�:ݰ���r�87?�U����+�o*국>�c�t4r��[��XD��ȷ�K-��]Y�:O��0���IW�,�h���;|��6z��b,HHK�v�k�����HE| �[4�~Ǯ�?�3S���������'=ϒ�J���VƴaoPb�x�5�?C��_�Џ�oi�.<�%���$?�A��#�T����?��)�WuԅK�9�g�0V}&߳9k���SJa+Nk�;O(=��߭�D5w�b��`�i	kdYk�Hh����Ǥ����r��[d/��u�0��֔c�zPp?9Ik1�R�.��x1��Sy�w����K��e�~onss;Ӓ��	v2�����b����l�l�:�2�|=�]��S��D�����fф��3����Gĸ���(�E��cm�w5�7�51l�+'���w���[�쏂<h�qB�r�u���n�G7!H��К�4^U��^o��',��G�:qR�-�%�43c��$��u3���+WO����3Ce���&�|\W��J���v�ZB���|�+r��j��H��$�N�Ds�Oh\.���pTq��l�ב!N"��S˕٢z|B��!*�η�b ����3�h����8fW$�_(����)���{^K: �4:ֶ}�[��2�<�ĥ�0���������B�ꔢ � JZb]D� ��c���F|��*yT��ʑ��%ܑ��V z�ʝ.�D��p��s/�$Wj���۸Q���f���)��&�{U�#��e)��/R<Ep���tb�.��9�]#�{�s~4���a�MH��P���o8M[�_?,�O���X�����o��+F&!1*|�7�b[�P�Gk���j��U#m�UWm�n=�l߫']�H]b���K~z�Ν,���TL���X��qiv��ԋ
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��Y�H�Ea�0o���0��C݃�ջ`t��݅fNdwi��Yek���&l���z7G#����}<�TK�}��~6ea��m�_`dGl���W����aȦ:��Xhc��)�^jnZ[aL�*���\�W�SAmO���X>���Z̀j:�6֥��6S�e*WjQ݌�D$<�݋����^�0�A��:�o�Q2�	X�u��V���\�	p�t(�F�l�#�~J1�H��������� �g�P����-����:jPߣ�Q�h|<l53�8QW@^�]�W�6RQ�W�m����&R��%��@&1����}t��E��ҏԇ�p�8������P=�Kd����O�ԋ	h%w�\j���A[����M���F���yoBLM|Z�13L��~�[��L��@?+yo�wz4.�.��	j�F"��"k�"8M$��Aŵ�S>�����R���ZW��H�6���[f`�ݳ>��
\��[g����̛���{'�kQSh�qi����|i����S0Ii�`W����H�Tw�}d�,�?'h������D\�P��5����3��(�Z�;E���*�O ��lh�F���0V�t7)]�cy�.��N@�b5�x륺�/3������N8��-p"��E�����r9C������K�����s(��������7F]5���s`��6���ӎ��N&�Lꝧ�c�Ҹ���n�U���p�b}�Y��4�Y����
1��Z5��y0��Lz?�7ʶ���Ff/���I��숙	�V�e!	��qMA��<�׋B_�-T�y-�(\x��|�����%TR}�R�3�k�碣����"'W�$��dMu�2�����%cgz��ڡ-��z�F�L����}�K��g�ߐԔ�O1:��@v1�S���c���&#5���_�ھu��#��{ �y�g9G��6k��0�t5�v��vF̜�\�������~��҄�p����F��<E�䯭|����_�&�]���������<�5��N&Ң2�'�̡���e�d��k����.�r����Z򘆤#�B̚��<��Xy
Z�G�f.T�<ـ�Y���U �����j��v@�ׁ����a8�"����+����܊�
x;_�0jΓc��	�Wx�:���k�0(�ʧ..������se����@���x	��,/tl�����8�Rp7=[�8|���,�½�PM�.�6����h`�o�]Y�m*ξH���	;���ü�q�Bx���G_�=*�����8�g�q[��zOB[2KP`�x�pa��+@�yی��zd��b��c������־����K�n.�&b�EZ�q-WQ�GxK��S'�YS=PD��f��N��q^�#���nSP�)7�(�2O+O�#����$;йb�|Di([�q�ю�GjN���F�R.-��]�g��]�*ßvw��|C�7�mV��	�M��H��-.��:�
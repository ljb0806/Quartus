��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��Y�H�E*��K��-��a8�<�L��eH�"� N�N�O�f����Ζ0z�{m��OH!7q��(^������,�<��LRfUCHj��}d�Hl�RbH�7"��	Ut��=��G����Ra!>���2k��t�Wvz�{���N�wSPs5Bl�Z�Վ�hG(?���� �Λ��i\�mu�#T6蝐s�i���(`Y��2h� ����-���c.��*��;��>
<�k�m��a�n��}3����6(B0�����m?�_�
���0��Mt�GhZ�w9'���xXN{��QCq,�i�7��rD��'�������J���I �I�8�]���׼�䝼�"�?m<�N���$�K6��k6|�B���e����Er�{?�I5&�Ɵ��g�o(�ď�g��!tC�Ķ���]_E�h���r��|7v��|�cSK�vtQP.AZ�*&~q�bء����[�r�Ny�;3?&�0�&^S09܈���\�c����¢��GUU����bh{X���/Il�z����y�<��3�T�H?����5b*P��!#X�Q |A�ZJ��S�c#ڭ,k�&5+�om�P)!��E⚁@<J������_�t}�UzD,�RXh��as��kf��//�3})<$��1�ζ;J�<v/sMQj��I�:#&����������,�m�������J���H�h�/ʷA̕��4�52���h9(=W���>i�b��9J�(ڭv�g�*��2�Q���j��s�d��8�9+��؝J. ّ��Yr��:=]��nXgJx��c֔���GC�[L3�]֋/ɹ�?�5^����ʈ�|��ڊ",��"
b^1ѹ	M��'��EmL=Ҋ�RO����ل@:��h���G/��v�����xE��
�[\�^��FG5��f�������v�KH,�؂�����r�s/�y��ǡ"桫�ٙV+�X���L0���7�r�<9�ʑ{\<����K4�7�Ft�~@~�vu�b��n/�$��ޛAh�`J�˿�K��S�H�����$��Ff�[&�H�:�������fL���/���}V�WY�g	��jT��>�|U��*���$h��0q�A����4>���B�(-d�	@b�ML�uV�<��MWe8@0k�@s�!Z�.��7C��j:� _ͽ�aX��b�q,7��BUk)��"U����J�D�{P�
,��wRd��c�G�����Q0��.M%
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�t��y�]њ�/�p�aM���Rիv�S����]���C8Sd\��!��_±���	v<0�7�9:.>�T�s��(H"��q�uK�&��C�f!��C=|�W䩺rH�,�#�wF�p�_���;2C�"c�4Ov�]Aऽ�8)�Pid����P|k�`��ѯQ�y�Ϟj9R�B��́��}�\T|������3��9D��@J��k����I��m���6%��VіR�v�K�����0�oD�����h_�����RCW{fH����E��	نe�r?�2�Y`��ˀ�7���@F�gJ���u	: ���˴�:A�u���hڇn�M�4���)���]��>��u�?��	���	����D�/5��(�1RP��:ʊ��p��2��_�2q��f�j��{��^G?቞R�Np׼���b@���	dZ�ɟO�`1
T��y���>��E6:f-Q������};�Yo�Č����JY��p�x+�&)��޾r6l'2��hkt��-ZΥ�U�M�Z� �`ƌ0�Xڤ���q���v5��,mq�O�k�}g�z��:y+�O�b!m��}]<�ųl��p����DOϡ�=��QA�a��8�\���ѝ�ط���O�i���5�1g|�*�X�D�&��>8�IOge��U��a�*�L��-��3*2vd7��c|����H5y�z��XP?����I��!�k^��s0j뾅�_��G�6��м>Ցp�`��Q�=j��#�oDA2q9��yv$s��۠G�v�0��JZ�ї3������1�,�-�(��k��a��ct��段��=���>��Q�Li8��}E���_!�(����X�i�/� ÓU�W�#l�9�����?�|4#g�ܖȀ�b�����Ffb9u�U�%�-M_,�63�v6�.r�z� �t�l�)��(ZFr�bΌ�Q��J_S�`�v�.h`PY.��f�w~�]��3���-�g�$I3�+��V�:�.<i<�p,1���;�f�@���u�ӣ��2	� S��|�uPյ;o:�!��i^�2qFgRS/�!A���=�)�%/Jg e'�X/�'�]�p�8�S���}1�e0��C��B��B�p��nOf(,75�1���j����6ֺ�H���3&���QV ~�_�С�PM�ݚ2h~x=���r%	~;5����'O���O���P�0�h�_+��/G���7�hӿO�B�P-��#���C�Lr�f��CH�p,q�g?X�	�*��^�����Su_��t'xႻ,�QWlv���߹<������ش���ѹ�s�&�辇���z0�&�+k�o�Ib����1�k
ҝ������`vԞ<�����մFT9B�=�&'�Ԁ�d+��6T%�æD\���e�ॢ�¿�#�Yu�-̇�����������;g��[?E�R�����q�U;i%���n��Ǎ"�\m��p;�{b�\��7"��%
���[��;����!>��0��xC%r.푾9H�K<{V�z�[�P-�� ��ptóc� ���s�6���Y���c�$ܠ�M�E%�k��� 
�%�O�7��~#�ͭ�S�"Q)������*�����04���.��
z�� I��l��2b�B��#�/G;p�*�+�v���	��*m�<+
n�c葅�)_�`�3���7� �u�� {�A��oT�4�����X�����(�ȥǎ���n.�|bb���3��/�C�h*v��#!�y����ˇ�Y�A�I��v�eP�x��f5Zq���)�Z4.y��j�5u���ڒ;B��QE��u�
ʗ����Yv�T�g��]�jn�:N,FU&���@�kh�dv��l�6)��}=I���s4*S~m:Oy>g+AU	��4=x!���[�81��2�R�dc��,�(o��w�x�U����_���X�W@b>)�"ɑ�9�[b�}�ֹ�bE	SOs��:��W�Ot� �� ω�u5�Kｍ��q�f��ڔ	�Ҙ�h��埀&ۃz��'S9�yS��\�p���y�#��C>���-i vr���G���s���ܵ�J%��H0. ;��u�.�O����3c�~]�29�L����	��~���2�Hf*R�Q��|~��!��=���z�)�D)"]�t��w�8�J�1Y;�xĽ�+�N^̹�N�@��	�;TIB``*��u�HX"����A#oPCG��wN�J3�1J��Ӭ[��������ב�t٪��\�	v=0�Z�U4]a���"nj�l_9�r:�n'-��6��o�����b��^ն�]�xnb_>����KV��Î�f7�'���x����OwR�ݴ�3�F��4<h��G��X���קD�VoE诗e������xǄ���\0�>������ϴP�=g.*�ރӤaI�|��|��qXw�R{<\A� 	�����ӾJ�H)��z��Q��פ��P�֬:�h~�shI���Y��K�k�V�=�1�	|݀T��:���j�.k���>/�\�H쇎.f�Rǆ�IA�iY6��
o_c�5��rv4�m�Ӌǆq'-����ޣ����q>t�z}�V�x�`�BO�x&�=.Q���N_�æ���m�GJ���Wչ]���+\г0Jj_2�Ӑ�.a!=$XKz�H��}UN��ѩ��A�zNn��%�l�`G�C`�h��dn���ûAH'&���;�g/�J��]��srΉ=r,F���$���Ѐ~�0��|�w���i�cn��\��P:�KN��*�u�� ��9q8��R��$!����g#�w)
/���N�� ������:�q)�Ί{L#��`����o�!�?[��&�a�,���h��ԙ����J��i��,D��o��H����l ���+�6Y�^��U�;��uԒ��I�h�F���f�׿8!\W;�����S�5|T����P�'�]�Ca�4�3̌�{��*��:�Z_�Z�Fpf �����n�"�y��[J�ۊb����g�klBom����,5�����{D��N���?�ϣT�� wA�Fܩ?���9z��>뾪17�p���@H~�!Lk�2#Z���Vl{B�U��qH�X��;j5�ү9в��I�S7H�퀍���Q���Ktq��� 5��)Р�`�	�tqP���7�i)ĶF;��du,=�l�e�%�P4ϴ7�R���wZ�h|����ņ�g��9��>s�e�:����JtG�Q�=�F��]S��O�׼��~<�k��@��H�^ڢ��l��M~��
V�Ⱥ{���\�_
�1�r_��j�78�Բ;�j)
pmO��9]z�M.X����f �n�s�g`7Ę���|�W��� Mi%�1�M�yg.��D<�d%r`�KnqS��,!oC|�
I��9)f�Ԛ��Y1�,N?����=�/Y�]�t���Z|����}Nr�����H$���"s���u@u9�!����lM� @gi�iD�f� ��_D����ܕy�x�w�����/��<��\	�q>��v�MNr����sd�RX��{�7 Y%fL��刟6)᤯ùz�D��DƔ(�&F����)�#q�+P�Tu��C�����X�<MQ�D�t���%8i63%^+9}��&�&4���x�Z9Q�R��@���Rc?s+�������K��4��x��(�H���x{�5%�<3e��Fc�B��]���`	���X�L#<�I����ĖLA�O�E�U��n0���~�o&�0���*�}'	��-6�;�
]���.X0�]2�7�iE/a2���PY�1����kk̠�FJ�W3���7�^��Ի���뷞��ܘM��pv&��{뱤���2��T\�р~�w�8�u��+"j8�6�/2�|�T����g�
	6�s���H>�������R���YfK����)@nf�/G�z⒠��j����	�p�?f��K�����a/�?1��[c�*�2��,�>(�!.���߂1r17��)<i���{�	��ʌ>/���B9=B��������Q��ey����ն�L�\kd)�#�)��ʷ;;i,}�;�0jU�O?���%6��V��`}5	v�-s6��T4�/�ϒvn�*&�����7�3~���Rw��Y�3F;f��@%��i�F���$�wZ�v��%i��O�.��:����%�3c�m|p5]�;t�����!��a7��[�/�{��=�!�����J�v���2Qqv�f���enVXN>n��UE�!Q����"w���G�ʥB
�>�8T�ņ! ��7ְj���u	a��A���&m���0ea;Ne��0�|���×�4�Eoթ�i~���KwmDߎp���՟�U������7}��.߫�e�τuS��͞BQ0�q'�-D�y1D�M�u ���jɃS!��!��d�{�)��"�����'\y�5�����nO�&5r��/��2���l�lo�o�t��kG��&�Oc��ȼ��~%��^�|�নfdA0�Z���7�ÎK��&��W�-#�,�ϱs<�o�ѥ;�����iK^-'���ᡇMK�`�Osލ������dM� �B0x�Pc��AC�y�
1�ەY;��MòÃ�v��W+�����'� ���U�@��P)���p��:�T/zSp<RVϬ?X&��˕����ZzD��ˀ��(nL�$��Ρ��ܹ��)�f��(C�,������oc�P�7|�9�n~�9�/.�����'Ă��"O�9����!˦��%D�g�c�>�^?d*.�.U��X�exHI��)BcXϚ���C?q-l����m�tL=	��x_ˬ��ƨp�o��
o�ֺ���������4��zTqB0W�g��n,ޑ��3��Gp��6 �'�b���«�t�, ���㤪���]e!���1Q�G�5��lt��Wܠ��9�_�mS�)N��`>xyC9WϘ��8p�Q�ߞ��7�
j����{���ms.�r;������w�ZGu�K�1|�C���"��>P$�4��~#��P�bQ�{ߎ��n�����C$V����:���2$��Z$�U�)l>��V��8m�u`l�|Z˭�~���Lfz���N}��ǹ���pNe���#��Ï�w�f'(Ol؏�,�_��mR�s�z)r7�q�朤H�1|�!ܗ���S�`j�fCDN��n{�j9��i(��~3�'#t�X�}k��{�jQ��ɝ�Ck���ۊ�?I(8������*m�ģ���>�}�:y�H��X/lZ�zf@�~	o�J>^�^�S_@iY�U(.T�h��n�R�,/��&�I�鈤I�I�M���ND/�����ʹR��܏Y�%m��j�N��
���o���,�@[6��NBrƶp,��щ�z�|F�ړ/:� �ˉ?�E{�_�͸��L,a�aDr������ZM��aTRtB���?J8���y��p@�Z؃�eN�R�ั��=��S�ގy���y�L&V�Jf��U��bQ�i��ο�������m�p1Z�@��ciŵ�03Z��7�)�'F�O�rj:n�X�ﭦ��K��7��nǿ�I����wQLy/�e��&��_�`��R��Q�o�:NΑ�@���JR��������߶	��5d�+#`޳��{��o1\*E���X�f�p�=!揬�Hp&�<1�>��N��A�oxH:�\ ���U�>|6\7��kA���9$�cnз+Gk��0��Y���O<>.SB�q{�T���u~�eb܀}u���^�)��wl�����&�*��v�	�k:�C���K�e�٥�W@���h@�w뽌��<U�u=J?pb��Ë��7�	���d�9);`��
Z>}Ƕ�+�3O"[�z��6%S�^�SbL�����4��=�"�
"��X�k6��d_^�a`Y����SG����`�������n�Q<�� z+��.�8��S^#��}G�	���x5�k�k��_���[���9��C��rTŅ@ݐA�4
s3�.��bi0:S!�gLM�$�}�b��o?�v�R�FR�]�h�&�3Ò�Z�������Ӊ̠fq�ߑ�����v\�s'[�T�dV��&��<����BЙqFu�`cW9[$�����1��Ň<<+eY]�,�WA`��AَN�-�)�\̷�m�ƥ4���]b�����0���y�LvӺ�_��H]+x�M����;�H��1��,���gO|���#�h�!�������/=9��2����{H�>E�=\�g ڥ��vG+�>�Yf�]��������"Ge�����^�@�ށ��j�+�#�� :��s�ݓ��<��hH��(���DZ����@��$�����zǹk�P+��\&��r����U�p��S�8�4����EpX����L��.�KB��ܑ�_Au���N�����6��d�z����64�j�)"��%:��Js���;9�ز*^Q�6����&-��,��ks�j�^B4㠸�U�C=)��q6����>/�k���qG���2b�'�n4�=�j����Υr8d����AܬF
��W�S�'�4�4�������п����J�ub�E��Oº?���ٳRa����J������1���7�ڐ�g_yn�i���@�}��IL�i�Y���` ���Qq䴔;:����6��F|�R��(g����ó�W0ePL��6m)�O��L�]u9�����@tךɯ��B�X�%�b��1a��Cw�wGb�v�N+�n~1��`b�,�b�4]4��G�8*B���E��u�Z8���qQ9U;Vl���꿹S�8o�)S�%o�8�&�0=].CG��1�ǁ�ekL�X��{O_��Ha���.1X<���y�7t��6��i�Y�*k$�r��m�AE��L�N�L��$nN��Ci ,��[,]yB�A3Gw�Ǽ�jm~8� �kX�|�
S�w�W%9�d��c*6���;M��G�:B�V�>���+N���5��7���t��q�lJ�Y�dy�#.��7zj����Ȯ+F�&J��[y,��}ͳvSOK��PxaijZɽ@?ګ��;����+�s�Ӵz�v�#�v�͆��:���_��h����P�9�S�j��s�z0|-lNn!��)�eK�%�����;o:dbE��Ԍ�qղ~˺���ǫ��/���ӷٺ��jɾ=����������y4N�Y��t�(w��\�,���4�3�c�������,�˾0��O{ROk.g��%�~L D�i� �@G�i���b�����4Ԥ~�}�x�����b�KR����`�/��`��-^��<-b�IުI<3���6�,������bl\_�p����M܏M�1�δ@mM�J��EDO��7��*{�/nt� �h��mI;#��L�,짭�~�����;!?��@��>�����T�ό��A�6���A�t�7��M�d� Oy��*��N�����e@=���O:���fњ�D�[$͵�cls�˜෢�l�}_Q��J[QM;�@7-�
�އ��� Ғo���+�	tZ���A�~�,��X>�o�T���n}-Ӯ���}�5�h�m�EB�X�&s�f#��|�a�ŉ�6p;G��~��	�%��$��6���S��#��
�a{�}Dfe��ͯ�B)R�V��6!3X;��\�Z�ѠZP�"�HH���=��#}x���{d�6�i+��@���E�#M�T��9��/�˶R7���`��ܭb^[8pkH~�������f�FAգ���+����c�]�)�U�W*Ǟs}h���p���;�l�ɿ+7t �t6M|i3ё-�A��l߼]6k_�Wa�_&�l:�g	���E��<�7~a���Kq�+Fƺ0�}*W���t (�O��"j�����-NGWҘ�b��w4[�"��x� n=Y#�ڊ�4_Ͻ��-ߕ��ɩ���eKs�����[��
��U�N�9e��~�&�W8��;�m1�����2��K��4w��́�N�W.��k,U��D&������� &a�8[lM�\gQVEK���o)=M�p�8��|���	����V������Wo����)<b�� �����mE�㍰���g�%�F�jG>�/�2W��F����|JN�4�[����!a�zL����Ϝz��T�ԙ��C�aS�ۿ�_L�v	R��-��X*��+������L\)-�n?�� �z�,��n�ڋB3� E�@�:O/|�tљ��|P$�,v]_�B��F����x���@<���.��k��+И�N>	(���Y@cvĞ"`G����d��騘�Ъ|���u�A��u�b�NF�j���ī����FB�tɅ��r��p��m���z3�^�(���(��#�Z^ɾ^�)�_�A�X`]�0 ���'�j����>��V�bU�_������N[�fYGJ�A&w"n�q,��gN2�{�r ��#��%�C������^իͣ�%���EX�2cWA�-$S��R��?��W�����Y$���AV�cֻO�TЋ��A��R`^6��+����G��^̯n}9�̮rI��Cb��vY��l�M�Y'C-ւk����͜�gd
Y����;���k��Ii�7�X�O��c��&$�0!��x(d���ٯݴ(����Q�B�na�*�"�ɷ]�<DxA)mw����o8^F~�2]ֶ�u�ֹ��:6���
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`�����T;�x��Zg���)U�b����\C�]ȧ�n�ig���uWg����Gb��i>������o"V�SdsR����r�x�����5�%[x�
�e`J��:������D��%�֯qd�����D}`��н6a�_�	�ͯ�m�B�jpG�zy��b:�1v�cn��H���G�#T���n��-:��L�L�;Ha͆{���{~F���pJNG���&�P�>ҿ7�Hefv��po�ڐ1��R����J�䬝|�-�|���/���'O���l/��Tp�i��7Z��Zx-~�P\`J�{*c]��RȾ����%�T��I����$:y_����_>k��R|�!KXEɁ+��J %��:v���5I��k��뱨{Kv�?���O�g�ii�	ϳtm�5��Ū��=.�Vƕ����o��<ƚ����T3�jL|���� } �� ?�m6m�͚=��RP�l�)Y������~	�a�+]��<�9	S�.Q��kd{8ދ��4xRq{9�]�b1��ȵ��Й�A�'q���������EԦM$���2�ԇ�*�)���
M6���l�/R�����1Ww�%��� ��gn�z�b`�+IR@���%��N왹*҅W����&�%�؀�pv���$�أi�=���L��Ӊ�v-��e{��M��p<�;�?�[���Ql�33��SB0�A��*9���c�O(��`���4}J���<t���b���˴�J��r��U�D��[�[@y�ׅs�y�N%
��p6�����T]���i��3�m�덭��߾$$�_<vZ��/���{r��_�ύ��`q�;�6ϥ�+��߹�g�I�Ҙ
!p���U���꯵�FT�j��!5�Z<[4�+L)�|�
>�� �E)W�i+s���R�`�GIе�� >��LH������Ѩ�����ܣ�Ԓ
�ˎ��|��G�����p� nL�C�>��*[��4�+�\��}Io��2c+�{��MS{X�p�bs�Yg:d���͜@�<Ӫ=Uo�य��*^[����F�v �XmXuʛ�=d�GK�����2jV��L#����P2g)j��������MՓ�?���e��RQtB�����c���T���m�K[lt�÷�}<y�m���Z�Z.d��2��[y>{&rZV����tR��y&:�f��sv+ߝ"��W��Z4��e��tQ�y�L��4��xkC��h`� s��l��� ��X`�%�_�`^��*U��(��2��J6gYwV*�_�	�/�R'.����ͧ�ΰP�W6�\3m.Q,j�u��b���NB��q�n�.lI�9ZKV^�+a�?��Z �pF*��9`!(���ucO7��?�(��^{k;?Bn���'&Gb�SgЄ��X���8C�����?�,����n"m�ڌDi���&"S ȖTĎ=�n�E�Z��!�N�7u��9c,	Zc�̂�������i�Z�)-���6;��Q/<H�!��p^a����Y�0ϥ��O���kHݝ>"Q��7
�!
��4�	5^����_�C��$G��F�920��JH�@a|��A،�x�FX����-xTɽr�*�@p|"l?�
Sgs�Q
��~)�
�~_����Ȳ�IHƬ��Xr{?�����
m�
3M���w�s/<�]��. yV�� j�A �i������T&�t�����(j-j6�jN�Q��XJ�̑-ֳH�?p8K�ϕ^ߢod�+�~�zo��ߐwJ�&~�%�?fF��f��p�=�a����ɟ��b�o0o
���+&�Q?�W�֙�p�w�I�4*Ac���TML�1%�N�tŋ�w����	�b|:clE�̦UwQQ�`t�cR�o#�W���ɤ�ړo���X�;.#��a񦠗Fߧ#���ʪ�r�̺��a��:��S<M��g�qɼ�~��� .M��� +��jaK��D�@����*g	A�ɍ۬]v�*+��\���S�۵��1��ϵv;��&KI䦠D�<7��1�ĝi}t����>!�TN��Ҽ�)��Q~�;��/ yN�mu���x���R�#6���@|W��Z��?;�����x,�	���5V %�GJ��,�-�� ��Aj[�g�H�6�Cn��q�����=��(98n�7Xh�٣
��\��.ۇ���ѵ1�qI�%o<��u~W\��l�U<�h�zK4R��&'�����3�{b�T�9����cb<O�.�8e&�	q�=��T�ttgDJ|�[���w�n�4����1�f��9Q4)Q�-�!�m�DҔM��Ȫ)�{��\���cµ�i��)�m�ĲҹeEU*!\�V�_/'�j1jU�؄OT��
o��,����[�E���E1�
�gs����� ���Cc���ll��S�L�{��6}�9a�FR�B]8
y6�Ί�g`[��Z���\���ߓ6A1��Ֆ=�4d�����d�ƧX�ȓ] �í$����>>�L�'y����RxWy��n��V?�j)��V�-r~��I�`��lC��w���6���mS7Z/�KA�=�P��y)�Sϥ$"v����0��W@puzd�8�`��c����2��1��H�TW�u�C����ʅ�C~ڴ�w�2T�Qn������vƁ�)�FW�$�ͼ��f3�ռ3Zv�RB]����qp�}��oN��QRC;"۰�1U�\��,i�sm��r �r�y�g[T�?����N/2Sc��J�RM�/�j@v+~�8=���8�m8��~w�A����ΐ����yW�(@�Gtp?�Wm�LgX��0��]Z�&���� �k+G:ڃy��DG��,3�M�CK��ƭ�*d�a�������wcaf���:`�bf�͸��s��8sz\*SZh*�q�V� S@�p���8v U3B���6����}�C��v��Dv
�{���jN����^*pneo�7�@Ve�������j�]7�{����H2J���mڃI	��*ׄ�/�O��5�1�1q�������ӽ�]�/���[8H8�����rH:4vq�>7w|�b�Z�%M����=9 ��(Q9��q�eɫ��S).��ֱ����uZ̈�js�g�[*GM�sw�7�7�ig�+J3���s��(��/<�D7i��b�w���I�r�-]||�+|TBO�ۜ�/���,�2gC�B�=�f�1i�����CRV�֡����jԔr���������f��.xq����9�x5���ct`�F�"�^rO�]��v�� �~�L���*/`ֵ��>vS�#�QЅ�4�z���[3,晨�ݑ��NDH�E��g_a�f*��=���æ*%]�Rs��w�mS���1������"�J}��Fyd��9[���}j��\w`O)��/r�Fz�@g����Z���x]$���o	��})Y����A����y��D�l��������ԃ�6@:7B�9x� !{^�b��k��p'�';A���+1����YQ�D�J���E7͌"�=����0�/3K ƭ�4b=N׼����ktR������MV���eʥe�q�&jg�4�_���Q���� p���&CE�+-����(+��)��*`��>%y���O=������s��2@��c&A��S�92�/��΍�^�/�鋸� ��7#0۟uYo������pdN� ����(�f� �گ%&0pP/��=�9��@m9W�k��4z�߫���˗R�U�����\��+���p�l�5�	�!��5;=)NFn��^�o[���C^8,�H���nm=W��L��j��6^l��(¦�U��3#�8d���d�� ���B��p@�(�BR3We�	sp-*���S"�{ɇ��̨�p.���|��&��lXRd)^�(�c�$7 �
�^՝�^Z����G}�l�x�4b-CC߉Ld��3�Z������(���x�<y8Z���]��	5f}�Gf{�%)E��nߒ�`�J���rG�I��)�Ū��Wx����O�¬�bD���d����\:�;�y��T�u\P��Ӵ��ѵgY��-@�F��fd� �^�r��\NQ�x�UR�B���A!Yfx2�0A�-\�;��#W{�o�d�bd���t�8+Ɗ��8ERS-�\ۓ�
_�)>Ha�8#@+��57f�A؝qA�s��c�3$�&a�U�ο�%ƿG
�/G�P����0��F��U� �������Ãu�+�W�E�Wn4�H���}��I��O4�%�K�:~�EhY�0j�Cѓ$�䠦��ħ��"��ֺn n߼��n��[���4��Kd���xe�רUZ���l�[�kPR�5���#��%���AE �i�3�4FV�Lo9wO>���c�d)��Yl��]��11y�F̒�1^
��a1�H�Sk�;�l��"]W>�a)�,g�'����r�A�X:t6��J��N1|9��#
`) ������΢�P-;7`M��8�z���6��Ɖ�9���B��YauA7Nؽ�OY�;��lxz���o�o�l)4�cM�u7<�sGD�mv�0��,rϤ�z*BgD�Z�Ӏ���	n��L	5�H�}�G5�<,���w���U����(2f�a5�N��v�E�s�Y�D��m�S����Ⱥ�k��[�[ڸ5Hv�H�{
 �
᷐j�n�g�O!� �?���X�45�V�Ӕ�v�x�~ʤ��c���W�k��<*h_ש{*ޭc&t��,�nh.m٨�q�V�M�4��1��dk�i��f,�Lֈ�W�M��ؽMe4C�e�nfb{ZxX��1���ɭI�h������6)�yW�ր�ֳ� ;�	l�h���yx�V�)K\P_n��l Y���,�IȒ�E��K��yf�Wͭ��d>������,�5<h��3�!�
4{8��~����,X���t���K��.�O,<:�쐛|�D��L��������2d(�g��8���f�&���q�����*f1K�'a���&=d��Ժ�u^-@�����i�nR���k^[��z�#I6�`�\��&�ɺ�u�9_3��ʛ`����
u�*�F����P��KԺY�Q1�g�nL�4Ъ�MB���
SEl��9h
7ي)�f&��!�Ndf�"?�q}N�[����b�r��O���	 �#/L��|�M��j �,J��NP�2炓�L5����˜&�T�G'}rM���'�y���J�0�{�4�k­��鄣st����PB�f@�E�𜠧{��y�̡їN! �Н]��t�P�gvgPS4����վ���.-����:�K�F�^�}2z͂�%q8*>k��y�zk�����.�mu}/p���y�2�mc�o����������$��!��F_���?�����ݘ-���,_�Y7}7�CE�צ؛�s�.����!�q0߸��|��$�쐲�[9�����S�=�^��]�>F��M�I��>yp̙���'OY�nh����h�.�ᔈ�I�αc�^�����L�JF��B��g�K+iS���y���q�7S~ZY]G�i�z�����Ӱ�d�<HP����v����FX+O(v5ҟ&�4�V��ߧ�;��yAvJ�^D8���)�Mr^�'c$��ojA7i��N�<�b�D|[93�ʱFK���E;-$��S �.ޫ<͐-��}����ZpH��`��R�-'���F����nh1������H�qqy��loȮԃ�Yy��%x�sO����5� �CzN�$"\��$����|��G?)X51B�-~'hO��]^�̌����O�?}ð�ʺ�,���{`;O�lw�M���+#T�ܑ�*u����Y�=t�P �� Nmi�����g��],9�yW�p���'/f�B75�h��ߛ3_���ظr��#͍�G1^�o�w N��H�AgVh�u]�>C8f��6�fc����vS���y��݊���F�&�b_X�V��1�<�}�TH��eS ʉ~�&��3	�m�?'zg���ck� ��k�3�BB��1VL���M���6�'���E��Y�������iAJ&:ͤ�5�ra>-SSz�A�j�L���bz2�������xtL7����Isg�񩰇�6���>�}o�d"�-�����x��R�͛�L��JQ��J>��{���0�(�޿�BE��yX{ێ�'�繽�|��U��zJH���J����4t�|��7ۧ����O�_[��b;���=j1�S1�a�Ym�돼�a�w�ߎ�����JM�+eE��D�&UX������(r��V�e�����^��3!���̘W%�Aa�.��E�bA<n�4����=qx�+�$�\}V��7ݓ��<6���DD��p:z
6���V��ʃ���Ag���0��#�Q@�����|�� ��R�_�o��as����!�P���3�n'S>�-�p�$���S���Co�`ږ��3�~� ̵�$^�z08R	��g���������7ĩ�%�:�]�Q������T�hM��~~`:rӐ��{��HcI̧��CB��+�l�_n��(�]Ȍ��^���xL�/�^7WǗ*�U�$�Y�w�����!P��c��b�٦R����yQ��]'U��d�Y���0P�&ܤT��M~��4�OJ(ʾ_e	�Hv@ͩ`�75����ݚ�vǒ��U��� ���!�M@��9�\��G`�����%
R)w��;���ݔ]�Cinc�"�5��@'���z=<�0��d')�\�f��I�r\۰�.��3lu� ��94�@�=Lz�˲!?9���2ԕ��e>̟>�Ѧ�Q�V��?p��Jg=J�H�L��$S��a�7�3�f�~Y^���(`��
�;�NZ�ں�lߞ�Y�����RKJ�V��2ԯv��M��ߝ�ec��)w<5t��W��d��F�cx&���kP���8*h�%�F�'*Ql��{�_�v�F=k�_�LoA˰r�@4��%2�m 1��>x�I�Ԭ-	;��5�8ÿq�hȢ����,��K�G$Ж*'K_"�$�ޕ�2�dA��V�������/o�rj���g&�4�yC�m��(�Ӻ��S��15�	��ԣ)���݅�|�痫U��~(EnX�fP�$�zn��F�����!��-RS��Z�Q ��B��{|O��rJ�#�M���Pl��g>�F;�h-S�Ƥ�2 ��/3�]��l����
El��W	��C��+J�Wrj1$�ÛI��r��D3�d�ĉ���[-���KI����Ӯ�vf����-���h����-Ui��e}�?n�q�	������)J�v��/3{��L�L�Մ\�Ò�Y/\6%6q�[~Ϡ�`ߏuV����O8#l����<�6�&��]D�a�SO'L;??	�MB��L�~�Zk���Z��s�Qn𙮽�ku׈6���?��fQђEKp
$S�CDT	B�Cs�|����مE ��P�Ⅰ7�9�09�_X"_��\u|E��R>@һo! [��GuΙa���^��������q�������BW�9�?[����Pu	�����V���
խ������7:�~O�&��{��a�n"�S�ѻ8���)���X�ˌjD""����8���5.Mu�&@�p�P����i�v���ג+��8�>SD-7d�1QA�\M��l�R�Hq�A�o�/��	��j`^9/(�~.T,�?WY E�����j�� %j4:�¯��X�60"�1��~v��rIH����D�E�g5�]do������Bґ����_�fl��`$0HMI�&�QZ��2�c�⏑��ЗB���CR�ވ!��O.�WȢ?G����u�T:@��f��w��/�!�ЌE.jf�2(@#n5pɟ~���kr1���Cv�Еl玩�.�9bE�h)`����B�F#M�c�f42m��i�=T�(�ī{��Y)S�^"�Ob9Ĥ��Y��/U��U���oC�{G�R
A
�1N�s�e���\I�Z -V�\�$�e���B���~��i��OМ/9����@#;H�3�#&��9H�u0ɜ�~5*WOF���:&8�}��C��Z���G�����#���7�$¯��(��};!��ҤYM8��x\����CSz�W�Zı�Eq���P�!O��L��U[�S����t������3�#�T?��!�
(����c�c�Yw� �PP�=e�l��ݿ�v��������r/jA���~�"�`=��
���@w�Őm����9������*�*��tfRՉ}u��r����:Y$Π�KDK�O����;�G>&�����D��������Tck6�Xiv/]Ƶ����"��i�{q�P��,o3�!_��$�Q��c�T'��5�$�l�cz�9Yب�6�6����F� B���1��xq��C������I��Z_PKL�2�`)V����P�I��K����&F9�f*	}�!�,F�������z9�5e&�2S!�S��!O-��҄�O���@��AY�&Wʦ�5��
��]�]��m��*R�Ռky¢�u���H�	lj�-� � ⦂Т�W�r��l�8{�&}�:qx�Ay�Ka#ВvQ�+3"�'#V>�!�^��6M�9y���L���b��"h�Gףu�`Ҵ-��/��o �8N��U�RzT�o>5C��,���Y|�ͺ${<��,���&f���\$DG~</8�r�7#�G����NT!bX�ëPd$K�l>�K���:���g��vM#s4|7�K��Y~fsdYV\��Q&_@�](Q��������!�+"1@�]%� r�gWa���I�2��{(rI3����M���(c����(�")�]���"�h��\m����� ��B���F9[�v9j-���
�C�Z�--LV�(0(P��.�H����!�At-�"�Td(ӲЈ@)�K=w�	̝[����]�F�b���Gg-���g� G��@��#S
��4�Y��r~�l6~D����@q4z�^����ŉ��H!/�7�S0�UT������n�:@4�p��yx�=���O5^�X����vG�6'���W�QS+�D0i"e唋__��³�P������#���Gک��W�ڎ�\n��=��A!���hCQ��Y�uk5�E�#f �/F�o,�#a�dh�y��RfϽ�m zZ[@t=b�=�z��S��3>�T�iG�-a#7�PWA�..�n���*s�NO�I;�3M��^��@��2iS���@��֋RY3�����J]@�A_M���� ?�p�7��̫�{b}>��3h��f�n t��ؗ���(j��츏8�t�"@���r������)��;��.&YÛ�0�^���dd �mXb'T��?��n�ɒh�+>2sXH�o}�)�KX�ê
D� �&F�Na���t�.Y��~Ҫ��K������6Vo�Z!���pd]��=�d�НO�ZQ��8x�U����Ø8���N=c|�&�U�\����]�-*��`�O�:Z�r�{VZ�..#�o0�ӽ̀5m�l2τ�?�]VN2�
�#��N%߉���GI@�����p����Cxy���ɞ��o8�������;Ժ����6�x�b�WdSa&�	U�'Չ����3����T�m�un:��7�5��O��񬹩�I&aG�8c�B��G��`[���S����"?~!��i9����.'����M�p֔���4� .�!qQ�#��oo��\��1�]}�,ܷ��Dh��~4L�.�E�.U�B�t���2�W�j{3r�s����NȧI�P�w6`̤�:��k]��qV��Te6�����.D[@���r��Q���=���p0���V353���'��\ʗ��l~�� 8]����^PU1"�Ow���D�[M�a�Y�T�y��%_3�Jj�&��)"�T���(÷N⃚2ݬ�o<�"�VX�S�֩rڧ�x��*��,���[���`�J��o��^��hĒ���UBS&-��c
�0ZU�a�,@����_eKr��\7����
�����3��B��8M��l��k:D�L��֟ȲQ�\��I�`�S��k���r4��|��
! ��rY�̂�F���<��o�EX���#߈L��e�w�.�LG���1��i�AO'"g�.�	-po�4E����x��̩0#�#��18D 3FĠ���K��s�!�?�g�Hr�D��)~#��ܯU�H���ی���o��o�$�O���r����U\;P��.rY�S4��!ؑ)�ൕ�m���A�;Z��$]N���I���J;��>i�����R����m����##$�S�?��\�R�������U��@�M��I��BQc�!kehb�	���5�n��.�R-	�Mђ�H�ޏ��0L���Ux��v�2�v��h��=R���ܿ$0:��NR���"�ɴ��Na�d�Y�
�'�# f�Bnr�"� ��$��߈"^U9Nz(yHl�
�k�{J�E��K��4��A�G�cq�KK�ȶѸ�a�`  ���#��}z�mR �P�N�#��oT�B�dk� 9��)P�"�o�3M<����]3������Ae5X�+�$<�;�-њ���@�ڐ�yy��#�N������h|�m���4���W�3u8�O�����I� %x��թ�N�4��|A��RNn�b�a�~����)�s�;�;D��Y��&�>$��㱒��&�
VX������(M;-z?�`v3��e��kQM�v�Ihk�f���%~�yn��}�QK�bp$���䗳8h+�R,��5&`4O;U�U�q��6���׍r�����r�N[�'�[���E#n��j;��W�p��6q�j\�=Gt�q���>N��23�E����J	�[���+��O8��:*vt"�I}�:�|��iU�qmlh�@p�kc=��m����N��vؑ}c�x�^��8�Ee�Y!� zF��-����4_DK{�J-ލ�~�X���V@l���D����,���"Hn��u���&h���c޲+��]7m�2��xl��=�S|T���**�^a��*#��C�/�-�H��`.�lI��	2�z�M�[��p>�Vܝk�������>�hs��k��*-�l��I�K:%/�Yg�6��A�����A[�~��j���0���8�wC1�1;�\ ~f�N�WMnj�x;�aIc�E��DN��J�$G�9�ܐ�߃:y'�w�D� �L��t��`NK�}�5������.�*�iӇ�i��Lp��hF��KP
c9TeF)FÜ/m֭�.`=Ծ����,�}B����3;�,p�W��J8gß2�H
wO@PG�<I��@R6��մE�6q��[	��e�SV�ڦ�����0� ��P\��[�5uη�(�����vտu�iJP
���!_�pϺq�}��M�ՈY�[���8OS��[u�Դ`�Ξ��ڷP��:-�2XvA:���y-�P�5��F�$����[�p]8~4����B�d��]�N2L']����pj����z�K�#ebҋ�����[��ml��x�9�8�>�R�v��/��y�ӂ��Y�Ą�X�b <S^�/z�����"�p�*贒EY��ԏjI�����k�Eo�B[�Z��P���.7��|�|�~�����c����Mg����Hw1��j{Zw!�^%<��$�`V7����RgXe}/R�`��Q��b���4}��A
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��F��g��b��O�|���O��9v��ɇ���)%v�3J��z֭F���/U��T�G_{Ԑ�
x�,�x��ԫg4�(x�³�S3��J's�h{�l ���^�Ս�2����F�&n��|};ό�r���١ا�5]��ve#lx�0��A���w~�S�FUU{�^F�I���¨��q�>�Y�0���މ�H1nP���rL�hBL��V�������l��1]��a
�B��Ħ+$E7��{eIW�����t8����x�����X�>�i�	Ƅ����~���~��Bj(h���_��K{!��^\~�1�Ud� 9�O���m�py��G��a��&-3�\ch=� q-��T��)�ɽ�\�3��D���_���'O�wvC?t��Y��E�f��B&�����o0X��q6r�1yPM���=h �z��-q���.qU�T[��
�e��i+�F�Ӈ��4��`��ݲ���A��d{�ҭ�f�T�� ��U��n�)f�rDw7+q[���='ܜV�l��,gi����&�����E�JP`�@�vN(����9&�Xya(�]2���%ч��z�a���B���v.�:�@W�j����zVɌ���Yӗ_��V��U ��������8^&H�/dC�AZ�ȼ��	��Yv �.v¿T�s�
���44�	�=kL����1���ؙW���*l�hL���� ��'�����K[��
��"Ɓ�FTw�Z&�)�8�ȅ�� Trj� �GD�� a�����|���M��߆5ǥ�z���
; �[�B���h-���iC���Qcp��+��#a��.V���c�D���0��>Ҿ|W( m���dH[���䈷pM��K9#�&��\�2r�Km��J/��v�,���K�S��v\�Ap���9�@aqVm܅B�Ȕ� %���S�a)�lNc��ȼn��9o<n�V�����ڧ�}��W.!�)$�jN�(>$��!&��Z�y�.�������lB�^�*�v�S2%�r�]Y�Էacf�$B':�Ft���hl��ȂA���F�D�kD��7�ģ��9�ɏp���&ZމH�X9C�MҜZ4��D�i_u��}@���� ���3��N�V�EL��2 �T�;�>ڃ�H��~��V
}]�"�ذ�Bp�+A;�k�t��ppV�tiތB����2x��{5�`������w��&��P��0e����F�+A��4�I�-՚V�]W�����ǎΩ��(DD�x�J�HTmݿ., 9��H�9 �g�A�ك0�������̘V��py�h��lS-]e�3U���q�M��c#P�������X�� #�ƭ�J�>�ܖ�o�����'�u�?$q@d)lr���{GJl{k�y*Xg�"��qN�և�'`����G��X���9Cg�:qT�.�x����T[W-�ݩ|���S�7ā���1��`�|����dq�
���>iNd-���N��v��:��a�w�Z<����Mg*G��5���?�'	�O3�����H�х�ekio�*x�匍��D_a,1�sV�ٵ�����VM����U�o.l�(C������5N��1����Uxj��;���tm'��4?��[=�k�,p��a��
�h���u���	i�o	�cI����fL�XLIZ�֢�A����M��0>�� �C�c�Nɚ���\���%A �c*hm��ʐ'oa�����c*w�K�?i���/�����	�뭱�q�a������|�g��b

}7�9�r�؊j/�;�|��Jۺ��&χ��_��v�My�vCt���TՆM�@��;S͏f�ʊs�U�^$Q1؋K[x��3`����]|�z��|'h�^�U��
qbk>e�_4[�W���Zx!A3��a�� �4ݎd�x7���%�p���*
8�����<�m4���*�����H�V�����-*�:���� �#;���-@bi�D8՚��'n�ey5��(�����UQ���i)�Zdy��Šؕ8ߛ�4؇V�V��h�"��!n޶��#�Z-��:���җمE��[j���@��u�7�Ly���۞�o�*zx��<��赁1��i�s���L��k�]�B$7������Uls ���H�L���^ $�����.ٞ -~��Ƕ�����_=9̐Z֠	�˪JmI5;�W�7��
�
�O��|Cq�׿oZֶ�a��	������}��&��eɍ	9L���6��w����'�$��{/��l�ˮ��/���n���14JZܦ��oeit�����E^��-�;��Zƕm�!6}0�aY��қA�KY�8E攉�����<ҁ�o.c�g�ʀ��l* �Cp(�u�Nh�)�<�U�e�-�!D�B�!I�<+�0�IBݶU"�����6w�ତp~`���v��8;�Wե���{�"�)潵b�y᷸d���g���YB���*?}�x���0� �WB���=�]�����X��L~���s�uk�k΋�Ts�l]�@�aCB���4����b��[g��/RbkB��Jk{-�:+M���@,��8�3�ahsz��`5�[��zV��lRpvg��Q,�i)�)p�a��E�sR^�HH����P�J�xL�l�z7Y��?�/�z�ZR$ޠ5��3��t�d���j��#�.h]j%����	bYȟ`�BX�Ahb1��rچ���6(	$���6L����o$��\̪h��I%�Ǹ'��.$a�?P�F��-��H��&�+�U>Ґl���y?K�p���v����OACIK�ō �T�@��p�U�Ea5 ���UK�B�{>!�w`���\<��&7W�@o�E�`�7��ZX�l&���5*�<ыF���Pv3q�jo�j��d`|DKU���gxbҮx��z�?_~o�[!>K�ޭ S1ǹb�1��u?Ύ���,���R��e�y��[��^��KV��,E�8g��㿙;1��Ҵ�}ؑ��_%�1Y���S�zݸ�T��1�՗�j&_z���`.�.��Pv��_Q]O� ?I!ﰅތ�@�$�|D�h'P3"]�U<W��hBWz8a�>�.=j�U?�|Y��=�V2��ۂ�;l�r	H5��=��Tk�Կ�R{��><�KwlZ� hyk�>a�1�Ev���ހ�.��f�lWە;ݓ�1�5/l�g���j�����ޢ�����?�?IM92��Bqg��撸Q�a�A��eg����p���`�a��`���k�@�����Z%� �1~���v�{�8#O�����f�-F��W�c�V�n���F�.�z�5������5���I�hؔ��y=�T�~+���/���L䌄2÷�J[.���3촼?�ώPn����m�?�d��^I���k��M��Ԏ�Plط/�{�	jۆ��=�?Đ���#��>ǈ���"��{����{��T��7��
�l��ps���l�0!t*��]�ٹm}?��@;�iBo�̒��n��p�F���q����2��ψ�9:�U�X��`��:z�DO���l�͡��a���$pg�^e�n*w�����US�< E�2�m�s筟�Y�)�7{�^��4&�$��:��D��Y������.ʗfw��Ƈ;�'�nA@���MG�y�X�z�{�T�+�Q��^3B�<��b�_9����#���\�;er@��ڷ��u�����%�?1���~�/�� �":�I�Յ����?6	XFST�	��F�rM��>I����s��;I�;��ۻT�4���O��9x�^���@;��k	�CEQಹf��B7-��F`��ݲ���wRߌ[2[B��~P^}AV�D��0A)��1�O
�����Ҫ�J������3C�`��6;\:�%��|4��G� ��e��L}��mRNB1
[6Y s��z��X帷~�1b$a����F�l;�7�B@	^. M��l�\�D�"�#?J@2����Q�ɘ�Y���E�<�[��ttڂ�g���ƌ�6(s�}f�i#O�t.]l� �>�t�v��/T���D)+��W&�ĞZ�7u��%?���Æ���HGR8��X��^O6"��rϜ�>�m6���^�xPeδ��!2$ǚy�c� +��AF��VT=���q�����J���*�?�� �-�|^O7��"�Q���z���2���S\l%~v�$[Wi!ɫGu�w��P�*�h��_�} {�V��
�G���W��.(�d%�՚�hR~�c�P�!���H9ӗN���Xi1e�p4S�CXW��!���~d�\�w���	0���I<�#!l�0�	��X臱E���+!��,A�i"�U)W#Q��5a]��ݙ"�˟����ġ����&|^��YE�D�VGI��'�ܭ��k���b�	�]1W(��m�u-x��)Sr�[5q�[�|�TyO�O�3��;�M?���E 3b��.�������h���6�mnf���w�z��@r?G�fm�4��%��<��o�D��F�.���[���"�t�ȟѡ��CX��r?�z�u�&[ЍEv=29�����L�E�w�(#����B�,�Lbl��]�n��?g$�H���r���@Lq�K��(ц��x���z�>�T�'�H��Y& ppIz;|�v����,��%��dAe�]�����oK�f\����<4�X�y����$���@'�(�,���v��ҳ�ּ.����>? ���$7#z������(���{���n��l/'o����	���c��,�Z�ym3/�=��fP{>�%-{�Zu���n��UюB���w�!�P3�������e�Ex�d�ܔAopxM|7p.&I�WzC������]ȫ8��~)whԩݙi��蟃������Sb}kԄ(}�~;tSt��h�z��b��㕸a�b�D�"��,]���
�=L��$��/��S��?*&���g$��#�|�
-�&��/�3?��eZ��!���N�H1������+��ߗ1�LH���̍d�\��#������"c"�RZÄڠ٧C-1KL��,�U���
(s��e�"? �,����O��(P��ڂJ�7�{�u�W�����ɭ,�ӻ�n���F�Ց�^��v�!�7𾻄H�Y���
w��*>+��rL�lGQ�)m�;�g��_�e	�gi:�Q*�=5J�-���M����#o|bY��d�]d�v�{l�/8Bk��.K��L�Q��χ'�p1ȓ��i�ץT�+;�]��4:pf�}��8�Y��;AU,����)f�~�X{[#@�v�nYAu��9�a�k�3�2�>���u�n�1#2�aݔ�4�a���O�9�=;@�h���NK+jCv._;P-9�*�>��u9�Mhdf{o�@��o����/cB
��e)°N��H�"�N�(a��SK�Yt$< �:��-��J�Q0�6I������BRz���ꀋ��W!	di�x�S�
�B5#Ȟ�q���ׯ?�o�'������H�m~T<�ҭ-Ӛ�̗�w�3�9�b�f�氉�t�˛�ʧlf��EV$#�UXf�.>�"xU ����r}^�d ���U�Q0�J�:
2X�R��OS;�q,h�yzը��]���8=Ҁ#7�U���<�8fs��Ə�f���5�y��E���"�b�Wۤs!�/�p�Ô���h� ��[P�����h��� Cf����	ϴ�Q����"���_�K�D�w)1����d&�.}���}-�P�d��3�q����B��#�K��Q��Y�H���F�"��_��Wu��� ^���e\��w�B-�d��� ��������҃�#.����[�w�f|_�"�*Z5�x-�``��8_�ǫ�톭�W���e��lo�h�ri�{?0tp���RB�M�5F��!�s��*�-�1l='NP����C��c���>a'��=ִ s�I�G�e�R��h�S�R[��n�Et�N��'<���U��S�6C�y٨���*mEq�ע�7�SY<��i@9���ǖ=1��v(C�GM�e��ՠ;aW,�(�3{[�ź�A���Bh���G?�5c8�=Hz9ެ����w�Q��.`u�Hwd&��Ô*�U�F��W�ꥫ:z�kgm�$����!*���ٓ��E��Ji�l4f�x���dd�l���΃���d�I�ƙ�ӊ*�I���u�i��$<�)�F��Ä�E�)d}��]���@�����`�����`��Im &օ�� ��r����!Ix���~)[�o�E1IN�v��8��*�_�|G]�T�ٹ�U���qVib�c�Y�B��K:�y�aǨ�n#�'��([�x6s��8���[��{�)2
�HS@^@Pa���ki%9���&#V.-k���) ,�0�HJ��dڿ�;F\Z<�+�@v��Nʅt�cO��>��M:�o3�oS��IQ�̤��R�T{�Ǥ��!v��)���٦�'1z��Z���@�Zo,���J�����h����)���_t�\3�xء��=*x�eF`F�9��qAn����o��$����o��Z�wmw�"�b{��$�%T��S����S�X��g��E��T�v_@qɉf)�B�TI���র�כ��D���R�X q�(q��g���k@��>�Sժ���Zc���Xf>��]���_H�Mh?��R�9��0F�]T�i�~)o}�mN��N]q���6�
f��Hq@��/������9�>h/X!���HN\�nd;� p�T�h�`G�"��
�xU�8�U��Hr:�׬�џ�l�ίJ>Q�t���Ԟ�M�[���M�Lb-�I�O�������$g�V���`�j/v���3:��tM��R�D��N��E(A}?������%�R�/��dt��{n�S�l�N�2)��H���e�cq����A	�W�
�O0�#�3m�{L����T���bqt�a3�C�.�~���5�}��LMN���#v��T�r��/��Y����,;9&;���2^L�c�Q1(��q��'nM����!{��;#<f��!_���F���E�d�]�KJ���Ҁ��%��3{��$җ"�J�d`��3	a��;qA�v?�3 ��^
2�t��@�.~�883���S�K~�2yt�$�_���o�������2z�F�1V#��h}j��ǳ���0>#�)n�z�pE�w)� ���MMl�eY� *��ϰ5|���%�i\V��s'|���g�o,/;�����,�$	Շ.�i��c�9���VjP�a��/�O�Wk�?��P���Pt]ޑؘf1A������KH�l��Lj��H<��q�d�8{Tڧ�LCg=kh+�i�q��-��*�s��zlob�^��C�7�����?I!��p������{�N�����+���8������0;����U�2�U����P�"
�k�c�y��?��]�/�5Wo���7��do1�DByБ��l\>���w�z+�JEv�l�	�'+}栏�9�R*���'D6<i��˹@���3܎��=��&����\�[E��m&S����u��H�z9HF�J�ׁ���Ms�"6iT�G�*���J�Ji*O���k˙g�/MC�bZ���U��n��A#�X�z���x�׺��U�����.�"6=�8٣nctBf��T`'���~�kuLF�]o'l�����������L��l����@��1W(.�.�>�2%
�AX��w�\��f�'�D������[�f�����݉a��%`�8�����+��w`sYT{<�� n$�д�N̬�X��U�b)u���Jl8�~}��iK�'V`��%���B���	J��Jb�!��"_�*���l�U�Z���0�#�m��e�Lp��\�������cp�eI��-�{��o��{��oh��S[���>��,Yi/#���5����9���'�[VP�I:�𲕹 A}�+���	��U�
�4��Q�0O AΕZ�H����R��PL-k�E�l��
Q>B��*�Z\�{�<D�<&�@��E��"5��($<��7�����X3g(����x��#�����p!��kW-<p��O�ȮM��F��Z��FȀ�6[�W�~w�j�Z&�w�I�j�g����م�Yg�#Ml�ft�A}�X�H;�7`^��箕�#�2��=���	�/kx�	���Y���s�1~I)��eV�02u�o����&�]g�Z}t�X�^\޼&����	>�&���:A�Z�1���헨U�{��ɛ�����������!=;j�/�],����O�!�?�0����HO��@q υ�|6aЈT��u����(�+�;��AI�]���,k��h�:Y8�������=��s)Z;��ubq'o�s+t�����bl���K�Eii�i�Uغ��@y�턞��51�-ט�������E� �șu�;u����p<��*�y����ZW�4����sT��1�5���@Bj-��#n<!<��!i-��5����`��~�W�\�;�c( Ӗ���)��h��a´mK�o�6+�Z �#Dh�B �@2�mVRw(-,��c|M��b�`泭
�M�30\��~�����[����D��<�7ұ>
H�"(��S�i�]�Wk�w����8��V��E74�-sW;>D!�b�^ho|��@��?�I+Zm�f�^z�uթ�Xܾ�L�,5Wq��c���^��jC�t����d�f͆a������k����;��ݻ���kX��Z���0g=��GR�vI�v.��-��@h8���yR�+4X��]���޶��Qonc��r�7ҳ�	_w,���3J���t�0��!��p���$��]
��wQm�KV�P�!�W��[~'�fU���J�#��|��]��D-Ŗ�W��qҥ�r[|i��.�~0�3.�u�LB;�T��/𰰳�S /:�/N�v9���U@�Y��y ����e
պ��H��o�݆G� [��:"j�9�k"���K���LV�q��Cw6 �!�*U�6��e�⛮��<�}"ԁ�3^�gB��\f �Fo��Wg$n+���ư$F���8�Ⲭ�A��7���r��{�{�~�- gz���ӏ�m/�/?lQ.9��zo�%�m
�+�0��^؋�T�=Ƃ'`��%"��I�ʬ[:�^⎓���_���$N����y�b���aE]	�Y�r��\��W���M���dS�\Ņ#��yZ;��ґ1�㠳s�̈��bA�^$Чؼ��;�����(�k���_�'�ַ�jI�ETD4�%��\#��̏�g�w�)
P�yi��!�6���p��t %@$��5m_�a祖PM��}��R�u�d�3I�S/w�|B���q���Nv�D oT������9�}�5 ����:��uJ�Q��4���>�R�}�V_� �*�z���T��%0���WУ�ngs�v+{I�d�MX�ʻ�ˎ�`�:/:�!���cf�&�4��v���S�Ě�v �*L��^��qvJ���M���J���/�i�,8�C�HݶK���~w�zg�ܮ5���hٌ��c�;��~���j�BI�G[������*�I��Fl9�����1��=�8��� �:�&]�����L�0��5B;��@,���g=��ͨ2�L_xf�
k���X��s�S��_�m���Pchc���ϟ��R`J�[���wj h�gq�kP-��ؿ6F�!9}"�>k��tbM^���ܤ?t���\S��驅�Ԯ�Q��[6��� �>��Wr4����}H�(��6"(B�#�q���պ�3��p���=r�E�tO,��u�(��O�EJ����f�v�B��H��?��<�=w��q�R5��m�|G/LDP�*y�{좹^����J�#����:�*j �v/v����A	��:���ky�d�<�Js]�|]7gJ��]��r&������k���y��(�:|^� �V��B�M�L=� t���v,1D�m;�◹����-�ۉ�@��-������H3�<����~�A��Oȝ2�:�#�Z}\����[c_R$Bo�<�0I�a�?2�#R�ߋ=$qJA�sP�O�O��n�$�i��f��g#�_*�gj��95�rK&5x���g�$�=�� ����+�v�B�x]��w
B*@]󺀋�hgQ~�7.��܎!."a�sF桽c�ad}+Qw��<B'-On2�ӥ柈�!�4�v����uNby�J34ӡ""�Q��g���.�eec��$u�F��g�F�T�t��Ћ�)��'����V�E��E���a�UM���s�r�ǳ�E
��A/��ј����Fo�r����K��5���;�K{����5U��+-���p{��{~'�ȪY$��w�G��+<��^�<�x�W�v�Pw
���lĊ3�M��k��z�R�C��)��y�E� 4�9Ӗ-�����o��<�.���*������+�����q�=@[���B��9O�cr���""92	qU*̯ EB�^��dʠ�"�m�)��ݍ����Cj��<(xy�o�:S�+�xf�V]]3�)��������6N��!;?�M������y\�k*�2Ų�1���B��Q�Z��[�QiQ�j�C�_�(�4#��[����a �Hא^E��ԋ��6sȤ3��l��IX�z#���'����;�u��nR;�׍ҶD�;�y�a�vD����Gߢ|�n��y�*	T�p\Kgj�a��-��{��E�S3�!_n�/� ���'��JG4�qM�K�r+�<H��W���;G�89���$4R_�ڈ��d;:��m���u�]B���G(�u4+�?����x�%�����z�
�t���,�YB8��f�������s�m��	�jA--p�����6撻7k�ׇ/���� yb�̤�&��#'ZlU|[R�i�IX���7�����Bf�'�t}\������%���� sA-}���U���d#��1�X���.[�"Ca�TV��4t$����Q��'�zy�zӥ&�A��m��e�r��1
�]�ѢN��]�R7��Ѕ�Og������7a��[�a�οZ�:�⠉��n���<��ۜ|oh�em�5�j�{��K�`3;1-�������V<VJ�� ����1/��K�{X�<D3�DA����[l��C�&X���3�J�g ��{u"��*��k�ǒ+�h���Aä52��*{_{����t��R������-JP�o�&lCOt��Jy�a]�G]7�8����S��m9���'���}���\�)���H��0��mcӾi3d��S�t1�NO�X�I�� �Z�������z)nd!��s��s��
z���ԫ��{C�;̛L6�D���[XIR����Z�	�<�����~NBO�'�Rr�a3�(�����g�6<�$��3�J�s61`����V�>��P��i5+Y�.���ÅeJ%I�r��*�����&
0?���� �n�D�q�[��2�v��6Pw�k�f,�o�g����]�t*����v�_�z�)��&�R��&̘��q�E;���x?7�'�-��d Us�(�#֦�n��J~x�t��@'0�F�F_�Vhyr7��K��m�6���M�"�;���Ţo*&@ҢT��������Q񗺴K4t���1�/t�Z��C+V��_l�?�Z��2_����3�u�F�7�ijE���ƺSֿ�tJ���Xd�7���a�kz�ɻ�2܇*n����G�Q'L�
�����b��z�Y�L�����h�UP
d�A��o�V?QN	�՗�ʡV0��P7���L�j78*3b�pԺGU�y����xP�LA����;����q�s�ϙ2�	����b��@�>�;G�i��%�@��N�ʁV3bi���혇��*-��`�ґ?�"� �g���T��)��@�7o��C�/-��K�Q�=���h��:��DͅB����w�2뎬�������;��W��pS��H\��"y��=?����0��|a���܌�#�ԉ�������F�����ՙkn��FU<"W,���}�R�o뇣�A/?-5������!iڪޭ����M�J/t�kEq��*D�i������)5�T�1U���NY���?u�,��T�u�g�؎���F��"�ذE�[�Q��/�Gn�+9�D����I�l�@�/q�F�v�>%� �il��2�\֯��NH2S�']��j�]����N��pZl�
�ePF������u����H(zh�����-b> ���
�;��9]
�lA.��0��J���ogO��m\.S�DS������X?+~`��t��4��4`�ea�Ӝw����<_c��+l�hM&W$�2���J�y=MK����SyJO��>��Ȥ���=z�_��go�:�����0l�U�ܸf�%�F�Ey�O\�ǫ�N�d"�fB��!a�4��kx����FH��ŵ��b��h�Ȋ�R�?�~t��� .K���6reIT}rT��͞�ӿ����w��G�+t&�ɧ�_��1��|��@����A\������=�(��P�c
�?mp>��hvx�8�e�s����J��ɝ�\3�������w�	�y|X�/Lf��^���O؆C�O-@sm�v9����9H��bI��B<�w���z�,�^�8%�WCCGݷ��J�Z6!�#m�Nk��Q4��|E�CY3�����@<���kn�<(<��Zw�F�	�yH�Zga⭰GGݤ�m��c� ��8Mj�e�m�;#��C/�bht�����Ūw^�I�ʲϹȨ����1�U��,���ⶅ�l�A���~o���	�cC�D��7�v+�O]�`u�0�"�Lp��X���c�Me��r�\���WK���`����uS��!}j��L3�B|~_�S�mp�����b(t۲�ܕ ����sQ�֪��Q9��N��	��'4Ӓ�P0D{�^g�z��&zO�I�hyp,���m��:�.v$0UMNȜ��8d�SRF,~G�݈*� �����D��ohRE�GS�ţ���Y�b(B�řo��<˪=�Q������x����B[�}�m_>��G��EP��A®�ދ����F3'��Ǽ��N\�F�Y��c z��T�������F�.R���f�	�8Fw/�e���eI['�E�
¥�LF����G�*�S$�Foܧ�:�E�"M#ݸE0`Y����TO+AL�Y�P}��ym:8�b_ �ڇ�F"@�yƌ�h�;`���͵ح���(�S)E/���h=3����~%�&�8��ug��ů�y]F �ჳ�ZV�-j����4�θe��	_`l��$qbo,��:p
�]k���B�<W�bŒ����0���@Y$�a��ku�M$��︼�0H���n�Z���چ�OW[���[z���]WRG�����5bc�����[��Ui�G�s�9����ݯ\�:o�B�K@7Bs(1�+� ���BM���U�Gh�`·�z���:����m;Y!�'��ȝ|��؅p�d/����}�1+�N>��� ��8+�����d�\`����ߊ��p ڔ:�x)�/����������kH�;������2"%;���l=�	l��K��R%���sQ��0N�uݮ�)K�/���&��Nj����k�`�L����9M��y�ּg���7�ͨ�)��v�QD�:V2��b,�0���٧��-�ܧ��k*I�0���@���Q�X����/�ݐiR(���K�q:���3�"�;�I�ϲ.�Bf8MI�ih@*�]�ǋ��ɔ�/ ��m����hs��k����Uhwީ:�4
j�5�*J�!ͤ�|���63��d�䧮T��@�ޛ̬��Q<Y�Y3}{�
1z�[n����8�_ ü� ��#�r�s�P��k�ı���v�3*:q1a���]�8&A^Y���"�~�}�6�M��k,�,�p�'0�&�yWt��m��>�T�p�/�hŸ�z(��*��V4�U���]n��S���6���u�;csMа�6H|��ӘB	���IX]0��o�W����I�]ǟ���4�a��^;	B_�q���X�a���J�'���O�� ��q�a�<m�^2���N���D�<��+��"�A��r�ܒ뇥�@��c�ZG�K��ѓ�u�w�Tbm 	�*��Q���ҎSΚ<�>� �m ���f�7��n���ƹ��)��־q�ٳ��Q1n��9�\�Ooz\a��R3F���\s7�,ɧ=û�}��z� Ʃk�	^����s�^ʯ\�Y���~�۵�K^��-��˯�G֚��h� ���V���ݭ�/+T��v��|�.;�f[�{��K�$�p[�?�]� ���V�~�uұ�ѐ����r�Rg � ӻߧ-��~�A��<�(��q:�]ɰ�ؐ(I �Yj#8�������U��������ge��z�����ӌd.5֕���(S(d�q������/Q|&V�)�����{K�[�A�CBUV8�k߀\�f���&��Si��3ޠ¾9G�o4Ѽ��oC����$�f������N3j���쿗'��^�U��t�V;�i��>:��5bY,��Hz�X�G�������,����4r���陡i�y��.Bj����:���9B��Mc���@�������?
E�i�[�6KOٶZdt��~oz>:���"��;B�p��O�)�T8�:b�Bg�d�IL�x�m���VX58z\}����b�6w����M���.���*j��E��M�9(M�x���7:���~��ԩ#�r�@=ӯ���ֆ�ƌpd�g���G�R�H�͇ȣ�[^�C���n�
����¼LN�ۇ,*2��n��vޮ������`O��؍��u�A5r�H��vG��*pP�aK�ƹ�Zrxy2��A�Z熈��Mt`!x$���W��R���`�=���;q�#��w��|`-��y���D,�Q�o�/^vw�����0������f)�~LRY�l���<��s�tb��,���X�?�:���ҟ۞�`�$��3�9�'�G�lX�DN�l�6Rn�fe�C��U硏1�A��'�I�CA�.��H���ل�P�9���o�{��I��>A�^_�a��\�V�b�Gd�xK��>HG�#C~�N���*�[ٓ�3�m��S��'T��H	�DaEm����=wh媄��`�r�N)��Z�c�c����!86K��e�i��z�(�
0�y���F����%p�hYPɌ���,�H���&M��-�ul�:�;��2|������F%�M���]!NE���T����`Z����/�Z�O��+���Ǖcq�C��s�~��H��%T��
uȤ@e�i�w����Ni �WG��:Թ	ô	#�S���V���0�a�z&��aI��42PBQSY,�|A),�-4��lh��b�����g����IZvO��G�LX�,fظijK�Jv���n�3��N�C)�l��BH_�q�e�0P�t�s�8O�����v�AN��'�\���<h^�sD/��c$���W�[�4���z�;�h���b�g�}X	^Y̝�S�r��9(�D�;�m����Y�Ξ�3F��o0�0Z34ꓗ��M?���3�����g�l���Xg؉�>�M�y^�WW/�qZ���A��@��.�i�m���kq�b�7���M<�����2�Į"�t,�҄�@��z��.2|��)}�
g?�Ѧz���q&*�����ţ�,F�l�4��g�2�2����f*��5G�Gt$n^H�R�7BӒ�t�%�K��Wh1$7M�����*@_XFmWQ�p)�y"���|�SbMN����u��(���AW'ϻ��c��޹>ُI˺����ߤ�n�{�b0��vs{��_�`�w;�6��ʙ�����o�q����iN�M&Qֳ!�O�� �
�+e���J��Du�	+*N��Y_bD��$���x�=�O��UJ���nƐ��C�7ŉ2Q_�~��/�ςy���'�v�&�+����
cߝ/���y��I�[dbje}X)2Zd�g���o�	�� ��j�l�=gBB�y�g	��h��<6mE,<Q˔�8�-�$K�C�4��Z�	��ԉ'#4s7
�v������'S�0y\-���P���_�q{o_~�ćҭt�%��u��B=���RK��7��,۽l�+�ý;+@���n�H�ن�AI���U�cKy�dw;�L�1|$O�E�4��~�j)�@=C����"}s���=�p��@����bde"]0����j��i�4,������e]�AǙ�����$,{������[C��N���OAA�m���"���X��/Z�8]�-I�Kg͵ȋ�!J�v��8�����p�W�9\\8��u�dK�D��v�"ذ��:&�9��%�O!~��� �92τ�b]����g��ǀ�ŭ8Y$����2��%�)�\�w�M���q4��F[��~IW�j�!��@��Ȟ�܅�mQ�!o+�X�mT����GY|n��I��?w��R�o:�C7G6���E����;��_za�ZISN\��$�#F ��N��f].��zѰO�C\�Y&U���u#�Q�N�ܱ:�*v��p��ͩrX²)���p�]KS�!�%��}_��5]D�~
�����c���e��ˢ��8��b��+�=+�'.,��ơ�	5]K�E�!%��.9O�q����f����<�d"�X��m>A��D� ^�E����CO��!F"�/9���.����zG�#��#��G��U-Jɪ�|b����JFF=>1�����
��v��'�f�	̵=��?�W�jlT��I7[�I����|W�e΅%�Fvk��UG+�S�zM�(�Ӄ7�[�Eo�F~��ݤS}��뜶|�=u��O�U�o"�ɷ�H�2�QmC�g����� O�Q:N��
���Dg�lv���d�M��7�e�Ŭ����-W�	��`K�=9$q�Ǳ����?!�a���i�t��кB&{��{�{H�b�c"J�
o�I��J��R���	���ِ�J[�`�gnW���D�J�jҎ;���b�-{�+�����M�խU ��������P}ϣ�@�$$�
ӥ�@R��qz��ZRYP��I���Ut�-Uxcm�8h�m^P�<e��,�NKJ��|I�x�T�>8
�R�����������\��K �$2�R0;�=����^vrI�#Qm�U�8�_7߼ޣDp�T8fKΤ@�El�x����������Ya����&W��Cp����	�D��p�d���6Gy�+g%D�U��5��A�|�8�,/I}3�|��Wҭu<�f���Ɇ]��Gc�.�W��qʆ�c];[tm�'�4B=zs����J��ٮ�V�#xR��[[��Y�U�3;z� ��B۸�7��
l;�o��)B�	�_�Q
�`�X�L���������z�~�x)�=�|�B�Ϝ��pO-��~,��_����^�0��[/8��(Ŀ�TF��}TU��ޘ%b\��s$7']"�N����F6ՕwE�K�4"2�S�\�\�ݭ��A<'_��ٸ�~����`X��#`�<"ˇ���Wڶj�7=b#���SF��}�a���ۂ@���e��%���+	~��,� �6�SWW-c�qޮ��'{���]U������^��X��oC�L��ˬ���~��
��ⶐ5�2I�0�ɟד�F] a�!��*i�D#��-���&��}RL���/�IM�Z��/�u�#�&������Pʀ�a�����I��\|R��!����$�L(}�_��h��عɷ�������=�*�TA�,2��YZ{?������P�)^�zPϿ�uXF�\�3b�9�o��}�q9E�Z�2�Y�TZ�ߛ4b��V��@|��O�<�U�c�'��Ԅ�xSI���Zum%�#+�Ŗqp"����w:M�<�q �BvXw��X#�݀�_��
7�I�����)�lY�����uYHt�E��!��.����S�9GGM��t�� ;}i�Đԫ���8�x�O5�e����)�q�v�U���Q�QُS�2G�M.����Y͕3�Bh������8������ �ah�i�/V��]�"�a7w̡N	Q���^��R8�[L���F�z1ٝ܍��J�k�V �$���JZ
��;�B��:������&�g�|*����Lժ	�x�̓�U�$�u���Sq�g�a���Be�������ti7C�\p<%�%2�����'��o�f��F���A�hh7�\�d��Ѵ�,��m�$�� �'�Z��B����q
^�,��{
����$&J=�ܱ�JD&��Of�Cı��'�S��m�f�����o �#���Q~Yp�u��sG��C{�E
]��٤�л�r���?�<��"�ZP��4�ųֆ&����h�x&�s�#���1�+��c1��D�K�`�r���x�x{�����G��R������؝%:!�Z2�	5�A��r_�>Z�G���>Q�I��7+�xs@L�Y6뫝B2 m,4��ܰ�{��Ioz.���3��G�
�D�/˄[�<0�i��j�`'Ė5"����ݶ���G'��|W�i���x�ǇI���������󽇲e':�D�M��ȁ@D����%C��]?��Hy�|�M�mҸ����[�X@�~��5��hv��'B%��z�����vue�b�XB��͊�z��-Y�ѥI@"��P�-��o��꿦WR��>��L��#�J���9�Ċ�޹�T����Gj�������)�Ӷ1���8j�|Ԉ�P+=��*s�m:��4�"�E�}u�R-����A"�c 8�F�~Sav,�^��y�Udb;zf)o�?l)F8Wي�Kj�� )x�c����VP�3��%��L�lޟu�IeΗ�R]�ȃ��e�.�i�І���I��I5 -�1c@�+��]"���Ē���O���ic���j�dyy@��Mzү7�D��ژ�Rd�ڛ"nJ�7�U:�qq�q+���/eTx�����s[�"	�jƬ�ug�.���[L27���>Z����Z� �J��m��3z�4�xD����M�$\(������C!(�������<ڎ[1B�����V����wP��/Q�i��eR�A�O�
�lW1���! iA1��y�F�<�)N�t���>W�a5��a<��e1�
O\��R**�:� ��=�� ,��;O�L*v�`���&@�u,YP�}sl��9�Bao�����$���g$m"<=���p0M�%��z��FB���N[[:�!Y\�s�m���e��M{�R�^�9��F�L���)�\��&*�Ԏ��1�����s!�����]&��=m�x���)P9Wq�NЄ��m���7k��k���Ũq�)��~�䋷ЪbZ�v��Չ�Ȣ&n��]%>���,��p5a���u�QỎaz�6�$�R�w�{b�4h�_d�_5�F8���X?����.��������j�W��Rg�ױ��$C_�^�����D���H.��E�+���I��l,�����-�!�������1V�΁��ə��L{D���L�ZSQ3���@�����nK��;.�[�K�[�Fb4�Q��Dc޴V�c�U[�����M���ɑ:�R���o�K�lvL ��F��:ļ=*=`�b��-��ϵC��� �yϋ��o�)�Э��!�]�������f�Um�s�C>!I�r�7=V��\���vc�g�k1�T$]"lI4t�]d��=��"/>�rpu�_뇐����/��E#���m����Mn���2r��s���&CKɮQ��4��K��X:��ˉFL��#K&<�t�يLW�Oe���o�ÍEq�������ܕ��=�A&��c:uv�j�@���~��&�Y�E�0�D�Hٮɸ��t5��̱t������gኗ��y .�P~}�YI�nez���_��,2�Fa��@Zڼw�?=�`����Q΂�?���b��B�:@^��Zʛ�&�G����� ��9�sC��N%�O�+�Z��D�d�vd<S7�Z/�G<�(H'W-[jX�P�S\ƹ&n��U�Y�=޿!̄	��0���N��M�� zD��n�|AeO����7\�y%_`����%t>�\��Ն<s�&�4b�@�%N�W�<>�︾ow�y��o+����G��}�di�tE��(q�|��*b��eT.Ij��aWG��A�@4�s��"�q
��{������6\p�v�7�s�uݦs�����U��=�`��x�z�RK췧&�S�S��������V�d�w��b.���F]o(9���&����������W���JRV�N����2���d.v�[���v�#��f/��n�A.��EX�~<CH.�	�A���WJ�k8x�Q�ُ��f��
fRsY!��ID_��txc��� �>aXgO����h �=���=��ZqNC���[����6�
_d,;����P���L� �a��7�h�d�<][S���n~�M�Y�~�$UL=	�'�m��#�	�̦O�P3�-X�|KU��%����,�a���H�j��ܑ�'����wӏmK��^��>pfJ��n9��u�I\����ngZ�G*�y�W��?3{�|�o,��������U�	߮mh{�V�Q�qoٍF5��g!v��,�!��&]`,שH׀0MZ�/;Z������a�4?x�r����%�<@��y��څ�o�w$B����$�iVh�}9VӚ8�
���Q7�h�|�p ���Fܩ�)�C�i�dPPPaQ� �b-P^�8D��ɸ���ڟ �}L\T�u��~��A<�,� o��H=[����q��T���﫠J?��C��2x%�5z���NZs:.�]>��ǰ���c��o�����V24���
5�G�i�=Ӧ�{L��QH�4�P�DnR>S���]~@�g�$�l}�PyW��3�]�����S�sc���u��LJ���=�Ͻ3{��6��Yr� 2G��9�2�jŊ��߽-���|�I��Zt�� ��?�1(��8#�$�����ܧ9ƥ�IS0���0Kv�9�S�
���9w�o��q�fo1��IT��4��S�����l����\�%�(�jBzҤ�e�A�v��*���U�T���o��bc/����ѷ7���9���*����I��
���[��H��]�@���?0�l�de��z-�G�4l��g0\��p�_��K���Ap<ŭZ��ڀQ�c>����]p�>L�B�Ҙ�ݐ��b*qT����2�q��&���&�~�FQ� ��@�3Y�9��P�E�k��1����Q��Lz�=����	N��F�ηU�5��"|v�0��v�M�sL}P]j�\���d����)B�5�dL�)��\|�xJ&�Tbgk�Z�C�]�*�� �B�r�_����x�ศ��b##.�Y�kOz��3��X����P
E��@LI�/��� ��鐚��&7��,�d��5�qb��.az�����ʯ|���%RX#�5,��!��^�k*$�G����Mxl�w�ӱ���/�K�f�N��$�-ƹG-���3b�%8��|G;����$ڒ�DE�^Ĕ٣:���@B���E"�WՏ��4����E�FK���CB�h�3�һ�o4���%6��x��0�#�:��{�����5g��^~hIw��`
.�zG�Ҿ��{�m'�T
4
F�ZY�hю,fJ�N�TzIF���k�N��7�����~Kʔ+���=H�u�Q��/+!�1�3���7�RR1a!՜Ǜ5�}M��T?zml�_�:�t�e���. ���5#��'�� mcˡ���A:!�u3,:���}��e�P��(����{-�a��q�c.�3Ǡ�������	�'"�Ĉr�)�v X$�h\ފ�i˿Q����seR
E>��c�������)f�I��/�n����;�ء�,Ǟa�U�j��n^hD$z/����ζ2��)��ƌKD���&9�N���A)z��O_j�]�Q�r���bXy�wW�J�K>�?�Z9��
en޻�+mFj��VQ2+<�z��D5}�p��Mm�G�L�^��/4������H�XE���=Y�c"������~�Q�g�m��B�~��-�_�6��4�mؑ1띹c�Co�7n]�5�T^?�2{[
��l<�<*�A�;}�^;5�[�Y�|o�ݨ+W�(G�R�a�6�d�t���߇��@�^�[=]�!�nި�Z&$LT��#bG�?Z~�#�T�Ӆ��nS���,���~���A�ݎ�#��x��I ���@�5{�ӄ�^���K{�T
��7��[w�9g��n��{���yy�NDX\���!� Z*��K��؄��3'��Hi����[n����n��Vt@8�˟!���>e�"Z.�Z���C	���'�_X�f"3�)$ɽn���طDPݫ����\gQ�����������)y���ܬ�T�P�-�X}+��C�X�Ńn$�}��\�1����Ԅl������88�$W��!U�A0��F&��^{z�Q�Mc��,����Li�B]l"�p�=����� ������t�U�0,�N3�/� ���բ�<�H�����[�9E2%`/]����K�47M����n���N�1���k�i}s�նy�W(�%hk/Rk��_��YW�ڷ�S�@���!~�(���Yl!�f�^v3� e��"/#�~����.xM5���a�\y8ZH���)�N<>I`s|�0d�H���E����)��
'���nۘ��R�-�ۚ�5�/}�_X�E,A�B����O�o'��� ��C�@T��fS�L�8٦�K[k���_����ҎY����S;���7�@��e� "�����i��(����ܦS1��hD:RBMI��oB{���#�j[a\HP�>!��w�pU�x��%Ν~�5H-��G�>+���#M:�ńAS0ڽdc%��FR`��p�{0G�8�P�a�R�x8����}�U^��20rB���F�}ĕ3����S�sY�^OxdQ�.��n<g�a��/�D:X����w� 'E�
UU�F_*��𬳽'(h��F<@�_~Z����v"Zx���iu���U�S�6,�h?D�z��:����#:�C�vW[w0�ئ�\�_�QY�j!�7�=�݂�7����ʰwZݗ�C}Eyɨ��@(�t����>:μ��UsL�7�
�x�nCPP)3=�]�?�~�j7,�.�+�I�F���C�a_�-e��w�"�oF�m�C�JX�]t��Ԝ�W)����3"9�Pa��J%3�o�u�7%�����D���C�q��U��O���
��`ԃ/�<�w�	�'��&�����']-W���N�����EFZ���R6�n�=�"�A�6�'"��M �b3(�%�I����Z�]��ڥn�07Ǯ[�?*����J��ɣaq��~�04�p�
H�3��-[�@D
��1�x\�ǲ+F��l3�Wp2��.�����)|�������=��FJߊ�H.����H"����j~�M�Bz���^r|�E]1��4c���2���m�P��ɶ�AC=}:1�,O&������,gY�ѓm/��Ś�bGO��´�2sX�@f�t�H�	̱��'��4�{���L/"�ۄ�k��u^��ELOFqp�Un3��T�Ҵt���E�}�h��:���m�gDNs�f���ȯFb�)�6����a��m�$�8���ƺ��as��,s��f�e� ދu�ʻYm,�,ʖ� �y�ƊGi:8Z���A	8��v�#ԟ��	-d:s���y�+0񘀀}���1Zd&N������E�^7M�ܵ��˒9n�c�7|%��O��dҺ�wrWa �.���J�S*`ߵ���v����ۈ�qU�%qKJV �W�˘��r$�}���}��!98���W�\f1���&��>���Y�Z֠:���t! ��W���i�d��������Xo�����@�_�P���R3��6wP"��Dk�����>��!£�ٍ�P��i�@����Q�w!|�#h��#I`��7���@�1�B���ɂ؉L�W@1�W�z����Zm���} v:��'D:�/�]Ӫ{D��B�w�D��L�������"1�t��y��x�u�؝�d1�=B\-�>!塢{��9�(o5��s�d��[�B�yF,����s�?����_�T��C���Y�}�p�N��~8�9�:�Ԏ�)�D� ��I+��k�<BcrO�� ����+��Iߏ��`k�v�勲�=�"�B)υ�\����d�]aa_W+I,���{��ETvM�m#ʝ�Y_���LH�m����=�usUl�Z�XI�Ԝ��8"���,ii���}G�GbPq	�� �%W��jS��?�_�v�3^Z���p h�	Ү��瀆b���F*
7�� �k1[�62���]^2����dXHa�y0~Nɞ{$��s����}N(��mY5ho�J���C7Vs�QJ]C#c@��H�s���6ӂ�o�u�<2������U�&*�inZ2M~R���}�k�D�f�����!	"�Q��E�D8[&R���&���4
!1�+��k���������mNea�	���X�"�HipYL%w��d��nUW�����1~/��+�����F5��~e+~���lN!n6�Y�%�]�T�E~�$Tf��t���������~w�(+��hu�i�Ϸ���u?U��/��)8֬7���Ʒ��{o�k�z'~ߕ����s�"`tc��#N���^��_��9�ޥM߯�E�3�^|
=�y��A��h
2Tݭg�J���E�'L��3$��Gk���I������.hf�9���1񜫥�ڈ����{-�WG�*�L8]�z��Si�N������<���1�.��U0���LJ�(F����gVq�����5Tޢ��h?q�����_F��?�.�^NX�Ǟw�����R\�SwX�&�U3�#�,�Z��};�C�1���I<hHKԳ�$�(\������֕�,Q�K��`^�S�y������.�uK}.�]&9G�Cn���qLL8G��ý4T��?��Nu�S�'�Q-��8��^ܐzyeޒX�^%��X�������#�8�I�A��/���%��;�Fʎ�/��L�Ϝ���hTdj�_TcFW�&p�۵�/(�nbd��V��&��__t{�E?\�O���kb���i��`���`�]��)��,�B�Vy.�!y����LI��{N�nP�Cd
��K��V3�8w+A'ya�N�:�	������jQys��5��� uX�k4P��7�!�+�����V�X�O�e���Ǎ��a�l�4{��h@׹r����=5]4�`%���ugu��w"�%#���m���,>Vć �?���ޒ9���\�}����`n6� 0�`�q� P�ɼ9��'��R|�(Kt�t]�,�Ž�����9}R=�����K'!l��{'��f�n	�~GQ�/�C�Ջ%CW4�,$7������x��� �
5���G���Zh�ᇣ�2M�
Sk~!#x��׬+���z�[Z��c��+�Z���@G�eZ[<�:����N��2A6P�TZ��1;�y^��'��u ��	�@��ޱ�
v��;V�uR����N�nuN��ؘ�҂{��[
b���a&p��ē�,K�6;��7s��H�$[$ݕeU�����(��xs�ŘHP�u4�{S~�����^�}��}sVĠ��O�#˫2l(L X�������u#-�i�����'Z��'�@������}e�,��>⸿]�;�!� %�_�oe 5e#�-�+���$�$~(_Ƒ�C��1�0���MHl��a��-5���ɢ0�&���-����Q��+*g�"��<��3�ؘ���
ၼ7H�ݾi&T��0�M��J1�\cÿS����Η/fB����H'�3�f�os��+��>�A��-��-�ꠜ^.ߺ= ���D��|,(''l��o����ZUB���ہ�����Dz�'�2����i{�Q�E�S��M�E�OYײ��IA"�6����pg�Z���`��N���F�?ߓ�٘�F�w莎�W#�e��]�|�]~����Whp�Q��̽�(�����sA��s��oS�.�����R�8}-���v׃;1Np
yF��Ζ���3 ��p�xQn&yfP� X ϛ�p�<^�#TM�&����a���"�aos�'
�!Z��)莭�F~�ܺ���9��r�A��`��0��܉ =�4�B�V_:�^WW8��œ�i��;+��#�Ɔ��4vT�gNw1���+�,n��l�~�<T^���z�1�6V|L^�c���m8���KxKqS~��R9PF�߁���&��P�<W*��$����N3��m��mlT�ś��靗g�i>�HI�"�M�����=�	
]�#?��.��.=��w�5��@�B��{hv�ŵ�(�}����T�����^G�"�1�E`�D���� >����i�{^�.�G�a#۳CSb���}�����El6�ZR�߿�-�`x��4Ϫo�e�Ȗ��S}�=y���T8��k�`L	�KT���8$�y�:�ω�s dY����4r�S�
f�U��1>�DԽ�����l�7����:�\�@Q�r��ATA}H2��,�-�m=Ezu޺��->�s��䰋�]�p��>G|��|��/� �����z�u���J&�[������a�i�+I?���h�ZC�Qi�w�V�&�
�}�DIN�(ļ*�$N�8a�Ҥ_~��$�,����C�j�Qo�o)��5�y�b��*��'�.�~S�a�[��~9w^���W��r1*��R�\;XaA�ߊ��hєR�z��3�x.��z]f��dM�g�W��4(���+��b�OI�S�ӷ���Ҡ�����ߎGa�wȬ9��E��&ݟ��P��ϸ�4�fG�MUWcO�	@���d�aG0�����OԻ��M-(�2�"�^Π�N+�4��L����p������"e���
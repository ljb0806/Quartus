-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FCCYWog/44A+6K7XFF10doJJ7IszOxAYo5trKoReF+KDiXoqM6ATh+hlmSTTyvODtyYj12d3e1WB
2AolLyvqBtiLNy3jNaoy1tTz7QCEBNN2NQiuTjgMf7PxKTJp5ned7ujmWwiFvrHEOH6MTadJOnSu
S8MWisUFJnicSqO5EYLgpQ4aZX23V+L8rOnYfupT8i89v7qHBozfkcTPy+OuWqE6C9A/McTO6ldt
6IMvTXHmuS2qGi5cfY/6rESBJl9bU0HMJAzrVewH+FBcViYg5alq0F6g6UHae5mzZL2wkmJrp5UD
Yd9VkZuRvexUVbv15cF/jXFRfO8UgjMCSDBfUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2736)
`protect data_block
Kr9/JHWx8EdvWtxApNCCmrlChgF9Qk22P1YWsHd+2wOjP7Kl5L8RjzIaDuijdTLd6+uZpEQIxVVp
jKqM8n8esLFKbmv4DM3H5cE6lqynsAEPTbH/eSP0d8BOc1aOXyW3LnG4H/WkR+XbuD5CtqXdN97R
RPLw5dORZcfdp1MPVDQ2NnYeWYd/5NC52/kMR5A3+CHTWOPlm4oyWVdaUQSnNS+h0puzjJxQC34r
j7H7dGabkGFjTFLwz9dy+W6Plw1i7SBxCXq+YllRhXPTLqXKrksdPZrEQ+LAdu7cfCYLduzHQcY/
hMjpudAYhr4D4nsxEvY/m956IWocEK4+smeIwQJC9uaqmsQ1Cw8aoqiMzqGA+sFCyKewMwzit9+S
098Wf/Hi3JrDUC0HzCzjrYTgH/M/RIKASKWvy8mHNv9InVlgz1FdY9aPUByxYhWJsijjGaFGgOSM
QGi8GwoEUDaGDavHYLdYxHe7gWUIxJ//cF0Ejw7mg2+6VE0MgQiB7uAChhU/RxDsN4ZT8nyjShJ6
X2n/jMMaar4yXw59crTg1yH0Ezh5I3WqVt4TivaNpz3plsLHnS1YN57EqgDfCaHWiTAbbXwXl5ev
zg8mCoTiHQl7cWBqifVOHgGK8dIvL7CmCe4ybi4G6uR1QZKRvq4eZgG/FXi5BeaaGR0rD0ZqZar1
QCQMzgZ5lGgADJWQ1pjnHrXr7PHb2IomR/YsdrRoy4sD0pvr50mYqGIpjvH5fkmSos51zTj74gXX
rZFtd9ceRI726HOKNKAVRE8skq11ORy3EEYDPpIbC/8uya7+tgLU0XWT9ogX5wC+3s1u6/IstKkX
YP0LHXm9/gVEF+v1IoY51WtPGA2GKPEPS4+pDkrsIR71aBy4/WVQAcOuVjXh9uCBBKspqWTHL+nQ
6BxYlHgNu2Rb2GT8s1tacgBLuQvLnkY2RSC36NqA+TlLqYFd4BxC2+dfLhxO8rWBAOvOaq1F5E7o
bd06ax/r2AZkpoKpFKX/KJZ+l2UujBoOERaqon0OkblVhF+bhe4Zev4+ctQPd8GAar2Thsz7Krug
5VwOa3fQD3fCYYkPG3Kn8KCxHMKKfrDp5RWujQEw7nOmI9RMywB/V91DYldRdMLPujb6gZNcG2dV
BKS9GvE0IiahAp6eNbk9L0ByLEkIeV3+vHQRrVHJk3Uljm9vIUmKEsiyN/2ye9kMjPuvWkeZN3dJ
tNidljEjiSLBE+HMUSTbK27N1p5kgUe7UaazYFbu0SgFzo/f1uNXyctZE0w/+zXRGOlwQeY1leY4
oDQXCWRcVlubXjJeSg/9uVPtGEoLIqzYz5xZu+0X76hdmKd5375YhhSYutDU0UjXE5J3DwGiyuf2
3NN4mVrVZz30tZw+VApv7QRSMBzdg+s8XAsbSltfXzcy4//kc6n+likZlXT/uvkgZQ5ibNthVRfQ
DBBv7jX4h1QR8xW+sp4e2o7Fy3B/rNjfCa5LGuTuRBfMg4iM31l3aJ5BkMtaCUSVzH5WqIuYRW5x
2mGxucx8qsGh/c6ZzJR3CZjIuhJVxq+1DwwBVqGqAbVOcM3hA9LSkmSejYwTvDd29GXnlFDrtoXr
tINXPz69vTN8Qd/yL1m4q3YpDBh2NgjFfmNU3c91LITe8cL9CfojH7vktYCmuHOstjU3c41utTDy
QRwHhbT2zxBDsnC3P1DiCJFsaN+w/M+fJX5MDvJXiMGvN/kx0Yq2cNaQNaLGpL3HzLIWf7y0Cnj8
TJ0Z0er/icg44wPYQ4t1GOdjituECibIG8aC3edSSMj9kkV6Iq4Dm3WSi5HHlDnfYlRVFsgXYrRc
nwVrqRgcyhCMiPs6LdH5BSGzBJY1gCWw9HOn7vqBah/TP2KAhQGfD3gmE0odNvfrYq3WcQHZqsoY
SWmdZLFKS9YUGVCf6JgxzkkWWse42Uz/XWEj/mtRYSeUZftqpTp4bsg8VNuFMn2zZYoVODUKdUYB
apHOq10guDjpXQqcQrJvhOjq7W7zu5higabhfTAckQM6baVn+oFQ+T3wunjnrGdOOGdncXG0DJVU
hHOLh5jPlsYRUKrihVlWmgWs6Nf7RdA5+bPOh1xumkDmOouo+IMfI7EGsjZAjy/4BE7EC26eqXtV
eKQrCck1F2Yhnn4Va/WnXOOKeGy8yyGn5fF5EUb/FuG9LFoWEqW2oltQydgy8Rp6kHhEsGY92Msm
+famSym2ofvqGkFI+Th35kIVHhrtxPwYjSpWV4dR+zdlkN895TqSO+91/ujezgofbOf+Qjm8Nyhm
jz8uUpxvSFl0QLB9cvoEU4p5RXA0iIKHQNCehJ+/saFzMc0PUI+yxPdBQGsQthG7I0hE8fS3m7yf
ps1ocNbUI7+f0sc3qm7uKBops1voBjHz8lqVEuNQUkh0qNz8TK6r2UPie4nnsQ02NPqpzG24+waJ
VSq9XzazoGNMOakJoHa+uk1bPevoNi7wMhOaCRuQORaYF+R1Sse75DxL9BdyshuOd4uDUnXMQlqU
vuSyRuV52jwrhlDb5BhYlr7ExoK3iauFyLE5JSzgLn6LLk/CqYgQiLBbBlJVPe/d6CjMGq29jsSp
Xkvl8jI4O7lHG/2aVyfI07hJf6KMSOTbIvRZXd5XraQcs5DLEcKZDLJga/bbIA5VTzLyVepYWnCP
iRvL3nhigCKNCtSqdS1knXfIrlgr0rzNYvUFGH5t7unH1UzzxTLFOVLQsEeKSon1V4g3Gu//OxNJ
mz+iLr4KnewToS41MJah7Hi3ruc8ny0t6CbJ1v2I/35QPeBkAP0E871sw4QXWI0H5fdn6M6qpoyb
WxvgZv3Svr0QKJWDxqHBSEfouitOVtPQ0ZAYnA9y6Dlgk6UudO1xZCGA99Tzv3m8bfq9TXL//kIk
x2MnCYEaNHUjcRuyfRV7NQk52LkBCHPa838wAJL4CbZiuwiapDZ9p7/9DUS1LVpXM2Cb3zzvLtck
vu20m1Oy0TF/E13w2athC6ct5AiMzssO6Hw6dG4J13x6jzSroLppdv8x/gDId8P/t9MK+ky0wNVY
YiqVBI8+wFpqIXlGFum+LsuDhcZxjUiiAv0BGIQbBQKxwbvaz6kW0Cc1S1dLch0OtkOwJavVMhSe
EkoNp+oNjB3/baSP/pvO4wMbDpiaL7sZJsDpNSc/RR7Kax3JknawraQRnnSOy9d6lObY67tQz/N4
jEm8syeSp36eWm4ASLMiA5mD3VMTkXyeyHZBNZia4ECj9wTdphXKFBjbpaJ9wMcOY0jBKrXh7g+o
yzVw/TLfbCvHwAi8DLZyYrQLOgrLG+sISF8Bb2H0xGPCIVCU2KFsX5QRSjzNzWoGfEB0WP4hx9zq
3qyLi9H+ysuqeqEt7hgOCF+zVlfzxyrpQfZMUN+nDhNoOn6LPhCMPP9JHLurSgqLiWMkE9VZ+MDu
UKcftQPvsqXkzRmFuXJ1Vgvor0JAYSbO85iw/Qjf8hF2/+eMmN0e6eyr7qB4hIpzGD84xlAbFdix
gjp/bZ+o3mKQKsympSxCwNQ/5NbzLP+7BbvdABmOc6AZv2RHxT0ImaLPMkEqHf65lT5+bxG/tkZV
ds/ETDE+0dk+nTJrtkDq5/mbTITNNUKKxLyOeAXXavXvMOdyKVfzVwFSQvMgXkVKTSxsrho06OHq
`protect end_protected

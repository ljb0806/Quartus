-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xy2n9Ms5CkFNx9yeEVbjcPaqVkP/NSodksgvuO2wmT1JHwCeJIXGI4D8AuRPHpDFyvA7ohpEx4H7
9GYqojH91XMLmi3kM5zsH356b4Rj/nROb6TpZ0ovvwRYUpUVSzsP21I4VVqgE6UrAbIUqGFNfeDg
GWvgUujAf9O32RvIQnHXWMrxUAyA2X+YshqJYndVy11IZry6d7YsZAsR5H637JrKpig4FTzC8usS
5xEmQCgcx9cxc279O763gkX1CNGQDHZ6faaPw7bdKADKa+Es75y8vTGbDzk271k/F3ICVOiCAwNF
x5NIvmrzyElmxuLj277wNmsp7S5tOjpfSPbRNg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35728)
`protect data_block
Arao5VRgstVv1suzLaYIeFuARuwMhPHRvO7k6galNNqNY/82sCGBb7q6b8qYPzW0W7haZNu8Mm2A
woON0de1hnIFSiPkCSvmXaiidnAkP1YV5RsYEDuL2AhE1gNFuZT9Dd25ja2WnER30UjABKUhSVEt
G9GmPbXUHmIz+2kNYOzs0VoeydbvIl6606U6aaUfcIj00q+E3wPye4k+yc9mjxBO9AgyT46PI1R6
SF3RhsRNTz+GVf2IN6f7jm3c5ZlaCJBKVta/sxMzYk7S4q1Hu0VBjnSOWoWd7mw32hdCMHp0lY9N
amcSYMUfeAJ+sIJ2H4MmYqr5qRTTUftGULVyLsAAozyYBTtJZ/BrYRc4K1+e4+V7HR1VURh+NVKu
V/4wJOTiDnni4fVvDly+x/UA0/DU+3GZF6dtRveLlpg7eATrLyOdMvs2+Tm7XmrL+MZj8QfKDTii
3rcFuVOHKVdKRYazy4SDDw+vRDDqgGNH9YL8aaGOsTvi02SAlYVO+L47mdX5fg8CEmUqolD8+cEU
x9Pn5I5RcUajsQMPm2DH0PQRvDG0U4raw7E0SI8s2C/6xBntHpFdI0rptlDrqo8FMM2lC6iNka2f
WoAd2VSlNJUB+hQ5UPhgyBOh589l8e+l+tGUeHbfF2Wv4GOpVzIHfLBTJB8ItxoL9tkrwZK7LniZ
7scjuPfH0jfxS5YnrAbmAEE8GdpnoAMDidtX92ZxI4bX76VWDRX4EYijPdOYycX5jP6hhEnkA8Ib
ePK2kSZteZtFgUqcRkbKsAZwhUBCYr+D68i70mtUGL4SxhqdVwbDrYj8AAHZASheqrbp49GfmLNA
MJGwTNwgtNm6VYSc74cTbkWpzd5zGBD3K6af2rqiL9B1FjIdPd8w2SUdqSPc/fatHZD6v2smU9B/
t4Kyw44hclZqCQdi0b/tPfm/xmLovVn/CgXeXsgs7pnsj7y5nGmNvrB2WKBRqzcgdKx753fg3D38
dO/8XJ5awYIz5vPr3X3peRpbKRWf554zo7OdRp5ZAzm52Z7ZpDmUG4YgvOYbh+5xVhWcu3F1D9wt
Eftn5B2WljdzRbeTYDUlorX6u4FZRGdXbDDCcUCR7AeOyguryWZSDdX1JjCAQ9GqPLGCtvT26WZ8
EPwgjFq9h7Owye/DZzE4YvpPCREdVAZsTv1bOPhPksI/gsQ2fwzgv7tHdFUjSa6dziIawg1D9IWk
fJS9yGfn/A+V5ApRDTIwSLeYGqpaM2q3dGZ0B1fmGumFE3I82alKR2iIfuLKuANrVXzT02d/WBNx
j78zBjC0ZkBapilgNrONiHr/yGxu9IIOEcEB28jmatSJljBZmEBDQEveDMThDzBxrfVaXm9hLgWF
QJf6VBPbrgQwShtQ9XWKfQ1o10CMici7dKwB80n2QQmqb1+3kCdhR/eiIEmKUzilAP2mmBctgPtn
RKNFj9ec8jaXvk8ejjgvBaaS60Q0n1C3dDGG05Ul96yMd4wN/hbpqcjCpHGxf8F4XiYWTn3kDGqN
CgoUsPzTct7bH0XjaT8xMTlaZJDokOfQsHcidU2kNBHeDzSpEk3oWf1jAuUOJ8ghOCCuMtJQh6AD
cbGWyFqwV9VEmcZmB8w0PS+/jHoAlu8s0xDC4o4qxjv5MeGLy2KMzBSmtABioXiScf26O4NurCNt
EEaJMp60i60doh5Mx7M3EPEHiLMxLCzK/fZp37eUeESaBe88Pjwg6rIQKHb1v11JHDf+B1bWLapw
OBN2mjI5HJgwTIKhCMIo3AmBfUM/uzz5m63nPQKhdfsB6oR9DBcd8PrLH2CQri12HxEbedCBcTco
Il77RNDC1zjWjm7IELoPL9q5PWwb06LhxTg9uGUHino1IaDUSN36PcUuXREODPM/PDgjQBHt6PC3
erpgy3eWuiHfqXtatELyWusUVi49xQyvo1uO27Jrmvd6YAKl8j9j7Tzh9w13TFPY/HA8AIzvByuk
ZUhwJF8cxd38vd0ptzf906XrujmFufyCRMF6IVUDMmW1dq2Bs+yclMu8qBFYNGScqVLa19gCqPfn
YPMU6PInMYQfpF+4yU4J+CZyC597ds9Zsi2sU4yCc+4L9ahpKNt+Pwg9XX9L5epUiY2tQb3Gdlwm
U+2pxffNGrnjV1M+P/x/dvU/Q4dG7DQZ6Q0Kp6ck7JSHWitVJ6DcmCzUxE3qhZVMcDlZJikjCOJK
OPyQ65tCEfkj5+RBasyVYi6lXePDam6xUSV/mnH0VXbQXhEGVeG0J+rs5Wb5rvOZeworBwzV0TJ3
T8Lf74MpVzBRUg6dCIP2IX5f++PxDMjzjjhKlmQFzr3rSQyHv2H4Rcx8L0NuYk3ngYi3s3p1huJM
MPKt5c8Fxoh1oOoQZXEnzq0bilGwvfr9kKeD8aSngk9cTmv/4UR7ubsRlqp9G4It9Wj0HhSThkpP
LHXFD0yReDj0F0PrJ2ISJlsSmbMpWRRT98O9uOQF3osVJxEvXLS2f4Ei7isHCehL7qwv4UDw26yx
Cg5074o6XE+X9HyrAaDvOCsAmgZgoirU3cJeMhjv/UfS4Mv8SuUh0ut1qbUMqzQWyS39zkFdFY9L
sA3kVLCD2KjPFNRNevQ24+sIj28TM2mHtnkZs6bkKZzbkAeu07vyJZAXS8IKbw9S/saJ0+u5BSdT
3OQmVkHvNWjOU/fmEO2hAZEO7l8OyujFLTUYMtKO+vbeg5Yfyjf/33fB43WVwTI6aqnajI8sdw2u
IptjsGaU8iAkRagdVN/36Jb09/3nroarOIQvs3QYuRZH4lnfAb/DNSW50LCXwYpa66Y69jIRL9Q8
W2d0HRjOD8mBq9nvbB+4dovirUHcDhPRgXU3rqmmwH+pwsCla+kiLz3lyendpi7P6pilnLqwelpB
dlB2vnDgWzAycROE3FAtUghJQ+A1B39mdRnjjgxdoprmiYxgLUTxp1U2YQPIxC/4aUDh47eqXd2a
u7V+ZvY8YI6trLSyzMu87Mz3KEhF8gS5cDGm1NBiFV+LCmQLosmuBRFWyaklOjylDQl5xAJp9nMc
+1V35I8kk7fCCGLdYZ+wBL4WcoHsT4PO2iHNL9GfEf7dIGY+5u6+tLUWQ9CwXIfaeR7rbDjKZmIU
UgBP+OfnV+XS9r2emwdujij4OpFYDOWaNDWJzbud3Thm0EsVI/Lm4hBBJj49QAhN6+uQOG2VT9B3
MtuddEEbEEgKgWEdB1rDLYwO20Bk7YuS6MV8mbqQ+m/3dr+HN7bTNj6zPdc14IGpx7dfTDLkJyML
2WCvKSx7tqZtRf5w7SyrxWMPEtOiBc//tCgC6yi1RvVSV+cfo+/NKAAHNtsrU7QTuh6LRULilcU2
JhVAe17051pJ6QzAI44T1lfcOyRhSs4PdVaM9LcrPbLibPRaNzodkj+BUa37xz8Zo9JHn0TbBTuD
UJFLzNH+b2Wktfb5HyBdiDbkZLHA8PhcCKArcmdVB7k4QZAy7lR7M93M/ra5jVdTa7isBRxoaycS
Yj/GHmiGegqYyEt7z4rkgWH41kAmpXn8ubxkkEuT1jJXf7VOnpKoLaMBgfWMCioUw1uk2wwdSSWa
vNLiREijCp5PQ/9tX84Gr4wA+TXM3J8AvEi4W8TlUjWZf/7WoeHoMFQjEQKz7u2o+kIvtgXbZT2y
L0+rC+c7MHwEEop4TNEHETU5ZFBTYK1YJfXnWV3RQdvT+2s+2UajBV8viOI/vxAkjrk3EnPo9Uqx
ZyuyKamhfCS8y89RBl+fEe7V7lCTAmax/qIXHdkHCsIcMqY/LGvsNGpbjZ3VCCQLilQR7JIaSkQq
LDIgQ1YVkHcB8e8Y/XfZ7DYyrXnnLzfIwRK+LS0pUE582lRWt5BDaxZRegeBXxFZ2Mrfn30Fc9jN
tkkjCHl8NnnHHvAzLMaoo0JANALQPBVl67zR1uFHLzYAkrz5xPOrAkvwDTgdIxnJaUO8vyk2rH1i
H8yiFRy092kioLWNEtaP64BP2vGDO0uxFcu1NTQFML4IMWHk1JanE1Bjyr1msKU7FAri0Y24z1fk
utakHDCtFxNzTRENQWg31CytOtq/OcEgWIr0fGqdVONgabyWG59F7JWXso/lX1tzTsC3j7qG4B01
OAD3bGiTZcV6ExDjKRy79f5/VAM6xJilKzZLu9af3MOXCAc8oLmoIhhGP+ht+u7f7C5YIggFUqSF
6rPP8ny/K7UvbvtNrQcVIxUaQCBYjDN1QiSW7qMgkPbgLCpKhdJCD2RzB7p2ShnhcSXSb5f74LHO
7XZrqtnVqFI3zB76det0r5cD03bjbmcpFQsDoW2krD/+jckFc/h7g7VvKSqdHGOYitFiSuvCLT6z
z8N3RB2maS8TQh+YGIixMsKUZpVNy/rYXXpNj2ULBGeUsfcyNptnRx06b1KJRazxMEzbsGPdtBWl
gO2gyGZiR5Qo8Mzazn7czxS35AqXToZutEYlf6HDmq0M+//LnyCg0CAzTeRleM/tJx35pQPbfAd8
o9bQaeZhWBsmLJ3XU5BF+pqzOZnKeF5wPDlFvnt391DLApstTFP0fVWqr3CC/zRVyUHwulTCszId
sEwStZ2OplzlZfbGNVWdSNMhXKZmVJ84QWvbA3eWzDFkdsF3ntr362DC7sRsYYk/i3KW8s8Fl80F
qJw7FjJkbAkLXphCTJ0oDH6Bw7QvjmbBM5Mw9GuHh2sWlfpD74DTFLOFcPlN2d4HrQOfB/JcVB+1
0HgDhFvjqj6EEkz/haFvo5F35xhsovyG0onQZhErbdvcjs8uHfw0URpEN5Z5RZh6qw7y6pmtsBRq
JlWTd2iCbM7rjbBYfdhFQ/Plb1fCgNk+LhANVY8HG3FXLNDbOHBLcHdEUhcbR4QGGFwNeUDJp/sO
ke9debjtrs/O1BqCYIWhAtxgayo6ZH+3X4JTMBrIyJuofk0+VIwxqIfVr+j6QqrYv2gELvzCC7cJ
jrJm1fZogJ8UIThvqq0NdJo3SEZwUA8KZk0TFxNhrP2dudXDynEhgps+GAAqu2BW1TyAcDK/GZrc
uv8nVWHmOuIqHxbdoUDwLINSQGhF5jhXvaXx/VfVLC+4yzNlCDk+ZAj/obSqPqquEFQJXGsSpzNf
t+tO5+5GOXkBPI3gYVrjbM850oDPz+63GpafEGbqL5FFc4MbhpQqm+vWDhSGfb2gZroBUGC94BgZ
pdQsL3c1sLyG0HbQsJXS/kNNs4g3EkZITu4pKI+hwdgs3vSK9AnzAOP7DXwUXvMI3a0+aEBzYlAw
136rzucFhu50u2/byDezbNhGhf0WgjeOvWpuVNgT29E6li/SgQdv0S2wWacrNvZvHRph1PZ6Htvf
x9+bMKnzie0Y5ZTwXKWx2+WzF6neXKrFZP0QubKTzc1f/NgGN9EuHRqSQN+/vK0UmUCcKsx6ToiW
gAK9JJfPmkhH8VWD3AGnwHWkFNUAB+jI6FVK5pYgsl+gChjjWGrlOG0hi/QHp6asriANw8+pQgUE
COtSXyZS7reOWKLx08DFKYcccHCNiBfBAkiD9plt8k4JIa51YFfKL6PD63Rxn/SHDgLZZWBcKDbU
g91KLGwosMdVEqYwxaipfrDJo0F+gy9izh41PWyix6W7TmU62FPzr3w9zjfeamriUIwO4Ezn2V4x
ZC2ROmOhZwEA51QU05PlVph67chhbWJQGU76BZTgd0ewNWQQSjGBPJI5tHVdABr6JSavBopxuQ19
DAnJ2IrzLvfNx7WTHHz4Xhu3bwvKp9BKKipBNeUl+YU18jC1jNCdRGLZYl+DRSlBvOm0wrHMGLUh
IHyazDLNF06PRYwnSACcr/O+StAA0mG0CuEms6MQlyh17hYfou0d2NfwBW4VhurAnD3xPSFsbMnq
M7VHYBmINudTAraGkHd1q0DszFbpCqwrly62yri5Rhg+nFrQjVFNFl36a1rPepjGNPW3SKgwpalO
PEhk/doNNXxu46jMo7fnrtHvxTM5m1POvWfAGIEi0Ty9t8YJ7+etCBR0oyOvbITzaH8Bj+vmEmTS
+cTZpJ72f85LD912HGcdP+RalnnTjr/LmAFQUNoutT8heIG8X7LAJ2UvRLEaTOhWBvULZLZPFt1f
K4R2qf/kY7gIcfHk9J8EpexMdcsZszPvUIf4MleNm92+RqSaFrxNx/Lw73VihSUk6JNnaiTVpfIX
I/SKnYZ7j9A3bML6CxxGRwRrNEeOiV3ixTnNcsUqyi7jC7AeAYfj46rlXE1LoSM7JV0Ca9IKCh2p
cUTvNlcblWhHkYUmPOF/M2Lp/B9S3hMDamlM/mN3hk/O3yd/7cxfAH70p4uvWmWgHOF13lg75c8K
ictKJ0xfPiwOdmYilGTzlVjhScu53JntM75QJWaXk0LTYtSPg9lJNML7vgP8IJfo8TAs6xtX76RR
vBSMV3bGkmeo496By7FNjrjD2ca3aYzFmD+EY1OOPaEC0W94zO7B+xXrQNe8iLApXCtQq+do0hv1
POciqCeGSauNkOjW6P8UWnfWmGUxNudBwpG3obPzl0whRJzwbg6/5ah5C8tHhLP+R7Okd4UQsfGh
uB2bYwXQwyytWXxUJrC/0JrxPBX8LLp1A7DTuDH6EFp5QmK/XKsQ7Mskio5Ug0rSv76LHyDDxu+E
Cvfw2LLqzuY/ZWzioUJ8jZzw0q9pT/whtuPXougfOrYELwbH6zXZC2APQRU8TjPkyFTYW2HWtpV1
GMxV16vXzu4OtbIRNlBXTyU3BWRlrTpEVn59fu4SF9d7blpeJij6VbGh7TAnJSq6/R8buYEgC9Ad
h+Romt5eQ+wL18FKsS96OALsWW63ogEzngyo7bwKQCMBuq+PbG1trbivXR96XOPzaPVXhwXBcvdD
jIkPha3JjxLk4sNafUE7u2IT5HscjdGVr7abf/obPbHoBxq0bYSYl5LI3JvAT/KlRz25ijQrwDgM
TWEVUmPxTmbLg/SfMDajjZs9q14vd4X9sIAfrM7rAAy3+7q2xIdoY5TKzVHBhD40xTHconlEUPm7
0SMCfuLQ8/TMJ6dT2sgIDg9Tb56SQYJH9FlJDfDoPkXUyX0W4mMfNjyCBFWDMRMomK8tV0ITxb9Z
KVL+BbmgiAOTV1TF6GydzmNV38iEKFI2YrxLPTR47/R+/EwPPJg2USwdkOoWoxRFJwXFRPCu7dlv
Zh7+8k1CiEKZnLnGLIKyav6QncZZ2ydFeQY1maAbIcNy9m+hNxaI1aOyBCmuKinj36JevT5uBzHY
bVk/Qqc2oCcMip19zbsxrUU1Lv+unnC6oiOeoo0f3IsvVsO3HGgMaz2Eww4+2Td+H4AX8umw1uZ5
+GkBhzEpTHrbhsvn7GHVPdCXoo0xeEMNyyxZOOCViXoj6v7x9qnHCnyp5KTm5njUbUaAtPf/dO72
wWuN9HFXkla+zCZozm6dII3L9EtnVslpVciGs64kMsDLh7iaICT/AJsTtZTUSyIZch7KlBfXJIya
Jzc/SP1uVonG5WoIRFCd4jB7ieZBXL9FVSz6aSVHiVQ5jrZbMvkRTzZ2HqDpLLUCgNrbnTqrjZP+
5fXunBXn/yUn09nWNWyoJ/XNJdMurJM2ZSinTtQcomBcq6y74sG2eL3X2aFvDlb6/ytCM1ZJ7yb7
viJ/bNIdrbILDe93uzFphnp7+67DFpANefjR3sgTrQu0WafqtBQ7MYu7kJKDiSiIFg0L23rO8oc3
TdlHFjdPXFrlB/qn/mZUBC1S/cxepyDrcZ55OwBVu1bJoyOy5nqKq/j/599Z/+RSSjcYoDL9p+Cg
Up4nXqZgDRDJPEwyUJlE/kDRExjRIY7IJMbMU07IFb9BoHpxjpOm/5LrpjeDA3G6tsXZ8eBebM+c
/nlvEb6idWKBSmZjOj7cNFFT/4JqQJvCKI9+JlRSRaMbvBoYmpvYzGhcZMGbmE2OpiVB0M+2hZ62
OP4rcw2dgNpH9RhVa8IEOnELP8PZJpoo8amEvlchuJBzes6UTh/x08jis4jYZQVMH5V+K6CKBoGS
xXN64tZvYKMJW3EEyak7EVgSYaMTzviE08C81t9jwgJ7No/sVtQOU1dZieTbdMoXrGyndwsBgP2n
jIcQSv6KX+3PZFFlwRVHxYVbEPUih5LxnagNXq+roIEWWlPQiUK1UHfWdC9fbgI2HQtX5nHgU4Xo
Hu8u/XBS9h18Hv+8rpLVLz6jytEZWKq5tUEq3zX/Rsf4YNeModHzo7d2z+qTOsxlLpCAbx86ftuq
lOTqWI17SVlAQElkkErePhr7igY2XesLt7rhdstghcWvIxz6aHgDvWVgnEidpOxDQf6sbIaoY+ZR
DVHjU00o2ckG2dHRR4rTOUwfmmHIZ5s86MBPiijFOznu0DpQdF8uTpyNFI+DAYqmjxaYGaGkWjbD
4NjjmYJyvCMIGOYGHBGjocoYnZNbqRFh+leAWL2X+kzSwVdXfQ1N0xf7lCAu8yG8cTxDXCA5Ajov
uom6b6YkpwHwJPj8NZ9LVEkJXYlRyx80UFYB1gbBQhSIKPZOClghpXJ3SO61OFzQdfDDNtBuBYwm
SkUPbzdjUZVpktYjofs0syKtF4rm2onJq9IlkRfQYISkNW33ZWUTTF48QjoSHZ+Fk0OjzLq1yXRC
JQxFK/Mjx+1+IrrHsl424dWAC7z3A/UxEQ5gZrCmJxB4oPDdCF4jA1AqA9bcnCgH1Jkjy4GsfQG7
xgC22ZDc4q6YGmCN57/zc99JXWfFo9pXs3S+3UucWp2mjJOhP+4BPXE/Eug+W8Vcaetr/KGUtOI2
Y3rfCW4yImfUyWwfNYf7+yL8flKZsB0SFY3U5hn169Kn9ceqN0R8Fz120yNF8j4nOQAbwlq85uIh
HVY+5NzA960sWY+VFii3BHdKYdzxOvLa/Djzhace/0wnCTfw2GNzOoc7ZGxT1a8zqVRvGrpBFbSY
aUxgXupGapTPoWKmHi44+g2ApLC5y6mE0acwTHrfC3CcBT3tWEqLmRCX+9PRiZJfNgCmuWC3BVOS
UQdw8skt1UvclzRKhWaLQ/uWnFTNZ+hUv4T5pl03GtEf5Vx6yeypGCxf6LAPJDiSlR8sSjAeCLcQ
sjkKzUEiF3INFPBrnAaTWXy7h/MxeiRm5lvriu41f/1glbmu5JMfaNwpqP43UKY140Ae10LZXOdx
IkYsy34xrSsQb25p9dftzJ4G8ez6KyiCPPLhZEJjMHbAe2Zw0U8fG1sHZVrmqVrJQ/MiADbrZ+J2
omydtDnYUGiKh31xfTYy2T/KOgdwEoQY9gYCkZ38oSoukXhxGoNTgs3sfn7ksy37JCYEIVmmVDc3
28LY9PYmX3FBJtWZ50y5qXydQe4ln8jSeE2+v+bsoXxl2TplOL/1ZKDCLNh/UEF3EPoPJ3PXGduB
JOpLisz26hADI0IuP+YPpRw06GzUwwt9qijLdN3eMQ2dDnFco0GnEwfnFz9k3SfUrbvd5lyTWqcq
X+tgixe+42rDAGMUxii4ImsT9fZ99VoAWxTY7YlP6OA2eXemsv++tlaEXDpZsgvIDBUgjUytFIQW
cKYkP5k3T+a5+4m7FWMLYlU9f5Dn11ntOhAI9Z5lwV2onnREA0aaALlbbfGu69Ng3iYThW7f8Y5T
sd9n5WjZlkZn532tNSXGhCxcIDmIPUBXGkFS7gz366ZUvY0B5vJRJVx+Db1yHVyZg9aDLWasMXLm
rUQSk2SRlNs1b5y3AzGn+UhifrW6s9u2Pk6/cqghvJ2k4RpUWkL+HQVHtB6GLGs+zklX04n6+SFR
N+Nb4hGPzLknhSy9/lns0N78mAurKAe8EPD6nPGE6uP0fzFW2NcBkzcJ58hgzn9DbN6AlgFHM0ea
RRDy3HJwFuWuipVMNVl45X9RUa6jiIuel6ao6lPgxlyqznDIPjxJ1vUOYvubeYQLvbqIKppJNOgW
N9Yubd3Sj9Pe/DonLSugLkp7RloELs3DBOd8jGbag5681oosEzC7WO4G/hVlfZuMDh9INObYVWrE
LpVWeoSV74XuBu/Vf1n6+GehtA8oLWCP4NAFm/UIzsQvbwaCzk7szXPo6hlA+AhKVWycooMt1sDa
0G3chckaGHQ6rUWnp6gSa5FmxLeTsnSp2w1DmbhZQ4lD8lgeyAnb1m0mOhM+1lsPpWP2bOqB07Zy
GaEYV9ySbTAUKnvzNwy7v7B4b9t5CVIFNPtJvoO9p/0khZyngphgqoWGlKKLex2cvwVFaTBLciyw
fEZY6QIheusXFzQffcCDARHFcoKOETmpG8WuiPqjYJU5270zzF6pdAXJrp/YFTwzck2Bhcef+5Hg
cY9S5VsewuEhdugHQaz9l9woAkd1ghx1YvLRTaBcMyzbW/BeqZGDj+/kOZgKtpJOo+YRftZ9ax6S
xCqyyZNWCGo5I+r3FZf3C6ybj0YgLFTdbzqLKgiQjn2VP2TlpCX7jH/yjApmNOAlpkFmB1Q8HImu
g/hSgzyp1EwfNNqwRZ47CGhnHIASg6nm1mYu+7FkZ4mn/zIhrR7aH/b4jHIwnVnYjWXicPLFsOk6
60bAGD1P6dgo8LBMGUOfCNe1ZI/Zf2Ymbi+ynsCDYzx53onZT5RFEHlr/ekIvprwlogUDmqel/sd
mmwjb/vmrjoq/ZZ3EGuJI0YBjaUBBZdbuuhgfgt5rfmwBr0njWKmIR+6yoIa2LNksUKrDnBy5eGT
GkQKbyCooPiZOkUn7eG4KSxE9kNVCufNzpVI8WaAuM6cP+cAj3OnbRRyUvS8uUeJDh3hgweImTMq
v/C0IKShgTwhG4M4vEas2N0/FHdyGdmlOA8JFfVPQrMmJopt7zMCvM2P+L5w7hUqU8At+jUxQFUY
mO7b2gc1KQ9kU2xNknwQRoWhfr/6kUrf5JgLt3UGOsmIVpTt5EBUYqnCqfycvnDU1L2QmU2E6dL0
4MCE7hcJ/QxCJw2twpCY9d+EzlN29W3IvTgVhl6xcatyLrGoIwLRsJFHFur5HTJGYqyELuKOVYL6
0ljTVeYs26oqPa+bdq6FwJikc092riKParq+/mT62/EvPJr+T9CWdQ6VTcS82A0DL+geaa9IfF1l
3MTVFgWxJMCu79RWlsLDIKHIqQzfSqlkmIPkTJ4+H9GIIQNiiIPj51k8YwATVmXYpFCCOaFwSZ1v
a6Ro4Bd9V81Z3s0HTAPMkSd9VUAD/eXSwszYybo0/OoDjNPPK7kJQ66mFk9LgNDiDqcMbJrjCSPM
+biSipuKzHvtkdhkPJyGnWogyQqDsWgiaBTzqy2RyO3blWuI+QdMEkvu0tVzUfou2kiU8vUt3ohw
OzDviiW5p6TV+md2fGR5FjRNS0t/rFxTZMVFOIudlPAVyCwzXPms67ujAAh7vwpSAAT5ZOXT3lfE
bEY1dUgajtK07ad2cwPrng7WhwPZ4Sld9uNU2uOZrjnIZtN5ZbcoZTxfhDe40Zv0nEGnkm1R72Aw
h2DRuITzoaEK/BwxiMYSGAqdMcLi2tKzcMuoKEAb20VBdVMIbV5nBqK94WJHi8ItKzwFWwyCRQvQ
PZVIWQv1IrSl53iyzG3iEcn1jxKK/H9XjPpqYncf0dxv4ICwV4jHInpUgMhn2EpykaLjm+0Rin5j
Ublr79dm+UOzQ8ATuvqxCNSbm7TNyEg6PiKSlbQQYnN2OpXhAZyarxpmrWs9QCkT0qSdUDIsBafM
Lt14DxPUmAWdJ9sKZwyLj5PmzCOtwgtEK1IsiBgKgoVNUcS1XyjM2rztX34Fr2WVcadLjbypaqJt
rGjGaNFZFEfz7FK+qJnVNCJZEAmqc1aPbdB5hqAFSFsFTCGxQeo8W83aXAu/jFhYQufnpZkhRI0X
55Im/bbqDJ27QfVCKMylMeqIVh6eHW0ASpRGTyWM+LaRCP7cI+DEt3rNWVS8j9Je8KrzZE3jL7ju
lo7QLxoQUa6WBZxF7KvWJHYJLi4G0J1XXAmyzo8RBlIu1xessUWrYjNNPQ5eaNopC1GZ2FJOvCxq
6e3Bvuf8zhaYCexHjdwtAbDHHn02Lb5dYVsfPGo3J4xF3B4oIm3SehU7MS2cbIwvEpCdT+nBEY1t
nOz4RN2/2t3nV4/xRBFdlD+YzLxRFpxx4pg3H6LmzzoGlSBXZMs1skBgwF6iKE09Rhb8Ij2QMEdy
g3Rr9PjlSFpyxBEe5ksHe7MBC0CI5vgj3noMqs7zhBWIq43d1w5lRcIz9Nx+uHNulAqJYRfpBgTz
twc+N47vTnAEAGDKgQOMBtOm8fbEDuKipKYELLqmF/+VsWeURNLyAloAVjwn9pcuczY30dG3+9/X
FNL+LpTCxXG/ivspPuIFS5R945KDBzqFjAjkafrJCbbtP2I0STl5pCP2vmO+PbpnoZ2i5mHUx8HM
tVQBEQT4Bn11s5sLTlzHKGCTQ9jClZuDkb7WU7k3J/0UKV0YNm6Z5fHH/uiB+75y16KPZpzQh0JP
OV13sLkm+UCDEya5PuDLyODthtckh4rog98OhoTqDpTj8OoWX8ye0B/iJwaQXaOD7Hx0QWV8YrkS
ebSgLxfULAs/cSUD+QePbQdmALEMkoGcA3UL1csnqPaH7l+BUhXpol4X034z8JgLoWkm+n2qYicZ
IFMRzJ+ZWpeoDWg9sUxaUFJbCzpSJEXukSXSZ5uCyr1p3JMJfKPATU5DdwzPlMSzltIlL8SfgItR
1/WhBTHcYhEfZREX7CB/P629IqfvcE7OsHWmWDwu1bfYD768Xd4E2RhMQtYZHazVgklVf/0sOWxf
z+CMOtMIayIzkPzmumkKAaZwZzhJx3LPhaDI65KS5ZYpwPvH6cINhKOH+YR5nN67pcRMnK/qRISn
s5Hcq7xJAXS+PNbDdO0+LnH7MfunSTeSWXqQRT/6U9Pujqi/zXw7clxzxQugFWeZ2I9ykrLm7PEE
c1D6gVeIWSScy9rLIkqCQ3MGyOlzgj425hao7U+8NFXRyjHIhsnSGuohnO6dYHCmIGoMjPlqs7FY
UXC2VVYtHLAJ0bi+vBUYMntbMlFQIhjrTjf9nNIioF9SLisFKDIQyLQVMmWJrqBPWcSq3NZ4+Z7M
RaT81SkPGFffY+SIurIelDrxUsVn2xl+hRcOhs3NNSGFv6Sl74BcM07FWftP1PPCVKV8pYmYXTZD
Epn1iG7CdCmzT0jzRcG0bNkBKqHK96/mOhjLacmnLIAS3hTZEJXzZSaZ7SjA7hpHUV264ckxFuIO
3xj76C0qbuZh1U4cUmEPjKf0UL+xVsjZ55lpPxmVflN21sfXfKtq6//Q+TLM+y2/hBOmPgBMbmyv
C8vorw/twNv7++63TOtpW7+AUBhRsybnrmnlIn0peTeb8nljYxM2PCD+0WbhwXRuH7FVM3rC8wiA
kEnQUB0PZ/bYbQUP+gbFJomffRSlPzp63H1OP8WSTBlSxHUW4ltbjx4A2NPtDUhqUPCq+qCxZQTT
72iOREcVibwD9zvEhxtJV8+cVJl43qrvN3bS/KvLbGnhMrl41f5fOzRU3+8EtO2lyoy9G9YurBTX
2yB8FNz4cSe6iOYMLRctibG5dp6WU5iMqug0FrUbGWyJ5zLxebO/9DB/m1XMfGWBNisiexz72m0Z
2RhpcLh/oSMSghNZqVnevpp8kGXSN5iGQ22XvSbtxzf1gCG0iJGxD94He2ZQ3d5SMqYF9sKoXyZo
c49Xrcz+KU1zcn+6VXLTcIXAu5BzHE1QJXubU96uratiGeHvJ+pJVzO2I3hjn9UyXccnsT7ov5Ow
NpA41YnATb+UA6RDUcJvZcjBu2tsA7z6zG/7Pej8G7TWGogGfWtQJKffcPl6Tbytpz9iCUFzT4nv
vyN0pmTt9yn6UDVsbBKOiHSqNmSAdkxr5Rud8V3X1PCrGr3D8kBhg+aQI1/9ZjtXoMYp+XN2KNfA
RboCennzO5bZT3CQTYEWve2OTvdt7FI9Zo5nRb+6Tm34aUA0EBLLULZfYscADQ9HXLMG0VtldBQx
vhdoqMqFKm4xw6Bo9Sojr8VFZY3f3oERD9BZ/Pph73AVWfg+cX0s7VGZbgm/Tc+7Fa1tob6Yo3pJ
AByPrYccuBuVI0gt6b635eFVawrwjqluUAgeIdgQYHg1uOozGpcili/8UXYnclrgN9jCbLLGO/y2
rmZn8tA7IdEpFnA3oTR15nRxT1bfWPn+YTKVf09DIWl69BTLsaPwz2nG6cSRccrwyeU0uwRs9FtF
xnk+E8mOKYb9g6BpDyZ3/3BU7vlEhU4VjK6Q/zQ6u4ryYSN0QuC0Q2+/f18ezaLsokkc45X1I0Ro
jJw1MsXXyFr6PudEjV/dX1dr7Lcbh+UkwAzXDRfqlKzQCyaOkduwifTXh5RdxratyzFwEjZ8NAE3
Y0QWavnQcLPvnVO+lYDz+cf0Orra6Yl11ALYobJmFu3tH+S304qnQnM08yQXN6rdyXSvWYb9F0yd
6jjJ/khEQ97/mghQwWfby9BU786ViIfZQSCF/EWdor9Q0EIFCT20IMTG7fsyha6nRMSVXR3ktpuG
UTny3RsaaQGBbxZk/tm9rQzp3H3XTx8xCExHQR3QD1Sse+SczSfJ/A2pilhTaiOmVK0ATvCHlrcA
+E2OHPEHW563eDGKKpso9WmKgf7xlr300JQ7gWAQ0y1DsVWuuNUdvvmQpvSC/7FUo2U8JgNaktFb
/YUVk6mD9Z+rVI/WXmUR0/l5wVUHrjbSpY6WiAKqB52NBQr0+5xF9l1gbNyJV9odgAxBCiNw/RtL
Qak67i1/H+U/vhiT8Y6pUe2O6HVDjGs+8DeNSH3urdrxiz+tvUEpXVJ6BUxwXa3UgzS/aaIpay6I
feRPUgzmsIDHuCHIRgyhlKjt0EE84EjazI9CMOtmYmc1i2ivndjNTCYs10AcKXNMGJKTXA3k76Th
D8e2hISALelLKiabQfuVj/Nm8nf5gf/ahyNKJ2FbAPmr+UinFlkJ/H3IcK4KIucFOErAslshMueo
cAmZhrEIga9t8iT5Xu8g4vIEQaTUvHhwXgBbh7+9LiIznbdl8yLtabf1lPSwT0CVFgZGRpriEM7U
LugOFTOUZhVszLaMjC0cPvWAr7a9TcMoweldGIiWZ3HZn4o7Q5RmXtmbGbgntAt1fXIugOGveS9F
b1+PXEhoeYLVUOcWg+BDNTEGibqSg+LNWZ6ENlm0UiwPOR/F6eLYUK5VNDyNWsFrJzRCx0yIRdE5
0WK+n6TWNdeVlnBI6S4slvJBkOegATHUMj4QZXJELGFNmU81k7aWyeJ/KlytuXGP2sFgMReNziiO
BVAhDPMQxpZh9cLwZXvxuiaTHGpioXUxU0L4VFWaRXOC+8sYQbFNydqGz4t9q9oTUnKfPzsubMKV
INuLPxCcKCASltQVV17nr+gd86gpBjM3gz3ZaYrxRWKrIq8dPoRQl9Kdqq9aCLOiz3AvhYssq3+F
S9pUoGrJKTbqXu1+RtEFxm8V1TeJsJC+F+Y7vzofAoaC9IkQhoS8V/ggNv2XVSoh7AcQb4HylBwP
luzV+vDhgeC1wVhYUfe8qlKL/TgDeQkSyCdYvzZTPxqkGtu03n3idy1NpQXheTqg+uxIs/1Bcxil
pUDvnSTs961mtqVkN8vXyaujPQNnpnBS4Fm+wjBiyn24EhGI0cDwZLWkr7p39uSMtS0dT2nZleji
6SWaBj3NxjInjH3Q/vm4mwJ8+SoxlJ0pf9M6//4JOtZl1tSsQ4xVmFC5kJ8iqzmzQaepsOfPmfCV
iyMhyNGt2qfi1SH4GwEJZdydqsPMyaeF2Tl/Gehw1/fJioMaEBRX+wIDoKbdihiicRYuCOVS0W+q
sJ6TFSErG06cEgukqyIFFnpuNILRtJaW2AMUI/cQzxuxoy0C8v/mY0LnvQghaOCpK7xxn7z9MoVH
4iJlyPunPNtUQHY+47BxfoPN5Y9Znko9YxNMwT+sDiagfTvUkfnH8A5DtwpYo8bWW6necXYZqdht
pWOL70xmUngEPIe0xWVuPR67nGvAaC9auZ9/0eUttETb06gloN6eHyTsoJB0+UD3lDuVQBKdkLDm
DSrV7loSwHoICcIe8QcGNL7MBCKv9HhSFCP5BFdvvxBiGTGl1HbPbVzEfB+YIMeUvtlhz34PAOjZ
8XyhqkIuz+E/shIUtuq3UkO68b5lZNmyx2pTIS1r2EzPi2KjpcI53JXMzAtAU3OWOL20XNBFjTXC
To47lgPy+2lZi0sQEbPIq7GbboQ2UbWtaNjubN4DqOVPE/8gG6uywvJfSy4V3JBUYQlF1aRawZZk
1oSmiIRrW5+x/GVgAjkkVXKNxTeNe9IFduM7pGs4QnUD5xrsinAu3HJ2evbKLf9l+hnIeB9TEy5w
6BR41B/3+CY0YYgnTtlDFfrMAFPI6hqnTFZ9/EfIZzdHhbl/rr6jAw1PepnRvtS0elZU4khIzv/u
UuGf7gcWSpVrEgd/H/n3bzjystvv6BQjUoDSRZJ0MDYkwAgpwwR535Jnet22k02H45WHVUEHO7Io
yS4yIHpK23KMtP6p2rEUD0cemPbyiGkej7VO1J06AHLAa2wrwDGDeqz+cZIQRqOTag0z2J6OEwOK
wrRXUmO43rIYgVD7Mm7ynJHLFEsQ/BzmmmAyCZw7EfRthsBeynB+fL6mC1hDtVJRdVkPjXwqWklU
5tWbP56ms/UGniB3dLgNx1YCrCk4xmdjWJ+3rI9n4sWpsZmxPJF92jgcmNzgA/zqSprjpxI/QsYa
syLUfgIJ19I3ZlU7AsB9OSNW4jDI5Ok9vypQHLJgp6Uvn7gRdmvSWVX2cg2ci0YsfFLjS7UMA/q5
g4m+BbujyZE1XT5aq3Zslc6YRJ4pYsi/jRvr1vv4GI+BizYcXTEJV9yIgwPUzKo+aFFfIfkXP4/z
/7BIN1bOwONj3JhqhWcyihCZHXTHepCalH0ensobjzRhODSMIYLAiUpZve9tdtrWDQ8gKfXZ08BF
gcfGr+5uoOxcC10zxFl3Bh0N9H3N0V1gPHEk1Ya2G4zDDtWtgOKplbZuEc03TwxqvjAJgTvKXv40
hz8ANtm0OANCCV2m4mwgWNBYPxV7QJosXbRaLlo7gcw9WKrv3U4AcWbBAU5hh7QkH4IfAQ6RT4GP
gsKpz4LeSSuApStUr35ItbwidzcFcDq68yFGTUZQtTSkwuykDeT3H6hFBnOd7B6b5ZFEJHqV/U5B
rZBo88PTWg7rrIJYkm0ekrdMepbYRatYr8I6xRbQloJowjiKVFKTqWVahWunFQNSzg8MBmYxL0Q3
+DhqY7DxQbpqwc8O5XlalUrM1EF3yUfRaFeiRcMWZE2jj8M709P7uS6NY2ADIdTO+7PxrDTZe3Qe
w9DAkFQUKWq4xjHRe00z/ZekGlQrRRG7pp3Q/2BDayMbKdKs2ozn4gUFtIwbBgBuTdPSBvUfXGo3
iMckLh2YVA9pXoEKldAwid4OpANOsLfb2qh8JWYFzQltsYiorFjp+Ls89lY/ztdMnhmYNjQv6lAn
BnZvb99pw9J3YOaq0tCu3FJ+tQiv7DD269RE6D5zxzOn9m0IzgqOLf9cZjJLHqRP7xEMs07rRvJO
Mrm7LK1HOVxJm0Vy/3KUNmZLkHVE/D+zFFLYRFQHuy6Otkk/6TD8ZAIR105XwoyidJ+HUdHSn/q4
i1fx432xEqdSZZBMX0syDinBY3q5ycHXciLUpKEZTm9m0HHOY7+aRVSknzGhz+hIWL41XzasttKL
L+DTFuGN5Sicbhtp6vM2WSn16caecMWJTmMRTRsFrYT+M6VoXHwnLeRN4a0wgytx7gjw9lHLeGvB
gjYKctXm068R4j3WxYgXQKYA6zWAW2vHH2cFU3qZ1GH3fa1g94mdBDfo5q0mC9PQVomTlOn0XAIY
kIiqepQuNiK1d71kxrEnXVcVVjIwuahgLAymKqVexHN5WpZxnOxgdWiRQzZW0GdJHm0fXyiphccC
EpIobNeWbHgQE1hAC2HTS5Juqd2MLHl2Rtv+lvNjsE0Ueb5i9uWR49jR/sGRz9rbDIWDx+y4W96W
r+KiJOW5HLDcYxGAb2ruyoHKilzqNuECTwGq5LMH8Py3jZf088FhcsszlMgcCct2tXflbpzj3hqn
Eb8fJPpoHsBvp9EeGDQ/awMASwBambkOItKHM6uxkrjDFyiHNQ0v54NIvBNMdNGyTyI9eMAk9K/m
YCJU/r1AyDSKN+iaLmvBtQgMra71cfSJe1YA9kwwMZttmwB17JmpTHJvAXrdTU/dXSZQwjb/EbvR
QcvOjLIUcZyrCDNBw1F1XKWwhkpRXy6io0IqxocO5ujIW0l4JchaIOkd4QmS5G9llEzNM4eANzL7
EjQI+SXULuGhIHgXmkHzcyk2mcm4tYH910eyVVW46VY4LJ9s6BMTGDcGAWq5Vd2O9A297oDf9L1P
O+I+woWv/25bua9OGK638p+v78H7CX2ak6fxjtx4egMSCcruMlymkcp4CVdGC9AuYMxMxkpnMEK1
YHWl9vfdkxI02dG5Y+ccLdyPGTrjCwadTZ5XwgKbqeCQBD2oRskt6mmmG5A7RfUO+7YXxLS8M6X4
66SG6nu3WcIWJ88aFuFPdqNxKuYtiNwvUr/YE+HDhsuwTFbNa6vidK0w4FqIvdyVZOCkUaYND++4
YnNiwqCARbLVscfD7YQtvcZUlXQmyK9AnNXGbD/UUk9DraJY+6sAch7kREQ497MCgEljmEgv6b6s
Mph2ju2uK2KpihyzFNnthK1sH/g6MU2wuVU2XnZa5RZZUC5m9FkXa+qjBF16DQkCC/O0aNt19RpY
M8ukz2MDV1FxPJQyLSMBnq/LS1LsEYAJrpwfXx9NGwmEBnPAdOJ3rtLHKZDvcEqDp7b3bfHkJy9E
ZqVzypusIZXIVWd7cigY25ohzSqqrA6NXD37Lq7ra8PaTPmoIQFu3eNDqOvAGYO+mvcbgjT54kbv
8STmEC7osrZVdRJ+aF2SraWu5bp7CGOuADYVbG0sSBPmzew58ltHjQykRMuLEbX/yk4wim5S0XnP
QR3gQSYj4fQdXK55tRG5JCqd0ZJoMmCp+CmsPO1C+Gqdvib6ASbRJiq6uHQ+7sEYnc5CtM+yHUTU
nTgSTPCmuNm4mlqxLVpFsSBByKJgbjF7OgB+ROhHASh3gSGMXJgFHXHUznNLtCx1FzN/mJ8ySg5b
ztOfXy0T0z6yzzz2F7SXcMDwKYzrhp9xGDX4WJ+l+bCBmsZtn6S0acoywNlN6jzJcyC70xc08H+i
EsuCgUW1q6gUklsR0XNS1TiJne/s2f9TOhish9QIzLuH61aHYLTxwFNr0ARJgVTPzozOb+yE0MG+
UAYTDwUlwc571F3/HAASDu+lLsFxIOd76q1/jzs9hpwI0/IRBfxtZbfoS7BO6VuEihcqQs9cspwq
y+xBATgoN0McGTAAQb8pQHNnE/Bs/GPlvhX07/cSfRdEQ84m7rdRIIeb2ZxtdT7p3Uf3LwJ28grk
t4NlWzIf14TydkGwqdYNxuYhFd5XJRNNFlYmiEfJ4bGxdBZUNbrsb4I7E7wVNUvaIXvrInvSvtFX
z28WtaBXfZ9g32lvKyaz7aPw6oTNCT6h5wuFYDsr3TBh21xOMJBDX/AQ78c5gzUfw75Ll4pZ2DTh
NooSkB3yUDWpqmCVxmQ0Kq9GMDlp1uRVx4/V9ZcWjUcF9NnejKD6KayiMY0DW0RbDYoXx15qvfoM
cW8Fp5cu4RuvMcE/9HHjuYWlTtyliTIKFltNqaBusq2W5KZlJihPJS48B2FQmW3DNupaGh61dxg6
TDoPub0CdFXX1FrDQ005JwJyL+4TTyqLTGxRjswqXtJr0Y2hkWDk6GNouIs3XBmdx5TwG+2Z6umh
7s3zr1R0jPmrEB3CqmX8Awub93RUoNTEMdD9H2GFSt0kKEZSpJsFm861lv32WFJ+t7LkJOxK3fdx
xcVo/bZJZZG3vk/jav5NkieFP7+9y1uaY+u11KszSi5wvZ5CaRclZ0Tc5Np/la9jGHf+Sx/FtBu3
LFpG5P4fk96FSx7zzu1xyEgqPo3LbVHwfLav897ilV1KkDQQ8p0MBp1GlhmD0BgEdGQDq2Rci+21
AoTh7kIdhg4I0oWcCCtrwXcOjOZjYZYT878LkRNY4yQJGnWN8++12FF2hw23f9GOQwFiWn/q2F20
U8TTQQve5OhQ4vinqQDPHe9O2xDBHJm845w1j4XUYfbzqZUGFpNvaVGXrL4ZOkQoQM6rkvbxv9wM
0S2ew9EJ8Hwnhm4/nAcWkDN9IQATxLPjgOcXH07OkWH+fcrXdoW6cBSKOJsA4qpNyQQdubvnlwGd
VpAfNZqoN3W5//c58nFuEl2LAF3XroihjTVegnz0TnD2fSkP6eIuxJwLU8xjdzZivetmh3RM3MtA
R2jMqA/QA6rTRsK/bfFpeqIFwexjTo429sAL2wPT7Sn9aJ4ACPoc2d+JGjViQP0/dXas8jM0SZfu
RL1EruT4FCa1YmX7nNzk2CxX+Q6hBNIC4nwYiifa3sas3CH6wTiDz1pBzmc8CVU/eNzBRaO+C72K
cvO/5Sn884kGPUdyacRuxKQAYa3I37nzVI5SGyHHIJv1H3Z/eltnjF+oBfrhZBd6xCL2gI7r35L2
aSAMlfX+uiDTA8T02UzI25leONeXLDqu8EhGXpY8CVeBSw6FSv3R0FJXx56qXpuuzJiR+Xl5+wjB
DNE172nGiZOVn0W2sgpg2NXSOlz14QK4qOD43JKy5hLypx+38GhX6EMDtY6t39SpsWxymJRruGas
Nhgorm4MfL4v6BeToXjLdQer7Q/k58+no1EqvNtUcxq/tK/CrxSjtgLbBoKSfFjbMiMMzvf/IIvi
6i5iSnbKZOgGS4CwtmkKx6HxdeF4bSVM1wEP4mukMH76XrtRMVvP8KhKfl3PsfcNenjVCiWNkesw
oCGcga1ZQWd9y4gAv53y2yARi7u+jjuyQillTdNv0h9Kn6bcdmW/2RE2zBDIJAWnutzNEhXlisvM
EL2uOJOfjfdtJVqejCCo4Vq024hMpFjzVpp2TpG8ahi4HWpW2gG8MR/x+bBLFsseCCXlXX+Y08ad
FJa2xwdmaIcOPfWTNwydUEtb260JdnrL/7+RT3o6CHubpon/f5xM7cBdLB5MSw0Mk+56szk90lc6
mR4C0Hj/nvH40a8ZAvQ4wWJ1kRr38S5EzUkVWsb7cMksV6gwDUqePPjv05PmibOT/uELTSQwkAHo
F4tjpLL51JaZqSo6oDiAs2WNHuHeFFHvGUJxusB9yThKj/84vpmgXBJVCVXERwoRxMACOfdiYSES
zzXTFSpuARW7vliGuX4htTZz+hpqHmDRWqp8svv3mKGpm+YJ0Gw18XN6yanug9zYjpTeKXi4gbyM
fwc6UWYPBq6qQU8xtop+avBw/qzv6ThVsCPEz0UW0GnX8tCAIMt7h+Mnxxu3IKvkiMr9nyrc/aXl
oNrT0LM8q31XKe5pSKnsRLANN3Ro1cRjbgGdhIECVJkKXqKUOrRrFCXFFHsTU5v11a9MbtEPKAh9
TIidkjDE9xW1O17CZDrVzNk3V/qdkHYieaDrJFgvEBtrDq45C8Pw+U659JQq8fXfXFSpdylLe8Bi
ZmuVfR4nr1uG5PHreSSd2TdwFLW9grviayhZnfmbntwTTL9Q7XYeDluym6DNlzwgEGiCxlkMfAOr
5Bh2HLVe01QQEC+btafSq21OUFrnahTiHEN70Ih7iALdI8R6viopmNx4DYEdkKMj35iP9m/e8j+X
6ShCWWO1cp691iFlZJi4qgKXeY6AbYebAt/SF8WGsx+NSZVMVoLGp5mNcowJTdRleAnnuKbBoesA
M14ro/BSDOA2d5kj/1Bq2Q+ppcqYeiItYfXXfFho2EFsl98Gc0deaMmXsGyoDbZbntH112X5YCTH
LbiVivFvJFvI4B0R+9Vui220i590cYBxfRMS3iw1sExV5r4X9uJEKKIkYJ9OJILNbBNwGmax878L
lxCtWoCmvf41asnJcU6R1VHjU0UMxOxmtGaj67j5yPolwPIZOFmf/EKz5aZ5TnMbGoEe+KOhrvXT
LATTuWRtvxkZ+EWZdQHwEMAj/Aeo01LVDGYZeRLM3hevnorBchujoY8MwzPFw5UQKytGnquu/mSH
arjCRjgmtoc0k24havPyNrpgxWV1ayAjEBsHUciPSnWSdBilhIu+PWXp0+WyamWERbWpsNiusu1G
kGqC4FOGJBLIRYL2OEYlaRnekeU0vRF8T44c7u6qAY5tVu2svTh5GgrkkQoxE33L7nf04m0A0XwA
f6DbP656FUlkXcHy6Em1ChHdE0etZprFaTgXnb5dcAShn9iFS9/ifY7KUN1xD/0vm0AtdETTbE8r
Yvo0Q4/O8fhy5FtF97B/Q+JhHOtudkMzSxU9wFQvcAGW4sHMDvXvMrcssInF8jx7XrAjhBu9x2TM
h5p7D54jMcU+s/UfgIL3NIjxP1NDJZ5KZhZ0u8pRxAz+xs8deDYjgQqOVa+51A50y7T05j33uwSY
3uiIgolfV9i8QdB4WhDRYhzX3luMlAxqXeg/FkKhUYks8NoxiIBZvzDs3C6NWzaI4d8aAJplmAp9
cbE7RjfreswqHWYby2rkBZr16LxodxqYyE4ElLmaoioKjhXIj8gg70ia1ycF4UDy/BbAmRmHbUXL
50JqSH0HBuewVpdkTH6X8jxrkhQ3qNUBM52lPbIYSFJ+fQT942e/mxA3+cpgTL4oHWQb5dvsaJp5
BedZUJaKU1eGo3by3kDagwBk30Gr1a8f9gps4UpBC4iEg7r2M3Ja7gQxxYPS5JysPQqfGAEfPcLG
gh9abrgLp2WK7JQ2P+D53Mu2s73cizGqQ9/8OTF6dFg7Tb3xBOsSuyH+jgj6y24Zg2cf++Ir/cnH
d93UGaYk7KrXuYz2viVxje8HtEaQt9WIObE7COlzqADHiIkB+qvRo2jNTF4QNAmPqdul4jO9jdOu
V12mi67gYYDHg/T3arJTEJzYxyaAz6MMYqrfFgMVoTh/qirRINAXsdOb5zLLtvpjIpfu3alLI3TO
FHYNBGyO4r2maZKUlhzF60icaolJ2aezYT+0L3BFxXbkk2/N/+E/kg4Acz4YNljOaTuvm4nY2T93
uQBkf0TyyLsqPJlpeeRwW8WHXuYOUo9KKdMhSRvZf+VGKa3rJSOHXrWhoyUMVJhssBdwiyK9C6ci
QFpPqGAzFe6tvNZlZI0RiHAr4DuMmpJtUgiJO7OkvgmoSTuD1Ay9rH4pFyCL/kFNp3AbY04jgFlL
TgU5aYXJmB5qZlio26fMnX6/VjsMRWb8o0/LHgiRkvmGGqEkowO2bCWZoXScPSh6rb5evICqoarB
xvqZElJ3Hzv/cEeZ4NEetU8nFKCj9DiB9JiNKF+UHrWltV7C0PIwFQfnCnaBqwQPec3y5LHPdtTj
EX+nTPMxXewE7+kBwyZP7nMIi/19L8Ax1+z0Se9lcibKoRMfskpQhRePX9K0fwfoYzR42VCRW/bm
rehe6SDb2G4mLOdlg9Frf4eb2NuT4Q2WL05rs4RFNPdkByifKZ5a8uAlhLJbzyU0OGmJc4tyePVB
yeFWrq46vILJul8DAH7Pt78N9romxOKPZDiyYUuK0IZrWWNhgRRXN89cF6DZkg5FOe4f7t8s8xT5
tKJs3fes13e9cQqQmpos8eYcWcHVn8uD4PXF+9zIb2ZVELIaGx8kBz11Y9DbTqUBXAEg1EDKWfH7
BATr0IFVrhA7qGitnHbI+21STJMIbVlyrfb5siG7n4DR1HkwH3V3ayc294Da2V6iD2RFy1jyzYd7
egbA5i9/DMkeMFYySLrr5FVD94beO6o9piVgLyHe+PXRO0lrOWp7GTDM/JIDooit3Z3NNlqFQIIa
WsgC2zoudEHhQR53OiSOdZsuy9w4BhTZGAcwyqjctEucMSA/+C47FUPsb0ADyRar+buAagZPxgAE
OcKN1FPjVIBVQl6Rr/NOmJyOGf6/P1JNuLzj9B8LBHXGxpe6gHRQUrJnfQn/47ikf7APJf13v9m6
LykBzq6ESadAtAWV/4zyaEP36FOYuHbCNnzozzPGfM5hzAtCnjQuLjpRufFBnGeV142ihQlLulGI
+YNrRXIf7D7Yh5YtEfNvGUQa2VSOYNqe2kwHeE9R5Qc00qf/MK4AYko2FN8vkdV1AVHIyhkawGOm
zFLM8QY5O9zocMTP2ixtuVy+LP3iIkengXHpK6JMF0djAKhssr7C5OhZ7wZR+pixUVhPD7HD7R6Y
ryb/472uWRrFXh/8AlZeZDAEBstFPV9R2fBN3MZquceNaFJRJBBrqz9Ls3QjXyZjCbD1gIDOv4Cj
jogkrhI0i5Lt31XTaCYmDs1BkUDABGTVYym5gQEv+AxYSDFZQWPL5yyCtRA6tW7sk/X0rdm/TS1o
/7x5W3+8U7B6wJEeDEXZMKmN8ZF1sSXswCfgstFiA4u/E4C2MdIoEmC3fgMterskrZespph8O6Tr
s+Y1EKoW/OU7Gw8WtREnOPXZD1kHUT8iTf59wh7GSqaBl0c1cQcW8clLIBXZ5PceacUBdeWbo0YZ
yS0w6//G9hi8QIAuH6R9yhOy5Rzx+QAMNWWbvds8/XFLbiu6AAGD9S52B+Fkj2PUKa0nwnlOaWrL
Vo00X5GDr0nxefd6+KmdeAQJf0pjQktoyQ3+/yU/L2NfQNtMEgskekAgvg4GHw/158at0O3A51nK
6AHuHqk3YWAChd/s8v/OZT0oxZtQor6Tm5ORHbr6ar9wIZgpZHz477UEqHzCxZXYwXFPZ66v/f3L
8YdiwZUfGVpAHlLKzWTk02gETJ+4F88Uok1+FyyWcHqcGh1O+zGhM+C6R+x1RDZzsmVGVV7HTZMg
Bz6OV2Nfpg6jSIO68SEnSWo3JcS8JndDB7z/NIyzaXYBIQrLG2kOiGrIC+uz+W8FD/1wqoH6ACvL
T47qvpwR7T7kBfH4jChA4CY1VNCdB66jgYxBe8s0+7b+cXeUYdYjlG6s4LQRsgBiMorNAH8tRUrU
xNrAzOXLZRryO++blys433NsLGoiHcNpJjSfZWXqdnEYJBuhLAR7B+YGJMQlyDjJsEGW8j6mpqcy
5ThJxo9NMtmHGcQ7NGFWuGQY0NpSGAMr9JTAdPyDfDmDWpwyrjtCTR5YVNVyWoGNkWwb/LN/dLdA
QMe1fUTYmStZk03XJ1FemRwHNLp3Bm9lSp99T6E2IgvjpiEV+l2EJ17KZ4fj6HRbA60pyEm8P96h
yySHXcR1sHcCKO2Uys/CppCgVqYdX38zlIYC4JZrhOJlGYag35r7NNrkbwi8nE/jKzVZhRZkW6pn
0/c/2Lilo1gr8itWLGGUW2Z5PThJGrkiNNhy8PSlwTDGa94d6iaBxC4Dp0aNWT5iVR/zQOu5xM67
ERSsJFzv6OxBDyN+TOra2mxGSSLjbP2kmOVGSw6yG1LRjDAAjeNil0lawmgjDpYJXT7Ahe7D2qsY
r9ZgCKcj3cS5+mleoWACEpZzSs3bhpWU0nBg10YYCDizXtz0wiknEsJTVEl6oqhoNeOz0B6svhIV
5supuE+7tiCt6tD30lw9aHfGqmGENKDdXvJG8DqBaceenyT5f06Aucnxt8XYQFVMRgKgQh6fMcZ6
y02pPuaRYQYYt9LtlJL+SCn+CfGcXhoZeZ1krtLtfNKMNM/6bSeBq+1VqhWhnfbZqEqNkGI089p/
EEk6x+LTW0DGK1V5CngLKFfxLLnk8mj8mPc+nGmQXVocsF2dU2kSJBVRkoy75GP7/gINuOfE9tAy
8CR4Y2RVeB+29NcwdgV92gzq7ZyPzsz97YcNaqMFa+5q+gnudS3N0UPcoB+Aizhk2pO3aSDSHRGm
8nVr6Hig9SZ0/4uhXXSn3rccf074ZwCKthF7os94BW5Uw2pa2Yct3fWmq4Alq1Dowewqj8MZzl/k
ROTzoGZkVy9RFTzMEmhDWdkSgkVATAapSI6JUF+t6t2nYNTgaARy9WuopeD0SsuPnEk5rVIQqsCM
qTIZJzLW0ScuGYXS+sDXVTGb857Rlpnr/uyoYtT/XlPAbB2XKdroOJfMU4czxPAVguru5iCJaOCp
VFZS7sH6xlnmIQ9dNxtZPoK5cw+jJDvpggLR+c3toINOdASzeH/FFGvah8nhR3Pb1b+AGiKWuhap
dY6QZ81jBdMgi3Rs/1jSNN8ulgvUCF5meG2/7fWH6ZFIXrQv18sWZG4sve6fmibveSRkaASvxEqi
devPHTyuAPVJfCVw22S2gFgLMGRAUn9J61jCj4vIyU9MKdth16i/zk1lQOEhysppvkrQnK/Fa+9G
YnW6luop6qWDodoIBSz2OqDVAWH2WyOLdqxtzIzVHOm7ghQSNfHuMAz9kkva0TLPLZCJzaXf4Nxv
1S6t1Ha52b/jRCglXpvpWfowtpn7n+b2EWNN5VuYqWd0VkVnWbvMXwFdgyEMS73ymGq2hpuQ+FKR
t6R1gvP+XTmWoEkixH+2dIVyvpzWoKMiUScZDnoDeb+nXizLYGZoVlDU47kcDNG0oZR/D12i2u9M
ps15hnxMkKtcAVm+SWsGM2Mkvv1oitft4HwMiIHgBGmofxGy1Hw+20c4LUomKg0Ec3Z4R1dPt6fK
7G4oNHzMeDDyjUTZ5HWmbgG2c0vnBq9wppzwMI7eaUazihf45DU3frj97cSk6pUWp6z23FwyW2qm
/JDVOOS6zaSJJ5Vmv3iqx4t29A4vEHblQ2HM38LXWfLsJIxb1aMO/tlH3bm4+Qeb9zl9CYtjFkNF
L186sSAgDUy7qaczRXE8CTJeSyMMXc6z8im9p+DClRLaA3dHFo0vAj7pqC4pgTod3osNzOMFgkJi
gcN3FPl1VJ1JfJtQ8I6ZHaXTTgRzffCtDzSaSzUTOYtaT/bmDf5enOpuuS2VW7aj75isNhRa3MhQ
S7tP9fXRoTYj758S9hRMLCgoeQer3VWNN4j/JYw4OE4MzpUXA6Qa7Vc2m+q/+9HuvGHI9FIfJ5AK
5e1UE3RRilQ/6GyngjuFqBIzNHsQJxV9NQblfBlfNsYnxJqIWMGXjNd34ll9g6VGsq9/eri2abp4
b37g5bDl4ZnStiQvUGYhYrsQ6Fww9ZhP9n9Qfd8T8bFm4DLBphb6XZjkabtHE3aSHMf24KE7itBr
k1LWypeF4c/b5eWStuB7HSXVo/fkKyHa7oI/jqNqe9/YD9hwDV1ioGFT3m/GVxiEFGLzvK5aQLtC
a4rL4DVJVs5YGMumDRhNUk9Ktg6e+hIqw5xw/2sGc5EHV1b4Qze+pmAQHD7CdqNW7Gtle+OuAQ8z
s4jLmKNjYPDA5M9fGGe6RALK1DlFvuWa6hJzEB86am4ff27S9FBUIvLiUMhNEaGlQWnpG24ipUcZ
tGgmd7ipQNuwRi2UopUDMlryq3x4Tjn3T1uTSFVUjSCOnIiMDaLpmDXXkmsiSinvX49/pmD3XrLr
BP5p+AvxOkkS3VraKTVYXCfmZQik8bwFy3b78rXyBh9zT3Ez/6MJ+bOCFw6g8ZttMppilpNu0UvC
sY+hqyEFHjnDVv1RfBOcB3tuSI3GpdKuI+GzkLeRmUniIBryTKVPw3iPM5As+KfFLSgD8Z10B6eh
6njdjVIH0jpMFOLPuzRZQPgvcYxH9ui6y/Z1RNyc2oJtyTuxSc1UINXprrKDGhEq5hoZ9rQUslMW
P3x5CtdzhV9iXtiYdQDbmQw2XWULUda9DttraWb4yRH3KEVkzot1v5Aqm3gDVez8jIUCjpNxRLb0
1c0CUGu3WhOwLfu++c9Jphn8uuFQ7yTgj3uLtrslY5bls8xp9zxqfZYxbi5KxahytcGEhH+ehB38
OHRBiSTag/PheGeH64nysJe40gcGH79bXznvQtxazivycxeIFvPMBPW7+3oOx9f+O4TRj+trPMDJ
V/BLSsoNl4WyY02xpK8PHsuHAIF21puiATHqimb2h77/HF/ucXfaEPALoOmK4Gag+9h7ySkirHe3
sMukWaHKhZfsXkaPTY1W9RvWLE6A9HEGZi6+VwD0exI5ED1EBAX+rhUhv/34BtHabdDyKxrYQ21n
l7+OSS4/bEJYzd3Tm4io0oDeMt7inCXPGyrL9YrRV66NomDbXNNkuub/fpnqLMLzokQDOdH6WvUj
Br3rl1O9glOkBNgT+KoAaRU9f6/nuWw/dFOMDYJU3CPY0QJEsS++FYR8gIah9rUMu7pp7Y2uK7Gr
83DSWxA5ax3NXrTw21Vsxnr4uxJuyNoFIXvRcoJCDGKAmM3gwdNfqgJH1v29fyqdW864rzzSceNX
iXcg645lldfvtp7MgRJDwQmAf3dURjpblAGwnUctXhQ1UI+SQJvyGbLhOEiho2FRamO2/sBTCV0w
CzNgrnUQP0vD4wLgYEhwDW0JwP7LDVrCV3v0vUtzf7I04y0ZQMHisPPUux6KrDy0JbDnkN/Nttfv
I0UbTbxsQzmKPknq5Ex7/5sx7Y6WRwZsLtz/ckdAzXs4EMEhmEsSsxxePm8D0oDpulCW/s0Q/kI4
KfE0LiQobX311/iN8YvMNZ1d0kDgbriD6oHFluIUhT5GUjuQqlDF/G/RMD34tDF2rt10S/R7SfYo
E3h1dKNMzL1Fuk2SFlPoRY3pIgQ8qlREf1lZ8A5zKzAhVlHOxRZgzC9VCnRbf2j7m5R9fh/2UIwL
ZaPzHnY/wDkID8IVA4LYUoVaf33+IlRHm74SAHX9/AeowbWRGXGJjskfuHwjNTbZJM96zTRKUd+d
eerrkZ+i4ld2HtQ3NW4piwRAIr7CyjdXCQvGNz7PrMVsOnX5YdD5EWmkzFhPopHS3sVXdUVSdGKj
RBl6pwpDZXm67BqzZQZaBLX9cikDS8GuZs/ta1spP3C8j9NvqNlRjHdp5W82OXjPfYE3rk2kZJtR
yILWgW5gU2cPg2zq530FuZpReCZlhU+QlNK4GBheWw+rXh6mBo+SMioG4OFkvc6UwlT0xLgZ7LCE
zXKkS7/krP1QfLryq4QN2bbQ1+UX7smQtZ+Nro5ac0knCTL1Nbq5JTSOce6m2r+78ONBNqkD91qS
a7Y+b3wctruTwcYVGQAhkONH0P2cPl2DTR9zfNP/j4JPFxriAgQT4NfOrQG3kQHiL6Nnp93Ttelh
2SjikIOyUhUhWrNSqJw9069pSyHPqSIxSvIVd4RXNsG7O9CinSaCI+BUKWmC3RhE4r+JEMg1uZxQ
D1CFk5As70R6fikRmRiy0v9rpaS+h1s/PF52Ssm5pmXqnh9VEIn1ibOQtDuMMPhOa4lPbcuu3ewC
Zaluce+ktarRN8gKoAxcJUrSZqc/NckiFA3QeyaGJpHSwmb4AfBrFY3qeoi+HzBonXJ1txh9SzTI
HIoini8xpMbCtdWEYL7i8XPPItKLoZSHebTJMws47Zo/9VCDqZXUsJ6JoJVfdQMBtSIbbzCDBZLZ
Xb8IxOXSKzAATA+3Ndka1+ApaAaGIq8/lYFG3og6whAaO5H2DHQgN3RC0ryLqbeSxW30bMSBUHqq
wtGndpTWfwg6LpawMG7IEYHZQwg6hDrfzxsf9bOIn0wxOrGk9RZ+g/Ub5x0JgJ5bG2sPBnlvGQu5
6JSFt5Mi+GPbOfsZMJV27sGT9IjauFuCla/yxmS7AUFq+OL4+cEK6G+0DZwBZfyABvQcLgK5w3IG
xzza/qS+UucaVEUfjwzLbqMprnaDEiYGYZdovP4AKBUqU66wAd7/ojx1pNZCMd7rFT9g9R3FEGzY
h5CSSKq0ZHicn9iw/Y1nn2jqYBvddHHiCyGq0LKMyY6gY4HnZKWLIWCU6h5FnBou7Nhk7RZ3RRkN
YnSsUhU0g+sceVflcBRVLi5sYKBQ3MxaeKTDuvq7I2KO+JATbEUw/NKFrRiEFNFsipwnY8c+RRJX
mSrTQ7zk+B7Gsys1tOXI/e+l0pRhASikXpa9nOdXtli0AVM+GU43Tv87DqZG86ftI0PVEK/at7RH
ZrZU/uYi1h8dC1V+on92NDyy1Aib6W7PyMH+00isk6kf1E074RW5P+3vGVzLGisTR2xYxVX/r03Y
C+ps/CvuWZOIGEJcKnN+NgeGAlU4wWYn1tB4zN6EVBCpjZhY3eMly4JZ4YujFRIzLhZVyq5F2Crn
WldiddOKBOFPVgWxAXb4Xras7SDDVPDTVGZEsNZW2USMwlIO3Y0t0vz0O61DI9qoQ6znHigJpO10
j5Sas7UOBfB1iDN4Osd7C8PPyADQnIKx4JQGvp+zwHk1AYgQcq9Vk2WqX1HjFdXPD8VbGaeXrsBb
7i7CifFdxRGDZBIPhD/OSJvJX0eX/gJ+3wbq73S9HCurUZiuQwr3lEjREP6IXn5+h5JHvRWGM/L2
CDGQIW8HHK4QV9h+/h/a/P9GXfWgXLOS/dxOTh9gzQNPFosobsBrn1bghW8t5o/xFPLfY7tfrkiT
9Zz7TcNkG8rnZLg+JS6vCVnNG/cGnQvPSOC2IW9dJyUtbf7DssETG7phwIWBaN65PAXuukMjMr+a
eqp1NmnlmB0079KCOwt60fUX5YmnkRnUCMwu2tbvNFoGcNgiNalrwzyEngRIUk58B02yEwVox4Jl
ik3crQ8AwSlyEkYvEN85TezcfEruln7Bxre4pa1VQPNZWAvfLps2WMxOJDjgjJwjFzATEHefqYxU
8CsbucgDz+3e41wZ57A3HBKHiGiihveWkE6aoGz9oPM6cRpKWzBrcw8Fdg9y/F9BE09Zc+0Sm8rj
bCuPGkoVMr5QcMj/kccjQUNd/O4xIJ/ei43agbccpssoa6IuAEOQxVvO7M0xdhZPa05Vds19x5xI
Dm5MXPkdMOlZ8ociFbGQxDk4HMU/hX0kincvZ3ydxcLWMiy6KFVfPLr8leC8SndQuqmhcadJoyc0
zanytF2OyuWvvM5mKNnmPm1axNA6anXlOqwxIJEjr929b9+ofdvPKJrC3vCummU+TmABRaMpHyQ9
Vsq9sp0FT0sOJ9qnsjnbJyjVNyxXslSY6bkPZ74lWbeYw3A5pquQBaDERakP1a9W6tv4WjRuxThe
Jm+o5IFNinMYXIPChBKhr+94/+Pz++7jRYaWxUPYeJTlIIVHoA6/afBXbkQlNpelVMwOyhIPnMT4
f8ewa7C1Rxl0wIGAHj2YjMQBXw2xDPUOc2+5BuwE77J9BYMaAREGjk7K0D7Xw1xjv0N4UPHVKRRC
3hP5v+CZzz8IlpKWjT7lGmMIzAT58Zm/dLNUAzd7zvJMORhWnwIcE6T82iq5NTi0I5jPUx5h4Fca
JiJCHsMACA4CTj+KglSKFDuUPs9FuN9qGdmnUfY0rKvTrYb9xfty2c9oAl0VAy/OJbg16NzMID3V
CYgljVjxlWa/gm7C4Vy42waKwpt8vyus8GzDAM/mn3GHm7E9j3kcHscxFw9A+L8n8MdKU+tnoz8D
r73U7q1Cp9HXb78BaaRaLOkYZaD+cTVEJfKVnadWCtQLJMUqg58CEAviBK+pJCNA/I0U264IXDC0
s2dbWHkHgG16xFjV4JpxVIcOZMb+qWi6+Ai4j/YUypM8orUxMG0kvrohLRHAE1itTXwSuZ6JOvL2
bJ1NQ6RhnF0z2P8+7ora4plic/zfP3st5htMX3uF3amYtLwvUKm8FWlFYgQ3VknWEy9d14WMfOib
UdqCveSZNheMzKdFbTS5Yzcl/bmYi6tq+yAbX1SSnNR/uYnGCzr1yuirI9wxdBmxHl3UX0wiBW7h
80ab/rDRRtg29gOQi/AF/Mor4Y2cIxovaIVQPo2b92vc3g5kKYVCb/Wn7/fQmOQ7MrALZ3sAR/f/
tpI1yiLH8kKmFVQQZ1E00SkNFwZm4OQe1JGGf0i/tAIKH6zgvzdkdf2hHMlwgY4sN1zS5fvXEfvN
0kqhZzh8cAiR2AEbNecOEosTTlyLF+GU4evLl7KfauOa1esYzuiKTZMyEWt3zQLxh5q/ZcvVsRcs
xFAaAjvBIVDI/JatDvuOKjJjQt6jzuy9Fj1zllr8Ru2Z57L1yiYg7Zq6u/DwXd7mDwVJWd8elCUp
D5inEeCXLLTZiuhViV8XkgEJmkty0OnWV/dz5ousmr3kY7Yib85AHQiXdxfDAkF5LBBjV9JVhlWM
iz5HUwsbIU5TRvjLY6fSDw9iU6lXh5MuZBX+M4C1TTB6uu/EHq1PzTBwNsztYEMJiUOALDv/h9dJ
CUxQZ7wBBw821LYJUi63RblVI2qP0fjc6NSY0gXsxK5Zmqq0o68YsgfSzJJ9NywFAhcCz/x/h4rT
iEj6IqohQSv3FMAKNiDAonmCz+3QUZIc0qpB1Bfg9fpmWQxNxbPjyq/uFF4Uiq1qvqJM60g/a1x0
Xx200EcIwd5sJUsLCUT5DhapnfeCw2LF8o1sO4mwiO5VisxekJoGAIHfu7mo7xGi/im3clGSNJ+Q
2rPtqtTNVYozrEXPP5NIjdsfU5y9XwbA3LHlaPca9arv/Bne/d4qoBLlNw17ySUk1NZZXxSZ0l0y
yebsmDo1B+VgENTEHC1d6L2VyUEMisFUg3Q+97pKPNyIEGFCOLfUwCi9l6kuH9L+wmz3062SO8T4
p0R6oFoTa3J5No5jZr6gbmY0XNkmQmyqAl2fx401m0D1/iKQeQxNKOr2ZWCzQCzDlhooH7tGZQnH
4a+RKRifp+0W9yv4JCxfyavnD293tDrC2kXdgqBS4DqR38b1EburltFkSoTAjWNA7+Y/JCzrcE5p
yoWeG1f3u/jCmCi9AL5hjfzSsNE1p6DbJfk+iyME/N/GgtdD1su2nwfsSx2282FnTFd68ALb6Lkr
Lf1PzPNpwdD11mKCNVWNO+cJwdtkbCIx2n/hVJV5/ZXJHDrFHHE+sm7by/gZY8qoj5eIeCVvkoZq
EimCVzqYQAUJUD3TR2y3aNyBH3k+Jyl1t47V2GXSo6ocmfhKpxMeppzehsd5iS+wnCmgafpWFE1V
vJPDOERERjgD/DTmovFLHrR5pzgJ/E7Upp+3f1hsf/BQdTquLcYxwb/wIxixcivVtCUi3vM1QKCa
xXzVk9FhQVZiLTUCGdgQT6+x0t58XMfF9REI9PB0V9Pn4PS5yiZgAOSUw+urSVkP89vv7zeqw1Ds
UuHAS3iwKFgRWxydy+EuDFTagV/khOq4keWdMmfmnS0FYdjO3GwfJPtohw00ad2WuuygZjXCTjNU
qxC4oC9W9+z2Obbf9H0fFinM/KMYZ2DUSbR32AjIYeH12TTJNZ19mvThOF1wFdbVgM30eBXcQTtr
8aYFzA5e/GIhyYX3WY9Ke5ht+NEwSEfJQwDvujuAYuGszgQpTgsPwlLgGEzYKSDeH9LNxqul+j7C
8DWpXqt1ME+P1okifwP1ewObmq4hFze419kunr8C8ATmdSOk18tB8h/ceQpNLa9VSna+Z00vxHuy
ZT1IkSBUuT8Yt8rh+xJfD6Jjh/a0ydzn5PEM2rNQBbUumNqfn4ZJ/UpYAbi5ahYlIGqI/Y8yclxU
rjl903q0fX2y8gjjHxpr5r6KMYYD+C/Io4sksyWC+EBK5zcMy1oC+OUgYwiHegWc8CPWriOcfX1P
hQ2NogOniOT8e5ev7GGFCv2HVMDPPe56y+pxJkkBaLYAUtKAVKDkJ3i4fLXzmzfIBK6JWU8RaUWX
2cSRFeJU0SEHX80S9Y6heE5b6B1WJ6f8cFtfG/9r9D1pObWGg614Mo8gq5QoKxyFjd0pHwMP63nj
/bXl5hwBsPbH9ZHVMMdpJikhUqgaU/7M04k3L60R529X4mflOMuhe5hCNMp8pCiIV1kVP9UlNeL9
UWkeFvZ7vmtOhyx0B9LnTD5JCZy2COGYEHQa/QBEkzNce+Zn0I1VGUZ7P+Ed8fLnt6ZD+vhXkOdj
cHaAqtv/2ISrBLEmYEd+SLSx+gOifV0dAwf07QZtiDmGDTrfWkHqEKIUKEP04BWqo3t1JnLapmeU
9w1OQvPTDckNtULVCw+K3HpqGc2wbQjTjjbbXwhc289K4D6lstj1Z/JxNCM0NDajLAJp8sImFDBW
gRywf9Dez3dEZeGR7fN/xgEcywv9EmNvYik9DuJM//XaFHc6jgXavD2F9vJKELg2JC8eO0syco0W
HCAkCd16sSJIs8v+30F0uJt1u7RyU+9g9VgC8DLNNlj18DXJMasRRGjSfRFmR2DmeQehuYLVdoFd
mEBwzEEEuyUf/SzwDI9cFFr0geKCQ0m1K4kCHe8XClJ5PX9wKDewz2FtHyqyUULxG958K5J1ycZW
HQKgwVTTWVnIU+ttxQnZke59i+6mNFRmTuvO9l20YdtDKYIRUk0Xzqu2uK3P86muwqlr838G6orY
hlI4PZavxqqsyM0x4fUPAbpt4taeUF//1DvwZ+3Pq80eFc1shhUYfXR8/tXahbBwGYQegRvjdesa
/hklW+iYAT5Jc61HcjHIvdfXXen0TrrP57EsoaU4WLimnKJ47C6Ssy9G6Aa9IlRfqVQlmLoIMrin
JuyYEHZ3NTgmxoCue6gyYuB+FGRHTC7Hzf55um7THnbrIQDqxZqKlKJcCfKzRe5FwoYk7BPeLMZv
bw2g1Ws4Xd0k7khS7Jnp4PMgBqQe1UOBLyIgQa+xFzNcULx7aGbU30UAZwsj+abRdzj+6WvaXvXj
VTWdkSjwmVQH7QTGM0+j0oRSs9Z/Hd7FQg6SttBEqVXBWuj4JP9EweFLwse7taZPo1geBt9sfhZp
IPoSf6brkIry2hXmK2SARNUWkDb1TkpwHok5ps+aQNJw1JDzjqdBICElfhxdZw0oS4pyxbZ+MqyD
L0NaMbJ2afaCx8FsPyc31y3E67onqxuKIbVgeu8WCj7fsdeXzJdTVhFrvSvTc8s1mGe1q7gGyXzh
GKW77wI8yTWM5dHQSPyjPzykwrVRD5he66jOe5rcrgxxWbIyvrjgx/cANOG+kk8+upC+ALXWsCnZ
uzX09OoFUxQ01/SxbcQN6zuTX2bEYZDB88Roa3YNuE/aDoI8Pl59qkWlP1ZZ7AHZnFgcCw8y6UKF
ExcUhp0dprLF9S4E5DpshFfiIizIxfgsU65t8jJtHdje4mMupH5FAsGdrvwoLOYFKHJHMbbjoiR7
mj5WaSLflg98IqnDVvAr9stzr8n5mspPkXwtCXl24LueWSaFdD6QUYb+EJFBtFbpyhL8cw9EIMl7
hyZiVkYBgl6EBnWmyyf5OsnreR8gX7oLF9e/0DGWOkAlUg1lZfD3lDYqdxNzqwfVRMeLlqOvr60V
iTUkPAhgmgi84NTTSBtY4pBt/WrexSTq6d+6UGKBlj89ovSpRP8OBJlyE/v0y84sJojbq2fyE19J
sx+yRUN1tvaQRmYhmdfk3AgxLLNntRsHRCo0A3F9HO8dEplSvvQJFJ7YhOZwehv0G3lz/VxbqZoP
+FQtSA3aAz5IvRqwCcsDLK1q8lIHezDzJBVEZtV13JT/mpmaqDW+EwpBAiCoouCY2VrG7PEdFHXb
07XGJdD68Me57VLF01uxpxhYL6UK7+01W/M8K62bgtQ5gy9Bt4ZHzMzKT4RbhiLFpHYaEJ6BY0k3
Xz2TjgqHmDebVdWmGGkaAGhRXj/UPyNx98ktQg6WxCdAkUikYSgCYxC57Vw0LzVyLJrBfqiRn8yz
VtpvGz/c67U0MW9/JCuqLu4qh3iPSSaPE2DILfzJv/0oJvIMsJG2NpWP+pXEHIdyATfPfpFNbTnL
xEZEjX1apGPti768YN+CwbF7RH66O2gPSubbYl3lClRHnmE6Q32DzMNkcoxeBLxqfekZEyl2PYyl
mqqcQJJ/AEEYNQuu2MQTxru95udc5lxnPWqYGLwkoK6F8ls/QygK42M/VAeMgmlPqHS0yfQkn3Bb
GRtNgW++DIDSiOiulwHN8/VLkqClGE250pS9Hzmm9ph8qORChHHjYWMxuka3rHQKf60nZW9RLsU4
H/QPlNGOvyi/oHPn+8xoX8V4kkg7mz7nkGjK3ymre6bxIXnkoI+GdWbcR4nXO050nhblXil2nV42
YE2vUp7nGUg8zBfa5LQck9Ecic4brWM+T1m0+m9ML2yH9H1DM+SvgY/CVzoN1f4+fYn1W7TpH++1
pQ6TDhEGSQFgFXTD1uJ099zKGzxQxrfGAsXl91oQttM/XtowaQS3kW9M4rGY8J9ce3exKH9o1C7o
CuJBYrrLfW/tIoB2PLmRQMVBUwBwHis1LI5ssvksbX9HF+AA28MmM+7fjKuJOs4H98Aq/xqAekFx
MYfM/KubP+xOHVI4WD6F+sdYluI70EPuGjrZegL5/3uNJ0kSjvcJ6uCMl47rtsQ8UmNpZZWIpgbw
bPg2fDVGoEvdfz3wGEP8UuHYphXShK6izHfsYgd6/iS1/On+iCq1EMe0sOWopg5sZg2zLWEvHWrz
8a8lBOckVXcUhX5yUb7YGwKdaxGFdYSfvWr6t2pz81dmQXsw96RkBPmiXCupCanPeoS5lmWULcz5
wjhsIbY1JXFM5/aiLla8gcyOXv/x11q9c1OottPCOigVh1FFsSADhsAqpYKR15CZu5njok1khn0u
kXMofu8NgipaxaZqASftQ0uX5ekspv3YQMOF7HCdjUdUgAFVk4OP1OBONIzwiq7vmmtErzeB0TRN
juhrFru8UOXeVyKJHnv99ixbThV2iUUTeEmQfiipmT2VC2FkvRK58wx+0V9OYXl/n2+MIjnLm9qg
1RVy9O7E6Ma1TLStkPzEO0IhvXUALtc637BTgtPN+JrnayeruTuLHHj4vONTfUF/cl/y5xx+f2Ha
JPG2E5CnZPFE9+3QmX/Mls9rxvz7x9fOaZcROhZcrzEv7EGKFmx72KXWoTEqMLNs4H5vq1V9fs7v
eNx4rLVgtqIHGVt+n3Q/7KD7/XmtMsECd2I992BL6z2G1Nuziv2/jvHulOuGll5UuzAWOyP8mWqA
xciStQB98Y+H7jGhQ2UJHayexv8GZAEgk60jwEWcp1EogGol7kB4QqtZ94T3P4ULEEVaF8EtVwH7
yxeMOqoTy4tdlkPEkj5711RurcM9bJlFmJ8pMVkEvEZyWdLLeEsDy10jR0FICiz0qf+85IHyTEWH
YcmTU+wda19VOaUsdAGWS6FTVl3ZxUO5SvEZMlYVH2NyQglW8WGL8PrCTZ/O3dYlykbsb35Jk+yY
2DKbxhOEzP1Rb0UZOR0GmI9V1naBCrsK6X2kMxlSTB6fEFlkamHRrNMhWOB+Z4xmj9Oyw4gr6Mze
CY2Er/MoSoCxicqHBWl5ITfDRD6RP2l5uq1Z99iKr9EyzJ1R1LNIgdHscjTyS5fl09cl0UE4vf90
xxN8vFis9j7ShRICTSgYd/pc2dHXPa4yOBrfnFZmG+EFrrwaCVKjwpRgwNrtI30MmjKA7cL64FBK
L1MkbGBi4TTSD5hLuIk174mPp619UONclA5Xfbfr0graqzvkAL7Y3E5K8HO2zPQ4CfmVbwoWvRTT
YMfXcwIUNjCuoC4Zb+C6JBQhDMSppJZfrSKSFZaY916xM4cAlJRgN94VdVatFxLJM5ALVMiX+HsA
0MbrjqShWo3exxarYzjK2aTmRh7iH0qpJU4ljekGySANTVYAIFdMyNJab5Eh+uC1iIPU80UJUhVe
mVFsTi5F4ruJeYernKQu1TuMTlD/65NP915V3WtgjXVmKYhF44TS3N09CoLZDg4TQOf3M80msppR
W7PShNQt31gVpp2+xv5zrxEeQ3uHEDb/ctYg8yPdyHpPIkRA9dNDz0sOiOwKq9N2EHYSdU8P4UfH
tqJT44EeDJCVTmqOBosBlyszKVLHx+bA0luQLY3mgugGYLZZt90Lwkm/9TPAXk8pE8xO7mpsJpzq
bmkvU0yHpeIGGYewfJ2iVMsjMmIbF21zm3OEs/a9gvf4VN29ZHnhHp3PfOQXtjZqx02i2NGkldAW
Kpl0M2ipzH5+zG36zPQOxLcGuaPa/JCyCf8meQc0is7gAkGJhp3n3uhS4enFQCXGSeGHpsznmrby
L/iKhJvfLZ4Ia1zoueNaJmokI9gwdVFmsfy52DksKzBmIYmR33zOz1Bf6aLVUpaExnw6lf4OlIg0
WnvxopXH8sP/997Ym403BZjrXe3/qcUNiVNRF83+o5ocjhjID/wBseCIgnxj8QdlCCbJKSQLfPCG
lM6PuEAIYgmmQYtupjsdXRoKzwH8eX+AgOpTtGEfbuBwOst+nOs+We0uYCnQbW9zz1nlwjXIQS9X
ZTN3tTXQp9Jl5/6qKkIP8KaZGmr2kxKC4cWg+JN/S8r/3r5X3YRvJ3GOzbdBWOjd8dIxMLozEPs4
DWuAEQptammpHW4IT5W/SPmwvaFlMDhyXYETk72/+RkVVbxmpx7kZ02AGIZMmxLDBqRdi4YZNs+N
HaYpThMtz0BKWSncg7u2ZHXdjASj+Go3k5bC8el2uKGccM9dvUhW4aUxJTTiTxyFd8AZWcgtMySQ
ddw/J0RCVKPd2QoZQtIFTwZ3utPfiwpsXS0YP3JGEUpbwqEq9omcOKNuy/6BA8OttMLP3NjLeg3+
e3/y5V9ZcmmpKm8dAGkqjNvT5SGsOrp9c24yHh88DmP9udgS3gfSEU6eXs/1Qf8KbMTAKMLI1t6D
pJfjFsbxZhR6yrGYtoQqCKuuGiRxDmiUyBHFwAuyGuRAIOKDE6mYesGbVRVt4q2IwyYbOWXsDnhc
pgKj+Nm7mlO5zO+qFG2TutH6DH40UltC5Pf/7Y4NmVi0ScexPr2beeUzuGMcXjHSbaTT3CNJ1iH3
u4kOL1XmTuuz9RYvCe0BKs6Bm3SIJ4za1pCvZjT59lxV1WX8JRtPCgqPego1orq0IVskhi7xKuur
NLSLsv/dtzCbGfN+LOLOGDY4jr5YTERIgr1UFa7HrQSNUaayF1Yk/Wn+rRg+5yLeraPuj8sW8C8J
HdcQxFr7JjzDWjlMU9oFqp9WzQERmmQl78wLQxoZ9NpkUGkIVocJNGNOh9iAjqr+L3c6UqXo7+l0
6PL8xiDkZQuAWbd1GV5n7XHeFoYfkAJNFy5jID+nLZdQbwM+BpudZKA796jnSkyhTLAEj/X+pVpF
KY3E1V2XkfWk+0bKRj/gs/TGg02WItkV5P2vST0yWrU0s22NlDASXoNkgMnxRVGxMmCLPbh2l6y5
8bXg5HWKIiAvq/R2uG4yZ4jqkiLc+6yYgh6P4giHM+61kLGAqbPepzYGk5/Qa97MjXGmbZck9cZ0
iMsEaGdt15uva7BlYuHEy0ijuiVQPEImowFuFvtkwzTlRtu0ou8OBMpHE35aS7vU6siSl2xNDV82
fP3wwO5h4JvMoLTavckveRS38aOIdhSt8c2Hy0nY1acDwXw8P0mlOnlKEFg3K7NKFdGLphq5ohTw
+x2IWeu+xzST9B/Crkpg07xPAuWO8UUToZ5o17JnEgn2bhV+ZWatg//J/5TFRUVkuJZ/T/MjHQ6t
uw882rrA0kgSwLMIC+LHFuM70obeJyZdU1uywBXM0PdoMQRkKGJFBkDGGdmt7WvQrc3nTREpQV3r
m05Obzm2zsjAs/Flp4nwNeTRaJokwzeobcq4Kk7qBY5BVsce1V5icYYImqcDaDIBb6EPiDAIkvZ7
uni+Covi1LwAUfseD4O7zWIf0ogxbd9E2vfBDWPGvXqxqhHAZkuTO4pELyXByZ3Yb61g60+u5PzH
PLdjc2Hl75+/G3WTL+l57AvLrCvBZYYOqjem+vSgaJbJ8eQDDl5o49gcL+/4roKMt8TZZYDX9TvQ
tsjfd6jBN/revZaZIRwy0c7/Qy9TYJCEtrbpz/9C3sPpGbbPc06TQBA0XkSwDO1F+DwoyU0T+Baf
IR1wujTWgTdiInJb9I4OEByimKfupNAUMWGhGhyIhSJrNB9sUWT6wzgFIYsnHrnBC491xEshj8jn
qGznydyD/YgtlK4Ll1ESqYHBiE4f1MIoYj3GycjojDp80Vc7fFpfmcPh0QiASQdF5jy+6Yk7WSwk
B6k/wAV+TVgb9lZS2je4JbrIbxqoRZrP0ifoQl5iU3aC673vgxq4/oG63jo66JLqNGJY2dVKS4Nf
XloweTwDCRKU7bUQFhv8WsbdBzu1tJKf5znjG8tqsrEstl4f+8y8yHzNk4VkR8TBI/4OLfW/cPNM
KL5JYV/xms5A2IPMCUV9DM7abh7v1IQY7kWVF/W3NRcTEH5wvTNRADxGHZjWyQG7H/Nt+EOkJRTv
X3ItSDSsd/Rm/6tMLN0dRUW8OKXfD63wuGs9zN6EKHlLRF2Pux4MRBtL5wgCq+9PYHK8faS6LBxR
MmOVt6+ShzspP9O6Ms/5v0T3wVkzCgr7H6d7VfQzydYVSs3kYJ0Ei7jW8q2sVqEuzBnPCKR1IeZz
Jyni8pEjUgQCUohWzMl8TNS3DFl/zq0GYzgvH+nxROzCJx5QvQQ72V2GCI+gZtbwnAc/BiebnFXv
NC5wIvq/qTXBtDTAtNPmytRJuV0pQg9fseeGXuHv8gDXx1aBqmAZtbi44taum4DL5QNY52m3ciKH
jEWdjHVsAlFxFH57jh0xibzsizkQGKCJ4TWArVFk6QiyYWsc1mObVO3DLNTb2zFn6PLr6qfSTolm
LaLclz9tuNGR7ETWoALFzkxK9X4He0EslbnVEq92zczt5XGYvO+KhrbK9QW9iunB/7PasJahXF0X
DsX1JPEjjs1Axr/XIY/R7mjlLGpXY6toCoc9lzg/8gnbf43uTG3KCISHZxExRTDsw093aa6dEJp+
tqV9CgJUNJgtBN9jUFsbZ5y2t129xwl/4pmawrck7oj79Bi3yj3PI21olcwsfTdEfOEssIrM7YY+
yyb7UyJkkieijN6XZUrBIOCgzn7qF03ZR4u70+BWX/Tqc76MxF6FVPEdZsihHRRYhSgKrm+OUvHz
MajxRlB/SZ/t0O2n9zomA1XsAdT4o766Uqx2ycyDe5Re03N05jNN9M8amFpuAqIvUXSyVbyAsjSP
8qQfIGqvu1UOz+KAJN05+8QOt+9J0XIlIcP0XxKQokofg2K+GKEvEe5hfe6VZLyKv0PUmVFTl8Mt
Ux+6j4gSjAmUERUW5UCjzFQmpI6Dqrn3/hQApXSCI4GRDrXHyNHKthATJkNfwl8SWRPu1t7HTeBB
gnx90iURTaq6VbBcmC0E4v7dcag2ljaxrbqn3w2trWu1yfPm2eEnJ5k1/OHrb6NItIEwhGJ9UHo5
+IVFMaDSrkC0SA1tGWI9cd18WVDClblAUyxFdzBf5tD9+IkZvY52cfzjBDtg+iGvZ4W86Jikwswi
6pjRx43OKimjHjB2/WHGGODv55m13nH2Vv5CrQh9YhteiXtnS8mNxguf0gLbTbFbSjERYwwZbO0O
WLEtl6DurF+QACZnq6kEQQMsXsceVfHjpohve8tWnz2YDX9fCcVMXp3nZFbf70bsKMBKqLiztxHn
SKKn8kaOlK4YeWSeX20Q97FII6HOjmHRQ1D54VY4ZuJK4vErg5Og6buquEkDT1NBSptCM1PBJbTD
dntSPz1Y8Rg+mNbN5G1vacj52AGWSkgUyrqBvTlHFbBZV6B17MnvRHcbT1cWTisE3D2tPePD8qkA
icK/4qyvpVyLHwui7V6NK+srZqU3FwR7nqsVR9dEBof2EWgCxm28hEW+k/MOcSQEimhoDvD2rtrk
quCKQrisx/Hz3QrlB2LaZAd/gWy3s39X01/Wb4dxbDTk5iK3vKAeT7PxMRnvEVY9amdENOrjx9nG
FKAF3P6At/3Xl9r5YHxInkrzsvcv3YgaHAvkZ3BpxCbh9OpgzBZkQih4lud7M6dtossmSDjOVoeV
4cIuYpy6hKNlCTq6QtfTwX1I02o7S2gLxLUG1APz/dyLmo2SCzUoNzE/t5Ccyf9Y1jSX9v94dyYi
2gCaRBk55K1ianUYQpm6N3Uxib7u0rZaG6UnHZwhsd1xZ0CSLN1pSWYGFhXSCy6OKYRVCV0O3DTv
CWlHUlJ7Ucnw3eCysJ/SFDpkF3Ln5ozefoxYXAbbgPXn/E7qfT82YuHmkPe8NE63yDGqA7jNCT1w
v7gcGqMhE3anoBfzC9Up3Qp9+K9FvPRsO60Eqh4fsY6bvt8h/K8ElqwyzP+qu+li7fEccogCPbM4
SDU34y/sDBX7B2isDdVK4CwWpup7TD6irazjgsWMgWZZcfsx1o+ouRRQLAdBJiq/1l13Vs/LS0vT
uottr0pKHk8NheqUNAsvQHFBaqoEdCjmzPRUXb6Q4BJp850kqPiwX3ufWvWSYHSQ8eOcJ06YkYDp
tvs/yNuRHgxVS+sM0N5dk9r6v7hsbGEG7IB52wgqITnj/j2GOqxCyY0m75OR/HzuzVYqnh/G2Sun
qpIwuqYZwaw6bUF5wshX2ty4y7l9Ege+Qk6LJD7IL9ssWp97n2dRQqlRPTZUIajkLjhmY2+e8puH
0HPgadv6GPAAJxK+E7pFRYLHYs9IppWSVI5iG5IErXPDUi9wt44fl2VrHPfjy4CROBBVi1ctShhi
ZU8hTtltSyQ0T10yRMo+eQ70gXmVEjKOR9KnvLK57HyJZd9amoLHKCOCcPPpRMtsVepLiXXxicRF
Pjt6wW7oZnUnWr6EIb1BQTC9dwVuZsZXnZjnyuEuGG3VekKW6cy9XSYbGtjqEvfSTNFJhUnMooaY
utd/cZaBAYGDmLwmzy/BYsElujHNhUjWV2JHWOb53PoObbjtPrBsc8HTXZ5GfHx3cYPOql+ayHda
/RiRwI5I1yB06X3yym3tJW/mB5cYcu6XONXQH/jiDHJvkpLk4i1Znym0DtbV6maIRovSOzmhTzJb
9OktiCo1stKiGVeHRpA/c1JWJHrMSHmTq/RWB+RhByxMvqefO8YVb/uVkLK+5ioQap2W8MEqaSXi
dw1XZCsJC/7MEaU/VWHEbhUiKF+gzZXgcDubPfUw9a+Jqsrr7R9f5IIhm7IrnhIjib0GlzpU6rRW
8P6BglkriERBMcZM5LTpvkmkZh0d7H30WUTny5ut87jr9/lQyxQCaqDvaOaCOR1/wrFY5tXtzRfO
ZaZwmxzTzkw0fyc+96f6VzdQOUU53SPvASj1SpueTP4iEsHjWiu+CBjmbUSi6zgZY5YXV9nPZRvE
MwYRBzx6YOeradxLQ+henVagdPdL9Bs2vjC59QxMF0txeyBmoPbqbNOSz9URsQlESHZJUHKBs9fd
RYFThEeQ7fWKAF6jfr5U6UZwiFYRNnC8l3cGr/MP5ZDF7uOlI7QLSEyIJ2ooYkWlQTmhMihe7Xuk
bbKt2nBXWVjBLrGVlHL0/uW56+a4OSPyZaK97LNu3P+V6AW9LP+2gqp3WQ7oVCO0NWwrtOQLEKAr
S7NDrSPgaefEow7hQ5HavgCLHxMgxi2ySE5W/g01aW92A3Eh1l88r5YJsjqwHrHisR6mEhEvGYy9
NSfUA+DZ7qQDpjCIquaIA//tksEo0p1ODPWA/NUFjDT7VA22Q1Iyzwq4Esbmv5RVjCNA01OEbhMn
o/3uRfwsGnQhPXGPVjR0sPMNPmxz3JFridCGJmF7Z+K7fFYUTuDCTY7/1eO0Kntj5+GNeOPX+lQM
p+sdr/sZD7TRtxAgFz9iPY0LEroNaxG1tKTRvMPYNpsc9+guk9PYYDGZSRoRY4FHVzVjPB117k6i
oTFlADUVS0i5GtMqAiT6XhzZRJgeEvQS6+RKNKkPlMBkNbga+gkNxmldrtrzuepl7EDe1//KU9xd
gZFVmW/YO/FuBKZLUgCoD3+r9X8iV8JDcMunQcA7rK43lyjAWt0KrgQkNkuvTfHW3CcbQ1YeY7RY
qV/S2qPiUsWsXKgWrQwgxwmG0/Czcs6fG6XcaTuXjFO+AslY7bQlwTsh1KIjphYdcwNmOZ06bcwv
jmEjW1PHHhUoyyH6LhcVHtjmAnTioWsaniGH+lqhOoxg0HQ9jM4QzHMwfWPeVHf9b3B1NmwkXeav
QkNHMcDgGiWz6XTNGK4eM/6mYmQRFAFJb/8eR4IvRcrqx0NEAWVSC4oNDODyTEcEJyRp9wYu4U9+
Lc/zEidlR7uTOC5CHHmtvaSRe2/JeLkDVY98msCxvdZdilQpzwK94Tsf3EVzS41ZJmjcd9Vuok+z
4MRkhzMLGRXCOKZmLd6KQFIlWo3hj6mvtvjBXstksQrSwm1cwcsMpFWPUp8P3we4k6cxt4Q7c3Mg
tlkD65WtMiGEKvldq2K2oy+x2n1LCmuTJAGdiRTtleUuFQvp0yA/zfk4cpCoXfrUThrsdNQEathC
TG3OVmOJMHqnAcTxhWttzNWMBkuhh8KG4+ocaxwizhQ2h4OTbSGSQ2gj1WTcxo6avyHjDGQSZveE
YUtCMCqxGhRntfUF+ATYRnGyy0zR2KR55SBetA0nMcBiVMlrTQr/oJEdShGLN+jJlRAPYIHAr1U8
TXN2KGmDZjo7AGFlUlv1izC1LS9Q5gW+kRsvEQ7ZKYYIXcUpLgoda+2yeUPPq7jY6BSkd1T5Yquh
IbvExeaqZnUGfH6FNghiwRrjh8MJcz20xIeu9bvCuKV+QkqjkUz76sMoIfyOmAMHbmXuC87MVcoh
Q8LSQU9KFpt/2DHH42X6C7r69x1HRm1b+fasTHI9URyxjnhs4lR3HI6hN+ospbtwBAlhW+yC6Lol
5iVmcPuSyrB3pGnzedPe+ZBtyZoBlX9zdHSXn12Lcl57T3J2vRJJ0Asd0QLbU7zD+Ud4JPfpJbua
fn+9MbjQ56IOs48jGtP37bSJ3O0RReJ5pnB8NJoyCP5wudHGRnQ08+K+ycjKnbBcQukuvjak8ThH
t8u/aF1AONlnuEvFoNbwscQGjl97t9SU8bmNlISsGx9XZYkKnoNfSgwiv/h8nV9qKed6LfibRBX9
erSPxn+iNiAG7iPgZ59w9LM9W8aIqxrdB5yhWvZa9nOLFhpPWqJGzQvJLSJQanpx0KfjOHvEuDh0
LtHZAYTZzZljXUmgPCsplwrIbPJf0DA2Ocsq+F37XHY9iYhh7BzoUU6xtUcMxm0hzfTeuo7wb86N
bCNMvHZYzsGBrKkPa9iRSBQiX3s5WfuoInmmQfXsknssYLpAQNFeg3Sl3MKpkpT6FJoHb0Q8iixQ
PMiC1SKPCQS/1kFiPyDMrcN4b4oLENQIk18D81NNvi6DPync/6GAhsjHagq55hQiDzsVTlkMxvPB
uwH03AJiG9JgK6x393sObFgnUADh1waylgG7xEfYf2rOXlGeYyS27aVs9yeu5KWbqhBC62l8XOQM
co8esB2HZdAnLRU183VE3bIkiOgjNCcit1aZwpSYWLpVomr2KjAy8TwUeQ/X3gDrBfewZWfkJZQE
/pk3EkIAiznghgexxo97WOnlRguaBE3l4mBmgeZjlRrrbJA5mpNkUnWoJdwkcHz5W131Inmc5iK5
H1KiYNSxmDgaVmOvZFMecu574UccLwdvvNwosBia6HR1gab2TbE/korGG82aVDexmh4apZ6bploR
4sbjnmqetj6VuNTUKDISBEFNkUergZ7Fp1gGwgzkm63JnWgljLdWJRexQ6PtelYSZ2AL37Axq2mS
VdAworn3oJciVOkTerzM75t/H3H8iPdEMXiiYlncJSergpJWFG4ox2CzH2lS0jLcNTv3LZdGPgGl
j7v6WYMRvhXLSMJxuOjQt2iWT+Gd5atDcPFzqiJSom5arL3CrC3CGuqR20AisAzjqB+4Cdfe/hwT
6qX8mE8vH9Ptsay8J6Wvj2XIlGY9E2UwwajlvhS003chnto3neFgNGYfB400X2L/+l9e30fGxAem
Q+cDDjaEOlzeVQNbW7R8+tNgK3TBT6rqtStfy9+Oy2sbAJFMY+fZDpG5PwPiAZa2QfTiFogy7VDG
SgK1y3/cn77DPsAzBWDli2Mcvi0oT9EIZQNJFPkSkgL1ag+psjA92QM9zdnzmIFxo5xjPjlyXEvm
Oji+gVclzfioWDey2QFzpPneYmk8Ew3DHoLj4mYwz499jpVJIWIDQQmQeYBN0ZAAshA2lK9oOaQt
c21EM8AzoxDmi6ImzHHFSN/bYwBxwofmxrt9yxY7ZPQYfhLA55p57urlcBL8xNOdntcKvNEWXpTK
v0eGAHkaUId3s0ckZTin10HgJPo1nybORAy7aAdIu9QqFqEMHnLuNDHeR7jcoENsJGzujMZA/THF
pTBBT9WXdWLaPkhpPVNFNdVuoKBgxNeS7A0zjWkxNDeFOlEfBnfVkSUR2B071EtdsBKP9ud/WBNt
hM3nRTDjYMpm8Il5GgSPOXb1Wbu06Lp7jVOpbjlf971idJ+Vl4vgiZdt2cc+kBfxmDnkRjSY2DFo
FELF1nOm0nu8navEvhHDM8Qzlibkn3eF98y7KJptZNyPG+FFmzU+CgAOqSwtvIQeFx+cMgwJC1p9
JKdA0Zo9mL5oCuQq5iFVsp9zeeJN3U2xB4mny9I1CHrEpVsRtF9vy4fe5hB9PHQUUCqoVXVRE+6Z
kkgMk7xYa5JV9r7+Koo+8yIzqt75pxHnQ5nrpetkYOnanKC9tiItvmEucuwfMkBOCqfrZ6dc/7sw
ozB5/RguqptYWsvvhmJwQ/iq3LOFbKbUj5pmdDAvT3an7pKYTgkKEw0fmyRUw52tY8iAoSEWUvL7
3EEjWhqm1/V2xaOn6JCwiu1SsugkpiTiJm82hdpBBbBZanKkYsIsS5rlKkoQPkLjMezEFgPAijEr
b6ovD7GfFhemDjV7QVJz3cGdK5GbcdkVVsP6wUhsCtNiuZ8/nwjcNhYL9ZFAW8RO1J2MaqHsdvoH
iuNzS8CRH5dKbS8sYLJEArG7dm0KxshGssBJCQymyDkskc6fj+k3y9kt4SZFXwAzRhDGywgCvbsn
7UnRpgGlcbZG5V/qNno35UTkSwmYBthknmYIwofK3igb0WlLym9QYrtfSY+yRm0DBIs5F3gfV7k0
aiDPntNKloi1GMQwzP91zwxvd+84yphuYsqguxwRlmxVoHYEsKIMKokZ7WJK742qowasyyFi0cLH
T5aZLRsWRJ2O0ffBjfw6SccVZUOYeNhNhb1XZyX+S8NZr4WB4D2K0URJccMAhNl+wf24sja6BSag
WEsMeKMBKk5j/5B9p/0eqQp9tA2qa4/+id7xQM2+T+gVOn8BUgGzezSr0VoJMu4ZJYBpp+PSATFn
n8tOufbPAITEK0fbjkN6hciLChvHBbBM9OUwf6EF2PvIq119eY2QBmM2k7UySyUCJsylPAElrZcx
aZCmlGy2+4W/JHIFeP0AigTnU+Yi/rcUvQ/Y+t9uHU2q9cEqRPnB25bHmJ3q1g+sBsnio0U3Qz84
SWgBdb/TfVsyy2kesBr+X4ScxA9prc2VbjgClAanHIl62efuiXVPcmkvi0+uWLC07DD0xiux/RQs
vehc8z3qqPNNEsIBQhv9e8tkJEvgbt0G90RXY94L8Bo68QtyUwjQljTXYddrt1yf37rpQODt+hBI
a4NpSMTaiKxQlgWg1m+QYME+UtwJ7PNDRMVijIMv6PMGAc/Jkp4yrRax4M5bJK7eVRHtToyRFKEG
B+VsLVh8+6hczhUsEtQUC5vB/vn6qDTrqXK1+pFfj6qoIRxBlAiwC8Lz5+QSWujsPJDpkc4ACZ9A
5urEs2wHMKpT3DU1RQmgUQVysjTe6ABUSPJCxAjS3Y1i+qM3oxYzRnUEu1ropPP59qRR1qj7gayJ
qKeFZObdi9J/n/yTI7IFmqVGACoQd7yj97eryM8ByqwpuglSStAAKa7tdaKdBz24vPwzOI81LkFq
a3KIFBs35Kw0SNfrwuVcd5fTA0O9pJzCb9FSfhu+/VuaopdSvVimJWoFjgZjdQ==
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�BE��Cfl�����1T���o�J�Q<K)-C�`��on$�-�V��)dk��!#eo���<�+�,���ȮE��Φg'��ʥ�G��?Q�~'sXOUh��>�c#�����S*��d��X������Lw�-��]�P�X-����#����6�mCJ������)=2b&RW��*��m/ �@��"�I�� ۘ���|���f��fu�H�H���,d���HN�[��Y�<�=��1���_�A�KW_%�[Ո�6����Z��^�8��8�G(���]Ü��\M��>��|r��=2r{܈�̪7���W��Qz3ZR*��1�s#��Q>�j.���s�`��H�p4�$��E s
���s����7uf����T�k!�_Y���-��OI��?£ �q�2K�`�96�"�p�"t������M�lB�{**C\�O���5�~3�z�Hh����]z(V+Q@8��}����I��=��(��O7J�vc�L�#�ei!��
N���;NT$gi3��-r�J&5�'�U?`���I����EM32������{)���+� Z���է�g̠T>�����9-(��c�IP�ٶQ�#�����
��m0��'�ݙ��ǻ�,<�UhWiˑ�h��ZF��ʋ�yLJ���tT^�'T�s��w1���	�Z6g�E�UDe1oX\c���DJ�=�bԋ��X�
�r��T3����뺦?$ ߧ}��H����i#�;�.�_��M��p�5��EA�t�s\�w��c^��զFӋ6+jm��	���u+�?�^p�r�ı��N�v�������Q�!���")��!Pd.���&��o�,ko�3�+��r�R��鈧�s*��-!A�?pȡ�:'�b{�V�LE@���%9=��j�����G����"��m���	*���]��q8.�ݦ�*A��D����:#Z�>A�#���̑��{}���Y!e5�<���ݣ�� cF.V}�����,^a���X���pX�RV���"X�ף��%��{�ړ]�7�����h{4.�d㳾4�^z�@mCQn鳖@��9������΋
�Z�d13*��wO�&�N���/O�:O���	�d�)��4����D�
��9A��e*0\��r��93s5�x���x����W��~�>J�s������'�q<�#�4�Q�_�7�����Q{��OLl��R'Dޣ]U��&���/bet��QXZ%�%�K�I����ćoڭqMD�n4��Mjw3�fZ!Ӌ�#X0*�Z��-9��K�UX��3,!�j9�kt�N/��s!7/p2�y�f���Ջ����5#j>��,F�������I!����z�S�D��&7��N��}�/��̼`mvGq�+q�D"��s��Sx�йJ)M�%���	X�w"�1%V�|�d��lƟ���2��J��s��2��.��i��)���i��0P'���p((�$	#9�~�	�����=�W�0@�-#�����t&�4Q���d��q@������;wZ�0X����ь`��G�n��(U?�\��4Px��@4��[u�.f�@���-_혘2N�i�Q~Aw��Y�ʑm��s��vB::�t`���P��l�d��� E��兜hCs��֓�(@+��TO�%/V�l=8S��7���ڐ����ه��j��|9����G�ݵY����ǵ.��!w�� �C�2ΆՇ8��kqxNl�&�}g�-�Ō��x7�.�
���~h�G�L����YBܪ�
�#B�c[�QP��H3[3q����fr	����C��/_y�`�Ӳ�n%J��F�#�^��!yK�[�5{����.�e���_0G�R�D���u�o��:�ex�?a`х�{H8���
��̅��*V�`���6�;>�d��3�nB!?��d c��*t?i�*�hoa=�))'7��1_P��ĚnPހЫ��-L�Y����5%� WH�,�����8�W�K��vYb�7�m�M<@�IQV��M�gT�;1�[c��H��c�	ݒW�zf*�>vhtލ�QG��z�Ԟ��!��X^�k��Pˑ5Ψ�Иc�������2d���Q��f���P֩!*�[�6�kXC��s7��<Do�@�yF:T7<�g��~փ=���yfu���BI��rbR� Ϸr�0��Tr��[��%?K���O�BO@9�B�Dn1n�9���Iq`J�[�p�{����S����	����Lu�"H�!���$�"������PJ�=J��x8�J�+�Ϲ���l�w���hsV�I�Ѿ4dY�ם:S�H���p������+��P���Qyv	��nQT����ԇ��֏1��E���-W��R%\f�M�$�,F�|�Uy�������#+�؊�����X���2X���/K��6���<Q�w�i���6c�}>�6ܻ�|PQ��|���r�ڒ�7��J���9�=�z>��6m���O��$:Ѿ%�A=��Jb@l9�e@�P��ׯYu��z����[=�!~ 4p��͇q k��q
�����%�ȣ�rkp��3���b����G�T�>���O{D���A��}��jH���<�N1X�&ކ�w�0�2[ҋy�MX�R2Y	Uq�@J7�Y��k�6��'u�žZ�[cg�Ǩ��Q�o3;�Wd��~��ay�X�߅����jnCmS���
?5C�� 	��N����c�f��y��H�	w%��؜�:�w]1�b� `p\�T��9����q��7�Ζ�ڌ����`�t�)y?[��m�螋���V=��j��Ԣ�9�?K�3��v=&�� �_��>��Z'�H]�|�C���	�0Rl�4[�Xɍ�����ބz��]��Y�l���p��z[���Tݾ��:��=S{��]�B?ħ����7�w7�9��[�� G���F�6o�I�q�NWS��Dw�M��A��,X��P|�F��?��%�k[yz���-����oEnm��Vz�RւK�H�w�i"�{žx]ex�X��Y6���o^��||�,�d�q>�luoڼ���'$6Ѭ��;�;c��*�<�Q(l@�޹���G�"�P��7��?�1{�����=PZw�$>�Jv�v<��B��luRN�/��w��8���R'�����=�4/
z]�İ�<�鎯�}-��&o<�a�p+\bW��lh@��,���pǛXZ�V����6�aam=�.�d]^
3>j�9�.kfW�S��)X�o�^�nrϚQ��$$�8.~K>9��uQ/���Q_2ߥ)�Ø6������yM^��7��`"~������.'�e�8Gۃ ��I�˽��`��yi�VC:z�7�O��|���r}���[��S����u;�<m�-s�I2Q9]���S������ KjP�G�iK�o�?�䙯e4z��b}|��f-�Ⅺ�i@RyǞ�/�d���8G��Zӝc��:(���G_Y9�� �-��ū�8���I�n
h����|)1��#r=V5@������}�<���x�k�Iϡ�K�~�~:����D��Ab5����b1X������l�TTxn��K}��0pi��u ���#�l� ���Տ�o�n*`k>2��f��$�>E��=�����W\yb8�e��͘��W�ʸJ��	�����n+[b�t�[�bRl]#��sCΫ�ø��'�|�|�� 셉���A4�YZ�m�@�0$��T�u�bR&ݴp��Q7�(}r�i�h�?�������s���v0��Ð�<^0�3�媪!�h�QF�i4�cgd��9J�=�+ޭ$�o���f.�Gs���������*=l�\�@c�I�>̭|�����쓊Hg5��sf~87ku�Q��O�w�����?��,:BLn�{&���Sئg��8�#.sF�&�fw����r����eV�I�]��Do2~���
b=�E�P1�y2``}Tb&c&��Nwh�m*'!?Gj��� �M\�M�/��u�6���\��C��ÐZ�ʱY�y]�1^`���eT�\~tlA�}b}�)�_��Uh<�4�`�z�~���'̽��O\T����ƥɻ5�W@3Vǻ�`����"�3e�|F8�W��B�t7�.��8���V��A� W��
�K�R��V&w�v.���
9%��y$�]���Wp���{�@���nx����&��n���-����ʠ�&5�l4�7�*�Cܴa=Z+��0����D��� �c�8U�~X�����h_~j�����n��:���pԭ[[Oe��ZX��2���,�<�[�l��R�a�^���V�.j{mG�}��ƪ	�+)eH���X-�"���4.�0��Zv�څ�Tյ!�w�P5F=n�:,e�����B��b4ƬB�	V�D��S\E�����۷gb� 23��(�N���Q�e��s���X,I���R8�uC��FP��-9�?F�s��)�,����svE�����=S�!��k��
2�Qp*�F1:jp��;;B&�b�{���������󣠉�Erg����)!A��8e��j]`�5����D^e~㠇fX ��x�f�s�s}��� ]K��[�^���PĒ����n匲".�t���iE���p�)+
����%#8G</S!�x�}3[�/$)�u���4D�5̒KVi�Muhd��%,5�2�t��#�l>��c�����gM�!ׇ���Rnāc��*��X*{gv:��@���H�)���,�nמoh�N_	�.��X�?��f�-��/���n7��-Gq�ء�?�D�C�բ�M=����t�i�jBR�/ݏ�fv��/�;a��.��^�â�U��$.�#,�b4x�΅��ײ�Q��ߙ-�?�5�4sW�e���:��@�G�-!�]^��pg]��f������˃�@��g�<�P���Yxב��]0W�i;��-b�(m���P�8��i"�L��j���6�H��g�̒0�21��r��&a0�3E1�VZNi�[ա�ܓN������a�%���L,��o��`���Z|���{�iN�R��ޭ	A�sUB������Aqڥ=�pW׸@�s�Vq�����$LNJi�E�$Qj,}��7ӝ.&�KؘOr�V��Ee�6=�浦�(�M˳ �,��h� )����`�C�g!q
�!?�c������Ƌ������jq�®.�Έ�[au���]� if�H�ȇk �*!`�����ݶ�	+�P��ӽݚ��)՝Nz��%�W�6�k��~�2��C��$���T�lo6�X��E�'���Cg)��o�����`M�f��?��1�d8ݠR������EZ�E?T�;�i+�F7��/"ђu����e���e-�Z�9�<@�xR��3}K�BҲ��-KwcXp���Gڵ1Onh�do摯�s>[$Kt�-3�d�!����S.�<,� �3ܾm`���_�����R/�i9��fP�d$�f��AґҐ���oƯ�[�NV��l��Fte�ڏ��֞q��/DŞ�0����[�/jc���>r��:ol�?7]d_4��)[!��zx�_ҩ�N�;*�T�?�W�;w��0������ܶ}�I�*��7[�����;C���*�7/�0^ʁ�� A�nJ��USp����9�cm���{�a}M��b�o �J�Ըj�~�@;�"�;��P_Ѱ����e���&�U��`K`�������}Ez��/���j�'-�k�	�'W0�6�^�g������y	��0I^���k��xH�g�v���\T�����A�$��sc������_�#�Ս�5�Hf�r�z��MN�]Jf3d6?$��WM���p�fKڱB\���]��������ZB�3�ۗ�(s���z��e'�'Z7}�2^�)�ħ�χL[U.�q,�|���Z���q� iW|��9HE��u��}$�	kq*e26M��Bl5�����.�E+�mX�7$��m�!c}�k$yNҾO���'��,8�Є��ھ���S@I���Kiʹ]e4z����\A@��r�F)oA#~f׿p� Y�w��������E��TV���*z7<�1,�2ɰ<�g��
��m?}_"�g�v��R!q��oH�����*Q�P���~��wZ��Y�zU�9�🕴Z�'AE�Hȿ7i M���e=�o+�u`2#`�<@�9체�u��9a��f6*�Oٔ�|�v*�^�ko���J"� 1���א�N#�
9u��D��'MWw̥.�������P�T��x�.˭s�H2���xB��R�G�%��
"���5**�f�%)��3��ޢ�j�T^Z���)�1
R�H/75{=�}���٤R��@��濄q"_�.s����H��DMp�Dz��2J}_v�Y@^N.��qW뢪܋"k�����ƶ�Ҟ���� ����Ѡ�Z4C��u�$��7_b8<%Uݬ���*���8��c:�
$�W�uUfj����g( �n��XX���E��\E�	G���;�P�|��wS���Hk��U���]��-V��]?y�,B�ى�sګ�W���yV��"'g ���	�%��oɾx&\������{�,�fm�*K <��F�Of��q��p�_�.aJ����f?�E�:0 ��޴�-���}����$g�ZQj���o��'�	��M�32{�#�h��4�&O%��&��P��]���7G\�j�[�ύ��:>��`oЕ�;r}I_��4� ��2|�L�������<3�  ��*�U���������!#΍��RT���a���
�d\փa�Y��m(T����Y93f����R�$X�/���&�|fU��1��M��a����$Z��V�g#�p�6w�>m�!Y^ǿ��Blt�@�,u�νc�� �%�8a+�',�7h�+��Qp����3��b��$��8��*��Q73�b��_��](/&��[+<t�[��<� ����=bE�R�2�Ƥ(d�xV��q�@���8�q�5z������Q��@��4a�an��=e�a��7�v���GS}��s.��()4����+�0������E��5�$�F��,���X��Ј��78�P!��)~T���8�`->�`�+0c��GYZͿ[�m�EZ���Q-�m{��M���\��Ef�h0BS�P�"�\�8�ԕ�h�;G�gmb��S7�⟨��C��u�H���(�A��MՆ��� ��(b��Un�Őt�k��锗	���z�����&3�ga�9��c�6�|�$0Aw�)i��p��*����IFџ�v9R�d�˨7����V@<@D���Q_�qk�m	[P:�|!ধr�A����b��$i7'M�?�J�bCA�ٸ'm�%���b:[M��ڰ�������L�c\��^��$%�[�KU����qv�MT��+�J�q���NI�D�n��%�b�v�w��S}�:�K����^�n�"�� !x����� Z ӹ^��~�݌�JG�)p�E�-h��駣*~�Þ;s���&�"���|H���vQ�u��Z7�X1I{X��m�opag��j�6)a�7��!���>�3r��-a��Z���7�C*C�#@��T��fvFt�~�`3j��s��=�'.����}�A2���0�c��r�Zw�9��F�WdQ�� @W)=��=3xֽ�JE����i���o�m����S|�s�=��, ����[�z%顰���2���
%����������+Ɉ���6 01���A���k�l	�	��e6S^z�9�Q.Pb+E�5�����O�U#i��G�bL5�B0��-Fҧ=��XW����T��h-A�<�ddmU07#����@Y�}��3/"{ 2ja��Kh�=�,�5l��*G�1V@�����%
c�&\���ڞrq���U�? l�]�o�X�.�
��"8�,�����dh
�]�{����L�$����CC�S��cm�R��K��7�4�%�^�|vMR&���cI2k�,)�^-c�#��'�{H�.k��H8�4̤O+`��f����xKP֝���:���I������N���{u����»ȷ�lュ[�Q'=��m���l�`� ���reE��;<F��8�x�`�3�0b<�p��W�[�*\�Π�A�ߖ]o�vq������X��+;6!D-�3��-GS3ʹǇ�r�
�#Z��ͷ�W\3k&�h_{���
��b��ޕp-x��񂔢�9���?2�Y�0"!�؅�2�_�f���&�Һ��3S=4�gz��Փ�w��;D.����48� 2|K8#�lQ���͑���AΖ����X�	y�'��i�Z�&aޮ�Q�Ew@8QF���~<E�q�j��26��y)s���d c��6�{K�O���]�d}��?y��N���h�2��.H���^���.��!�M���U�ǌ�:ɱ��4�[(K�l��P&=*�%ʔ(� ��a�vZ���
�ھ�KKR� �X�ܹ�<%�w��̪�k�+�L��)�(��>ٞԷ���>����i���<Nmj A~� pJ����� &�T�Pxʇڬ�ұ��T��i�[Lyg�՜?(غ*���\e�Hk�؍K����u���#����A���4NxF��|�D�淴=�%��f�O.�9e��T�2 L��^�/�\R#;��v��u��ɪ��J,R����ǃ�_�1˜u2~)�^�kw�Sl��`��E}ݽ�Xa�����S\���M�}�*/�gk�)_'����%�����7���s,QU0'rdW�i[���By� XY�jՁ	XH�gS$d���zhN)ƾ��7�]XJ��EnQ]�*�mQ��p���4dHAgN���.<��y�����IL�v�s(&\�D���n4!�6{��� B�cB��o z��u�5��y|_E�q�þL�?Y(R
7�Z��2���)|Q��:��a�.M�U���hEo�K��+X֦�Y��;���w)n��	b�R��zG˫����o��WQ����j��;�D% ^��oz;O�د=M8�6W`d�!���fd>����78.���yß�m��pR;ZD��@!nЋ��M��C�EqY�'v�Ѯ}��g��d@EPѻ��u�w�|��+��y��o'�D���s#�J�~U�-\=��q�l	�4N����uR�b��>���_��aT
�����Yjt���d�l���f�����b*P�X�Vz��N1�˸	Q�z��}����_����_�|u�eǯ��l������(��d)U�d����W����:�O���3��Yz��(�H[$�K��Uѫ0n_�!�#f.�M���?cj6�D��:V���S�hU[��no���@&�h��#
&
W4���-��
l�J���[�aq�b���w��楄���r�U^�m��$�Y�OG6GfQ����y���M^��h��XB�spo�0ϝ�4�"��[[YM���+�����y��[�M�M�\�./����MbGmHW�APM:�0�H~�����AG�h��@��.}��P�Bpb�b��uܚ�5(�ƻ`v0>?�f^{��D�y��`5M��7���$�P�H���V|vz�3<X�dyS\�Q|2m�f]MxG�a�s��0�>Jb H��׽�ÍCC����J��wk������p���'��g`'�����R�w��5ej!�]6�\b��Nbo %��jwu�Zz kݖ0�z�yDm�m�4�K��n�|�1^��Ѻ���I�N��q	߳Լ��_�=ָ���lp�Y��p2�}M��g��w	e������wZ8�__�d#?����2�5����z���'�|T� ��� �|�S���l�����ٱ��Ȕ�Bp/�`՟bߝ�޳Z���ya���4�T����ַ�� ��*ZD�+��j�F|��&�(��b���wx�	��g~��YP0���U�J���X#v�	�i��*&��\����Jmm+�to��^��׽���nc	�O���}V�RTS���aP/0}���a3��C](zߵx&�`ݨq.l�df���鐒G[F[�}96���T������H�t
z��F��&�Xzc ��KТ���3:�q�n�9��Z}�@�#<jW���醉�6����Q�8�a]�$��&�@���ɧ"�V���.��Do��R�p�8=�ӦW��lQ�wX�����H\gc@���-�8 2�YG�
(�0�|�ʌ{�"isHi�J�i�Ȧ�`Ԡ�cYc�cm�b�5}��aͷ���Wb��;W;ɏaoe��{ӄ&�P���}{�]@�{.��D8eW���ݘ�X>��}qe��#,�ڽ9ͱ��c�nM	��֒G��<����I�V�wM3�v5� ����Ñ71tQ,��\��0I��mI"���U��%�v�l��f>�Iq=����}	��t�g���dep������?���i�!�j\���&�'�/�@�x�����r�C����9�Fe�of������l��=��8;U�T+����g�w˥�&i��G=I�����ij<��F/ͧ��,_Ɣ�.�ɰI��]�m�����ӍK�x��2(��͍,k�2��ρ5�����d%p��'�%e��ZU�kzmg�)�i&N��2<��� �yj��l�.(�+�c+������IF�; ���70��-�U�rN�v��I������,�1t�A�f=>��6_�(������[+�����5$HG�>�{����a����� �uLg��BRrD��f`�}!Ϗ'*1O���}�+�h�v<��حw�%A?�Z��k��+�T� L�O(��.�KI��|��6A��]�����	�Q�7�5~��\'6�idk�������~�����	�g�=��-�Ǡ(�n��9b�#z��Q����|� �$nx��y��&�bՂ3o(�aSC��T�<��tW]J���ڞ��Ya���_�1�W_�{`�t����Yw�#�,;�Y�2.°�T�+��*�nY�P��\���[j[���es�N �ݻ��:o7��qdJ�ʌ���+�l�8V�x���՝��0o�+��m������q4����O�����"�3O�<��p��pK}^t�U�מ�b���>���s��xJC���Z����U�/��1��J�ݑ�3�S�'�����c6&�'	^�,>7�]ǌGN��JѴ��W��F�	�,�6����+fݠW��0hW)?��o�$��{��!}�ߊ@4�$[mb-�E���ٺ�p`�ڢ�0ъ�Ry�<��K�%B��X����c��:�@���4D�c ��C��ę����Xf�����y97��&+&y~���۞��Jۯ�a)N��ۜg��5�&Qq�X�a��~˛��������O`��ϐp�[�����X�$q"�B�"�wQ�Ql����:[�<�d�b⹺�?���`��g9!a;V����`F�3�=�i=��r)�� 8|�X��=�$b�Vg�W�8���A�F����e_�^^T\�CJ0c��
�n�	�?c��~�2���ޅ�4�����L�Zp2�`�!{�0=�C1Y\0�fYP�D�K)3��(@�Q�ܞ=����GO���M}lQ�ڶ�#6]���L����ܚ�����);cx�U��}�I-�_�߆�^�T�xdà�3�����N�_/��j�}�լ����S���&��q,�}��89\�W+��~�з�DQ[�eg�1�Êg_
�+c�V-#2^�N/f�k�cd�x��bE.,���ǃw����Ahg:4�#s����ؖz�jZy���4Ǧp$��XN�iS/�ɂ&�.��y(�׸L�x����T�ђ=����K��_���ϻL��%t��Jb"wdI쬹W}���z���#VO���؍�,�Α>t@>����13�0F���=ք��(�k�S�!��c�60v���K:hʽ�D��YV� �ө���1��r=%<�U)��R�P1����G���{�*,[�Vݎ9k=Y���!�!�( ����u���(?�!�D:t�I�4�%JhZZ�4��p>��''kpn-j�}�T�,�Ĺ��C��^Q���K$[f*E]%�C��Ġ�|Sp���%�ǌa.�,V���a��0܋���X���;vSn<�n�&o�.N+��>���&�l �vG��鋆o�e{F�N����Ii]�R���q�ثaW̚6��REՔ#�'�����!;��tZ{��c�ŚgxOT���þ�����r�F��pD��nRbt�-�N���$�kA��rJ�Yi�j,J�e�;�t8��1).�|0χiXХf���C;���$_HH��rO)���*፨$'�&��I�Nd��0�s��h�'�)�g-�&�=��
'�Nk�1wg��gz�W)���|(~0�|��ӥQ�je��,G��.΍ٷ0گ}%H['�:&���#�q>5o�w�=Px�����yl�l��l��/��Ǯ��+El\�g�*RQA$-29��>+u��촻_��	z��26d�;�y6��|��3��WǗ���<�\�M�t�y��Rh�ƟlO|���� $S�il���w���7$O�9+G�ܿ-�SڞR�خG�-���2�/�x�����${��x�膦|�x����s�V���Iw)�ʓqw��X b�����|lN�3Cr�7���N��|
u��y�  
��Ag׺u�#UL�,"�:Ѣ(���4>���$U��z�w3\��s��T{a�*�1Y����<�v9�aKo*��L���T�;�=�`���`H'����>ʧ��*N��.a��0`�Pn>�2�=r>o(\�4�3��[�	��;�+$6	͊�]oo����5� ��.��\�6c��o��tꗯ��{P�U m�
��n�k����F9�1�������/��Eg���6<㿀� �厴�Z� Z9��1��
�]r��7-��?l�lz(���F���Aà�xְk�t/n7�* ���nO� ��j��A�tyW���!��BI�ʃ� ��w��L��/d��W��4���mL4��Pw��J/}nAW�� �#��sj������'�_�e�
sum�˃Nv��t��Qd�����G
���P�{y?�Zw��t<DUq��o����4�N��Ŭ�^��SN�	3���X�h��Q�%
�ꉓS�a�d��$��j��r�^v��6�D�jb����TߞW�V�e��E<]Qj���(K�!{"��(� ��v j�
&�����1dR��@�	�ݿo��5���&8��:T`j��)������*��9.�IF�r���f'	�K��Bd6-����ll�ɁE�7-��+kgh�m6�9��<��zg�[�)o�t+�3*���w���A|�Bw��.#Gq�c�.:nU�S[Rdo� l�ɭ¸n�G.wb`�~,;����f+���;��T
vl(㵇Z^Rv����8��_�/'c ؂k�$���+��# �!�ls��������nA	�Pn����� H��ҷ)=ǝ�llk%��X���.��u�u	�9U�>�U,�J�96��Q�{��#(���RZt�N1�es�~��6Q�ry!�M,���	u9�$؇�em�y5��Z��Z�?�.��/���������G�b�>I��?���'Jx�xYީ�\W��ҳ��[�.�N�&R))��;/����}qS9��3�0*��WU��Ѣ�1KN��Q㮁�������sL_�BM���E	i�R���g���5n�|ҳ��!M�Grk]�4[ߋJ���2z����k�ԊyX�2ԇ���~�CX�m�*e:��&�o]k��-G-ų��RE���fQ3Q+���ă�V���~��G��"7�>Z<��ж�����	
mL=�ajWG� ��g�[�2��)
�-�Y�n��9S|�U�y���vS�B���-� h�v� �
��>�=���SD�$.4B� с�*�4#g��'������1TBŗ��b�����Ci�/�r�e��^ǽXρAߧJ��(�6�-uF������蘅&�B;-x��R�~�m��"�2O�Q��.�do�OQ@�~��	,91��^35��t��ޣ��D�4F3�i�<p
�WD���~�9�	����1�mu�9r0�N�����<M��J�8&���h��&��ձ}�iO�����[��_����(��g1je�X��+4��nY�>�����C��\i����KБ��i��ܹ*s	��c�mO�ʸ%�������|�V�-�؜��E�N���Ag�M#@��L��/�=o.o)潙vҲ�yϳ?������U;F�j�8vS���1���,:��7��������g3 ������e�b1~L8t�V��*��!#i�!T�֏�_҇Ԧ�,�zd��[���E�Wnz����?��AmT�������|e����?��#�
{���V/� ��I@��,�&��\�@@c�}zqvAl�^$wT��/�7sF��Pޓ��;��1j9%)`��IY�mw4&ʓ���
�!�u�H/���ҥ�(~��x:�Yh�hd�ު>
�:�dA���b�3��'N_��MY��KÂ�r>@�-�Ń�����a��~�׀e�o���iv�R)�R�K�qg����D��$�VϏg9j'S18�"e�W��S�P���]�)�`��!����I���T�h�Jp��N0��352��"Te����s�¡��8��
nw�� _o@�I$�aK�*T߆\	��@��wG���Bh3J%�E�ն!�%Q��Fx��T}�8&��3�n�4�A$�%"ƍRc����N<��־4��D�m]hYCR�N������	�B��4��W5����"�yr�ʐy�����|X�/��7����Tו�"P���Z����z��۾]�Hw�f���ǈE��l�A�j�Q�\K�Ew�G���>S@��	%K�ӎ�jZ&�����H�MAPtam����]�\�fT����d��>qV�J�Jޤi����ݪ�Z�("k���xk���?o�:ʌ�W��裣���ȫ�<;UY�y^#��[���X>�^n�Z�Z9b����-�����3 =f��H��l/TK��P��Va*�~��' �UM���XE3��$"��"F��]��Mݨu.��>����k����Z��@+���;�v�>{�х�\�b[�)�>��-�����S���Qj��Ba�#s�1��x��\�]/c�	�6LQ��Y Ի1��K�[$#X���m*�Y/���t�ՀDE����w�Q�!R����0&L��*�w w�J��~�a�Q܃+�b
*�*Bbd~Hu�4�Ok-_i���~��,^L(;w��T?�L���ǧ���Y�v�Y}�]���s���K�}�״��6�b�J�ҁ����ĸ�<g��{_���f�l��_�$:r��D�y�� +L��k�Y�2���:�z7@P|�̝�5k��kdw�ࣹd3T����<7P S��Ù'����d�=�=#6�Q��~�<W�X�'���9��dfGpd}��i(2��a��B��o-��G#�m*��=\�Wt�td%�|��qʦ���<4����盘O����� kv��+�Zr�!����4^��c����ފ��i�D�GH|A;\nY��TQ  �!�eZ(��K��*���.��2D��A̷!�G�ǈ�c���x������z^`���R�]5`�V>��{�̥���?��j�2����MF�t���X \�|N���[�y�y��4�(�l,�)+���P!����S�$��[���-�6����ěi����N���yt�U�s�-�q��	s����`�� +�q��$-VkWF7�F`���O���wN�2�|ʮS�O�9�o=���$�D�^҆�ѵ5ܒ5�((R�"d�l���.����B���ؼ�\
m-�?�m.������d�,�ކQ��G<�2�����f�H˻��4�X�ncr'Z�	t��(�Fa=
S��5�ک�^�Ĩq���D=�\*,ŊL�O���@A�ܝɂ;�J�s��js��B�j�(V=�ժhC�͝}N~������W���������9�1��ðM0�==��ʽ�q�%a�c��Q��K��7�w�������u�ɡ�(/&�y����82��lyH��U)Nx���'J�a�����D$�lL�ߨM)H)�c_��K/|_-�SC�o�i0�w�$Ni/Q|�i>z� ���N����>�x9�E�	�E�֚r�I�����{�, ���I���ķ�F������~<�/u`o_*[ce�)_g���?�:2�w��0� d�[�Sk���:��)~E��r��P�Q[�A��+��?�:�J�kj�'�k�HaI���.*�Lµ���B��9B���ȇu�u)��3ngYW�M����$J���Y ���E��32~�&[�K���Om"�X�EVƙ��n�����G��J�,9����-�o��SKQ�P�o'�$�r@���DݷT�F�u�}��l�6�C��͠�R��mbby\��������d�yAC8�GL�$��7`N���+��R��s61���ٌ�(�����(1��[�=\�B�ccbi���"�KrBI��h���@u"S����� �����t)�#h��q�>+���.¹��V��JX��ۊ������˲�*t�[��Ү�ckD_;�GE��j�x9�9�ъX�W��#�R՗�Z��Z&� f��s��V R+��6ｖ����-�:	c�e WI�{1��� �|�i��@+�{�俒1��F7�i�@}�Y=
���Ɋ)��9��q1��#�1����b����\5K"Ft̀nYj��T��k�����bd��!r���r�.ƣ�°,��wA0��_2M*Q�8+[���Ynl@�5�g$&֟��_��?���J��C�x��RZ���X�J��^	�l�46� �M���V��T�&�n��Uk�-���ro]�0������\�qİ�@��DB��$��E=�!�~��قd�ұ�/�S_Cm�O�؍�=L����蘉4gi�xq�����6f���x�9h�=��V�Ú���;�ء�=;D���b�4��zx�ؕ����"KƆ�~It��x��H�k�J���S��Q�МAaE!��)���ƴE��1�	�>�Y/:A�w#@��nz� A��9-��<!s�ZE���s=� !E�2��'�tV�WY��#��
���{@R'�D���7 `�!�'�F�y:�*��}nt�'ok���Y?����O0�ջU��м�S�W\zC%Ч}ܠ�B�.a�3{��l�S`8�����?�������ņx��h�4�E����n⬷*r�=abm�4�tS��de������y��.=���T�G�M���Y#�'ԺA�^_5�I�����0��&�@��z-;N�ɂ� m���b�'�1^��XF�yr7`m�
�3a(��V��=����v��Y@d*�p��FX����\�m-],�VB�g��}"�ޮ�h�Q'��w"�Ser�9�n9�c6�Ȃ��0R����9���#�Ԑ�� �^+�IAD��>}.��+S����@uw�W��M}���)�P�pcŀ��� �v�u��Ѿ�K��]�����I	���5��^q���>GTSWe����;�ED�ܽ�U�*`L�4�JE��"q_�W�".-��x1�ԍ�H.�L8w����t��Q7�v�9{��"Z��)0%k��=�I��0�"SO4�~���]oi�'G��՛����j�3�~n�,�k�C��c����Jz����Z�7���v�| g�{�ǳo�k�/�Μ,�y�"}�8��%t�Y$���Zmزw>ǅ��T����
I���Se�>�|���F��9�Q�K����@r�;*~&�1MT`����H�<\����U��A��٦��5�aż��OLt�@.喎�8�inx� �!}�'~,0�4J�L�k�w����#�9%vE���KU��@��Oό�Q��̒�#:ZV��=��{:l�?�?���t�7:ϝ)�X��B�<m��LG^��+�ީ?
�<HE���>u�q9RB �ߟ�{�[�PѨ�3�=j>�<Ո�a�@�Hp���#����h)�!������/	��Z���5C�^4b��U=�6�ij��|�/��'��4���#U}�b(�Dd��8�2��Ի�Gˁ�H"�@�
0�����!"m��� �{��;�a0�[7uaGs�����8�Z�ؾ�ҧ𮂤2͋�Tvg�RJ�4t�$%�C�9�4���{���p����z�[�2t�\��(����[ea�k+��J̋
h�)/o#�H��b�L��	�ac��Rj����3�\y��<h����ڍE�y�tg߫=�J�yp��\��D;�E�i^���L�6a�jĽ�������u���PBV��Ύ9q�'�]9��@�'n��ą�fs7wWh\jL�	!����g/�4���'�G�ػ%D�G������x���N�����_A$�"�?V��P��l�t|��q�F��Hj�xV�n�-fg�z4k�Dꚭ��S��+@$e�j��ȶ���І[�1��`hr:J������z)�ۧ��T���-�p�����Qǂ�C�����//�Jl%Z��&Jr�L+g�e��kA�b6d\R�a��|۩���T��c��/,݋��A*
�����ƹhGT�5�g��xҲ]y:ҍ��>5��u +�-t��aE2�:T�bQQ�P`�����_�!W�>�
��h�a5�&q����N��3�)����Ε<9P:s
-"wv�Gii��<�Fl�$`_�VR�`�ήO�~B5L�K����]�@I@\=(s(3>B߬�M[����S�B;�2�)w<�� 2B��d{Z�>�M$�}�F)�ra�pwV��xpX�2h��p�``ݾNJv5Mٮ��H�yK<~�J���� i���!Ik��Kzlq8;@���/�[���f�ʑ.Qh:{/su֖������r���J�8�<��G�B��ދREU�Z��I�b(bA+ڮ#�lO�ꃚ��i���	�T�o��ӂ�AKZ4~�*��,���^�з΃x�����~rF��5��x���Х3��r G�5���r����n?L�n���D���>zG��'Gr�����N��Fv���K�E�
�e1��S��ZIy�ўjmp>���:<!w��.��ŊI����-�~[y�P�R~���԰I�WU'>�	%��"��8���9�pmjO!�}YN�S�#�ώ�����.W�~9H$L�l?%���s���zF;C����<(�ݠ�������tS�p� &�����y�$ӱ�b<��o;oJ���3ʏ`U��
��^��
���Pe^k;F���۴n~��U�
ID��
l(��(�k=6$�����͂-�M���֓i�̅
���K�^�c��`�/�X1���]�䘔�E��5��*��6����*5
��EɼM�1��qN��*��J�QH,N��5!u�SB�"j�͉��\��E��>���ÓK~-%4��U�N5 ����#�xwV�O�P�c�_��|qaG�Af�i'H�'d�}S��0�'�VL�`�Yą[�?��L�5G�<��ӏ���2η���o��U=ҿ���a���2�+o-JSR�`�S�� 8�� 3���v�m��,�Ɔ9֏�?�7Z���'�*�It��c������(�/ڀ�Y+#�z���:w����O[ľ<��߀N�$.���L*�2��?
[[�T!����y�PP?h7B�$o��bd��q�J�T������ϔ"a�ʼ�Yט~���J0�7>���e�G����{�o�_�*���S���}�����Q��S#{�Y�.>��*r�5�_]pd��q���?���q�ǌ��G�r��ʰ=�������&I͋ڑ��m�"C����QO������(.	P;�,&)���$�w�'��ӂzp�x�2��n����� ����'�)v�eÜ����b]V�m_p���Q�P�!zT�C�:[�&�^���ǍX��+��{���ɿ�hbX���[�7۹f� 
b{��������	�q�� y����@t^�f���(a6���Q�T=c�q�e%В�h���;V�v�l����l����O͜�Ff�F�  �#�H�  �:':���[�m�W^!��u�y��q��X>3�!&L�,*�a��T��Հ?M�/��X��c�P+��>ޢ�s��P��H��S�0��t��g�&+ 5j󍱆����܂�|e�)g9ړ��� ��\Ԩ�L)�i4��
��q��U�ԌA
(R1N�$����8I5p,"M>������]�`)��B�$��������"9�%r��iMȗ�3��k�!���7��e�w������������#�Kd��F�f���5ñ!:���`,@�gR���V�c���f����*y�%P'��v�F̏�_I���l8�iK���T)����`��l�:
���T$����h9��gC��8���ꖚ�+n��~�����E��J�|A�L k7��4�j��O�F�LZ���d���iEW��/~񁉗T��f��&��bg�:�=5<�j.��=u��ڑm��u����n��3�˷�T_��wO��h�DW�:�E(�y��)X��`G�����>p�Z�u���[�k���QC�2�l��xuz]�W���/_��(��X��=����ηa��8�񸨿��gv洌��p��^jb9<�*�Z�"u9��t{�
��3/J��b�#p��2�M�*ű��yj�|=���Z�6aܜ��KK��0�W�Y��;��E�XU�X�ꚸ�,,�~��M���@�����=Q���*���ьBĥJ}��Ƣ�L�]�Ig�s�������Tl��������敃��%F�'Zp A��e���{�T|x���yƃbl��_�5���c(<Q�,��
��\�Æ#��I�,��[��9>0��:�|jy����Bl�{��@����fS�4ʡEؖ�r�I�����[�&!�f�}q���'ޥ�k��=[i��`�71�B)L���
lo��A��Qfx0Pw�w�ս�K�S��8)\�:&�k��RD |>I�e��dr:�;���R礯�x��q��W
>�:l�'��2y�#cwV14�KH�QE��D��ھ��E�����?x��t��oW^}7��&��ófX1�� e���?t;��h�$�k>�)�P�\�i��������DC��Nϡ��Z9��4�\d�� ���a@�Q|*H�"�y�Lʀź���Q7
!��^�H=F�Sj(+N�ֺ��F�-�>P���U������T�l���C����0�3���;��@q�FC�	L1��C|^W�2Z��7��*E���VX�f��e5 ?ֈB3J�a?w}���5�ٲWZy��2�%��!��']��V?�4=h/�_ i�?:��a>L��X��GE1� /�bvE��̇R�Q�&���Ylp��o�uUO�ũe���9[��E	!�߭O��Pcj����G�?ѱ���t�+���i��{�?Kk�j��2[�P���	v;�n��& �VL��W�ߛ/����.2jF���^T��9,�h�p��������"�>��;���Ьf�?�@�A%��[5{G�XC��,�.���=5ϧ�p rn¤�j����H>��N��-"����H��2ۗD��j+��a)E�ŉ�4�d[FfN)a����G
|���b�1����.�UA���^|�tuey�9Cj���5��rz��o/Ω�T������b�6j=����,��Ԧ�>pM"�0��7�{Mo��kh����R��`뾌ݣ�w�s�� d��%���N�K3�G�v�t�Cc1��kaҼ����]#Z�!��@���v�ma5�X��q�EM�M�[�- żR9�R�֟��טh!�Y���<�k���e��{ޭo�L���1�E���J�g�,H����)�Ҍ����5��GI�TVn	Y4�ީ���M�}jA���)�S[�Ґ�ℏ��'zp��R^���"��?�D��pa�ab��g�Us�*7o�ՙ��?��O8=H_�tx����(�M����&�p@�&����N���6ǍH�r�Pw�Ec	�ƶIX�z�G��gx��k�{.ԲJw�Xk�;|
�N;LI���h|[�L�*G�(z���>���q������q������ਐd����_Sd��r%�|qC#	�ЦɜӨb�*����b3]�DI����� ��f�\E� �t��a�U��-�8m߂�}u��l�4M�$�S����U��g���ڡ�[}~����)�7�
u�U�Rl��փ�z+U�kJV��-^|�MڍV_�a�c�e�,��9�_��	66 �Fv�k��@3j�)ʷ�-x��C���e0��"�۬kf���0Vwt�"�����+�&��囁eky�Rm�H���<f^�{4����b�#�z���r����"��k��C�u�?(�>�#ȫV\�[3��v���a
-\�9$o�`�!:����.'H��񚥭���4n͆�h���Y����%@p�'R�L�~!�o}���\����	&�����|�z�H�89u��mؔp���w|6�q�eV�(g)�}��^5�<*�����bi���#J�H��h)$�OIk��V�UK�7��g�����S_>����3'NBo�R����&�$ȏ.���Q�Z��O�":SU��/:��O����1u�p�I�������+��h�9��:ÝE/�M�~���U^)T�iƿZ�K�ea�u3wGcTh{Z�tz�S���S���@�}og��H����\��3)N%�oEP���q�®8���QM����a*x`h:�P�9�BN��1>�G�7�5�0�R�0�?�E�@<Π0�gv�Sm��繚O�U�5m��'�%(�wHD�g�,@��ʘ~O�N=�8��;��B�ߎJ����-x�O�*��#QP�8N�?��ɴwu���^��#-6�M�Tcƙ�̶^G��ő*N�ɱ�w��\@����7������e�+�b�Y}p�$���8��HC��B�ֽS�\)w,�[��F������j��9q���0��Wk���c8�P���-�ϫ1X=���7_nCg%��KǷ/���;�`4c���Ϧ̲��$n�e�t���y@E�����l�!,��	�&�9=�F!i��ϰ�
)��Wr�������cۢE��(����o54 �1�H\��+����yM��V��1�?��f��|��D�Y.[�E93�S�Mc�u�8N�����cp}�X������#��1f���!d-����f�kI���n`Su,�GƐ�cn�R�钜K�a���_�H5ԇ�]� 9��/L��j1� +�cr����P&��������b䳭6ۧ.]#��)����b ���9��1��(*��n�0׋_Y����3h�8������a�>�H�0�SD����?9^+2����%;�B�.e��B�
���YtM%]�a�`9�E�$L7t�W�o����뷯)��-1>�� ��{M��c~�y�xR��+��P��I����g�	@�h�)x��E���!%�����Tsu�f��h������a�Y�7�Y�s5|�+�4�)�a��%5��ΰ.h���3z����pz��>bx��0S�$��˴y��L�����z�M8���W�����Qlvj�LikuPڌ�ܩk+ٕ��ۃ�\H���xk�:T�+�\�^�N�^��uD M����J5T���(���
��"R�
H]�RsIᏅ	u�I�]0��}�p��b��گ;���t�n��#�����6�\�,kf{�N*Ԣv̢�� �\�T{Qq+���b����^�hS��D�g~	�8ף�����+�{r�G���Lk@m���y���]o�^���?s�u858[��z>�(M�����Ӣ$Zi]�2;���w�P�rY]��Ի���S
�6" ~~*I����{`؃���1��e����/ɿ(��a�n�6A���|r@G���jL���p��R��}����5�l^��rd��!�Y�5
5�'�"PN����ˊ��=����PAy|ϳ��@�!�K�#��5c�9�b��?�o5�p�E��D9(����y�[�m�xV��S�I �g�&a�Hv�2��PkX�N����_6��1�|��w��.�?��RUF��f�Ѕ�5��X��c�#6��IG�	�]c�g��7��y&ցH��?�y�?r��L��{D6P{�e5ޡ��wUX��e��(�mKV��:��N#�.ٌ�*�F� �ǺІ��HKIxQ���|�O�(OIJ�M���z��Ļ�ر�����d��3 ���ą��}�Z^iNU��2�dh��^j}�|u,��+j�z"�:��? �d�/�+�b�5���=ǯ ����cO�&\����"2�i����m�7 �_ב�H�][�˶�����,N���Χ�=�N����9X� ]2̎�UA�jF`I�<q]���L�
��[YG�Ӫ��ӕ}�.�d��l�+�D���0L����דyJw��9-GA�F�0%���;bü��}���}�_��V�'�.��@��3��I/����O���]�6
[[���S�/%���?����,��L:���	�b�r�n��#�?7����� � Pl�]K2��@6���C��&��ˉ ϟc���#<���a��<mX���܋��3�_y;o�$X�EP�c�o�ȗv)Y[*Qp-�,�Fp��������/
j�;sѪ׸'��7��I�#:�E��_�����3�>qZH��v+W��OP�d%����G�P.��G Ut��I!�)�;�dõGלIX�q��T�K�����l�1���{�2k.�#�չpӔ����~�˿H�yo�U��q����o#4�O1�e���)k�о�=��Ҷ���DgS��ǵ�t-m1��h�c��T�N�T��?Z3w׾�]G�b����©�Z�L)(N ��W	a8Q-':	Y���NE�S3������$kF�\	�H�@B������3/�K�	S��uߤ�m��wC�:'H؏��E�@��+�L��]�">�m� �8�W��մ�V��k6s�
���iY�*�k�wMrz��a�9k�P���/�(ڈ�����Alo�u�XU��(��췭�ۃ�%��x'�GMDC��L��F��#ڠv?��8Va��^���ʹ���UjF?!�,*�΋�8$�H\������A4�V P;/|�>� ���~F���X����������������bռF$�L�uy���,`:�
Lk���G���]����x{�����T#õR+�T���>h�:%��ձ���w���}�D��᱒0a�����O�WN��b�S��M��h�\`		�-ܪ0�����	��sw��O]Fn]�7������;��9���+�#{y�':.]�s�t�������T�%,���%�u��U./�X�l,b1�<��MY+oŅn���waX|'D��{�[(L����y�50"J8Y��QX�S���-�'kZ�-�/oߑ�i�0�_G3���~�W�,���c!��=�K�_��v�oa�* >9�M���Mp��J�7��'��:
؊[4�ql��@h��H�G΀��`K�g��p~���w�m�"ɈO�j��|
�=����:"��,���&�[V�>��b+�l��ٽM8��iy��
��s6J0����"�m�s���ݡ2~���ُ���D;��e��'qr蛠ªyb��o��:����&-˙�>h��c�A�5,e�p���&�H�����
v����!h��$9U�MQN3��B��u�������Z�뜳�5s��NC��R׉��ǂg�n��-�=��>��������}�{�b ��sy�P>�� �YOףA]��<x�gYNz��,&:�6�̜0�7�+�#SZ��D���%�:[w�c /*G3e �����PP�!j%*B$�]*KҽJƩ�����~�-1gsޛ1�G�~�/*~F#�����~���/*H&57�_�S�{s�J��s� ��Ř��wi��}���C���*㖭eFx���,(ܒe�F�ۘ�S�#{su��ۉp-L���^�]�t1�%��I�g���g�Z�Y�I~�ܗ}��<GE4J�v)�O����qUi�ܬ�w��r]����_��S�1`B�����ݔ�.��dh=��Ӓ�r%��[�9׵ȡ�2}��|�an��ϝ#���f
��x6�U* �ekz&迥��&p����mN��}�F����3�T���1��ŷ[K��{�U��/C�A���2��^����7�S���9�&�]ˠ�|b�|�ސ6AB �a�ܸ�/	�qs���2��%B?'s�{�)��$�����08�>��"����kq�|-UӋ|� �6�4q���z �ҫ���韋OvNg�A"0�r�(�0�H"�������^3��pypyІ�c�Z�E�>OHVtY&�\������5Չ��tK�0_^a:�l�~�Ym��
V�6�I�'���Nve!��O}���M��髈��w�Θ,gpԟ�U<��GC��dc��g،m�}�J��u�Y�R�m��X�i{+��wL� �a�&��A�0�Y�d9*�ɣT� i*ķI�;�_��U���tv�D�w�3�Cr�⣉b�Kށ�l�@�Ǩ�<�=�\��,�`���р�҉#R7G1�Ӌ���xCD7X-/�`B&q��m�"~B�K��_��̏���y9��<>3�WM�&�-���k�p�H�O���A ���	:����|�P�+�7f^R�`,t�������q�-߅W��=*CϒA@��H��6Z��6�1^�Zʓ0O�K��f��ܧ�pum-d"�Iy��.�W��C��g*<r�#�Q�+7��)�=��и�4�J:��9��g�sq�v�D�A�-h�)��y�Ē�X�0U������&&�p���-������.��l9I�r��%"�mΝ�l�bs��Ȱk��3G�7,�/M^� ��w�Ӄy�[6-�^z� )SF�υy�yՏ\!F�$}z!bJm��W�h1�!��G����,�~�j�bz���rB��?�������<m����5m7�4�]`^u`$-��\���kB+F��ڂ!��Q�ɣ���r�Ћ�av��zp��rc��vI9c؉@ B�#����86T���P��IR/��������@5���$�|��r~��E��Eݜj�v���ud:T(-�/q��uzBTFU���:�Q��l�-�o�u�a�Z7{����-p=ke�F���N���*���^�v�5Ԣ>�8m��s�\:;�;ΕS��ɆU���V�c�N�gQ�8��^;2�.��ϴ�*Rv�� �������2��8��Z�
���V�PWW>���*��8�%��f]�ָ�R���+G��0��G��(�+V^:�k������W�Pi���f
��,h�w� ��˾O�m"�^�+lzg�A�ǐ���_c���zE6�$�g7��\h$��,3��ʂ~�r�NK1����O�gAP��5 �ٯ��:�s)�0��l=�ݥ��ҩW�4w��`]�Y͐E������gժu�<���g��<ob9l�NWr/*��/3�%�m$�s3d&囫+Z��d�m�\/���-����)�J�q�PW��K=����H;�5�1������S!}W�;o���"3&Z7�����!FJ2����T�Ϸ-/?�~�P���b�Zq}���U�P@�q��o#�Va�r_3���O}%������t]f����|�r$<��Ս�;Ԭ6t�7�;���T��]ք��0%��)��ʥ����2�Y�����F��)�2�,,��hF�·0�������} ���A�3��pz���O�m�>�P�p &3KE N�MN+W�hR+�Z��灻���~h�8V��b��$�d�ԅC���A-������ӥiC��+�s��sl�" -��檢@%T
+]w��Jfw�E�N��
��@7�(�lV�_�1^�v#���xB֍��ȓ����I��:�c?*:[���l�Ѐ$feX�Le��g�]��S�@]!�T�i���*���z����N`DR
i`�(�&��֩�ڂ�k5����t�3Y�|fD�%m[�X��_
�I.�����|�<�elX�&�v8�S��R32��^h��˰(�$�F�k(:�7�O��Bl�'6����~^]�wM>Sjq��\y�)�G�9���c�cȬ$t)�/M3�d��N;��_HȪ�z�`�����?'N`�*��@��+o��a��c�*φ���a~E�I/��H� �̲�X�2�;���`���W[Y���T�����Ǭ����\�{{�!t;���CQ�_(�Z��z��{���v��[GIm��Z���|�-	���!t#̕�D��ԑv������e�)��*ofi:��"����u���<n<.���Rs\���BQ�c��L��ټ��ă�	zO<�\�y��R�Z����쎱k�?��Ԣv.�}�`^�e��<0����[�a1->����f�[r�wc�,C X�ė
XT��b���놷��ͼ_0B��|cM�Nb=.L�ٸ��6�<��r�b�E�
ϛZ8����"�3j����꺁;~��~�����5�R�%�H�ڪӕI���8˷t�ΡKi�,�y�C�n=��X~���Q����Y;n�%�F�@��E�$p��tJ>C��.��ޤ0�H�5HєFy`)���R�ש�~�#�&w^�H��>�:	boNuy��oT�+�U�"��sm���{�A�S��'G`�S	=\%��P,����'دb�j��f�܏�8��`�
=�+��	�kֈ
Qqp�b�`V����ڜ��l;_��&��W���$��I��r q�&��@:�}	(gLAr
fK{�/>QcK�k�=�WF:�n�����!-!��
��Sʋ�(�է��y&�71ԁ ���b�R���6�;,�.+������Ar�]l���1��q���<��b�Y�}�|�#=SŐ���޸��8v�x'_d��M����'�<�����X�W�I8�poJ��B	��ް޾��̧�?�ؠ]
��yC�sl�y�e�5�h�R��l-I��ot�!�����r�lᝑ�^�>����]D�,/�C�d۫ˢ>���&�ZR��6¯�Ϙ��&�Ac��?�^�b��'��eJ���RJl]wK�\�� ��|`b�D�=I�#�fTīE��Fa�m���%�B)���Ë}�%���� L��hZ�^0*���	���֏���ů�,W3e`= ��1`��RW�`б;zAz��Vd{��Ѹ��9)6q_Uh��;
9�{Nvv�ީA�*������dֲ�Bkr:�����������	(��X��AQ����B����O��Zh,����$h����߬��-�5�jG�ב���q���_��MR��,�����Ґ���X1��!\�] ^&�Hx��'$����AYmc�D���>LP]N��^fm�d�XQ�W.+��I�Q#s�bPp�*�_
�������U]e|<e%�Կ�&0I�s��<������N"X��o�����k�t��@+�
�ɐ�xѦ�<�V�x��~������+�D?��n��2�/�sJL��d�������Vw�w�(�Y�L��Ѿ	8��{�ؘy4䢗��#xD�e`�Ts�#$y�6vƾo���-��9�+�/%�f�&�<C�]���
�0����
�0���d)�6�#���g���ϐI���itV��7=D�v�d��:~�B��I>�:�N$�q���ßw�>����:�k���=7j�t��E���O� �Ռ:��5p��C���{�Z�Uqk)��RY'G�\96b	�Ja���Qה6�&���+�򙯶�lkI����(zAF���6JT��J�����&l�-@�py�%�^����D팈Dʉ���Wk��i0	9gU���{�_5,���qp�&�߂P����],Z��I�� �twS��L�{�u�|�a�d��ַ�EÒ�K��7��T���W�ֿw+wh;a�1Y�0�`8+�ɉ�{S�k�=?���7]��E��svS�&`0�QP�~���µ��8��̌J8������9Fܳռ4%�<�7�������Z	��LVg���7�J��۫����L�$*e|�ҭ�Ɠ�d���p�ƕx�u?9�c3裐܋\*ҹ�Af,Xde>`��ْ������y ���&dN�I3��V�МD�I7��D���x�S�tK�]&�(�Q	>碮X;��n�BǪ�T:;�.��,�����p87s�WF�jp!�x����6L�C���Ǥe��J��.�0������4}���y�ȟ:��E"�D��f������J��3�J�n����si�{�����S�6�H�Z5�m�a[r�I�@�����@���\Z�e�{�h�W���t� �����3�5�H���n����{
l�Ⱦ��O���p�j%��v�$]�'�3wM�?.�Ν�L �'S��Je���%YO�F�4&H̃T�*���pODd�A��l�7��X�5J�HŅ�k3��W�P_9«���ತ�"�Y�=I�@h˙�YY�+ZS�]N�u��^��Ԭ�_�Be�9n��ꀤ�ynTc^��#�6A�4Y�o���T=f�a/��H�*%5���o��y�K�J�D��W}'�Ƀ3�����+��&(	6�9CK�p/�أ����A�H{߽,]M�*��Ze��'���׻�{�_z��,�(D�-=c�Ncjqq9t��4�I#f�V��`�N�9�a��W��7�$�l�*�?5�5sk��1o�~W󩤤�/#l*藕���?~z�=-�o�U(@z��2Fј�x	T�-	��l� [\�҇;���339J&	7i���B���G�D���k��p��)��B�-ވ���SHD.9Z�'�:C�K����w����f,���8���Y6���,�9&I�2tv�}�
L}%��QʘD{&vM/!�ԕ��qڤ֟>�q�u˩�A��l81�`��5�h�됚c ʨ×��P��Z���dwce�K�"�5�x<?6�^Ů�L=B<N��_��9���^���r0ʌ�^�7*�^����)�>��H��5�B6�������<�Oy���o�x�.u"q񷫷�q�u��l������z�m�*"E��g_��*E4{��B5j���]AR	p��c�|�n����n3�y��J�'@�я�d�@p�p'6����_A�\��Ȓ7ξGH�2$Úp�P��WîR��/RdJ���q��*P��������j�#0]tp�U�;�K�Ow���DP�r��uhdÏ�/VLI��;����W����1�������t�T�C��������Kqv`9�8��bߋT�c0�" �ymX��3�B���$��F�(e`o��)�q�oo�W�g�9�@ϼ��G�I�'��4p���U؈���S��
�0�
�s��gR����^�	9A��Y9_�E>� 8�S��߻�>jvgR��I<'��	(-�ڧ㿶T��"�A�i��A��/�Z�.-�sC�����
�A��_��:����c,�Af,��AU�*뾹���s�=o�v$Kn�v��ԥPB�ke�`w�kP���3�V��`���@
�`u�����?�1cN���B�
�V���m�IT���q�a�Lhn%b,�����:N�c�Q�W+��Gg��3�a>�_J	p���`���#�#��q��fZǷ�l,�C��s�.��F;|_?�X�*�[��k�aĔ��h�����k��s�5���>[�R�kY�2|`�N�Qh�����>���&P���$P�

��;���4o���GDZi֕�N ��������P-��Vܩ�`ӄ�5$�����Q��Lw�+@͒�z	y�QM��{������l���@բ���"�r��]��[��H�	[�C^�i�"����ڐHQn����\��Yv�9(���fM֡��"�ǜq����Y����oY7@�.�9�{�T��"���rr8aٓiqjh�W|�v�a'���w&��܃љ����#XY9��_[��+��8�Ð��J�/����� P,�C��o�	�	���W09s�0lҟ�O?m��02!Q��)T{`��v)���ڧ��u�%=,�J��C�FṆk������<$��t\g���	.�p�5��7��pҸ*	�x�UD��[-��_D�P֘K�>2�瓈�0�?|�URboAI��\��`?h�'o��\J������4e�H�q|�5zV��8�T;��%����^���D�K���t]�O �\��g��&{����"��|?\>ȳ��6����<��bUbM��`z#����@l���K�|�����)�T���$b��Qr��ia�&������2�i�E����~�&��۞���9P�s�/�-&x�G��1��_��"_���ӣC�2A��p�	LO��	�!d���: ��i=?���ѥ� XTv�[�R8pH�N���ҍ�����Yf��=f|�G��ߠ��QL��I��*О?ןZ��,*��0���7��<���gw��<������T�+إAzX�:}	-N�Q0�x=R@�-�o��~�W��Y�}`d���:��"�Oӯ��Ӳ>��l�/�7[>d;{��Y_�� Q��!,�U�S}�vO�t�v�� 2�_
�:>ݶ���lڜ>�6���aK�d�e �����e�-qu���8�>���
�y�e�!��2 96�G
�*��ۅ'�`$~�v4�(��Os��9Di�9H���P~h�Q|v����!�[����t��<�q�`�!���<,�2�X�7y!~hZȝ���@�Q�*t~f\��@5��/��4���W)���G��T�{s���Q���珈X�`���7���`b�YSl�4�]��*A��R��)�Z����j��R�t�g���n,
�YKn&�',������$fK@GX}?q�>�DL���Z.�ѼX�����c@WwB�����kyc���ERb�G�Z"��p���K���i�g�fz�v,wS��w��CO�pϔ!�س�牶т�1�y��?��ce�k7ԁ+��V�r|��G2a$d���i?&ǲ߇,��$6��l��X���A=�h>gf�Rg]_Y�m�|��;�f�|ö�-O �.�E  �������7<���U��<�l����U��!�`�hXck?��(�::��ޛ���/�2+ǲzߕ�aa���jLhŝN[Ɂ����'�����{o(���[a�i�(�̛y�X�_VYрH�'�I:F�C���|Yt.���̿�:peG�z+me��=��ʉ��%v�>�NF2_+�E�����lß���}{#��DHm�~��Ԏ ��k��0�4���ٱOǮ�w�v�c���G6�?�a:���U�J��@�d��l�AA@p����GG����=�c�Xp�-SՎ�BFօ��x.���/8Z��%���:���+
�T�6�Ә�4z?׷�^3�9|�GMз#�����[H�%tj ������5z���qc��`aȇ������ފ��w� �;E]�9�#�_�?�]VW*�;[��U6%�_�(z,|���� �bc�����WJ{i�~5�#��'�p�������/c	�~'x�Aߝ-����6�@����jﶘP�����T�՟�LIl�!�F>5!^�-��LK���⏂T �ݹy Ƞ���Vw�c�8�#vo�D�p,�*O�[�ǋGW���~(���v�ׅO^��֔;�}��
c��^��$��<�@��i19�)����Ǹ��Z`�<�wY�O�r�!�J�j�jh4��޾�!6����=<��ό�d6;/��pi>����a[�����ֽL�m�v<zw�A��_�)x�`ޚ��H�I�!��{	�� 9������6���fnς��|�ޑ}5�Q)�܅��KdԸ�5���������K���X��gI��\���APY��:�:���j�v�{�xn�]��1��B6��A��p����u��VCD����b�9�� }��I��C��A���O�B(�R\��Y�^�7Ä���G��)JZ͵�,�d���x��Q��2��b��
�{���@�#M�wSj
e�>ꡚlFPvY��,0��?�����@�>����Zf��jG�|���=��y�m���d#>�n>�pY�m����@�����A�v��S��U��o`�P�%�0T\�.72�:���F��S����2�K°�
�r�w�aCp�ȣ1 -��[��Ir»cNb�{�}��λ�qg.@m��9�B��Q��ߧ�L{����vaO��:�@?.GH�r��ۓ*��@�
�.q�|6��?����+*�bk5q�x���`�(�Վ����{T���%�q�ElQ�B����+\z��;����U�Q�����_�l�ɏޟ��{��$���:p�	�������Tz-��� �Pz�F~�N���wpEj�%�W>�X�&���{���;�x��p���j��4�.DK�+KFV�B]��1F/9�7���rKP'0.! o����&�%��u�^���&�WL������U1��,�KF��DVT�#9Y�����W?�7�+��X#�t��8��V�8�\,��?N����$qI�a��'Fp��O���K0�Yj�� �ɧ�A������ln��77&\�F��(����r���SZ��>��5t���iwn��8{{��$��i�D>���I���n��$���g<�e�����޵+��a�y6d�~$�bJn�C��}���*w>+u4�� ��"	*��H��%H�8v�	֍x�<d����vc�u:�N��GP����
c?����}��	�*��u�d�Ԡ�����Y��P��5~�����M�]%[�~���� W#�	����߲�&���I���>��G�z�&{�1{=��B�8�M���9��G낉�b�
�����ݭ:b��κ	x)@�[e��cӁ�UY�{�۷�x'wᒫA������}��Y�	�H�nⶠd��5���f�G�+�����Մ�g��?Ć�{�EfUeU�_8_ߕWl|K�%4����$�,��)g�ɮ�Zo%p��BfN��v�n2�H��?g�����J�^���iN҆aW:�3�^9M���d*G�-,A�+Vp,)������c�ii=�ͺة���,| E���?W}J."H�"��'#z��*���4�ad���8`�6�I�1J+���O��Yѣ���2������_?3]�*�~o"��}z4{4�Шe���U#���^ ��}�}k����G��a�nx�C,i�tZ�v�(���z��H���1��_7�������ӡMi���f����ܮ�#��+�M	М$%��D�� ���*g�IA�Q���>��=�ک��<<��q���&PJ����7�2I:��3��L>ˢ�v�s�4�Oz?�ԣB!�%�^[�E�ۥ��t �VR�rQ(C#E���8�<�� 	��&�M��]�q~QSZ+�]�U�#��b�l�ֽLs��w�VLLwɿ����C13풫Õ�^�o��SNv.�#*"+8S�L��5�� UN�JIo,�N�屖7��hH�vw�C"
,8�dCҥ��w��m5��5����ߠ%JI@��֩��7K�D��
���@�r���hw�bah�6�u7��Ш�zNFH��
�,�l����U��l|�m�@5p��n��J�Yp�m� �R?R*O`׬9�^��2f�4�P��$^��b�)+:��:X��$-���!%�sV.p1��>�4��Uqb�Kg��7�ufU����`?��ݘ�����8O����(��G;:ɗ� �͙�+E�D�mG-|޲K ��﨎P�N�9��ב���	05+��E�����+�r���B8u�1���.n�H��	M��a����i�p���Tyy�[�c�B��E0�~%q�d���Dl9��S��e#ȓ��aV�1�:A���Y�ܱ��L~�j�c%4`�?q݈u�Ly��<B��K�o�M�Zy�U���Ȕ�:��5�b�;����No|��9�|�k�E3=C?&#Ȓd�'��X��ȹ��^�� j��=��CO%Yj~���v*�cac�s��[���.Y�i~Vx'6q���d�R�OY, �/��/��ZZ�����l��'�!nA��I@�\Ӌ|8�	�.:����%�t��4�TX��G��B �,l F�^]���t� +lN��z,�PR�ǚI�D,�B����^"��^q�b�d��T��?1rg�EH�u�<�&��8�	�9���X��ݏ��B�DĠh���>Z�=q��6v�b]�2,`������I\��.FR�E�0�C���Y$����s���V�,=z�qd���K��044��Zr���Oފ�{�Z�X���̄��p���e�ٳ��'��f�@e^����iND�mޭ1c�<Ah��k�%�v`L�C���n�U��h1�Ov�=�,��S�S�B�xA��Lc�Z���7���c��ya#^�ʬ������6W������x/v-������m�`?EO8��Q`*�4fb�3v��~�ē]ױ��?�����y���w�:����~|�t�&��@.���������K�b/7�ރ�m3�1M*� [@4N{�L���Qـ@����UDdw�5�cߴ����*=�U�}�E��*���y���㺊pB�A*5�
jK*Ƌ�I�D�ۃ��GǊ]�:�0�<_��o��wzOr�?�6��&0ˊ4cRRy�#Vq����P*+Yl�a�ZO��z�W����
�fc���\�+��
�Z�K�Oxף}]8��dN�4^�?��k*�WqSMC�_\�T���������&Ń�hE�]��@�ϖDp���ǶK��~67t�QH4�Eԓ�٧�o�׶/Hv�%���g�g��\���T��S����̅��8�5.����1��Kt�:�:{���@��r��o���O�`��POAPF�Hs���aZ�C�2�s�Snv(��g.΅���x�.���TQB�Z���I�� ��
h�T��t�`5�A�GoA��)�zYhUfIJ{�ۮ=���X��b�����]�P����C�tl�mwQk Hs�k�9���/�\�W|�:�+{#Q����NG�y=�ǩ�.�ӗ��vBe�/S�,��L��o�_��H��P��v5$�X.����9d����L����n���]�!Y������G�
7@8��v��6H�����p�|S�����i�"ӷW����L�Ɋ�;:� 40�8�`�<���R�J���Bs����C]� �s� t�p���Fܛq'2��TԻ	{+qҤ��
�ڄ��T �s��mN�@V_�O�6������uR���a*I�R�	��ڂV>U���;� .W�U��U�����0EtG��{�ue~���9��rC]��f_�4���6��_|$������ѩ���6���J����{}�Hܯt�Tޫ�B�w���Y$���rf�t_GÉ����c�d ��u�qkUG]��|�'۠�.'X�D$C��R��$�f�-3�OK1�x��|d��Rnx�n>j=sY�
�1���&V��F}h��;��9�Y�e�Z�l�7�5����q�+9�eU �x-2�+V�4|o�%Z�ݺ�=��Y��[r�K��OLMYW�p��Z�hpbzeE������*�z���d6����-!��L�W����[nm��2�����,-�B� �R�h}�J2v���ޘfa��HŢS�k�yq�W
��rJs$[E[�=�>l���?�6��	:����?��CC3�ԭ2^4�d�p�m���}�w�@�H���UZdz�"�G��6����r��|
�Q�NO���4��*���}�VҚЇ��{K]O�T>!��~{���d�x�3hX��6��)x&�>+E���4�t5��*d�U�ӷ��4Y%쉧v�o�`�\�W�������3)�p�����
�1��4�';Z?��m������-%�t5ctyd6�N+IcH�㓉�لpW��q��&���4`����i�����?�)�	�)��}uc���'������þ��goJ*����k+;����'׳�έ���^�Q	��q@?8ќ0kٕ1l"�H,�-y�m	��c�{_�Հw�T9�����j���rgR�,��%���6�X�p�E�9OAZd��mmH����y���@����+F��Z\�Lr�'���9�tQ����$_di��YJX����[>Zd=֕��܁��J��>��ׄ^�4ђ��~9�&����~����7���h�Uϰ^VSd����%Dn!��ib*�%�be�n0h�В����p�;sTˁ�4�p�L�+d���m�k�L ��?��<Z��J��^1�Qn"^�������Z��v �b>�<�T�����:�u�$���N�����AAb����D-92SQ��!��K`���La\ݪG�t�һ>$vL츳��̝��B�1y8�[����}CLh�dk"��§+~F������$�1X-*��?�<,\� �t�Ag��M0 �y�	�w��L���lp^-ŕe�!u}~8��μJ�@w �&t�w���H�D:����ϗ�r���ˉ�_�+��Z���������fO+lh��R��E��ܤ<t�;J���}����>���QM�a�j[|��.�|�G��P���ǆvߍ1����˄�z/�.�>x�/fʭ���͍fy���dج���W��K[ﬁl?'U+���i�O4=���D$�p��$���+�p��E]�5��l��2�Y�)B����<c�ʖ���4�7z2"�b�4��/| +���<_��^z�
s����Չ�1ī=�[E]zbh��6�6�lwl ߹��|Lk�������s?�7(3�[��f�Hp�9Ł�H�o�Z1�+�����҅tQ8��.����?&ɚ�/������&�c���q�E�#�%���}/ژNk��Gr���g��V]+�H@f�v�u4��I<'MK'}hfFs�ox5s��}�`�7�C�Ҍib{�/2���!���_�A���U��x��G_�ϯ��_��Oj��շ�.T}��'3�"S4�$�Q�����Mt�����x8�-�#mO��[�z����:�3�����R�ۨ��x���u�����g%�� vg��7Q2ݎ��Ɍ��j}#��w���a�v�i�p���̍x���
A�paʍ�M"�w�UWG$�}c��;�Y7��J��Dt<�~tk�u�҄���6zu�UB+� �v��%{�듀�-��|E��#9!� �}�Tp�13 >�Rdh����UNI�)�	5f��~7SB�a�5�5�/|qy!�o�m#cȣY�;�R�	3m����tʥkp�Z�z���s�쒑����2��ڣQ�s�#g�7�;9܀^ō#���,Sӫ|�3p���DS�>?+����ζ	�E����R��6�x�n{h2�E'hq3^�	�ЅR/g�	�(�7M��.���@��!��V���&�� ��e�='�U]1U�&Lk���O��f;��_��"�]�*&k�\�����yZ�e��F\�ܹ��o�М	#��+g?Y!â��̓K" ����j�f5�J���D;�/0����"��0��4�~1�̐�Ot?:�����e�ejm�n�Zs��K&�EH��7��P^����e��&ڕP)v�6��B���>iDo��x!�w�S��;ԓ��Û�HF�Z<q)�:J�M�D���q8��	_r�����T��^�~#���m
o���/b��:D�7��\�QMfP�Wi?��	�C�0�W$�R�c���OD�I�[e���3������2�|4@��b,D��N��1F�ʏ9�f|��@��hc��T�� ��R�;���q�)oZ`�ә+۩G�`�ͳ��S!���;5]�%rJ��x�r��ޟBr]5�\�-���`A�����Q0�,(����)㛓�`�z���odc��Rx�R�8এ[�}m~A���Pq#�n���s�$l���d���n����
Օ7w募AOĎc�[5J�D=�춛[����_�Ǎ��9#�>()q�B.�g% 3�Q�Bb��Ua�����&�5���-��)��9���Or��i�]/�ݳ_kH*� ����Yn�p�ӝ��߾(��aLՌ�ت}iP�a'�����z�U6��Ff�ԪZ��Ǉ�^�#��3%5�$D�Z����l��3�!�Q:��^�M��@���En ��V��������R��\[�h���QLX袭�MƟ"��x�i4�v�K�`;�����D bU����+N�p���%9b$�� �i�_A�-P@� �Y���/���]�^���%Gh���0vЋ�I��$'�?+�>�O�M1O4Ú<bA9�4L�}CyM���!��٠|~�Y���>?��M��+q�+/��[��_ޥD��`ӣ���'��H~X�z���g+�N�jh�Ua 1X���A#���W߳��o}5�:"�-m�i���_KK�q\+������1\���^F����j��O_J���;�c��t�^&n�P��(��>�BÝ�#�cja��1��tc[��h�|D�6�-���V+|�8�"�$D����2E�[ݭ�m5Ӈ��UTCK@J9z���?f������$�G��=��J��.e	[�7� ��enz�gW������k�Ϯ��KD�HZ�-9\�3s�TX�Vw��>�����$�82BNj*�婰گ�M����
`��1VX��n��=�z�	��/9�ih]�Pb{�T���YhlX�̹gr��SC�?�|�>�j� D�*�<�N��a�Cd�����(8 t�2���.�Պ~��S����}j����HŪ4Dc&��ޓ)j/WSM�=��8Bo�|��watUQ@�K����/��U(��ҍ��4��Yȸ8�;�*�eyWZ�
�[n2�Y���N�H��:̅_c��R�B �� @��[���Z ��7�d�B�8T W�"�ijgG|�*�Ǭ>�Fs(�a�f�mt�$ �Fӱ<#�������Vy�Y��.�s]���b�9C^@��H�61���{�0�܏v=9���Ȇ��f	��"��s˦A�FV��6Ƀ��}e��ѓ"�d�/��Lє�����Yи5	��5y[��|U6de�J�P��g��
E�M};zH#ww�b����i\'�7ص$z�?��|`�� ������?^�dPej�ZI2�I/1���:vQ`�o�����"��Ba �#���<�t�l��kv�
�6��P�~�.�]Ml��<���M��)p�����a���ҁ��%��NvP���~H{;(��r,���a5�B�����(�n��R�b�L^�W�ӕ��F<բ�6�!M&iVd ��"����]p�oy~��M�n\�y#K���sM�z��L̬�<�s.{����}����U�*ed������K��E��܍�>�b=fH{n��/Ha�^��kT�kG��MeHL,��~�|��?�OT�;���8�~U}�����-r��:ikJ���U\��ISH�'��ڍ` ��~�d#�0�UR<��/�P.&��1���� �|LH>��/�.�^����S�.�V�JeX�ey`���� ��ĉ	�m�M��+��rG3�Q���)b���u��_��B���T�9�&�V���w�I���u��iP>�7���)��O�S�pcH��4�<ƿ31A@�w"�q犪�B �l����ec�}0ħ)�Fl�7[�X.Xol�kr��o ��gL������Nl5��O�(��9���y���gXZ��MNiߋ#3�rY�W��n�X��C'W���M,�8�':��g���f`���'�\a�A��ٍ���2�����Ч�W��.�rn(��pPZ�%4��Wb��,L���<�$��,܅;�:����N���kSv`gpP��r"�pVP�Mx'0%-�<P�c�$���2���tiV���mk>.�8h5owh<��Y�k�)���~�,�}Q�1�q셒l�n\�ӻ��T�v)�{ۿ����bK����c�J͸��.�v�2�BC@��!��D5oV���i8��{g�J"mv$���ũ��T�����܌���xհm�|Q�%-r����½���پ�%J'��"+	ʎ���I��?��>�; �Ҕ����Ml�6v����R��T&�љ��ޫ4��/|�*�Ӑ��|T�E�L��lI����$Z�4���x	�����3�:�b�PXpqL��m��������(�-��e��U��Y��f�93_��8�䳰�k��	 �y,���z�x�/Sά ��o����?�@tv'c-~�t2�ŵ��$8�L��K��
�Sg[m���x{ (_k�U5�L�El ��$����i�܍���Ÿ|��"����'z��\������T��2��>���tb D��xC%��l����7�6������Q�.��D���%�{>�A�BY?��H|>SR�\���~7�y�n6�_�xч�b&�-����%w,�歞,.�� �
���]`�M��3�&RS�L���B|��S��	xܤ-�)�̤&>*u"`��>(�Yܓ@Y�u)�����)�">��"QxY��!R�M�R�x��I��Knō��eϢ�n�J�E*�篺<�,��	�8�����h?Νi�^-[�^ �Yk�d/M�2O/�����X��r?XS`�G�Ә4D��J��ɫ?p�����5ͣE ���1�U�~���/^��xIQ��B$�թ��$Ҙ��qn��2p�/��M�����afom?%)>K*�X�ρn$���2���KTO�����B̏�t�G��Rـ.�P���KU���^�Z<c�K�\��<��<���m5��#T�_�l٤X}u��[\�L]�Ǣ1�pc�X��Ⱦ�Fi�$H(�8����X3ݯ�<�E���ǰI��4�$� �[3�k?����^��.�I��X�#T!538X���8i��AbMM�Il9��	�E�p7n��Sr>��x�>���@w�K�H�������1O�@�����ü^��E�Z�.@c61��$syX�9di9�b�X�5�ɕy��T��d4���眲Ѻ���.��+%�iD��-�F�[�3��93�p[��k�k�B{QF4��`�4�{uC��2q󲜪�=E��������ӏ��]֢�'���)s����)�I|����|�A����?-��>�sF$i�yr9�Q�gV���O |��DE�OC���;�����n��?5�<E�H��>���d{�Y����`�;x���3��wN�SE�#8�h�Y$>�v:���{C⇇7kz�A7]�ڱ�)���ak>�@��F���D+���)Av��+ƏV��!ig���T+��W�����5��p�t1)g����F 1�IF��ȝ�
��m���m���seV�ane`p��ԣ�]����=��RY�o`�7`����w��s�
M�hl��/)�!��qz=����[Lb���"=Ή�<W#e�XnY;�,y\l��f��-���߃E:3��Ԣ(S�dL]Ǆjl?ZI*��E{�R����]����U�\+U~�;�u��F-@nv�	�)���&o�6y��W�t\P*��m�%�6ڮ7�f3M}V����������k��a&�����&����8�:��8+v~A�پ]��f�����eۉ���O<'|k��t'�䓤ȡX���&]9��U:>�Ec�Y�G����!k5Ĺ��B�\��b��|�bv��Ĝ=���3�gDf���g��Z������khXx3��/3�1�%aQ �">�}��1e�m�{�A��i~��հ�Z�c���d6@�O�Y�z���YX�s$�aA:��T�~�֡6��|�siWg)
��,�2���%��}�/�?��V��GP-יJ��~v�k�~�̊V�%gIј��� �Y�2��R:�q���BQ4�D6q�q�0��hL7t� ����bY�~x�����\�N5�>�e\�j�����p�����F�PQ����r�t����
<+G�4�s�� ��/���>`�y�I��=�d4�۔N~Cm�d�
yqo�b�|���q��m�
�J�S�H��#Ȣ|Љ{G����ۮ��t=�%uU�P,/���i�׈�Vx�%����Έ��m���|��2~�PNY����d��VҨ����'6=������B�M�����@&}Y�\� �<T!V�Ycu@\u%�@3=
�rF%J���ޔ��)���-j��{���@��j �}X=)��')r��.
n�u��`U��ˌ����\s��25����y2JHH�L��Q�R�q2��n*�iP����q\�d�#e�X$۾�cf0��)Z�Oށs���3۩�+���Xǎf;m�X�!�Β���ʮ#�@J�q��k4���)ZS#t����Y�"?%9]:�G���K1��p�����jc���Fjh��FL��9nf��#����&���{t�H�� �xxu9���VW�|�csw�3��08i��,�@6i0�|�|��|+�hhG��Y��4Z-���mS�O�x��@J)�D��\l��U� R[�b{u_��
�Xk������M�Zm�7�fI����}Kz)R�Z�ܴ��kV��)��9|��d��3����*����=Ek�%Jx[>]�/�
����A�'2Jh�hxu��B �����h������R���΀�م4 �h����v.�zm(6�P��o{�֦��%�����9���m�*�3sX}6�<��`*��+�>�~�֨��DH�$��o���h��<����%���B0qC�Ӑo�˓����\|D��(0����@0����e�"�0#�|T��1���	ka��&�ݻ�0<�2��A�(X��X�D{�aנ2���~�u���xSN|�AK��ٱaE�Sh�)#�o�!��Vpo��°ˇb��D�{�>�ϒ`�����+lј�4�%����>�:O-�x�+��ܤ��AKv?8�b7�8�/�y��y���4\qnu��EDB ��WL��I�9Lj��c����7P�=b��Ǐ=�$�se��J�[��zÅz�`�*j�m����=�X���~in���PjP�W�s������N�f�|�Y	��k�e(���'=`$���1N�{U�z阿�F�42hN�Ư?�61��A^b)�G̏���`U�p����+P/[�>�y������YM�3�ZF�ѷ|��������s�Ԙڼ�Fk+9(�n�g��|$5g�a�J:�R���G��md�Oa1��ەsqq��_dbp���A��k�X���_�{'ɤ�� �r$r�+���cj������׿=ʍ���C&��4���1(f�Q�-�YA�j�W������[�\X޼��h�"�q�!�-�\���X~_�h���Pzԡ�6�����zG�;��@W���i�D�X�P�a�K1��ޖe�����+5Î�2������V�ʄ���ԠW��R c'���[������x���c�q�$;s3� a�Ď8Q{�>N��+_�R������n�-K^�G���8u:
���u�?�N�����'���{Gz�V�ި�Ɏ}�� R��E�Ac]���{���b�X���$橍���	gB䏲����&s��Tí�g�� +�*8�8MU��J��Jꭿ�� 3.Њ&�Z_���b�e�<�2��{��+���!8n�E�hֹG� �b���͍�,�R2�����tv�8P���p�	f�bKK��3NQ,0Cc��z��H��`������b��Ґ����b-�V��s�}�Т2%���M��9QQ�\���ݿ/s^��={ec�9��F\X��}4IM��4�j[ٽ�h�P�1[�+���}������R284RZskR7A7c��������36��9�ִ��Q��J� c������mq{Z�s�a����I؃E� ��&�`�R�ʄS��0��h^���L=�4ϖ����@P�@��k��<J#�=��P�ޜP�A	�J�����-�*I��x#�ߟ ��
Թh�a�(p�gТ�-��k{P�u#)��
�>��|ۜ~�©��U~)/c��U]d���EI|��O�~�9���Pe�n�2H�5�B@a���e�=(%˭)H�Es���� s�2�d���:K.�$E�~Zl9ڧ�J�4��K�����7%��5�pB;�6ۮ�z�������7�e�G�0���À�H�
�����	�|��T�u����z̢�%��I|n����/�{�S�A�2K��m�%��e�7�7����q��{d�9�(���	 ��NJ�;����e���W�^�5�6c�5���ˠF
�(�L�Z���1vY0m���8͙v��P�]�9��{x=���hRtX�"F�� S�ԙ[���TU��>�_iZ��Ҭ�4K�Jq#�|`~�������O^�m6��
�Ȓ���;�wEI���-�^TU����z�3�+��ۻ���)X�0b�o#Epz�P|f���o��S/r
�L=���X��#��Z�� ����sc+��S �c�S�FwXC�]��s��	�N ]T1�Q�N�IA$+�����`�A��Utf4��_3��$��_	7�@��?c���������#2w`�-5�R9�m;<z���\�hQ|u�Q���q�_v��g��+u��9�� �_��� �����'��2�y��~#|�z��jA$�59��*��& �8.�	ð�t_tɖ-�ʁ�Ɂ�MGN5y��?�ܙ�Y�;�2���� Y�P<v�3�R9|�1#0���%��0P���0ſ*"S봨9.�rER�)u����k�_`��k�k ּ�#�� ������Kk�&� ��2��m�@o%������2�<m��0��'62����wS=�Ϫ�lk��Q1ꥋ0�����m��;�b����~d�>6�8�E�E�}�kȷ����'��8/df�:��3��
�t�:�M���ҽ�4M��")q��gк+"ohpo�+YZ���{�uB�Ԋ5db8e݇�U��5�?_�����PhD�7[�`�w�n�"s���ObH-�퇶5�	U�v钽�f�G����_nhk85��VK�,n�]$X�
b*bd!  ���I����a�9̷�m��F���y>��|����v���M�쇄�}F��tiY%��V��T8m]�.t5��0��F�� !w�@В�_�ap�z�`���ciCN�êǰ}ܕ�T[�%���`������
�V�wU����'��`����i�U#*�c�B�u@ ��80��@xB�+I8�W{u�攦�c����I����P�9�m�Q�=ۅ�rE�����甥S�2��)�<��ΐj��l�,��/�tn�)�jA
���K[z_��P���Z=�2+�!�AN����k��ݤ�
��Î�c�`�����5m".����:�V2MbE���I���O�+�!��Sm��J�1%=�皁�A��W��x�@���q�*���QR>�̓18����dQHޏ�����ن�y�����*#���}�n��ᩕ�[%�q�(�؅ikk���J��x�d����|�!8"U&T>�"'�d�ȹ��� �pFVEd�v]���H�+a��dk�\2�<����mUv�M�V�8'%U�Y�`l�7ʶ�/"+�����!���Rр��4���Z�5u�P�9ͧ���w��c{�#˂����*Q4���}
-C�j�Y�sޕ�Z�~�ANz�kv$*ް+F`����X¤��n�yO(�c�  ���pT˓�����Qĳ:���ۂ�G�K�fC���~o���r�h� _x.���c��|�b;�aV�K���k�	Oث��u�nYz��?�S�OV1"��VĤ�K�mߜ��hʙ�N����?����k�!��(ux�ho��]�@
mrk��"��.O]�-�:�H��`�!7NR�A���l����ir#]T�3��Q�~A��Q�U��wy[�NF��l�=Xɭ�+D�+L��y��M=D1vǶ=P6ù��g�e��5y#��W���h�<�UX\�%?�����Uz��1R�Ze���,G�$��ptU!GaRɭ[�B4� i90H&�w�rkw���L��lj��輄��Ol�t�'Hf���w��� zI�;"�.w��Щ����MԤ���]XPѽ�5�̐�GI��L��	�j�J�/��.�GrVk��gg247K�²��u�ē��7�����RbFF���g���|o|�R������5͟�	u�Q
6�O������ؤ-���Rz�V( �D<;C��[�3�k�!����_U���)��'V�@߫��g��iX�K\R��)�3HOY�`s�1XS��73�Yᰳ=#wnM�:ȸ���}��Ȼ7<���.����fZjK�.���?�s�iJe^���
���!����&:2#�4A�A�N���y�-F�?~1�G�`�kh��`�E|��b#��HHB����Ui�����oe'է<�R�/e����.��w7A�z4#��tI.���d4�=|@zTG�p�����\���c����Jkte��#�5	���b�dC��pM�w~Q�s�vP%�gF?�Ջ�ٙ�<�.`�uKD=��z��  ��CF7C�n9�%�'������,3og%�㛁��~U0�r������%������I� ���mI���Og��r))'&RM���L��9�\��z��}�1Qh��|L�6A��]C*Q���r%�e��Y��^eUgn�)(>���?�jW�q#��(Sh���`��t�R��.Y��q��`�O}n+{��ZmS�A-��Z*���Pm����?�������w�k�|c$ȏ�n�z-���a��_<��>A#��۞!�� dJ�v8�1L�ŕ�[Q|�G�a.���	�V�K�_��.��<�a�|Õk���k#�f��5ҕ���l��	��5@��I�-c�����9|m���&��ɳ�d�G���U3�,f�R30T�| G�&D-j�����4%ORF_�+���f�y�S2�\*�Y�u3"�	 "]_��͈K�ze���?P����Ā9�F�ٿN�T����M#8[�c�̔��u����	����JY�	O��|�R)��?rс��L"�����bZ�iUJ@ʝ����둕���;v Fc�H��2jc�X�O��;v�j�K�\5����T�븪�}��V�A�]��'�S^k�ޤ�������9�7�,<��p[5�j���";Ll�G7�U��o���9ѧ7.��Z�j�{�-#�T
�0�K�|�
b��*�J.ɴ��c��2�17~z�,�k�iB�<�{W�PHd�5ѯn�)���<!��_�̱��M���[��߿�ao�M��P��G,;�)^>�EQWl��L�a��*�դn"_�˜���c�{�M��I��(�v�Lhg���F ���:*\���� �ZR�^zc�������MI��N�FTzN������� ��t����jڮ�B�-h���P͆\�]�=ܠJ��A�My��0��4 �T��yC�5d,݄�M�:b��0r_����!$6�d}r���;��XZހ�U�"�J�=��<�+�=�ˀtg��5(D�{G������R�c�׶�v�N�aV�6x=�MBW\�G~�FA #�G.��X��r���^&]��MBD������mB}a�M:�Y��3p��cJ7����Ñ9ˉ��	D�_LS2}��#�xV���x�=KJ��[�B�	;� ��3!R�j��a曧f!�.�,��l�B#:@9'��DH��߂rp�ƥ�?�N���ݢy��J㳎�����K���~�[!��/�U��� Ai����3�X���IF�~��Cd�����wZC��.�{���.O:����
��4!m�ڊ���D�
�A�z���U�@g��{��) Ĵw�u�_���l@�h/��kw�������]x��'�x{߰cۛ�|#˅���Mghkd �W�҉li��1��		��G��2�r5,��T�]!w�Zlr�^������=�_3��ǣ��>.�磚��w���ډ�E_�ƿ8L�Xt��8_����]��WO�U_�e�}f������\����],��0!φ���������Tޕ�8u�w����J�aC�EVC�������u~�����$�X�uΑĲ�@��j�F��t"�:F�R���ɔ�bR����7qj�j���R�Kz��pF����6����8�9���1�ݐp"���R��#6��F�����,9H��En��R�	�mBI��d�}����Y�v�]ۺ�����YO�������.�W�<4��<���T?l��=s�a7f�*1Tn�����d/x��������`5����KbP����erT˘lq)`?�!���,���Z�YJVs��b��己1��1��]�SrWV;�A&�ގ�=���� ���q��SH���ʠ������f ��/����\��)�T�V1Ő��4ӄ�1E�����1!�B���\�N�U��.�ݼ��e�I-��D��i���!d�%�����e�`q��� ��= �?�K��	�lHԐ��5y�@� (*�/�� E���B0��vRF�[*�sU�{��*�:�F7�MX���0��B\�;k�A���_��!�B6�$��)T��s��`�<�S�	�V���<�Y�J�"e
�X�c@"|�Z+�H�Xrވ+�?}�fq��5⫝̸��i��V�t���K�rD�M���-g���l�9p=�J3����b ��6�p�Ct��L��#��O<9	k�.�"b�w�_�]c�2�m�U�-Άn��t�j ����D}l�������Q"����}�x�-�'L�H?`�`�Gr��rt��&Rlr�n���A�ۇ�����!p��s�+���}��4�B*��*���ם4�Gm��D�U*�������#�b���l��)��#_kyw!&�9�6���j�s�Ȩ]��[��I���p���S��;3b/�������5�Si7�wi�4��2h7�X�����	��@W��X/NW?� �̦�J�Q :Z�й��h.��5���C}k�(��2x��t����!�{۰I-�3��!�]Sm_�oz�؉��w��6$�������V�y�.Đ����5�wz�=��_,ܴ{�A�7�yK�S����o��0*�$�
+}k�O�"�6?��%�R=����T���yK�U���Q0e����k�/P�a���V�#���$�ܙZ��L3�.��~�6�l���32@ٮ��Cܒ�R�[�R��R,^w�f)�X��Ḱ�&�;�0n$&��,*{�|�Z�x]��"���Ѯ ����@;�Ln��	��mJ0B+��:�AQ��Q(�{WW�����ؿ�1d�c��9��t����x_͞��m3�Ì'G�Cs���e ��}Es{1�o��B����9T(�|;"�BO��n��B/!��az@��C�Fc&��2�H�}�D��w8B�?T�)��)�:��M �����!��
�mLK��7Vvc�N�>�(�M3����[U�H.wKeԝ�/RS+�=T������X��P��LҒ�/�,s	���Ih���R�`&�f)�˚Y�%5C�]P����X�}�rC�h�)Ȕ�ϓ�%?Z腣wpؒA壁����p��w�nЛ ��V���^<ׂ��+n�hd�6�\���C��_J�P��~�0��hU\�>��\P�MN��ܯV����u��kQ�3%g�����r~	Sj^���]�N,�h/�G���1�p�e�^cМ�n+�Rʌ�@kO�Bs1�a��~�g{�SF8IցX���.�r�\#)(!(&̵!�e��ŖU8�D�	�lRT� �:|��W���xr�O��]���?��!tE5ch�]�]~~�|�!���L?�E/0!(^�U�0��/�BKHǈ-L|�L�,�?M�Ӎ�`ͻ�K�<5��Y/2��lw�Q����1�WH�X[�����Fv[t�_f@�-p�$ޣ;�;�/_���U��$Լ�}(O+=�ti��!EږbcQ��Z��b �B��Y��&�i�O��gLa��vB�o<ԙ�d8�	��1�-*�#t�B�궴���5���ƥ�L�?�|�P>f���S��ڛ���B��	<���/��!�Rs5��.���	��&�h��!��ɡ?�w�s��e�E�6"O��C*�G����I'cs�;��x�扽2�a�	�!����#�%������݉E���a�
ʑ�Xo���qX�d\�8��հSckA�0bY��+؛��)j�L�f�f�(y���s��y)�F��b[z�ۡ��)��d+���r��6^�:TMm%��f=q�n˙��|�F �Rt/��i���2��a���t5��:� xO�I���i�
Y^H2�9�:|/�FV�9_���.<�lG��5|KO�n�Pb9~�X�}�ߜM����VO(������h��`]}���,�S�%^�zN�����N{E�����Sւ��̊N�:���hon!)�^eW6n9��f�2KPk/Od���?��a߈�|�P�~
�9z>���zYt+��G�O�;�@�����P�J��TVxH� �QF�=wt�85�=vʟ7�9l�OC�\�K^l�%M#���k
.!fr��51��6$y���p�[[(>���A>�3�~{�Gvm�*�r��2\I}�)Q�d�����N��c`b; �ެƲ������p�1�^�GD�r���p�^�\|H�[����[o�fH+���@vń5綠�7�x�|����Np��(�'n� ��I2�;��9�1�g}�י� ���~L�a �3[}�p��:}��4��ԫ�n�ν��o�F)�Mi�GA
��UI�E�^�|M��u�Y�xa٩&v��*`���D�<AU� �������D���X@@��C�"L�/���"�f�b�1����Ѹo�]�1.���)UQK��ty��QA�D=��]�g�4O��,s>�.��J,?�:�kG�4C�����T�b5�x�W�h���o����|����)�N�� �IDbXi�-ɟ�
�h��:|>����dhR��
�OW�lv/�X&�yOa��,�?��4�c� �U��Ӓ���'-D)0�\�H�D�u��a0�Ǹc&*�+���@�&bZ���C�����VBP,�Cf0��!���Y�x�_݁ˮ�!B����-'���qym��9�[g�%�%���a�fKL�y�si�{(��օ�e�G_e����5H-b���}�p�p�</��x���˄%V��%���C�<�/^����*�z�� �݀2}&8D%��	Ϛ#���!���[z��,'�t��5����~kzhR�{d�s�[.�R�&� ����B��I����g?<A�o.��Y\�tYҦX趛w�Q�r� %tN �	��m�k����"��<"��w��5�Q(\���MH{E1~hNC��4�!����1tڠ�����޻���������t�84��m�uN�A�f��h[��d����¼����u8@��/�)�_�Is��̱/�p�,x��[M�����������?5�^Q�sj����p��������k�E�ʉ������G2�=�e����/{ �v"\��*�Q��v�7\1h�/Ƽ�����:v��}�j),��vm�e�����4���?ȃ��X����֌J�vg�ͧ�:m��!Xꢣ��A����{���]�5�䌰b��~4�h������6��P*��Q\�L�}�͂�p��☙ȃ-�hѻ+��{�Bi�F��=5�0�n�F	��Z��j~�.����ۄo7���MA��W���p�2͋|�	!�z��0���UHw���Ǚ��QJf)�9ά�G���_"۷��hU�&?pL�\�������{��ghH��ۄlR!A[ FX�=���	�=�w�7��d�*M�{g�K�������?"�q
<j����I����*����{jUR�:�;t�*��:Gg3�C���'͠%�*S�8�*E>���W˗XJ�.(��P�����?9�����F�Jϙ�a��GFG�n��J�Wº�>ʉ���th�۾[l����@�NG0�Σ�����T�6�@B��ΎZ��e��a,>���ȹ��5
(�����	�� �3jI�%u�Yw�ε�ɷ���\_�,��l���0R��t:VQ7k��	���a��|�=��ˊ��go]7/�rV�q �����2m@���Bo�YU���Y�c3	����.��n�dp�����+p8�^��B\��=28�_N{`D�L�L����V�T?4���7J`R�j�j�K4E\Շ���>�Y[���`����:J�!�t4GR1]����P�h�lr-��\;�����(I�]�{zA*��s$B��{"�i}c�z��I�����U�P�Ů���bq8�q�1c�N _ȅ�tI�Ō�A�~��LdIa&�������W+L���Ir��� �P��ˑr��cd�Β�ti��\���W���=���Nw����@���e��B
����{M�����l5�X����dB��;&FW��O���{�3"ܣC�{����~�Zr�8d��qZf�jK��;&���Q�n5�s���,UW~�5G2�# ��x���kv�G�I�Ii|�a���q�8��E]ﳪ� ��g*0�t1#2�;M�5c��I���Oݚ�_Y�_��q�91޵�XO2y3l5A�.m�cն��N["�C��T���ga�]�1���hLI�:w=7�w�	������b��T)���>��m��ɭ����tK#ݺq����Ч��R'�حX����	\%�\|�>����2QT�M)�����������8!r�7͆ȕ��9��3N�J�ՔL�#3����s���ɭ��������I�raK�(5��6C��5ĸ��by��g��H����"��gPX���A��� ?�H<Z��'�)���L��VN�T���c1��!�P�]����_�R �]�i(wi�}0��a�/J%��`����ell����Y!?d.5L��ܟ'�a���<Vj<Y�JM�q@X`��:3���)��;�g)�f�����dq&:%q�TD:^���T�{V���I�=�t/��_[������Q�A�	�C$^Np]�Fd h�y���nh^���C�<B����I�S7��7Z)��21�\���*�l�ww"-��4֭m����;
�(� 35��Z��>��,�m�AcT7"�)0�����c�+�b�kXBQmY	�2�e�l�_(ި���J�k��ݝ��Z��Kv�&0�A� Rrя\K�f_	B�{��F�ȝs� �_A��8-+�:坳R<�R.~��f�3�5F#j���A+�] ���=� �wϳw�v�Z!�:�]�uz�����.*𴁾�#���>%����	������r��ז�����L?` ��<;�k%��C�_`�����8<h���w�0׽�|�<�����i$����27�Ss����װ��m�|	����!"��I	���#
/:[�z��P�:[���6K���"���`�y
R>��;.���isRl�6
k��AZ(�¦#�b�>g >x����2y��jZŲ��͈�����r�-u�W�T�9\b-�J�m�ׯ�p ���:������`������J�0 ��E����!�l��[؝WVo�|��^DX3���`�Z_�sHA�H�S@���)J���j#����M��42��3�Sگd���Af�x�Ed��*yN�>���1�}pk�̛��[}��7ߘ���_׉��/���H9�Y���i[U����,6]Z��G�5�on��q�0z��?sE�w�,e����+�`���*/R؏�%��B+�0FU�eiƝ'���T꧒0�T�8gp� ���0cNcT��LNԍ)�b5<��7�B������7�b	ʊ4���T
y���7�I���+�,bJ�{�¨���	�|f�Ov� �NsZ+H�K��MYL:��	_K�ÔKv��V��o N*�ы<�,��f
?r!An�5A-�K!PlU�
.0:1dsg�b�%!dK�=�*�!�<��Q�d��2)�i���H�dA�����t�/�\W�>م���˸ MhO&|�t��h��x�Ώ�q�u�j�Q���,���Q����iky�.�(��4�	��ߜ)��a^4�Wt���u���dL��f�)`��S�7��m�O����=��X��M�^�r[��o�q�NS�����A�aJt�/��g	5֤��M�2Uť�&�~a�s�������Z����L蟓|�P �~��]i6&��tNH˦�~Q~1�W�A�F��T�<��E�*x�G��PrW�F�V=�*�F٪�oe�Z��{<J����-QKs�n�T/j�-�mS7�kA�x��;~$"���5x]�8��@��@;LI�qll~]�D)XN`ʦ�ʭC�8����8<��+Ow���ȍm�&YT�������q���J�`��	�EQ�>����<8�I�?��#l�k���)Y95�I��%C� h�L�"!��8gӟ;�Tsn� .�"/`䚠Z���Jg�\�͚,�n�%�F"� P%�	�~�X��M�f<c�W��Mz7�D*��9�ȯLc���ⵌAWLzKR�uJb!v�-si����F��WswR&���%&���kJBq�M�~�@���6���椐L;k.���^Er��e�2&�\�
�U�y$l�0���� G<���[��Aa"�~OQx[)oP	aJ�ۺ�D��y�G�5�q4�%�
P��
�N�fi��qol�Gs�}�#�Jsr�6�Jj�4o���Ƅ�lq���x�W�ױ|e�&�T�N���1����P�7����Z��{_GV,Eo�s ��و�$��>��)2��<���Ѿ�|{�%�Θ�2��]Ƥ�R�7�T�40�(o�z�����1�ir����P����r��n�Y��0�本��T�Y�k�&/�� Ӿ.���}G�a?�{G�l��,X��(╫�R���N�NMI�<�?GLH��*d$6*�w�qT�4����d�x�"b����]�Z�������7i����Iuڶ����tq���ʹ�Q��[�������}�`�v��R�B��M���a�g;l�rs�����t3��K5��zM�ּ�c��z*�ȧ��s%2Bd��1@Qu~�P����؎5"��I�j�5��i��>�@��Sb���j+�؎5�j�L�>ćp�Y_��Ԥ��!eP�����:��A��LHW�.�0��7��Ȁ_mm�C��`C?�G����AC�}D��=�<��T��:r��.&z=/d7�����~��H&?�S�!���l��ծiJu�:f��	e�a��Zݘ�<;ï��]�R0�9Q�/_���i�p����X��8������C,�^h}��w��� `���W�w~#��"�3�v�r�p�^�������(`�e�W"��J?bA��^�Q���@��Qۼ����Oe~ۚ�(BöR���D�q-g��'�9,������&��N�m���aI��!��RW	F����Ȍ�����i�-D�|�$��4�+��f����-'��sdl �WS�ۅ0A�@�c�>�*`�.rJs)�\��V�q���Q&:u�����:�ꫴ	������ຼ�r_L��ŗ�%>k�6���UP�=���~kd�	�w^��\�c�g6���`s����,#\4<�1���f_�p�|�ō��5op*�t =|������"�h�e/�h��D(�����/on~7�6�H�Z��B"�t�����V.
���B> �77�r�߫���h���-&$�t���m�RBvf��{�T߻;���-]vV��?���0�y� �xl�M�]+�C��yL؁Bd��l���͵�lt�y�D�|�@;o7і7�� oܠ�t$F�������F�j�5:����$�:�ã�!q/�#5���׮�C�RπMč�
Ԯ	�@�Ƌ0I�X"��K�eF��� ~I:�K�20��a��N
F�8�\&�1�r�������H�b��|W�[�~c
j1-b��M�#l-�7!.JWŪ����쩻.�V�WS3��C��! zCs�@U�I����sPŘ烞�����e�W�P���x�,��Mz���R���e�S�Z�R�<M�t��,ᚻ����L겿qL��p�r��� lbNOP�[Vk�4p�W~Gv�@�C�>��p�@�W1mc�F�:���g`��/��vg��dp�l"�|=="��2D߂X��H��3j�T���=�U���x�#��h��𜋲��&ꆵ������X%͕�YUg`����g;�O3�wF�C�97P�H!i�w��wxʒk̶�U�7�����וea�bԚ-�j�-"2F>B�M�A�3��2���Y�п{<%Ki��n<�#6�\K��-��^+�@�0��4�.%t�xF�s��,��ǸzS���x �b�Fb~7�<��x!��f�D��ۤ}�`�ʾ^�f4�`]��/:��P��NUx�x���d�m�_�<��Z�&%�1�/Y������m�~xKM|N`���<��Vx��$�)����C�*��N����m� ~Q[�aZy��%Oݴ(��9�b�'�6��7��T��y���)��g.��s���W�٫~\%Q��[�A�<ag{���qj̉���0���&/IR�T?@���� �LU�g��[�搟?,��@��m�u��'E���?[��;)��:�������t��Q'W�O�ct���K�Ѣ�z �uS�Pњmӂ�ZAqq��>�i;@�hh��;�����F�m�K�"�d� ÿ�	{��P�~@J�<��p���׀J��mW+�nԈ��(�u��b05��9���v�2�D�[x��z��߭R/U4{�\9կ2Z*�9:���T����M�(H�MEL�R�ï�.����5xͲ�� ��ޗ��_%�b��-O�ޙ�uTRJ0u��v\�U���fS���iXR�$��l�5GyQ5J�u٪�;Z��ٖ�7���p�2߫��x��NP[T[��~{Ih֤oD��*�Y�o�&N�HՂ��� �,΀�p�܁�hy�����0C�ki�gl`�Jx]M8�VlŁ@yHq���z�7��<}��X�B�����}_���W��Y!_-���)j�i�����-BP�NEa���VP��a4��T��ί������8�]���O��a�ʑ����m1w�w3�o���s���������t5�r0��p����!DX��t�OC�B��O�]��^����!���,�i�һ����.�"_�*>�[vMzéK�/z�ȇ_Ya�RU$�D��'�e�fV�����HC�2΅��&:f���k�LժG5�=0RI�e�$K�a��߇�1.����A�;,��f�*��_�[1day�Ad�7�E��DʁXP �������p�ҷ��_��ǫ$r�	�ʣPrǽ��0.j�e7}��}�\E��~�>V���щdy�a�$ ۢ��F��%�Dc?��v8�/q��6l|��%-kBա%Z�_>��Y!��	n�=n��%FD��b�&x;�(x;������ļ�0���*T���gqb�	�xlB����z���?Ch�j+uR,V�L���)�2S�W�O����ѕ�ރ��b�%I�kɍT�M z�3<����ؔo}IZ"^<�l��I�/�W��-�i�M�]4���Bo�@�^�/�yVo�^e-$�]����������o�h�]�j������:Bu�J�����Sp��J���#"����04x�x�v%3�B����'���ݔr,�)�=��^u��T�L�5P_,�Yp=����#($��U5�R��1�+��y��	���.Y�49<�+��b�Lz!4��U��g�!'Lz�9�������t���w�;I>���6b��H���Q.ߵ�����HrPK�>E��������K<�j���лLNC��x_|6���WV�A�ftb������m�eA�yN%̨�4�>�&��;|˪%DQG}ݖ�z({o��ۼ���_M2cSO^P��@����P�r_��a
QD��R���#�����aAֆ{��P\E<u���8�8!jx���C�q�JŒ]j:hTeJ�����"6
n�h/m9]����ыxZ'|�7�K@�+��fTqY�iNZ�Ooε1�*ۣ%�c'��,c�ڬ���s�c��gme�6fvUL��Nl7���b�	@�Q�-�5�pИ>'V����rO�u��E�ڸq�4|g����JC}tB|�Tܢ���f���d���3�1�=�H5��@����C��@�)��&0�"=) ������}� fyv��b-II�������N�E����5���wT�'I<|�Y�p�:�~>���M��a�J��C?p�<��;�MŤ1�|R����ì��a8g�0�� '+.+��b 6c�6�����ao�$B�gM�w��/
x�&(��QG[*dN���U�
�͋���S�p޹�d���>[�,�[rr%j��g��!�8;������͗�Ƒ`����p}��.L�+[�PY(u���m��Jiw��`�B���Wo�)��V�z�nF������q�r���f�o0y��!����l��ټ 돚f�2�KQ��s������?��vГb$;JJE��N��� �J�Ѡ�~�.|IFS5�.���5Y	P�k;���?e�qlq(t(���u���nXcO�4ɒ��c���rE=��ƛ��%BD�D��,V��9���V%�Ѩ�CR:�P�ӎ��/J\.Ǻ�`�`W�]�>�����#�ͱMX�x
<SO��o�Z�kr�)fDD���
㸓��h��jVE�Pˆ�d*W�ю�aj����`��9�� 7�`"�JNv�]y���-,��䗰[9��{����h�$:B; 3!��$ݲ�v���[��s���� ��X �s��Q�՟����t�C}��ױI�2��'·����R�pW��P���[H�(���|��n$pu7�53(Z.9~�S"fz��sd�i�����W�7�:�,y�AjE:�6��w.^�+3�/&�c�j ��ޓD5��LN&�I�2IE,� ���s>z�4Gj�шe��D�:����N�h�;jh'�l�Ho/#k��D)�������o��>{I|�r}!W�{�U��� �g��΀�fzy��b��$BpL%+<"�=���W�7�㧬�V&��;b�����o7r5����d-���өɭ������tzA��7�����T�����4��]jCA9��.���=(u�4h�_w��.o���չ�x�4,�Sv=�)Aİ~�
�h'5c��N:9�2�Pw�, <ݡ�<ւ%�X&�;U�(���lw��o/�L�<^���4�k�5+�M��`��wC�T��;B��3 �Xw�D�d���53ª&�`��>�z����#]�=�l+�l�x+�FZ�EƗPo�?��
l�m����׉�cǬ�;]yc��O�K��p��p���5�P<��P38P_.�����B��n��aW�>rΪw�l�9D�{�ݠ�L�>a�X��ѸK`�PoD9�8����,�Xm�!���F#br�܆��b�@I�������J��`;T�zS�m�:S�1��kn�syϷ�ʽ��v�K(2�|rc�:۸���Lu;1��l~1R�_�Jl
s"4�?-@i�L<����(gƤa��bh�x9�
_� ֙»qȟ
%�??&���Q������X�o�����oK�=P�~b)GX�ߟB&�.����o/�$�K�r�,m@r��+���LJK��>�R�7ݒM͉�X�9��U�$>|�nne/q�^��{C@���
��'Ý�W��(���V+7�rQG�#QS>�%SM�'%�N{d׋U����9>�	���e3�:Ht!I̍���}���M��&%�&�4�MT�&ǳ�.�E;��='	�,J���K��>��Gx@wC�Q*^��k��0j�#$�to������ٕV�&M��%�}Etc�����W�&�w��M�Domޕ�BӵPT	FP����v�%�\�H�='\��vM�8��^$4��;���T�/SU:�o��\Mcbn�B����dP�d(�L��$��i���nx��,�h���o��:bϸx�-s��˚����f�#�{ԯ�Ϫ��b�]V;y��z�6뺖P��A��~���N<��[�[H:�[�HV�>`/q�1���\�>�V�sAad���_�Et�tE���x�Z,]�1Gp� ����8#kH�����L�K�����h�ՕI���D�S���hT�{�����NK�-�T�����nݵ;�,0�"�Nu����#P��;I��V�s^�zV����n���g�ĳ�hŨN1�|��e�=t���(����|!Y��O�S��v���ME)���H��ff����$��̰���}��-�H m�ؠ�O�v��[�AE������y��r/�K�L�B��t�B������Ҭ^�c�?��`
�t�KJ9h�gȰg[#���hs��b]� ��sveH�]����
�0�`2�Xtx�`5���jw�!ٕpu��UMl�ݫ�ϟ����ױ�<�Gh��\�O��w0H��u$t���w7K侃u+�$L�*�?SW�c�{�-SØ_�>�t�/G�5+�䱥�O@�ӝ������R|�/�f|Q� <�Sq�T'�H`-ƿV#�#�bz�Z���6�ڟ�$���e�j�o �z�Yjr�\8X"��t��A-��g���Z?},�df<��6
;�0�+�:��"z���Ş�Ħes�+�-�P弜8T��vG�ϕ�4�ۧ��Ss\@NUl�2�A!�z&�nLQ��Im��g���ă�� BR:�#Y�r�*|�}���
�/�`xt�"�
�g�3n��ة�+Y ���C=U�@Vc�6�\I��	���7��M*�2I	 ����_�6�aϡ���P�J_���ѻNǢ�q�I���%I���[t���$��=����i���ټQd� �Ϡt`�ee{�f����޽PpӞ�xā���'��VM�Wz9�Bju�/}��zFG���qU��FP��"m�W�����w�Ś������-�货�Oy�і�evV�孷��u�R|�������,�Nv�E]"�!�l����qD�&E0ߎ(Щ�>i�@ٲ�4�O[C���P��U���P�f�u�ß,�`%,��.b�9#�N%�p��v
�f_�w�y����1Ɨm�?,�˪��OH]��*�C��Q�P{�'=k���Uti�����y�g��L^ȳ�.X@� ���x�����Q/��V!{�y�l��8�vܝ���G�n%��\	�}����[ҧ���}߃�� �V#��<�+����r-Ӌ�Ƴ�N����J�.��*&R!�yA2�V0^�,�Y�]u'�����U`�����j����Xp�\H�[,�����>�ޜ����)b���K���)����̈1qa�U����u#P���2�� B�������H?�6�Q`��S#�;�-�~B�U�{��݃�b�I�t������Lż���O!���rV{���9��x.�����W���>i����C�Kd~�J��\��ۊ�Wjb�*��c�Q`�h_%EGq�Z�Sg���좴��k#���*3p�����*�)g��r<��H�`��jd��A������,��t?`S��2ߋyF�Wr�I�@��pq���2�ibx��Nk��-��D����!&|_�I"\������BP�iF�\�=U)Pˬ@�����"^�-X�ju{]zh��}=�X�'[�X�Bo���#qt��=�lG��]�W㓌����7��Z�4�ǰ��_�3�����'fZMń�g4m�ŭ.�U:�t)R�ӄb<��}wI�ԝ�!�CeI���e7�?Bz��:��h�� �eVdd{�*����
*�|���b���
2�`��s�c�x�u���<0d������6�_c�
Ų�����A:k�.0w�[�k}~$�7/+�=ځ�ǧwY�Y��V��.�6��Jc�����t2��ak��1��^�*�F·�t��em?Lh����䩪;(AU!h����J��:x��Œ#
f��'y5~�#�[�p՘��s�\3	r΢Dy����$����n�L`i���i0;�X�=\����ˊ�祻�M��3��
�fp�ˮ��Tra����J]���0�/n_n�h��cN����π�E�v���^��SX�a�}W+���o��Z6u���9�᥼�N���]~0�ΥU�
hDU*�� 7��^owbO(o�KU��UnUj8C�A܈gx� ���㝩��N�L��oB��W��3f��_Dk�ٱئ'�x}�p?LK�=�����ڐ^��T,� m�$O�=`�?͡� �_`(�6�*�m�D��j��Eʤ]c�S���)�O<o�l��4SUC�ϙ�9g��h����.�{T�٘��SLPw��Xb�va|�n�I\SGE:��!�W�j��)�3W\��Z�L��0'�K�k s�);ǛS; �`N5�e�6��q��IA�4���?`ڇZ%c|%�O]7
�!�Y ��ז����x4f�]-y������Nɂ�L�n���.~���@��ơ�����/ꯂ>TD�{�7#?ݬ���J��Kb��Y�Լ6�e�&�fxM��ǳ���#��xk���7F��a�||�嶧io�4BƆ}<1A�{r9 I3��������J� ���iS�g%�%C���� !*�}m�{XTc�0?��e�j�g�!f�u��OY�$�r%�wH7b\O��؜��%zC����WjC>n�(�>���C�r�;iX�j�`�bR��ZD��"yRZ"�SM.�)6�f����qiy��t3R���q_JFuY�	�y�� ����IO����@{:��jb)z�""�@��q��Y�8�<ܪVg$,���	�ȼ��=I��]4g���њYU�ye�p9�j�T�Xi��h����gNπI������|�%�{m�pCHaC�ͷ���Ĳ�]^��T2:!8�F��Dh�z]��!���0�r����^s���a����	 sAxu0��~}�Z���&ԇ���O�ǈP��@�<N)N��%9"�V��N�t>�Ȑ�v��s�h{�ʉAT��_k`�X���Y�o�w����ݣg�$ `6l�.��I:"8����E<����gv�nPcDʻ_8��`��m>ƾ�R�|�d�T�����X-È��҂��W �wİz�͸ܖ����wT2�[��;	��jcU����Z�@�wB���k!�YJ���Î˚��n�Q�RdX$�{M�Ȃ/]TF𢳠b��W��|�v	�s�	��MÇ���g�I���9�#��%�5��kN��}i�F�!���>+8���wF�w��ty&�'`#%XVU�A�� �ٙ>�Q�Xe��'d��3��%'"�^yoD:4�zg�gs��h_�k��_��Z��B����P����G~wes��:����3L{O*��." �����)s#o�_��
�$�P춴o�Zd�M�����S1��)~Fnx}c;�>�07�wt77� &�0�.����2�`���
)9�JϷ��E:�	z�D����	��f��
@��ߗe�2�q���7V�����Bt�?��PĚD=��I4Z�3DI������՜N.��L�O��ѧ���V�|cpz��f�jj�|"�7��bo|r �O�O��,9���p�Ũ��[s�Di��@z
m��k�m-����T�,3g�8������ v�H���4��E���d�\��R����$� �"��j�	Q*a9jrcc��"�s�������z�d-�7�P��,֍�'\�1:7��,8 �c�C ߨ��Ռ���.Gd,� +�yL��h�� 9��m�����=U�މ��o%��������i� 2;w��+�К�⇲��i�<B���4
o��h#v�3��Ҝ�F��Ml�K����瑲kaǷ*L^�[s��ԍ��� d��n	W��o���=:3l��1��O-6���e�}8`����T�[�2�/�Qc��%��C��kP�
tۺ��A�:~3�������?�;��f��C1`��jހ�խj�ޚ�kiz1��Ю�(�|<����s�����Y��'���E�Z��
`��ª%	~f�|������+O���a�&s�{�Z�GƘ\h8b$�k���!HJ����xWSqJ`Z5bs�)�4 g�.Q��tљ_+F��CZ:�7;�+�`K��4�=�*�'�UY��P˴l1�|�M���f�.�K;f5�ߞS��cOh]�j�3�vI�V���=��yn�oh�H��.�v{�1e�/[�l� 6��T����J���i����Բ��C�_n�#��+(���E��8(	_������?�b^�j��Pkn�E����/~�鿿�eoAC	����Z�t����~g�j/mG�c�2�D��)��myB9�S�J:K���MP������̫���mLHpF�N�5�q=��h{'��g �%l��%,�����]'��#O%z�f�0�s#�z���0eP0�T�@�52�L�N�b��,\.(�5�QB��6ca��������&ړ��	9��Ɍ����V�����lІ�����j�J	O��r��>]���zp��ncrx�F��W�����W�E�4�8Y=D����[�={P:��5��f�"�[̌??+�q�-�{ʨu.M4ha�O������6T	�r�";ڻfA�Ѳ� �B�g��8��L�j�ؕf�U�KD��;�dR1���� hw�'�,�B���\+7��G%;س+"ĉ7L~x����H�{{�o�����Zv���`�=s	yGǀ�j���:0���ԫ��;W·��F�tԆEb������@�� �F�}/��/_�j9l�q��@�5!������#{�k�	�υ~Ʌ�[BT������^e�?�L�����B���.��ŨI��Y�b��h��<?)��]׫�.z]I�3�"�L*�&ˢ�,�������e�K�)|fc����uwx[�R�ī+fw�e���)���ܘ=� �g�+�s>��=��1ƅoWL跻?wZ	)��MgyU]0��a��v�IPɧ�Ts/~��B0#
�^w61���żm�����_�32,��*G���(��'�I�ݮ�}~N�飍�$�ڶ*;B,������{�}����oyh�@ ɨ��a��c6�~7�r�4]�D��R���������/���e9ō7�(�_����^��3�|B�J[����^׎B�H�f�fJ9�?V�ec�hX�m�r��`�y�A!��	:�H�Id���:�`o�2���'2:�i���1�C��V��i��{I6�M�����g�]r"��[����~�J!oO���j��i=+��IDM�=�T�Ͷ4��ߡb��2��j�M�q5Jb��nB=���Z�g�	�
H�x_�t�e�3@��L|�_$3k+\H�i���Zh�qTd�^"¨-�Ɖ��H�@t������DM}?u=2���F��֕π{5��J���^�e0v��·�X�s.lHq�<%W��@j�0ц@r����L5�F*%F�:���d�~C1��;�P׎��"���T�%^�ry&��3�8DEP���	g��ꒅ���=H�ra�L�-����� �yX� \�@I���ls���h��{j	:s2&�I_�e����6s�� "����� �UX=�?�����冾�)$ci��tH�ފR���N�.�u���դpV+�ʵ�}�0�Nx���&-^���Ҽ�N�yX���c��;ܒ�EG�ۺ�ר,�;���xR�Kc�͓��|�;+2j��evsm�%�Y�v��Atp/����EE���-��"(����[��� \^	��C�!�0:�Xjn�i���g���MU�a����u!�y��G��N��� S�#�8$�(�ȥ��~�声��7=����[dOЖ���)�ea�+��Q��{bƉ�<�xL����3���v^� �Pţo�1���bUhL�Y�����<r��u�!x�#��� 9 �UM�ca�v�6�g�"-k�*�T�:��c�������e��Ù?����\��}��1��I���Xv�P�+7��lo���C)j��@ ���w#��W2�
�X��*-��v�7���]�+.�ތy���wT�
��(�`�XY>U��tl�����n��O܍�Dߖ���B�'��n�<_�/��S�W����@�g��])�}�
���5��N�^��� ��sⅵ�N�s1��n��x�U��.<��zD�W�Um}Ϯ��Ҁ��[X��4?g�R��"SF%U�_`e�C�9D�`c��e�`�^E��l����vaI�:�\7�0g�z��R=�'l��n�Nk�_c�+��k�uO)d��@���(���kc��Я}�aku�lq�w%s�"1��/,���?׊�3��~�ͳKƱZw�!gtꁮ���ع\�t$Zͬ}�"Es�y��s#p��~����ML�"�ŵ9��M �A)_�}܋䰡@ޛ�9vk
_;U4�@�ϟ��Tc۲�����Nm.W�������$Sk��Ų�F'8�d��@���Ε��*.6�۪��j|�
|1�ŭ��=�&^��d�B�I�g84�?;��S��٭���H��y*�Vy#o��c�dbD�)�.�5I_�U��Z��+�N��:�e�-~��˪X~�hY./$���Z,���1�z��\�ٖi���{$��wSU�q�n���I��_��s!�e��1V���؝��Ob��ӥw&�]o��3��5y�e��b��V��ޫIl3���S��g������\Oҁ��G$�? 
�1ޔb�fH��,�=�� H�8���0huJ��05XyUmS�^r۽�m�R�(��uk���xԶW�t�z؞�b��"�4n�Z�wC��[+����}n��� �slwӨ)(7^�92��	BKx��2�ڄB�O��T��N���_��d `���#�� [�[w��Q�](��S3�g���d:��2#����j�+�7�w�t�~"��k��ehw�U�vtB���Ne�hQ�F����A�hu7�������%5�[N�>{+$%�`hzb<L؛�����
����m�=�yz<AJ}Ng!� ����q�sn�^L|�s߁y��kZ477�u�&/Id��EN���f��C�3_�Kn��ޞc�x�o7���zF�Dc&d�F�?bS�&l��p9�ǚ�qPѨ.�G��(,Yְ[��a�x���"`���`�\�qC������(�!w�b4K��Eve u=y�3,��J���Y�1r���Ĺ�l_��o�j	�{(bZ���
]� �J;��a<��@.�q����[8k˘�Q6�p?ixd:�N�,"��1&\�?�������J��o����M	�!���S��s����ݜ�u���\N��܊��:T��e������`յ*��lw}_I)ATȯj�O+z�x^vQx��Z���
���~�z�%�e�B=b��"s��F��� ���Og e�K}Ń6p�����ƈ0�m�O��x[1�8�Zޒ�:�kTD��ׯ+�C������.sg�)�?��Z���_���,� s��� i>kNw!+�$�+C�Vp���H�[��^e2��h�4�n�T�ȏ��"Ѱl�7�;2���ў�J�ku#Q�μ�#�]o���20�����l}y� �Z�F�hg�M-6�s��M��D���\{�X O[�\�K�W�E��U�(��p!�?������3�Y�ِ �$n�J��u�$���#N�y���r��޾�	bt	�<�~����'ܜ)��@S�XHY4��v@,a���Z��M�~��_�RP��>$��(���$K��C��o�d'`
���ot�p��=�U�&���^��PZ�Bz���|>�3�q�e� 3�Դ�`�H��@�jЗ���Di� 8��q�V��_��ɚ��⺒�L����-��P�rn����	a�v�����o�j��v�s�iԆX}K��TDT��{˄V;��;�� f�C�T��GGLW�N��-�P�\��S>}}��!��W-+go65��:�.���k�*5"�!Mt��W�����cC�#�ڐ݄/��nK���p�m��x�s<��B�4t�tE��oC���Eֿ�%+94N�P��H?��y��6����I��(��[A���8�)�m��2���p���r�2�[�S^ؒ�t�jE�i���2�i�-��*Wi��zĞ�p������v�Y;\UP��R/Q)J]��8�o+˷�i%���9����g�����Nٴ�,n�p��p���z�*��Ȗ���_L���`��^�
=W�!���ھ*��GU9o�����n)���\6 %uH%Hg��5�u��=�3��7T4����$���[��#`~��*�4F%d�Zy��Ř@|oV4&ݥݜ��l��<��}����l����,3p9j���|���z�����g�*�*��� �1U}�DC�9������S�6Bpt��l�ڴ��������t��.��3F��Amn�n^������e`�=�N��������'���m�y��kl�pM$gt����!8��O�g��C�5�`��P�vj<�o�@��Qni��Wf+��zL9W���vZ<W��o�RWǠֳ|��wp��Υ��:�Ym]:��p�-�j
KW��Jp�#>a�|.��SCdŮ�z�c�=�2+1C�����N�m�d\>v�d���Z���ee�\!��2�T�o�BN�mZ��0����n�$���5|S����Bʑ�͏7���ٰsc�Y3�写�q���dpFN� "�,(�k�]����ש�C���`R�b�^�%O��
;YtjU$�9���c�:�7�y��D�{��C����/�Gy�d�0J~�HSO�B���ws���BG<���~2�^X�v�Rm�6�y���aex0%��E�`F�վ��ye����Џ�܋�b����'��xUy4bIZ�Z ���cS���h򶼗-���K�[HT8�ĂXw�8��+�8�D�{�	5��Ƭ&�@B1 �U��x���'D���T�x������b�L��>�hiP"t��(F�y�QǱtY��=J���f�p#��J�[\q�TI�w;$7MV�Kc�f0������w -]�(�ݲ�Z��q>{ؾ�����>���`��f�Փ�d]Z��	{(������^�*�-��G>�W|�����V'Q�K����;���}�G���+��Ζ�١{��sL��-~70iVt�ao������ɮ�C�t���.�-8߾h�|C'mêi������m����ׅ�"���z�{�N� Ol\�/�ử�,YRr�6�0^)��{p��X�Zl������I}O��ы�"����ݙ�璡*cJ��E��Lnד�˩�G�(�X�,C��7���ź��v�w(Ϧ�Q���)���J�M����|goXP���x+��������Z<�Sc��<����wM�3졞����%[膁�ZUޓ��ʦ�{�녅��N��g��oi�|?~�Z���C6�_)��E�o9+���އg,��Rב��Xve�"�>3�g�YI��I�Re�*��ȩ������y~P����:[V�pϙ�p���ܣJ[Р!�GB ��J��?UJ&.��6�&	tW)���i*Dk��a�]�H�Â��S�\0���4/��:���\G;48m)��Ih�O_^��|�;Un6�v�&12�/xPV,�H�^<X?򬚠�����L��]	�ի�@��Nx�fi@a]��E����� M<t�R͐�*�XrK�jq�X<�%]cp�+�
l2'�蒑s���R�jh�f�.�u;�6`=W���JY*�K���9�=�VH�]�$�����D��3[H�Y��;�B�����ظ�[�:Q�
sO��cy�M��Y�R����h���⠶���0����:�e�ճ�v��@�{���:���[�D�/	Q�1*f�k9��"�����R���y��#B�R��r줹'k7��W���>�������/5n�cS�2+J�3���yT>[��嵙�����^J�k|���eO۹4{4��EN �Gty�^�WеmC��&��c��Eh��ܚGV4�$�KM����wF�n�j��q#�p<>�{CJ
߳e�xL������U^�rZ�R9$y��~D9�
L��wN�*��p��S��e��q���%x���?�_V���0����im���rwoqB1G��H}����l�p5D��.���	���G+�	8�c��҅�u�Q9��'��"Ѣ<���
��T��pÃ?���x�4u^�cs�y�%qU����G�k�#��T�4��r�m�2��������m��f<�ﱾ�l��1M���λ��*Ys06K�O���q7�l^4��p�i1�N6M���Q��~v�Cȝ
<�3$D~ũ�E>ؿ&�bS���5C��T��u"11��'���ҋ���E� ����TJ����P�&�1�y�ln�;0f,:|�S���Ͳ�H#�:�
?`o濼öwW�p8�BM��je �_ω[IH��%T����drؽ�~��xC/ъ'M�*C���*�c�L�Վ�k���� ��@��ޣ�;;W��8�{M�ݮ$NI|�u*�_�s�d,Y�ɳ,>�!�	�r�un�O�ݰ�mW?�s2��.U��T���4�.��#�e^l)�E��D���?6s5��Ǎ���.P�͑n�Nj�%$H{��k�Ў:}9�"{22EyM�oA�]���ǰHK_;��Z;�Z�=6P�˺_�,t-'��[G��h�����|�3xZ?���O�~��F��i\����nrHX����ДX^�	�h�s��W���u4^��ef/m	���qm+�5G��4n*���`���3Ɏ�ј��ז����8���!ӵ|I�\��x2�:p����V�
n���(� �`�5�y�GbdB��ʶ���3�5�ZRT�W��`uM*����pX��Ѵ`ďg��)�c6��꽼o�����n�A��o�M�~P����C�~`}ENti��;x2�m���\1�I���܀s�z}My��ַ����]¿���%%�[r5��?��q2*sQҟ��6��2	L1=ꡅ�B�~��A�.�m9�`L&�v�MG1�TE����@:�Ġ��;�L�{Y�Z}����x<>�_82������:���;�w񳠲��Y��.�1���/�c���(���|'$�|�c�-������(Iq��ty�$��:}���6�x�"+[]�YW&]��+A�	�[�x|M�?F�
����MIKè�;��l����ǉ6,6�L<�}3�}Z�DCڕ��O�d�ݴ��o�� �[>b�(�F���u>��"I�P�A}��zj������G�� �*'�bL���V(~?�"Μ~.��&D������ ���u��j��!.�j��MhA���/����[����Y��V~Q`)�/�Be,6��r�uT<$܉�J � 7�n�V��rB(K؈�žf��x=������s��Ad�"��y���c(�n����h��K��c�����4�s7�R2�En���˴��U�FU��u#��z;q�X��bvXM������K�QU�F.0a_S��ؾt��/�|-��D�J�%.Q]s�4���x =�/<>�<�����,�ձ�y�=&��i�l�kx�� �s`��f�d��*AJ)k�5�=�f�_��%zw���C� 0��"��Be"��K��| C���Uc���,������5K��$h��M3
	{��F�p�]s��T�Pw�o;�_�1��S���k�=�97�c�f����vrW�m�#���!�(M�nϽ��i�VM����Dh@�3���ֱ���6�isj'�:�%�>��q#T� $�¹fU�w�8�n���>1�K �rQ�KJ���4��R�	$�]���w~y���c�k�
?#"�8f:�u��d�-*��{)($\��s�ͫ�qz\�����ZW��Zsէ��]p��e8�?�-�aS����i�S2�#�]q�4�}1�Tb��۫�K��=t��栆q��f��@�����UBE��z��a�Z�!��"tA��z�W�	څ8����%��p^���`�P�A��w�����Y:�/������l�5��њ�MڒB�|�!��5W���B2\��L�[T�d�d�g���'���%�{J����Dj����:��>`��Ʈ7q�K
J�a�pQ�ȓ�����(�(��{�v Vo[q-�5٨�21������=� �����)�P�`�wq�>&H��u ��\�^|�9�$W����>|Ǯl��l�j�?�'�P�2���P�L���eL\li��5&�$����k��O-��&݂��y��&
��M�Ȏ]�GP�Ѯ�������σQ�{d�ӑU��a�?,�Y�h!��Z�z��ٴ�f��b,�u�R������XD:��E!t�+	��.�M��PĸN�X�\3�+ME��6\X�L&p�"!��}���\'ee�8�oc+L�v^�P��o��� �{�1�b �o�#��u��7<	fu�Y��2k�y����r�K����:��{.�^E�����T��iz�痫P�����0j�%5[|�V�;�"z����j2v���Yh�Hշ����!�k����-�����Ĕ���ift��m�����{�݁bm{�<���yI��#I�o�ؙ����|�,Nhːb�aR�"�0ߩ�I�R����
��/�LY�	��7�'��p{fc�� Xi�QF���A:w�(�#|�fw>��I�;��qd�9c~%�K�V���ۏLe~
5�� ��I��:��v�/i�E��|����g�&&YE�0��]�;�e���[�o����|Ԋ1�����`��ܖ8�V���2�o7#$��'������������p���A'�/�
nM��-�ᕬ�N������12��uy�jvҟ�l�]w���nrsjN`���A㆗/&V;c�K:ό΁���oJ���0P�w`;ix9�4��2�����
j�f���
�$"���v�$���$�w6�ɖ�,��h��1�A�g�0g"B:ÒVdA|��@Ykػ}Q�!�I]�?���s)��NU�/�4B��S����ů�,���(zJ2ݒZ���6�A˅�ރ<Z��L��٩��?o�U����%_Z��{��p}�*�v�i��ȧ��Vw�d����64y�@y��e�b�ϼ���&p[C#���x����٘���,m�Q:�'O�w��wE�<zX�ť|f��c��'	v/�*#]y�'H� }G�]�V�����%%ag3$s�{�[q��x�4�t���1�?"Q��g��(a
1V�W�-�� dٸK_Ѥ�"$��0Z�S}�'*@��ڪ�r�?�=c_X޳lg�������F�=�dJ�ՙTc�GMD� IF��u^Ϲ)#���CW��n@�H���Ӗ�XᄨS�q��A-�}���x��n��@.���i�w�wI+b/�����oP_�R^��M�����å�r�bY��c.#��!���0P��:��x���k�W�K�Z<�V`X�(ʉ+ ��� $��хH�q�*����T�$V�ʁ0�:i�xt?s�8q�_�o�>�GR�i�W/W�����#ƑQ+��4Kn����x�ћ�r��0�p�ͺ�U{f�8PO;)�Ւ3e6�?�����>
����U�}�
�C�5����0p�9Lz����S�g}�Ǯ,
��A��Dd�55�!���>5=����w;/�*��A�/��>��pU�_�=��
��V�8O�s��T���>�'�A<d;�B���SC��E�زW�Z�e3@j��nY�DP��蹪���� F��<X_d����6F� �����ίD8�9�wmt��@.JݛR8�6ޙG �l?g�Uj59�q�Ѿ�@J٬KDP�ߨ�y��5a� 	F�O�p����^��Tn(�q�A�k�a�������%�e�z?/��G8z������o�\���cN�0H8N��H��;�	��qYW!����rm��_Ֆ\ĉ�|��B;[B�K��6	񬆼� S^��[V������x ��QohC6�[Eh�C�tG���]K�\�����|VUXt�ݑ���>��@
P�|�_��
J*vɖ!�l2���jw���c=?�Th�Ϣ>s�v'�rF�8�}Y؃h�;}�(L�q)�
� ڬ	a��ݬL<Y������^DC&��T��!ξG���y�����������Z��	���Rڤ�zߴB��*6�'�Ƈ�D- n��Ν�⏗�`;��A�g�c��n�C��{6k��ׇ!o�"��ʤ��dg-�2��I޸w�����W�n���&4u?JeD�
 ��'@�#k}k����C �j
nƜ�#�B�g�Ğ���C<[�������{BC�L��}�Q�����
ҫ���5%��	�QK_x6 �*{����%��{�Zp-��Q�l? 0�e���l�9.��#�>ہx��I�l���8���4��� /@"7{yQ<�m���ѴB�!D��� ���kU���e�c�~��iL��D�/D1�e�V��w�O� ���/���y���2�5�����r�/x�SHE�b��!��0�07���xB"=:�ʯQ�w�)��';�BW5.���ˌ��clh�G(5�����MCY1{i��ڎ�f��S%Z�pϺ������Bg��A]?���j�I��0�սM�7b����==�����<k�����ڐ]����������b�Ӊ:o�6��i>{=�4�)��N��W�D��=õ�!ZO,�ź��7����qEj�/~���o�+�x98fN�B��]��~K%�1� ���j��YS��K��������"x���D�?L��_>֣�Y�.��<>�=�3����a�.�	����3�k���[z�;���b��j�h�;�5�"�!�1��x����b���'�0��L��e ]p���5�&�z�N'��+N��Ic��6e��S�F3��P_!��1��>Ń�u��l�lS�:@��,R�id��8���xuR�u2Z�o��О_ƂV��ݜ���j�1��ss�sy��aT��0e��q�}��}�uF�e�4,I 0}U
�m3���%q	�� 0ƛ�E��V&@����R�a��Ye�X��>C'
(�21�驋ͣ;;���g�t�-!G���qwa��T���wO�V�La��RF�Y�Z�����')��N�+���kcIؒ��C@���X���E,��,�1m
�S��>�O| ��WIZh
q� Kg���i��[\�S�j�W��0�V�i�}2������ěb{tn�!���ɧKl��,�uƳ���T�E#���K(���R�N��~tr�Bz�B���!����`�#[Jz���U 
��O�L���eBQ�?��,�9�8���:�N\��j���g�;�TsC+�4vK��U(�Q�IӫU��3��I}�j�UL��zfi���NO	�%$���� ��{���F<��Vw�d��f94Oչ2�|)�YYH���ҽ�N2�q'52���,���&�S�̨�f�y��v'�o�n����Q0\�,��"0�'��Wp�=ۇ�t�X͑ _�G�g�|n��]�xV-��`{MK~ζ�p��%���r�·�T?q�1���M�Cɗ2�@/�t��ȝ�����R�W���P��hu�Z�ˤ Ïn� |K2[?2"�!N�p��R���(����s�ghټ�*��ٽ��u���o�[�b����}��)x5}�)E����^|w#��GRg��~�~��X}+�1W��v����.Bƍ��J��A �T���U�f���Ԣs���p�i�<ES*�u*W�U �`@�H�%^������&�2�JBl�n������ร�[����e��)+�%l�J����Ɇ<��(,��F��'��Hw\��rm,���ql[r��g�n`)��4N�*�bY�a�����<v�B��K�ʽ��TbV)�Hla��؀a@�� v�2�4G�T�I�`��n1t��}S�_�����f��<����s5�j�8�Y��u}��xD��]��

�k��l�xq��V̀o��8��;I�k����iX_ذ��}/K+��=����-��[�.y���Y�A�_"I�U<���R�h�iF�|��gP����Fչ4���{���&T�H�;CM�68�c�t���3��N��^�;�0L[$���KԪR��|��ה���!g7����&�-!o#1{�;
�=H��$FB���#l��o�m��F�czTT�n{ 	j�+u%_#�����<����:�P�͟��' ?N6s��	m�<�	q�+'���s.]޿�8��?Z�ݝ�+D?��y; �y�O��+'(��T����V5P��F�t"����Z-_k����T������x '!���'9Z��])�?�wz_�_�NCw/�O�PMeH�H��+�J��g�<Ԓ9�ZO?ln��0a�mZ#��AˇF��ms���Gx��p萹��x�5l4��2v|�nE����:M���/� X6��2�n,$.ć���8>��d�كJgE��`�\�?�$���d�~Ul��j���J���+Y�c�ڊ��1I��1}[���@'��]·\B�\U+n!yL����-,<�WQ�;K��#%۟�rT��f����/���8F�7��=��Y��~b��m�l�\E��W!E�ߞ���n���Tz�i�I�s�u\�[������fQ�pBZ�B\�uJ;��f0�����Ķ�>6Na�FB�m�N��xѪ�8�=
����-z���-A)AZ\Z�"��N�� ~���fYj�"'6�)���@K�^�k���.�>�wp��#���{슔^�i��K���H�i��?0�s!n܀�l* аP/�*�MX��3EU�5cq�#n�,��ћ��:4����g_���4����4r��а(��$l5���!��,�A�b�{˅|�3�ҷ�ڶ7�p�CR�H��Ө"��X�Ks.I�	I�.�I�8�DZ���2Ѥ�l
��D�P8J��J�95���^�b���5�e,`cu��$���	+g¨(K�|�Ď�9 FAT�mW)���)|W�@���G��O��W�������"	.U��P܇a��q��o�b{A�yu���"��ͭ(����':��7��A�<�i�^d�Z�5�͖�;�W�e��Mcٚ]�8״��t�#�l��v�8JH���"jt~� C��V�ϔ� N�uZh*H�y6l6���h�N�Q4/�{�/�7R�k0��Zۑ���z�����~,Weρ$�l���|�0���أE|�^o�u�SԌĎJb�}*���P��ϐX�`���#dڼ\p�S��:�4
�2цtU��怫���6F\ }[{��WG�����[��=�l�aן�ìq�����sZ���;&�&~j��jL/pf�vf�A�ډyxll�v���� B�wʠ�'o����n �t �'�C
�;l%$����/��1A'�$��ymA��2�a�W���QD*�_TEF��ۇ�5S���;��_q{Xs���� i��xH�{�ӥ�����.�ے��x��g��$�HrQ����p�<��*gd�E�{����X�"x5@�1V�]g�n{Q��\�0�����ܺ>�c�|+�5~���Q�ؗ���Y�����<��j��]�8	ږ��l��mw�N����]����OX�,=P����X�"b��,��@ځ�S�6��
k�G��S�=�̜�PG����?j����bz�;.)t59EB>����������L�Jˏ�G��3~��ͽ����0��Dh�^Y<@s�[�UKJ�H	�zu2g6�82��:|�	�b��z�o�nϼ/�.ʭ�Np;�Rq"�s�Ȼ7����T�QO�}vfP�~�L���s`��ƶ�L!8M)��vT� 8Noc0�)��E�>�9�C��e>	&+{��3��!G�~;�OF��4}ݭ5�D�xuk�}*)c�H��<~���;T�fAnJ�_ ��-O��H����'aI6�y��B�7!nXKX���"2<s��4NG%�v�=�����p���S�g{'W鰄^
[����3}=���ۏ��_E֊�r6I�H|�w
��!��ɿ3��3�s�,X��s��BZ�A���P��_���Nz��?�g���_��1����ۃ�wխ�M�&r�),[�`%�X���ۆ���\2�H���
�Q
�W.D|���bX���v��٩����z��Y)�)�>�s���fs���c��B�I��:>E��9zi���!�.�v"A��i�Ň�J�c����ZqU&����yx��VY\�\��0�����9�h]��54�n�l5:�8� Jd<�*1�g^�	��^���Z��\e�i�-���Y"]Y�;}ݽD��\����R��8(.��L���	��x�)Cd:��%�Ƅ����2���&X����UE	��`�NS/�����K��U &��וƈ�[�b�XHUl;'�'s������L$,Ǩ�~xǌ����O��-[�3��r@����E����zI�-�S��I���(������R:�{(��?�]Vi����3��6���uדsSn��=��\��'Ko��a�6�|l��;a���趵CR���>NO��z_U��U|L��Y��ŔJOz��~Lk<9(l��@�T��#XT5îf�mt���Ee�"������rw�}E\���h��vÖ��b���9�+���xܫ����eQ��Bn-���3�1Z=�V��ȸ<������q�Y�5��@�3u��ǜ3
@[ȌIf������R�#�M{O
�Yc�ȆUo���s���E�x��In4'���n�7�ż�ڰ�2�k��B8��Qum���.�1���;:j�(N�����|�I��j�ݒD�<OfV���#��,�����>&�{(��8�m��_8��N9��A�o��%/b���߾�f�u��1�>�q$5!������"��mz1E�H,����1יj�n,>Q ��3j~%l���_������n;��.�1'�5������cn��GK[��V{ ���WU�)��*V՘̦a��)9@�g�<A�85�p�O�7IFF�6�@�H��L��:����B�8lO՜&�v<���O�4��q� �˚#�ʠ��)�C��h�#�p� x����)pR�:'n�3��y�d������+ ;:�7� �3���T��瞡�]�ʍ10!gI���@�l�VPn�3[IX����1w����Z9-����9��)
_ڞ�����vaڂ������D����3CJ~FM{]�eݺ��"ʸ,� �Z�^op��K�sF:�o5ՠW㖒���=��ou�U!��.6߇~�)��;��1��I�[C��[�I��5��q����g��0� ����{N���']��{�툷D�e��c�%mq���J5sx6�h=��%��À ��z����6x1��Bx�*"a��#H�� ��(χ�#ru��1(%8%�qF"���f�~W��'��~�?���X���<5U����&�+��8���y��Dtv�n��:!���姺�H���H���� +ԙ�������oف^��"'i��6��#�R8�?�n��?
�(7p����<h�l��1a��%���{��/9u��:m�Ȇ�4���#{�Fz�~�Դ�B{���e:ch
S�2zy�����מhvWD\���BS��(8����]ƾI�R��԰��D�K�Njq#ǶgKlz)�	W�m7q����R"��3� �W
'�x�������C��f�~��ejeTk�w�FE�y�1�yy���֕Z����U@�����Ɨ%ս�8%E�!��E�{B�R��N��8�
9�f0�v ��t d�y���."F���h!V����!k$_��$����'�Ԓ��!�mp��_�=�bF�?6;ک�n ��# 7"�3�=���+�?���:�|^m) �ӍE��xi4R����]�*haZ�6-�^�a�!��y�p��M(�~���Ơ&�z��۪���7o8&wl�6�-Q�궩b�������Y�ӵ?y]�7B�h�I�vQ:-�V�|���%��)bUٱ�Bf̋�4L]|J2z8�a��eB���_��z���<��8������y��D�ml���� � fG�y��:��W� ft<%-�[���T�ϰ³���(c��lxx��B8�b�ȉ�<F�m��3}I!�"�~eB_��6Dt ��z���{�_:���OtZ�4o�݊Q��t9�7���z�t,l��7��S��M���Rf��q��qn+;�H�r�ˑ���[�DGT2.��p�-�E�0��g�>^���A^�R����™/��(���i-B��ֹ*�.o�q!ۨ��׭�I������c�(ƿ��v_�#�ͬ�AA��(�
�j�c��=��T�{Ūo��]ϔA_C�#��#p0��+F�[,~��!�bVۖ��DM	���S��^�Ub�v��ڈwd"+n�����ݧķ��G���7EEG������s�.�_�C9���rwC�ȩЃ6�3ڌ����K�o�⣤J	?�<ן��הy{�oթ�R��!�Փ�A��&�����3	���~%�m�;�g�����H����X\�����x�٤�@��P	b}�R�Ji��l�g�7B�m���n)�p���ZBWA�,d$WN$�S{���ihT�ށQ5^]�;�LK~*�c'$�*ݏ�x̩�^#=��b�JI���&�]��f&M�ٛn5zQĔ��U�|�i��j�Qc/�s�, MP�9 �k;m���_&]�s��8'�w���Ы@r5D.`�5�f�K?��f��0�L���i�ؓH�T�W���_���b^��d�,�#�(̼�QaZ���צi���y�0��R_�uriu�ΣA���� �R�,3�5���v��Sa��tE��j-��XB�11ۮ枘��5%E�]��Y������7h[�Z�=>�L_ù�gv�Cx)�r�<��=�U�/������?RaJ�l!){!�r�@oO�4b�)��q/����Zt�?^���G�F�n�,*�3����3�
�ǂà�6e�RMe�az��ה~1�̩Pn���<�nlO�gC�csa#�o���e�8�(q$H$�uy���(���I�c(��	Q��R���Z	��y|]��J������ ����<L���S��YdѭXoDN�w��r�Ddp%�K��Ts�X�T�Z���\�;�&�K1�(YQ�vЎV��G;�3��¡��Ի�~�X(0��0 E����'��}M�˘�!!B�3V�4���.)�.]ؚiG/����?v �>����Q�����ț̸�Y��1 ��j�p�H������K�K�K��Gx��\6�B+=��^K-#~3�u+Y���Nq=0Q�p�Xږ��\v�`q��a3
�
>�-3�	9�Xܖ�]�b�K�/%ש���f�)��~DVtvŏj\����Ҥ2�IP�t�����y�:�|鋖�=��6y������iV��zVtA�͸|n�J���p�u�a�Q�s6p1��r��k��!�K�5�F��!�5��ѯX�a�#��Z�9�8�(�G4��vl��E{�1&]�E��>��yx���ºj�aHRr������\Z*�/R��� ��##"�5g���(��	�D���r��4��(��띾&�20˪M�M��D�w����`���Q^լ`�L���Ւ2iFSۏ��n��u�]�lO*RBT�֣T���7��������?�S��j�7Iۑ�u����W�*��J�?��E�uY`����c���F!�P�tu��dr��/V�Qӝ��Cu�㘍w;ia�O���|p���R!��kq�ξN�Gx�O�S��P_��X%�<�C���Ͻss��)�͓�mn؎���K�#����	�~��)��k���i�V�5'{F8Ӌ�\�Ì�Y�P�U'���-�-M�|��VO�A�Q���I"��Eo`Zh��d��G+�T�������&�"#f���5�ď:�o�E4h��Z����?q,u{�c�X��0o�tb$���`g ��Ѩ}����D��O��(v�;�m�D8�&�1)�n6�F�ϗ�\:�B�Ra�ק�,���~������|~��C�~�{"��a.���6;�_�?D��AZ����F`�O_��G��__Y�r��������Q^�Znrq�����n�Z�)��_zg*����>�I����f ��e���8�C<)	5~��,-���t�=#����Ht�%T����w��X~��QW�J��Ud����;��U ���r����+��r�:\-֤K��;��z&�v���H;������`���s\ٚ��C*W%<c�T��=Ll?r$�;�מ��3ɬ��£t^-L�g��'r{����m:$]\��U�`;.]��>]ǧ�/�v��yv����~�7������9��4n��?�Y	/��{�0���eO9���EK�������{�G��@�)��Ί$p�ׯƁ�[�Y�!{��#�]N&`��D�-nMv��j�y0���q慼6d�N��F:��[��~"���2��ĺC�JO q%e�>Ȟ1����R�9#~S?I�	�����l�d�*_\�A���a\�-���G�Dw�V���Ö�Ya��*�\1�S��{��wn�-O�(�D�a?��@$4�>��y�h�܎<?��.����n0ȷ���Y��in�\����*OM�L��뒔L����)p�Q�e�fҵ�y��#���N[��J��e4�W��e�?/&���1�f�\����kAmUL�Y��Hm�I%I��1�2h|Xq�vo����6�8�/�*W�2lG����[ĩ���8����1ߜ�M���^"����ur-y|�v���}0H�u%�`�P�X#:W�-0�<�(�N�拪��-A?��'YEaJhLϯ�����rM/%����,�E�����\�S�#ܶ𬮱7�G]�_��{61v��:n�R7 ��r�(
�uQ�� W�&ض\CDȧ�%�3ƚ<Q�r��Ȗ��?���F�v��(4���AN'S�����%���X'��;��'+�m4�X�T���_,�������%[���pRD�}kԗ�����T���Z� �#���qV���n�t��d��7�g"zÊ�P	��������;��\�2�Z�@��bˊqY�˪>"�0��z�l��GL�0M�����NiC}pw�I��L��-&�	Gh�3#,E½̼���Ud���r�����w�S#��L�%�ʵ�����>�����-6镅 A�i�
�zz��(sڞ������}i�D T��˨���=�:I�~�4���.4�"2��=ӹ?~�
�k�P5'�Xl_(��Ż�	>!*Iqi�N�*�:�9XOʪ�`���c�"�9Kݸ�d_~�#o���ѿ�J�`���hf5�����v�³?�������P�IxsF���k�%5�E h�E_�bt� ��.MSY<���[���~�lpv���0��N�V�>�~���ٲ�C��[�r2e���W����B�Rl��'��\#\w,#�k8�3D��;N��.@t	9�!`'����=��߄��S2�3�u�g|H��2 \�6GF�/`6��y,10BI�)��%r���0�&�����`��!|`��]E��1��<�=Z��&[#ͫ�-!=;W;(����΋��?W�S�F�<9��2d�}��t!q�H��ƵX���W�,����S��o
w_3�d� L����(O��fN�.�}���y{�i���f�>Ҧ*���y���Py���L);�JS��"�R�:�/ۀ�NՃ3���(8X'$�I(��t�1/<��!��z�P���g{��ɕUu�������#$j���E�`ʮ(~��'C	���c�y'x��cx��#�R��L-�\�6h�2�Hz8xM1�D[b��uxChc��(��8*5@�		���,>{�f�y�{8کY�T/��gɕ�:*,$���`a3��9Л�3���k��������Z�c�~xh>ق������y�(��$�o��S�
������EH����'��.O{(}`��ي�4���;W{�wf:i����cO"	�G��Q�@[���MR���J�c��^�a�V�����}}����R��;�
����uR˳���q�Vd�����WQ�|�[8hi?��>p%��0,�vo-�b(�*���5�	d0��n�*a���%b?N��W�ot%���0~O��ia�+���nsh�Q*�Y��-�8s9�w�#�J�6}Uqͺ���3�G/��y��gŘI�E%a�3�K��m�8�7/]���&Ng��h��	�XNձ��=,<��U���-��uk�C�%Қ���Xj��fs�Dk��6]�� ���]��] �)Z�\7��c���7Q�ҟ�M���Z
�eE���(Z�᠆�%�7.b����ԃ�3öil����O�����D.�<ܡ��Ƙ2+fmL��1uT���'�Iև�����b�36֫��Z MK�ƍh(K�'�%�N���3m'��-l�*�nrU�Lo���ۭ�}>��]nd�솗gK��=�$���]F�z��٣���xI;� ��h��&X��/��#]ê����?K�c���=Ʌ���U�����V����j@ �ǘ'�_Y�y�ԯ��џx�M��C��}�����Bf2d�Xh�����k��9z����X�8� �Q����ayV]���JL˚��vp�;�׬�������B9?Uފ�]�JR&]?	�i��
ws����K�jC��Ss%wn�ҿMF�yz|��]�՜�"r�@Ж՚�:*@�3)�)�|~@���9�V�T�b�l~�|�S�Y&L�5���0�v��X��՟ �h'�p�����>�Mlj�3�\��;�`#7��Ѝ"�,�����S	{��}v��֋��|3ɻDl�*v���-�n-=jrS���)��Ay�A�Q"�?��X7�w��q���L);������T�����$v���+N��`��e���X��J�GMz�M�$������{���qo���܄�.q�����ޥ]#�U����\�N�7�D���/��+�:��h\��{I�5�&�}T.���2⁃��a��<�(�nt.�)�i����D��=k��;A.�$p��P+�s�jϗ�����5)8鏃�B'��$�O�f��A�Ѵ��~��� ᘹ%�{�hQm:1_�*�	��%�7��I�I����/��<\����ϡ�ǋS��i�d�y�Aa7�P+Y�%�7��s��D���}��ƶ���5Y$�N<e�C-�)��t,ڷ�d��D�Y[�-�|x��i<�~ꍺ�闭�B�²���:c��N��K�h��F;?Fn}Yu�0����S�'��Q�^�����w�a\����f���\l���]qdB�� �������OO�����Tg{*���� y�E���Q�A�\|���P�l2�U�.��j�@:�)R�Uxj�j,�<Ɣl�9�0B�T���Q'U��8
��k�6�J6�U(��m�����]*}#���ݒ&s<K��o�{9���W������ݬ�G%S�9����W_�鳚��b�_eO�����HE���I�"��nC�o�o���P���Ժ#پY��D��5OMN�~��o�n?rV��,����n��%�m�G���R�&^����FH�3�	��0�lk�fM�kn|���h}s�7�3�z��!k�y���5�\��`�5�S�[$�$��I�j���c�:K1�?F�+��b>�?��5Őt}7�9�s���ȝ�aɛ�E�;3C���G���J�02V�g�ϪR�7ɔ⹽ @����A���ρ�6y 57ּF����	�pp{�)�+ݺ������UE=��죆k�I����*����d�zl���UѠaT<6�?A� �Ph	U�2A�԰�VJPׇ�y�}�
�~��~�ff��;r�7���"��{�;#G�zǒ�n��9>z[��M�U�7%!��1�U?�U���C�xc��ե3��K,Y��P�7h<�Oj���5I�j��ɿ��
���]�11�!Nv}������d|ǒ4���OmE9D���]q�$���)�s�3��ɡG�{�_3�¿�X{ɟ�������DĆ��e(n��97�Y������_xhZ-j������J'#m����@V��a����K�.E�+���m�z.~�>(�3~)׊Rxt���Y�0�9�3�;�ή�=����:a=�� ΐ�����%����#�2!�γ�~z{f.�6�����u���
�K��]��4���|�RL�C�R���S8<���[�F�W_HK�ؽ�.E5up�x$�<l�=�E7��9+R��T�x�$�WS��j�5�����!����ͳu���X�e����4��)����8R�`jU���G웑f2�Ku� T�x0��vZUh��flwhű�W�J:?���s���3搭k���8N��h�K� 2��Hų�}��Ô� ��xC@d�_�� �1lY�*�G�Ncc��S�s�>���ĚL��_ac?��}�N���Cަ�g죏ON��/��B�XQh�6���"e�,���z�=�f'����]�<#e�aBR�K/Lă���Ϩ_vҕ;��JWA�Z�TPY�@��NUw��hnZ������6A\>��V�ՆNV ����w}eW*����ª�i=��j�%>����FI��/is/9�ەKu2���_-�f�%_�4Ӈ�h��y'��XYϾs&��<���'ѕ���XY�� %-῅Z��!ew"�⳥�v���@x0&����홗Z�)�W��r���2�z�����^�%i�@e3J젰�������ū.�=�n���??�u1V�>�w�S��%J�7�@Rҝ�1����[[ܩ	;�^��:n�u�V�p���pN�5�b���k�3�j� ���e ;D���<���J��c@&W��|~MR��/��f��,,��DDC�MO3�kO�ؿ"�IXZˢ�u+d�W�F�p� ����H\�Az&������e�M�uM�B����\s���uJ
��`b�G('W�I5�&�r�b��fi�ؚ�,�qlusI�X�f�[���2���0tS09�7&���^���gq���>�C�w
*Z�����G���M2���i'�9��H�n����.+���'���N�zr�~ö
(E$ً�'L$SW�'��ׇu��~ƫ���W9Z��D��	�~��:}"@�x㺰:���n�&PzB��Pb��t��9�@ \�$2\e�7�}��=j�S61�!^wEv�q0��wE��<�T��=�c3�<BI�r���	�7u�u��K�J9ӿ^�W[��n^�!��q�T������O�嬎���j���I����jj��Q�E�i�������Y��	 �\#(�z^����O���;���8T8+�EYW��T�AR��������D:�A��ʣ�ЯV�ir�&QEG�Ё���pբ��0e�O�������� ��7Ҕ����?J}���Q��=�7KF�h���K)���p�mY���A�����4���|G
F��G1� q5G:ٯ�䫮�����(%��1Ъ��;��*ĒAt��!D^cxؠ4�8_[����?�%��S�F*�R�{��],+�XC�&�oq�gU�I�@G������2�A��O}j���2fk	=!�iIW}^I_+�l�@Ru���b^�����_J��a�5��r�-�ȸ),Eh������� ��L5��J,�A����N��8���ZR�E�9�y+2�x�Ya�|Edd[���2�}��FĎ��w5'=���x���D�쮅/��
5PHYk��)�~�$�hG�8-���P$�֥�t ���1 }c���)�r�m�1WWǡy������}�m2A�XW���Y>���A������:�i��B�B�:�˶��/��Qc��d4d��J=G��"9i��k�H����d�,���T�bIȢ�DX������-J�t��� 1��s��9��{����e�ml�?r`{\>	�|���V�ޫ-W|�:��,����T�z� y��H�k4/j���D����ib��uy��ţ�a�v^]�Iq�.I��*�P6��M���nzؿ> �BJc�;�(�2~��5���q��S�ºD��!� �����~w���]o�-��4^#A��o�+��T�2����#I��d�ʦ"xg�@^�s��`'=)���\�1���B���|��G�su�]���w�e�n�u�n�ү�zEP5\.�5=kW}KA�%5��@�?�C�~=^O9@	�+q;�y�5w�9?��e��@O����dp7%\�VL�f�mo�*���Ȋ6�J�V�&�D��>���$dBN�^g�)h �v��+Qp G?g���Kp����lF�p;u�o��\^��h~`��[OBAя}T�چ)��F�[��'M~HWg�W�l��P�_\_Y��^�M	d�[3#�% �L��hJ������$�b-<����V6��M�6�t�]l�*s9@�C�v�{�T3^�.�����=�C5|2���^l��Ne�ޓ�5���X���;�!hT�a�࿨�����%��4tI6h��=΍��������4.s1Ovy�>��Xy��S�|���������ˁE�����h�R^����7(q�oIs��s��j52����*�[E3�X\`�I��ޞLSK��~���$�ּ�.�FQ5}��hN5�/4����1A��ӽf��v���IK��xm�?_t�ɒ��9���"�FL��?J���G��{@ Y����-
��"w�FL���}��wA��;����%ɶ�=������F����qVn�h&P������h~��5*�s��.���Wx�r�<�/���@K�~�l�L�o)�%��6����h�}t#J��`�
�����S�_�w*�S*�����{�3肜��.R�O�rF���{D����or�c����/:Y�}j&}��*R%�@}�ȳ[yN�#6��[��2���q�}XqD�.�/_��.7���9��1��7i��4��n�N C/J0�[8��T�k/\F\K>e��,�f�Z��-�p��/!?E��G���M�P���~J(e2��*�@^���bm,�=�a�P��>q-�=5��"�yڸ��: 瀮�T�?�P�> �Lщe�D��$Q��-~zl���?Pd����yTsW?Q&��҂2����K��-/I����ƀޱ�@ӯt�H|�8� �3i���9�cظ�<�,h������ �X[�����p��0O4��7�.jvG��=�!�����HXP�i��2�T�t�efݷ�t�2T�����?�/+6����m���a�v_7��+����d@�/��H�����H�c+r��y>nY����5q���z�(�=�#���p�����)эjōL��q�{�O�N�
C�k<��/����r
��t�d�\�F�pA�f�%��7���6b:��0n��zGI1��i�II{�g�L8lh����g�x����2z$���� R8ޔ��`��Ki��h=��`�J�ޒU7��Ydб�{+���l��&s��[v��F�k/�Dm�Ј:��6xԛ�n_� <�	���&ͫ�N�vZU��Ѥdq��:K���؊�W�+�I3�P[�g�@<b��
-Mgm��`-E�&ת�	h�P�ϻ�_{b|S�V� ���#0�0�o3&ǋ�D�]V� �B���<f'��s_(�9�����<��F��)4�-���ط�5[����?�R��ȝu��H۰k˥��:Y�u�t|b�	�ټ{��;�
���/�@R��ރ@:m����Q���F*'e�S�L��~�ћ��-��%UA�׋���i�g�S�ه��*����y��9����)Z�,P��}���*ߊbI�����[i#�������g�	7�#�>�x� 4��ph`
��nI�
�B��*z���f�����!�#ۜņ�6&^���a�����wY�[��38����@]��(%?�q�)��ź����ۤK�Z��U�'�?�4-����ek�a��'+�qkm��������It?�h��ؕ챶�����٩�n�߹7���p.�� @ΝZ�1�fB�Y	cKt�m΋�$p�����S�F��/�/��A���vd�S'����n�2�gB���h�HU��'�V㥨�F��O�&#꛿��=������9�_#���K'�@�˖@�~
Æ��8�K�MWj�h��T���������
�>j����_�T�!-�2P ZƩ���O	�1��$�Qfq�v�@[K�x��X�n��(�F���Dmݴ��'���_x<���=p80��9}k���'���
�����2)�&�P����b)�yM���ES��u�
���Y�p·�0��D�[����-��Z9�OW�l�p�D��W�=�:���r}1v��oj��;s�E-���Po_�]�\�m�����+�h���^>��At�����)$~5���'
^��<�A-�Ll����#;�c���T@�77R�%GV�й�!4�p�Pn�u��4a|{��"X~�`�����"@��u�����ɋ��f��r��	��W��a=a�!�jB]ĠH
�X$d���+6��ya�+vc9vI�Ul;����5P����h9;
��~�Ȑ)I����c�?t(B��0h��C��J��lKK���1�o8ɠUO?E3�L  S0�5nѧ�5f��>~�c�G/ȼ&_XV�,��Ґ��m*�����:���	�>��R�h���j�[�b��'9cF��÷،6P4�`��;�sUu��]%��(A��|�)vԂ�K�<b��*sG���١ahC�i�l�Mt\`R��tȈ/� �`�c�W��e9����D���Xk��9"d<�h�@^���Mi�tWͳ��Y�:�ʸ�Hg5-`���-�&߆�����[/��:��6MU�`6�*A@�ZgW�i^���k!���]ޙ>�=ulQ`���D�`��}��`[;�{X�Z�:�_hɍ�����9���gE������	�lF�)UHs��A�w�Ho��NC�����6#�Lu���]Rםq�.��E9��W$iiM"��9D�{����H�@˜�����},(�k�\xW��P1�b�i�P��x]BO�˛�g`'��[4��#I�~l��k��"�f����t��D1l�P���Z����Ut��m
���J=5��{��S׷���i�bԬHG&,0� ����f)�޹w��T\j��_�^��Lh��Y+��sZ�)�=�#vX;h��`��o��n2NN���������+�+��W��_�V;(|8P�1B#��)��[�_���p#�ۇ�.v�x��]����ذ���P���a�3]� ���0ʡ��[�8��J1V�~�o��i���v�90}���l�@�0�!915�pQi�+��<#� 0�MZ ���؋�Q>ݫ���f�O���C���@ c��Y�*(����-�x��������eЮ��(�]�: t����@0pa�:�Z��O�#�5��x�!�r,��*��*_���=a�������(P���0��2�WLzV���k�4�_6�dU�/�+e���۶�<ܥ��+9`_�&�t�E�C�(��wQ�@��M���VS�Xԃ]�3�t�j�ı��s���hNB"_Il�����f�SR�{b>�J�
_Μ�~���\{wL���1�kW���������!��+ Ebb�͇bG~;����_���k�<�PC�=M�i��mC�..����DZ
��Q2��1揿o�� ���{��NЁ�L�)N�.�Ӡ���)�]*r.���� 5d-8� ��;��s��������^�u�]�� �O[��W��g���W����˖��u9�nI0@9�et~%���e8����Ĩ[�ƛ����'���D4�	�V��&��	�?����;�C]�z����é�%�m���[Crɀk,�z��|Wp��_�4v�jU��xH���z�4YM�Z½)d���w�D��\����8#�}����!��F$b�*g�է�������_�;T�n�~�����eF�Q�ƹ�D*��S�J�p?������X{�v����׸uȤ�_;FK1mQo0H���A�j��b?ۙ�����wv�r�$�/��FG��	*��	N���p�_|���S�X���V��ܴU����P�&�}�D������866MM��Zl=�lUs؛k�GUz���>����c�ʜ�#�f�8Z�@+n�е�����Sq��"=�8I�w�{de�6f�T�˘�+="���:+,-��㇒�U����;�<���o$��m}��5�eF!�9������fΚ-9�r���yEM��z��L9�.d�IiX�j�,��Lĺ~y���o8�Z8�$)n�P�V�9�,>V��3�������@���(ɟl����Ι�ӛY��H�k�Z�%A���Kğ3jp!�1���0F��j~O�G�D�->�
bE����yǺ��f�(�Sx[x�x�BJ���Z&I�1>�k��\)��P֞��a0t�iٞ.��-�t��6I2�L�]���ʘh�|T�AIb�!ڸ_�A��\RT��0��B�r���j����[��{3��w��D�
���$�^K����+��;P|�8j��.)�����_`�c�zm�Z�E���E@�a%z �����0t�z(�W sy��>��E�d���0�f��{�k���N��gQ��9��tX�<�
-���Q�3w��E��7#f>{2A�\��'وe���(jg\BI�"Q�h����S�t��٩~l�T��2�g��#	�H���ğ����k9��Ӎ��_��)�x$�����f�/�(�d��$db�����3#(LW� 5� ��e��e���
Z=l�����3�g�m�����'�6ϛ�ڱ��Qi�Qث��'_��vxZY��wQ�OHM	�2IE���^��Z�Yex[������N��R�`+ͪ�y<2��h�����ٸ^���H7io�#>��T'g�@?͊E�yI���i��_ w�s���i揬��~hn��a���콁�ﲧ����+=� �w>�Aja�&n��:������f t;h�Ͳ �[�qw��Wk��f=t�������y��8�J��\r�;��������I�ۏFj��f�D^���3� "�����`��TQ�\<�I�R�
b;���~ߔ�QRwP�E;⠏颿�~�)b��A_C�����q�%��>]E�%a�L#6.���X�2Tz>����]�>�R����`�9���wZ�/����X���,q��MngI�!	@m��w{ L��򞞿�� [f�:�V�����d���t�Q6y������P�Jz�-x=�w����, �^����aW�5��]�#M��)���]Pb�'�=F�[���1�u"��.m�Nf�8nit)8�]"���`��ġ�-�)/hƲi����6Y'��`K�S��c��<9�Ev ǘ�:�-��J��tz�1\�%'���G�o>�G��>�w8o�⡖|�SY{�F2�����C][CJԽ�����Y@N����{�aܻ�r;ͪ_[�N�zM�@y�쒹&	���<Sl39�ۃ�P�.�	�[�3��F��Q��ݙ��)x�,�|n��-ܖ~V*E$H���5|����RS�#/��E��*0r�@c�0g��XX�q��0	\��`��ʢ��B�f�`���3����ߝ~V��Qb5�.���v��y�qD�A���v���A�9oF��a?nҔ6���<F	p	t��C)FK&�o����A�#dp4 �+�4�G��O?:�OI�ȃCz$ث�f�T�-���;V[��]�*k]#�)�[v_��NX��Л�4)L詞��:��BL�7�����A[#�뿤�dT������즎�4pA̻�lA>ˌ�"s:1(,����C�x�����7�y*���n�o��~�#�J�<��|5���4r���*���v��5�9�w��N/Xw�TjZ���	�a�����^�^��O$q�'q\�牼��1�[70��ј���ͦ�_�(�w;�v��Q��<�d�!��x'����E1��j]���E,���E��Y�,k3�F/a��]�E����	��XTZ�t��Qz!����C2l�2�C�𨯽+v��zB�%��D������S�\5�i2�����-�,6ɇ�s(s��ʒk\I�敶Y�d�[�EJ�r����o��Zk��ҏՎ�ؿ���e��:I@Ė���d�������a���\����Z?��=Œ�r�J^'�LtR+"oi*!CiT9f�e��K���j
���'ɸ"���V�f���?"P-+�����Cy����!r]���&���Ŷ%>)*� ��N�Tn�����pk�L���$g҅�m�,g�К�kV\��^tf��`T�'�p��->��kJ�E`�q��p^��3?��B�;�� ����7�k�~�>�����6b_��JY;�c�mQN�ލF$��ng�|Srձi��L'�  ��:,�p���A�g�a=M�qecXgtҏ%��]�p�8�^��)t�􉣆�tap��n�: U�=p��|͉T�/�]n�?	$��6d��^��ae��v�p�5�r.c�z �����\m�@�I��?R��I٧k���E�y]�]�SgY�okR�
1��9��}����_]ū)�fȠZ&�*wګk6!�+�z����h��n*8��oi�� �[А�5�K�bͷ���Mk�r�u���>���]�?��ƭ+�'���$[[>�w�R�G���1�����G��_�%Ih���襥t$ê�І� E5�	^��̜z�~Ṷ=��I�*�i�$�Rl�y��)Z�L͍k:"�����[�97d+��Poȑ��������B���T�cЯ~��6�1������_n��LJ(Me�@�N����$��j�9��B%Ol祐e�p�'��XW`F������_��{[O��}���*�n0�F��T����>5q�Y?� t+h1#�����w��H��2t�dE�C��P"������]�ܝm#�ir�+C�=��������"�O^0K$������P��
�:ڬ/���J�6�Mg��}�^@R�'���]AY��j�놉'�ڱF$�!�,��};��ƿn�Z�	�E��0Z^�4�#�mnF���| �S����j��2��T�����ޜ�k�F���%c����!���8]� (����4� �ffW5�=x+A��)�,����Y.&���2Y�������3�Z�4v�%]f��Ț���v�`�ݒ�������%Kg.%(u��hk$��h7ӵ��T]�ETz�R;-���_Y����')���fxh�8�����@;����3]��]z�����Tb��uqB3������3�&�ؓ0���lM��V�Fj_� w��(�����^a�����l���J���C\mOO�|*<ᨚ�}96�@W���Eq�ҼA%9I��֌��[$���8�w)�\�8����E��Eї�TE3N�1B�4V3�]��A c'Q(y�	E]��}m��Cvk9<�b�$I������8D��_-��K�$����9��=�P��F�l�/�]g��K��P�����[hp+q�8�ۃ�*UĶ�Xe,՝�Q�c���m��?k�y��a�>�0��) �bV�������8�T-&����O�R`o�?\�Ow��6Ĥ����.Z�2	��������9	���ZJj$�Q��j�'����:�<Ȼ��0�,3뺽�}~L��V�'Z��,P�[<y_�!-{�O���{QF	=h�����*m����j�|�32	�j�}	>�y����R����N���oA�gPpu��~� z���4�cJ��«�S&4�`)^
���w�|��r��=u ��=q͝�L�^����Ϧ�U{������fF��f
ά?p	�1��>�Zښ�s����^��~�����9�&2JuЎ��UGԚCO���3=^�6*ġ���\�G4��v�)6��w��ڼ}c��c���61$�#���gC�d?�S�m�̩���;���7��/3��d�k.*r�G/�,�A���-qm���Nl��W�3,Sk����1J�χ���2�[�����X(�/z�ޥ���c}heoZ�	r}\Q8�H����CU�FN��1)f��K�N��*��od*�ԳaΓ�z,��z5�cr�z�.V��iفV����4G�G(��O��f���t�ĕ��n���Д�����lb�����iϛ�uvEQ
Д̊��6�=,",�O{c�T���7Q�Y�J��4��H��o��`ec�8��z��z%t��'v�LVo�Z͆c�>�1`vp������a{�$]��&!��܋�zSy��j�&p�r���0��oׂԔgk�avz�m��]�[lz]�js�Ż+O�59f̟S�z���k<��U	:�+$�*�@"��ǋ���D��;K������m�St��~Mu��}�+D�b���2�MwQ��/�<A�:��K����$I��!��:���[/vђ@��/L	fd_7%����}F��-��9��2l!yݩ-��� ':�%F�E��v�)��o웖D��~�j�sI�W��g�>06��p��֚���Jp�y;�I!��8�_0�H�Gᘋ媬���p��Awн
��`�����e�����2�ȝ�������2��[8+Gi�Y[P�)~�6R-���%��c�Њ�d��H'îҖr�@�{{g�֫$��_e��a�tz��S��Qs�A�7����U�%�b&:t�[zK�k5��r���n��^�=o�ȟ�h���"�T���-�u��I�b{���#8ܺ�B���1e������u:�ZT�5��K|B��#�{�9\x��%ΪkM����gJD��xP���%R[�T
���Lz��E��U�8�Z����k�e����F�G(�/X�8ӫ=�x�Y6/����r��
��hO:pS��ޮ���VJs�k��qT�����~��s�"��OX$����l�iݭF����t�w�@���KX�Ο�\ڠ�b�̜8�}�c��	�Z�K1f�m({6������s�N���O�_5�]#�<P�S�b�i^�0�xձ8��zlޡ��YE�!��m�ZF񎼾��մ�x�YQ��O��]΀�����$< v�kwk��H��&s
�\����N����̯cU��'���)����o�cS>:ϳ�YzǙKi�Y-�j���(W���v��~��4��ch���`�J?��n 1K��0[��zPo��f�7�	�3^�kd�2�D����'8�~8�S����2yv.]�τ�WO�}ڹ��=�S��C;��P���?a������Fa�Bn�n�>� � u,۔�d�c<p���S�.q}Q�g�NIʍ.z�Ɣi�nG������bV���SL.�f ����ouc�����8���t�R�51�;q�B۹�F�ܚ�؋�n�ZQ�/�`���.(4�в�GH���f&�����gQ�m:�%ؾ�)Ɉ�]g���>4\�ACt�[��[o�t2��ܲ����~�����Y���[JA��k�LI�Ol<��ߞ��p2�]0)�K9����Af:��%� � Z�50�/���0�x?�S�^b?Ty�����2١���[y�Q���^��۩ |��2���s�-��zRD-�-uQ�5Q�/I1�W�2Y��c��)a3��KFk�bv-q2��y�۱���9�eq �i��i�!�Ѻ�҇���������P3~�<q2���xyCz��ϯ4���\�zI�Oi!�-V�eV�6���|��r�/�3�h=�������k���Ot�$#G������Ƨp����uDnҖ��x��$�o=�,At*�Vr.�|Q�� �'�$����@��D,��� ������ڣ��"/Y�O́�Q��["�|�T˲V��N&��޶��G1��?(��K5m�$bp&H~䴳�9������[��Y�9��ɌТ;�$a��d)�t�9��ɍ{�|�z!Z�̕\�џᩰc-?=�i��`�OĞ'dBV|����ԃ��btpJ�d��i0&K"T2���F,��]�s71��GSEI�:%�pe��h�BPOQ<�a���Y%�>��0#ۧ �����K�O2�-�����GP�[n-��,g��t����O��ܶ���w��$8^$x!��s7�W��n(�de�[�io�9k�P�t��`�L��cg4��&,H�7b2���T����0����S�T���]��G���'^�L
�"oy�]��%.��fSG	�S6��^����A!�O���ق!��!���<R_�??JZ��T'z��^-t�.f���ϩ1�w��UQ�Z�&��MdJ�n�2���5=�$C���罬��j�$�3!�G �
���kC���;%�$d�B�������B�Lʒ[������N�a��1>M�� �?�Ő�5�U̖C:���̆*s����u� @�S��f/BP|\g$ �k��,iaT#��]�W�@��N�+3�(��A�;Ë�/���B�݉0>D�¹�K�\�|��㍜Uo<�o���ر�g΀,?�4���T:N;��W%�W�KB]�-�u���%�~A{��e]�+'X/����ů+7ڑ�6T^����7U}2�Ѣ#���J&j�����T�� 嶦�{tn�m6ߺn�k,�1�,�o��k� ��>���ʟ
�栿�61��z"6�2]�Mx�F�n�u�����p�C߶���~/��6��jF��3§NG��Z2}f��uaK��e�c����{i�X#���6��۟e-�
�"�1��6�~i[�(����D|��r9�e���x?��d��ν����7M��SNGe�^y�@n���Wc�n��>��O8�:�Gs����ю,d���� ���^��;����O'��j��|xt���"���{]� �m%{�H�=):~��ɣc��A�G��9�~�VC}S���
l��Jz�0��*w�kN�,����l��̱�tػJ�O���*�LFO�A�.~�W�+��I�T�V�[�)Ue,I$.�a�c�Y��p.�c �.&����Y����
�t���qiDp�3e\	���?�K���(OQ�+�Ǝ�c��+��J�>޸��ҏ�d���k��y��ܕ8����O��y�Y}���vT��x�l�J��tT+��#�u����3��.1l �����'	�2���A��jjߣm,t�`��W�/ ���P�����/-�;`�K�z�B�v.����^sI(�G$[�Z�ǋ���RC�Q��&���BGh���Z��hK����K��p���B�L�Q���EN�T����<�����B��kj;*�>�[�0E/&p�������
����d�[��^Z�M�,����õ0 ��j����Ѻw!����FAc�C�J�����]:,�߅@fE�D�vg�WH2�C��f�������9]G���rR�z�������.��|~7"qme�{A��Y�Ŕ�|�m�q��AG����A#����0�3y����f������:g>MS�	�@>�י{��#H�ڗ�R��|Bq1����KDDȚ�n/�E���r.Rɍk��T87�U>ρ�3��GO�<���08�ȚH8��Su��Uh��������da���l�_Z+8��(N?���� v{t��R���BO��1���ƭ�����rzi���z�ř��+�QB��C@�������M'���i��b��E�|O,��e��G��/!�D�Vq�#;�>l�U2O�k��ۣ�%Ӕ���K-��У������3f:ժ�Q���c�c�Z<�}xl��4�Xx�?h9���S��่L�0������yf�9X݀�grď��f�_;sUWO0V����]�$�<��P�c�Z��L�ش��Nt7�:+D��2��Voξ�����[��_�!.y5f.-8 .A� �T��u��ugdg8b0YR�.�:��1��9��;�+���
y�P7>��i6��� J�7�ܭ�ͺ��;�Ͼ���4S�_�S�j9�Y͝s������h���l�D���]mA|����X����薂�d����^;dWg,L��;��i 5i3��������e��<�|�W�O(!�y��u^�v�'!q��i�c��B�&��|�*�?ž�Ht����s��L����0�,���j!���Ą����!9�ӘB��w��~�)!���5�����Z�#*k��V5K6ǽi��x/[���������r�t�(]1�#4?pl�(ZvU�)���4� %N4�hQ����8���1mD�)?��D�DZ��^b_-wb��"�0_������ձK=;�)��;\.\�Z=T0h��f��ܓQC��ޱe)!=rp�t�u�?��h�:����b�8TJ��=��^V�6���<^vQO�a���+^���'�fO�dv��(�Wn��ܭ�uƷ	��<�(�$Yޗ\�lTm�I�#`��ʪʛ���_T�WY#N�פ}���M�M~��y�C̟�w���R��b{;��=ܸ8qF����V~������
���m�@O�U�<8;���R�P�8�^w�`�ĿdB
<���p��r��l�م���^�X�/"����n�V0�(���uwMa����(n��8Nϯ*W��X��,��+aHf���Ȋ���3�K�l�Ep���Y���!C��GNF�S�$�p�$��y}�)�^L҇���B١�V̬g� �3N����,rY�z��iy�ৌA�N$�N�^�M	y0)f���8>@K5��ln\L��8Ե�s�!������an)'�ȷvZ�����xff�l
���}vz���/#
�E�fet9�sKB`�����Q�F� B��@��Z3;g�(�҄���� ����w�{{h
2�u�;X���^:�U>3�.�G��HIe`��_r��J�$����a%�,"7%��7�������qB��������/G��t�q���f�xM�-��G�AYw���gq��^}ad�L	��`q~���a雤�����q��L2�%���k�!�rsU7)N�l��a�hE�dD�<p�md^H-[ˆ,a.�����kOz����W�e��z���B��ꅃ�Bhb�Y����O��n����=2��A���D���ũȦ���L��~����.�Q�[YO94ԟU���Cs�z�:��`-&�>��ns�3z�x������6����P'�4�	�pT-Ī�.�\Y0��q��_�Ǆ\?_ր�?��z|�H�_?��w��~|JHs=������&�Z�����-^_�$�Z�>0�`�G�ezW���������0驟���sTT�>(\�)3 �9k=m9PY��۝̦)D#e�'��m��.�g*��q?�	���4P5>���Ѝ���
c�Q�_���DS��<nȘ���n�`=���~����?�v)�7VC��X
�"!D� �+�ӉjF��.���]<L&2z��pT�q��Q=���Xp�+�K}�֛-VB��v9.��W�k,�h���
.�B�+��h���E-�]�@�v�On����y��c���~���a����U�]�]���N�Yi
������r�zZ@����~���4���U�.������^�����A�D���n��q)?ʗ�#pBxT�)��=��G@��R_��J�gJcYw��gX����/�0��-ЋH+�,�ܓ�RO2����-�9��Ҋm	�0��%qIt�D#��(���Y��!�_�0�#�'�NB�����zA�	/OѥD�@��:���n��֒G��fxL)�E�z�!�w��5�����1��P-d�nj=$��������W�c�V�&��X�63�*�\��:ؾ��C�R�Ϻg0+uR�@:��ƾ~j��k���v��mx]�$�9��N՞们�H��hm����ՙ�"Ͷh�r�j>�z���JL9#�Q�~[�u71�}sq���`�O���C*+%�<J8����S�����k=����	��Kx�Y�^����w���mh��ybL7��
�x��{{[���b�;M��J�U7��1�<�H��f۫�΄�[�Q�DKٿʢk�K`�J9y>�G7��	�%Q�,B@2�S�M͗��e��Ս3.}�:�F,�\�p:�N~�I@��\L�y��I)<%A&d�"(\����2����#�
i�*yD�c|T-��n���4g�r����Ymw��o٣�>������\U�5��v�a�}T��-����TQ$��-$���J�v��xW��ӣ�����x�`�E:f�g���$��=��A�j�~��tc`�kM+6�V�z�g�� �4|��o����~����0�'eh�2�1' !c��c5B�=� �a��zb*g�=�|�WޡSJ���4�曣$��\(t�j�R	�1��mlp��{��0�CYWVc��"L�zZ�蜹��1��m�S�\����F�_VsD� ���>Rn� (b�H����Ɇ������_�R�{~	���t"	�A�\��'R�"��
mP�P|� 	4� ��vlY s3{o���V�#����.ފ�-4��֏�q75
*��坟A᤾��&_������E�Fi�2.�>�{���1��j���k
�g%�B���y���x�N�cN�)į��[�:�ub @\.V�e��̟�)�υ�c�}Wz��y�o��}�^�ɛ�,�[J����ï�Y�!�>��A_�����D�ʶ����&ݣ�����fc�|�Θr{̻���͈]x�QF�5˅����L�\��>u-<��3�\�>����K�M�Gvʢ)�}"���ْ�.$q�% Md� ƞ�Q�����k���;��������mz�iX�nL���i��y6sDO@�˭-�������C7���!��<���-�&��I�˟\m��:�W��3����K#j��[D�ܗ'�|�oQ�,�_�3�|��@��	�á�°@��ܻ��KBT�0򋱯1�Ј��yI����l�(�~GaC�ޱ힠�s�V:��D��=k�� �yU-��[�ʻ���߽�/��_[���>��~EZڈO��Vw�R�r�]�t��L�P��ĭʄX����Z�o!���u�E�V`S%�08?�N�u�Y�șz��o�O;�x�<aG�8��2��)'��CgVW^�>���`�	�.#zuDŔ����-p/8�p���J�%x,7��&b�+Ɵ��bDC����V�@��0��҇�l�h��j�!��r��K����}1R�]�r��2��,0+�'�u����V�y��.=*�y��0Q~"ˡ��Ɇǃ]�U����2�����m�F�*"�q���>�ӈ,���m�h&/��*�팏Aɘ�����%f�֞,U���B�ހơG�{�����ۊ<ȏ�8�v��No��D����f.yxY�o��0��?X�@^���9P�اS
uL�'n3������3ݏ@�|�[�yvF����C1�Q`��Ґml��
��cbYp82@�e"�����/]_��;Z7L�ds��w��5��SЌŎ��l/��U�U��_J=�]Œ��o�p1�r �xb����P�%�a��M�'���-�	ú	��B��K�*Gܦ)��뼨c�F��:�.��L��GvZ�bR��uۆ���[����9��iZ~�U>����ӳڴ��?�ap<+0�K�g	�T.�\��5���!�f���l�$���\��S���˹c��X�Nl'��%^����]�E��|��X��\�R*�-l�rDM:�̌2.jx$�Ā���V뼎WIB��p�C@��L�P���-��ޚ�Uyp�qWl��kx��5��h��*B�ձp<B`�D���1N�q��O�H�2�����o�1GT���5�����>˔�Hi��\ ��^�z�ݛ멟�_�R��ո�m�-�:�F�F���C5�4�����������S(�k@u�d��F���\���LRN���P�p1��D֏-�N�q��{�0ƙL�1�F�4\Y�'}��3�`�������#k��x��"�,~��}�:V*6I������q,G�A9%tŗ�;��0�� ��;�#-������I�-v�m8���qw��hF'f?��5�+����Џ.�y��)PGP[��U�-��Ȟ�!��YG`����a=&����LJ6�;Q�����`�X��k��ƣ�`�;sC�9�w���-�y��xn�ltņ�/u�Z�?cH��m�1m�u�#�4R�R5�z�*ȅM�/�_h	%2#xa���ܲ{�`���E�x���0�]إ`q�Q} �qur�,��w#��+��Z����0{`o�k�cv{��M�Խ���~#��+"�2����T6����yL
5`�T��X��?��ʩ�F��v�!��~�F�!��e�)�~���)�(���J_8Ig��k�Ui��z�����?���^Q�ҡ	b���_��v�����<�͆�����Հ�]9br�P�C�pw���.v���dݫRD��ȧ�8?��E��>�xρ"SJ���Qh_�O%��X�j��:a	
W:}&8�(OE��I�l��Qgu��O�|
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uUppbOwVST/uo4dgs2TlOO3a8r12qMmOAvxQpPkGTIGb54krruLr01IRN8ZlB6ZWKmCnCcuOUH+L
o8lwtDewJ8M5E4U450vJvISWXVsepBi0Mn7jB5cUy3iwtjnzzU7QMjR1ck14yhaHs+5Vw84/gEFH
qaylQod/9Yf+lygMSIMDAw28ItwZf+r1auwtw2PgMW6C3Na4SNFZZStNBaXYXDnvRwIt385KSPaI
iAyDQCvnYcX40UzDrprkaJ8+1WxUkPhgAWN/GjvUdv13+yQkFVKYQ06vlSG0gZ5dfcxe8WxHIRGu
+9X6MFbSfwwMkqQRN/XMUy6yDBzDNPUeAUkEJg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20544)
`protect data_block
N+wK3lJtp3a4PW148APEaNdh6Kp0kWDvKS58yTQzPqcVQLiAQQZD+BKcb61ngDNOxT4fc+Iu6d0s
boupV9mJduf7H1oVRedxZYjLwr+nT8dC1+6f920ghFgT03YUJ7LZlCpbxnL7CIBAhEthjw0mXzGR
NfXjMRtfR4SDhdECrBXiYgnbsQe1vf6+HxD+iMK2gbnohVkD7MTqhFLFo+FJN0WFCsqtc3PTck+V
uwfv1Jfd4XhXIvYZrsn6kepQW8nGJ8sziuePRebNvtk22hsJ8BDudRoIyn3GNlZs+3NZ+WiZcyOy
6Wkpn2DEgnvLMbYNOSwHyUJNf+4cvQbXofJych0NMshD3uzA0eqGPct6JXSr0rFjSFnytUScsldk
Un+xbmAqoFUd4cfSXpwe+eEc7o2qJNvKE8vtc3i+DMOdcjNLlBRTuHBOyQUmHtLUJVSLCfhYJRjy
9fpStYs4B0Dg0SYc9ue/yexhIgvVesll3ZQ/6OvcCh+xaRILkg22N/J2GOsMT13wakodz6FbxqUS
btM9XQFBfC6PW+qMSEeWFfMmGygXmsenomiWbNomaSBMAMqe3/JKIgn7E0IpWAwI0pNqZJziclxv
LRNqjOHxf3PeQCPGMr/NV3LHBXaODsi+7lZPqBupa4QWKk6PNWEx0oy4UnwLuruXKfQg5aRdbyzU
du5TR/CHMLRUCY4sDRCeU2SGQyUOXqm0aNSIDwBDntEOBcmTSj/slm4JM3IAV9KXzXVjGwDaKbW6
fDKgTdAmw440Gby+pejZTD7OuaSboS1XAAIjpD6RiJ1MBX3tqlhxNEC4ICDT24ptGmV40a4nuOc2
b4SRN/iMIlwLVBw05Yaui7hDjQ2b4qmWyuYTb7XPblAgfW8ZC6eiqUSRVzykwYq/NvIMySn5u/XG
M4QBF1+WECCdjwHGhXUPLzojptw5l1siI5EhEB4ez0pGVwaWjmwFnO66anqAEgZT7CYa+zs++7Lv
g0iKul+2XKpqo27QlTqRXbRVouPygCSYQBrgb7/D62atrDBKlEqZKVRcNJWObEs0b5M8EDmYaG+3
ev1NqAyWewojAW9nWNk0OJNRFqJvho3i7bTmvmGpUB0VtbpF/R4gfvpIZf5pOjat4SrFq6EkLNJX
nW8+31zQ5LiYZJDY9zgbGBSE7wzG74eTndLgecTOF+7CedejVMp7XUbpm9+ZRRcjMkJD1OKL8vmp
YzXsW6wMoFwtPPPC3QyGl2KGYWtNDa4DRlSg85VrkJd8IvYB32ebtoRvJBCtDJMPzee4Sd+xCGmi
h7Sz6KjakXRhzE1bOkw+VqVIoDDn9c//vrVHEba/n1OKW0+g5wfsqj+ClXUaYbLYEc4Qbi+54H3N
qvWYRxDHn3tKDtY9SU8QzjTYPucicyuUE/xA/PtFokYYOSlwgu7QAjCdmyeH82ZDHe+zRj/vIlNP
+beZQ/Z8v71UHmWJO0h/QbFwsJiRK2RtNHjyOx/OpRipyRHq4tNcVBq36UhFwPpBVzQthSKgaDpr
3S8kdeMwF+Fyr0oil8CbMntXbRnuDaGyDhs95yreUdaOsUlMgmmtFny+f7lUjIbS6cAAmLCAfGLP
t31FXxLaSH3BjjIrwtdxykcH5EO3IH78l8MLBEJGE6GRiVHJLtQJEet7FLodUh/HlQ4L3Kq8FIWp
iIuuAxW0Tb8671QMmSKWLEnZZoxVUO/1oPjNfpcYYUlfxQlW6jJ//rfTVFqZVosn7EhgRUVYdRx7
zw0QMPA8u1ZdpqMviR6aksdb5ywd50lB0aOUO9J4S1TI6GryyDkHCbZlPJ4+WOKqLt4xpj8hTpRp
qm/AC3HxRc4q6jCnbyHbykvUVRmrfw9c5LKVDWyeDZG0z/9Pv4yRibUWi50foeqnRXd8W7UAErL4
vkvomgDMu5/547QvY6C1XyDBzny71ISToMaa3cZs1H3eJItKhaq1hGdMg1dg4JVm2AFXkZCitOTx
oEwSxVH/z+XLBl7UKdoLseKL9KNa8QVQp7Krfw9Mjxe4A59/0oem/k1PdPnrmmxktsn7AFp64UjB
TjftRk4EktV/5+xulRzndOsyMDP+QqcqGHKjMdNFvY1bRDJLf/MNQ//Nz2QbzS5FTGjwCFmDciTa
uiPe0q2sjetMUZbqlurmlrYB84iHTl7SiWBZyEgLC6sDvHwHw0uHGs2Y7qqoYp8PSH4FM07eqBDN
zRTXV5WhnoJ4st1k8rEkhjCRGgWJiznwIDqykKosXDk9NBsWW+5UvwAoffYzTWRPS9TwXXlLkAki
e7gQBNSP5bHkqOCPUVtKjg49OfjbOghYkuDCpF92rmgKBBRybn84yJs3/VSt6DZOh23RNuiNu0ti
03/NyhRhxJaVi6Ce4e7cPYzLJwZ3SQtboFwnxjNkcXo402ls9VQ7ImtddoKPcQGJlZhOItZBVhdn
39UGnZKhu+iE5goscS11rLMwYLzT/b90fsaiAwRAo2Zl/nhQjHSRvPls+pHKOa6Z3QTDeqZDjStS
fp4ouIeFXw+9mPGDe/4ekyaxcZ2Vdi9bjA+53x7btnzY8t5rPsm1TlOE0Fli0ApF/+8tdRxD/Ekn
ZpImyDfex2dLogbxCGIp7XCpRIME7XLQ3QjZownf01y88a3AGYPFzFfzIdVEU2xCq4r+ibL55koj
027uUPht9vrFTvJgMYYf2LhzxpNxFMjOnF/Sozez01BzmR+XWq6MtxyWd+ALfX+o3Qubwjivm0g2
gyic/tGmlVjTtQEZ3/7wu5jI8tSZ0Yh5yaQ+OgfDvW5bkcdubE6di4LHvLJV0W08hdydZDJXHxcZ
A6gdOZL5fyz5BX2mbAJoiO7CtVubS1NSm/jAh+MTp+KMU7iN+tDmJIZ1HGhpheHs0tmcVBm7PYWA
dmwlcFpdjXR8qHtCByseOSH/imj19xtl4L5AMiw2C92NxTeu+qX5aSfyj090/eGlkhDpqcmfsd3z
RSOZeK75jeUTGHLTC+yQ2p7GK7jYprVkI4HZdUdTfm+OmEn9NxHkSTd/WQTrKhCJP0kOIEgTGJ69
+MWCm75loL82iw5YjTa32sorrFXW8WNC5yKHb9ZiuCXKXyW9GUxZqWsu5afzlyTS5loKlW/PE+eT
6GWWZEiGisJLHFPrR5WrqoH2lFN/85jUrO9N/jBO/1mWIo+c3BLaJMrIvZ74GLHjnuRGQMjoh/eR
NjQ7UDoj3xQBEWwgydOZkWozzvNMO6TGekEkY+9WZOWTokDKq47LEtO8ZzVkoZOqzJxfffbXMp0y
Rteq6KZ79f5wpF3TNX7aBNF6Lu66VWzIIm1E+n01kzAIMYWwcBxQwhnkWtkvk3G8RHo6GzOWZCpz
b9g+TAbhjFcDXEtskZKNEwei295ZYCN66IJM4h33JspAQy2/ilTRSovAefIL0W1Ewfi56jVYtOrJ
r19Q7d0hux3qN/oAYywi5DjAvdYA/UO+9hhjNkAJ/+L7cNNuFwLFxd8c6mEXDD4PgZKFMtgyzh0b
fPir78/vXjM1Oyw0wa03WE6eI3hz6XyxE0Y52rfTnStQsnNQeVx71lsipTPolxkDdR1ObT9KFC6L
cBz7h78D5Y4RnRCH424J5ZkvEueq1zSMOn79kWHvzvmkmUE3DWUBYF2tFF25HeZJGlpEu0Ys2hb6
hPmV4njBbGn6zKTuBRTszW3pHxnb+u7EUAouXnOZmEzolYZ6oRvGVaQl5D+Q2A8rGjrdbt+l4bcB
+2Hthot2ZJBPdxsyZbwmE383jlUrWjZMvl+vsT1uXhimw8fY4FECGc/TZ5Ks1CozkSeTzERq6lcq
K1q2G2BgBstGlXGcYmnzS+UiIAk7t1GN9KIk6UTYNYVbXDf6WQ2P8teL0TCdQ+GpG2gKb5nPt1Dm
HI+S1UjhXdGKbRK1QnRzcJUazaUX+WhAmwDkfDQ3frlgDXuRCGum3ISAmihxe1c/sHOaDYaeNp6i
1L0U4XfGz3aL22HwdHJYlAONhM7FBx5NB0yn7E8QcrfC5+fdlB+YWiwcHJe2tw5KGhLlf9rWWVMZ
0m0E2gt7/ZALedxIvNiFYeP/M3sdJSuM7dpoPmh/QDTkg1F4HQuSBn41nMVdmcfww8W+luOFo+DZ
5+lySJL/FD4SOYQ+U0R/GCi5YkvgBr0A6JOXlHjQrH1uObUurKp1m3kSUD0I8PM3n6eLbMyC2cwb
QdOtiBf1dH4OdPhqkEUmxLwbO/si22uFTLJx8H5q/aQSXLjAIXvrwyl5TCWEHAkHzLxz1CIzxzSb
zYcoxU4jrwUdDiXkhNfLIN3v7wLcMsjmijYi/gVFOBmhb90/kcHI6IuLcGZdLXUJ7lGsYiZHwvsh
TPGmAvkrEiYLp6eZzK5aJvObZK1XJQtayFY+VWDR0XPSvUN2NZB8xkS84y3vj7MuGpUUmBJvlmBF
EUfj8y53v8MZMjT3zqtkD3oFCDrWBuEsp/yqSpsP1udrX/a5hWNXbFxVizlmcIapq/OPUFNEOozj
ydq3fAyyBhWyFmB2w1wi7vpUMrm4ANW+TGRCnUhshXnqWs57oniHhtB1rfB1cNHZ38KS0UUqzjm4
CQziU3uOf4xr1opAcTBdJR3JERTqTr1b1Dzgiwt+rsU+GfwWg5r+eelFjhi8pSz2Nr/c10rXmuz3
fYwg+PKGGzRXnQHwUcmzpHXwDjR/Gd3aci/rRoqPrgpRWiO1DYAqE2nZ/kiWeYsPzI/t5j2mezar
AnEHmDtZAfriR0vERcDDrTVDD4N2xRazFe5UyapXj+31UbVPtmUPRIiLw9FLLU9bFHDB7M4OsmzY
e9ASDi4oWRyHGyG8I/r7636PKFAZroKJ+agmDjskdNhXqZ+vVS4bA9Hjp7/GaUYFqyC7u6HRJBuK
JDF2AiWOYbmFsAGZ+AEQ0Ush6zNLuyBuCsasEVRoqwSD1FCE43Jp9zfD773+pPtVhTCCW0h+mHSR
cfRxeOMZDNXhB6spZB1mafbRMyLdDYKUos9UBNpK7E/GzL91+y5u10Kq5sBB3hdYDrPaDkmmOWIV
GuJDYXnu8X4gHEGamn/2y15AFsXd6Y+FyWxX6OWxRGlzhSDziKSDh5Lmyqb+ITxgLiufcwtypNPz
mTJNJnWW3+jnuq9KndTH13eYZIOc0CYhxoOfmk9HWCRmKqbv7D8AOZa+ZM0sT860YwuBIvTKj1B9
a1onbPqmMLGfKqKAyAnvxhcaB+3TOPRlAx9xrnpsQGvWYsOBBPowN1N0lGwxxYhFT8sw+YYB/5hU
f1e9bzZmRWQJinTOSaM4uww8CEVDIyoyLklGp+E6iXwDf9fgnHRQX9/bH5s0M6uFu+YMo1NRtAZS
PLUa3iMY8Amvz1puBwGiYFvlJ5uQZ+0ZRg6QO+GV1usjg7XpbBuQJbi5WuludQtxgGkq0u+mJHoB
JhyTQfHeLoGeYvRy035c2QxPPuyPqk9Z1OJRvjnrAXbqHdyDpI+uE7CsXIPQ8/CLgqG5bH+f3ftA
/t/8jkGMtfBod4CbaP3ArN/EUyEejT+ZBgj2JXGsbEBbs/7h8aJVj6LmbTZZHCAJWeYADLZMh02Z
MDdzITl1lmsw/Qgv6TOzfmjt9xR3TTGMwbx/sCtAmnsydfZvwns07wXdKY1152XybBycUAUmFgGZ
XUoL6QanSKK/GxqHzBTOGkzgVxDRdkoRJuDkW//DHuBkjFlcBGx85JMwDb0PyhVyZKAq/sdRiR4m
1V83SncNzqJNcTgm1NLDZyObXnFNx/tBUrMtT/lJPENPxKncWju1X/ZLpoIbzNoM/v42MOJkuxkK
/MKKL7p6Zp2CYhMfizXvvFDmaw68XLgjV8oeBDxqTvCee3DFuHzb62yrUl0yrMMbGXosHwmih8uV
tQlHkQoG4NRld86xLRJq2cF/s8n/W8dmdTDmz2hoRi2UI8Ja3CMqmDK6HMCL/KO2NGnSM9ZgDcW2
tBj/bA9Zb/khJOPxPrWgS32VpYuDU7gs98WnEH+1H0IwA6kPnX/mS0X+hLHwa2E+rHP50SB2mkfC
Ussh6oiivBWoFcq7xqRwRqH24A5rOzrtx/AgqPq+og6HlbwS4L4H1nqEvi+EwyX4tiJ71gcCcLab
N1MexKNEZqRB8NgghwpINswTmlMQ1ZDbeV1VF3uE9kmStRudq0Hf4L1PEZaMRdPPaYJUcaF2kmum
JVsAdXIzUiuq6WsYchrnIouLnOvgbmruNnXT3WUK1H5HtIIoYo3+TG2EpKjd3w1Gd009T1GdMHAD
NwpZfXfbIxfTB+uU3hY10AhmoXv18AsHRSUkK7JRVGMwnNFHJQMMtmWO+KdMM3LPr7g26um7Phy3
uDHoo6qcTcquDp5qh0Wna4lLaDSzSteS8RbJXWjTRts8vMfayNLBbLFdfG5H9QPHJIy0PV7UlOzF
J91zU6KsiujQG/Ucw+oDVj7LjFbJuui1VYFnWWsKOkPbQ8GjlKrXCXUHKYa0d1pDPwqBGDkNJWB/
6WfOufnU5BUJkC+bXcd7aTxqUZpksuH9SmxHFBS7vHEU9DHon4pl44129SVAOG6qr90E53o2/6Fp
JBq+UZeE4uh2Cp3dBzOs/z9y9WyJ05oDFVfw+JO9PrmoXyTHXouq4lCYKkwTq3P/nPpw0FzyVtyy
qMs3hYReyaNlDJMV4/Fjn6wZ5Srqgxj/y+LiDUR8Jv8vHhNjRMoLkvsvXDFqELJHfmQu2CnouwD5
uRfkzpcR5zEnWxzkMubtpt9RWjSeLi+BOKBbI7suD1b+Ibgql04vuHPBwN/DLFNbusIe5kf/KkRt
5HvYj6S/oP8gXcXNNQgqdwbeKSOBxRGQJF2Ys7EIDW5NS3hLnwUM11duSUgD58MIlev3iCBcTwr6
H5yYoDcdcDxt9gcuXGchIB7piRnfQOdfWFI2bidkX39709ToJGjhqKOUvrhGYtgJDEotR4+to4KY
Oek1BzZGGm60O51JJPOAQviWj+qCPKx5w7tFR6nSJhiIFO35bcWDuV6dK29lxg/yPBTCuausDKdD
B5YbiFpRH6e7i3PHceVPJwkB2EnaPdAqZWVbj9bAM5f8y96fvoDiw/1wi75UEhaEZGsyQXQuUHbh
dBy/WxN+MTI47s/JoeniELlM4VZ3ze8uqmU1HfOXQ+g/kGbPYAus7JyaWYL983ByAczz3+w1c0am
huSDNgNLvYZPZEUNUQk/fz4pkrb+fgnm9eyJ5dxipLsgmEJI/zZsPpt44wQeCyHVX83XDShUMWUI
1JxrOR6w69AeuknU0oTCBlIS2LIlTs8gw6yKu6TiZvfnTrUvVhqOd5/ycrWs9VCEfFMeJhWasNzs
PoSYIHR+Ixvqrgifin0oVr1DsU/ZfMt02EHu7mnKit5bsQAh3axEaHRVGf0ynqVNZJlwpArmCGBp
t3WjcnYr+kJrD176GoDx2ibCHrLuufPVzB1Hhv11aV6Y+OYrHKVUH7uiQQwI9VtlNtcqnupekTnJ
KWgdpagb40owhv7sqf34ez/jGcrmHVCV4Quqq5oqhvLPsLiNjDEjI53PNmZ39HUWxjRlTwf9/1YN
MA/g0dMwbXGOrY3/UD2qChpUOkLmbkSaGV8NF4F14DErFrdLWFy1Y1Y0hdJ+vMXvsEycYbRnPveH
pAyQks7sEBBfR+gMcp1p4m5Q3aCHOZbrAR+XBb/HfBrRno5RkZ9HekSWuELzejPyywmba81MTxFH
kocEg3MTdUQ5SqUhMZr8XtGXl04Wvm2BHMY0ow3g5ZpXAAo0e+29ydpu9Zm2S0RyER6rLpzYv9fl
sZM+zG1JVs11TINvlYLFnIDXWVlZYfMfikLs20v0Dd0jGeR9G4q2HZWYkIeI3HpRYdG3Z5N6/adc
IF41BnON3vmyZ4dToReXfZbonqcLhZ/uvtBwGo4JWl8uEXUeVaI7buu9GPsmpqoeCAx9tvryv3Bk
g10l0VZlprDgEe8t9NbDGiFBSCjIkjyuESIOvuEFAGkjNAIkM7gwGzRaDgp4USJykoULqOHpT/fD
NzxQ3RRf9xsCdUYZmQgVm2lLMu28rCO6y8mVJfU8gJAWJm5pjyy1jfe8QAvXt1v1ltoAAo5gVbFu
tuuRRqZa7pxuf2dgIuJJo1+G26dbZ08JCqB5CpH1fyfFzdrGLy6YorwHSlYv43MRNSJgCiyqYsbZ
Aazyj26DFhNaqDxCIB+JbChtYDki1duWX53NMa5FzbukydrcElep19s0kWhLHreVBU0mJh+QVfnP
k0bpAEqa5jOlSA6fR9KxWvRgGntF+MIcHAXkCzOd2vbCBQQvCZCa/yYu5502oF7VlEiEgPKpTi+I
ZkHdlWMQt8AK1vRcDh36hWDvXPL7JMWs0aHQPWeGcYA8YqdZ4tADEB8N1TbKYPxpKnxX24LBfuxj
E4zb+J+zlhW9LkJhLOY5uMZ/Vqg2N4IJeBqKcJzgSD4p6t1CEzYnxzFy4DHaRyVw7JMgh51jNIno
yVvSyArFnG+CRugG3PXeMi8xnB78yM6MbZvmZJG5tAwuUyHmg1HvJkl8kjiUTqUKS5+oc8ht5gcT
edwEq9B7d+AQE3JlG9UvWxzJAU21BlAwr/JK+rz+80XyIcdePiHTFNIIAH9YxqxV61TFevMIFHnH
wS/BGLETdXADYjEKVgw92KienNOhlWhEP++xgIN4gwXGT5+jb/Cpc6jGLf/JSC/oVZoyUn329sr8
xXw0guPnOv0AFxOO0tUknVKzwUcdkxU1iBFs/d9J26f1bfERMDlBSuwcErl+6R8/XBFvzY6LEsrg
7kdMCa82eau20TzWWdTfWtOa5/R4UudbBiTQZDLlHhPiFZdQdqYiuM04Er0VOmZyl1AGvcv4n8F+
SObPMHSU05LJQA9KURnvs7RN91+YTCDGjumjsPPhdJ9A4yHm5dVHs7DEGCvhHAj02MKTn/484iI+
P1LlMNkf3ksBHmLaKyKwEV7vOUKoO5ys8yqb46Q6H+KXiWDr8YtH0Tt2si1a+5Hc0Vy31qERGxiy
384oqRLHOyXCAjTMrNlll/cs96kUeuvJYXCzIk8e6seXiiTwOXbvaIbd0MEecEclbNpp8cmA3Xgp
xx654UMVyI7JtvQa/7q8hb8i1AvdfJlUav9DP/C8GZJRQopvUjB3jqcQMdsOVF9cmVs6J2HjXV1S
e44ORtZtbWlUWzK7hkBKpC2UdUqqzvvZzRWzoJIHSCJMxKKVYSiW+Qdr+KUsnGlKg3EwcI2UaYDG
P7tfl9waA6FYn0Ebhsb0HmNLhvdkLR00pGwIi1dpgXCHbiY57Rsde6b1/MVV/M8d5PDgyjsDD7Pg
ALbQQGkzz+RbExUPL1GSw58nAyHvYSWYBmPsSwzWpXeouxUPVdQq+5zTdTdu2Z6DMZM09TP8tYjF
G2+h7yQD1DGIYYSgWH06JO1oM4PtJOLLyfjmC436eJaOrE+dbmovlvBZkJKnbakcs8fOkZGbCXzM
m3tSNDyly38Vv2tv/E8+mVtEDouT/1F1egQ3h3aQD+99kwCDcZmTa5KDu3ArYKHINtOTqWMuNY3N
yv/6q90zJBgN76dUTDZpT1qKwFSITQeYr/4M+VfLtvAzQfR9+LpkZU6fKjrbQn8tWfk5ZXlrPfd+
C38GcXa0R0CRgs4uPEqQW+om0jMNuXpylhyCDZUvnHuo1qCcsbszoqOx1NOiGrGlAq8ko2f0hUix
aivHZXR50QDolgijRghTZS6SphYGYjpDxy1MKSrHdsssoIqMjUPmZ1On+fTIm+nSfUsM7neWMt4U
zsJ1pCzpyP7xF0N2ORLNGBhE8EyrbOnZQ2IAIxuRNKPXbJM5KmV7rda1BWDaTd5BzKk5u/16/5vU
CEAHOHWMTuFpD+I/oB/TBcjMasxLrjKp4bplmrtpML+EQBpAEn5lGJmHtZLvJ/Twwz9Y5g0lRucI
hGRIPsvpQJAL2c8Dop9ucPga/lxJAhogDF3J8Q6oWt19IQg2zSeEkJIVGtGGXsv6r2WJ3GbpAFPA
kROgiKzZQldXMlqVNecZtP+Yn46LI2HoYAhCxKpAf/U/616TJ+GEICPAkbH3aUFnrompaFgk1a0p
zqT1S8s4pvF6/xjNWRQ2X0TuwtfYZulR6s3qXMApIXalLR5GKRaCTdnAiUEohnLjrNpZMY0jbBwY
ZKK9k46Gfo5AKMBY339pVqugM/uWtjPkReQ9ToGO9NclfbBOsmjhV4x5wWLuBKw6snvfjDFqLJtY
JCQNeHxvFLOhqZ7XAAYCaLBxB/J/ZVv7QNnK4L50GUHqhnKfpg1ZnGw6CME1aOBDmUDna+gqvKtD
98w+XeANtP0tX0fNafB9ZSPOlFvIyeIj54lvEq7PGOin7RiRSG+wBDzb2gxyrC7gwswF2Ie2p3Sm
7odHOqHgUQG1vVn7404WTS0ZaIp0JvT3lqic0qFAHDd/KQI7EKbkYRE/ruCtcWHaewzQ8iXADeCq
47ZNSwigL3S7p8hHVxIJ5aUfRIiMyxtkVOrGkj0VfGeBIZGsuQAO2iSQIIHnS0p/TW1ALGz/aW4/
o8lMv6bkSXU+CtJljhF+UTPhcYdJYnldv7YemBXLrwXrEFSoAJRln6/w6f2wgVsPVsoLCxYdjjSS
XR73mhl50pMOhwYZxg0H6saexu8HqG3FQW0FK6LYiOB+SZEp7kcThzApmUtF8miwCHe/Gd+S0n8a
igy+ZPwD93n7XomJiY045z4QnhetGno/jIVllDRVvzxd+S2ylhs7g3sSQJWWKtnlTQFdUqQHloAi
78H3gn/seNCmEtlr63nLFx3+lLgLI6VG0JSVvIW0M11B6U/N4GD97jl3leZTGjID6Is67MO0q5/p
Nea+HUOWPBuJDzh9Zg4Bl1UoPzlFz3NX3iMtk3U433rp/0sOdrBHKPT8at8VYVE+YQcGfXNm7sX/
tQt6WP68NB6R2rngbZjn73thxc42DjegGdv+2sFbA7vfowkqmAUWyibdLhSwVvDaEXryxzm9x4wm
OHjVKn6S2kLJzqYfKf9bzOrYmEu9EVIzlsU1DokJvncFxRWl/R5yiLR4olTkLyJOGRXNqWwZhUvW
eUxWctvjgPfKsFsBYcqHIIVtOrDNi6KVIF7/KcqlT3SYZTUWLHwF2Kr6R0LjJTPS1lAhv5DqWT/Z
fiDbFYA2Qb9GNn6OW0hemR6amfwQTJRBze2RBKK/R2SBjXpaF4DvCqsn+xDplQzYsW5+6DLj0aru
Dhrk2ysWgPUtuWUWCAltobcUrCRtLjMskwPpMhj1sXqh2t3SiX663oq39zwUU4rew1MEMUye565d
E0jGib+IBoQ9DCOlhQE9MpfYm06zrWn+PcmPK1OHSY0D3AjVKN/BoQN/neVUbIgSM7OMZqjTU8tH
/hgx1qN3Y21X3Sd2uLETX1zU08qM/mefGaquNrCR9bB6QK+IoA4jq0ClNP3CYCxPUZd79ni2mO/d
iN1LhWHAIaSnQzo611xoeVacEDOWKECqHRGfsXJ9kLh/400Pc15GW6X2KaoKfV76xhWFK6vlqNVy
xbumXPb+0yf63iQuMoBK/XrZM369/mYIlDN//3OrTE/P4nVVcRZH866RaaWJIzCB1Yoyd8xdC926
94cnTv7BUP0C7Dt6ZVGwj4uRblKd3jRUPGWHp3PRxD0fvHTkGxkLpO53AezTpLNKGj0JQJ0FOdX/
45394coLBJCSjWE7X9VzuLMp3WQLh7dF+e1qwHDaAsFBJCiccMVXVnYAQqeQXT0OwGYBENvAx/P8
FqfSBQ/9M8/bknZq1SuzvitWcfUKtfWLw5b1NtRIU9SxtRlhbu8Uj4Vjg7oI0vm/UcB/gPVpx5A5
a2v6yNAd6KbDlngukjDoPHDMFbYgd3Ch2nb0p4WT7+HGiY4zeyNDwVnRTkwyX5d9NPIum7Gi+EV5
bZJrj7jJOn94ooO8nVhfwKWb1zivszXt1V4n9tqQDeaNhCe+dqIh55CuPLOo2JLkfpDBjcZF/rBX
dMw5FEXXFmkY5aPB5A3fZyi9DayvSxIDYMW7OGRFxdJfbWnWi3O2LFF9N1L0FivJeZjOSAHVntXb
9hO4JnjAXiZeJdt8j3eS0LwV8e7AKCtm2/lIrfEdfthQqUQ9ww9kEzxYfl3Fnm92094i5Vx0w6+w
vFCvcJeLwRbVOTS0DBb8hPfWy18hgcVqeOqQZ97UJJ/9IQkzO8Bhm2a9of7V5TDxkJ26Yox39t45
pu2fnf107wdUebmf6THPDbzHnLIV0NS6IRwN2gVzbqJ9V7BpH4MjjmyT0P+ujATV/dXzHxqMt2YW
kzag8jZLGeAixC71fTi6dEg8DXkkvqVQ8FprVFgoaf9a1qkf2OA86iaiZRGXszOCkF3u3Gy1TlkP
gdeF21yIiyCXbrek0UobGzVoF1NmsWhIkVrhFO4UgvBVHBfN/ug2AtmTCJRs0J/7I2ziDTpq+tge
017VaG4tKx4ZZ2f0kZPn2H752Wpo1eKY2TaYwk/tlDwx57tCk47cbX34KC4pBjAgOR8wE27OpYUx
dnxrZFYmtIdB9fO8x3WyB88lih5MMa5ImymAGZmq6CghO57ALuvViWdxO81uRyPyq7sbusKawsWg
POyck6a0zsbQfn4VRpquOMBC6rgkDamSgvR2a4RLjLvC2rDopm3e0ZkfsxAdVIfLv67cS9TC4/Ej
gQ7in4nk4zJQ3h9kXH9OdUYjavwMS55q4JaP4akTHXxcHUCNFc4BEHwbgpdtcQ9jYlEBfcL2LLdO
GKnRNk9gfoilJTqDe1tCrwF9ley0PPsPJl0bF+MXqN+fdLrIgq8PUeu5yI+BP/joDJ3Vey1h6lD3
NWgd0g8EF4mVkASnnLfvi20yn4Lca1ugBvI9sJtNX8CBj912r6XJECo3QfC2Q45Ag0VCl5Nl32JT
cS30Clr+JFYOSfPDdJ7ICPUiH7EhcI3ySyFQpzB/3Qo8RxyiQVc3YV+BYKvSd7BXhy7YelpUtcUe
d3lEiMCNcmySNJBIfET2c2/h1HsEFiW2/OiPFZ0Uc9gxT+Dtj9/Erz72PUrfO0jtdm+3Pi3PhyYn
cPJKeu3JRQaILnAGdlM1avBnJ3MM/eeMpnWFj/6tvOaWiZhrv5qvC+6UgZ7NiWYBHHCRMs4ZNi4b
6MIAwxQOe/evvhYrXoF+mHrhZCrC3DwlDgvDu2tjn/6JDydGrK/2Mc4Q4wJ9emEhDC/5d95augtS
OLO0Rf69huTfeEojvbkEM5GThcGma1uzryvzUxIUnFzvq0jz/8Gj+MD0/HdafiIHx3TJpW3p4ZcT
KPv5NeSVyyYwZDyTfpBh7bdEU/2p8qsQY6F5aAGlNCa2l+lDFORZ+s200seTeLQTnN7Gif3Ytb+6
r7+3Q0qMOGMR9hKgU3E5GlZ62ldyb4/ph8YLElpA3ISF/U16GH9w61G3OjXYSmfb/O2uZA70cHX0
a3rThQqvmakopRKtXk24e2ETSeqDhPmSydtxoEJpcRyX6RVl74mSDvtYHbe4D0Uyuham9Turvd3m
Yfu9k/PqkvHvDPuHBf7V0/0x/bjg6YavKc4r6Anv6uT9HryIk/qOE2p25vEkTxaYzptqculn6PK1
7S13kte2E3JqU4JBQodGJ3sPjuBoCvtXnqdMnhJdRmE9fnfN3cpvS8786Ofo9m7p78811fI8XbtY
N+P/EdTnWbNI/2mAI/QOAe16iLaf5NIcrsCrU9RWG+gkNQj2W8uutpSOQeseHvDexs1cgem55iPc
Ts0r9agmLvIHPkm8BUADCMXj/lDU30F4EQWD/U5l7iSAtktqBfhpgj4dU6iIJB4KyoUo0+/+lyhk
DXzKnl+58O9J2OrRdXFYPv5/bntcj/bY0Md7vGzLcjMX60iF0CN/ke81XQPyAK51fQ6uK5X9OnsZ
b2mV1ZusxRrJa1+piUjNT+9ugJjvfo5nkBa8T5E9nHhYiAOqU40heUH4KD8GslvBym2Odd2NJpX+
dvL9AxmcK2hLZSNN+90st/BB4O7EHQwvOw6eIVa9v+D6Lmt7HxOWQiG7AWm7GmcThn357YkoyXNn
8Me5YM9OOZDulxhlvmP815th2cQAxgsSmvoWW1YrEbU4lwK4IoS/Ye1zTY6U8WukBAM7wIAinS+b
yKKX100bzOlC1y04PU850mKHkvJ+Gm6qE0nbh6ubUvTMriIBTKPm1kFa0Mzk0hzDKZ2uKxlLVJd4
XsaQCbOFmWdbzPb379Urb1S5qTmXvQIc0u1RdglqyBnge7GU6tHjaL7kD2kUusDvSdvqdyWSHArH
AMqjoQ+hb+IECwe/MBFvJYPIQq089O8JaMle5cqTKgp7lIcJT1lYmFrNsuQbQcfZ70bmczKivRhq
RLg6diBGTFUCClYyp/aUJ5VLEFzvzdHgLLKHb4d99c92O9kCzY1zcr26B4htfkV/9n5orJH0yWub
jI7vcxNj9p/2zOa43pJW/H5gTvxSLK6ye7SniPLSnzqx/tx2aZkQbYblZEIJlIdZkpMlQKEnfCpD
spuVDXefoMe7iiqpv4f2g0YAZdCtWEYu4gBzP1a0sXiRyVYBoOpB7h4fHMcnSk+wbw0R0vbWayUn
B/kWF3H9MeoTcxd1tTIyjraG5PNlip8DCA3jYdvB0dKcQOwt/pIH7Pz6NqH4U5u0EcjWv7fvFbEg
jKRSSECagCh+pkXvpGjT3lMTVgPojNOyXCLwQykfXRaQX3K59J8g6fY0gZgXB2NUU9iJrzQn4DJ9
yQD4xVGzfLCqm317uU1HWZot+NcSSpxvvx4mq45JBm6m9SuKtCR3MjIt+SO9dNY4q636veWjvuta
jaj8rEHq2qQVtdS7uDp9wHC4cmLRYEShHhJ21vNZGAlAyo7l3+Kt6LrD7QycQAdtt9a5ktVVRXRO
3R6k2kZH9DIKAmksrIYGU7TXDDjdBTzPcnWVMQJydLEnKitkVSsyt8vMEfbV4dS8YIStA3YGfUJ1
Cuaqwby0kjD9cpNJu6liJg7wrhLIh1EsXF3t6RoeA5uePwtWz9TyZc0KioKO7qOUmmS5uiyRL1qM
/C8QGo8FnTzrven8ENPLLKkP3a+XYfKr+y/fPjn8jD90L8gvQJLW2aOAzBzVEd891iLeEuJv2iE8
GyXb6ezhKzLwKQVV2j3Qmgk3u66DVUXSmXWWpoVQE7TYDO/sHtG1C3dqK9BSnfQ5yVnS9TGB86KJ
REv3TOlhqrDGGlwTGrJ2d5Bm72d7kiiPqYmmrzISFpX7XfQA6hcxqYjCHWxM8rUkDLu7T6KtWmkI
V10rJoUelcahp8HUk0FARZy9VOZUkupwPD8VOGIo6Ede1pg0tT/T6CtO6OGl1bh2EeTs9L78zfdW
lw/EN2+Gkp3iXUWvyZY94Zyj4pKyiJxpIpyMTZI7CVijU30P4fYSDgBc4/JLzBy0AjuNZsguKB9A
CguN+s2uYbvfS2VsqGl5AEtj3u9F1lSMMsWHJGUEeTY2BeoBd8c4LgmSD6EpW2revllAXEt59hd2
N/rCUX2vWv9fZNbunTdgVuSXCy1IP8cEoTBtQ8vgaA8OpVbtHgYxsqV0B/UyLA2gLSsivOyfJvbW
ZJm4lM/YDAfIWTae4Hj5xVD50R0TvcS0iVBxX8mEP1iMBMM0lJhJl0dbxlfZLtJuDBevM5gKuxtk
Pe88f/uRgj8MMSTIiNkwLzrQY7S4hbGyhG4tkHqM5SWIP8Fi3bY5J2vR5ekJLwmIh9/bIBJMqpCr
N4n/7bRqU0aoR2XE4qulBlf26iK/Wed+IOmWSDLuMuzFbYcPwgtm6Ar5IIQvBXrKCmL/a78ymhER
dw2l2nDvvjm2lQWKCXsK+LRlGbitNJk+dIimwMRUG9HVycxxl5XbjJ5gpIee05O9bgJMfpWa+1+Y
49ni0PTdj3TKHfyUbAnp9FBVBRa0tOEgL70Ik6Dl0lnFelDL46CdfU9psIp+OwzcnbYQHuos1eL3
2JZXVqhhOhTq253OR4eMiYRiG74msGxMaopTeMHv6WpGnkmh0si/UwkZmWJ/elrxwE3X2tKAmxhn
fGHfgq3O/5bYoUURgmdHLvPUWYXkrJEsLUVniTLYCW2UuRPJ8tOVspgv5hdeYsOuD6EvX0VEg/nE
oMZsiqsd8Y1k6UenWGh6bl0W3uk080fk1Snq5wY2QCY084t1i1V+Wmb8OK7sFW3f001AqwIhm050
lB4zrwKY3nDzzcAOEx+hQBSWXqc35ZZSjGDkkhMRZLzcoVifYKCLKPSgbDIb+H/zbhxAFYNzSG6t
RP4Bmza5dMoC/yMSlz3CZwhOzHi9uJIairnxrbxLNa+jox7PPTtUbhYZK1HWNYdTLQA/egBt7KXH
qX5nyeibbypQ1G+urPmdm8r1vvsbPujAM5n8U1QkYDtd5AwbyIi/kbiW/cAf93v7M9s3OFoEVOeu
GCpg2FkIgkuG4Zl1vodJ3PwU8BYeVoZPbpqnoOqQ1+GSeD2LMH3zDUF1TAS4suwXsvcjsJnmcW3b
R63dLVHPJvUJt8JLVsyBNb0m5oGsNlxAZlrKfsapVllq67doyCF1URLnxjK0TG01aLB98KM+oBGT
bIyBa7OQf90FlJgz4TmTaO1C3FuA8K8sMrzSlxP73kbwY+S19m2c1KarCRRemFs7bUge7qh2XY5M
BFkPvXs4kP+6Sm5loCBEcrstfCcTxuJ7PaEPszir2rKmEm6ZgGK2GsNul37GVyb1yu3+iom430Kc
Dvan0LxZFP2RXm2xZAsWrdc3on5npRCXqcGY+QasYJPfgTdd/DOVCRAvIY4Q74zQYaZyW2igW/le
98AwPB9PeCoJAOCaCCADut8pZyI1+BHqiH9GaI4xpnYlD2x74ga96XkvAXF3yr+IduTbcadIctDZ
lCfg21hZNf2ESGyaR817yYaMGniW7kOeAg1IpttkTh8BhkP6kthl3//tk5LNIkljNW3vCraI+MhV
yMClNeK9rBcyRFsAGM499wZ5ub3cqotuXsk+ID2yYFfsECX3WJivSIlS2QuPNTEs912Bb7O60x6R
uzl9ZBGjDn7UtZRZlNLzye5+xjsfVEB46ktQFMIFgip2BYgalilSFpm1R0f4FEoR9vOudYgH6osn
+KBYKtr1h5nVQspcz3k4E2VqvGIKhP3V/IHPHd44sv5lmJ7LYXBOBKjrkNuvUr/czsbramcGRO0B
t/ptI8VVJumsAEsolyB5T3zHVnLLS3m82AAKJJAnNr361I5+oJ5wMx30EaXzR0Bd7/aNs222+U8v
YBe0i99aW/Z7DhYKSkV1x7H7a0Si8lsXD8MRL+R12sZnZBp0Eyy+B+li1528ehjC3lWgXZO1kjKA
f27AfyrMpUXrAubT1jk7Ex/HFholeZ/m+IAsPtigRuEACd0WcqaZ61GsjyOinjYu+uyqYXqxyQQA
V9qn3iYDL4k2+0y1pZmP7UmnUvsZQxg+LQZz/TH75E+4AS1szHJ3cwbSEIwHjAnOeCahkplmtE0O
dvfMtba8p/CbYBkcL1MXDqHGjlbgEs6C07IXmkKoE+WNOtmNGLTc3TfjEjzJ68jbJM5xQejlvkr0
KB3f/4QtZMBxCRStHY58HSHfarQl2HBqTQ84YkaigDmLNZNu5sDXlMrEw3HMjvrxe0fHsRSlgIgF
ReqxoUhBAzQXsZpVdMfdowLjw68Fx6wtZ62cyzD0VvMNm94SEU1tQWQIKIFuht9vAAu3Egq6mNtB
yhGe7qj8gE5d78bWEqUSxGgQexTGzpL3/H9qiVmcoj4AW4mXAtyLmH2yklovUcUQsnlGTgnPqifY
zxslFS97iFFXw7HSODUYMaw09iur4+JayeUczGgLDL8RUmyf/SQ7YWEk1v6hzxiil+wkQUxkNBOM
g0cB4k7kg8KdDQjAbC60oiiwocvPq+sWIIBPYDcjH3mpJ+7xxYIF4IacFOT4/+KMGlVB18DXl2Bo
cSjDdeigF7aWsHMU0hf94Bz6++XXS9d2fMPonufOqi3Chbi022d+BH/wswvJTz75zDxflsj6gxLJ
aJhJUCBYMB8IOI0f7JI+YjAEEtwAZWEYv69B6qfWPY5kz5bPYppKKlLQ3pDk10tJ5NBqgQxSxU+8
B9qxR+YwYWa3d0OMJeJYG41SOvDhZ/Gxk7ArAofHICebHpdRIO1Id7oAkKbrfare9qHz4tW7xyr7
OWIWJDmmdDwlZ1AKByLehA19Yup+OoLcAjs/Dmr5kZjD0qqb2A3BSC8lHWJ0+tkS466FqHvA9Wqt
xk8yfoHRmegxcpbPjdcxHV8dji6l6cQ1H9ZwJ1lvMccDOHPftJWmYEH4VmPVemiZE/a5VWEH7COe
82VEKQ6n4QMxGmhMRSOFXhiA+hQwN/LurGuWi2GCFPWnXegxvn5blp3Nb0mLbN/AzPwvn5eePTVb
au/LwKqYaSC6zzTqHTOUo75tJLb6qhsfFdeydoyIW1KzrkvVmy8UClVOEb/xC9HNdsW2Jsz7dP4S
DZFEnJ6OxtYD6b5ATI0fqtnUBQtQZvIKyx5xJ7dinX6v9YF0pTIB876+myLOvfK6SOIme4yZeHA8
06tIvHpLdCYvOBRlDWDtR2FWP3+F87k+D0TMj1KwWRWxY4Lp62nLaEJcPlPa4fKVkft4umdEhxj7
qDkojOTfk0teSr/xkAZxwy1u5vreYo18pfaYd/9EH/TOMCmzpLlZtFcyMWc3NpKsilV1iQO3cJpz
jv6Z46IWsmeByucsJ3l8zfrRaP9LF7srqP9kAKUa6u5koSCaRQGm38tmqBXmKY5irreEjbgxl3HH
Z/uGh0Nesr7BvIs8XHT5QMi++IFFZ/6lPl+H1EvLAtXz3xyBJALtkaVBi6WjdoNmLiHtWphYrmyv
RUAy3Eq1nTS0UllKvQcGOAgfLtUNK1yd9zLSlgI6bBv1CJfUQDZ/GMQ5PKJo6r1PIQRxmL0k3PQx
wIv4dB9ue1xd2f23irXpIoJdwKua93zFOX9RtmQ1JWLOpsjL/tOOZoaNHy8loVtIfYQObRrKAdAk
oERW5fHiozCdVWt1PkKH9uVIi/zN22F13TwIdoTKpii1VCA7QcSC21Oted4q+Z14w3B2CohIosXV
g9jR4LgG5a42HTNWvBmia29ws/4xCrkV6kCoLArmQyvCtfDzs5T4Gfi4l4mgG5N4ZdqE3NrtsoUd
DkWdM/jBMO7q1s2OZWvwQbKDthU39OtqlcoCnBbHenH3P8dZByiBOiiamuYSGlAJgCdcfgXbqGQ/
zeVXJR7oQlaDKXzpI9POa+dD1QSAy5YDCMMPqdqoC+fJjut1yXlWUU9TVGc+MCsAge+zZgnN++fG
Yq1R4CBv/L0jRxhxtrgG9wsTa7w72yZZvQ8ZfurFXOnNGQ3Q84d6F5lJbjHAj/vFjlzVauv560RG
ZWUOuW7staebNbZVPCT5H+aRGrZ2KHjqdUnHjqSGkghmpB307zbFidn49k6Y3yZppurcam51GE67
I3X708DeB5VeMgRMEy/My+hKN7dTRNU7jr7QINsaxDAOq+GOfEqqL5mXLuCFQPNjAz5vdC9tmnYi
THvreCzfm5oA9O+SNr/iMtEIDLNVYgX5vnxq9dToiyZ0wrrqFmavVx1VWK7xFwFK0qcF6U4pl9i4
69+7Gdon7tkBbwkSeOB/rZ+i6MRhx+ywvnfJ/X4TNUkw6MTXqfMjyrLxwCbPB+LsNddqMaM6wnCd
HTwjWk1Q0+PsZ0OJ+ekJsKci83/vOkoQdjVZHgsgvnh6V23ZUU+lUDC1WDSlqjMIVfYsQCqFNpNG
pS5bj6r0cqieiBuzOsVp7Ok7p6/DrYNJm6zfsfc7dcAQtT0i4G3zm3b8VwMWQbaq6dPfzD9sAzf5
3M0IVKlgiuUcK82bKyiQXBFFKiJ/8CbLj3FlNVqPedCdfz5yjCW2xJcPAUdArNlawXK1wMhYUrq0
HzR+HlnFse+qmzyPqPma0Nb420lqRsaRZ+HHWAfIvuOeguJqNtMpcH5EAmFDNYDwrGCtMfttIarx
x1buzF69uKsXVdOwlbo+ABg30pEsZEdF8jOoL1j7KeOkNNFp4fhuo+RT9VCaYpJIA0qdorbUvq4n
vroT9bpgZsTKS+otnr06mUpr2AsAAisbtIsh3+RItYSevZgEPdNevQPypcvxTmoJkwl0XNVM9fPr
4D/MurDGzeURZQlu4sWjk1uoubPjQEfy0nYPsiGc4YEy09yH0UUikNj8PNQMycZcef75Ji1KOjLg
+eg28J21siQn3ZL5QxB63qCOpMJv/wM8bQQgEYiXTWCQTR6odE6zsqoYwnMoKMYDJzzYXuBAQbLV
qtizPj2W4mF0c9j/wcn9WKtcjNclefgaLh1v2YkNAkoCiPvXhtx/R39sxB06wa44VcvTKaNOe16T
IZ23eLXT28HBIonMxfoZaxm/M1NEpGwYYNWxIA5W2eeuVPEGYEDWyx46ZYmsk02OT2z7hZK4YdaX
7jDlOfZBIS/N/VhoYTlGrH7uDoRwhv+4tNwIb/CeJBRtflMWoUhptxEhgYBwtCZMXOhzd0NwA5yk
wjhci+zEAO6870XRXn9cxVnTTGPF527MzAhLdM3vmvbE69ZtU8aehK3wLX0LuB5jAUh+IPQcy+WG
Za7vgPsLXpP3xoBGcohrySUkTy3JB3nqTtuCQKP6nUm+h7aC8PKn2WCJLEGrygoCsEKwgKM2SGvm
VkIOi0XVpENoiWe7V6cvVK86SI6YjTi+8ckxtQARsbyb4KdFPIZknjwdXcSRSev80t0sNmM0RdyR
n1EtIEcPDMvYnO36eIjwfccAip7aU8bJLVpZgGmzETzFsd0qCvrWqYTUTf3i4WqPsQiX+Sw/7Hxu
/vHCDrI6lbRfLak7pmeFX9TJRW2enH73K4EqkkiIwxF8I2NkUPIBox+z4/8tfVtN11ziILkUgzJd
F0ruMAl5many8FvPWvonAL7CF0CVcDsojI53PytWMwnqhu4zPs/TgXVNByHhFxcuatAvUoiQw9Se
Lvfn1B0MZiPSh2zPgFwjcFJOcwo0Y850sygXTccWH1x5HFd6ms7ZRdVzrsM7uXk8xnmxB8oubn9e
yHGuvyAfvyyXmWXBMDmkY4RKBvz8goo3JQ8QDw6J7Qw608Y8+4NZ+lnrnXy0l179zeJRQ3YDOT96
nPR9GqjBUd004ks/2Bg3beIHS8ZxAg1lfS7UOePG8CuxjXPRVBs/+Hb5Iict7p75V+N3kAOUB2g8
kVUgx16MVVfRBoz/ISniQi1uo0gpqhBQ3F3u0yXQ5VqmboDsKKVcdwSvAWK10J+jrM6MgUTsGYZb
oSJ7/mJVhfGFxc5gYP+fJvcUhoxbU2T/lg7c/cdZIyv7/6lSPeb859T2XkdM5d6YqAc18tCX8lMp
xovZGDQrC8ox3nuAdu90SU0DdxSF5QFkW0sbWwHreIg5uBDqFTcd7q44iHmPVDlVHTfp7ZWV2fGi
GyueWJ7u9yWwuc1i0KJePURvvwbUVNuQih5zal9NtjRNOV69LQg3FOxX3HHh/h9Et9iVx0S/wggh
5N5L6I1njNjc+9q4Fr1mKV/TZV4wJg/96XNv4O4lS++HRXMve7Erpu2H3wSqUBCLvBEl4QnUC99f
2HXg5SUorhwmQbsd3kOefYGmnKIryN64K8pym98bQ9xxVCVidSMIBdQTPw5hbT+qlPdJdtcl+Nd+
+sFEqkQHV45zHfudKjl3ke1pOBwFu1uQPevutD/lHaqC8Q5min8VGjBzkjBaMiuVMb/QHdp4Xah3
5HhWvN7eQQJIMnupdumq2GDwHK/b7HusJyvreZHvxL2Q/2R98YEMeOPr428IHv0l+uBCOZbp9Co9
85oN51expMdoouQfP1RLJMx6EQEKXFgyyNJk2ZmRmUe9pbcwGEEPZJ5PWpjoa3SQUo8eYsYqpVK6
tUfwDX9CgtR+RTQpL0LxXEDgNmRXi5NXAMtdCVp5QVOhTB3EdPBp4U/QMQQmacOeuW7K65SDK7za
5HC54vyXNhRXHt+59cJ+KhuQfBO7a/MTkQvEj7WZmSsoR3N8bjNC1Wfle3Sj0XIt6jH7ofsz2HaI
7ahUL4uITDRvuC3aMTLjCl+W8+PE9rPDxy2NW42CqNewpC1ISACxBhpQsPTDcDGWuGf0dkzFRBBe
sytol6OaEI+O4BE+Koxn2h8TbGhDEAGCS5nt3Pp42OVZkCeJWHJPFPNHgDnJ8y4+QT7GzQlXsR7N
Bz6OF/C0VfoDtRDu4MQqwGnJg5xo4AxtGbDl4TVsdVzJDiqDs8LQcNcuEhapEzjlWpkHZN+ngqYf
H8Li34PAGeJNBXb+YFDbLAgotO5SEDQX4fUywNJDf9oW6Y0JsnsdbbVv7uzNo+QE1xCfhh/Au5wG
IKiXT01eWKy6IDxMypd9Wl5LkD7E5ylVeT+VCOlDvR3TFv8J5qeAGv8WucZfwxBWCBoTXscCkxap
nKF6RYQEk/XXo1UPYiIVSA6y07CiMgwjkZcf+ih9fYZDPk+VR9g2lVUUZHAxBHTlJxYBZlyYIefu
JNYkL9EFHNcPHjoC9sPVx5+idm3yoUfn1dib07ggO/sy/Ur7APZSrxdYoYabeHOAX8ghefYu79ol
jfoS2q8d6SLxPVQCWq/uIB8yXpW/2xhy41wr2Ru5KrAouKmd3Oq/gmLYTleJD1egQYSGr7zpRJ/i
LTneqpbIM/gmL3dqboY7seqIxHk0dus5uSmaZykUCAlftKMpZZ9588LJxX3ZyOR3LJvniiSEGqvd
iLQe/66l7MA+kwZumPw1CTV5q4kznBxHHWsCtBaCsCk+hNGiZw35k9BWIddMFucrfF78gIIW2n/U
PBauRId0RIVF3KovP99AlECOagELj5t0lxWEd8MJlS1I9H/cz71IK7Oglk+T22XmSe+w1B+XT+gJ
AOqjJHhWVLOwu0ddgY30GSYC2v4gJo201iEQmwh93akovR2T0QeXQOWkukuMgbGiDRK5wjW2tqAK
15la1bJkSFAgSSAfB3cipYLBa678rry+70lEU4Kk2HdWwXDa6AI6WdQehg+k5VsVSwtbGFo/K9lU
mW6pwUri7GwTUb5o5DVtteycff04JexJ/7PHcMO2Yp2iNKOTEoo1NOUTxnXMGk/XDy22t6qx5LgH
eZymuMhOYdee9rrP+UqsA+7FKy4L30PkQcG5KJPlAptvh/qE/aqisCPR7BR7cTBRGSkYPmAstqXl
ai0CI9kP2M3fzzVD78TdYQA0hEUhW1fTQfhGg3BCNV/RBcMSN8ahDBVMok/uwM2aaKNpIsa+QF90
AWmGhu70FLte4evJo4+zUg4AJ8qy8h5XLcf4WIvTovU8sttKY2CTCFLC2AN61YFd9F/eBryTF+aM
6XfvWioN1c596drid2BJfB6tb0+DaCjX8gE5F81SWiXh6FZqoWRCCzNCX/n/PWjEwOMZMJ8dkWq0
4/Cf1eKEJ2H/yg04ETCws+vBdf30xnWgU36poorlMwZswms+Y6X1jbRQN+mxF+rHK8lDnStsQck9
NYbXSSlvz/47sKrWo4MvQG4suSZNYEfIT12r0tszmJMDETRp94ou5QIdAHJ6bkyeObfbGlFa6cLN
pKGoywcO5H4mI2MY4Oi0j42//OcHL7aGrzpXrKa+LJ3C47wzU8S7JrBcIcRMFF++rLSTDum05nPj
rXl9Eiot47Wz8cgjQ+sFwjhmv3ycbJajEnjOIO0noGSVbGfRV9ncXVObLvfjGoAPYgJgWl6YX5kI
sn7IwrnlX5ieWNhh4BKCOu8+AUeZt0MlLL0wRDqEJBQMRSeV9YHDDtfGtb15FwRbyDImPbYUTgf+
jfz9UnISlOs8j+aI11gq6L1dFaZZq4wrx+oUfFQ7AVUnhjsCGoih6Cf4S3gNr7CjeJT79M7ka34Z
H0hGaykvZQ1rO2A8cK8GuITr43rs7zfq7W4RqA9EynBrVu0OS1y+avwdy3SfCnilSrUqeWqDGFu+
hZ064HhT/NCejv60G89sw634iSy67mPQCJcUFLNICaIwQ6C1+bJ5ECjFMHS7tg4nLmU67NwS6bbU
jteHoRtf6liDuk9pD0vcsfHeujnyde4lykfkk1+1mp6sneAE10txPlz7guSA4Odz9QRBL3u9Xh3L
han9i7qpfxLAOdgQx7pysOTCgubozbrla1QK+vq1LmST516SX5bxuD6M6kqljxyRDfjR+MBq0oJn
WhkQVuphDj2UNzl/MXdb+0xKQWw1HQr/KZeHQJYS/lost7N6cttejI/Wlw8G5KC0uJOQn5+KNdIB
wrFDub8S9c1kAAW0SawQ4OmqW92KsJRtV69e57JGDWbifWnEbujUUSjexCXgDpra0kqb7QmTrxfV
flV5aARjT1zg5Cx/u6MDJtkZmmLKxOQv/Lcg5ZB0OVetnetBQ8rGF5cph7C8YyTZYZl7MFaK6Nbl
jEziCKHYFXeHjI5u5tDBGDdyhz9Qp/RNgOhD9No9VVCPLmkDVgAOS8xKd7Y7C7SLAAIoXIPE+b5c
++zXPmvVqr//NisR+GYvtq/pNjVCWv2szUPlo1H4/fxF5gNx1U15GheLzGcTyQcwQnfS5EGBrv7E
huX5i50NthoHG6Ec3kJFCWGMr6+s83ndB5HHcjH8SBbLqZ6c2QVt0HizDoQFjeblSSzD2m/NC57o
88kK9eeh14YSNcsor4TGRQi//XZd5ATa0Lw0ulyi+b4IFseX60KKGNd6yFhCPKJoPSN8KQoEEQB1
gMxDQ+GTG7P20fEtR+wt+EE8qKGpF59crBw+EwJ+izEA4crfEr16obVMd3bKni1JORrliLl+Y1uh
nLP5iEE+G0n5868DMq2vHYszsm4vexHstDwpyROZkoznBsf1LXRTDrRZVKc9LP9DAmS+ttcCPnhf
LCQeqlD23NbqXORGSCv5PMjT4678irA5kOSZqiinRgFbJOd5hYuwELmYTgXTtNWYIUOTpwF1yQv7
foesSl01hWY1EFAbaSZjAajxZ8ZvtoSsSEN6hUIby+kYpSc0FL8sWoBhX2ftnjK0g0cVvTlJesnv
SGiIzvv1jMKcaUXMsK7hluCOuzzGRo78T1elYhxXR8Uj6OIGkaAd91VqcAUZRh5A0zQYqMlq71fj
NIfJe5OgJNHDR7hDub3a4gBSFUgmC1Jk+3xnQLWUHn/YrOyKfx4ArVu4HTp3VRBX1nq/QQl/uOAu
dKdeKQS8Od+iBRxSVRDODhK4DUopbCbbxUy7Byjif/zszgAJB1KUOqqRkBWDCyy9FUn5o/mLlZYE
wO0vIXEJ6ZrIJHNW7XhCE0yp0wImPbk531tvVybhoHEeR1PlQzuegtvYH2bmaYUS6zuiAwmXJEVe
neCZ9CkBkMcVfmzX2YaepMq+MDCGeXwoBvaQpKlulk0SJr/b1tFYRbZrBzJ6cD7jz1SgtqRI1tfp
IJSlyTH+k2r3La7AHWHtAObPozWS6owfVo4zoyScBwL67OWeUMWHj8suPCRqvL6pX4Y4gEOiofiC
s2DkWmHodeZ99oQMobbWlJHUl1w1rFGjXVpxqmhIVaOSXAHaxlsTPdtfi2QJmxSOrxEmPe1e897F
m7uKcl2e9HpXyVzxFSQPfgVxOkINU8z853QwjqBNHas5c9Q136C1Fv47EkNrOwvoGU2dh0JqovXR
OnvyUwm+RfLqaVuPYX65yXLNYk/vaFvUqVotVlXz4SCM88e6K2INxipaqfds6nGHhtLk038E0jp8
ow+xFV4SHPTBrYlLjQNCVjZHOxyAPcNqFtxH3uELtSIYBNTcKJnsC95dqfJX/qfvyZKh/31klbfK
yrJinxS57tGHkkNa9uvunXFMbvJ3AkWi+lAYhGhpZ0FKFof2GtXWDxop9eBhQN7DXwWS77wu9X9c
9r+xJWz4w39ms/PU+H37AzlocYujPklDQ+K5HhcMHeSJ8p9s9BiJW7NZMZW40FiyPF5MQzZS6CQj
pIz0GlMfHudlbt4jn36B3f68aqnSoU/IWKOEzvr0HvLZCncgFzh+VsWWxJoVMXCU1mtJtE1562zM
F8elWc6am2UaRJQK6npsXbswu0pLRjXDdzf9+rRQ71dZN2eFbEEFor5VKvwG0qjIIW8rFk1vA4fd
CEdThmMAhEv1eDPagch/qyVLQaJq4b8y0ckatFWPWkWQHoO9v8XkDl6ZrGt7PWIrwlSdJnjrOnJV
gkF+6Vqyld0otsT+BlLwtcwlhKmvrQiarno2ArFfmGr0MG6ruJtPilYjkTGmh7U2RChS+d6JIL5d
xN0q752FoCxcB9zhmP335GSOMY6vSVhqBKkCdfAs5BSH+LHc77MfOr/ephgu0SQPS48icbMnJFaC
Ax7f6ompIstutEjMRzmiawS7XkWzythUxbhZ7zCDXqPC02LKvStCIsH29DNbZtGqxjdWFa1SYBr4
I1QJT7hFVqVtfDzdDMYjYLmR9UkPTowWJHAwC4FI3G6WYzKHrKkQOhEFdukNk4vHY5XRq8xtKTmc
kIE76egBkzo7RocpSZAu0GLwJuqV4cTgqZOma7Ih38lXOBKFbt32R87YNrJYVRrfv6fAv/7UwIjF
91+uVrI6CIENiKId9XMN+BGOzJQXFcOjWHZKiUmBBbN0kxdLcyRvc7KanIbggKPubAoUIIouRa2l
0r8bYAy+oaCogzyqvlFnntXmVIJ1ItzuI0gH3c3AfhtFrBfgrrYjKIjxUNw5CFXt+Z7NPoTFuYnn
BwX+jcR5bta8JoFrPYZTL6sd91Md0flMQ9DJlPG9W7Jqu43RLWLmfHt6pkBp3p32WUvky7mt5nvE
qtFSxCD8tB8tuWq1DkZ0cDJFLhY21wRkrJAMH+hHiTAK53qn5ApgmyGCasAL7WU3UG1dYEAwvsfe
RjT9bBuN1zdBn+UvKr2Z1uyYHJJnIZMBEMw2Z7Fe+ibObSQDgR6yGH/APPTQhLheDz12U0G4siPk
O6/gAfKMNGF2a9zcB9emW9DszHn2qc5bkKc1HakuHgtL11bvRTau84IcziHDHbPKM5m0HTk9BmXY
2gQsSWoB4SLWrIfOJHAVw0ClRY8xV0vV/SuJ1m6vS3ZftJ4iW+Dy90jAL92VYuObRrKlop+NdB9J
e9W6buXjKwOm90l+RF3lwTqsq+Fa56FJfOKSEdIXWM9Tk50Mn2nv/lJiV/fG29Hj/jJHSYMOOD6K
oj+RatY39m6+aQ1UkRqeeEoPnQbeQ0aWxqQU0IghQXW0eaupd5Il+Uf8GDqmlZk+lQgAsZUEvCIP
0D9c9bwyClQk1sBaiRpuiuqaWuWGNzKRUgzrH+6DuvMaK9JSj8osnLkQvW83BDhuuzdBLtVJRrVY
rnM2qm2HoIWo1HhUVfbYx2M2nLuK/mTfOyWaEdJS1wXPJ86zU8Zr5C4WT0fb7vUipd1T6EAlxRnO
gORQJhye99jUd3soMYU7/eDv9ONFimpwE4RErA5abJXEhITOuLC9Iek7ulaKOcxWvpAmJfdvAroN
n+2LyM3Ak0oLgLS+5pgGxzVoSbhyMRYR
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dvURQc4jzK8jMGJp+AY7Vi6TjLNUg5b+iMcQCDcQ1MwjAMXQcFJ1QB7UY021mulnnU3itV0UNO5D
DZma+9TJGs8fFJg/0I5oKcGEqWclUPwoq3PHWM4UpQgGm/GO8w/0F5bgwCG+FJwHlAX+0kn8Nz4z
fpXia9yCR0ETAfTTg0hD4ypbtrrgp4eggLp+7ZQ1IWmpkeG8LC9HO5v4XxpZ5P7rJcW1+OHrdpWJ
ZS9uV87TG14d8tBbU84mkIgnPr8s+7slNFWlL+9+1t2uKKQz+zE5Jp7KRNjGO7BqdebwQqlkxLMY
T5Ts5lFg1wslO3XI8PtP97mPBRI2EXAwieJ2uA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
rFAUyu8Tmq3LPPCM+80qKjUZTL7kyHc8CfUas/+8+qukbDFwkx3pillkDQBA26Bc+TmaNUTLLoUs
pzcg2Qbyd8a/mC3919EaHtdACyaNsYJdqqV/e9yBOErWZOWzgMSMkUdQvlQkdFQ+uMPwptPZYZFk
aWSpfGcnjxEFw/tmAuaJzgG4SoZCshsj7v0plRmBNy8cBAc7mS4zdRgVyzr5VDUUTiE4Ef4phYuf
9my93EsDOPY9/vVGJvebZFMXSGA5U6EJmOYa+qpNNTDTLF9E5KWaKa11s/MYuDO5SuKvszqDpwm9
e2VlKCUGcfWShjeGFHhpysTe+lL9sFqGtTN4cwUDhBWfT0kGVAeugLADLvl5L3tTOBS+IScL+fMm
GVLbCVJOSt/3lBOrZz22rJq3m81icIdcrX4bz03aE/eHekAcwtajJhKNgRurq++klwIIvko6T+t+
/CDHmBQ+2j/IiXf0Lw+Rf9KAcssR6K7h4eVUnV2exfrn5/ME9IeX8K1QovHVSULEVf4YmumAqjXB
0mUTqlX1RZVO8fJ264j+kAj6NQ0NdJLyWvXPhf2v82DeQ2NZ/5o+0UWj0rRuZa9NssGZFf2rp8Kl
+gPf5ZXLqzovZdnf5UZdcItfoXH8ag+aptBtZbyz5jE9vg9jR6VplmcLhSLRYBTWv8q/GQgoDoIF
QpUUOVXCifVf+ij7sMhzopHPIEj/uIAmgmqQGLnMPkUsNak6Fhcl1i2xxP1tqOS+BAMSSZ/DhjFr
wbLVeJ3Q4/grF7w79LJfcNeO8uO4FIXDmpnqOGWKiQq8PdSlyz5GnjL280hQbxQ8S8Uee+UfUO5b
QirS20V6Ew6xS39UquZ3dyMtP7d3XXhLJx5u0dx+bfOXZIwYOfYEn/gC0PDM3QIb+Su5Scbc/2lZ
vkqIspWR4ufZVCmEeFU0PPvToNpKqz9yWybPUvqA16zoIh3wZbUdOs6/sVwuthiTaYZrnqii3h2G
0o2WxcjxDBmyCGFHmPuIvObzpyCHmrWq3fPaMaCbydL9NAy+TA0rls06UcFgiJTavWmDQnUqqGba
M03R+sfXpMNxQMfMRoBeALPw+jr+g/ui71utZBzm4JUvwWT+nFTYvoJx/HH1qoJjTBVLUUSx9hgm
IBSlTu5ZY86KYdLIM50tHIihbFGtH4icy0/6r5d0I8SaidqdM+3nYfLULQ5+PGAHoBrRCN9nqx0g
zI7cOtByMOlPagR0CuoqjGh7Iwo9aKFnxdL21mmqqnFFeDuIfE4rl8Y7IWVgD1un1Rj3qFhzVtud
RGWDQZBZXEmSm9NfhxA7WddVqFasi8SqiA/wOO2nOm11c4zPUtNeGNk6MyZuGIrJzt8/Hhqtt2f3
1VDbhRKlk3Yb6J/tV1ljNVD0bMFcuwVjMaIA0KAb/8vHm0BZLYbyPAcz0/oRvgtY8U2wX3MhuESS
4pHLs+AxtEp5GKPuPNTDEkB+YGjxot7mFvLYwlyZ2LcUutOBHIDuOFC2MrYW6uboBcEYvnN/aHH/
N0lU+P4vfRna2OE8QEMf7070Gl4iucCzfuC8GWPfobUkGaT6eilBe3SZvVK+SOIx/NC/Sb5IDARb
dHqHk3UVX5SB2qFi3Trwo4mQKNcFU+oXHuX/M+7Wu/eHRZCG7nnxwZlGJRsjk9bSg1zynJMmUDM+
VAM++h5c3bKeIAABtU1yjCtAgcJNSjWhieuOTianiCEkXVvqJ49FechPsY8tl+w8dJ/z33CyuSJt
cKdtlNU/VzJvdHPLQuFy74YCNYxGmz+kjJr0ZDJmdkVt9gqRXSIVCA1iiHtfrDLcoE5AXNj3lx1N
dgazPPhRAxPeYPVSGsUuxUjrDriWGati8kXgHFltEhh/0PrXj6Vq1u9KkcfC216nc0lJZolPg8H8
7ZbFwgl4xtBbLBtmjjwZ632DFmLlB7sFB1rK0NDUW6gepyNMAAuUJJflrizHc03BXfpnYg8tXR3f
rXdErWe/VcT6lS3RARGw8BMuF6w5m9rq4UHeYmQvwxEkU34iYOeHxG6kNnvmuqzgAnI5/5whkVK7
wy37OfP2cyrOYpGcT+QLv8UGlwUbfLXJWbmLYCXjagRPgu+BqUbdj7mOCEKOEK0K3Of0TadvZOD9
T96RNTKv8EmibLAIX24Z5+G9vB4iOaQrq0QZAi3piQeZ/0l4xx4Qi+kF5/S1UljMb+/SezefjA0h
on0XFnX3eydLp0xpi3QY5eJhkbUNojlm9kBtJJgBQNfR1N9WbL7BWbRx5txP9cv0hGFdJWh2JGiG
p8+Kroad9uivVc9Nr2U/rVILhE6Vqyiufg0Ua3+nqfGekGRuwxNVmuukQ6HGKJfvjWL7J4yFIPgC
v5Kmv6pePZcCBScrR4JDDi2wfPwFXHDz23WVWf25qxRlHYRn/mgeT5cTQ3cermO4teqxcThOptqN
pndH5+SRl6fdljuci7xc5uB2f2SnQFu826Lt3yv5UL2dQvh3Owb6uYoE9XYEfAk0KVBB2n6OFhb3
ogKBNnTPaxznsdiasEAyOnk9ErY5jPp6WEpSbCrvvau46Mtx98K68Byg9bR5S71IVIu9KCPJ7/M3
xEcPor3DdRp+hxGrSv3BFKOdIrvFLahq/HaAYCQQZ/hwFwYnw7kdDZQFCFSbFrrWbZXZdDd1h6R8
GdOGsjOY1c5zb0qbImRQKZ7VwwoKgm+zTJsxhSMhm99l85sOGN1rYKrzl4M05xLrc+yBILMnQXyS
2qrEPOQzDkfV3EnFYaFZIeUrAip/RGnrALXcv5chjAGPQt5+ujEhjzAkD70Z91SDvMQdHgilAoYd
p836NgFaU3O0yjeY3WWcf7m7sSSKYlr7CMRNZRHN/GM8a0DHkhB5CSc+iMkT0mlo4BayO6VAhTk2
lmAJlpHcqKhovRU1/0zCibDbeQTo3GMxnlTg8wC35BcsVpfgJZEtE8FUN0VuapLdYzRM90I9U2pW
5SWst3NZ7VzKMcPx8zCput21FxavytZhzSoa8sigX10yCGldetJgUcmQbEVC+wrWDB4O2v/LOWeu
6RmAzjV3vATbZdA0/RfXZIfxqAIPmnw1WBFvOJSO+iJK7lVe4bsbG2dEXkZqjlhLt/J7AMayqVIU
ltrXXLiiN5apNaRPc3RS3MBTRqbBU2OL0Hk3BQ78liBLDMHxkHMLu1w5EcJk7qBjbBcdanAkOHKb
AHT4111OR9Ekd2yvlIl+jkyspGx9W1Z5KiCEoWwGSR8HLdi+AfYa43FtkGVlW7U3Xj8Imp38Muoz
o4RgHoQlQ4XIuvNHI7et4Zr5oDTNrmhpSt8ao3/FJfneVNBufKAAMmQOzYngbN/68wssufOxa1ay
1QmIg9sWfb48SD5DV837NMTk+CbG4yfVd6uY4rjysM9QB46H3nevc+KjAZpmchUUya/ZfDHdFMlV
VC5mUGNtBam2ge3VQY1MAawhdru1bZPPuRFd7i7HTmCaH2WesFxQo1plRRDCXyX/VuRZ9ya3pDAG
pvUelL0aWu/GxyLemamDPWp7vJ6EVqPofzr7sDFknqpL9kIpI+DNX+ETqbtNzT4JMh4CP13qPaEx
ioykXU9n2QDlNe3k6H+v5rYCVr8TrksECZWPIO1ubjoh/mNBFMl1QZeAsBra00C1rmN7tCoLn+Pc
WfeFlzwEogXkakGe+qJgLHPL7UsHK/Hgk2YS6ujPDI2VDFRycLUZ/TtYCSvkxRnKoTKY7S5GYEB8
5O1EBBTRAPAtH6pcz9OuWU10hnduPR+evu/0yD/5FzwL66ANXejWyHziNRYKBrQKu9HDQMSMdFit
XIsnFLYFKMoT6ElcglxhrIukjOXDMx3NoXjftHR86RJnxkAptlDBDBkGSr/WsxMVXaFqEiJpfTNJ
84tJROh+CI8hyEe8nJEiEpOEznSqSMwO216IDPVdnkcAxPiyf+Fk12LmANn+VbAi2aBJ+Z75FuFh
e6iaEHKfeclE45MhVbUhf09TtlGygiThyt7G6yvRDXXdQQwLupeZSlEMto+1FNkS18mO2S6gNEIk
QDZ7GXJZ+nuDzESQ3RYr7uMqcHThuthO425gwjWeha7BYpD8HTh2uIOK6Yvl9BMapOBRvnvpbLx0
RoNIrB0tG38KP707XQxfIfui7xffjH9DqnxPBmv33MbDtPlG3upzgXdUomlqfOZl65QRDSa7yoE4
FN0YFyi242cRXXztLfq+cn3TtpIhmC7/cGYNBDdQgAuYaB39KWCVAQ26M5dGTrM2TvWE79c4QD1b
3QYGisgn0NVyQwHoC82dLjjAbufIvtpczbgcu2g72Veyx3oSiIGWE9ygdq8nIBvk14tb4hx2iiM2
dSFzUzQK4T3t/zTCNNhiUs5vox9wys9Cr6f2pqMxi6XZh1gY9uP/CJZO+RJEKgT8gymQOEHngfhw
8LPgPJ6s3fVzcAY2USxjswIU+4aWwPIYRk0wJNQQumJrrdKoLrNClzZhWDsQLlKRAiY9IWLRaYQX
7jJlz7vzKlFDMOSR7vaKvYaWahuh/7WFjHreIyb2u2qUHpiBwnzFbIbJSSgl93zXLEDCxLORmn93
7+6ZB1ZEXWqCiJcl9yQhCSqt3jfKx47H+mBvF7XB7d58FXp9dlEsADXvSXhvWIlHlS6VbQCjR5Mp
14G6Py3y54MgSr6Rp/EwbwEbHo9I6vieU3JcmiSxFbhoihM+zV4+YN81yYMO22if/7WVQJ5SFGCw
xCyiBd6P/orRCsflhW2I3R9SeTGrkrokVIDwoKPcVmwx7KNLgRdxQUzi6q2Gna1anFciLevDxcWM
xkOSe13LUWP+0dGCj9+3WQ+bop43j8ljhs8EdfEZbU2oohQOGQPT6/urmrde9gjHQgwZlGelYx/H
bQr+PhGmGvB1C81Xs+eFEVTGuQaUh7YM1NJO0r9zWEMZRY41E44+KHR39Xh4mOlXMVRIWAkHec8G
RcyKleeuQUJ6RimBgCmrglf4QzThm0p2BRbQ99ULV58N33NG94jw+Y8MuZ5wUak+pr23Epx3M9DN
04C6CA+TZLPY/b3Ksbnm0Jev3PjcxzRXpBZi+praUrWXB1uX2xwYLDsajC3FYVFRCUyMftS6Te5F
zwm/OhZhKieRAliYmc/enWsbvEyDOMmgJzQ7XjUoDANBU9sHMjykI3P3rdl1t+t79C83om9cmd+l
AIJ7FU+T3zTxFvP7Lw8vYDNNyg3IgPDd2Z3bvAVIqbPErmiCpKh81m8gadw+4ZZeI/ykQcKPQfSJ
X91404+JHtlwkjFqZDqveW3zJM33ehA0J+CAxm8S2ylhokvZcc8LYYOADDEJUj/a2/yW0VgKIMJZ
/38kTBwT8rVKK8PHgrDfJhiVZUc4bEUL7Z8G75f449ouMZk1lG3mSgLUtgQoa+oCiRGNMGXCw5e2
1GAz+IVfUeyLuV7MnEbmCIbPTBG07WCJN33QVhdktMoxAnWS11meOlCyrVWYl4giln+2Q5/2EWQ8
FRZzk6pm+v8HRKchwd5t0P4wi+cWe7J58Ih6Q6GdWkak87K1zILus5Pwer/RVgQFIU6F1c826StX
U5KIFg4bk+SxkNXWgHAI0Mi9SOy4+FqxFJ3AtdZt3KtNX9F4pQJOn8DCf7+ZufEa4LFEFRYR/oHE
y1Ekky/3nVGx8TGLZ7tmpjEDCbTO+tXKQba5u/EvqmmKClOvFxLjkiJYvzEfRGBN8ewoV0Tg+jXW
t+uONhde06CNhqlQMmAlM1nEVQnD8DJPm4oBh9dgBzCvC5W00r1p9PAVQiTfeMjMjkO7LxSa8rAq
0An9StPEQsAtTNN2DqUkuiNB8DTnEUcae8KT+WMdb6KuUxdwVmffPx14poTq/dwWV5++4i+olIb6
kHCUf7r9lZaXp5aO+5b8xZckngrzlIaTDuuXhHUQ2TDNf0Boq+ml6YQQiwmwZC6lMSn3ytEDP/qf
3CxsyjYt0IxwOQa1GbkXCdIxdndtm2ZSpl3mAlhZj8B6zZP45tBdd9XRFgYu0VWnf/Onpon+HhAk
W5MVUIYGVZXHZPOkSAMf29XiqtGdJ5lpnhdvg+Ik0/kPAV62ByZz37KdOeZCQP6gmFQYPnnabyoJ
fuoaxAKvV1YJ2ahiaF30wl7FxbdnMOgbWsiSgb4XnPnpsL1fvna/WhsDOdPEcCQTUjzdlRDj7tJC
K89C1aiTIOgP7mEDVvGD6c3do3imqvXz/NU2iRVcIAGoULDvabTedG7XXfatzasBjLaVJHSytt4G
QhZZc/GHCBiGumXBmmgoEHYe6StP4u1P+Xd47vqphny5VtwX1m+LPxQZlE8Hl3UrWqf/Cj612Gmf
3ebuVaRoaXk9E+6BW4Vp2nuXpnvvowYy60UCTcOy9wcFX6AVhzLyD3k1aC1j/gW41jyzQysY2rfa
64Vu9X7FBlV0Hwt3L5RklWEvnLjb0WvCNVHKHiaqLzjJCGBJ7WaGif2rA2A6whe0+BAQTB9vfzVC
1PD2OReqPGjNvvD90yZ8aa55+b0hrumib+3G1vbWFRwIcudYAcVK51gV8OOvDI2QuPBGKrHtGEOH
5BVEtIBmQuAr+hFYz+Ne3+MvnxWEonAWSVqSnVhyvdlc5IXpkA7RMoJE6LqZPDpXIa2K/AdqTjUG
oEKL3fVBz0EAHRpoobN3xwNhg28aTpo1HLAeF/PKoqqlcdotJiaXGWmow0PVdGW+FC+cHFuhzncI
rwXzmv9ebn9Ig4ksYo4Xw8MhQlwVp3qxY2SPx0mYpZwePTHGEJ6zxxeNdwDLh+mUHnF7gt8wFTpR
VOXYbsr1ykGXXMj2POBP2sPlqoGbSD4HnPp1xyWfDnYZ47HjlZtCGDGaUjZRRd8DE2NN8pQhuUon
hjDMX7oU8OHHDGUxl+YPRpawkBgMMKm1eei4jtSU97x+AikoNFWlun9T++TSoLx4GTPzyWyKnh7m
A42InLeK27yaylD0js0IwjRgFgL/YZo8LBwD4NAbHHv3Kf5fgFQYqMd81vwZnLeCqagN7mzv+ILg
cFLGCZBhShzmKOXu/vm1YwFdsb/hA3SQ5yqC1/aw60frE6kTdh9LtCvqC6nxYWXlAz670NHfVkKh
yaHkYj2CmTqlVCgC0smDUzdxhDo7gRw1O/mHjnXFUMp5cgt6FiiqPYnwUFTjqGjq/ES9AnCHZxRB
fJjNmP6oQ88XeaLqqZx1u5NOqyIzvwJoeySOuvWr6JrT6r5mAPzfhsmYdFKkPxdpf0oWK6yqxGUT
oBxH+JSKraUO+Sx1wKznxDJ18v+6r8DNFhEHQNVmsuVJJhSLmpdPHHogxMnxFdcmKb0A/ZiJAF4i
yN3DBGT1Y2gRYmDxrnO5fFWCUkmTMX5/GsAzEqYMsbLbB4rI+X/hw3qH0bXsaGQ9L7Gfg2Fb004I
IiW5bZparClxAmNOvd7iAA+oK8YgXBcQlxZSz2LFAR1Mmf1FD4UzwnMShma2e2Pd8CVxuqJZHODC
5WOVvLetDZ1ie61boOgo6lVgCerUANGNXeTBcGEf+gQYgTITYuthw+JDbsSV0HqvBo5gm4Ccc8Rq
WKu2x30cCWFBSufYp1r989jSzgd6bYwz21/s3pc4byJahQarHS2ppOx7120XRtAuEfKEIpbLC4x1
zSOkgT0xBwaT/JnBktM5LSFYo+fBoC/jgh//lNOuC54HOLEIGE25my59CYpl2HwjLU4ssyOQI2HU
iatZSpF+JG/zXA/Zzxgx2hafi3DHRSmzKyw0sQokRc5Lr36t1wcXsNgyUnDfSuIzmzWiLeDhQW5f
ZsM5/dZU61DldVfz4OKOQM0wYkUCNujGlsgc+sBL/ZtG6xskkFpXDG2sWDj4J++V27/VNHg/tEXU
HWNYeiS6bMb8dpzGmlnKzi88raQxztZLg8HeTd5/pBtlv0cdeFkF7DlqZQ1GrlK1QlOteL5A5JNS
Scwn74L7i/X7zPN/eUh5YoUyk0Mw2llDcPjkyIVVU4tNWrGaOmxhZ0hExmJpPK/acpvtS1SVS4tD
OkhSOeJ6M0E2WZTwzXPInult2z9Y7XjSw+C/VmiBvz1hLiF/AqsJjuJwTW05v0uRjt/1W3zxkb/p
rhJGP2hKIiPZAsx5LibUKs4hHcf/4THO8tH3z/i7RSIrRcScKnloQYvgP5RNuj7I5EPLE8rJoqIE
cwz4yPhnYhIXi7LRcBkGmtGw5nDkSDQBI0HtZfymLi5zv6OLNrRaOowK/WfcC7aUkKLkztefF4/x
Ga42YRzAWCLdXmvqlbHEfND8j5Ky+wKL9mIF1ABQt8vCnNENQLI89TjUdxVQjEB1yLh3p6pzv6yL
2FFUIvgrKhu6oNT1xSXdLWZHpACOZlqlJbf898djmUWGdGOAvyYhiEcJrszXxDFG5ZUyFNZsLc64
QIDSSmgCY8jhH5lUeYqgsRghi0BKMZoECOhl2mEDF3JZMBK47mHzexIHl8J3XR1OEPZf+ZUFgt4E
UHcvCX+/g5b5plnRNkivPEugA/4XUFlNVVuaL386oBgS/mTg0s0ZYyyWfYsG4VJQTWjE0aUqTjf9
zTzlQR2ZbzkzpqQKNiEdw15ryxs+NVW0tvUaF0lvaf8DZaF6eH5jVmkZDuQBaDpXAkk+DhoSzmif
3bhCXkfd/ALDz2EDmUcAhZKIRBOZlK1cGTM5GUYo1IUcnrZg/fCGsAukrRxggOU6mF/Zi9hrcKwK
SDo2VSLlJGYLLop9HYd+gkjcwpH+XAGvnKFKUMaZdrGjuWF4r64vjKQfubh+3yCvWijYVh1pJif8
k9IjvNaxSy3xFMXrCR8qnxd5gcArBuBNhU/gmMHXEgPJW0JOjo/hqj2KP4vO93qnAGrzKGdY0WFK
HavqT4Hndu4d1//bQC6nMDqzZuDRH4QdGPyeNSfxAlWX+8t1ZlfUuxw8ayvXzTDRkAVqW0zjeb1Z
UGCaXk/MMovXhlb2M4bQI6ZU70JksrW/nP7o4ekBQ3OL/tKPhcTG8qP8ZJg+oDcAyBH8cdjSttad
p9zimu3g/CEWlr0+kmyZptoZe2KLZUkvDLtA+x5K9BnWZglvigfii5pQLKxHbn1GWOHpnC52MHP4
mDjx0iFP/kcyQ2NHu6c5ZUq5E6PoGbCboQ/bvt0jyWaSK6Z6Qqe4cNnm6fnKm5uph+67oxPq5yAR
Xe2fKixF8bwKZpugO4FeCKpWOzk/R3qCVim6Q/ig+veIh3zXSx9LwBCDEliBWCfY8N5w7b1k3EwC
CwxlBMf3ZahNsbuduRDMswDBtuwq3Mf24X0ceS3zGxuCOqQf2DTTm8puMCknpY9Ri9Cx5jF8mjCB
R+NPityEulG82G12+8dpU0MaOJof2XsWkFUPZdgQQ/qfVipGJZRr4Z2jTJllokkJdhX0Wi3Tj5Rr
hv5UyoHOXEBlUTco/AsGLIYl3IEl/gyfLd+Ua3LGKsHUB3hlS3xybMY79oyMDYS52K5eEum5690t
INaBgn2519KNbTWssrErjAoBf+MWJx20BHZ/cu2G+TwFIMHoK7mQbIxnbkIPt8ApZ+ClV+xjZNDq
hN6zKHcwjDtvxSu0IFpIx6FmIiCE6ihYI54qOzBPI/uJdKilsgDLYit39EgnRVlWfbCMh2IWFLQ4
1L6Gb6/DSrboYTMRfZRrNrwHSs6imDeDSlGKx7AsO83sG3v2jXdFSjyv5ggiy/Iq49LWRZjtugzM
Be/EKWpCMdKf4Md37Ygrd4zWCE1MC4CndlBNGA0mWUI/vtFjfveiweItLuKXP0cCr77f8ob5sq1S
zGsN8722OznELTbnE0Bw+6ZbTuLRCFMwTEi5fXWskV5ShlKeS8iSMrXvv0I8IoB97SaQsLieI2yY
ZHwN7JAULe70kL7S9ODQq4ebe6/YLG34no6qfgQrNAR5Yd9wBNpB34MR6ZTUK5kM7VUsbepp8XPL
fcN2jNyy62RjMdcF7p/bQpRcgDAKWKiBxET5lizvlw+kLFAtA1lXseFAcY8cmMpca+Tc+nUFAUdi
yaM0zgZmdS218QpQ2E95/CPuRIq9t1ImnqWk9N6vEp2/+10u6KaddHyO1ypf+w4htKhs7diSE2rL
nNHjs/x/BSB+XTwUeifvqwHYP/qrGI9Cf6BFfLBwjCvxvoqTydqrkE9PL3Vnos8dZHPPDu/E1cAm
g4y2y9EjHzNpG0sVrXdHIulAkFigkHU34HAZrJHcz8/PHom9PMBQ4joYX6h1/XCD1e/b2EvL388S
Oeq6uFISmnRxgQMAsY53lOw+dvAZoyudUIVQDfszZW1Cl8yOUq/vnymIYx2GsvhB4+xy4Skmlhat
8xvOkS72+2t218OKmPCz1hZ73Ie3QLjVrzWyz7P+cfdFppQeuZwEbpP6sTlldgIA9KrIlGktfNrr
dhjMT6NYhb5cI6K/gbl7n6uN6u0s4JCkEciWhZystjiiv4AnCms+m7L9GT+1sOKpreR5HCIlt+XU
G9rRT0uMKH7hAUrWtYhuPNp2Ukmw1nBsMLO+iO9HgDcwv39V4kWwBDPr82Qglw+p0Ph5VN/cqSoe
2q04u6kTAByjoH8h6Rt7n6n+bDBvMOdJRoT2NdRFC2hFYqoA2ypOrB89D9p6KWPaEZkMUgdL4KDY
wgeOfe1ps3KoILFXt/B5ODmdSYGKXCYCIjlPpb4rWkgnvniZZnFxH90XtlbO7bnU8EhhqTgbIcuE
E1u6ntRxLjVPzqRAL5SijZD+h24dT5KqB+yt41nuyXqGQN4wWO3m/3s+At+ce9EcIEyXy5oZeo/K
/jCfuvxlsCoJ7ZzVeU5o0dA3jPPB7r/6O+QR7EGFUaI2IRduLAYa+xPzdbrpuHuyTAmr7Hd1brnu
LOGp4U6Uqidi1Le/exGx/QjR15AZmF5VHfqqjJUPy8Hz5HfgvZtZDoO5ottdAG1XJYuLYeGOvNTT
m8WOlU9XW69Tx8c4r7HLTffnuhY9nqVxc0BJ9IRdqno+Gn8K9P9ZgYa2U1aiPCIkrY7ku23wDgRG
OLzCaOWfvhO27q1522CW11/JG+R+X2NCjCRWzT8sVwG/AQpBFuFk8gsLmw0k6Q9l5CLWm/QoPk0J
XCUgr1g4pnbeivMQl43VvO1arYgqKpi7yZyy6ZcCmXQ0xhuhLHLmc1S+N5L92oRHEN9CP00sQWt5
UzKbF7+ZPg2XOmj9RbqQNlcQzNyZ5UQZ0QZebqID7Lk+OZvKcPk+QIocyYh7hHsY9HbZV2YGFX1m
axZuGi+xeTMm210MoR+ZdaArOzA2wOPSoY8F4JCvwHiuepvfNmZPNdyQsRJBJPOm17ExEXdyEgWb
XsGRc5yTaRVs6FKulr3ZHuVv6TEhF506hsCYAsELnNKYmgb10uA9QeOU8FhwyRJt8grrvBomOA4R
OwLjulMOIW+oItaT8ChQXTSrl5EHK7Ts+WJvsCb1knCihoBbPMMA2hKMYiEfAOllnXrvuJeRvKJH
tqDevXNTUaGjmgC9puC0qsEDOqHFMfSbPmdKYOaIqxB09kjI5Ndx9rQOVL6tpFvaQyW9+nCo9Vig
Z4xuczgh7MhDbAUARWAIRJoLPXVmNlrzbCKIkLPsDNc+PWurXj8tpcgcXebabOoTDb3iws8tkCE/
HXtAcqS2AbygbLTYwScslgGjKv5PUE7dhF0HLGDEkElfRMT+N712sTZxSlb8EfigNZLHl0a0DvQx
ViudCCNs8xeSZWgE11OF7zSoFx2ofw6a9Jp8CB1Mv2UX04+xKJZvU1HcR1sqIsdDVwSZwAlNRRld
kLdp3X1swwzQIgA681lxA5LS9eWQ24aJV2B49d8NY5Eld4E0+bceQnTp14ldYhXso7hVCHFXy/FW
M1pxC/lUgX4Thg4IVDRwBtW6Zvpti1582rwP7Klen9D5LAm3mkqEsX+x+XUohdztAXyYdOG3jJbS
kmp0RWH7iC825PYG+rYFCbA4Xk4yTPcrHixRicHvvj3x0Yqxyo1IjzM/IDH8cedXXaYf4ZzdPk7I
+ecGMjL5n4VARcbuhLiklAVUT5hBywPl+Z8EvsTUM4al6Y2HQ54pfQLj7d+h8xhalLXgAL5p8rM+
t5x76W0DkYGollAmXaYJCsfL0AwgyclPZm5SoGlh/8n7gmwN+lIU7QTaYg2Ezo6UHh0f+oYiZaQj
cTo53DpiN2QEuyfUSM9BaEmD2HX32IR5iMRwAIhoi2pErFqtB1Lv8L8FZ4RNmlMTUGdUWhCJk3Xw
VlNGE3Ko60LlBlUPqNThE9WaZgQqR5Yq3i2MHJjEYrissap++CO72nYrygk06tYnI3niBdZBHPco
Wpj8nr3rivjFzlDdYz4Q/EhhDpZirqtVbhgwUmNwxXZ/swRQvG+3Wcx0SXp3Lx82FOHk2Q9X4MYK
wXLEpipDW+HLAFPRYwzcrH2Zh8WswxHa9PnlNCZX/5/81BNb1F5GspOwK+w0GAX3ndL1uj4S7iAu
L71cSu8A68+b+V3dDreuegYTtmdixe2HXdVYsVEztURm1Jg8IGiWCGHRTSrZF/pbsnHTD6VFB7kr
Lgj2KKY306rycyVbUPyouZSVsWY4mqD8lxFwby4uGepSW1DWvqENGg3vGZDbTM2FaWCkYQ1klVVw
4ufcVZ6kN/1C6PO0O4V+ujbNTY+0DKDL1ykXKfppufuLkepV8xHZ+dJWbd5oFOeuFyCUMb07RxXv
J0rkZa+o8nbxUzGahRdh+gprNmNsDlfecaDfHQQz5vMYvOxXElSAScyUVNCHlozSl4fMPY7LR57L
pPxQQLKFUAiwm3Ri7nZ8/nqXWb8SD7mreAioznjkzgpLN69esOwOaeS3+ABmdAZ3ifJE+IijSpXB
dPf7W5469Ub46bzxRzwS8x/7o4L+cbYzCtOHI+lgjQPU66hXEKK2dQpFsC9Z7M9HN2duiZ8q78IP
t/ajxewD1Mrd/1IFMQAbAbWU3deJVGAI5+SGNsdkwj0DRDrN+PGAfKBZ4ghF97M0nTxNDRLX2Ffo
wJZemHzlPMWvFFD8CWvF/nXPpycSNVSmuPJvgCTBBrsq9EKpQHeiEnaIEZPacrTO95brqkF9BioX
aiugg2T+p/Rxag9pkXoOlYP1pjjc56FTww0DSm02IsuJgBzkdj5XNi6wGc9eSqZBcLzGCdgjh9vl
/52tI984C1lvbf3sI9QzLj8+3arOonEetRdpE4tf7N8R1xMFSlRnwAPH3ydvTJ5AjfPEPjyQobGV
0AXcCI8MF0xeMCHxMgNy4gDj3ghNh3dFp3J+lzWzFu1KlCBdV5Dqf77N9j9EvzQdGvqHCDdt5WJH
Rbf20qkMJ1uIGnoE6mTPlKggDBTerFHvVdT031zrfFBkXDcjI2q3Dh1eTA7+7xUw9kjvC0VTVGXw
hFHIOpUy06zBJYNa+rtV2jqafqs47RR1qenikp2sroLU+JEh1SwVSed4+dKcqQt8AXZhdntJad/D
OMEC5Ygx74ZKmA8gQfKBvYJbWDXNlD6Zetbq8dK+my+0Kv1OP0tQEoBdG7M/K68qtsWRqaMK4G4h
oCvZHnaOf7vh9MugtnjfUQrOvs31ufdg1iBlxIdNqjm6nVvU/H79RWba44zRsOEj2Hvhiq4qYK/w
y4C4LPeHaxyMazTpKLzhsFrowICNyl2sgjPcofZc6ZVu6CQG2W8g5aYeZqTD4UjthAfgYBamDK0+
+u8fzaCYYaG8yD3d+A3Jyxq+dxF9/bA2HVEm1CaVYyDSYgtA1djc6cDh4HP6qu59GNYXxE0=
`protect end_protected

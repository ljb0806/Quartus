��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7�����������	$��BR/�`�f����=|o�hN�<Q��^0Fx{!o �<v��	 �[���y1�E�Tڅ7I'��7�'^#��́��y�'�a�� O�KEʇ�m����@��=P%#3��(M8���p'����U*9�����J��Zm�;�}j8X)��Ӗ]?yMm����mN.������j��p�]�H��%Xg5Ԥ*�X���9y�J���\���7{�f���]V���^+�F��6��?k	5�H��9�<���w�at��a�oA[3�r�QA���R'�`R�^�鷃07���)ص2����d�\�跮�:�˄�	
���A�6�o3��/�i�"4@��{�?a��s�OMXvH�-�ϊw���՚��r�4N�pZJ�U�y�����yp��6Uָ݉�	l��n��T"C8G�����m�>�\�BK�J���^nDC���u��,D6�ਔޗ	�T���O�}:A��^�
��Eɉ#��=6��P���q�����#F_?�~����y�Pt�"G��)Sfg��� �),�1ɕ//��>��WW��"�U��n~�.0k����(����>�NO"7�C9�#L�E�����L!MA��02��l��-���������>��1��N���3�a���\�'o��\�{D&���E��q�ҬJ*���m\���G���N����vM�����7;�ࠜsQ�({��D��A�De�2.;4�T|�
�2���oq��9|����r°  �lR0Z���M6'��&�����y���a�y�d�o�cv��^eD]�)�Ö0l�ƾ��:��+<Xa�o=��)�!��T�RX����0�Q{�����nd���8��̡p��c�^bQ3Ë�\���<q���B	 W�UcQ��Z��,������܂r�\rs�A���9ti��vA��������&����I!Pi�vw+���i~�I]���lL�t��"���q.,a�R
����Lۗ�d���g�Ef�t �l�{����3b	?��JBPQ�Xa��B�Dc��ߟ�f��N
�fS�o�\`�_�H���G��g�k���!�9�bx&��*�Ȯ]��6�(X���O�^��a�9���+�>O�N�o��I]�ϔE�yO�Z1�E��/��j���JdTa-lUh.?`�aî$C�?~J�f��«	���棃3�tmji"6q
吻�iQ��u��aT��C�dI���^vo� ;�^.׭N���`������¿]@���]\{ xu�*H�E*��S���榟b��mQ|�o�ʘ�3���O���!-�~���B/��~�GOS�-F�=K�d�4'_v�Z����󎬟܀3ڲFoзi�D�*�,�/�.�2c}LMT�p�#����;�:}�,��O�E)u��#�Y�.H�g'7���{�ů���
.���J�?ɩ{�~D�^�>3!��
?��T��
~3����X54Oۜ5PO�%Av��V�W�d�t��oy`�#����#"fC:�{�����/K1���{����	�A��ބk'��L� �G�� ݰN�"~�L9�^�_N���w�|�ދ ;w�y����z�<��B��O�/9�]CR�?ocP.�x-��VWU*�}�!�W�i[���{�'k�� ί�q�0����^�-�֠�GO��4�l}��t����BN�M٢�u,)p��	5	�X
���5�:�|�撿5q���	���O�[�����?������%$ٍM�Ӷ����a��@rXΦ4$��5%jHq�������o�,�����5+U�mk�����6:�j�ܙ��q��B8<z�M����W�9�Oc��tK�h���W���EIQ� ��^{;��%a��E^%�y���;��>�b�/֖�|Cy����C�F�+5�dڙ�}~�%�X��L�Y��I��e�5���#�^Ӻ�m�f��-�y�ΏV���zK/��5ڣ��r�?ƿQ�>JH�!G��{~��̏��L>�����7��6MΊuE\7чe0�6��Ӵ
�v�2��e�C=�^����$�w�� �����)��%@�k�KB��(U�TWӪ(M�5�j]ё�,�WgB����h�Ǎ8G.3^Ы�i��B�q3�;��l�������dn)e��
�m��M��{goFX��a���P^9A���ef#5{-N!V`K��t �3��� #�7��E����a��X%�3Q�[YٜH�(2{1��L~��c���xM���2��2/Oĝ`�T�|������pQ�
��=��}� �uI�k�y������۷����n
u�# �W<ʺ��5�h������J�����H��DIb�;�ں\��3h,���o�`�p����G�\���|;�Q��}�?:�×ܬ߾}�^%��L)4���`��Hv��yl��MJWT�ŵ�ײ٘j#q����0���my ��1���n��#d�p���%?���k�~�� �,���:'uqZ�^�"O���\�^���l�J��n@0��@x�',�p��i�؁\�=gE �-3H�S$�� ��Bp��y�~j;��/y[h��Ҵ��,�4�t�/Vֽ`�K�x��γ��Y���5��4�wDe#}P|��ρ�=��Da���'e2�&e��ß�g��ruo�;�z�1q2z�-Q{9���y�2��d���Y;9$��m�|i���]2>/�#�gy�ҝ�)�	8�Ɔ6S-���1���7����b�O��a����SVT������Yپ�6'cܾ��$D��i��c�!�>^]�v���>^���Ej;N7#)�gMc9W�`:Z�YA�Z`���
��ksȢM[^�3N��UR)(R�l(b!g~��亄Z��f�6��+�X�!ғMHW���'���?|q���4�I������eU�� �O� W��PƁ[�Fq��Ǧ�e��?����YAU��*6;��|�q�M(���M~���``�U�������DA��!��&;��q�Frj�8�ϲ�iH�	:��wC�]�_I�%�1Sv��)7�8�X�jk����ԗ���r�[�4��Nv��>��-@�C���#�I��w�nLޯI�Z2��m�W��Ao�ȯAL�CNU�Pwy9��I��U��T��_mט3����C*ɐ��|9j\���`��b�xD(�݂h [�I1�b�ͦ�EK���o�-���<+��z�}�`����i�.�)�T��W����K��������MD�:�
�^��v����n���'�sa�k:>Ŏ�f���;�T/�{���#�>���8|� K�]�&���W������Q�^���y���5��Z��uvg��2���vS�	�z)���Nb�$��m��jmPq�ί��UZ��S4�h��l��l�|@j3�Z_����2�`�*���>��6��z�Vr���ĥ��LWUV�~�'���q���EL��kFJ�2}X׳�����H*;��R��އ0xʽ��o�~TW��`zF�0�U%���)Yٻ���q/�\U����Y��Kh).����C�ڸ�_��#N{�?
��eS��
�-��-V-�����+2���mjD�i�R����[���"��[+�+~�T��%|�_H��f�Cn�5j��ɥ�h��������r�&<���Ǻ8��q��+�>�-u$����"?�Z։|���06N�k�q�f�?0�wΕ�2�A����r�������b��P2��`i�E�Qt�	D�5��|1���Z�,�aN�>���>�}/���_?U���D|���̹U��l���_C�q�r� ���z�7$�-�]��]�-���z�AF������<�5��Z�=�;G�pНs��!���m�DJ�cid��z�hڧ�s���8h&�䓊�_�Fs����/K~��s��8�G�d:D+zI�^l��܀�Ign,�/{'��:����ڐcc��H
��P+O��i��u����ō��lt�Q�=���)$PD�ՂO���h����0��&u��yJRh -z���t��e���U6��De#���쌻A/�-��y��浿�����G�Էe��A�D�iw����<>|*����{m��' ��:���ZR�R+��I�
����=��Wgi���X��v(iP�z�%2A�(��x��F�F��ʃ�a�����Qlȿ�:�S���D#N���h��W%7gr�XR��SG������ƛ�Fp�Ś��[k@���Qem�-�� m�V�&�������yJ��÷�[��&z�%�9\7a�dMՂ���[53�>�Xm"��谵��t�=�(�!b�;� ~*Qեkt���{`�nM��獑�'_���m���&�N�ȉX��F�i4��sf8M���9��$��pkip,�R��V����:�-^���/V��W&x�#��V���Ԟ�~?û?��MO���&� �uŎN %�mꯘ={A��r�/�.*t�a�4�^�L�����:B��t��Q��:�߾���b�@Xt���'t)������S@mrX���>`� Y�o����0��|��q����%�0~��c�S�p��1D��->U�kYA��n=�*��=���þ�*��a{d�=��֩&2�*f�3�q��=R4����t��xX��r��3^�Um�w�A�C���3,�u�a��oM��B�׶He� �l'��B:e�&bB	O��n�#^�s�z]B<|���~Kr\F����:b��W;�Ŀ��첫)I�$&7v�y���_V�rfh��h��Sp��o�`l ��f/g����B���V�Q�\�-�CS5����+���&1���S>j�nM9K�æ���g"�׎+M���ݚ	)x���/3��f4��1��ͥ����UJt�u�V�Ϸ��.Q��#��>����+�����`�V0���JI$�Իow.b��H�9���L �;.�I��N�!���-n����+��EUH݂Hɩ�1��|�v�WvTۍ�I��P�k�%IC��\������;/�?%Ѽ8l��27GC�ISh�3����s�r�-ܙ�x�Y��y4=���w�0�r��9���M������-�iYr1� ��q��_��z�ۜ��u��+{u���Ь�t�܀�_����g�����4�]������d�6��gܳA��B�ּ����P�t�Υ�p���<Nk9��8F�	���_SŨK!�jR~3�G0۩�(~ߢ����l��jC�q%;���!��v�W�`�6�D}f�<���^P�S��\{�#����9���R�/�c���@^l���ѻUO-i)68�pʿ��ި=@`e��-�쌓������m2��M�G�PYc�iq�7d�!��2����,&*��1�J��&ģ��n9��W�H�nQ����i��7k ��D��3��䶮P���H�h����ퟝZ*37����ު�X|��g����P&*�\5���}�34>�z�������_����kԞ@���,%Oݧ�h��0�<�>��$��T���K>6�o�Ű�*�$��md��}c>�D�%�]Y�(H=.T]��A?���pL%�+˓1�E�*u �1��J���~�I�έ\G~�5�\��FU���}��)n˃yj�NʣtB>�^���#��'ϭyF�4�Ć��r���ӭHU�x�j��]�6�9���OC*GЃ��FHFFK�d�n�����_h�pZ%1�b|	o��@}��st}� ��)��w�K炁�8�d6iY�l�s��w9j�g�E����t�t�s0P�_ !�܈�?��V�Q�
V{�(�2�)�[sl)��#�fο�*�в�{ p=K(3D FN�&�u��5J�55�"$��Z{
��2��D���~#vׂ�ZL\�\�L��mK)�r�=���
�b�`L^�T���/��W]8�����Pˤ�脏]L?t���R�`�q�S�hP��]��Dw�x��>�}~��~��[�p�n&*�;Lr�����tM��S��r�V�Ub��j�U�n�)�:JLYAlZ�N�ɵ����H>zb���KSKmG�F�$�߼L��z&��ƣ=h��=�O�˜F�Y1�_�K҈��l�R�\4q1��d
:�����Gq����r��{a�I!a��+Y�e ��S����b�Y�����9��xlg0�f+��ؾ�s��Ѩ5V�f�I�L��/&����s����}��)o�H�5* ���@z��K�A�q#�9?O�y}��t)Hʋo��R�
��Dd���Պ���64�������NJB��ُ��/:=�Y:�9TՖ��W��}/�V�F�T�ɡ�l�x�H��n�~�~�ز��#��MH��z���2LB��ѧ��`���@Ԯ�;Zz�1����}�����cz ڴ�Zl�R���H|*ו���͹��n}06},*	������T�W��k��-��v�1����T��W�a�4�A|C(�dO�56χX��72����{_�э⊴����H&�-$!�*����>QG�.��YP�?5���e���_G�����{���^����;�/������|>��yz�����C�����&};����
�q���:EB�6����ߐLX��OT4<�-�A*��gZ�0�����|��`Ş��8��-֔�Ԫg�RG���*\Z>N�n�g�F����Ӕ�1 ��19�C��1���AB-�nF�τ�b"hZ��YLl+���f_k��"�0������) ��'J���e��Dg>��V�1��q�3 >�zJ�����\� �@�����a���f���Ae^K"!x�f׈?��b5@�Ný�������w"6�+?�;i�1Z�<�6�y��.j($O)��m����z��%�8=vF������F/��M:B�F�%���6P>���HG��v�~;G=�ֻ�O/Q�J�xc�\X�W��U����	�S�Q}&�c(�4=c�!�9���XFP�hR��F�h���?�Jx�k��XN��&�]�$���Jq���W�Oֲx$	+������ݒqs�
�L���̗	�D��3RmΦ8��3,�� ӻ�rG��]O���g��ʈ�ƿ3�/1�!�!~ ��{�G���j�������[�3�]7�%�B��-������B�s��ݥ�5u��=RNqgݷ5g�� q�t��f���f^Z�I�?x�9����о�4���rou����@�)�
o>[CWVL����ͧ�[�s�~�凝�ȩ�t}	>1Я�J�x��{ߑ��	��+Q�9+��q��&W�U��u�U��G����Y"d��=Ҙ�,M~&&S\"w2W�	�k㰡g:�\dU�.��Q��i$篕�$�/P��9���XŽ� �ܰ?ה��T��A��vi�ߡm��~�A/Ü��d��Z=�q�u��#��k�ˉ��Y�|��(�@�h�JG�v_���
��cѲŲ�p���JRy��<-��a
���7�7��s�6�_����+`�V��I!%����#G&�t�m^��h�#��y��l&�#��������l�t�"1���"�:���{X�B�:M�����o��Vݑ�D*=J��O,Q���4w��
C�2�g;�W�L�/#y����&c/��19�|�'��:�I���r�&s0gė�󿑔�l>� *n��ܲ�3�3���H׉�-|o��$�p	'���J�!��d���Iѡ�棙g7�ۏ��!�ء0�E��<c
S"��.��3�K��f �A�6���T�Z6E�E�*N�@v�8u�(�e����͑Z�s����X��	{�'��,>�KT;G0O/p�"�պBc�x�*���|;�ل,��˚�=rd@�q'5&��!��������:����rb�+z�L�m�r��B�}��/�X��Q܎9HO��}�$p��=�B7'I�Fo��wR��$*�f�#`Y�F���p�bPA����~���Zߐ�r*?5�AW�i����O�o^�͚�m��S���?i�ݘ;�����%��0���[�=��1�J1I ��I� ^��խ������(�E.`�,H=�t��՞*��k2�33r�!@�E��؃y����-'X���h[�}��
��P׽��ο��@���`���(�9�m���s�W_�������ă�����P�a3ֆ��7S��=|��5|�ٛFU���\�@�J�#�x�O!-xI�@N)�L�eS��r'�#IC*��Ŏ��(YJ��.u���թJĨq'Ѝls�6�����4�x0��2{��,|�ZS�uF�|ʬ���4���կ���G6�=���FǴa[����f���I΀x3�r� 9[%n��"��G�'y��k	��?I�#�d8P��uɚ��U�ԁP�%�^Fn���	3K�W�����(Ě��0&�|��5Ũ�&ON?*/�7���/��Ȳ'�z((ADd,��0�'~�N��(�A8d����aՎ�xs����}���Ǫ�VF2�9"�!�R��{��B$f��T_ƸC�]��\�^��Ʌ�r�>;�O'Z�8���{n��Ŀ���Cw|B�FT���
��荰
n�Bp
������L��/ �Ȓɿ�.��چ��H���DѣnP��d#{a%����ť�B��`���������T�<!�f#R�;)mȼ�����v<�u������p� 1Y�8=N���G"�� h+UER��);m!��N� ���V�$8��Kc�'>�K�'��i[)?BBL��9e�T'Ƶ��(�y��
�xN%�_e�Ce赔���t���>�g�<��RS���E���?���`���}FE��K��S��'�C�OQ��N�Q8�.ퟚH�߷���� 	�Ԗز�{G���~���?�9�����TY��ߠ��;H��9�����@n܇�$.�҇��K�:����l�44
��Q��z���t%)�ājXR��_������L,���
�{u���?>(�M�d�>��,1���f@��̰8iy܈2��u�S�9"��H�Y����7��_�w��ܛ�5z����9��6ihw�+�[}S�4��w{�O�����̓�U�\H�}g�p�������:�u�I��e[�:ɵ�N�gJ��oe6��O�p�B(���[Ծ��e��ʺsW�g�� ޤ;�å�=�8U~�o�g�N����6���)�/����r��vɘB���B?�<Cq�����DN�`\I���ɿv���IX��߼��L�l vw���{�;��ǅ�\0IF�!	��8����j~�9�ixK���g�Qh|%դ$ؾ�I$�1N������0���	�o"<�7�զ�Ҹ	��ݙ�I�B�=s�R���E�S�x���3�HӲ���zE�V�|WNvm�L!B���;kO.P�P��3�w��^���3Sh�  �����:�%@�N��nf�Ua��ﶦ�ݡ��-���iaQݥ�!������tGY�qDf`�T�5n���6�{%۳�䬵�X�6>�>�MVS��<�9�"�~���;ܦ��=�֒���4��2���T�3���BXX��h&?G!w��d^�N���fPz���S������ilJJ�L���t�қވ�f^�>1"i�.�����\��}�V�o7^����.4�j��F�z&d�F�:�k1$�9�X��''}'#r����7U��x�'vZS�[@����+�'(��ַ�����J ���������oL�R�ޙ�&rt���� V�r����c�a ������nD�#��H!��:��ߠ�V6�(�Uđ�&��z�q>	�6��ټ�A5�Vn�2B��-�����d���kx
=�6�~X�8��(�a���~�Crd��NVo����#����,��.y?�do��n�No�1����r��W)�]��3�L��L줏4�	�����g-v
n�[u.S_�9ȡ��X�9��l��#_�Ȫ�v�����7�j`�0��/3rsb�%�!T�4*�`�d�����Y(�h��$�G��r%�A�A�Tud����$�n�F�V���Iw/o���(J�xj^̆�� �.�q�H2t5�L�F{�����S=rn�B,���f��d8pKQQ�����DE.����=��y�g(�agfelN��X���������-� C��g|H@��KG�����wp���3J4"���3�1���fʬ���9�P��X���D��xf�E�۔�2i1�)�P�oI[(�Q�u�J�����;+m8S�yT*Ƞ�U]�1î��|�T˜��ތ4z���Q9+�F�F��(�Ƙ����?_�����@b�S�3��k����ȸ��ف_���}�<=x���Ϗ���y�Հ�2��'����pNA�D���ͨ7����$L%�G���S�1��� I{MF�kK�ʭP񒈀����j��� ��Xn���� ��H�K�ٛ�C��ZGTT�j�G7�g�� �/��'`�Zek_�]�����$,ƧW��V��A�֭�}9�4�ŀ���� yk�Ї�3�,���\������J���Xh���c�^!�+*�IJ���@�^�6��c����;&iW~i�)< ,��%r�?�  C����[����t�����w�9��iy�U<Z����{S�rF��T���@l#ل���w
H�	@�؛��]1d�b��f�,^�9��]w@O����|gs��V������uFO��:�}�_�`[�����vk:���~ǀ�^��Vc5������j.@�ϤS"8^�߀�a	9��)e�O^];����ԡ���Ru'���+�-���z��%��@`��u���m��.�TUΫ'��Ѷ+�B+Vp����?��vl�]���T�ث6pW��^"�l�`���3��^��,7�-k5#	n�ϯ*+b���#����n��,nNq�/�"��J�p���9���=f��O����-�����6���)+zJzև�Ǎ�[�o(�^�(�x�wn�ң��vt�R0��sp�Q��N>[g�N~V�/�;�I+����Έ��7�G�nuN<B&�0v�4;gƩP������Tzg8t:�0����C�5}�u�"?���ݱJ���d�pj��c�R�O9�O	c�(�PNLI���ػ=�r���Z�j�cl���3y�a����l���Z�>U/a�����&Vi5�;/�,o �|�&߰��)u�I/��p������WE:D�!��G�׸�r���]3�/����QE���1J�=Cl6�^�NB�R����iv��h���Q����[-�>e%�����L��h�,��[G���'�.�x�Ck�v��#���Y�77����*L�|"��g(i��+��eax�'�s0��t|n��F�J�E�̢&_�G���N*jj�8�S���dx�� ����d��4���B���j�.�x������j^%�����Cp$�IpO�.��:���D=����)o���`�1�1��j/ð�	��Ĩ0�-2}�^��s^�ՕH�ȸ�V�3Rr�}/�qN�E"�h���)!X{��
/���(�Ĝ�vm�Ѭ�S#G������^H��1�uo5|��1�0�B�)q��˟	��Lʓ*?Y�-c�R����5��S'>�ù�� �؀i��g8�V��D	$[�h��L3I�g�m���7���Ӽ.Y&U��[����C�n��t���u�B"�p�E/�0F]�ڗm{�n��H��n�?�7�;j����=*�j!bo��]x��1) [h�
z��Ֆ�G�B�Y6��	~ĴU����\��(����Z�v��z�[� v�V��D�[!��^�Cznf-S&���TL.���=:A�N6�tp�@Q�P�!ҏ�Iaј��*W(N���3�=�cU����%�Z��D���MxG��L� w���+��%�� ���Bs��*��b�4N��L�3�z�1nTdY�C���Xzx@��q(�����lKe�9N�!�6��Rin�l��O��3�ƐJ�ArlfK* ���������:Y�����w��}d��Lݪ���E���/O_Ek�2I]0F� w����!�_>N��
�ci�s�-�(]<�`\~F�(��h�r��(5����H�Q��?�bU�h���<���6N����SH��5au�UM���^`�ݒ�DDQ������l�6�~���O��~�qQe�w;�:j�����2I�
�O�V��Ht*y���tv��ꢪ�U��D�Ǜ�1m�d������3j6�����"��(&�X0���������
S}�e�����mP�l1W�v��e��Zu����� +��ڙD������;_�2�1
`�iȆ F�i�5��L�RF�C�zN�`��L�~)�d=t��4�d!�b�V9�-X�ӽ�^���P�W���X�����@I��"��yr' �0%3��(�1աS8��E��!�:or3��/��	1+OľD,����+�%�q�� ���g�[hj��!�����ƛJ�APM0S=?�y����4�;�tdz[9�fr�z���O^'��or�����	j_nY����rh�~�4��8ة���d����e�b!?����:$�N�g�	�6�����߃l6dF5�q��0�RG�:� z(�f���NMę��9Y�e�N���+\���`��۲��в�@����o���6��u�s-��F������PВI+ƬO�����VxN���R�������j-�[��s����;f�lPb�t3_�Gg������F�����+��=�۶���ON�E���j��$� i�]����~{x�m5>��Pm��Z5?l0���J�t<6x��e��MB�A����t�_���P�������t!nko��p�h�<��}�pA���x�p�Õ<��	�޾){L_#�|*�l����+Q�9�q|�?5Mx�l�WXr
@ӄ�p�E�����p��&F��^�{.b�3�f�&�B���dXJ���8�����HSQ�����[����E�;���4�C����A�����Y(xR���D�aky&I?pş�*ݱl�# �R�扰H�z��-K}YJ�����Ȣ�!�Z��[�α$ݟ��f���+����� �Y����WSW��E@��>���A��8i�!%�j�@MA�u�� �Wо�3Z���:{`��<n�u�a�"�������W�7V�P�}ؠ,���u�#���dX�pr�ɫ��0���c�Y��
�35�[�v��;��x�k�!���b��@w�vK���CJ]�d��B�9m�{��1��Ed�����YU�e�)��BiL�a���)�r�4�;"��"�_r�c�jQ�4&���WnN2���J�G��ֲ2Ԩ�p.i�I�᯦c)A�@� NU%p"�m�%��Td��C<2h{��4�O��\ZM^ݕ���b��ecq�R��#X���ݿ;�Z���$�v>��.W���u�<�JB��eѵ��r�(��-�]�)��-{e;�I��j���vF�&�@�g�^��t�H7�k}����:��C-.�f�U��J�d����p����)̕j�#��`�	X��J!�t9���J4���U�0��X�P�e��"I�A�g�<�aE�\*����"+��mF?9���kKmݩ�� � &���i%fr�E`�G؂Gq�_�PgJ�3����Rf��/��[��L���t_+���)sx�N"I�r��$��4��ܼ��GP����^P�O�H��f�k��G�R�%���������qsm��sc�I���"��+�mQH�5������hj���Q�ɖw"��H�<&�Q��>�6�MOW'^��P�����f�~�uez_7Q��F��R��w��})��V��Հ�P�"�AE��W^V�uH�:�s�Z��'��T}Έ�
���~�P�'�]o�8?�M���J����b����G�l�A�D 4�K��wp�h� i2^�֙�#�?{��=#���Z����d�X�^1�Gn@���_����exc)�f�d�sN��
y��לz����7��K�8���!���������H�4�!i#K;�p�����z�&\��/�}!?ꁻ��r�Nگ�u��}z8��`4ԁ�{�gП� (^�A��&�;r�U�]�;��ia[����7ɗ�-![�Ajz��E]������;���W�5�����]��\�ܝW�nR���գ�_�s����;�|eC�a�#�O�p����O]�}���|�p;oQ�I�=����=��%��*�Sa�cw�|��f~.��.�0��Dj����M�W[����˻��Ȯ�FTR�����i}�=����)n<WP��߳d@30����Ѭ)d4�uܶ�2��0���<\/�/���Z��v������hKZA����<���q#$6�2d��,��:�%]v��}���!�VSަЇ����?�	T�x;d���G���T-h���ӹH�o�J�����1�m�5��n]��(V=�KA�H����������-�mA<;�������y�[��c)��S�C��~���<ݧ7(G�/&1�*nj}t��͜�̶	�E\R��3��c�T�q��ĥ�����:`�͜g�_q�랂���4&�����m�<l.g>3�4�0$Q�����6�4���(?�Od�ֈJ�;"�D����Zs����g��G#)k377>2_�����s���^ܖ ŸE<Ei_KVg|V�8�Y�S�H=5�,TM\r�Yfk��n3��(�:5Ӗ/�ٮ�|����!�]�L:^�����v/���;�j�H�s�;`.�W{�|-ϥ�����c��p1
HW�DwXp�6��S��
F덕�,�3�B�	G����v�}D=�凖<r�u	�A~�-���d�}��������r����[�� .�^��QQD�\�rӭcdb�4$͌B��H���7�J�p\�	@��Ԝ�G9�I�b|�*Ig��>����)���'�&w�#���M�_���O�A��H���f`k�@G\�)q�-���Z�?���m�� N@��������iP���r]=�!�Ff/wf�2:�Dqk^���V�0쬴�5��NU�z`m[_k6��> _^�đ%�'��_��5E���?D#�C�quRw��'9�f]-ca��_�?d�t��W�	�P�a<*��.�}&@�ay_�P�qWU���!4=�t9��F�b�'SW�}����w����ǡ�2l���%�ގg�u<H���_�B8�
�{��$��O|$v���I��㦓<���_:�4Z��/��O�����\��W$-��7�I_� n�]�l����i=!�tf�#��Q��~OO���o��?|z�}K�}m�	һ��Q�d�>
���6C9R�([m~�%��:�i w�L���1㱁d)�͢'�xG/�u��T���Y�պ鎡�P�K�ݏ:�Nj��1�@eS&$��iP}F�ݳI�)�n��4�` /pXvư�5�`������r��J��>����>)kr��%^l�KA>�O�B��/٥����}-1;�"��E��#��m��� �8��ٓ��cxB%��W=QKj��_�fu���f������h��@��0��Ab��W�G=	��W��݀�ɓ|D�(�k+�,�{�?�Q���S�,���4�[�g�U >|�nJ���8�2�a3I��Jw�������^��_�h��!�iuw�w'�����K��qq��Y��#QS�ߌ�׀4���i�E-���t� X�򬈖���ypw5iL�Mj^�;B[)NrI@�i�ñ>ɲ
q+H̖���w�ق'����1s��{�H��v}�-�6�����'�ͱ�����>��� ���`\A�����-@��uc@.�A��I�)<����R�+����4�	���v�6�:~�U�h_X���o�ݰ~;�a�4X��DŢ�p�LWi?L�a�0�>��c�0�.�J���a�i�uY�]�Ll4� �+�����e׀�P8�Ռ-8���i���Gth�~�ʃo@�TRE�Q-�1*U�+��q�Ȏ��Z5d��_PLq�Xȧ��D���sI`?tBe�,�ہ����q��(���iE�"��?�m|���K4�����I_�Z�u5�79�f9B���x����(�TDY��J4�y<h�hh?
I��S�K�
с�xmS�9����:�����(0yK2�Z���b�3ٝ�]뫪9����������Kc��2�S�-�2a��e�2��?e��e�R�[oV��9Y�� �������٭!�ifoc�T�G0S�o_�tу����e��cv��	ќ%���#�&]�#�7&�&�^p��U,56���L��� ����� v� Em�b�1f�(Љ���/a�ң�y��E�dA�±c�Q.�$�f ��n)k馅	5��(�FSK��1����0)S����0��X���?��-����k�Y��qz��a6�+X�R��i��EF>�"�|&�s ���7}�
���4C�n�p_����|f��BӶ�Z2hż�����J�ۢiod�k��8�lK�<\|M�h�py/��۰i�VuGS�\x��[@M����p�O���
����Fr����z����tV�]�$�Q�z��cG�j#T�be�����t���PX��]�F7s��.G�r�� ��w��Y��>u$�SD��ճ<� j�|��1�
}D��_Ok���������K�)�5���^|p�X'���K�Q�j'�B	H�O"�I�q,���X���=F�H���\J,F$��F�s��Ж��/in	.�q%��Dq������øg8��x��� ��\���C!s�y9��K�{bq���*�kz)�`vH�h��=K���n"48���+@>����� r/�41V�ooE2��jF��?�)[PH �C�!����;���Lzw�$Q7�t�ߧ�y~oK9"8b�vY��kerz|���#)A��*[��&�d��|0���-^NY��<m����/�`�e%�l��@F"T�q����rQ���k�{��T���j, �MWr���b'��q�2�dgC.��xB�gJ�2s҅S�#�� ���2��&�m<[��'��y���{��=+�kF��@<�c8llL� @i�1���(b�$�~�Fӗ�ߔL@����� �����,�(s(�_���GrI����D�:r�$�6�
U�H|w�1ũ�����4:�fx���(L�����>�F�RZ�\1}�MyT�@K'\6';��Ku�<�'������:���I�|�c�7*=dm�p�s�s+D=�&j���W�\������������{�]�`��|�n��5y�yS�C���c	���?K��)�����<ۇ���$E�0n��F7�W���P�M��NN%��2�(A~�9�{�7��0�j!�߷A�W��4EYsg[���\�E\gհv�ClB03D���q^�/J�̡�=�4�M������U�":��5���D�$���'�	��T|�JiH�~bM��I��x:���jS<B��h>쥮,�l�F�N,`���^�P��ez�D���^�� _�f�W��ȋ.�5�*�pmOc!��8�b�]��-l���%�mPU#-�ZS��@u���>�	kO�{*��a��j���΍���0�&7�\�{�'�1�|N3q�P�o��O����V:�xQ�i�����ߖ5��t����g�v
�v�+z�Ə�~*��s���)_� ������;��!����c�N��e�lP�VQ�N )��[��-�(��:*���hW�%G��*qy�9v4��ٌ��|�leF!MM3��-���T0���\�(c�L�S��p���C*���-��Ot8!9!Z�kD��"���Y��إ���)꾙ݕ�M@�I�@8��9{�SE���񱶂�����Wh-��D��@#�"GP���ч��ad����q����P0���Lv1z��</����|Hei⎲wbs�d1��fƅ"�bb_�m���� �[�E!a���s���K'm��Sa�],�W7D�K���?_R�h ֫�$k�������)���	j1.)� 4��;� G�hq���LW@Y���+�'����A���N;�Q��t�VǈI�P�	�Zv�YMm�,V��/�d��Ym��I�-���P�E���&\�]�,���TN��@l[T�Bʩ�FCU�m���!9�b@�k��oq��!�Y�6�/���<M�*>�ѱ�=�8�u� `s�fz�y��S��ykqUi;1H��q�: �d�h�"s�/-�M��+:3(C2^�/��T1��Վ�W$��eӌ� ֧|�z�EBR����v���2��@Y*!�`��U��Hy�k��2�W!���?�&<n��Io��#��8���{�V$P�)��S�k+�f~ڒ���d�6���1'c&g=�@�L�/r�Ĝ��
D���� J����a9<C����5�T��SA�~��'�����O�!�YCo5<��J�f�<.�f$��z`���K/o�LD�������	���������R,�Z��ƪ����]��GV��'��JSZ?ޕd��\d�7`���udZ��ο�������g�F��oH��i.*��P!ֱR����p�ULX��D��D�Ss�e��G���ޜ�o��$��k����w��s�ٗ��Y��Ǩ��+"t~�l�V	�y��\��$�i�؍u,��e�Q¥V�Ъ�}"H_��rEa��S��z�Up�I)j^~]�:����h~Ƴ9�ʹ� ��1�tG
b����U�+�/��] ��'rA��e��u/���9� ����:�k�U���9v[�`30��E|6�,Ğ�ȵ#���T�(�V�ǆ߸ř�_VL���/ˁ٬W*�4T��;'_|���a����J8�'��.K�Z�xۡ	}�
v/[8��%BLd1��,��$@{@��7�:��IVΔa���Uv�+��1h�|��[1��I7��}7E�D�%2GL��Qn2��8� ���kބ��+P/yH`b(�� :bxH�I�4ʾ?�eM�0����v�~�ѵ�M�4�ؠV���_���G�LK��t�~*�<��*�����C&` ����^͘���z����eKK��VM����}ӵ�������lWfG1Oc���{Ї:@n���1 !:�1����nE����➷	Q��9�v���P{�JQG��(��	�%��%� ���"r�E3�f�Ch�l�i������F9 *�sv��� B6Z[���aU[[ТT�&�h���������0��ya������4tF�$dc�pC��i�.��e��4��� %�up�Պ�2Lח3��j.�Q��-�E� 
�3㳠�MnIS�m@|�u+[����.9�A�%�&.�(T 1�[��s����Zfz2#��#�a����!_s��e����ױ9��؇�+�frp�@���I��S�nwn��~-tEN_���^Z��,<^�2� n0�DZ��7�Jc]~$�8���젭�Z�E:�}aM��L��R3~8�W�Z�xӅ�߁8�Xl�d�!1�Vba������Q� �U 0Ԝ�z�����/Rws�g�-CJ��e�}��?6߬�ՌAI��P�fO G�ؙ���g&G�W��~��0��G*	4FF�X\�T_�.0�Tz���c>�>�QJ��Z-,_6�Ҷc�X|������Y����S�rf��@u5�j<e�N�]�?��k$�%x��/�V�q<)g�@�T=$��Sn�,�vLwM��F ������R��:`͋��"������V7E����a�?+g�)�6�]ȯ�����:�d1̗:����4�t����E U�*Y��e�6<���]�)�,�5�j�S �'��Єͻ�Q�@������i;� ݵ/n�'�J�\'vI-G��X�i�nX��(��)�8]kD#<|�a-�Aa�) �n
Ӎ8�{�W��.(�շ���c�]K���wicHN�׃�1����ʎ�Ճz� �������##�i��뫛8�6�W��)��U�+&�S�ti|V�z3���)gF�Ϫ7��cEu+�񀟥e��S>���/$6��n��_Z�����XV�RJƀ�j������{�<9�2�������������!,� y�K[MQt�-��������瞁����o�#�O�kFQ8�y�U���]zwn�,[�1���b�������-:�	Px�r�R�w!Ǽ���9KC����O����g%���<�DF��3j�*�G��A�k+�&�b�O^J����]q� � ~�s�A�X�Q�q_%lQ=�!=���]bC�3}����[�-��P��7��o�:�E�aZ�7����V�W��$���8��Sr'I��ᖢ���[��R�zV�,�ҤQ��c��X^df 7����ԇ�x�iq�5lV�>��`�QS���I��)ƶ�[1��1��[{a�d��{�;�()�$��3�Kb�
�I��'������<��Zךv�Q,B��2������u�ꣻ�<eF�z;!�w�{G�e��ˆ��V�28��胄���d��<�e�ǆ}xi�éO�\����W�l�@�V��7➼�x׶��Ӓ8-?��H$�"��WA�|*p:e� j�4�ܘ����\sKi󗏌��J��A�hel�%��v�׈��]j�$�Ӛ�0�H������B8��@F�B^��Nt�?s�M闿{�(���ݴN	�.N�%^�<w�I ��Q��`-�0p�y���>Lc����^�����'�tqc��r{y�U��~L:G��'��M��d��Sŵd�h�w�~>ح�3Hvx!��hP&����Z��q������␐��uh���I'����1���λ_"-����\@�|+��I���jN�"��=��{��u]��Z}k0 M�C&������zC$X^q1�+Eq
^^	Y&Z�|���oFY%M�4<2+�I��X�7�M�m��{��gX�'�|�kt��,��p��Pc����C��}T�@�����'ȡ�?{+t�`㎼�,�e��@V�%��%�^��0�aȝ�VvT�]!�3�
6
f��&y��.�qo�\�C���/�ގd'p�]c��+���k�����\���(#�˔�����e�ѕ���)�}~s#*_u&��3U/�>/Oǯ��X���>��@\ɝ�� o�o���uhg�p��ޤxW`���"ّ�h��(d=�p�`M�f�����jt�}��Y,,�!<0�..6��^[P�Q�4R�3�fD��<���bw�҇��KR	e���i�f�L��k2�����oQו:n뼌�3�(��* ���D��5��U�gN�?
L��'���&�h:�X�$_�W���Јd<�7w������gEA�L�7L'�9���<��4� �=�������ݭ��iD!��:���1wz�6�*O�#��d�ǧ��X$_�p)�z��\�	�{TC����4����K �80 62��U�rh��U�a��#������Mk�CU�j��"Վ�m.i��h�Sl* ��H�����?�����j��Ya6�~���[,����$o�yb��Z��@��ء?����l����t>T՟?U:^Pq�a�pB��i����ҵ=(�q`]i��ޝaq�U�����J��_A�N��iS��t��Н軒 ��AS'��>�}�X�g�_A��{*�K}������"�D�x69�F��i�k�L�x���d)& j$X�(��,M�k(�P�"�+Ed�U��辥LCV��
�O�'���4�`d��KK�n@:4�h+�b��uh;��x�{u�WI:u�҉��G�i����6*Ɔ[�W"Y�;t��h˹�&R5�-j�\b�7|ft�`�gq6�:!e�?��i[6�������W/s�}��n:V�ʖ�ܣ& Ҫ�����н���1���R
 -���������!�FF���O�(ԯr2�d0w��?qYr2n]~�t޾�g��;n�],�f�lD*q� ��P4Nimy��@�|u|O�?�����>=�[́!u�h�ql�N�=2��	���s5����g� �ҧ��}Hꫵ	�uٗ�P�M6�p��=�����J�YƯ9��V��Sa�SdG�5��H�w
�`��- ���n�|��i��^����LK=b���m-�-��<�6Y�3�}+�^������'厗��X8�t� *(��.,n��U�Ѹ�\Ȅ���q	�":�L8N:2��V��O��4����am�.c�	q8'��0>0;;+�n����s�=c�B	�մ]�a(0�VT�">K��a�z�vS!|�5ݱ}��eZ�(�U���od��bߡf��-��+��{�����w���N�p�%�T�t�%S?@d�� ���4Xq��Kl���u��G�	��ֆ6�N����ng�Qty���R���uK��?����n=���N��pQ���?��y͒ų�����w|�:J�N�=&徤���Ƿ�oHg9M�J�ǲ��p�9�{�~)r࿒��w3�����Q����h�N+����1�OaL�3�b�IA�L���~fe�!�[��+�L��DO���>92U�2I�x�&�_���H7�q�a�2V��H�68��RR�k���Y{��| j�+d����gc��E�{K�=��۷;��-��Nw�ō m�]j�!��^ʤ`���>6@�����##662ۜ�_���lY���Ƥ�w��!�S<�L���۾�D&p��[i7~����9��r�?�sٔ�����m����ú��鄅����Ӧ�jM�vFC��Ų����y4�v�e�������n�܅�=(F^Qx�� ���Q�\�m9���߼vP!�n��!XtU�<z��u�~�j�|�)��w���`�ǙV�geg`rk΂7�f]T&S���1*�DZ�E��uUQPۺ�>���)�Y�g�M*��V�
�J���r&^nBe�}����U��nI|q����"�3�4�����r`s����_���E�%]���3�d���8�3�`ƅbg��Ϗ1��y�$���I������qSl�� A� nO�����J_}xr���'e�d����9^n�_�X�Ң0����W�z�Y�4���~f/���1�=��A�Fs�I�I�?�c�H|���ńN[�1�{��������������h�F縍�D�4�RK��YK� �4�mݍEG��[��?�9�g���w�}N���j�I"��`':Ԧ��Ë�D9����������BZ7o�n�=$)�F}N�OV��#��ꑆ�N`�w���2L���g���ogZg��f�z���g2�jjG�^
�����'j��R�u�]U������`.'�%|SK�E�5�8X�����qi= �=���V�|<��.+�B�|Ò�p��Z	Ăޢ�3�Z����T�'#`%(�\ڟ��˱���Im��QQ0�"�~Mb����4	�q�B��^ol=��ؘ^��0gB��;��oI� `K�_}Ӭ���c�|���N�I~��H[	�`5��b�����<S����ZF��hWM���u�u6�\��p�>>�v��(1)�l���~�$�XA��@ߤ���<�#VS�ښ�A��������i��k��-���6�/i��L� U�&!]��y	ށ\�vY�l�'@��@ߘ�/��T$��|BV2>��v;�!�3��?�f-gL	��Q�#T��R��?\>Z��WP	P'�-J-0�#�
T��Z�J�`72;|n&�0�=L��yq`~�2�&Ae&��PT���=��q4�$+� tC��`"*!PP5̎�E���c���TRS�=\�+���ߓ=��lIz�����w^�6 Z%{�~�N
�-�&@XWy���-=-�}��I�Ӈ�&1R���<~h������t����U�dn!���ht�2�z3��z�r�m�Or���"n/d�=�l���To��aol )����֗�ڽ�N�������Y�T����V�&sH�L.ڕUd�5^32���"�&��A���Qk�U���>�~)	�&UDB��;&&|�Zb�m��s��`́S����(�8ek��f��=J[� �Ul��e�	��TH���Y��fnR����l���S�ܛ��kH�������Z{aPW(Lb%�y�� 2��L�X8�L�^I�	vK}/� G�vܞ=��D���v�0��^C.��es��h#8�߯P�����@�aҖ��[��[�QR57Mj����[>��Uq�ټ:��T;�����]�NkMt~Tm�c^ReDPm1i:ތ�k�R�$ـ�l_z��"�g�����ٚ͖#�:,n�Q隅8�r�{�t�s��ۓto��A����fh�������ק��a�����M�Eʬ��.ؽ5�7m�R��e�k���I6�{�2%u�Lv�q!�"�[4C�S���ܝd&M��/b.�m�pVg:�!\ʙH��6�9�a���6?2Ӟ��K�(��u���*FoJ�>�K���uv�`�Y��0��i���J��S�ڙ=j@c%Q��2�.M�.x'�ӉM���m�v*������;#�0��+j��������<�G��U/���u]���M3~Rw�����<��o�����!C�y�&���l���mI�Y
q�呭x�7UY�����ơ:�"x^�h��m#�q|�eu(Q|�p2���� H���I��}���,���5b���]@a� ����������p}z��Yf�� '�����:�4�C�P�p$Z�
=X��O��}��G�s�f2�Co��� �B��W����s�F�'�P��"��	�,H���M���G	�8��߭g���^v��u������ � N})�H+o7��!/޷���Q�ڌ�݄!_����?�o�[	i�M=�hZ(�ʫ��7���,E͔z�-��e����Cݵ�A`!2UK�\��хŖr���ǫu�����E'��vvY }1���3E���>;2���w��D5�Pg�nB� n<8Xu�20�@�-MBYC�WJ�h��e��ǋ�l�5�q%�0F~sCO� �f�14�,�6Σ�@�t��l]���AfL������l0��y��,U��g���ֶdc9oYW�2
�\�s��!��Vz5�$]S�X3�PJ�J�{�yJ1�ݟE�q��g; u��y��w������ȯ��"��n�*�����Nj?�xѐ<�@?��z9rS�;^��]L��l\�y_���矚	��mZB^����K�qR�M�\��}�	�z��} �
�]*'���e�΂�� �)�Ì�����ks��`��d\zýo�Y����n4����x�fٜ��A+�~Z�OpLjǙ�x��- QM�xO����]��ڣUk�3��{�Z�z0�~n�!b�m^{�t?�	|NL�q��Ԫ�cNɈ� �1�ɛR��`�[K
Rd�I�9�N<� ���K�\�Y�B�M�2�H�Q�Y�俛a��h�i����sj�F&0KPf�5�i�aLά�;E�ձ�U�r>P_?��J�
�m�D	_n-"��]8E=7ړ���`}���l_vΒ҃��(j�pƦT�`W�S�D	��eHfK��c�7�KGVP��̇U��j=��h}J6A���NI�Kby~�ՍPY~B0@��&��qeL��=�WK<��\h8�`����"b	���J몥q����#�s�U;�j��d��A���"h!*��$�y����{�oV�w�D(M��E\�I�v�P�ٻ�"� b\����	8+��/&U�,G?���3笭�d#<�	��(�L^���� Z��#���Xτ>�K�?��^	��Od��3�T���K��wO�MA�Ij�Yk��WH�G��
Z%{��S�
}�{ ]������!��:Oa�*�栟�u���z�GX<a��E��i�� %n̘�H�Ğ��k��� ��r�6�J���@p�z�I*�'eq��M��Y7SS��#����V..%�-������x�C�K����uL�%HK��P#�����EiE�(�F�W5�� ~Bپ��u� %	��B��ȵ��*F�z:'q�}��u���[�C�0}�-�@ ��=߃_�u@�c����j� 5aHn��]���oө�D�����s�VG����%���A�BUQ����q\�z��K�+"��<1dT���O��d���W<�J��	���΍?2��A+%y��ssA�Ƈ��y �M�e�l]+�/��3�m�W؇�l'����f��O���h�e>q�8t,E�7��8�	�H�C�5B3��������:��Gf� !s���@R�Î���{�{ح��fe�gm��'�!vx�Y�����Z˱p�}��'\vr�9�)�k�33�DVE�D�犗���%u5���kI2��A�J���з��$+wwdl��yV�>�'�hA���HO:�[�U��Dc���b;�g��l���ů���k)�RW�zt���e�["=�IT;��m7��aM7_�+�]6CiBa4:B�K_�8a���O�#���A7,v�I ��&
�1T�$�CV��f#*´�/�@\�,�
|��k���v	2��C� k����r{�J0P!�|�=DI��i���
�K�!��Td�t|�����D�R�m?&�)�w"?����Wj��6��R��Z��I��(��������b?FΑ�L�
l҄}�l�C�}��[q�8�<..5nt��
u=3�٨�y�*5�v�71��3���5z�tֵ���K�Ȋ}����������P�WT�-����;��]�s�>2A�� L�Tĉ��pux(С�_���_�c�O9�רt��1;�BR��p
iј�R�:_zT��_Q�;��/4���o���;�B��ٿ��OT(3@γ�.8UN$|V��M��J�ه�;��8_�����f[�!���|���*�n?���(�Jꢚ�Z�^g�� l��h�'$�P=��X| ��SV�x3�i��Sr��I<�	�X0���8}D_K�X���\��5�u��ѓ+��ȵ��;�TS�Aҫ�W��y(�~-��.� u#������B�v����2�+��AP~�R���F�kD�:l��&EY��ȸy��f'qw@9�8��b��;*H`�6O�����7�΃�֟���@��
��:k��L���F�V��z��#�G�чz�t��Njpf��u� q��ITw��rV���U����'iK���j2�g➱7�Ɍ*�FL��C��e�[z��:�c`�	��/�����@ר��6��K�b�9%�SF�F��,��߉j{6q�����,���a�Y��Z$������K<s+������޿���X�}����J������u�K-��I�z3!c$x`����t�q9O��-.�^�Wm{B�S?�K(M����@����=�74�x���6�#o@!s�̦�˴iw@�ʵ^50|fiZ�ן^1��6��mn� 1��O�w\��.m�[�>l�����G3KM����F�]�߾�v)S�[bփM���������.Y�1r��䞯sp~6~V^�6a���W�d�v�M!���t����x�d��|�F�
�~�C����@��ù����:�ِ��W���[
�3$�E���2�KY0��wi�WG1���	��P�w}��˪>�I������·e��~N�3�]��3b�A�Ω�|����@���c��^ojj�����'��C�I���^ۀ���A�8�7�ŢJ[�?���d���y�����4)F�u'8������֭����L��Q�����N�q�ez�iӈ�y��:g�����`�2'lw��D�׹�QvAK.�(���D�Z>i�\�@j˪�35
FF\t�ݱ.C�L��i�=�2���e�� �ͷl��t���q����H����)K�8'���y�����dA�pt;��Ul�H.��p�u�x�2��A�qIM�\
�&��8��[=���%L�ڜ<�������Ò�������κƐ�q��C[/Q�gqU�����n!�}%p�ݏ��8��u�d�&J�R�����$��Wc�9�~'$���,N��ԣZ�>J�8�@��0��g]����#W�-��TX�P�ЭN#��V�R�����i�&$?�D��+���������5����<�v\V�S,KjẶ��% ��0�9Փ�H�=K�HL؆PV�5��׌�M�S�@�E���,��nF����Z��d��:Ө�P�3Rughڗ��ZB���,ơ��@�S�e��1���7jY[;E��d<�ZT�z����5�����BdVt���=�>m]|U����m6K�ȭ��b�s�`kWI��M8]�X\�W-"��ǌ,�~ҽ�Z�^p� {���Gb@β�qa�آ��Dy�e��T��.�����u���@I�mtG��icG�D���Uw����Q1�R��_�V���+���� ?���1	pƦ�����e���q��K��I���z����Cݸz���r�������&j2E�1%n���,kU�9��w�} ��?��r�>2�f�&)�F�����՛{W��ơ�~�@`�9pX��K0�ZZc��j�?�#��R�ba3�)
�s�� ��Hr�.ETo3���I~>�1��d�c���V�9}�����2�4;j{Pl0��1�d����t|�}r�B]Q^���f���l0�l�{�i �.���|T��yG*b\9/мr�RC��wc�a�.��#w�3�C��9����$p.s�}q�����sQ.�
}�D��ʇ�%��.�/��\�}���)G�k����h6�S��m��igҭ��ke��l� K	IHm2Ln�p�v�q��>��~^����cT����4��(T�$�?eO�^-��lm�jQϐ���?P:��RK���'l�C�A�qH=��P��A;��}K���x���
7jԨ��Q�RD�O�J-�	6p��4�q�-w$W��X��L*6�Y9:�th�B����7�c�Ρj�h����g��>����,]*���|	q�@9�ė��^�Uw0��BK�\l��_�hX�n�o+J��'Ѹ�O[�Y�.l�,���<�p\�A۱�$�jtN��E�CDx�-��k%(��0$ ?�S�4[9Y����j���fWq���J$�8�ۏA��R�� ��^��^��hL�pb��Cw�K&'�����ǉ�dK�G2���C�Q�	n�����d���XXpW������!V[n�{����Z�IjB5{��p(�Z�UkO��Uͳz㺮���j�'�0>��<�Ng��4�ɜH%~�_��?������t��$�$�7ͨ��+4xغ����v(Cݮk	G{�vC�䧈��oMt
C����V^s��f��IE5q�ES�R�X�yڬ�}�Vۆ���̈p�,8����3�3�m��CFN�&U��H��]Q���L�eBfs�Z��p5��F�bx�{����X��ZD��+(�����A�Z	��$,X�;�j�2���jK7�n�?�5��c�|�O�[oN�Yl�z�u�<fccՌ�5��[��7�Y�=��rrW��I91�6��OA��2O!/�F�tw����}S1���hB��i�Dv��n�a���O�ӳ�����+�WlX�l�s�u�QN�8�׽��E��u�_3�1���H.#��C��x�Lp>d�"]�ոnwa2'�Ǧq�F���3���
�m���L��v�0ck-��jZ_�y�ѣP�
���*��u��=�q�ƎG������� l���K��:=���f䝳�\�B��Ԥ>���Z��r���zo��yB��Șя����))��q���6lE�q��m�^�$ύ��tf�ݦ�-9(5���q��"�p��I���zmx�XxŎ��DS�[�!���yq���E�J�t~ ��,lz�2��x�fӠJ��0������q{�
�R�e���Z�11��3�S�{�_�$Jی/�F$������	��,�d>+6 �;����:|�M|I+hv��I��W^A0Sƺ_�~�[�e�dM�|#��:|^l�|��g������6�D�L�����V�g)&"Q2 �S�̺d�@��og2������r�8>޳D4RT߉��j|���U�U�)!��uK������8�Bi.1�+��>0IV�g����a9�e�h4��>�wˏQ��*]�ӉS�ov)�R�h�M�M��]cˈ�u��9�n�AY>ʴ�T!�lT���F�VS�n��yx�ۦ�j��4�.�uI��'_���i����q��B�m�i�T?��D�����A�7�/���ծx����	̗'+�m��m?*5��v�[r�:@����/��F>Y���VRk�k5љ�gY_(A��=��1��6�د	'�tQбf�g*��K�$�X����	��s��ǿeO��w0 �k�ʿ�Ա�!wT���Tg&$�&iU~�nӳ���T;���O��&�)ϗP��
�6�Z�@ -*%W�.a*}b��_��bN'� e�\r9ev!��:��	�۫B-O�p���0P�k4��%���Q���[��[�ɏ�a�
��Nj��Bw�/����7��Z�0�,�gR�<D`�Kv_bh
z��/�I��H,]ʨ-�R�1�J�K=u�m��Tը�OɅB*yt%�.��/8�	�����ʹ��j��[�gr.|���Kf�6�GR��E��h�!�W�T�1�Xj���oֱ�r�rh�}ґ�Ԭ�7�rGPb�.��WFp��)3�0:������i�VL��9���?epj�^Os_5�<��Øh��z���r�w�V��UK=?��_V�9��B|4}�Q1d�ПY��mj�ʺ��x������oE�C���S~� �k�TG�-,��̴���/��{��ԛ]��ᎄ��X�wx�O���Yi\o��G��Ʋ�YT��ee(�&@��vh���U�4%�"�M"t{B�`.��}�Dn�{���7�#�����a����ӞL��,(|T�WO����mi��4��ƅ�J�)4_ۯ�c�|��?��Q��I���4L� �;4�����wu�"N��`�Q�#B��l�%��#�v(�,�<�}pz�'��7[�^����X{��jj�jC6�}�όO��^i4]�Wt �5�f����euZ��r�2Z���i�l>q�7J5�P�}���.����b.yw_�O�ފ	�I0��*�Wc�Z
"b5�r���7��ce��P
'�D�a��-Q��L��C������Г�G��\����mg�PS��)��2�;YZY� ���N�M{���&��F/;�0�9 �S���u}���r�9���de$�ԭ��5��xx���z{)�z�5���
.�Z�5V-�����Y��J�`'wp�	_L B��)�^��H0��6�Ճ+Ku`� O��sSQ�[�2� i��[H-�V9;[�y O��.1nRZfc�dS�޾���.�T�����3�>az��!����C�O��H����Q�K�?�u�B�l4���:W�Vw�� (�x(�����OF&�e]�ůk`� �|������J�߽�I�D��>���	�l�Ƽ!!bR)=a�j��0��uX4�3'�㈤�^��f�6|4�JP�r)�����f�)��s�kvI���LY�Np�_���>�炖C{{�ƹ�]�d����%��"��vm3��[�Z���*](=�����.�`[�I* ��q�)��{�F3��{��z�g�j:�(^�	m�`U�k�;6;F�m�y='�@1����6��"��I@[��a�#o��Ѻ��z]+c�a�ep��z]���]���COpUReq:�P��>�	����	O��T0gz���x�L��pY�/^Ǩ����#+��du���M�?��4�4.��"bw����}��i����V1��}������[̯�yv���Z	;�����0 �@
]��c��ɞqQ#7Ef�G��y�x�x48��k/MDm�ڜ�)�����P?� �8�D�e�v��B˪�˩�%^?��ˈ($��L�O=Y�-Ź�&�>�����
m�B��N��T�4V��'H�j1-Cΰy �kI�D��}����d� ǼaD���aO�1�-��b	�����@i.�\��a��M��א��Ä?�t\����l���L;mtg�^�S�eg4�>��Ft_jA	7?|���}O4WAU�%���)f@�9�
7g��f����'|�+�]B�U�穥�t�� Y�^G7v��g�`���%X�D�vO����&��$2 ��GM��*0��/����녒�&�d���x��׫_P�_-�` �����𪆘��Wy>�.�v��X�x���(���{��i�����̥���c�?�˕���9Xˢ+G�m�O
b�c��ȭ���0cG܏h�� �6"�UA3���S�֊�8���P_1� ����I`�a5����2Gg�=�##�j=�W1Ƨw&K>�!��Ϸp^du�!c5С�:�`og�W�6�ѿ�z��.�e ��.'���9�.c��{ۯ�kg�ڣ�-ֽ_��
�&M���7YxV����E�3Rf� �7W3�8�!�G� �<�ǫ@����>�`|�r!�8m^Pe�X�f)_%���vw�ŕ[{���_��ikF0��j_I��o��x��N���uG���Ϡ�ml�Pf���N	��NQِ�I֍F$���I�W�68���8��0��|_IY+�e�#�c��~��&��@��:�^\G�S�r;�R je�xF��d�aP�(kڞ�:>٤D0F���5���η4�����e�x*A;�Hc�f���f ���z\|X[��Ok�!ӓ��[�PN?ܧ�8M��ޛ{� �ڶK�'κWQ�ց�����0X(����%��՟	EU���N��8�4j&�<� 2�<�t��;+�b7�u�9S�������/܊s&gf����sw�E���i�KG���D�4�i_���5��I3�#?�����^���$Y��!2��!r��&҆��x� WG�<�I`x�T/QIm���r��7�Rʤ6yy7{��-<,�k�O�5Nj�;< �DƗH�	���\<Ss�:�����Z�j$�)O��.q����x�=�")�	��$�����3ǃu?�ɓ��n�'Ӡ��n�}�#ɳ]7����v-��>g��xmd$j��PA�&l��FN���2����U�A�G�t�,�s�Y�{��`ڇ��o�2�t=��	��u>X;���<�|:�h�5;E��-l��N��`�����T:vB��I�p�L���G�6޼SIyngV��.%�4��p�a��7��h�헫��V$�D��x� �[�Fۘ�D[wg=t�=Ǆ��|O�Uݏ!TL���vg��|AS�_Y	s�R']*�a���]�wD!*�9�:���t�akɝʱEqƃ�]��� `C<�E����\�S��B3�j��٭~7�y@歾�����%�x�elv|)�L�%<�\��r���������!/�,��e$�	�{ciPdҤ'�	�ؽh�떕�|^���7�C���9�1���2�X��|@��3���S��7�b�-*�wvO;�@w�n|�`����k�>���u�>aʳ}�~>�C�]��.'k��P��Mqr��JK�Yi^:�t�
t��^d-��Ž,�z�<#v�d��<�E�s�i�E����꩑9Xi��+�6S���m~���\��-��C�Jɖ�O$�w�@N���}��5��T��gқ��Fi@�?�i�7�%+������r��-���#6���uM|�}�&�c����\��&ҭ~�Z"`�e��2f����a�f�b ��G�u��c�o�<��h�]\����P����a&�Ԟ/���xo�Wٽ��҇9��ߪl6G�p'���<���naU���Qc�Z:[��cM6�)oL?���q�=.�
C��| %�@yd�x�h �:��
+r�ѳ��#p v#��K����,_�[vw.����bGHb��%��_O�)~G����Q�����/el�r���K�
>K�Q���A�\�@Xw������R�'�rX�.�[*��4ަ��8�6����u����VG�zd���}�#�i�`rGE�b�~'�����O�
�U�.U@�*!�f*�);p?��>���nU�u��z:{�8�\�y�Ԙ�L^��y�}e�@�lR�R��֯<v3�*��|�9��B6�h��!7w]I���o�3�����R�h�__/��=d��kj^�����02jЗ�$�*��~�b(�3}��6���n2w9�������|${���ZJ��K�����D�4���n�@j_|�u���'ؙ�a3?Fq�r��Y0^�F5�Yy.GI1��kM;z���v�0�kv����t�ő�iT�I�J�O�~��0�H�y+f�^�K��$,+)�\���R����vp��>ŀ$6�1X��,<��@j���ҡ��$ſ#�ciM��Ex�b+��󋩴H�8����f�e���N��t���M���3ߊh0(�4A��4�4xt��(i,Z��!�u�$ݏ�{�ͮ�Z.��_���#nBˣNsDs죵�:Y��x&n[ʟ�yy���K+y���]Uj���V7j�_�pOy���,�x������ �{>��%� {�+M��&����朔���c��1��RAt�T��8\Ȇ/���3'tn�@���L��Ŷ�w��2�Z.ѻа���W���(����(h0���~y�v�b��ΔM\c�z��&���V��,���v�7!����dsO��7��X��q0���
P$m1�>��]"�JzO��
�'Q�sm6��h�K�Zrg��tQ+�3�C����$3��V�q,�+_X���l�-�7<B��t�{��A/�f���t��f�<�B=%#��������s%�ǵI�u�ߔ;OvQA�z��XQ��Pf��_�}�i�f�Y WzJ(�=�*�Ew��D��*�@�G����1��Cj�_�"��o`��Z�;=�ҮσL��o��?6{��l�Ta�3u�7��pzQ��b-��M�dA���ҡ�n���z'��6,�%��.X-��q6Z$��j������v�љ���F�Jtٞ(_~['`�(����_Y���c�+	x�g��
v!����n� v���d�>�Ez���}�=�����u�|��G�|$��
��=����ŧSO�U���7i�5���N�$+�
ԗ�V-C��X6bcg���YT��u�T��@�<�
zC�Q�]!,ck�b��ұI���b���?�����n� ކ��)>|H�n��0���Q��ar�$�*�?���B�n���+_�� 
j��|~�6��'���S��f˞�(w�����]��C4��C�S�G��p�9"=A����㓉~2hϼ���������*�$��0��k�4�R?Ab����ZU�J�߻�=���z!
hi��;p
朢Ui����I(i�L�pFyBFs�1�8�4��-.�'�j����|x������~��܄�g�6���u���������	5%�͞�H��Y�6d����֬N�d� kԳ{�";�ǐ=�����}���hKĈ�e��h��.�D6�oP�?��W�ߏ���elC��:�ch�����D����
�P]��AvQh���h�4 a�S���K���QD��B�ƊL<,��ٺ$�A�d���u󢴅'0O��^������D��k�6ܢrFj`Љ����o&Ś�lP���� �-1;�������R��%���ښ҆ ��gk���&u�tj���x�*B����xk*���R���M^�cҕ�b}�9`\��.�ύ�Q����\4V�DZ��l^q����[�&�s���=��1�\��Vti�;i"fm��a �53�<�62i.��p
�=�߲N�&25�y �2g��qo�O��v�=�L��U��q-��vO��A�7_F�%�����j���nq ��lj��[N�<&N��3�����s�!���v�{�qӑ���n�Lн-_����)l_�k�\����{�-�2�L�m�'7.��������I�r�+��Fڝ�p"���)�*�۞s���:_*����54�r7k��ۇی�<5z�����J����9��!<�+�Y!�\zE?:C�����M�Q'��s��&�%XO����q��}˟��QU�]�r]�N(4F���mk���>�I�������kr�Sy F�qBAC���Ƹ��**�_3Y�·���;,=�����X��j���L41'|A�Y+!K�Yx����S�ʸ8�A2�'��&��Fm��C�Ep�]-��lo5>������Ŵوa����T@s�����i�)K���w]�-�L�N@��E]�W�)�W9���d� ��'������qVĕ��1�L-88=��>��.��o_���SL�6
�+�2;���kY�qtǲ��Κ���4b�����,S�n9�c<B����5_ꪞ4�A�6Lss)^k�����O�8���(��㤉^�ߔ%D�5v�B�����g+��3t��X�N���˂u��	�̈� �^�a!1q��ԍR���Ы��E��|����{W��5)�~��8��Xa�X���@��~�q"nHaa �q0�@�i��Աi�Ѳ�pW!��)$��CX�<ģF� p��+����:��9��~��`]SO��ɰ]�acYO%�4,��
����|=5�k螖WE����j��ܭ֦�Qy�nB�"K�@�b��Q�;���V�932�`I���}����+��[v�Z�}8N�����nt�8v�T�"�FT�<gSG����7��NO�P_�Np��A�e�8���֤Ԅ��{d�F!��nP��AY���VFMmz?/"+�~M&,<nDWZԬ�r�p���&%%4t�,K���p՘h�G�sI�x���!�\n�c&p*`C�$eY��O�W !��L�M������Z,LK�.����p����R�X�EL�U�*�j�z�o��ۿ	�H��z�R�!M�x>Pm�f. %�i�Qh�~�-��Ah|�'���ʲ��jr���s�Ayȣt�9��B��U��2�(����w�$�i����Թ�d�Ɔ�-�k�����!T�
r�K�ye�D&qn�ؖ�?��~Eg�H.+L�����T���.&Րӕ����;7���ѕ��I!'W�KR���IIi OI�t~'|��lwuB� 1����� H�<O�^S����Err���/+	:m���4�����Y9���z��=�쏌����#�3�/G7Uf�6!�J �|��hɉ1fKny�n���ڸߧ6�An&����w�����c ��iek%M���O�jl�M�D�!'��k�y�� J�y�q8}�}�{v)~3���>)UaS � /�a�ݥ�sE���0��Mq7�^��=/i
��['4r�S�ﮧ�6�M�U@����m_�	�e�*#O��U�|0�� ��X�e��	"p��B*�T0V�D�6ڒ�@Na��菼���e�Qb!�~}^_!���R�?G�TY�i�/Q��v�V�$�������;~�oy�MN�/���$�_�����{J����_c7Q�
�I'�i�9xGz��3i�%r����{V~ͼ�qr`� ӧcs����8&��@C<�v|�-j�5t��k�	��ܸPM��[�܂F{"��Ȝ��wYײ��EM$/H<+>NƄ��6s� ���z�,s�e�������Ai��ȑ�u�.�G6[\Q.vW)i�ڏD����-����#Y�[�����G��U���3e�@�${�\��ߖ�y(�vBbI���!�uws��:�ι�����d�`8�:h对�g݅V2�1JY��)^Y�N�i��7��u���[HI�7��m}�X �J"�y��Аm�'��6�2���;����
M��~61\U�C�/��A�t��x"4! >�/��r�˧Y�^.�W��Aф_�;��Q��� ��i���0�M���$�'��PBe|����½�lk�N`^�[t���c �� /
�~6Gq���%�4���6�N�X�Vv@�Ky��
�|�B�^���g#T���IZw�1��Q�sZ�.�� ����R�iՌ�8Η)���,�h�.'=x9x�"������D�>�<��h�@٫����Yɥa+��t��{���>N����i`��͹��23RRa�=��וt!��=L@9 yH"8�=�5�zЁ��-�Lͯ]���N�s���i��&�[���A���4+10��Cn=u+��1WT���V���3k-FG�C�,�䍚��NK��A��A�d����]�0���Z ����w�7n����R$d������Gs3b�7&I��_LuKv3��,5S$d7�^��j��F0��彾�l�߁~GB�������i"���H���1��<3����N\J�&��;#���v�X�Y{���r�#�+-K�Yt`�����Sc�ߕ��S�<��Ok�d۸��̼{nQ��M�R�)�|T���[=��Uq/?`Y *��m,n^��fd�˥1Q��"Q��iU�J��-�Uoz�C"����R�_;�C[�� � ���X�K���xmJœU�ϫ!Y����\�Z��tG�Yϐz���.���Ex;S-�+A�+�`w�[�4DD阩�±�]��gGhu"`h����$ۺw�戤�5z��R/X`�������U�6G�
�x���wluO�~�.X����?F2v�ء�~�]�{Z9��˿ @6�b��K�IqL���BEy3��qHz>RN'�i�v퇺#k�(G�I����(	tז���9��*�?V`���S�����Cch��E{�	�F-�X��L�5O=��΢Z���֛u��	�h����:�����Z���� 8#d�����_��h�ۉ[�q����Y��J-86\���� 6�>%�e�d:K���2��������F�EC;��5�zD�ƍ��E����M��:ud��  ��1Q��m~"Y,`�f��0C��#�H��������]Կ�ʿ	�]ߜ�+d0��X�9�65�s%nD{������e��Y� qE�
�e𬺈lY`�����4�b��M;[��7�SZ\~�R��]p������њ�_y����b��V��gN��Dh�#m/Sag#" Ӱ�E��9G���`����<l(��N�G���]U�8�9�p�Z5 \���o��K�����	֚��Y~=�+�E��C�$c��5ڄ�l�`X0��s2���H[p�ZF^*�l��1���Н����s���/K{�P���o��1��߱AzOwCv/���;��9�$�'�8WHX����j�= ��	�?��ҡ�ƺ�oV����s�t(��([�����s�j;0�6�5�|<��Ǹ���sxJf���E��+����)�?���a��XgH4C���z�>t0��.5���p |!C��ƂY�7V��L���w[�Rٟ�]�����A>���!=����� ��w����D%0�h�C�i��Q�����#��Cx��O�8��uϟ'�H���s�r!��.�gi$R�BW���Fjbb�U#��#�V�h���i�ܳq4��$����w����S(�Bl���R� 1���׽��s�c����ax����c���:��&��o0�W� q$%m�_},G&.SV�8h�~%���.��SA��e��r�t&Xj�da����Ż	oF�Qℝ�� !�����w�g�d��+�|�W U'W��T��e�ݦ�Y�As~�Q1�9C�L�<_8q��}�pm>�&��/�F12�*�`VEsWC� ��'��EF}}��q�6���-`�qLB��m���e�~�=gy�����!t+⾟���48��e��?�����	��ўe�}�4����\Ǎ��
��vpW6�E�
��2}�:�.�|���@&�Y8�Ч��1��θ	�(����\��|	ɭkZ����fj��X���7�u��K�\����pÍޫc�v��v��F�
Z�?�^�Ip3����`�����ؿ>.9ҥ�'�I�u�E���8s��S:-&���G�x������GQM�]�����(F����&K���K�25e��]�V�`����׭c{�����a���I{s9Q��j�b�<�����օ��4H����Y��0�>"�j$=ֱ�8+ugzU�;����*|������s�Z�`�۱�5dO~����|�(���M�J��{�?:ۮ�V�R
f�S\��q_��Q�?��y���d>���4{`�h|�X��A�1m���+?�pD:�a-k�{����C�g W�\Yq�X���)ԑ�[���z�v�C"I*�~_y��LE����d��V(���ia�#71)�Æ��h\��8�Б�g�2�-��L"��eZu����A�&�}H�u��h�F���+��wZ��^�%�~g������I��P;'N2J���U�Il�1'�8�\Bb��Ô�C��BӤ�A{�c;���&�g!
�=�1vu`c�C(�.��4�Hp�sXQ �0�s�6վޮ�c�G��n�R#5��gqfl�H�K���C���@�p�+��Q���=9Q��
�v|�i/�C�E�V�\rږ0���F�t�����>��{n���i��w�.���ޜȯ�m[F G&7T�!8z[�����Xxz�o\��	�8�#5��?�8�a��q8�~"6i}� ؉��\���Z?�?/��n�����ǱQ����UM�Όtd��[�|W*J�gr���X�����|8�D�x����ܢ��XD9����Fx몍�,�ư1#�� 7f�ؾ�1�V2A�S		�2�]l���&\*����'o��xC��$ K9��"�p�<=S�Iy� ���EQ&�;,�ȉ��m��d�Z���bEGB@>x�H�u�nEw���� :�D�s��$�NÒw�BѺ}�f�c��Aw=KF�7��"KN�D��?9��r���Y��	�6�����3ϒ�� .��
���5���{��O�h�w) �"ݽu��H]���C	ρ���U�4L8�H� v�e��T�&�;����i��O{� ǟC;A<��{�y��7���%� E}PUC7�=���RPф����K�ҕ�J|&��m�OL�#�$�{�̉�ʕ��܉�<��-��!8����j����M��;B�9W;�m-T�Q�������r�׹�������J	�OnL��q�B�ba�"�5��]�����Z{?׮�3�v�c��TV�+C>�놭�� ���p�R]0��$J
d��6��}����Z|�c�t��:��k7����^]M6`�3�W������y���V���}h��(�?)� ����p،�Gt7����������^i(�jX�N՛d����5��V�ˬK�Bq����C/ߥ �.쥧�����N5ki��P�V��E���	�#J�M/��:*�Ç[�wѣ�e�aǤ���������G�­Mt�I�Z�g�KGXć?ݥ䔎�0D6�y��J��O� ��8d��2k���Ś	��	�X}וjs[�7�I:kakPPe�M�L���g�,�@�$��NE0_��Y:vy��4�G���_l��!���t\ ;3Q�S�<7���.��-q��U*%_m��#��í�	 )�S< ��&
�MB*��H[[b��5���:�S�M'/�j���*�{�\k8�i���
y[j]��s��>%^�M���y��A�1�6���_
.�(�&���Ժ��3zO�<`�sѼ���$S�}��_׃:S�I�"̨Fs!���9��޲Gw�)���Dǫ�h2!�ϭ^�M��9kJX�J����P����y�����9�J������[FE�C}�~�Z'?u�}�p��.���؅����K�~�*���##�-�[Q����X��Z��V��2�Z�%�9��F�y���wd����{σ$�lL�5]�ol��rxTx����[5:O�4e��N�l\��Se1P�N'���otl v��-Sf!B�K�p�Y�b�҄�PYTJ|�� �E�?������r�VS��:�"e�Aɖ�{�rp81��``r��[��+��}�1��ݚ��+~�m 7�sġO��$T�]_Cz>�C��}�T�k70Q�!�I�PAB��h�u'�ߋj8���g��F�Xaf��B3t#�נ�G�4P@��Su|!�˝��@��4>a���k2-�ʝ*�G]��򰟽��?��r\���-_u�L[P�˫�a���p��IȹE"[���y��K1Xf_����4Ls���b�y��r�d�)�c�? F�C��������o�V̎Ak���S��'p#H�[7-E	��>U��){�>u�������H�ذ8�~��m�K�}l(��Cƀ�~���3��}�L�h�`�_{���ʉ�q���ޓ�3�����H�ʱyH@LtWB&�1u�S��R.bs�q����7�"W��P�����vEr��f�J�0�JS�BƱ$լ�������/p�ᄗ��Q�e�3��U�lrDfiۅ_vaJ�~�U�dPV�B����d^P/���FU�b�cs3�W���W)-��i�Y#�~%V��GŤ����QI�ʢq����d���KyE�&j��+a��UBin����)�b�=�x�<�C0�L��Wd`��C�=��{�,M~�S�����l��#]>�l�[�;�a�C���������c�i�;�O�wv�>�6W����o� ������r4�C�����M��U0��rS��U@��d|>p����J�&f|R3ૠ�d��ͅ;?���"R�,=�>
9{~�����[��(��k��z�)8�m��R�I�hڑłk�3QJF�	k��2#�î҃j�	v;ϑ���Jzh�O�c�JJ�d��w���d���]�\cf�E/���H_Y7���޵M%ng�[LT�tT�:m������b�i���f�C^a̷Ma>@�6�N^����ep�Pz2�/�<�1?�Y�$�=�1�ISND��˩�ާ���Wn;ik���,[]���7�u��%8�^߽���܌F�\F�2�x���s�+x��E�����$�w��֐g�鶗=�w%����wxX���KG5jd8�h��^�g@�������Dut�U��0�</�&7r�k���GqbBZ��?H�-$49D)�z�n�[ܬ�<�Hc�}B�x��ƃ*�fk�U\��K'}*�ٴo�$�)�������� �����Ч~��=�Qxwuvt4�|��=�=�C|
?�0F=����Ĝ��\���I��<�-&@�,J�@��Jtѥ�����<�w��͏��ϲ��K�9hmf�q˸�����na��-=A�FrD��"62�����ZЮ;:_�s�5~�
j������f�	h���Y�>�К����C/�Ra� �����ȭ+g���,��e�63D�)���>�oQ�D�t�_��'n�z��d��f���Kt$c��PQ��Y(M�x�W8����p��Q�񊵠o���'�DՆ�Il��vߊ����vȸ�z�?d�m� g�؅}fwj8O�er�̔V0]��wf��o�(`�ȲȈx�t���Z�R-��6S^U��|����s�Y����-�<n�t좫�Ib�S�-�2�}�i�܌I�������J��q6����唞�!_����z$'1_.bA�(�%b��Sg��`�~�b��4����k�]���lXGa�ē�L����S�H�:6����
�ݛ��?s�")d�Shm7(T�����c/;c���LN۰��3�I���,� DF��1{�:D��0��off����*;u�f�
�@ʾ�=_tN9�c}�����`}4p����`�nt�(*��d��<���*$8Z48퓁io�o���`OyV�(S���T�����";��w�H��`"���V߼邌�&t�P��KM cȷ����n?��w�"5����}��G�-���RL������ƓG���6�$þu;n���]ńv1�
�^a�ʎ�AX������/߇���2�����Q�jW��D(�X!c%B��y����c�p�Z��Q��3?Q(�,�-����ޠQFLH:����ݠK�or�.A�:�z��v���X�\O��%Q��9^ѻ��OlG��YI�������j@�ڜ����ڬp��/�Q��P�ķ���=��`�a��hf/��9����pc�I��9@��z gZج_��ҿ�ܢ�e6�up�����W��;��Bb�:�;t)H�M��S'-i�J��O�(�c%^��I��2ϝz/Dց��in�~�da�bQ�b)�b��k@�n���&�t�#�д�5�a�풕��[V��+�V���]z������g����������qTo��0Q]��^�5����O���OF��^�k]��#;�ة0��;��;( �S��|Щ��0��G;� ��sx�9y������ߤ�A�z��r�>3�&���� ��O��re�i��{���|��!$؏m����D	���~��?z�;[��U��3^#���SS��"���>����������w�V'��=͐3�y��I�0]oU�5��٠�T�Yi���T�� ��_Hi����7 �t���<POn�+�<�R?��C&���%����_�kw��=\W��$y�w.j�ud��/�-$# Uy1��D��S  kʼ=��
�������o�zN��6�l����p�F�*H��֨_x?���e����FrI���ݽ�2��z���o�J��m/�k�O%��絕�bD�_�lB �F�;, �����w71��pc�����r���)��y��=p���(�c���i��!�U�zW��������T�@�&�=�	E��Y咯e�8
ɭ�I���r���-�4��[ﭵݬy����t�����#�(sI�:��HZ1�b�:�H��0�JQ u�i���S�����}��Hm�5ty1P	xg�+�W]��A���Q�+�}�����4���/a�Va��(�6�`� :�_�&(z�s� 0s!�d � D�t�����xOc��5�YR�<�7�[̊f
��~�4نܲ��^4)m:�vHп^�X�)m���H�Џ}X,�.��WW�8���h����Z�;���4ve-�(n~��<�_�{9X���$LW>����6�z{��b�����`�y�ڜ@�ɺr�׺M���1��@c7�TX�(�8�L24�<�I�~�D�$ե|�s]2�]f�xmp��r������S�$
��U�vv�	TSI&��!b V�%o��(�G�V�� �����	e��^��O`�����9j�@֭�� k��Ё �X�p�`���9S��������/� ��#�D��sP.���TD�(�ZSfV�K��N�"<�����X���\�B�p_�Y&��㶸����3ӁEj����Mc�TG��{
�6vh��G������O�6C��ld�o�q����j�`�n�^)��IQ��S��T�y�hW9%��JQ�x�
��d1�����nj{b���.kH�
�қ��j*Ƣ) n���ͫH��˹�G�o��]��;�<��ZD��r�	7���0���,��G�yv�Н'Ғ�`u�ѧoZ�N��)��&��(Rs�S<��mՌ?%a��κxak�C�6�d{���yOį�^,~�����)#c��P b|�9p��h�j�x��Ԗ%e�$�۶Z��gNp�,�:VI�Ci��\{�ݡ-\�Z�M���O3��&򖰦|-��tz�%~�zK@�Q���7�9}���^ �����Y���y����2���ED�)�g�:&�mMnJ�ŋ�HmTG,�z�k_�m�UQZ���ϟ�n{��i��{�J�rgM'wd�H��}V$��r����A<�����,z���_���Q~UP�J�x��j���ö������P.L��$�]�JÕeO=@Of��?�,�޴.C"4{�[�l�K�#����H �@PS�$���#h }�2|���#��p_f���8u�5��v�w^l���jV��c5�Ԍ���)���Q��[�E��-�_>�G}��cN����F�=��Ҝ,���m�R9]P=@B�3>@�_�#��j eEdS�"�h|���,l�͂�P��:�~���;@��}��7���
[��>��
��"�n��� ����'bY��x�iڕ�z�"E�3K�1�X(���^�f�x�.��k�-gwb��J}�^��t�i�/P�R�a^HS���Q�y+���Ѩ)os�p&�,��Ne}fF~nB�s
�0�Z��k�x�h��\�����mt���K7cMC�����	��ӄ���Ř�����1��$U26��xlY��Ҹ��v2B_4��D�"�	 Eb^�ב�4(a��[���X�d:�Ǩ�6��9�^{����v�+�W9|��]\պ ���?��X�K����Lv�Xz�X,�x���^�7�N��%j��{��x��=7M�!�ߘ�[�>�#��FK��"�H���(���,�wuT̈r���?�/#XBS��u�ҭ4�	�A�^o�TK��FݵcG��y���ƜI�$Y�b6�f����!���U�fֲ�Yv�:`�O�M���D�v4 ���@��=�8�v���� �wc�ƃ��W݇�p��";g���՘4�[�L����*�����X�pYAQ=4�A��[�9%D2����xZ;3�EZ�dH����vwDR��9@嶮�ky5�ۜª���֪�L#�@.I
P�B�&�":����=��M8���P����B(�;ކ���ܛy�e����v��|L�1ė��-5�3(��ݚ�4�J�]���A���j��o~�;}[w�%-�^3�>fO���uuֺt#~�sQ�]�x�_��{uY\�Sa�|[�r�N�2¬b|�9+lT��N��Ƕ]D\�O�3΃q���My�����k�๵s�w=���`��C�7#������)/� �hKΏ��b��W�En-̋�\jHe{Pt�>�e����ȹ+�r���Q��Ä�s��6��Dį�3�*=sǧ�����8�9��p�p!��96��?Z�1�G�c �G8���g���3�V�'�f	+���\�p~
B9iǟ�:�=����)�c�>*�`Z���{�b^T���Q�6*��5���\{���c�ʰ��J�����շZh��CA��r����x��t�?�h�H���W-��F�l�ی/�#�������$�9��y�nM��A%����?.�!���r�#_%@�etr�Y����e_
~��@�W��Y�I*��O�+4�
j����$�:{�v�_u���)�i`WkFW�}p!z�-�7 �)�{A�[FL8��:��*T���p(y�}�5�3�m+8}s�T��]�fNI��X_c� �D#��
I]�^ux ���:?�X]φ��@bl���Xػ�!p��ok2z5b	"Y�*��uE�Q<�!��7�5 ���(�eo���"�;�y�'����&�)cA���݄�!֚q�� .[:MjI��F����C�w������)�GA� ��l�yd��9�ħ�R/q6Gko�}m���T��I������F�4P/ӌ23 �I�Xl��̌���|�kN���F'��_R��`��`��:�!Mݗ	7���ǁ !�y)?�
2�'�v�c�[m�N%�$��Q���%@KH��x�R�F�� ��ʗ&����t$�<���4�˯W�3�$��c���T�z��ۥ��5��F�p;`�g����ǽX�h���b�%7� L��=����x�o�my�[i�«�4��}-��3Pt 2,�%���+�/�����6d�QNY ��l�j��Px!�o-xa� ��㲤��\�!}OO�� �Q�n�(��u,�F�IS�ӞG������&�a��A���J'0�5zN���@�¦w�����Y��;�����Wn��6�;j��y�e�`r{(����^?`.����p��cb��;�訽3�'!%k�v�AQ)�=ʴ���#o0ppr�p����$�����=��Qo���e{~P�Ҡ�Qd�yz0)��G�u+�4�o�}�p��E(g����Rn$��F#~�<���WM�]>��0R��@Me?,��O���QJ�@��ä����:��8����t�"��z��^��c�)`�������Ѽ��fETB(o%�7�CO���⩲�f���ù� �U#1�!!(�5y��W�{C�x��드B�p�����*�5��>��_���C���#��p������i
���Қ�!s�K�����2��C^uQ��՚B/N��i��`�P1�P���,@֑�q�G��"�D7Ҡv5���ǰh�4�'%��2�R�w�t�-5w��f1o����c����^��C�4�V��7���#i�|�K���iV���EpZڳ��Agn�7�\�f�b#ZC�K	p�P���G#T�y�2o�8�����g�;�ao=�q�`J3�%��bؽh�A��*ٱ/�N��� Z�����ں�be �C��k*�{apO`[�c\���Yg8�"E�#��էet���^Esz�@<GkDi���E���U��Ո��fc�qt:HU��e���=�LS/c�t%��=tp7j+a�<d8'%�/y渣�Wr@�Ӏ����S�f}1�����6���5͆9���Xk3��Ÿ�yE
Zs��&��{�v!O��-G,0<�^w�R�}bW�Coɧ2{��(�^��ߥ�{��0�N,]�����jU�"�y��ڑ��}�K�AOj��:���D�%��^���9�b� n;�@d�_]QeR��CM��u��Zk�M��os2?�Y@�i���쏦�[��P� ����]���'F=ãu�h��1��2Z$���(iN� ����5"<y�R�@��U��q�u:0�E��z���S ԙ�a��x�	 ?P#@�ʗQh,�Cq�/ST!�G�㲴t�G.�X*J"��2?�@F�%,띚�%��r�?왉t � ���R�����N�I��U7U/�Ʋ� �d������Բ>�ʼ ��u����#�v�vX���9m0�%���׻�KI�$��N4a��%{99nJ?PfDn1�l#��.od79�_��+V�OG`��p��u2�@4%*��O��"�VŊD�v]^9MB�Q�]>���h�7
�����Su��x�X��t��i:>,1�!ל0͞�5���&���kX�N{�����kz�~g�p����٭^O�g�tO��n�MՇ��t-	 �@���,%�H
1参�1����	�������K��]�MM��}D��Z��í���1R{]S��f�ӧ�g���ڰ$[��o������\l
���<S%�	^�Lг�J�QC�2��ªu�=F}4t�j:���pv���F�E;8#�:��o���,�����*���/Cּ7�6➧�Uk�M�y
|RqW%"�[R!���M��j0}�Ç�S�d@�H��? ,���[Cc���?S��/���`�ˏ\��B�І���iy([K������񟏡��zd�<B�H�,�V,�R���)]AQ_�u�P�yOX����Y�{�qpN~��o|�Õxь>�ICӚ�����]��5]u�,w
��Y���hW����SA��ͮ�ȭЅ=\��Bu=D<�7��(�� k5B�n-8�2�h��؎�=����U)M��ƒ8�ӯu�u����:Š�̻�����=�&:F1�s�%�cQ����qZQ���������_Fyc�Ո��s��cB�M7�j"$F��Lks	RW��U6��j^�(��p1��o�V�]��ՃEv�HK&�,?�_L+���{��2ȼ�c3��S���XCf�g��d.��r���w(|g���ntlz
i�c��$��n	ϝ-�Fn�� �� w5�<=�ͣO��T^��Y�ݍf\�b�e����������&��
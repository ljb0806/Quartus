-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0dFk2RVGHUcUEyYRYB8bEARNO9m2pzyMB1OBwFnBhjz5rOxJ0yR0iKddyWM7JzBSl+Komj3idNkz
xByu6A0NlAytgGFQOWocoWVKouP3/Sw4pikIGP47ssndn/6bm5n/KnB11uOYjiFvcPaWY0UVOf4c
ChHoVGSGu3Y4YakaHSbLTw6ozDe9NkTJJQLjQLvM6RXQeCZVUl95MiUjJa6i+uTbOWX+0c0GLIJ/
7zmcoqYtkOQNMo+nEl8YJ290iJfOiBuubCIrz1cnL00DIHPLB1E4UvXAwrqX/MHOauTlxQ0Xq3Gh
Lwkz0jpufU0aXN6NUw2Zzwwn5h4N4MUlzhHX1Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 82048)
`protect data_block
uConoUkVVN/rpPrZ7CqF3av5/oCIvpVXHrebkcRHkMa8MgYjBtzG9mc9PdgOS9vA4iXxsPUBDXZ0
NcP2U6fNSqpqYHrTY4LXeK3B5HJ2GSANoqZDNVtTI1R+5Le+tMGIpibSU6oHqRRJSqItp1AcgAAn
FTYEzpw172QaadN6ZkeRFg9GF+pV7/PU49jaq+Bu8M5z2YfozE8B/+h1d1IA9Pau0pfPbM+Hr3of
OEzY+rlPpINMYOq/RwonB1BJFcc9HPGpcyhvdOfs2wT6XRXgujqjNMawBXolh1VwgnPIsMz862lo
1jjdTBJMAWO+VV0yygoqV1ppFZh05LkAbXB30VBAn9qri5QvL+GCuznTirS3y7a8aHjI+eh67B9p
qmoDbLGjSe98TYcZSJEsXFhVYI2xsF9dnHv+BJVf+dOBszbKV0ynva3VYx83/Apu8dwBH+WpvAed
yxvRvJPgVPwDkMZip3kdp+ksMHBBsS6+yGAUe+x1coHAQh7Zzl4hggUGiRaat4QSWowpK+PrHLLg
O5Rez//S9riS1vE0Ov7cbngxAj4OSpFW+5wb1rQMd5AAMDfcNvEnV5ksFwP5dI6s7qZuGkZeSkIU
4ipTISJEletvPcRK5LCic/2gyLvV7vBuTtEzMXwiWl25GBVwvWRmY7DQQ2lRYhu9o5ymNhSoWjtt
gtSRn8P3Z5V8LRQTJRYgYLlpIq1MvYDiL2bDiVmUI2Y2H74q7H3kk56tbcQQln7iowuepOfD3CtI
vGlfdBqZwTdwjCjgpwdSJJTPxYikKiMZ/btHCYKWu2Kn8LbLzsjAfE00Q9bmMWqvicm56moQ1qkh
5czaUByFl/+you51RdaMlXjvEaxMtUO8pPrGUQrYAMl0epYp6YXmbhGsXlztONwpDEvbKp+3FD6w
4W8sk5BSrl/YsGsxi2M9Wn9vcTa0TYGKbJGU85mbXM9rIvvj/BelGu7wVB3S04YgJp9MS5+3+Ylt
4rQi2kW843YwjtJkrQR1yLSxEAftaWlnJNM5cQd8X4ls+W5+tqDVvNgmwmWEIZvhHuBzfr2zT96U
mU9ekH5z8DofSObhDgitz8GhPIvFnwarnWGbfIBleq18j7u1S6mrfAD1v9T+C1OgfhcoKS83tYuD
jnxiqzzxQ5whvX4odblngUdpgBqWTG0FdWHgAj+zTaw9lWq30FZEmCvm6ixm5vsfe6VH4GysCvVJ
OSrq9Wxvr4OI1/3U8eATK2JGzzp1ziwXhG9pzrGr24CZK4Ih403trBT4ipwXvQkA5iFFtIixpQXE
6C0REzi9klPLCcD1DjpSl8j8UUa/8aeHLs7iuToDeKfxSafjUX8CC+EUMrKfeGXJZTOrCQDNxdbw
44OP7eEFyaINV0Z5SxbhTFGMHwTLHVxVBEkzdsW8SP96kLSs4LyQ3DH2xdHP/DCL2N8aj/GrYlMi
0/qLrsuigVo2EdueLSP0dJjDV+G63yUyYA8gIhS64oVu6DwL3HjgGNTACLZRx1AL0b/GrzgwLVYX
85zMB974lpTsEVsXYCKSOMbDreUtbVIuL+JAeYYcLfR2/EE0SqIONx79v78FVrVvtpb512qH6ogD
EeKXNXhKMmJZi4AOkVqrW6MRnsbg4qJr3wpNh+zqECgWABL9MlkU2pwE1bLdAiU3d4ARSjsGk6CI
qytDR6+s+MK3P1lKLMgI6e/0fD7ImfJFrTc9vWfmpTEwFWERStejUlHJO1wjpdE5rEHGXLJG+WWW
xayHp8IOtEhOIpoZ7WM8X5B3jhuYRSdUvgpXtOWXJxwOt/QCQ4EA+g7VYvN3LjIGgykD3YKQn8QV
EykN3ht35A7TTSwqfsHHTCAqpELiFHTBVDs2W1Yl3VNyk74XCXR7DUjGgW/gvvcT5XOplmlE6kD4
08aC3ktuaKFHOj7HYNYpCsJDRwRkN5jM4IzCmNubn1AdILcsIxGYSrqrMGx/kKAPMHDfzJDkiLia
WmfgTDz294w/KXu4GFIUb8RlIXxql2jNWTLE1h82rMUqn3nGRrpA2CsyXk6Jt1AUydR4WPsSfAM0
QWKwwPbOImwKz+AFRfxDb59qpFOC6TZCoYz2jZVJXo0vZkg8763oQzfQ8ORdFvZwLOhfnkIUVTgQ
UaeH5kTovqVk2GGKPIfMSSBFmIlMFKyLM2ifPD2KpRTTZkRBY/6E2yb0ypS7uAe4xhUBnoUZTTkh
3h9Ncl7/RD+zVg9+r/ft+7u/xZWINExCwQRbuDekZ9lSg8dRVcPOp/e4ooM8jqBroNCQpcvx6XFT
ZmtpA9zpbfxT8oxaZ590ZbMvb/vajoeylE+EphyB4KQR5iZtxJDmkfjmcCIp6DT/60wWYB9fE4UJ
mV9y7NROmLYJ0nTXrFoibekA7OIzzZA+E4x5IpCcpyOT9sifl8gc5GKXIU7Tv4tAcLIBwtFG3nXZ
59TdeYHwMKIcwWlxmU+IxpLNIYSLEiorJZ7LsxvxJ112YjFkINEZA8v6/e7A1ekdZtx9l3Q4s+/T
kJxJrE/gBDj203Of9i+7+gsm3snrd2AjOOYczo9LZG3o1KkTEQUaVq1PGAgL2mLpZxuqU3tc7lam
1EPeXNY2A81Sw22BMiOw05ChTEiFGZdL7wYgohx5WnZqOLzvO3rXIIh3f9yCbC+0fre5FGYRgZM6
yi41Mi1VcQn8IJWBfpO7QMW8asIvpbCGxS9GsEQuxSbJdmBRRNTCoK2rS9b6uS3qTnd2yhsnYrv+
i7yUp0fiuWPQmuQ8jK/iPGA3KJn/1c7Xp64L/sdWd2XDDbaa9JRcWuAzshs+CUmUXPdwjeu7U5j8
MWZFEncuzpt68uZXhmcrbVx60ZuTXMoif/wwmJj8dd8L/FHyFgoJLdy/VbZqR7HRpRsikMFJaeiZ
lBf7pATsKnp6E/89xK0FusIQen0XEYqsKN9IUCG5MP0cNepPkd1XM9Wnf5ie57WumpVZ67GAhFZx
JGQuJoh7zbFiGfcH5nFQfSo164S/0vTaGtQCk3QApezIAH3wyKtkR/3d+kX93BSBcffVeb73Ynoa
HzGZdsu+W3p825i5CVhrD/q+7AgnMlvIDK5tw8Ds7RPk1PJzgFzoGJG2IuRyGTI8gVEJN3c/yGqb
hAXiZqlDkH+5o6SycIacMJY//KhknaapjB0KkfPYbTeIqZqqb5UIWK/qkZwl1W01EI6Fde/XWZhQ
gM7qOGYTHA7Elvdwb1B3IIOT0Qwnf2i047heb0eSd36aTfL/J+v4QiNQOEY0ghZsR3eLEaWTJfMk
Q5A0P7XDcaVbZB15zwHhUqlgCdyU6EPHpCaQxyZjQQGjX7uKn9F8uY1goiPrFV2SZtxRk+k7z1Xv
wzTtuvtkP8fULjNlVVZZogL6wW+RRbuA77uJcgmL4AU7gZ3ErTGmUSeTY+WEeX7Vgba+G5MQbJWE
h+XBlPaA9XlgtxM8EZ3fQA+BTM3mj8cFSPQzkqemmPpAu7+9pqs2pdhcu2WfzGQcNfZOXC0BmvK7
AEDmSQ5FD22Kp4iDzSLkpyhczJjptPas+npCFRpnHIGywPRF+xCjl8HN+aax8ZSOa25ZIpcS96Q5
E7Ac94faQL7yot44ezRbBTlmQFLc/eE4a1yq1S9vMQs0mE+8751wajy86htR9CxuXN3Xjn3SX/eY
z2yjFPkkIf0DkO9hPRTq3+MrTTmY42yh8mqVqKf3oOm3+bDg1E0X1dTFFyFeMZGYoCDC8X4fdqvd
vAL/BF9381MrfPkWpEDDtbXRxTVsvDW83dcY/KYwPKRvCHgBGSuOtthzMdDdIfFY+DZiZiRNfBDC
W/7gQ9Jf4W2eWBta1209gcdF+GSegApMOfwQ4iIKTBJyzxjkocehhrcpfMDmR7+ES6pIaGuP7p6B
wOCx4J4r1HaokvIdrS1C7HENZOeDPgaSUAXYS1t+Y2+ELNrSOVZMfPQCYUXVMGcShkIGmLgpVgoR
z996sPlt0rLmaAiqG0foWc6+G1tWmXWLn3/z8rbIzFxDkcn7zhLWpi6cbYOb/ulvu+zw6gh1rCth
3DoDkNDMllwFEek1wEpe9c2kW+rUcpzHdacxSVKjAquWNqpYUg/8I3H4V3JIztwFSwpVFyoNphcy
wh6gGa3bRIiM8TMI0NRyjVkOW+yQN8lkLn1CaS9WeFGyo2Ti4Hnv7bPbIkMiQrk4qeGSspO40NoN
/RLOfV9Ak0JPbpaSSPnzfAbQgPsi8jDDmaNlu1ENviLlpiyR2JxgMCSDKKY8WM0DVzvBWPHpsC4i
TUWV/j8JeRGInT/CJMVS35eRp0h75HsfL1URNXP03K0yXKWhn5/IResxSpeAqabgpDzaYQNrXno2
Pykf/VDDxmxc63NL/nWs9Cbye+JKk8Pj+gRQ1vKOzTsAky+XWIzOGBm2scOBOcRkJGHrK0V4ZQQL
/PsnDnz38Qx0QNx86OBEI37uNB39hNmkUee9jo5tCfXeGY/uZhdb++n8qLZLa2cMAIwSrjlmmBy2
dF2htyCkj8OSy8godRyUPu0MBKd5RM2/WJ33jPgF9NcL4aAaChPcFM01UlymFW2qk2A0O7ieeyNQ
ZljEIz6pb/iW6FzB06W/8gYWKl0n4EdGmJkiLBd44xZKHB0x6lo6WgLZ7ZZxjZY6yOLI/FZCLAFG
TS3l6Rc2YZiM+v1gGeIHyYJKFF0fAMXijPxbsOE15DhusqjmxoL2LrPc5g5M1it1t8mHqVW5hz5m
tcOKEqhcp9rtAo1NfZAGbDYRBJAZmkOHDnk4hSedQkPRm2V1XRIpwuyi4fXdTjZ7z5dBbkmVolGI
6kaMpeTxE9JO0hoEv1SsLXAJD6D7hkM7DZFKji5LnB6ymhsB2gBuKpyvcIcUtbm0YPekKC8cIsVX
FlLRfllZYswymFX8/YDMkTCINeMVRDrxiYHJ+NdVnVHnbxewLKBmZxNh2C2EHB3wypixSzdwttoq
Tmk+x8Id81r8GJnjjcLy8tA0iBhfM3VvKuKuDiM8evxcro9xV0YdBMVifvaUs8vH79F4JhjYYGI/
hsZ/qCjjNHZjo3jGAa3gTrBefH1448BkaG09yN8bjkDcb13LOBEXX94iKpuWV+KbL6nnPmiOeaIJ
mQ6ylJuVhc4cS4rRFHZ4gtza8WvlJoBFwLCOVIzq72sYhYSksp9Mmt0E6HWLm1n4YagA9vHbmsgY
ygLfVpxrgIEbQxAJ9MaUEBjqs4lTHyLxdiP1FnIUaPnzZNwMtOsy4MKtFBocZht0S94dW7irtqZG
LK1IFSsbrMFV1RBXYsQ2QqMIW1fG9VqlGk2tmsYuM8wQRD/0U/RnLyaBRJXuXKyOR4rwmFKcPlUt
dLXhEVbsZomEdm7//RaQOXJJaw9z+TsE+nfWtK03oIhevc2G3RlcMgInpj80NwxQMdueGZXRUCJ0
dOZoRo+I36dGB05qepR1fjSVBHhKmU6m/VixCrQkZYUXQDXE2b7JCSo2SeMQTyjZUHZLCHVHyo8X
hq45+uSfCN1GBNS2ovyzuY6w9tZJBVe5/ivJlV2UGPb7q132hHUQE3IudJ1Rv/yk6zAoAdT9Ug1e
wCa2uJxGGM7rFR1/xiFAKM+C9tXdVAhqIsrg/nHvW8Nh634ZhdNNlsYDXeuuOIRXuQ+ZoIfmStho
w+uo1cNydk2/npIhj/5C9iEYH9mxpNeySv110C2utzAJyNCoc4vEcpZofDzBbgfmiVKP/qfift+m
LEH8HDoHVVHjktymQgHji5mtDnUcNh0/PwAhuJA292ULgX7ROH9PzxWF9MZZtphTznj6VNUkV1vR
JNaH1XeT3v8z8TMjs/do7Y7KUnMn4s7Z305Q6dlwOghwBIN/MxqfKYDAF0MVbsaK9O+OAIaLAv5/
SsbzR/obXHSGLgoDz/yYrHgcB5dWYuaN7au98ojY5u0ODmJSgFaeIDryoqwfnAD/sOl54NCZK1fh
9J+8jUwuYwXMyrAcqVQMUcmSDg0iYRy5sAwg7u219zZe3iISagj4AqwC4mH1Scr7V9tE9o7xzQEB
xVktH0O77P0Cl+A2tEWwiWqK0mL7GruNgcXjHKF/+uiy4GohzOqligXpLQOxQxO31mXn7kF4owgP
5tjBSjBNLPtkarbhfS4T+M8O1PL9LJsCYKYDnL3WkSrP1AK4qAkR19BTuCI7ZIFG7xTcLpZmO7/I
fa8q8Nqc82wMFL/vD/HiOIIBQ0Nrp1Xs2hrjHJ9Q34AqOnWwRrLdNEe2IvdCWtvO73q+LUovmnbn
qQUEtkyJF6WI3wC1ouB2p5xtL9dw4+D1zg8MflDUc62pUhGovgWXtsJUSg2HPgApmZRmLtBxy0f8
l1bPIyCBmD8JxztDe4qYrky4nUBDRKIHz5XeNWjj7mZNrPsLO2HW5Wspm1DApIq/nJS+yySSNz/c
/s2IaTjwrQuzP6hBBzq+AN2maFLro4lW0mbDODyEXenO7LY/6J1dG5NCLeMxbdQv+qW0Q0d2ese3
G0OpaQfjdtu6Lw+ZaiH9VKuD74Em8HlTt/g5oP2sfSp/MPM6qxVxdtgZlaXlkVKjL+BCcQXJDtNS
eDwA0QMvOTq4X5otDFLC33QNty1MhHWjrUNt4QDCqKBKknvtVFgTaKqkWo6VVCrpX8OV7krK2dxq
ASxydy8Yw0kGT2bkZ6WG3j0Gah4UVkKoSab/BrA5y+xMGfLH1rXtOfT4CVmkADZplJ/OdGn5oK1A
J4qADH1MSkbdSp1+hFUL/2uydLGF3OLltB/PmbKGD01jKXoNdcElWeiiS8lNNqUbGOQnYtf5call
QRgpqCEwSOYZ5rUzIFYFUQURupiKeVgmMLMr3ORup3GPXmi/boHeI0zWEWTI4whS2GZfm3Rh3xNY
rVe6pztVipZrS5BMVodzJOYzEFXc/J2fo9L99qxY7nEwDD/LMatmjUxavKgaZjHXe4OqUiXITe/W
3mElM2eUjh/sZbiLlnw5l7xT5hyojJQ0rol1LjtOgd9WzH1gLewbVKcxg1r2Z2lGgFxNmyZuaQUH
YzXI7QVWHzQ77FFeB13cFit/iL1LPHa1/HFBnJOithA3KL3lYV3T3eyic+1JFVFqfP26kicHtYXU
oRz46q+ysl+Uxdr+RZ7VuoN2D2yhoMxOTsAeyKqB4/0ZbxIIoKYc95PYJLtEwvqowuyn1NTz1S+6
D3P1AqMouk1SfDyd8u2aZdOCB7NIK/bxm778nYztFiS+leGM3dBhexQ/XQRA8enU9MRZLKZz0Ps1
wbgQQKWUWhmh2XFzJPofu/wD3ob+kN8GNEG9NvWOtv/lPNE80yq/nU1V7Vn8TUC/Rm48q5POrvOG
EqoAvP7Lb9iJFMCr8W5VXXlYg2u1fiXuieUHdZJH6KA4DvE00S9S23HCKLnCjX+GEsjTdPAUHPNl
uiFLucl4cFd4yL12Hb28VR6ca1z7wlUw3nExbYv9PuswQGG04r+93v0CprzQD5GQSDWolcUQokqH
nW/7TUrvB2WjIsiiUqAW4SgU2EcOhXMKmTRaEznfBZoxVxVJs8Q02s+EZoWb/ZzHQt1FSezlFl64
HAMM7B5tYGDQsKstw7PNhnPfi1mSPmFBqXNv5BumPQVCcAmJ3BIxqr+34w5JXxuHvErpQ7cZ1/5K
+GQh6WkS9VoFnaV5+cmW64sSgEkBEMd6FLcBW++fpDBPefIVfcexFy4Lcj3XKXL96HXLUPxuIIs0
Q5yjEVq+snS3msFfxQtWp3SFYXu5eoPn5IcaH1DAjk9vngq9fkTIL5c9aRmRDX5ETQzP+vZrVA+l
jyzRgqvGYWV5BQpWB6xE4lOtW/7iGjaGuF+wSqVhjcRxvDtPqNTZ8+5N5rOj/1Q2PGOmUmTxdHKS
MvG1HcNxFpqvQK8zqiEv/O/0YlMcHunLOc7hHzArsrR2K2jq1JoAbt3wirsTXUWf6q+rRyOm+bMN
feWaVBMDwkWGoGnsCj8uj8EFsnla2FtRMxooCwVf+P6cBBo9WtCN2bC+E915+ymxBHpxI1Dgij1d
/j6NYNn67nyZzidvrJ9ZYEPnlfROloEdsMIa82TCjtce6bVOJ/kvjbcT8IoRsMXjo9eaJy4IyHRP
eR014hyvaJg0GxrxR4J8pBWu/i3dNuHopTXV9zmMCc9k2JsPzyNZdvyoEwGnd8Prc3tuLHCH6sSE
OW/M8CN9aY10nIVcyYUDvIH1KfEdRx0EIeglqw4YZ/myKIRyWSf1B2Kv+Qfy/4vTjHvAu+u3yxyU
OqQuE/KvfkAqw1CgVoco2hRe0Rb/vNauoo6yHG0HK7s3ZK4LoW3/EIe4yRABWtO62cq500XgTERt
xQ0IPbgJV20uz0/hJboiS8CeYl3DRvTePI6Ozx5s6EVJBv9CRApGR5bKb5VawegIIe9G/hpgHFUF
dkWT3ekuzhnth/CICquNB0zCvI5uaQjeDlgMiaV+f77pLoavhgJG+UxMFX9k51BsrDxSKq8ky3zf
9fjYq9Xhc8p5pTYbqvsEYk7N2ZOVY1st5qYI3QSmllmr1T6oTf9khBHalqfYwLFzdxpcFJkJLPf1
UdoaGzv1Xf5y29Vyt89wt+Uq5qN5bI7qh3ipG2bKdR6BGn6hmKG6QYWazA/RclGOkI4L7NJbx86Q
l5AGfiJvMb4SNjiY7Vv/i1QHEmyMViQUNYzZBmrfzbcHEgYlSaXWexSjMTwcLCdAJqFbzJYIBja7
DmBL7tT4bsp7zKsWtHueFi4+rSfqBBX/b+AOGCW3grS5GnacJXiJHfSzdvHzub+uG1Zl84EHe9lw
Gs5SmS5lKeKCHfsJ+AALTVS9DhDB85mWPNzF+F8Hb7HoeJzoIyEsm1yB27usLGCimzfb+tUaVKJJ
z8YmSJLxuXQ0020tl7HJiU70GZlC/gQmZcK1tMUEEz/GyE8Nw75gR65ox+HO+XBo3dg8U6n7bI5A
3uo6LWPco6W+Vd3lGTw96sE5iMB0vYCfCk30p8EJMtK8xvQa2mNQx1x+02J58epvVhVPHNNNLSe9
Zgs0VNq7Dy5KY5vA51bedgBdAqg1eQjaaUkf/ndGX0iaWv/Tn6wlnYPqnIfEd4mH5aAFQx9IevPB
BOPHwtUz/+FLrH1RmUCrI8uM7xqseJRdSq1zh8vb9EyNy6BaHhRQH9B0jDYAH2fBudQ7nHtIbKRO
64o7JLZYKCMwzwNO2SyupYD5c6REfls/30mcUYuR6t9Bblo4DpEhmClAGLkHBZY+zjsc6d/Kx3Nj
ryq3zhxs6+3xedeV2EJPPsAUEl861Ssb4xwJLkvzv5ktvmzxEmflyS+KM31EVFoDthgkCWgvnjVp
HJNbW6nyhgz5uy2SErz6nLc1PmFgER4417atVpltf9BQweVNASXXnazHupkvsgLWWhTPZEwA8TsV
uS3mngo7H+ekdz0DUI666S9qy9n6ZyMDMgpPP3vKIBrfsA1u0UbIY0maloXfxZLQmOJ2Np8qAubN
buKgSkBJKdxH5URAUjR6xu4GyGieR52AmwrnUUTaSf2m+3QE+KIEY57pgsW7WS40ffZEkahJVKF1
mnDVUTCZHzBzN+iSNMaZ3I7jndQ5mfzIQNfBwt4lplvyE4+Iff0NEBW8zXnhR6keYPjtQTCZdSle
AcaPvvqRjLxrxZ30VH5yZWlse3ceCknz9g2xDE65elOQzwGBkxTlltGg1I20gc2wSIm437KQRPPX
IoBIvT8IrqPExyY0wIPhEUUhB+Ns0wuHhFvIYAopYV5GdoSJPGOu9/NSl8mo567w7jNxEw1owTsr
tMwxQvGf/tefAZdvn2XXUW1Su/2bWysEbdrZ6b1RuxXaM+ndJ6PV4q9dSQmi9UukyrUeYfcC2Hrw
oinRoc2SuXBqyTq2YDeO6czlxDUy+5HNPG/hdBlI2IO8D0YSWibWF0xH4bFfT1jXWF/dx1Ri483P
Jl8Wq8Oq13BItEILXhrEVcLPhKVJlzzkD6K/Pe8xvhB0cdb8scRnLL16jR3efJm8LbzaEA2Ucn5P
QIsug1HBYg9gKiKuSr/5s0X9/dHutw+iRgOLZfAv51Yy5hJIAuWkG+E3a2W7NKuAMmhKqlEfVsKy
aPqI+5uEKUNPNOOsFd4CP7ISauO4TQniMVItqo9sHDFbPooo62uH+/8Fsqdu8WAuDvgvG0ytSqE4
wy1Atz4oc2l7HK3FzAr4bF9FSGauPjhsDKDBbWiqAJsOvpn2SwVVzWDvoDq+tyXK5l2HiVPYhcWm
JSit2gPFSNI6OCvHeAuctjQgadgWnibnUjL6+MFVzNPiJ5t4rSA/2V6wtLDi0MAf2p7NWOKMu9PE
QSiEkQ7mLP1rrsRZULOoru9aefzjavJ491BVMcTk5Okvx7rWal7TNfbvlmqIiSIgq0x2CeMGOl5A
1Qkfblv2K1nOZdYy13lQu21gaSxqvasKv9QwMeNmUowfauanRM4yDFbXU2NYeYP5up478Nu6rYp7
vQJCyb3U0mZaccGcoPoX07AfP+QLT7PST9aF+JiL88E1cgT4WX80yajwFUHR8mklROfdd9tfLoxd
tJWOFtwbJPQgpgmXCCKlDb8jgTNEERzPwlwRY8jBHKj9Wa9YtQ+9mgdQMLJzbmaCf+ZqpBZIVO+5
skj92qmFTYqQUSj9RjHWCS354R0AuYmnkvDhyTzaeD6lbGo0uGla0T2w8D9ZOsnLs4iHjY8cGvhJ
k6SO4VgtoLgfHzjAfhPpkH8gapOnRHHfNW6BPZ4ccK3NEbze27zgL18geRDwNkVvLqcG2neORK2D
xo9aDuxnOJB29EDvw64YA1TiqAIGy3iDusfNI9l9BGiGGBQ6mSLhfrP01ReR0j/vO20YiSOoTD7x
38MnfLvTTeryTK8G7A/oiuWmDIY/3izyMvhUqlA4Ve++6ZK+S9NxvzUYsRkjEgEo7LTKWIaG9Nxb
tcebJdTwBiGG7Ww+VtYTZe1gqmiuAAJZ4NQdBMvRcEdaWpZiMi6L0dcs4d9BMn+yRvf6w67sNd0d
qeGme/W3+DBIVu31wwjYW0pr8FxqyV9sAjBHGjA0SZXyAi83k0wRqt+RjA5xQqCAzLhcut78SmWn
eqIqlx88Gkdp8KitDvOAP8jhyGpoEYHt/582FRyjCqcrZylYu3TLmJX7tqwJUSgyMEg2Un3uYwVQ
BulOixRSECB1KMxUJK2nncU0inAvNNcUFXCjtnF3T2waoJRYr8skyxWDGZuwPOjAAT6EQT3JQgcQ
USVLsAwObF9AKESECeQ7z9q688vp/47/bwOCA4oGWJj8/zelaRM4iR7ScXpnB050A7IaMt8hnU06
92j1J4//NLCD8ZAX06e92AjOILdKrwWniKS7xTBRaHAzGsV975o8jXGuN53L+9EB7kRiOndzr2Xo
epuzlLVbkCkfK8tlwffwcmkgijOuNriic+fvowTfOGygYpX9WvNif0hC1DIW9r0cmrL13Xvnynhy
ANLv0Ok2QsMz1ah4pYvS8DNuAK69TyWnh09DrXzt7ZWML0LaKhtdJ3dsi/Sdw98W6Ui6MxG4ngPk
ytVhgp7kbwx7rPm2md2o7W/PJmI1ni1mlWO376JadZKxQdcA/tOIZ4m4xAO2ZY51PeOEvrHXbYk5
Zo6coq0qb5snPXxsO9v55zUJmSlXfZm1imjZG9qWhtTQIniNUouIDRHZRZg8zMQxr3CEwO0gxl1O
Edt2BN7d6Vj5qy3uIqQnvDIpuYQy+chQSSsgkMp5ZedIU/xjJ6hRomhvKJt/xf/H313PoZO3qqwy
0dN3zlqfjW0F2grA43FflHK8qU8g2a/SGrPivspDQ38Qu6hsjAOeE8KsPwqy0rNRN78FyNqOS+Vs
1wZWKW04Q5u+6uFXVaiEWrv2ZFoMdFBEvUksoEN1CfyBO4d0TYEEIwNuUpPMVpPf5hdmZo2pBNRq
ooNYyLOHSZ3JLkMoyJ/sp849KSHJw+gf6xnt8nykiMYgYThCQ7TxDLJ9WuiWGNx1i5J18imiiJY0
+7KEGEkUImeNHPxsXM2CfQaSS6kC5iV6FaQv3khLniyeXwxhmo9pb8QQsoIdjv/n5WIK/v0zLkQv
EbPBzE209tQmOWz7iLo9kqwsuhGAca0jJCRosLoHti9090RE3lHIJBsSFkIpobwtc0SACEys47Ea
H9jSNUhiF5kL5giz2HhD6uJasplZgnbRKGZ7QKgb2EUEw+NdbH+qZaFDOvbnUDibOfwmBIX63ssX
Wk51EXelx+DQRhYOSj5rKBGWOXpve2C7Sb6KZFRMrWZeb/Tg+zFy8Ww8FNJDDp7rxBygBjEmcR4p
+WWT1g4tL4yASifAs8v3hpos0QmmaDjz6jVSNk7fqdbDAzePMeyKltZJne0PBEtTG2sETy2JUup3
VcIbm9zUbpDbMdV5dP5w3e5B84MdEH9XkUh9USbf/eiaG1l6NwxxOTpOxvjyG8NBsKmX4J2N4HNI
Z+kW0MA84sEIf4tMstZFqCVduCHZpGN4inBLYf0hIAvG9sVPW5ZcniugsNNoSEWMX9fKpmHxufke
96oiTMFsnB/vJvAhHNz5gIvyqnLdxtHjVOOrggH+IoFaqtp8ivL3kZRDcVfamU3efda7YJUxr/Xv
ZKsmum/iG+I0D7k19d+08JV+VF3nP/g4Vm+Ss6rMvExpkn7K8oUp6PYs6hR2phf8eEIIV5/prOjS
gRTEqpHtkcSa2J2VJNjWveZZa6QEpKFiW4JtazdXpRpyfBXuhQ2P0gWmPX6uMgusLzW2r2iWWb+a
kfaC2mPZgssgqo0GHl39ObfF32I7tfrL+11G5CMF9LSHmNiViNV2NrIs4hp8DgfuOtuRZ5OnQFQ3
l3g8VHcQOt4ZFJEp/8KYrO41uuIFqEbS+/p630myU6oq6wQVMQ0++4NA/Ts9qaiUfDn3EacPkXtz
Gy8bcrxihuy+ZAG2RR2addxX6FNv24BXT6Ltxpg3U3NNvrDedTK+IRM7typ6H3DrTtetCYgSA6pU
eHfICE5beOwkOG+yH0ZdaKt6DiSXJEwII9gZsRN1jK24R01DjhEVDkl8ZQycmPNMPsvG6HBca+5z
k7NrEVU7TnP5limm0T2w8fca1kAZvajryaoGT0th6QwDV2tYyi1Zbgk9vLZ5N5RM3jbGClHiwMKc
UdaurCAWjnilM+MxSOPL7fGAxKmrLsqPYvd8uds1clYq4Nuwdgv8d6mYwqUtyMETNJJKuho+3jk3
JHCior3XIZcwXhLuEB2lURhadklHDhtsHacFAc+/vftFqagJrQseuSdHG/cjgQnKFdXP/vDBFR8a
63eiooXsqMKiHPmVFUtT+cz2xiY572X643rxEI2PXyWE3W2Zd9AQRs74/CZ6QVHgBCE/xvXqDqCr
sr3/xO71jD0IlfLIXjDgkUGODeOw/CCPPFPKdT8O4O3KyfXuaIBgJWG2Rw0FvfI44PoVFx7xcNlH
rASx6pEXEuTjYCLUGodeyxRKY5Oj/rYyjTC1y+ZMurEAL0htwR1MRiIrvZ5gMGvkvfsNNMX92W1W
NpYH2EwBsmGW6+cIEdbYN5YajYeBA6fUzwiKZ7JeAIfhkFg5NRr6uuKzEzQFXVJpkeutUWGxm+v/
rd5WqPa0/lcH8ct+XR8VuUZunckWAVJS7lRf3tAMn6mcN3G8dMSvT66arJy3ARFniplaEYqKG69F
CaKCqsWUz2jc3a2YybN0GpcW29cHIl1jEPxbmCmmFObFbDdnkPlytI/Ki2kx9sbcpZXOnrpJyggz
U0RPkkZEIgltoO8JDHYKpI8peougivTSaNjd1RgyMcVSxJomtpJVnvEKlyCFCqNXkzQwgAD+BJXA
JEhm318CdGtxsae2hsTWJvEaV+zgwaM4t4Eh9C7N8NwkqfWf5htU/x3DG7/EUFFalSOBXFvVgaMm
d+rwRYN7YaEPEETg5CTcUsE8sLo7B2k6sk1SjcLn7idutydWAkQR5/FO1RqL07PZBd8B1Q9IvUan
xPexvtasPJF/7HF/tsFqaupX9NM4RQmXFKK73P8otQOsTGG7texG71obimDLyyTIx9sXrmacQ9NF
kp+hZnEFFfZOeqQ/uMbIOAn4N87DOzmWBgbx2kjMyarp3PDmAM1Nz9yFL+QALHXsMOuR71ghDak1
cRnTBGgpzDhtNd/5EvnRNkEFp4ISDDAzQYb4eBWeTtBeo1olq+ZlRLb/dWGlGZJ/FwRyqaGbev3Q
ui/3fu01CcJK9TRZ0ze9BZ8B8lxqQdXicJMBAEfS3Gyq5GrJC35prb4TCkjJhTCddAPLHeYA22VN
u/KqcMWfx45Quugjz6yxz8jBvDvJ2++qPt5npxdFDCmjCpjDJ/iuuU9P17z9PyinoDN+63Yrnu1K
fTgZfuNqhd1ScZ5Mkhum/6xHqkaBOGNgGvhtKXkB/JWYJRMkH8Rt9mEycBYN4jROnhSRgdy3fAYa
ojZamqzxXGemch12qsEpPz7kbwuo1XpmPX3PJx5L/ajBaYxqOs37VJOrd2sJsTRvu6qtejeqK6n2
e7M5LQP6rg3bJf3D8lPqFLxbFkxIf+XK5dntNL3czY/kqWvD0g7V5QUc1Oe63p8mYU7A6Q+XaNjS
mBvBU+613iN0UcyL/5fOfAj+wXV4s4NIm3hCh42xzIc8i62m8L8Z2+ayGHKVt2a5MQ34gmHBupsP
b6RBmCP2fdHvuP1R6FmFoT+xR+IuV/RyOrR67Df0MejzRv6kLkX+vmEYZMsb3ui07bSOD1mqAWb+
Tdlbvg0+RCg2++ccWKYVSwpb6h2yPtWPJY1WqVVsnQwEMRXfWB7of7pK5ze05MUEQWCwwOx580hw
TzH+oT2XA3Cj2jg38RwZ6CWddKsw3lLkxYb8ORiE1PNGz3c/8yo/PJA4GiXyP+Egj+r8eDtzQHzW
vEJlNzqyXj3eytlOgv1Gvwk4j4BgjXJ1LXhBK0jpSjyCGvwWOVBcdeCsJIk9CrizgvhdKgXsG5bz
z9woGcItzIv2DSsdr2fc3vBZEU2/LLqpl9KLnvfBwwEA7nBvFMYwKgk9doZ+MFw7gBrQ8JpOdtLQ
DtPiYBX2rbbI9ef49JN0leekSzUKJNZ3DL3vNYXIHmqj9YRn7K8ePGdSW7NzUVC7Qy/61CG+sbmo
j1y7YEDTwgTwUu/W72m2qPCxylGeFSM52u+KeDwfo04lAjppZTd5O/pvELtcxwZrEIaVPiYgT60s
SNC1UwT6lGFybAfuzznlu137PoVoJWl67jyv3Ubep+NpyWQAANj99x4FdjX7DW8rpoCwi78cAJNb
dPehfzgM4fsMdLlDXNL8wcEQ6bkJDSD31WN5FsIUuJxI/Cj5HFBCX9QgdGeJwHky6zOj0+sd7bUu
PY+aot09lefZfPX49nRW9FYn4j/44GWMamA4T3uhbkYroyKl9wI3JQxoY8tlxjSpQ1utRqD9fhlS
JiSfu+CR4WtRKHewiHqQ1Idju/OFEp3kyGESd08xNGYeiXqm6bJgQcNGNSGch+Ws8SDlh51+rzOF
NDsRdg0uq8cYPMFrKaSPkm71vCO25KF2ALtseDJhW8gIgz8WPDGDSJbEk/n6g+5AyizmOCiKNFTy
rzWsksfruxqJ3816aUHCV/es1tYYq3JQvVWXxF603721K/xJV3vvNN5qN2huZzvJkKY1iWp6VtHC
zFXSSHXPUov3ftVGn4RPyhcTOH3QFI+cPYP7rUgL4idhOa5Y5J8RDyylxmwrUWCnJJPmsKdb+yaz
CIzNpGj8QF0JHTcBqb/G9d3he+1zAas/OECat8OnB+GBojntN3bBm6KKeiRf4iEdw9cO1OIrQ3Y0
J8ZAy+bbB2mZkEh9IEv052AUF2roPkqeRKCe95jQGDdzXWcye8lnn4DLM/++B4j2nAxjgj5BW7mH
DOnHzHhY9RDTZdvgEtQdb7jOmUBUeudQRRaQQXUojqwYbPHSsVzO4JeTGebp0fBu3tKaJJ8VxmAK
BXft0sWKno6MifM5om+aqXjQbJZQf41RGK1emnoGgXxcSue8u2kkxSMi5aHwsqKp2FbU5BOcUy6b
EserjxZoZ48x3ItF0gtzRgVu49fUD/3MJwkmuVd6u1Of6jeW+PXJ/54hXZCT9M9qT41vM+RiYVHk
K1FhOjYB1krdMFT1Rstg/q34/VRVFO8DxtnWSt9fXWj1B3galt5DuT94lMGgWRuTk6+cjktioA57
n6hjA4Xl8yE8IxT8S2MQgc5nSFBr1j8FrJyFU3tEVgNi0ZIMDaBe3lGIT3S4XH2yLH9wqjy+Knd1
yVO2YrImSoxMiddjXXS53SpLZZ22toaq6UujSv474gQS5IKFLYNn/W7mstOJjg7WKFGtdDNbbyCv
IRIS/KZsjEbPJQwGOlH8pWIY5kujsdq3ROJhyaBIZrTYGOsSvGoGOGaX42Qr5yW7jxaio8vjUZFM
GDf7caQWb0PTFasxgCMo8ES53Fs22vE+vIS3O/HpNDJFVZ4hqTNQt0wNCz9RqqisRBF+QERmtyaO
lXY5BGwE3CrpdwrK0qbHoD5pdECaIT2LqXmxnGqaA5aJDLY/3L69Ss9EQeRCSXGxuuo1Ct7K82kX
gG6ur7+vJG6GiWV8J6CMvXTL7OFb9ZgTReHm+2X9N/Gwhm4KIu+xQTLc5LQZTtSAgQ90KnYQGBGI
g+1TKTj5Oq37MQyIefvGgXRv6nT8S1e+BN7CXaesNUBCVVA1VoLxg7hC8J2GgE9oiQ+Bl0cY1OMj
cX7dpiJKjN2vEKsc0/OW0njMtEJvAZ1ge5oMlsQQwj/lZKOLwKOUPSNLTsgqm3dw7o39IhXXJH/A
aKDNXJYnxQIIqAzvYWS3CP+BhF0BBWAOckn5hpe8hzkSk0pqSojj28Rm9lkWQ2h4Z3j57k/PRPMo
lR2Y0iUeY3QN2BT4+6Bz/1G06agwhNwOkpFkDegk5EGJcgfnY5EUhsyw0A+bD4FjASomXtwIbW/i
BPLAJXZCK3ZD/93QwRF6TDvDkXrUnEAzOOSIjGZhxt2+FCkO+DWQs3MK5iHMMeP4XtCvxsDPWbxv
+CfUk0++l+J/NyATVf+fl53etadIKhRnicA1uu7GaP0cyv/IE7pRjhZr+i82Uoedd4H5zWrEOWec
LUZn9aC3oj9C7+32D//GfeWPbusMgkrdKjEol2UcMaWewCjP124EKxAVDHyYkochAQqMaxljuRni
2CY57cfoztEpTihGUm3yizYQpsQKnwkkCNd1CJO46JNsPYilCLgc1O8F1v888F2FJhpAIBazxP+0
rxN/lDEQ/5/vnVFlDEUKRp8zzqEfrIpUJz7Nid6EoL1Hto3vi1rxUEgDGmpOVNHzF3YuZ4NOzOqV
iYNFQ+WmyDkHGYPDKP6ehmaXJszOJq5IksW//cqdZvKjxd9827UyjboIS77hLTAwqRdvpFgX3YDE
CznJb5HWsB7Jc3a2VN1mRgb8F4gYmBoGUn+D8V5MDUIhfIpjsBz8H9bv3yU+EhHt/OBTpiIJX50l
32osLOLTAlrUbVQHgZz0ZyTSNDCswOaiuNBooTBzKfVLK8puEf+hgehvCcnwocKaUx4AVMWCedyA
e7wfuRPY0QMQgahO3G76nU9jGDPfNOW7R07m2WFymygPWOjRTlpU8ZJSWGovvQ04pX5UuUkix3rf
uGPOvo4PgIFjPqzajNOxZUp7CHYTra4I/9NbBuBi5c+mRsUCZpBbmk40AvbkLFPdvf6DRvin+ADl
xAnfrvnPzH2Fwp7FLNWyXQPbYhGy2lP4IqYfBTcQvnPv0U7spsl8IwqMEYdqIZE4GGd9T36/Ovwa
EVEdj4sfmIwNbL7W6BNN/4O/LquswSgF4u/VYKQoTpZxUJ5OoZK+nblB+o/LBajAFR9n/yOPDuN5
48yHPm+PLyIBD12aMHNP0rFnKgdKdB+c13uwMV+mDq36I5OO/c+Il9OFIxLWyof8Pmq+CGxibTd+
dDnw1APQ033ZL8XSGWTKNKCfEQjEndnDZ73CyAQhYPSlDi3ZQXjOvxD7gdtDKp0lMMzyUQiB5cJT
mhd24iItoHUQIy9bf0YKKQKnyTc9ODRKqi64gXaURqMdKAWan1/uJeO8TXXgn1/wzYzi3jxFltMj
MZdDqGMfu0gCbAXXcj5UWjFCKbjMYVUWOAnWvlNY2A6cMLsylE2WR6ggl0cpzJrThBsl1gGd5A0D
TR0C0CYDIM1KevJsOa79of2KmxHcf6bjN2qNIDSRYtZLd1vyhAoyU6EZWbhvd32DCYNWfXHjnd5R
w5zQ2VwIZGepldCKOX4PBYG7Li85ze9C6Kud9MnsBj7aKnX50AUyKUWypIWZweryNtexSyRZ0V8q
ii4rEkbz1lccDHXGBQ2E6Ruwb0gnjTBPtFA0/3/RSx5h/S64W1e8lCOWyvLhI2Gb98GG7/CtKrZn
DhLvhpYnehlJSHPobNWVW8xJZYe8X4/xQRi+c5tJ/EaHNoLG2VSD2dOcib9PIvtAnH1wlguDJCQN
1rTFT0culO+C+h2BFBmr2TtisZtx0za1DWS7br1Q4bmgYwOuo6fVk09FBNeG1SMElUdUHXPkqnkD
mAR3e4WduiYrlKw6wT0h8JEtzNCOAkfANm2bZ+2obdob8PjrmRa8JAIRFvR8O2+PiUSGGVujtW3n
9YYGg30tmWvwTPaq62DfvvOXCDQehJG4P8J/ALk3IJAVk7+7TdoyghgEOIl553kI4aAcDlfHMiry
RHOVhd3LZNjhZJZz/A5gjpG+GUMZ7f4cPXauA2G9zo7hBXI6bdPNX64npjz7jKzjsCuXoRCKFjsv
7bREMopaF2EdVSOogAZTJuT2nMWoI5Czmb66TCornosLJMFFNHAF1+eAshTzfRwoasTuT7NYnHXB
MSVZL/aPrDl4ZbxVrQSpT0tZutvKlZG5B39/hAw3LNsb5TwuyomoiW6u8XdPb+i4NpDAwYCCQ+W+
E6xT0MSGMhhMUdZMAiLHRxH6cwxeBWOjUM4ai2LtBEYhhNMZeGI235yuBUp0axpYeW0So7kAwv6G
k8JsP1WYaWdIijpwfVbEMQG30eZIRdSfAPvocrTZKp3e+Fm8EAnn1XF/B796FKLCzJVHaW+oBbLM
0wTiWA0FEBJTnAWRJo9dTy77UXyaIRbH111mOHe4YPDVi52vL6PDc9dKCj3ftKEHc0fEVLIbRdGm
Uyc7aPc8RuCOsnCdR04l0cB7dQL4fXioQFhRlXHbfYsbytYs9GWhCj0CU4XZbTXu0jgNCWjxd7g+
rQpe2laKbU94nBfjA1lusPXQIn2yuwiT0/mY+uV6Ym/3yvvQHZRzVMi1xR2gGoLaZfUlgb3v/Ex7
uZZV9M3ugwcK8JEbw77z4hWFi/nwLbKfpNAIU+lGKRtXoIzNcZW5iZs94Lk89Rn0xaiYo64iKVXP
wdFCc9raDhEAYANcuiMq+/TMig9dw7shxv0edMhV2DwfR1qJ78FPpjLvywMfAeJIZ9u8j7vjVcoW
92PrQBmzPYb+69GbcApQQyWac+onHjDGT2AZCUlAv3i9/4rJScBtsUwNGCmU8Z1UvoENiM0RciKo
r9VM0aUYUp0vIuaQckWs0WlMe+a8YUNXwMilaclrSidCP8qHSQOiAwCQrXImsoEnPwh98vG2A8iu
eFf58yTnjSbVAAAAyLL0SqEbXd4+IFHPvwblKIyWE6w5yVu9zZxM/LFaUn2PJ222dQrZjrgPjj2R
D9jFNzSzOITlDwswDXRCoqKaJrAprjh8VsJh4f0DUW7t5LIfQkSdE+iEGonKR8lla4PSTgTu3vgo
PtDH1zyZpWZ8XKR6QfDu4vvByolCB5UrZFgXAA69DuE+9AdDBR/wbIKBSyIe2aBMecadsktl1XLh
haDKv5o1j1ZSmJPSQ//RSlOPflNM1CtMBYqyLnvpC5sgs3ONal0chnyCLe21wBUc+yDO7W0CHMos
L1D/QxT8uG6mPVQF6QBUIry+TNaLixuIxspRt9k8duQ+cA3fGBm+NipregbT8mJFkTpOzNeQ8UXF
k/Syorg+VAuI5Nu4zCtL3gWiudgIFixudW9j45YGItrWHouvsXxBoGia3DwOlxecY93MUs9h1Whn
4jKF7GHIF1r1lWXI+XfQRkKPele44mouzR6YfT16tpYi1l7VjnQemYA7gJ40q7+TEac/YC670FSj
SPnbLm9OJxctwU3XLX317n9Tn/MPPTRg/FMsajyRXMhjPiMrQNxjljfCGbAOZo02E3JIRYAMrxmm
28+9fhAFE7lHR302mR2StTkVWzXf0gpqvA8Uvb4N1haVoWViJSCYwgLfl1YLXeNoFIXL6t0W+Zjc
i2Z52PbXtuM/xkFrQi9t//PJvSGiS0LgHNhKma9AHREm03UNCreWterDeQQMlA31nslKeGaN8TCt
6dfEegQaSKRS/v4m8rp6y6NQrrJ9idy7eM8/eG8b+Y726/MyMYuK9A4MTT4qg0khp2NJbnKj3ks1
HxwZNAvYhCTtXn2UEffz427CoPndZVjWW4YaGovbenu2o8uAicuKcGmTVcXSvVOr3PQwHF2dB/KP
NeTNdTDlCFyi0zpWX7M+zG6kYhtp6w11xcqqD43Gsw1yKgPgEO4vbjnFwGMnJqZKKVnGbqAN7+Qe
v0Ugr2zXwhaFum0m44MISKu4BVmPFVMgnNUWvwqAsae3l150rXnHudEU+5DWtZ976BIw0I39DNIj
u+hDzPXr9x6OY+2TIrhcrqssGrGaeLcKIdiAjNLr05CEnNUeNnfVeFrCf/HcAup5aG8LlLYw6HN2
Op/QcXWzzWWGCs7Dgn2XSeM1jk+UhXZ0l7vHSvw3SVWsovmFtlhz/aswIbwcQ1IloCANtQGKAGVL
9KYmkNfSlTbgSRzPsKSk7N4xmBfGYmJpu9AuicU8c3aDoCgYvQIvaOfdx+kpoIEG7ecDylaMRpzi
QvArx1wf51rNace7iC/WCnBf/J1ZFqyRTKzYLDTW/4HPI9SaQUL0QtGSPljRpZ781H3Nj6aX8Ap4
tZw06MRbwVp0IhODiUmOFLk8H5xvU0a88sC1oWJO6dLWFpLkxdrQcypAUMdYApvhEL5Idudi5ofL
MhLoWibEdOLPC6j/8nnLhK4jAuf54Z1wKnCX3LOvbWNg/j4XTsfo2p3tBEjS6bFm468QO+d9Qhes
nmIXXxM5BXGihovHyJ88v0Cpi0uMVMFpFOY5qnTubY04gjo2KAj8ghcyVQPR16OtPK6kHP16tzQE
7hxFINw6u63feI7ONk0NCFaghaPFS5KgepfFdC94p+0b/LCo2WAmM7sGzceNwJjsKxuq6HC/IFlH
UjjTgCsugkKurhwOvR2vqDfBnrUHTKjLgaJeukxA4BN7CY9+CPLpvDBTLh0kByK8cjyPPhhZpWd0
8fKVmdOOeRpcDq5izl5tPfFmvfdSI2A614HeEHN2RnX2S9Xf+PaF4YfLFvNPiq08y0f1ALGXIN8L
QGfoXc0xkp0Y1BBOcWQ+qrOJi067HGtghuU46PvzDx9NMjKSRtX1sKBEK3TMrYVpZ8SgP/8i+zCy
9jVXMQwc94qwkNb1aNfZ4+E0xyZnztX7nHLopa3iDlZz5PIoTlHBG37ghfdPAVU+h1zZOYRUMFJF
1rs94CTSYEPXl4RgDvA0JgD68Ai6EIhH/gvJKvQAJYp8nXENeHeSbRWCeZ5yI4RDSJZBiNPT5KKq
/CnvNDIHtG+jUuhNCkqvgzWW1bvV+vZJxWmutVFpNXougcMM1cs+FMXMRkpa0nUz86b8zGH2uGAz
nPp5pggnsgIsx/5IrnsV4mnP1J0BaamTYPl0ORMQ+7g7x4NtKiprZtWP7DVRX3UAvuEe4UN2VpKZ
gdBEwIkDRTjfXMd3lTiUtEpUxj8DJx31PZWAQDL+CoXN+Sjn0pGLe9NY9CBZDggs1fUq+sLBvTuC
sWuVkPD+9U7xy0s7rEIVzYeM10K68epDyNOybDTjSAPqoVSb8pRD5l93Q4XrxFIAr/sBQg4HfPRq
ByzxXTtnmRfkSEjUUjdiHFlRxbpghS0AlGoAeICMHA4e7KMkqKlJnYeDBbXpav4w0fx8oQ0DG6Xe
zgzg+8kpMiq7QaVmV3zPU2NBX9TNyzwhz2sQx2FAX7OP215cDX2HhSWQvfuXORdqgOkIxHV7CwJu
c8aqvdANLZQAgaCo8DBfjzmdidbce6SoxeMvVPQ402VccbXBCI9oleGfV1yUPMKwPjE2qKsoE7NO
bj2iT4hrn4ymC3AtKcCzEsvuH8hHL7w+enieIEA/Khvr0AtqI2gz7iNMd2II/MbS7PsbnXxjA+R9
A12Sbv+slgMEpAM9zj9yUKQinexEp3IakXYTuJpis1CFl+wQAbuAzHSJ9rP9Tx6EY6arm52eHP/8
x34FYgRKPfO73osqa25qZY9VM7AVc3nommGJ+h6q/YVD6YGrAKHoheKEDMzAGbO2Pxf4K1tH9bfe
qR74EUokpQgbOaxFIGq2gr5/1jYulk6qb0bMvYgV6PSjmGSrhpnZ06HmBroD3CQueEaPjxac7sRp
Ddh5QzXf8KsU0bmH6/LnIZS1OnxTuid8/kjzC/xTUE6mkkCjYVSV8vZFjeM3kZZJs7svIBMctrCI
QkWyYf4PVdvx2UAnC+wyEcTDZX9dWXIM0NlnYirBBCNKX65QbmulMd/yE2oxRIXS187WPNhKXafn
zp7cSL/56STFsNMeWvligIHdz+W7jFZix7Ml6eFRUOKK7+4jqmwqhAvwbU9ZVGKbzMXOccWFUOO4
ACi1+RKn5wEBPdO0FXh/bDNTKt0vPbEMif992I0uSKafuOKyoL5UuqN9ZwB58reBHrn2ANZHyVfv
FolUYIiztBjWEZNMzOYlRBLXY4slefZzkwXGzBUp9e8ng3DtrUmjs5wpuZI5+OKikFS5jSOfsbBg
aoXQhkbRl9+TyoCpRTmXPGJAwvfe+OB2fzBh+PwNxEIBrrXh7aeTRLGRb/XUKQahbejgNzV+cJpC
M3JRvm69irS4qbq9ZhdOiFwYuoErsQYZ3a8GhLFsyu6eJ9EjGTZFE1s0yU2X8u7jwaL8NRbgNBrL
ujKk4GdU58wT1eTwEN04Bafxd9EGI96XY0Yl9+sCgwlpgtomTRE+/iOvgV9Gfo4yLzKmJyNIdxkq
bINhRoP0BUz3vHN8knLo/rzGJPTad4E5AtJUpR8lNW0XH2IDOf+SH6UxeKvSbubDu4SlP/Hj2zs0
2V+esGUk3OsZDABKlaDgkVkiynkEGoJQP+gH9g+4BpIrAgegH2ZwwHJqf65UmBg3LwTQe4Go+STr
0AqIqsXYiOWRWu2DTT/8AeizJNCry1H5pVSwFCDKc7icW2CR9q+HKd2JG/uEq3RbURuY0rX9lemE
taEMpS7HkYkSYma1G/GlnItoA1Uacfue+PSVIwUT1T6Ql8CBBdS6DWbNYIWOMYrDeEQctNJXTQ9B
4wShmUr7BCotdYAoDxkBp+ylbGTr6ZgqwwAoeyI8QZyUW2mi2AbIBqAbVAqiBUhBfE1RF8ySv0dt
x/zzMc5ikbSlaoKCSAL3WCc8QOI6ZVWgPM+VZCR2mbmCbs3liCC8gSKVJYvAvIwAj+LK0iu7FezW
48j0OtA9uDRCGuGUmB4ZjVP1fYBIYaAnVxdWeLmFtJqe6ZqWidKErBbMJWkFuxkuHesxPg8ob6j1
3KjuGJ+lFd5bM6p4nigQBs0qzZRY5dP0Cr6GY+BPb6lw9IOXf+sgZ6v47nKK8dVKfg0bi6jfNdmS
Eng0AgteFjoJZHvSk+ywBQ3HiaZWHXiObEiEM1igBWg9PaHsPBDqfz3WEvuIU2NcbFLoV9ahETI6
apaEhwuu9ni+notsx3WMS6B+x0if9gKNGGFi2WMRv39/FF3jCypOgbJ/fGls4lDisivJRejE64Co
IsNYepp2WPU1ialp43YaI75YsfBRkrf9u5Gnh8zwL4aPLRDeRv38BxcHgZoxKWRoDwohXmy3FfIv
o7/EqP8oNp6ZCGB5ry4dboxzTWNqiETKho/swi+qMLL/DJBMKbb2I9eYAoc5tB7r8jkBMaWgIXZb
SYbPxdf22BGJgI4pgNyELeyXP10WNW8FlAqfQEkruIMrkiMbtBrGMfNstkIzjtPrG3QpKdRL6TKy
JhZhtNUakeFP3GWATgt5IuQSd44qiBBp5HEm9cS2kTDIVJPFbskWiQ60rYfymxWBJHxlrUl0rjlk
Kzj0Okdj9pHi7r7RcXljCAL9EIznl0bARndJQ6TLD22fgxrxpxm5la9cmAwAv+CAykxlehnQORi8
M9mA6pkp0nLL9E+twZxmAF6UgOvtDohqpCOavVvRZGFvKfZjr+FkIturE7BDWbG/djQm15+2IiLu
MY/B6DjRyduAAkn1F9oKjkc9ql75yqQ51CUbgorLyVopR/dCAZSeIiIp/j0MdEarQV6I/6b0XfcH
LXuR3rcCJdWdEnD+0PE9U6b8KAIF5ZkKtX8Irr5aY1AjwJaLBVxe4OWOYLyN95FyOIa/e5EuxueG
rEcq9EmPSnJmnFu8eO0b6AU3NlIJOtKJqsgQJgO0YDwpfkWxj/Q+Pg1XWwsz1/Y8IiUi1+jkCt3z
gQkRjCPZlYwjdOSAnO3X1xvwk/xZ3e/IfCL6jR+R8/oXYVetIuZNQYczvNFQpYss6A3BkD8Zv5F5
uWJ5cdrikWsAZGbRlbS4i55QCZGTwK8/LAk+XbtyZ6GjL3GU3FRP4RHbDX4rVCTX1msphYu9YEIg
UjQa2WVBO5spp/rMST/MuCwuYmQVErQH2WixqYbW/kTAVeh4a5g5ZLhKrnTzHRHjHs18DKJsIQPi
NuCIfZxYRzCXDCpbGbjK5NXTP/Hq6ucGj9Wb02SrsbJpYXWQDGUvW0tKvzJ0/RbMa5QidaGpdhE/
1wwjMmwRBvKheCHNoWMcINhf2mjLDSb84C662weDc2OSR3eW9U3gEnB7IhEgaYN7hz87V4nQnI/Z
u3YIz7yXWSt8LRTfJzuecWvctSQ9CL2hjGwIEjHqmIu1DqPtWQG+EOAsgO2Ficcs8vx1EqCMScx+
G8iOdbSiCMc4WU8v6ABwS9bPPZaddYKSvhgWwr6lICB0iXgndJCTmrj/7zLzCJ3zGO5MCUTl8us7
1j7lJe/4kadxo3nNEzACi+7v4AY8JeOz1GNwPLZHiVXUcquROhC99dRqpb50alXKuyeyeb+t8e3I
CrLfB14YJFWU/5BQJoADVo9CfUDwvN5i2ZQYbJNXnCp9SQXh1dk35Lp2N0GV7cLJI21wmoZJ7aTx
GlJCHW7QJbON2L8zIYcY1hdMga4smd9C1OuNs4Si5EF0Q91to8EfBg+/FDkTirmpOaa084fd/sqy
RibQvy9hTZmJfAYn2e49OhVzfjc8VlSodbNGuwd/0wxg20VAKyiTrjZq+MMyrZSEGjcHYae+FZWI
u2jZccQ+jFprnyxRIURDeVDaslTJA9BRmVLeMhIQ+t1jVjJyAeRWXGWMx7oN6eCyB+4+gbvhAJgz
EmKVU9set0bdQvJ4jyosjJy4YqkgB0B846jC9YIEWH5J6b5aAGHZLlXAx97t49wkzgQVMiZgbof5
AADY5ry+0AqRAlYG0TyQIV9wDCvkdPwEEVLZUU4P5aIfnCuLJwR/o44fJylWVbTpBR3aL+bwTAzi
6kfa9s7ibSBT4iZ8RStDthJPrmrKcqEG/hwFpROPsv+fd6k/P7QCEm/ErKc0HffqRViDYOD9Tzqs
4fdXP9CPMknU3tS1gg3DxOJ3mIg+XgkatMZ67sBvEvbhU9l150o+2RM5AxFDRaSQKMb2UXiZYQkG
6NSIlcG16N3NLANlZx3sjatJGmalGC0hnNf+G2SLPrcQ2o/NoI/psevoozAP/1lBZLhJzh8RRwUD
WjKfIAM/YSzqf7z+E38KStkrhQDpN0KZPerzPHsHF30NaM+6umys9Y3zi/xYI1fwwtg0t+o6zEUC
eo5eyfMha15UCmSi1cbX7R9zH/NtkkpXLAcI/fayS23ANnSBZ6rrItPoBnal9+sHP/Mjy77zdYI7
Q8d1sbYaIzWSUPrkaM9T5DwUsvTkiFsWxpGAgr/ZysjwNAHFfsbZITBYsizTVP3ZMMkDRJD2x5/f
4JctguNDBxZGwiZ2+mGATT5OH4y6Gw+7SGRBQVDRGSYzEYo5EBriF1uDL/tmqmcxOeQr+FIaSl8g
a5/K+bcrZURLGfJk6e0wiyg5PlEB5xblkm/TnBb8VnGgTlFvZ8RdiPXthITUfJO3od2msYTQYonY
fN9XzXhSNeyA9p6aBvWx/wEGujTA4DAsr+rvdiG4cg/2T//BdvOKCw2Mw5ebv/HS0OM2P/bmcKcG
67WmBl9kSxB08PWO5kan5JiN2ncu4Jggx4xeSuW7FrFuvFqybwPlhV6eDsoDgsf7cbdIavBG/+0F
J1nqx/Dddlnrf9GUbp/uHHQJCU48+IhYNU0VN2hYU64xuSDCuTlUgqR+X+yhSUV72AYbNn1DHRPL
CVSlbHooetlWQcpiXQ3LT39V+xDlGOysAzAngKnr883FFI8JJBToHg7JiMjq8TkBaJRiQfJV9b4O
GZMVSr9oJnt32yL3ZbblvgYgik8RlOymEv4A9KNFUP9C34n8eKTstQh64fXw8Q4OsLOjqOFmpVXi
QloqJONpXAWhPSbFX2RrBR+5eMdiNUiVJjEfBZOLsKMAnYgw+ZU/wUhRuFLzkZJBXStpNiRa0EI9
0RtSL17VnhVJBiOP8HiahWe5nAZu/gtLt8VqrtHu8PGNBqRdYBS03hvAp8A29H9qsjUCHATZfn5Q
qpirs408ksGXkBZfHQ2jgFY7GAHvICFPfeSAXUHrmkV2B4DDdmpR8ew5HkT0w0/mIWSpGQib6OIt
o6/zWHFn2znWxJys7Ix67W6hwv9NikZU6dQLjnucxKFI6iYzjmLrHFJCc9s/8FRGPixP4rEo40TH
3Np3unqER1RkSLi+s+DPXn2lPEVX/Q72+QpBqYRZBdBGgzwdlzrqfdGScuA5Bsp5xcJ0Hc9N0xyC
vaGCYrdaqMlJJcUdtUFPBg//YWWdcrq+t7bwZqSUx40NrJhwhpf94l2ozMIoIbhAhntzmf6uXd2o
SZ8Nc0Xpe7NJ9rpy0SFcEvG4zOR3xLhX2RfEKBOq75Uir+BRI/Owp8P0U6UQJ2zG8Kkhf3zgDZRg
DeCYH5dVtCObC6IEMs//kRTZmcmNgX+3tdOoL0EMAlznDOT7gOj77vcFvdAAv7JWHlq8oxdF35KY
yNh37Gcz696hb7/J9sWO1+ILjALPur7emPgbi5AgncjWTcTyE2fGI2mRHWmpV7azGf8nxWS3yxJD
rZAFNyDUY2nddX0V/VR/VJB4ZhobYTktCK/mwjKO0HquSdZv2cTvG4ZYbYyKD9LQWVC1v+H998M3
OPLGJATIrGDMGcHcUTuYCyDca2/n2iCUOYZoa+rS507cvlm0Cvbn0iwdK/C4qqEMpaxJ6Z1I0OfW
KQHRa90JUepHpTUt122tFZ7qgrutPzKFXVsjVTJHNuw8s9d9YcW4zJOu8CDHmGXt7a5alzOfoCPs
UkI7XhlMc99rNqNM/OkXwT75TIpoM36U9DI9OvXZMmJu3zz1X7GEKxZ2S0nXrKxJCLMXpMF1GplD
fNi/YzhuExo1NaC/I3AlPXXYv8Z/xoZXT4eXMtSmBCprvS/GcQt3ayy3hLYyt4Qw3J9QBc5hJnTD
xpIaG93PfALe3GLRPOVrgArt9g/melw9HPL3aUa4Teduc22bzpgNTaPh4xdYQKRMvfKWu3WEjenA
JS//clYxx06xL6yDVwSmdPhPgDQX82BKdgIcLXgVxdx3cQSKsZ+IR3ZoqVz+xjb2Jl4bpD5/ofQ2
LdLWuB3VkBt5b50WC47MIys4O7aoISAHK2s8u25L6UoWQ/vA9Nmr8sjV4n9rfKR2VMmeHLhwEd1Y
cLwvCIjaCnhdNLwfOfczRyTcDfBT3Ebk7LK8G2Xzf3f9wejpAhSg4FHZNre1/bLVWrSKE81FINt+
cYXYGS8JqjEoIHjcWwK6YLE050emxXZNrH2AWXtD4TWjbxzURs19rT/tkQh82JTMHJa0I5TkleXb
gU7qRB5Ba6qJAagaQY22iXyzfDbs3/v03Fci1OyIQAXtn8Vcr2ooENW8keXIRhBCKaprScLn3vO+
VW1piy7Adfn+x+a3/tUpezc5b1DJ9+7Pwrr0Z0bHry8khGwP1x90KqJ/HzDTEYeEtcQXqoD+aGiL
utmSt76On0ajuhOR1Q6xtPCiKP+YASRanDuiwL51J/L6yBhBJ0hpiX+31hbP5srs6hGbhJ9TZJXA
j8UzIe/LUa/aNBYRIFlX7x2ZDg81WHyCSoiAW6Ngzz8ASoAe99nOtOxhN/Hbn+np2DCGqver8tNJ
KibkLsTbnldOdrgEyNtAeZfzIgUTaQmmQaECP7QKIQwdiSrsNd3JMkQ6KTe2nv7Yxyjm05zOMXww
d7LG/ODZP4tSvp1VY0xWlXBIiGhIN7tU0JwKZ2+GbQ19oZW2T18jCgvzTIZ4DhzDerc7L2zRQGlU
ZJTPsOvewzO5K1TxnnTzIgsvDfC8WAPkirl6nvHnyx44Jo9ieRPETXrlopxIRQ1OTJeCyN9mrF8S
BR4tr3bEQ9lg1fjCwz8OacKmm8myqOHrHPT2ZGrrjbntnPgdPJe6Jd7fQXmvvNVhMHa0EJSYXnrg
v0+xIsB2I1aIQPgalBHuVi+5JpIafc6tt7PL+xx1SpvNGOmoNBCHQdJJRdLkGQf2gwwxmOjoU2qH
CkWc5tiL6j2bYZ9gvcIWF+/wvwAYStIRs1pOHYqNmS1uQZ8v2z/iJKUsTP6Ni4bHXy7bPRRX0orh
Tq7XJt7GBEUM9MJaLCWNIz+JgCdSrID7WnkVC0Mv1fc/CGulofKJnZ2IITkrwH12obu6lob8W5Ue
vpQusnsLGj8y3jFw573+oppyn+dhjmNDXtyr9TDth8dFvQHaUOK5YrUh7QH8ZcHrIcXpmCwyjx9R
PkVceuuzmhYcTKrIndHXas2NUPDhcfH34z4ozwcBAxI0G2YQjYwSTgclTfz1VJNf8CcvkuXFDgYv
38vfxoA+jLeiKJCt1LhY7YKM3KtO5gxa5OeZuZhFUnLeJqEV596lyEXCPhW+ThlVkuvIuTvq0U7n
2a5Ao41CtCATAZ6LZkh9/DP3x/vzMD9kzt+KHT07sufnAVqTUBtEsMEJxRpp+G599VDz/M+O0j9o
V58tg1Z++qn3jqgTXiKxJoSvTVs3XypUgd5ImFkDQ+KCfkbyR9KURtxSqLqj0kVv6vo7s3IbCKQ8
gXKTx5SRSnd2hJRuLgDqX1jV7GSPmd0IDjEQ5YjgyP8hn+nsAd0ujVTV4LkTvm6Jtey6Zf0kMnql
NrtsCDAlXWHqPHiVCWBl5If/x8+WlpBjwDBD7S40XzX24LfBKgTPxeFPLfVh1F5CkanWKSXZl/sU
TbNd+EwEgmWWFAVNxRRAPRt9d/8HS+gIo3anlwKXZWDtLIDbmMIACgOyL0k9ZqSVdCV2hBGNZhNO
Cwq6estZBidDfDzVYkX39yy9Qak8C/86pGMGetOcjYE5v1pExakbZ9x1RIxrRSaTwOc3+qSLdJd5
2fLZHCm+nPgBo5GjxoVeWc+BEgX4zpE6aCLsTUYM21vWthF8HTXP8VDwQxTORbgpeeh/YsIzvSVR
wgDYmFCUT3kKg8VA5lMCXozuAL9JrXfZnU3yg/nqL+rWcp1nqNgMXJKRtJ5EntPuFUPh49OT6VAs
EkCOjx5DuJohAXNCXIxw4rbG6eHh1X/chv9w5uZCNVMyC7zjv3vD5YzZt2iQaa/v6WtoSP0Mpf79
svPCImq9kiWhLs+fz+qzxAg7pbprTQ4A/iS4qLg7mkJUPuGRomBNoeDTn/3eXbb8RhHNfx5xsj4x
0gSnMyVSjWijFbxvVKkF4aaBhp+lDgkSK8PpbTM/ByOvz9237QU0BYaYqnJ/vBDng10VHch5IFD/
CqDh5EeRlFjrEZNbA6/t767RoMU+nxWWptnii9DZBs/pbXXM5lhLWM0jh0VhsBFsvX72XetQz5vB
tbRC619wBxQQD0YFFqxRy6ME2NO6aInvokRF7W71E6EfoJGXPObk0mgjRvGAuUxB2flsK4YPu7+w
4ueDeFrFsCK40wD4gEdFqVW1lqU7DkTOLJUB8dItZiS73xC14euBwXXNqwp/OeZSlTzNjpjvmRCb
pQYhwWnvxKb8sFPAExDlKLGmNsWt+lpT5nfBB4wgn7d+uWXBrw64AySyz8dG0rqp6mX1wHrnax0T
gXtZLzWEWH4lL95EW497xk+KTRIDUOmR0bDAyArkoUmmfkGYIgkyirjsFtYkjVvG7tpCzFsCRTjx
FJRrvLhWPuXWTTD5oFqss41dj3bjMFOq4OgjFJHJXlWQsVjS+pxPdTjUQO5/7QrAvWm4zQd77Y7C
38tjfqQ6eXIi6k4YrQ7LRBFXddt5s2KruzYc2SsoGDrrHxFIgGL8YRpPYnfWhgmFvuirOBW7pd9S
csJqL2Q+D6ipIMnhpiF92Moxs0/YkgTDoQDCdkbolupSxtZrB6t9qz3aqdd00FYINbG8scVoxJlJ
z1y4ULoV8A2oWl1hc0Eh5I5QqIN9NlAtZpZJReTvhw74TfEkDYsiMOkALx5Xs04fLMOd92BTo5vs
/dkVkRmQQd2uySQYXQB9jVfSg7fB95WEHrFAdfkNt/O+WKgIAHnaLPR+QlkgQJuBKQzeYEQhJzPR
NS0bu1j78pc9NJUtaAewcav5NsbvS8gYnpA806l/jGTx3CuBQzgLBbfikwcZ41OQaeaTPMBtp6jf
LJwOVqXi6euU2NOF5ggPDn1IUS4eFL1heRmSAbUXx4t2tFwDxGtVshJoG+SL7303da4mvGKi/hjX
nPaU5tVovJ7upmUoK7EurSbqcbUsH0qkpfVQDDVTa721NVVoZy+lchNNuQKbeFkzMY3vfnHwCA6B
4iVafYs3yuRZwpC40URExaY9WAI/lppl/dK2J+RMBNIUk3qguMebLLNeexv7ewZXKR8s1GtI1/+F
x6gJAVYu4v92TyUyP18Q9U2QCxpuH9wokQGCLf43GBiv25xbtFqhtilhxQBGyRL2yf8yHd8NjvVU
sv5JcHK7ttSC1D73Bo4NxNkrIuF+8mBLvpDCwbm+1BM1XNEHgho9vAeNQe3XJGI8FOtJzmkJO4RE
EGfugMF2kvujf4MV1tY9p1ceTBu/jfKJxnlrEHIa6EiyOYTxcnUX+A0Zr9lt4X6KghYzHg2YtIM8
qgNbFm5XGAmHs7O17Bm1+oct7Rw9aINIMHtXr/5/cQBKxfTmeTVLWePH915tLF92IeJEj8HAU98G
3uEMsJbCqIaREUejkyjgabD6YJC0voWDMYl9YVFpKQFNIuq0qItgDR/Mu/bFn2fj7CwlZZzr8PeW
4LS8B/Fj3ixSie1G5UGNKNaDyQ3UHrEEzKixy+ms9b0/PNy7gUkXqddqpPmTWUC/Fvh9J1hu3ZIu
9tefaEVen45DShqsh3m1JnlkjtkkY4TrqTMKAI9AOV5lzHzIKmXjzb+jHRGBDk0uYEo8u1WL2PRA
f2aGaV2HSJejyzn4WqI9glAAAZBqPqQdHBwM7LjPPYUEs2hQaUa684oefhcDrlUaDjm5k/GzOKfH
JkA6lvpKeDOBHHXKG2wOvn0WFnWaGeAYnBN7NIqVEDkpYpejm0Fpu1VxruJzpSlEFZmU3NOiEsE0
SPsI1LrjnZGjHyG+TZTHTNihDhA97WMxZIdI8F2HpjsWbSzFl0Dab8mzZjuuZCqtENCpEuxrMw6Q
8iZ1AEJT5fv86mrdFY5Jdg8oBbqIxorM/cnPnTwRTWUgDlBu8dHV60yD/A7qsc6sR1KdSaNjEyn4
mdh8DAuTz1ByBbBr6Iu0QsJEX8ewy0LMpo2pX74YXiQRkvb7Fp8HlWon9T4fMoA9Of2NbKmYcjgY
u3AI/K81ysznDptL0OC3YJgg65CXHb7ILEbW1vv723ynSNps0w96bjZXkrhKHrsCECcZzVPQlLWc
6T+4GiI+o6SchuS9lZ8dXigkqZsE4Q4SdmPW/OpqG/ft3v65w2CdXqk0gkEG70hfzHGcwdFknden
Qn4nNhulEBuXqw9JiJjg+skkzyGsZunHr+/YI39XcsTYIvrAzbCfoO6MqUtkF6UtglCM1Eda/F+V
IDHQFS9fkrnWB54bU8//JuxWq0Yoj0hG9lK535LdpqwD6B2H13UU3kNf7+HLgmeI3VA+k/4XWMZb
32jZHIu8n5OdtwhEeIJcGRdOGng63sTu1q9dlaxvEt1gIM/WzXWwgqkV5IJeUmLAz1SGrRBz9YEv
NngMiCPm7XVl/chQQ3VTeNAVHdmIGvqwS/yx2/XDld1XLp05F8jkVNWhAGohkd0AId4SkoBk3832
SOQz5Y5m5y+fvYDzM3gqtw1g4UnSkOeGArL0/Xf1LY3yJNtvZdxQbvf5DjkP4mClOhcHcdXJe/BP
hbRGa9mUPCNjWU6wjRhmBaYSNukafaOKTP45Usc3xMy/MLAWdDSKtOUPVJS/hwQQrzqtG1aQkPlT
W+P+uJVzE3hVrRWXf7yq/7Gh1teCmc9hdLC+P0/doj5KXpYrCEi1IuK8Q7LT4iF/rjKBJ3xuIRMS
W9zsXy/6sTH8y/9jplfFW9X809ECVdj37WfhH9fgVU4Ia/Z3lIUehbaX4evMBhV19uyKsQICwd7d
d7bVHpjla7jPcsd2jNdq3WuXNwuGANVJsoKU3XiKdYsZBGqqZ6ff2mOW4cZz0u1JpzYvhqcmgkqn
9rz1TxlF411RioIiuEUBLVaGwwPse+iV7ARav1i8C5fzH2tWKCpGfAu7koipwHumzu9Cn4pDcS/S
fJFsLZ90hMAe+1mUOW6O/OSRe7R4sVnfUi9hp8hHn2QRKh7Bsnf/YHttCLflDumNte1JaZibaRGF
b1YYX/hSk6LRFY5W5wUrdOMAvzTbkiZT0A6Ysb/iXB2VnOlbSvJZCIy5LZ82JypbeFHX8Et9p6rP
rwxLCNkYVTCJyvt+z2zVsqhMNGi0LoQqbPTgMKE28Y2s/l1zVl5ldGyHLAoNPKEwlwz5Tux1vIHy
MohuVWw14xjJiRCPw7h8zm4z+tI9mB0miiz+GYVKbW2evgbVoe2gs76SdolV1LKoaKBMlBFuY593
1cS2ibSkUzs2UYk/9kzbqYfYR25xdotbLs2tw0Awyb0nWBkeoxPlPP/PDm+0ZGMB3WTW2ZXxxPKL
Cctw5Xo55k1vhVCV9A2GpBjQTB9HYOyN3XhZiNVls1c88T2E4pRY1GpRIWhBQ5KT/xQ5n+Nqu5Ov
x9Ddt3/pqjZrNUT+S87crwb8nSPD9vAH+SggPczqL5YDysZAIGPwbVpCy4NQ4ed4r8UEYtOBQeAz
n9Mac51Kgv4+C3b+14F8BtvsLMrA5n/FzTXejfxWgwH7FRLobqW5K3KfIUF9LorYFzEPGArHQAq4
sb2EkKB8R29igvv12D0gvx3hELdA9KEFReU4Ao/LUE61jLPqSgZG7qSRz4Ve+kxvcSworlkl700V
1oUBm3PmqSBchnvl1GIGnfLVUjZQWbkBaq1Hhu+TAIUwLQT9tB2GQF349ofqfs/wEpmqaqK/yntp
5pQpwVgQSYudUPGPqiPuJDxZT5pZywrTby9hvbWaR3GyOan5Ycm95ttZjkz3uJm2Jswic/oivjQ8
senDrw10b5VzeuLbjblfhKu4mVm1eWuG7U21xYe48t6H2qDicZVE2c3NGx/zF3UfS4OZtFbfYe1v
nWTuoIwScpzPORwntlS1hZFjBaP74hRxjuZy5ajpNzOyqdZ4ZNtsRZJHevZDl2RVmFmX8H+PbANa
5DOrQQotkihlTpvOOZnFK60NCvkkzVIerWNCJGewz9nBZGHRN/tRs08h4V2hs9Ek0LVB11hYOjKT
t9RP7hQOK//RsUEeJg4Uxsg7pH1T29kGiLtKhj7kdgVRJdkmDEbldd7TNVqnZ4M2gl1gxORXk4xA
WR6yQ8zuDGmCeaILH7rONrQOiQTLFfmK1DBUyZdOd2V4Os9yGMZSUevX/gtJHVcNrYBsbG9dNmSu
9MCE4l9emMeNOdXXaRU5ZBhpo5wCQ5StrRMClTRtTs9haaqMZLsVOHUdcCsC0MefR1j5LjBu796S
xKsquop5SZ/NMFwtBA+a1PvnJgeQlxZB+qkwIyno+gwu0xUUGTd9bK79tcUmK/xdbkSnqbkwQFpx
NbavExkmMXJ+ZXN4aSU0y1Ubb9v1XcAXDzWdb9xzOF2S0AgGdDEd8ibfDfCBV0g3vWuiqPBww7UK
gCKWwk60FuhalK7kWMFmmKm3KacDbIGKqW3HaL4M+q99QYLCvNKjHx6VoCx9BGgqUdblAfLYTqEf
wmMUJAk0vECKD4F6X3b65RjmeT06Tn46oomG4EHesBXnEYeH5eaoKU1ykVbIG8ItxpMQoA7IrBn1
ZhFDZjUjOSylr8glYVbXzAddetrKxmIDk50TqSaSEQdOIE66JsCIAplJXyRoO/rXG6JHR1CqecCU
QnrEVV2kBSLV4DP7hAXupLlGncWUEiBoDBai7ZaBjiEECA5sacFphkPogCDCr4u6vKeQ5njC5oVw
HAHwCz7Vz4Sznb+mWqfsVD+mjbNS+P/EEqgXm3xLaWwig1surNSeANAHBiFncJQQhGgbOUfDOJmN
4op+KDB29V/M0/csgbQpVR7b6qhA1iU9JqzpeOtS2mkG6E0DZ7DsYIsOd0Tr/yiETOS6Qq1evruz
9O/qp8U/ty5xxZ6oIAiEDGOaS3MzCOy2QRPYnsonSsUlBp/4YoFegAnobYUqg/Ntso4TgAF1BXlO
gXCskao0e+hQyVOkTNjkip1IYmtWKqG5FojvYhGBO6mdW0W59enUM6Q4DMreK9khUdxpq3p6TcdW
FZU3p+vp7VFlF0jFZzT3RnWnushJCb1nP3ikx3jb5FG6YNxEFHduG/IE6zhiCBBLo09wZhgKzRxy
k1fITE263dsR4BqHDcaCL1ShvdVxn01WjF35IFoSIDGuGq82hy9jH5MRHh1wrUG0EOmJuC5HmH4y
dus5jrx5LwCZTXnJvDGabu+BtsmjzSmb4MwCmOyAGE/AkZlhjBYocxCXp1FSY121/NiDWKPs5CbF
1lTvS0vL3A7SnoSjCwiK+7NPY30nKVCFs8gR3L87Yz1k3rAKo+6VYrumIukY1Xm0py+a9tnFQ0zh
56/NkvOJyA2V4lbb23oujg08DizZCjsOkNf7dbEz/Ce/JD2AkN68/XX50UcbTu2ooW3ROFOt2Hor
8PKgLfssgphGP7S6FPq9LXfdprM0fpYxUiLZ2kd955fpVGFv5gN2vLbd41UtfqIQhOGzZcd5DnMs
ZV17iGinAgYAOMrDOCShZtWclPuEz2BdrDHaCy05pdOMtma4qSrgT3FFqSa9tK8WZAo69pVgTAv3
HNyaHK5hDAgINX96ICfGEI3E2XP30Ls1nqERxE6oUMaFDeivvb5+LyBY92UhuUZ99M2MviMvfB1/
Q3Y+qWUdDgbxp0/suAZK1m6Fdxou7Ti8mWsZWYEp/gVNzf+cWP7djAciGliJLRY4lwzBcg2wh1sH
022SUlAXUKDTuesIPDNe33HVBUU/vx4P28IyCx+pfXUjwbbRlWZYIJZhXtANphNwdM2tsLX4P5iE
2HVZJCMJXjUBMV2SnZv1TNVTnPzRJWNevCJqHhfp6ObvK/y1fy4DaRFVyWjNLM1OyR06GTklY9sU
k+tWPOTSNSjCeDvi5MM89gPiTChv5DhI+gs813SS4KGOUq0LwYQV3PSJz/5oR+hRUyC1c8CLY5I9
9J24ReUuOhZWGHKdCHGFdji2ragWVVtGilhMakRcHRlvk9aHSVoqhZ2IWQEFm9eliHZ8JNXvv9Db
RKPgugLwzF0LaFc8NOzpeGaI3iqiwMMYriXrrLR3T58loxYFpFAQqinDHz7gAo1ydzwNkJH4hZL5
KfaMCxQxrUQK4j/7JdX9WGAouzdjk3Qb+AeUD2bdqmjarn81IyNIW9prywwCBPdHY+FcXo71QCO0
ziuuiZQKllWjSV8/nr6WESdvKUpWOoq6as2eWwCl9PbECCcU3B7la3ZXLYAia74hezZUEXs//yjn
Ik6IUQZHSycjjd5Y+3rEWGN3yKesj0lYKiW1qqnHmN+zFpof2GCoSE85psnli7MZrqUTVYznKi9d
Vhr0e0nGYHfBclvLUQixem5GBZY2aAcRNXMDWF/5OyhpE9kWwNWDfHVighX3h3vE94ZWQALul96I
wpZLeIlBq7bLlcc2J6B0DZm4P0C6DFYb3LmSAbI48gt9TZKMbLGQz2CIfGPERBwXkcKL+e5nbXlF
YMzKtQ8GlfCPCmqD1hyN3ye4BzxOI7cX455zY+YtHFSBqwo1kTSTT4tUr96/G0d8pK2U6pZWpIbB
EHT1mFtJfLaIJIfMO8i9yopO6D2cng4SKHnGQmYt0syWec8iixR5x8FbM0D3hCATszgW8WE3H6Xs
f/WoQk76OD6lsPXyRlhcOpJ92Sfo5mF3S67Pdx8IC8At8YNbJ2dcZpvxgrRJBNRWiWkkbxgKiCQ4
MHEV/XV5UIis1mBU60rYjQy7TUf+Bf6ZN0YXCULGkTJSqNQRYfcOM2VpO2OXg3LqGTLkYJvH9lJa
pbRyBKX88gdsJopMo4lXGbUo3H+jBJh4UUhM9NTm6/2JEKAoUM2EBDmKeErprW5vZZVVRZzYC9Zi
q7T1Am1yRn5xvDzmLAdA0zBOrZcr7DTl0l3qcjrOoR38S/JyjZfzl7I6Xfm50tmsuRDJ0CP5HtZI
2ajUU6Ix0xWbsis4CkQ88O059wQLsuliybJgB7/1cOj98lnQNnNoZh850kAI/IFkYQfNBeHJh3uV
xIIk8PVVJU/WFOHUbyQ78TIIPr2YpZuoyRdO9BOSiaYJITafQ9KvpXU3Do5N7Q/6K2FAg3thDgjg
cA1le8bUB4hXHfFuTkcLJ5akZgj3xDL2POX8KMUE79UhnmLWtNBnDfGeTSyEAoGxDuicBKFQD0tD
UbS78j94e4icMMonOibcGM+HP+pnCGBZAK8o7LlCczxJhFVKGeoSa8Kjeq5EmU9ciSkKaO47xmDl
HBWvlpS1CmH7U7uAVsN4y4CbiuYiNyyXHofEoCnYLrpqwpslxBm5g22gI1AVug7DlKVXfnyPAPpW
gk0LuDWPGp1NuVUZ7Dj7KmWFOJnPcq79Lo9UjeL+jA/fzuSDvywgUi0eAuxinj7g5ZNxkhxo3mcZ
Fb4ZWoC3u0MyqZwvlr1kjdXIrcnXunkEKCC7yKghNegC+ZkIkQ187FZhwlj0fXXrESgVNKuzWeRZ
6r7qnqnuTwquFioRsrenZhEtuXQtFI9M985fbjhBiwy5cDt7zfXlKEXDgSKG4pK4fnE/3LHNl22x
nN16suBQwaOo1+q/OiwdSPl0ZZKQ5/mvg/vziQlppHieiQwjyTtQWBDjtJAGqS9uzqAIpSPpVFkQ
+jlsqY7sxw+5a6y+vamDmdr4AmHHPH7EjiYLptTPltTq5m0QlHIaD3WQDpXcyv6sAm+/SkdsYzZM
X2Fon5gRT5BXVoSOu9N4TLAXu85scRCzzleBdCK9vbBLUqAVJYvmj3FHsRXLCUPvMxFd/VigdwfS
WnWwokcPl0vLMtEwAegtKv9Z9hWZyBrE2ZnLLZV3vMbxLWoIyL/xghPLhYUmFv1wMcteE7iaN6ND
qavc9gD2NcFJcsvgAHV6Zar9qlWjQ5MZmW62u8ltNnj7xuSsNgq2uqHLs8AMHe17gHLc75MBNRun
MEk4ISHzTF83lZfeyEsaYC70jTemtcaccT0kP7G+blKPlMj7NAOVTTiaVhfZMBvUZMJRNv6WLNVa
4SOouO/oxd45vkvgtj1KdCwoDT0X6BQxov3K8XRVSQ5FSCviWzcYx0TF6cOl8gcN5AJFFrdITff+
RlOHsyoAMm30npdWzYvQ4CJzq56HUtAvLGD4w+SwMqGMhGvbKhZvcr/VyhtMBze9HGI19uVzvh3R
odDLPvc09+5NN2PQycQ7ieckxQQx8MZlxGowvVpgLsORR5+qzZq+JPOuOPjeWMQK5QCPBOEUwWRn
eTK/ykJZm1mbzBxH46LlK/AqP2d0lzvZVVRO9x5lnQcI+EikbbSadM/2ZeRn44Yv5cG8ENykCrT2
cj0UWS6zIoFthxNT+X/yOWbqJZURmjuCQdQ7lMk//eKzszJ2BbUE8D8/ZxpSVMbcElNTtSzqRQcq
EarXPUST/RApcmopmhmHuxgk6PzcTooYw0EmzngapF17gXWxzlB0BAmFe9ra1fT2JLUz3CCzkPZU
qbb6745vltIyMyHdZuNns39Am5EVzGOSA/Nfnhoug5+8YUrQhd1Wprm34i8u9xKVK9C5yeBk1Vfx
tUC1MDbZ+9hzrXzGJZ6lyntCLm1AICHfnkIyrqgtvII2X29EJEaGppzz/Dr6r781QPPlEkcKJ2WZ
cXUWNo/HSH+9SaPdgTWzRadp1gqmmbGVcSIui4By2PQQ+PWJLn6jLJbL9ACA3VtpUKJoHzyeQhzZ
mKL7W0o1xj/YVmUT2Mwf2MEQYNVZ9jsKZH4wH0S0JhkP9j0zJguvTMiF8kNNaSeYgko1LnBeoMsZ
s7/zFuNxRk7nhs110N9+s+MEmsb9RErwgz8EsCd57QCySACtEI6QSzHr/4/tm6OJcjOhYn89ak7G
xSvfwc01KwfIm2Fhy7qC//rf0AnZSnUW4Xv9pAxZ2Uf5O4DShT4ZIMIDpJC41+TOPG71IZBWuw8x
RvfSBnq1F8rsb+uJuKYyQlSDQj/91wVt4ptuWpWNCWEuDb2nsPg9NRWHAI4MS351j0VsMx2Jz1vP
Gz6cZlRd/kSexjk4FiorTj4uwt/Tl5Zo2+w65eRo6m5x/Kb3FAtG10hRx/WX1pIKerGVubDyGCM4
y2prOMjn47aJYyslLNRvkrU2YwGR2nShVkHdkx1ibyFkUKjf+YqK6HBjxbOiqYLrUY6aGMwJDf0h
m6iaJWLFogzZN+vD6TPx6L1SesDa3qJpmGFWJB1VEWRIUZz/iwp+49Vg2dQk8cICXDshfeHkOXKw
kvtHmXX3LsEpiWkz03p4y8mkCOX82agUJ/753iabK72crsHHX51QKWLLedNpuvOHj4kMmeMJ15UW
zxPP3au9t/yCLpXPuvLZmSTrsauA/9NEzfsks8nKsgjByH0oFESJRB3MYDtIlbia0nOP1VUyVut1
pK5q4mdxcsz3pt2sY6DHcZcIxa8g7T2220YyPEG/wEUKE/NPXRyTaI35mB/oHQQtuqdt6sbDl5BV
sts6sDJPA+QR/n6x5C/H+XCRIF+Xhvqg/UZsSrr/BRJMsoW8lH07g8hdI8Qpqf/52nBBw87aOORQ
be3U8mq/H0trkM+oJyqGL0v6/8L5REEbBXWkQBv5J9w/Aj8+d4EF856jwtA27r3yQcx7q3cSk5vS
LE3Wfg9Qezq1ioiCBPS+aYIa57fL7/5c+7OoA2uIlNoTZUWI/ZAeskzgv+e+P164+ppfF3lDGZ64
zjzaIShwx9u3O1NopYxVk6ZUV8u7kQocTO1LCd8rDs3CCHNWYHVtFHbp96JQgZp+DVG96URYZRSZ
PVGXJdAs60N8K47B8+DWUMgJ9EaYFEtabuYQoUhsSAK9xGbc+Bwl6Tag5XHqWJindsClozbTI0i0
ySnGtDOr2ZKICMq0CVR0LgTtxVdHIiuoXxm2xA2314DVK+JYPLfCXehAQsSvASPbvZmY4mSChSnq
KYpFMJGuUg1shLLfI92Uq5Camfo5YHrQh7Q7vIhjYQKsHc5lFn8uz8WtVsLmb+v+OZd1v2ZpasyR
oWwtg6s7Y6mXbdaTasZFFbrzjZKDGjarZh+6so3BIQM0UHQ1U93KE96P6tibUakSE4V/v/bJ/tGU
bc7XPEQrD81u9bQwpe/Lfr6JIYP0eJxLTyQ81ZL+UlHR1cN9mt+5bnS/wr0Kk3jqyjf8btlGniA1
QUi6DEGIysgFFQfShjEWF3G3fXZWfptLjYvBH9tLCmv43ODUQgMJ5AISobnwsrPGZWyN1uD01DUc
S8gu/3lb2q7XE1/WQKp8aElGL7GDFtbi4yWsFXHsOW97CjtGhDN9IC0qcGgtyCfvw6K7pB3ap7cb
SLrN7yDIsQe4JCnPNDTcCb+yoQnSDsGchyhbHeg0PA89SNWI2CX3WjH8cSkdbnNjIipcQFnUcvje
ZTh44glhx4fYoQ6NoeKL0k58/kBXV9CnWCAjsYqSw+DIEJ2yrAhT3NdWZ+0KgC+MGK4zC4GS2IN/
gacZeQ/djLFCt+PQnIHPvsrZAp8gY03V0NuRmJsDxJf5nJUc+lxRkEu+uo9iA4jmOmuIrPQIbhST
K9fPlsy2WBWVMobhQKsdrx+ge/vJro3nQDnXcxM5d6Bg2MUUfr5yDDdEF79xhSUchjQVar1MKgac
90quau/bdTlLC4jBXCGxG8Rgc00nrj0LD/l7XwnoqLXtVEOc0umnb5N2fjcEMIopD0K8PMX0GLZZ
R2v9oOw7hVdM8vJ78KrEiV18g675S0SddDckBOPMAKj3Ni2zu4Bgk/jBjMXgQ0khlpWEKpTtj7xI
dovc7Ymln6vwGu0Mz5Krm8qoBm71Br3y+na7lNxjvx0A3oQWxPH406C7perZKquFG3lmMP54eicn
qm1SftmAlrEflrXW7fTfx1t9Py4/7UouBdnzivjvCxwvnEnkDGVlKahd4qEzUz+40UDboMEGUk7q
E2QURs6+0QDfoAz2uDttLAnGYqqvx8ddkRHbCCwToxwI3p0uVW15xt/dtZ69cbfvL3v49U2tnWWp
NwFFGKbikkf3rWkipsD4psCKCbRUdz/XwHuqfLz5pW8uLnBzbhKvpmGrVScDeA8DU3LT5QZHFe3a
jPyQfwlyRg4w7a7Kp3hwmX5SztQhR9q0uk8gusrkJQ2wXHXzPYCc4Uo3CRm3KjPKzaqL7EwhDYtR
HIp3wy/8evnoEBQQc99YKofC7CdbumXP0pvqrkd/uxXhw8G58hiuYTgJRGRj6IWOm49ku6moeijT
hIE/wERHEa5GNPqBjg28rp/WxYNcaGx8QZNQcPpRSgu3VROMDjA7vuyWkfVey+10N+o6oGExEIDk
hEPv/B2E99RboLbEVK07EhDuCA16BqoHU87dNEnl48dH/QQpd+Ih9DIjUsHyAAS0oYxnmqAcePHM
gHGoifyTlRzt73FOmFyYsylSL5CyVKPuRl0UZwlAMh0JSCDMO6WirpDsV0jcUlHZDtY3z4iG07g5
SSSP6EkJEKbPE/ARq5/IQt1LR3QB/juS5vI91x+nDcZxP3AP75mJPqcFis6jC5idtTedylsie+wD
0DMgf7ztHWt+/8b9DZ3KumOtsw70SgekDr5q6vrh2Rq1DSeSGoCY7Akx5wEnrAs8/zpdcxoSYPyB
w0DlFegofhulTqpHCu9WyJbWJcdUPjW32b7JnQKIqZZVkaasT+fNGl5K4rgTCtxLTzANNy/Yd4II
jq/7JwM78I2ewrj3pUDe6qD56gD3nW8ylCHMieKMi3fohwrLepgnMXuaaYs4bplD6UeBh7t45TsS
LgfjghtfB24+YYe0d8tbizSawHVeRf9DWugHhhQF7FCUJvt+Sf3eTysqU22esuKzD5tuOVERM5L1
BNkl/ukla3nloiWZJZIcy/kd1jGU8whmgZTcA260OxEAOvwzN+Ainx/HQtgD9H5Fw4S0KR5VC0vF
EJJpJI8qd8S0k+lhblSshx3l0qnfKsBcESA+kMRPBILeDD9eFyLqdn1lBm+3y/Frv3NWLM4CJpER
LHxj42jtzdFHVGfb648D066X4zUyg8GgaymPAEtGEaiIRzx5Th0EBbz6G96vLgoFE+5E/jJDV3rO
RCm9plR3++qa0hM+JU1jhsIuuSCP6yfbM0N2hfRfWGF6w9tel/gd+juWaai0Ug5F3uUBGYt9dLFL
7h5Yfm9dmSoecWrowculT1I4tlZYpnfacMWJx5J7Q5+1w+Qqfszb8VDN0vjdXkYkJ8BcZ1BVq/nQ
m6lY3ku+uzTgousqRIJ9jglRKE4ftk0rqkzEKe/IvVBV/VXWNBVuJHvWYg3DqnaPEh7UqJqnaPuX
2ONwuq90cY0q91OiAXwmJlVUQPwY+znasib1TGTr4hYklXzavRMqA7ijfblHuDmiCElGCxgAC21e
sje7IIj11CuEAU/XqBR0hCsH89BCe0ugQ/otIPOtFWAL4m1HDvoMLy2STDFd73/WmFhMw57e317W
BE+0msYsGTRQVn63V9CWKHsGjSkkSIvZXnKUNuu1OqMUtyCVaSOh7QJ+IY2/wFRZvQ2KQOud0E5d
FKnCkDNUHy1Og2h4bdGFiImxF7l3E+UBLmyxfm/+hCxHEtwVOP/UgofUdEEVOYR2MK3kkUx8/dT8
i2EJTYrRT5r/AzWDrB5pb+O6utfRU53fe6a3VQ2qMLdlU4AilAz8HRYY5vwP7NVbpTjW5v96SqLj
EVC2Bzb/3JzWzs0A3RImX+Zuuj14rRHIgWO4nqFyEz2zYlzCrHVATl6PFf7PlQQJsalQ5JVmMYjX
GSgnyRV1X9CRlJGpwzLvrQNJ3DReDQm/DTFXytaTj+iCB2FZezc+sOr24AdVCi5fbx3N64aKGLXP
on/GGiUe9fyJCLrBPnh8vv8jafNX8yiv6kWisOq5mv8Ffy6MwCIXAv8sq4sYzkPqps4LBS0FtH+5
7L/DtpwlsX5R/ck5WtCHdv7n7cE+bf9v4S/etf26a6LE5XcPJTVA+BHZc0SDlbkS7ZvkBFtLGw7e
eFdov5SbPDnFw8jOHCOaH68HA/RBCxKLDF/YZS3fKCPSqgdvZCWi+4LnS7F8GVSBRe87MSk73aqA
dzyrJKtaAxfhWwj9tWTjCQ0YIox6QvuUBeCxb0qrWpXAXC9iY822ijzL0latwLz9mQ/VVZTLIx8d
aLUYLR/sOapxQiXmz8qGoCiDkcD5r5FXK0nVfuzy3EAyYY8nRHNWJolMOI6WXrRfu/RGWOBisJCm
sPq9qI3Kq0Ba3kdSbz8+HHyZxnBNa3zbrmpFjDjFoUHPeSQIcsokxE1/BUN0aW4eNMf6957JMac1
s5Y7c6vqGoVDZ3D+rr1kXKkQfhR8NWLia/Owp6/C7/Dc32+Gqidw1ZCOcDtvpXt5c7BIl01AqjbQ
ebsLQhzQwaMfT3PcyeKEWQ8l1K0gHqe5u7P943GwwX7jgoP+6K2aduleHYy8gWIC6swEHOxjlvoI
jc5PlqMJdSkoIWzTEmgQkNJkMQboNdC24ZZJSUiJD5Ci7Csieslu8mFyumrEb8abXchIET1DfC8u
w0szwkeMOIomEYkziu2PPNlbWqJhXhH3Nf8qmOizRnJhMvk0oI8JDYUKCcYBYmV3Lcp2AySdTuK0
japkMeVV6QHgv7pFowYRNwDZe3oHP789pUBZopzFl0loMxXZ4dfu1J78aZwKLW+vnP4+3rY9XjZL
QsR0BLG/+nHJNPqIxZtdyt8mNdj6FkQm4bC2c8s0Nomy3W10p5fnAg6w6l6KoFoMEdbhX8sCU8r3
lIvmQIaFk2j8Mq8jz282BDSZCk5z/HOPiC9GMKlKkyJvNi8P28Eo3N8O1F8S4eVc1vY0Rm9HgIiT
Tae/CgaiFZnolm1/oKt9znwNp497UPP3mVVXQR5iy/YQtVdHk7rJ1xZXhVH9MyHyLzt7ufFOp5YU
I1v2s7+pvNX4qqQgzV/Tm/WszBNRW8wVQk5AsbWN+4VBfVlJMkre3Owiu3NFzRG8aRunVyTzzc4n
li+vlN7BJWGiwiCTwQfXUhiOrsLn/JBJAbsLq1xKKd+NRG9wF1AO3gIt2ahDOyyRsy2Lif1rsJg0
LwZDAoAZgg8hpOOjqVWN/pHIMhqaWDnKxMVcLEQ34zFWZ2s2/UpnASnNvXJO8j58O9h1SUISxf/o
LFC3LtD8tnBF1tCHE/rq5wxeGfbBBCcyyoHFVk1+I9I3onSTRIeyxcHk50qyeYSq7UWN0ZND1C7G
8tNEATEPruo2h1IF7C0UY0PVuQ4Aj2/FNf3dP3vta/1TRAsYhBRMT20Kv2bcyR5Lwmv+GH/I8QzZ
zMtNBAGA2ALJpPbnyFzcCM7ft87Uine+SZzoGU6izbrIkatPILA2Et4M/LJwWMnBL7sgEli7du4U
zkilcnaRTKKMnc+MlgE1tAt6Itvdzgv8034YN8F1ZnMfWEFbjRXxiyEGgybmg/75KIT6YuSlU5P6
rJJrf7JZmPZjNJhjEfTpEQr+bL2gfKGx1EZSlAGwMDWA4uFRJuOjwXpCslzSWr/v+S1SZPXrjlxt
HvYHwL+jqjzQVydi5ci5KZasE/U9pDv3GUAbkAVrvbHc5pznc/TgRIc2wBWOB2uRYncLPdpwjP+g
8kNSe9pSa6uZggjmNjrcV6KaNjMdSig0rzoIC4y8UxC19WjOFUVMXvplp6iE3wY2+9Ewg2y6BJ5e
nnZAlaRJDa8fe+7ox6dEBckffqxBLi2oQaC4GN+tP4egF6jT0p4epBqwacDCysa+CTyq9x4WwTFl
oirZKDo+AhVMYMqrWydqkjCiz7Dwdzzr0lFUslcE2wfdZbRapCxOuAyRT+rLqy0knWCFCszZo45k
RlLIzN59mKKlzXf/8P92V45Mcm6JN4GNAyA1Vy6oKEv5Ve2iI4hDAP/EUOvL9sJCsQy4BW1dnFuG
kmKx2FENNUIvmdRnkIohrL8xqQl1220ZSvnJt6L0Np1v/KkYmVHkzdyWOe6+dvOBxUw/Z3TcCfob
uU34QF+9YLD8YLnty6C+Y5DDh4p/NbcDzdLAjYu9KL7tn7MW/EO28KmyqzkxvAaAXrKKFua7C94+
36KjFM/X4MOme4v+bJbYtJMzSkYDAJmJar6ZCzqwmf+K34+zrCszJRBtmJyUCHrbGJO/kD9F3Ooy
V/Q4tmtc1dwskKARLoklVr3rpX803tpE4kfe3WAbo5+bCTR9rgRXR0batrDf4SmT9YTULqNRCBWL
Z/n2b2q0IZ1kpt5jhFQuYWm4nkhvKMhtljJYqtyGA6GxE1XXCu6yJDiqlhfF52jt8I0vsn29Tz03
NaInHt2zegZoklJO1gz2OtSGhJz2f1HvtyT6GYDONRjRSPu3vfPEwKkwf2P7m5rAtGIf6dXVLYbP
kkEQCEnAipNnELV8KnHQUK7+r/PJ6qV4swG7XKOu2nbCcMwsqM1mVm0kgtP+2kzfjVcftVIsViI3
XMRRg1lvtnVqWC7gh2XPHDWLyeSZBYhto/8e0sem/ezROo3PKY//xO8hHYPg7Jir5ECKa9FVLsD9
TXgyQR+hCV7ux9PC9H1zLHYx0KCiFy70ufIsYirPRTwTsOFF32ar1sw2eEkCwTF5lOEqfeLQxhQY
gFkqJiIk/FYUWPpvagw2B3RwtLDIwwzydrzOo9Q+COfJjNr9xbZ0Ox9n/5ZGAjpU3M5f8ILYhePB
IzHTlfCY6GNL+QlJLrakFsKODqq65h1OM9f9Uu+b3V7m+ZMs5EXaHae5Ia0b2Zyu1L4m96f5HUr7
9TeVUkvICcklsKSt0ZOMd+t0EkQtgLg/00oszQ/ekcPDvopvDq/zIcfyzyjd8F9iJjl99muouQ9J
HNj6E7wRmyE06MO9SMfURiwuoWgpC+tKVoVZRWSf3E29XW8t7nd84PEinymRbZN7RWBUcnd/nTBD
DvTohNRF59BaBbDPlF0bPlQoL9EMLZsXqpIgFJ4YJPCMqNXrKWsJ+rS/njhw8qsGLjpymxyub7fE
Tt8X60hsudW+9kpjcAsv6yi/F/LnXAczRMFELQiDXKkZtqxZZYvrOgqnMHuNPeYeL6tj18kKVfFq
RmXvtlPKZRXKmdGeKJ5I5VekkKOuaWYNDBCQDkQK7ksQuBITU6nfdVwGoOQ2NJYqnQLJeEaIPmi+
91n4ei6TLzsO8XrLYadVMlTuGnorleFR7wt5eVNzpuIC6hgD1DHkiV/PU0vswG0c5uke7Hb/iqS0
q92yQv2uF65jK8OpAdAu28su4XUWZHsLUDVqJmNO/2/p9nfzlCB2yx5fi/O88opfhTUxrSKga1hd
/Uoz+viSyQrXAsrUOM+HPqcIMX4utfabQPZlEW+ikuOzEmbtvWaf9B5z+cZ1WBc17KbnH43MESrh
Iizbglan1lUpQeIyWQQFwoG3FglbS0eN+8qM2ppBb0jdhvqxDHhCXA7w6VCx4I+Yl9h6jdoxSm3c
GZKphp1ZndNArN+vr5oz5ZeEEV5G/CskC6Gm/AQWqPRGU+3be0ICIVbG6FmOe0/BfaHaq8IBkqhI
bh+uv2uycnWuKZzoJ0pPej82WkmqII0Yo47uHzNaq6UKOOhKpgHaHDsunfcQp7Fr1Rgm1ymxBZPm
HSMFXBVVnKzoAjnrnp4eMJqmEkqiSnrjgEIdwaxLeI8Mh/7CtWznH+mgE9UIqGodEE+BEAzXxxZy
3jJmN5yOUQDix2nlMopjzxZ+8gwWwzn6Vj5dfTC8eZ4w12MLgaxBpqo72N+xeuWAtTAmPYlWm9pD
EtOoDN//byYG8rZdUbwrbScKz66EExZ4WyvSdFw3H4qsZrDmGmmbjBJ36Ms3OIjq3yfAlpuQ7TI0
DGDGedU/GP8VxeIdCX/gyFsXK6ZCBzI1leXZ5AMHMmJ2hJ5HTW9qfic6fWwrwBAlVfdeiZwSLdrq
ewm7fSM4mbmnT9xR4UrzpFGn02KtSqSQR20ZMyMI9XYQsVTfBrjbBkJcKSZaRBiqfO83c9BoBcuv
QsbdAum6Aj/4E7F92FpYVqZ5CfUGesuqFvIHLfmj0MlxmdVG0rXCFCzQXuo3LZ3QbTzq/gcP0Ag6
hlyucse5KhVXBKLHB5ePVLVlIEPWzF+8og2pECxR6i7psacn4pAilPcu4oTGMAp/kAN1Xq7Ra2BA
Kh5Lp/Et7IXTWgBoPajT9ackajU3s50o/sNy18LGBF1rCtsj5v67XD0JhCi3mn8VUf99Qy1ML8Ti
uubc7bzSn2f0o6W4mugic2QmerdaD1urd3YE7evzVfB3MbjFi6V5UJLW8iNba9E0O8HkYPpOnM7e
0ZpnRYJH8ixBnO3A2e2b4dcm0mk5Kyehh0kG0rkAfl4pluEpJEk/WXO+7ie+dn9nXsxM782G583+
AVJhi/9GlqxOSKz1omhNWKEKbITi1wBhEe+uptXrpJfwXwJd8Onk5BaUNeK/i1D9e76KWyw20AJb
pxhEOQ7rU++6gBnBoJp9CDivc1mxHcxQhShhT4w96ZpsWPWRR2AAO0DxgC3X+PEoWKgwH+GRJDd7
QOuzW3h6eDohjKzZ1w3jq7ZY8zIc+0jPqcEP+Pf2SD8xhNRgbyXyLGsmfwbnLdqZFniSwVd/b9mB
zL35hMU2h82/sQOjfhYKSq15va+qWwfTQu82qrOmMLvJCyw9egXSTvp3z8ej48NWBv7rXtiQTwBM
Vi8rAYPOr2TWm7lechwdjnlhJ0jNkXlqGAyrMHN+qRtR/pRw5f9LYzks2A44+cSw7WdjgES2AtnA
bc2aVUxeJDK8z64AYJPy0UHEMIz1gNNCfRZYLTg9I7lO3/Gh5ad3EEanMPwqfCKaDp3/oKRtBOve
XWPte82IrXCMQuXt30ubKA+PAXWcyULVAAgqtQvpozhRCFBqlKnCu8/cf9wFJe/DBnf+vTIPzxl4
XGfGjClhXR3aFUxLA/+pfokhyhVPWCqPLUGeBILeu9YT+kjEA2y6D7MTc0RJ3MsbNpoVPQ+92d2+
dFO0acPuQdCgTZlx8v28uIOQ22GeUrr6JGju1lQ1C+D+t8NhNm8N28fx6eNmhzKIztTvDcxd9aiM
U+N9h7cNwwK+pATwPl6sDTxn4N4BE78pmSIZLcgLm6r+O/17jPpGnva/KNw4WRhHkLxqayYnTPby
TUhE7ev8UELnswv6vZFYDUezSzuwO/T74sueqoAltnY8OfhOxGaaz66UZqwfIQOeA6q1dm6eGSPX
M6yG2LBmVWwqIzkrm01b8+s4qKL8l5I32TAuZaTl/vnlJgDWArh7hZyLqmEqrRcLJTUzrwsY+009
ohJycww/pDSTToKws0KZmH6rI2Kiu8ObM5xcB8KqHhW5NgUQjk6QCkc24oMXJz5aS9hgnD+PWSCU
7d18+E/ahBSw2tP5HJ3B/EifaLFkIFoK4gd+5H+4XqQFApT4w/k5/YNsquqogAsGwbqd5aGjQU7T
HVWh1PQNs+aPbTJgv7WYq+HMrWWO9gClMjjNWGWZFN5XCdM0PHFvPwQydwolFulx475CPHJoV+Pb
3d15cfvnSXKzOIUDUfekUfIJ6iP7KgKPn+QWBE0yOjfu4ZPvdi0nBkaIbH/LEhqX91P2DYPSRVyl
85Yyrfsa8HpZUPQes4dvpZyCDBy6j21gL5F8h01yU0p0/Z/4EAct64WY5E+EzhBXuMyIK+bzO2m3
CVggp9Ot69M1D8ywYLmas4TdO5M9Cu93yI9N0UlHayEEzS1VUclAxOFMfthHWosI01uREEHEm9YZ
DGwNI5hZuQYJc00+zauR+AiAt6Jy3+LzRAY9K8BIVJzoFC6po1+4bF48yNR9LZdh77M2n+W8PB39
7qAMMRm3OWdIsA8YRWjw9dOUCeIYj2hW1fu3v86nsb3jchcUptagTr68kUlRPRfq4ksecWSaBgts
ke6iKNd7XcxNqMsAuaTSlr29iaex5/gTrqD8RJ0hS6uAHyp2FMd2asEArgB1h4k25kKcyhkC3LSy
CeVeI8jJCRNVK8XQB9nt896DKIR+diPoEaxQfHjr0lCr7fd3KKu2V+iIjbldE5lUZRY6V13L9LEP
xaT9QD5IZXh+Exr2WEEerQrdjtPQ/AL9M34vo2tahT6OpvnZz11S4X3In7LEodsJqScuJNqIheTb
aZ2WLDJNeGbab4Qt9AMlVI2I6qgDHt1EHE8yobazpym/jARy4CHFU1f/9CsaFrtbXSnxftAFWChZ
nYgOD7iwYsKV5SG02zlNzqFbxG4kdvDKLh9eS4drFywEljjuS2de73A/Ygz+W1vyd/iKYx6pW+NU
oOid60bjvPaVWAw6EonHo2Z0W32tAzcYUWwQgHry30vrQAqECSY46Gu2Pi9MRQn04hhsHaUoZSws
GcN78wSIqAC12dlUSJziPGC6riJtA+QCV1/vgqr7wu/wdlC2VIgFmhA2sSU6SCjk7mmBngsjTWvE
slIri3d1b08p6V5DmZm0YqVEPDZVGiu+fXpKCTV2mLSeeCYcNJQ8HUX3vJx+5LxgXQvQk66lgNgX
S7jcN34iUulYvwLQK4r7gXIhHKG59eDiinX34dmkKntCktTJGWX6JwSruAGtpGTbbhLvG51W/Fuu
P7qlfPGJgomiCuLt6gi+rp6z8SRdQTBibgbEHB+YCniWBbTyp8qiNe3nLgcrQO0VBjwPJGcbOAzZ
X4IFM1k4m4+YzoXNs3JGB9UDIO1kMYL9NTvnR9EbO9MJafJakH5lQzd1b37FVkRZTb3bL5suFPS/
OwJIKE3ewNve9yC8Jd3yvwJZ8GWiOUI7t11zGWxWjo+espilyxfZ4P5tmoKkUgrXHYWExOthHq+e
Ba+GygR+HFhLUUr3NwNzDsGGAxhGEPTjfyrClOyO4SfqET6ApyOIqK8GAGJgQHpKvrJFyAGhQGel
jHz2ZjS1dpwZnrbSW+DX4kp3aRdUjGhb31vxPptnutmh82UqLAtwAoqzf/O37I5mZKzNN804CkSM
TjHFOdrGVTZunthsAxDPjK09Vj/kn5tAqmoDpHXJ0/CvoH7thowsPRV23r4+avVqekzGHizPFfCR
ZgGuwW0F3INc0o9TsNiAmfRuEWBWtR5vlzqeztgdcrQMm3x+6fQr1lJ0FD0UEZety+PIUiFRietE
5z5jpIHFEU8l2eS+G1VCYQ2pM/Y4ViG0CR9QEg7oZ2waqT2PD7XVF0I2fdLFeOiZJDAOQ2OqMHPy
dI/FwMVlgtbLKW2uvhswaF22W5Gl/E89VmcQHNOhCy/FEnQUWc33bfYwdc+QcJ6BCDx+LF0ZqVX+
y5xi7L/CJwnZhqzx1ksg3ChsjIywVmJLWDk3aqvbC/9XfLCx/BPXsazyUM+1fgjc3LfltgoPNYz8
IEBSiLMGIDtUe2GW+6kHZGfv7+RMxG6cZY2+GhLhKWUlhEs8qpQjdI1CRB6hACDylKe//0xvYc/C
aCsESgfUdTWjYUxPK89chIzo5SSe+f1WwbeGVRl6z1W0QIMMhVKXbx09WxKgBxR6oN+Vy40QYPjt
OkxY7zwq/33pfeRtQFvuLHjgAhPIEynFRtNm/tAbl2yfisAgFIw01k+ExrNIEXe3gR2Jgwtj64Pm
Ux1AypdFySIOisZl1a2vHHm1a5aYkioGk1SxJQwZ50cSbcfNi4qMWU/K/65kHfsEKxe3uj8bhcM8
3E/AcZ+rpmuwyDL+juQF0VXtz5V52R9NHXTtqb3aqGTjyT95Ejq8myyjFMzo5lB+DdCguWepHAhh
kEB0YYGy89GznephR5ZQ/o9gfbWmmXMe/iUmkto7GcOeOlbVhZJQhhACWjCNjnHOu+3VJW64Ftgc
aJlqZxlwoRffHNEUQ3Ua/AVz3WZ2gOlEV6jFLKwQ79GLzDYDdC1gZj42VpgpsNdEM17LCk9cRfKb
gR2S2KZymy0/J3ZOsbYSURNl+tBmcI0GFcbNbThtljEi9yaqGCmwv2KftmvzhPJ44RLypnTTVjwl
njExGwDnAuI0UmxrvC8799TTgUcAp/7R+QxxVXINozeCurhgP05yqJDsOG9GKzfgCaIHQm9yw54R
fnlepNq5PP6CdkGcbaeYYuAJzcNW8+y6Sp1SMwvR8w/e9isu4wt6CRDkVL7jt07BryPWl+M4rdRV
erOJouJN7nSI+WEvkSXNnBi0iQJTxJy3EzWTb/86HCQK5rpa8Z8ZkpS3jtl569yASPRrCbctPccD
hQqE43Xm+zIOlUrIPPS3W9v2k3ZATqoy8uWtb33XvIyq+NT1mi37oA4tMEOVboiHpqPoNTsLx0ay
QJCbhtVHt0p47E9AtvAhrjUijkiCWjqTK0Hq/sgzgH2UkPWJ4YXeEv/p7e6CWjMX9C5IqxOjg4+j
KYVmshztQ6ImkMPHxcEJP8aTUJ+5vklXxbsPm3y9+RoFksyW6MjM/xzLClbdq6ivrTfXijqKcBKf
IrOyvap2W0Lqcc9+qeZgJI4cpl/6dzHjqLG7Olnxw3iJ8bkzFui2NdcMP0Os/BMlmwdfpy/kpxYl
TyFOslBA6/Ta1fdzyRJgHj4NaJeEiy+VbFncRHdeFIgAf0NNwocQIUDAlaSnMsQfONOeDWG2j7Kc
pJvyyHxEUVMoevTLu+XUEghqCp7SPaQ9mTBnTxrmMn6kuyz2c/gV5lxzhlyHirtR1D0JOEXs7W84
WtOuSgcfmZr4KH931yaWDbQ5iIDy0gI+1dByMO2a+ie3psrGUMsOWQniuD+BFMbcKVUujnpkdwwk
4Ni2mcluxcJ17f76cpkdxzrIhxFbiAh3pSZWm+8xJ08XfqyxZ6c/MW459Pmc4i2xq0YrvcFNQ2f3
/6o7p3OqlBcJca0FgcjbLAm1EzewwUJ2fefKKEXjYFc2N99XbMbZWTGAYHtkR6ooQNiZ6pPAiGWV
m9ZrqY1tyLOAyXGF8sBvMt2Ap+/YEkQT+2X9m3M0PsTu44FMj+hjfPdIGGW+A/Xfb/iIA2zmSZ0x
RUkyQpLPPofZvr3OLXAcedFn55jbLozboJp0ZenPIbV95guNrMLwSmGxRmZ/jVTs0iQ7BZ8gn4GM
qhXyS1AHfx+quyuu52nOETk/xeGM6i7bd7CfDKJmUpyiOFvSOTcjqD//+GNL+cSr8h/Z2jQ5hT59
g1cSG+ZjkyDpRih6VWHuIKhf+q8eMoqlAR0Oe51gLbRU/spD2jSaQN0HZ4Exe3kmVjwgNON2crui
pMzP1JfQ6vY+jkz4hNopLxCYwH7XCmtFEfXrCKb6CCYDsUOJDq2OTKHjHLmQOocS9RP9f53bizYX
/F7Dls5EJ6QMjkeqngXvL0qOFsq9OcKMA41SkPi9JKaxgiATqjiluwf532xfwjDSjTW18QuwMQqf
z+BqkDecCxxw1HeBkU1HuMNZtxD2OBfzLNaDcaI3j6wlDX035ogviMlUF2aG1ChQCFzYlzWQE2+R
bb+EJeWH9btLCF9WYv1XXNucxtH1Fta2tl/7P6/QjyiwbrSL4VFMq3eqg2hCBrsPHsLXazN0+0MB
61qVPnnUYYtWctCzXKssGvMahTVtNl6zG+PBw9IWRc0buxC/nt6OPyZWwqRXBmZ23tLIM92riqQO
JwV+Zpvhey5KHXXf1lI3S/TfTas223pOC28l0vQUzpc3pzjD3xj0HA7mxQ3SdmGOWcjY1a9FVk5o
pay3haB+gMnQ066ixcT9NgQuFVO+1v6Pady98H6C4Z8kF/gReI4Tq+M5hA1I8os2SDkurokriEZH
vDYpJPXICYPtcwXDt+WNe1Cok6Ou4OOrMJT1vPIfiDbmFviPUrtliND59vwgWHGGk7K+la7xUi6w
zoZubhRcIXe0SPinoMOC1hzNgYCwNW3/E6iW3N+uhvM5+ql+dZOkr/+6z76s5LeTsmpK0qkacShr
W/PkPms+0bd2zoseTJtsvskUbcUv4AWHtC1poLzSbv7JpAqJaS+MuXD6Ny4BxI63q5SmxDDMcmQS
cIy8yOX9QsTPLh4/BqYwn7uy9CHcGOFMSMR9RAdMmh+QM1mNbS5yWIwjjSmBma66+TWoEJuH2jMM
HNe8m9Ex/qBCNm26UjqnXkbbdPpKNLvEEmUkUsjoMCHcljrE7f/k5IkaedA62nh+JWPrdjtkAl0u
8fQp7lq8l/2ZDBmz+xzeatlxN+NBoCmtdsmHSLjtOxDXPvU+vWUJ5L/GXyR0/Nn0xBzuV+oCSbbK
iMqdYzPV5bvxgAkTbDdbLnugPhK3G8i6Vjev2IHgMFIa+a21yssTVNdVjlFPTx7AGnlBeZC9Mxq8
FIhD9xG1esd1m072oQwFt24ub3eZk2ASWMqjEGdSllJpJAbrnQlBRnulzmfoL8vQdVslK0q0BJYe
/ldSM0pswmFM30yRqnEkBr23yeT/EMJYZd5Ri/NQEg8b0OsmOn5vci8mwekrnfPvpR248ylpupm5
sCtT/yVjkeXzjHaJQfflr2Ap0yIBVs1ZBsEDFeSsqCIEIBhieQ3rPbSe+vHTaFwUb0p2joFohTSx
ejBL9Ssp4rzyLcepQtnhi/vg8ukBoqPS8RH1IyR1d7y2Q7vPRcftp11a9gam6gVBoc2D34ra08Pk
09niKKfsSvZxeVw3MBh+kIc0asXoUacrV9PsTpGhHC8gLZRpCuoEHUtiRDvG0bODLsHg5XI904oE
4YIA0qDhkmjtWlr69eK0sX465nyARsabA+j8sHrHo+O7PCDdn6bG4tS6HxchZlrc5yMezZVsD7Um
1upGdvkM8pK5dbvTNjR7eDDYeIkVWnUfW9g6aT3fQef2m5YSTcLe6RoWYTJ98OoVn+qUaStWTwcx
2GxBiOZB4FOPiYZFvVCNOwkQlUf+TdWQCSoQ42oB3rax0OexyYbVtvep9wGkZP5IxdORsXFOBQbc
NWyO8WIeHcysN8XEku9tLiRdUd9/FDWuZnJQwdAF2OCU8UdLYtomXSXEtathMHx2eMbalGB9kjej
kWU653qkEX3fEAf3seW9E2WE4JnMw2uGNsZEdX6JzJ7mmufgt16niwr/y7vpDndGyGY2vLBW839U
h/rGUFij4hXtFxxi5yCNNZ8iCwuTsG/UH+Rl3tFVUa8w0+glknFcZVptbxpTLEJU0dmzcmEG5gWO
IaOPlxSnUGksSC8Am/tXqDErxDPgPvAEZw7ND9nEFK0tdHXQVNsJtJ0QGB2VMxiZgC4bCm8EIQ4t
3/yiTi8Evk7xbQEV6XsK3ZYwlGl3dDU7Q8MseIlEVJCgtKRIy0Z9mDhZlm+IuMD2OiaDH1kI3d+Y
dnFKzAO1ojFRrPHG0zPYs7VYfmSobPQDMSrPpiN44Y0TGG/o+2zvmxEfV4yoILAGLKduQDh/1nzA
Q7lhfxtH+/ALx2rKST53MDKGh1CNidns56IBPFoidzscZhmhiONrMMbrXhzZVZ1wlaUbz9rF5L3y
0hjmW/m2D06uTppoK82kJuh2e8gp+6VMHGxlAc0sEavb+wBpVSryWaKZFhz2ovSurO63zct03s4p
5tDZtXpOogYn15GLCPdA9TKFDXvnbRGYfJA3bKZZgnD9O3Jw3mplucyiIG+RqGkAkpak2V8YJYd5
VR5UpAkWGvaacGA7a3XQ2MRsS81LS4XPsXDNWkciuYmYoaeOzuNz/Vcmm7EyuOU8UVfXGuRI7tAa
c/K3LLCj7cA6Y7UgNgRdd+yFKiXstwLEwhuj2CmgkyLkzfZ3gAAnA3cs+Vzy/7WQUe5QhThA79B5
4EwX9Q/igDE8Dgg/fDCOFJwl8kxO1uiEz++C6nx9db84bz7mBUUAwq1s4BD6Mnlwj6tvjIBOZH/r
IAobfcUHuwLFd4q02Q9b5i07/93+9DpUAV7iGpf9dg0QPw0LtkOEVkRA/mB3eKVlOSSg5WNHXEt8
HeTWl7AuDyzZ11+FvP7FwIrqYFeE+IHtJJK7lP2p+C7B5ngX/21cUprajhzT7NOJxr41eXe6jcaL
hDwXNUnCQUsHI3a43BF7MRX7wey/mCySADeN4rSRNSq1wdLJRKI8T6fIePIiFw6W3jAOr0e43oBE
4JJUi+CYhN7TMkV6/BTVdZKDZf7IrWYrgAw54UklcD03bRjR/LD43+Sc1riJKemC6B7hh0QdZTjS
shyF7JNAR+mLST1TVf3eB/vDcqoZ4nuruaL9uV1qYPIN74rwQIKEe67rvg17/6lrpicRj07pkagV
CegicQ6sr98yk6SJ9v/vqwZn2Cy9Q10Q76OSg9ZQ152mn1c1yXGNrE/I7elClH2fnh4oBU6OJ1Ts
fVsKjYk8AggL+0TIqDy81m8tfIUxma8UjqOScafSqjsrIrbzBVKJ3Vu62+cnpwK+chp9CDyl73gt
8o4xmJ9tW/JyCu1qSTzizejAUygkMz8Jm/8XiTosudcYcyTb68H/hclgQsjU0+wkQlz7QKKwlnDb
+w6Wsr6tvcO6rtRmLNqjjxPhjB13hECQlUySToCWiSC0FbXGJYoClK7w4xGVw3ijU30pQGB7rtet
5AYSHHyodbzj5l6FGcBto1D+MCzyX0Cr3yl6v+pOq1eamgEf+wxgZNzoTG0tGPGLKIEQwAwhkBl3
tROCX3loqJLxGni4LycqwtN3MFvGLQC3nJbRUizLEVXrIiHT3a2XXekYjNfXmJTFA2YDKB4M0hz0
619sasKoGXC/Z4PDcPY0M9iA28kuDXGfzv2ANipoSgpadZeIqoF4nf9LZ8j+lO9lE1iZ/akUfiVv
eOzQmr/Qo/NorbBQwcEv8bSQfGlUP167b340zUYs0ib0iyJ3sHZa75ofukdTxIy4bZjUDRNl2wnV
9qHujNmM9sF2icbJo3vKTyv0hZ3Z9lM/ySVyJ/+nFdkUJKQBNIalmVDiC6Z3fe6ZutVcaLS/YSIU
JCrCZ21I1LSzbYzxa/3OLKES+1LTlTr+T4YQrozaxmNp75emyWS9lRc0zgtlMBSDyTDToiAUvB/f
N4NfRn9aJQQnZRmpvb/hQZkzTbD7KNcVq9np7a2zLb4q3EtpzpwbGCOqppRRrtfibrFcMydN8VTt
K1bLMOADGi6ANFlklgKU5icOgej/uwuj8ViUHW0MA4NaL9ZIYDxzSH7bNDr2BBGWcTaMp1cudguW
Ff+kKFQ8+OviiQ/I+/7hjmZnoVJvbv+YLBQIvdNqS8qylMEl/K0wxfiVS/RTd7rqbGMuRvT9ajmy
3YcpIBzf4zTbSxtWPUgyFi+PGpXT8KPWn/YAegvcyKgTYrg6vykcqzQytdAIhLvk37DnHVPf3sXG
wtULHZ33qHqaugl4kNwZ31D80HUg4S2rpuGpio3Ig5DGlftxiAPqZE2GDWWqJxxqFFNV47Yz/Io/
mDYURUsLwylqazXn1uJ2mG6hsS358za4QoEbPtbfbzielYYT5joEa/C2rFQOAUxxqETqLNMggwVg
T1ZGXGFseScZcNQghaMlFRiLO7JWt16r2TNM6/b70WFUOE0XvTH/cOFoYU/ujHzkRoSX1w2T/9M7
/y01/xkBdRHnbu3zVVgIPkSjXX0AIi14KDlwkLDyn0iziPDuJRmdGEcQbWwwPJWAKsR29rrrU7Gn
YLYPrcycPT9wzvOt0G7bdUHLY7CdiLAmH2kVLvu/UmuYsIVVFLJU1nvM0XlTot1wIZixJw9r1VnA
RprOPc73Prv7bC1MBGvCd8xXlyeQHQ+zEGr7akIPEUdkiW7g0MLJ5kvKLQemRq5EQac+4lX0pBjH
QoSEFzTCai+So7Hkg4TswBMq6fTCiSjOXzv8rT1QHVYl5C9aqA4iU5aPxfCZbyJcbUyU9A04stqL
aZT/BoJEHcuysnligcJLvlnkSy6UQO5ZvaW1lXqQAAe+R2aYOD7w/YyVtPPzNgqb+MBuBz2u+k52
GbtFbxy7B5eS3JmjlBsKzU+IoztDCtmYuwn2yDrOi2I7PHZjtNutydvt/rochHLtShAqOxv9RbAb
ctB9N3LCKtXQTDlN90MBcSUeQCAyp2CNrP7lgDJfjvxVvUzCcXzKPQf6i2eR4sbn2jkAtxcr+/KM
RO6Ti5prjHqOgldOYnSS0xJvq9RynjPsho7jTXGg+bY4av9KouZIi47oHv8bqENJROp/nJbCgH3h
M9MG0wY/x2DJU1/zWRqP45miR3NY0ZjyhxW8bR0TpEz2ytnySrMHxp7yLVRZLrQg9NzS/t3zS0eQ
/ZXFlczmKy+F9UyKBwL7mKn7ucSwvDlB/+3CEmgKOIxjsV0E16lUMlLHkw6cCw3Q1++KaD+bWEu3
V7mFgX1O9ebuUNx/FPJXU1sVpfzamJOuMOrNro9QVDWp1CIF/n+iXX2it5ZPFmXDHOhgmRetariM
4JsVm8CgYBQVLvVfaHM0Yp7UWkGkaepBLyl7tRiuph/PzATggVxihwul73pm1Fg327LGw+btxK7o
yfXmrbWQznDVuVMTSB57HYfqk78iKqjFl1i+Uq9mFOez586A5ycjjdIl98ENfWj+DG/Pse2JJpSc
5fXnrdHDEqEiOfzJzBiAq0Eed3/h5kSUiDjlHFnmI4zPNsihsfldfdzQGlC4wAFiLypDpPUSQjGH
2NqZljUO1/eTxLTXW6dpjnQ1SiQBRYaq2HD2P8D55LC5EIXvB+SFvsKZSry+FQ06WcJYjNL5Boqy
TMKZH+35c3AEbqKUH/6wMvrtCyCRQB6vIcaXbJrd2CXZVrZOnjkj6e3dz0hk07j2tcMF1xR2a4x/
Rcs2gJ9HkiX3B70lSDx23vxz/OzGV1ZuZoP4Fc6TTrvqeO0u1rRPYhNQv/Jq8/mWxLvBvsT1OnR2
5Me4nMznsbojoyOtKfsglEvUvU4ltyxb8u5rqw/5VAPCQbNoXgUHtZWN71Pkx0RlrgoN8Muxi4Cz
zgWEbVH/tYdx8uRRoEQ+/1VzEshEO5nGWFwL4YNEgG09E7lZE1Sa1iOmQg4uKIxE7BXkQJVkSc5G
vbbsAjIs6KSpIPy0m4TjqlF+1g11/xPiZQuGxoQxinWcUEQ/jlvOXLvc5v6Qdn+qvXj7gMhE0ogy
LMo4DY+YScbrCzModWRyo8Jo3oshND9RODAbm4EryfsYZPby6IC7AgGcrdbctfqrGblZ8ecqlwjN
UAU60HQwnA7aVIzlbl8yxagTlBXSloK3D47inySKZQAQT0khWE51zmPzncfxDVIUfTuKNQdNAC8n
5dmQpu4M/CMyf9QJ2ylVIrExkQqboU4Kp/xY2zTvgKi1bSjZsqnyTCowI1fJTExgOx0MGsenc16m
tEwqyvaDtEO1T0+xztw1/y5zrMbcR59WCAhgKMmkAJSVll7QPxR7G/pUnb6AleKLu4ki2UeCK5DF
PucVM09LkCFvPhvem87BZoY7/q2YpkOmZUgPnJoff07og7lz2KqABNlEzwvBJxxQPlTDZiGmgiFQ
CFHTVwUF40rn6FzK9tskwTiyIaAzjOTT77XRev1z0SggiFqq07WSpuaF3DgCayARoT0FfpnHzMmK
1cFQCsFTFXhRia/o1c198hntOIr7lvu+lG6Ru35VwGXr+gp/bC+jCBBMl+gMgpNKul+8Mxl2oXxm
9Jxjbw8XCqdUzB5B+EE3c3PgzclzfjH5DYYv5wWXlf2UvAu9TfcLOeVnom2iHlsZoEhMghxCfkIw
YSHj+dLKnuulk3+4oUvpGCqjZpJsOV83LUzX2Q1RsWpdj5FT942BGQv61LXykkw2rG+QBSBNxNHS
SgZt3Wo8suKhFtqb/dShrp8vW38OaUHwGeDE4ejCGC9/V7/ZXEwkDx5qNaoIAly1voo9ba7w3rWF
RiVpCncK43IA90BBNt1+36ZIMb4NsgQc20gX/MRwUxW4Vb1eLkHDVAe3sPW0L41adv47vjfJbW5P
In4ByVk1XxQ3cvAO8+KrrvH8WmMKOQ5oiwZJe//wfWtEOPdhtaDtQCHx1KWrEc4N//Wrlkif+i/B
ACxCSGSw1Fxzkb9UG0Gjdy7IvAAvVAVDC2eJx/IXeYr6mtTDYntfRgaxANfqb9mSVm2pFxU8Sg9t
0v2M3DQxRfboz4bSP+SzsX0olIi27usjgMO92ym8rxVKu2bAKI88C5yC8xCbw6QMm9EUoh65dheY
qE5xkw/lhQdyYQDewrBYpk4FNZvOgKpsgxFW7dDDDp2yc/28N0RDqlnaMkc9zk272LsGxPTXYfB+
0p+bjAvoh8pRLOwjacGgPWHYAAFurrNoXPQw8LeorfxuaZa5+IQlMVD1wzweq18PVMRg2ewHh8wD
1AMVDOV8ETggUasj1InyS4Jxaw8ufKTc393SQM+U20Ar72PGYOcdhh+9xf+1txR+frPJuriRMPYB
a9L6ggZ2LEEayIZCDoRTmjvPodaGM2LFtT8zcz+mFRGbYIlZxwAACMOwp10FZZG9ilqi9phgXADM
WQYplPjeaQJnckjdcPbITkvEb/MqIh9okpmr/D5/7qNQ8AzUx5gHs/NrG7Y9hIiP6ZAhUW57KVCX
1D218h9y5AOxbLhb4UNxXtjnZyda6tKSCz3rF4xIuY05u9DSO6EdFO1Q9i5wS+xMC1sBmwM0pC+y
cbUS3CR1b+Nni3XW9nrAOIElQ0DLvzmZ+iak8iht8Fmmnsgdj1azvln3vP8Y/eqaP7D0aXxogDLk
eeaGBpTMjRoYgVa53+BvyuB/CN7m1VcqdD0GYRLIG4B5c1blB8165Bi/TVnfopf1C1faML0caWOI
4J0lhWI2viTA1ULGbFF34DvVaBO4nnJRYCgizxGhb1HHumrpjh0ZUfnHbKjegd1O+nE0ZJmRlWns
N40qGfR6mFL7q3lrvEiaG/3eUtU7N0vxaBpOqJ1FEr/ZiQ+7vF/0jLklesC84/u6c6FLgn/QbBJE
tLFoCuLv/WVQXKSMh36jldN12KJbHDnv/fI2HkVyNt/A7KfqUBXYBQwtIk5v905HP6qpaNWHgHj8
ThicWPa9DBNTagPLyrULzbqdUqn+kQzt6N7VAq0Ly+6Md3/62x0Z5Grwe6xT7QzclFx7LlVzdHOD
q7yn7TMbCUCga7leWhrnZMWGzkRfzx7gKyu2CSpIdeXJ3ugu8H0astO3PSxpykeuWD4tVvlcRYid
Y7+ZEDoKMdEQLhHOLJaWIf+VPYO2WzxrFJWP9cTZcCgW7bQ83070XcQ5XY6lr/k9RkNpB4EstYcu
nOcSd9SnGtn+K1xE8jGv+CvEWws41suu/fnU8gaoBWZVJDVeYXucqPUyOa/sIudBvb1sjYHxu7hh
qzoAPcTe1SHhXFJepYUzr3kqnG0Y9N/67I37xv7JfnaaZtmPtvm3wWK6K9psvMjNTcMWTagEh+2/
lOBzNw89mgrShTpaUDRzJ9CW+VyZcW1VgdiejBXNh3Un9lepCjwU9LnBQwde5hvZX7hgCwwNslwJ
6jw+btSS9FWX6MHVL5zj8NsQzO8q57z2h8UAnca/rWjgk/sGVksFT1wkpX1O470nXvLLcgQV2ZUr
t9ODyyoE+GQ/DfqB0OrMxq6nyJ/ij0w+FKgVCd/UHFYe9Dbr5vsaqz7QCspjxDrH5WN3Csh/kxDq
dT5YPevIUSvJgHQ0KKVoGKGclxg3zOBCS9dJZC4KOK0Jba2LwWyoYt0dwDpIp4LG66MNjVXwPBuR
B5foZYDKNWmWG+JPTUqaTZZq8JBcAgb0/yUBGIOckURSYoqq6o2jHMqfeQAPBWd234QmiptKdobT
UcWxY/PvF5WyIDwVrrzcIdJsArv9XzQ9i538YYc7OuwjkujzCGFbTitCrxJm3bBfGALu9ZTETJux
BacHEYCkD5GX7lV1IiLO01udCL9IJIAtUZsmh8+ZsNRQYahb7ZFYef6ywbD8PCl3Ffo18G2hStkm
hBbjuqfXkrU3Sp18M5h04pbeglt92G2GQjbVMbm6nDqVVteSneff/2Z21tFfS6IdyqUoYKBmIbIT
EvfgcZw5ctaPSyVOtbh9Qws0ddRfBPctrbcqW3unURsatGnbJ3sOKj8egt5dxDKk1MB7VKdeOSeg
jH4df8dfiTOWul5OEInH/uKX8hCEybMc77BOBt7tVbf8hd2jmLSyQut3PsrPGTDpowIA0NoC099s
wFFN39Z3K14scLcH/B2z6W7TFs4s2WTS73o91HR4YXYdH+3QBudeqhJYkB1Hfc9SV/eWqvcBo5Z2
L3pn/dI/sK1l+kKqA7prbvCO0tI6fxmdb2zBrLXZ6A01INIrcO6EVdXvi3Nm0ujPwnMBkyA9XhY+
4ApGEws31fNVMDghE1pndyE+l0uBKDMMxC8QQulkU3K7wy/pBaWhGkDwxbbZA0+Y+G6PIgfRz6jV
he/TsMiWbZAUbv+c+MEaOe+mLnpmjup7QyVaOdlfZ0cGFlHmQ53K9O5CZyq8Pl3+52vVGShPsl5m
g3p/f1H/05h01VUtLCaVXrI1ozzRRDEDjRhho+znwHx1ndw3TD9CnzExEz4otpcIEk75O4fsWuFU
bclDI5rQoPZWIzOL+3n8NSb+o1Z9dIAKC+ZlO8JTAQFzLTqBMJlx7Gprk7mKp5MTO2t1d/rg1cHW
/MO+29Ro8wK6COIdOcMlfNZN1n89PcGPKYuDr2+91RXI6d+zgwyJDf83qJKixu56m/h1Fqf/4S4p
auDlKnqihH4BliIRGwAf6WJ6ZiRtUy/YUw3Rf4HydGZu9n+bbX2shU4KxAQ0IrYFHKScUkViB2H9
TcyjpREY5zRvUCEO7eU1QJt0eowC8tNbOAYqWU/dp3sHbTuYB8YwLfkSs3GpnSVVp1kV48lYLrms
YA1BOb8ApE0lXhhz4OZRIn63LPouNwAzvZlAdjdsO5m0MtJtoIjy60bS6XvIwzIX+4ZHqZhDh17m
Sg8Egu/thUj0UokCfxeNHsus+5+XjgLNGAZW9Im0FyWHBnUIxq2L0W3BcGTDs42hT3yxcU85xEEN
L7KRj3rGAWNh/Sg5UAlOtznU1xum+EbiC+SF/WQNl4dyQ2R6/5Hj2xQJjpHiSevlc9fw7Kud+DSg
YYeLKba/IIFCa0SsykMK4F6bDlRUQ+uD1/JMYU+CL9rdNCu1Z5/ovRLustJl2Sy4n23MU/4Np5FM
yXPTOejusuH1rZZwfRCK7IXQgP1pYvvbryjT+4yOb1+paYEHrBFUJRmG786DNn0plnXhct9BgFaV
fRuZsfTd3L4ujzfU+bczPwPIYAi+Yvhoj9nocGaBiJ53Ty4t3197dcKbLBtB7irscrgK19UMJ8Yh
m9eDAcwrNEfKj9L9IeUnofPRJURYOnqpH3IsBT+mPSOXBO2vjrf4Pvu5wuc7h3yIcGJ7sCGkL6uC
XMAckBys3FC/mCRr+VcI3jfFgZobBOaE7kCY5gb7AU6/9a0KCRUvCfmSJxQQcYW3mK7539bwiNXM
uvOpBugK+VEH3FbVi5xC7w104wRFiLU0AAr/JM8QEhhvnOJ0BOrxW4cHpHtipXSfgwrWH7zu5jsM
N8I2K99zjfrwUIZaaBQNlfPnQ0nTASmRgC9LI3SaQMxDushVP30Z/7td1i2YjRifbhelEfohrjzD
Aqruuc1xoYKMwfPRXBGJ5kaSLCDojjSBojsxOR0vyuQQcXBowqYz610LluucIIiKCKHi7sJfzA9r
DcyZB0W5yR2X2S5B1ytH63+REr+uJJGwOn2hZyayGA5mZSfO3I9dVivSmUFW1AG1ObtzBaolSHvm
Pl1Q/ml7D9DrHhfCsHxO5OYKNqXQ5vdl59swszyvPvUw2sNUHWC80IfhmoZRTTekdvq4nYcsSZLE
FeWYnLhl23CZAfjn+W89ATiVEdMzalRdfEtiI9R4iPfhLRhIrou8kb2wgnmNTkDjFTZvwYY24uYj
HZBwWyUKWYPKMC9YNpiWxmesxJR/SSekWak+VgXjYoDKd7eiPAyN0EYXRSPFbMsETSEmTG2IuaDd
kalYjdNFPDw3Hl9y/kRozS8xEMp+6mkcyWFd9QtqtTGOfzO2eyJi/lFsaf3uHTpo1QKOB5XZQiZT
YT+l/1uevm2Pftf7lty5vR/zAhcQgkOVBv7nf8bYQcT6WjmZQgZzhGtkkkPPsfkdOf7mGNqVdyv7
5rBcVxODOee0HIHOdZgiH6xDU7hqZHPZyq1WzJks1GS8EfRKFX8rsGLb8byidB3trMC6qRBwgRGc
mfSulGPOH51a8HkkE6f/JpsagG4ZkvlkEnayLPFiJOlFJUr8OCnbUPDnKCx2lqCzk1AkakgPASvt
b7Arz9jX7ZRq4QnWRNt/RuaH36qeIflaNHybhQOUOznCwBt8idLcoPq8pjCzvWARRUFTYYvDfF9N
eNrjbllV1rCfiLqZvvx3vlcWKc4ITi0A6DKx5dnasQd1d4Ritvct7bUIYXp2/5cOCHwREYTltWhw
KKN/3QwCyCgXBwm/h6TDDTgIlvz2uFLcz1DViTBk3KbmNQmTYEl6+1K65ZLULBzsnTBDzc4B7OQ5
GepiRPmoZqF+bwLxUztQWotAH6UQlA+ouOr5qu+X0HdE1MTYzAk+VwjNtbYbg8W3OlCqJCsyjC/f
+igv1Tw5eEbM93mV43nRg7GWt8GhSKUTvW6W5otBbQzI1vfP8pHbsY3egntRwncv7OhlTPD5Ghoo
zghnJWEC4f4tA0TBiYZu2lRGle5MUovEE9G7R7XN+ZCa5EmhwSY0n+w7yOZZXVKl16wJm8MKxq7Q
g5wANYe+OChQ+EyMPCKTvSsE6YtAExJetmYlS1JATgSczrdQgOnFwee4gS0JiK/Tz7wAresPgKQw
t5CkjoE9sZ0qozrEpgkiwpbDXwiONLjCd8/tYiqdymDyJH5leqKo9fMItvDrh1WC3UgSD0Hjgkyj
zGSdYaxioI3o8cgMxnFO3LjWuNm1aZrKYVCdhWkYimvNwdfGayfFW3c2V8B8NYbhl3so5XH+i+bR
D8p+BXdFNvbdnSTaolXX0zwUrgteS9g8TVSThTenYOMJ5iD7L7y1hOiwsVa/H/AOtNfaMcOd/DQQ
/svTfITRS8bmknHbDRGlQp31ePmyClRgsxZQqw22F+3+ee9h8AU7pDlEdsZ+OUIf2s7UZc8CvmHd
UPkWq8/nPUR2UseswbnD76mG0o9Kagq7HbvSiv0HC7EsJZi8b2HuzmvuWXKEWJQyc7fkm1WUU9bJ
zzWPy+INiwVnvLm9S9ForcuW6c0shaUmaJBNtAge+R8Tq/qsa9qFHS9TKeyj/IiueIIM6pMY3rA4
7Qryd5zIi0wZzJACMtw29elyow59vwTlLRodU8JYUBQFOT9IvumDSdoK33iV3lJrZfasToy4vKCf
SwEJqf/qPPTVmDiFrrRkge8RC7LDCr0yvZXLWsPEgZJZ+oYs7OFh87Pxu1fb4I/rNgj8MDvuhxaG
OdOh/bag9iRrAYC35n7uvRf1TkI0X8B0Iit8SdIvcKIxs0KZWq5H/03H/8KJx67jakK2g+y5QgCM
LiS7UQ/4M+V60s6/XlZjvxZLb9sRINSKwFSAydr0Yus+OjkI08bwc7xksplvcocYLeGH3OrYUsIS
1YPRo5EM+LrPm9gwF9Tx5XXVqxWmzwQ98AWxtiQdw4Zu0SbqS6LDkbUlOpqS7wEj6wiXbA/SY65L
my8AGBjND6nTI8Zm5Ogf0wBk56ljvGB3HMG8rlP172uCc2dZXMDQ3NLI+GEyx68gTjrrKK+o/ONu
T3zls4DSs0T2yEv6F7GSCvi+tAL3j/Dj/dQ5MpYZVzWHjgCFyyHtdTzsatitQhJDArV7YOAHXjTE
GSLK8VE6fQ7JpTvfiIqFRnMTH/HRmd1w7ch5I2vkdlpzxLk5OOYbRxG6k222sGoVlt5i2dBgRJZE
B0izGG3Kg6fNggYxOSrwc7wJ8XUiA6hcTnHSCLMZzIRVdEGMlkWm5690d6BNJSSPsYIgFhyYBfKf
X9XEasQsotyls/hoPKMnbXHBe/KTMrFpGKlrXXgyHovKIuteAr/exTGuRJq/qhJwy3M3QnQXBvGk
Af15Ilr6uwjRQ7WVkRqiQUOZrHIZEWX+CKhtdHp+tBzcEGBMY+vTD052FPpY/3RFEGu4TZZsHRhA
wKvtND2EcaKG0CazXg+1YEWj3Dk14QizAKojWwBSbDfMi3HDZfFkxLm0k1E+NAGPsyNrec6bO7z0
ltJRYOnTPkTb4v1JyGeKQyRgWdQVgZQwOVokTMT3gdKCAy0Kb6a5wvdPu22i0JLU9O9f5pYfk98D
/NCM0D2BkWP7aQhmxG8N86iCFbMGAgypM+W49AcQoJP4A8CoOjVdMbp3OmdUrdhzIIiQ/HjID/gU
SdO9VosUZBAaibJ0fX9GTiypkh0mqTZCw/cerzkKWoXmCjWJ5ziYrJsMM2VEXjJEOIWf4FynBFZY
YkOIRcezrEEFLWbbLk3JXKQsOhi3ZWAmofNfyPPPyPTmsi1x+cZ4CuSozFIYIZKEXl2YNtSKmmDP
Aohhh1kt82VSDiovCX5obnhyWTXzP6uvluiTmMdmADz4ydg3MtHixc5IAIMP5/4oo6g3SdJf7TVU
e2SGhatT0oDTT4ANq27K5w1mizNinMJYlNIGGcTFUtQYEKcUD7ltR23wjKcDDKU6+wowM+TNvb9i
jOi68n4557jCE9Uq6cORtJXbcmdiABSJjc37f+u2Y2GsRikHXn5eDbuZJDH8dLkoB+Nkm4e0c/mh
8k1MnZcdQnCc9hISOccHrP2FPPa+QPdfFIiFYsNRchmu/kfRm+KlpzQRRv2L5b7cODTPu0e/5O/l
KCWr2ltlIJkcc6h3G1Ge0K7ErXHnCNBOiaW7DN+7+hdczyc3n4dzaXbHZbtpR8Xogc77izzCmlzC
p6O5MzsepND7ZsSI6H11uOR5zaMfGHGSs7dBxL+6unLG5NLRO20VUqJfCrpEKAc3ofT6LkeIQ+2f
/32LRC+PnXmGVOckZ+BH+QfMbeQM1CW+4PfirqVHqT1NyAC+YSDJqVd6A+/x8rruAR2RvkMrYlE6
GQgLvav+i2g1Ld7FNm5t+Ed54lVg6lGEhjmPPrT+kQNJRJn6THLf7pc3zU45063YYrD4ZrAyvr5j
KlsamRcRpmZ7yXhs9i/yHYt9m5eaWuV9BBGY9hMObgrOFUVnX0bdUdUj/I+1Ilz9OJx9ORpg1G44
NFU3bpr7S1h1kyh6r5McNbOXYMcWEsUV3sS0gNM2gUbtej5mXvp7XbByOkTA0ilJG1fuVfxWT2PX
kDa4gqLb4b851LSEM0SXx697XxaK6+RVcilqZ7215voOANl/VMyDjJvsqfuEBEg9WVk+7La7t4J+
AaUjg9JVS7AwQcZ4yJG0q/ZzgNcKik+yxD4izMdVe2AJJ+DIQYd17gczj72GATIW2nrfQfSCkXl4
WT0b9Bvb52RQxJDr7mUA7eAkFuAmX74nBCUrgA/PveKK5cvtpRd+W+JGLUgOFwGY+B4amxddS2Fy
VuehUEohUIMw6MNdjy1pU9KHKzY2Qq/7BjbHTI4xoVF0rS1Rzw/u7Ism8HVK72kuSfdBVe9ZCwcx
9skp6VAEprIB6RgEgluqfMKb058fqwzAD33NHy3jhiVnYYFNt8H1fH7IU8rMJi5ho8Pvqf3sDCXH
haGu88mo4SvdhgA/FuX1gx4Uns/QIVLsoizigx1P4TbdsoJ0I2NCEl5BhZ1bABa3CctJHzKRF8HF
LMU/rHoxOWo+ArVCX+VIwykKZNkW8hpworP0CUuVJO16fpBNPmt+73CPkCTJHLH66hNj9iZDMdbT
bJYdjy+K2vkeWMMf7AjCkrEgBq3wAnFaJIYhSNI1bdLiRbUigw/0Ujoz/ZzESydnj+1DnipQly61
IBDqOTKLf5Rpl/n2wlKjTytKf6u9X5bJNJ3Xr2HHLLis5Hf0UQCeP6nBalnDOE0irbz3beM4NEkV
RFDblPA0ml381xBYp+aLbqSYVrbU/CG068pLVI7xEQWNTOwXnq6SPrArKjPQjPeE6zzxYFxd2M0j
ox46ZN7CTcsUcs5Z2X9mezbrfyeKVQlaoO8NV5n3DcgvwaRRxL1+7c8/0ubWUvvOyR14w6Kr7KX1
Og/DlbzQBzBLWaEaeFAj/IVDrFD3QfKkxOoyvfljRb8u/ZSsZ1eMuu6KLurIy6t4qWN38Kx0RoVd
jBgx06k9IsdFa/HdLbOJ3EJOiw288E5aWZPz4VH/uRVapCjUiVxkh/pSfGKccpDLAV1W9Md3NOzJ
0hSNvJkr6yxuWlLIXEQh6Jy+vNEYHOfsOh7SlFLhEEgStY7C08Aheh+gxrj0jjAVp2DTPNIliNTZ
Rp/kV1PDLWwuo3v7UUi6rYjb2ZN15K32GJ3UBM6yg3ya59kYJTr/lw7zEuEmB8PkPboc6WoXnQCW
f0gjjEmDluakzK0gl0D2C/VSvLYi4UBF7Bo7Ub63Vu7SLBg1anS5kSB0eWNRCUMlBaMnVHj56Kju
/LUOWItDaDfR/oFQPXCPR72UqBdgwPRQxPkJK+AwiyohKbtOrAbiyYiE+9fZ0l+eKG8puUb7kVnv
UVAWUmzzzGF86esfrHvGOiU1nz9Z7LUP69nVk/dTuxmb6lDLdEq2CM9aW5aQl4SgVpBUFNF0/Bs5
DOGBtuK/FyRGzK/uqe0P0pLqzEBrZQGFz9i4QDWXGz6uzKmGisa6C/DG4pLIb4d0fPu2nMKnF9q7
nxeK3tOlnAKN3UDdasy3X2GjHfSg8o3f3OucPU/suEqhUgtFOqf8Icb7z1ELoCnVXAFpWQxyexAc
r7TDXvwRVEdcLIi58BiTeu7b+2+BKYgyXNLXb6OfBD8GqxZQVXCC1XssFVI2nnl0JS+atbSEBTQP
xp3ApGuYCLCFeesHHw1dILcUvOvnq+yJHBhxgQeWBUXCav0t6R6D1DMo1dKY71uo+0/xn+aHjnvF
0fOAYcArDFy6SLab/FYPAK16cez/pt3mYZcesElMU1A3Hu06D+zk3nBvtyz/X1R9nFt21MTpVclt
0Vqjz4F0kobPSSghnNe9ircAE1oSfaxwgkZIacg5F9LVS9KHMCqO4zKUcwpzeJF3tZPFaaXhM0B2
G2Rje+kwlbjYeyjsXqzp0eBft4opnbzSq3jj4p7bUUn8+aPoYk/3aUpIgQ7EsVMZjrrGyQbMGU+b
JgYnUGEwRomWwpxaaLF3pNq1ALT0mBZIFNMEhW94LXOoWWXzQxixq8qkC/J0+e/R8iYE2OOI/eRZ
IMvDDAXCY97+mL/R/xb4dJLtmrdxRTFymvGxFMBsa9iMrtQ0rD0M2HGqvzCvXkYfFwlgdAlNAlQN
qY0aUv4uGHsbnlkq8GBX1sMNcE/UEjzDEpQLnuM391XMPmb5TbDkVItFEhfSRtTZBd0SqPnGEpeb
PtQcpA61qHAPrRSch5qhyBCblDoctXcnuBt/ruqyQeWFcvev8ybwNdyrvwdNcb6APlRfhqcourF/
ndVqiXeRoDA6Fwka1sQxpb7j4ndPUcSxQQvFFpjDI46viS3RTogTBItTlfe2iVyEmhW3B+x3Mz8U
r67n4w6WTAN0o5hdWW+9nhFViJfafdXGj0m2h1CthfESKgx7FcmxAoq+CFWqbR1KInwSQBYXoS5Z
MVihc2l16T/flQTxKdC9D1fY0p3Vy1dGNL31l2BPxEQcmREcD+EMc+J8M46/JHKnFfOTi1btiuOA
ld0ymvXov6ySc6T/vbFVRKGzyq1VVQCxt3WF8koIs3+TwhgLwvb0onWpuSrN42JLE+JiFNTo0Rbk
Uzea54F7X4+Fp/fDPonuCRs5vvjbuDj4+c/tWaSXnEy9vGO43RV0WYFGCC131kDW3aFpqXeBWZka
DnetL5LN2H9FyHcEyQyTKhpTdwWniYpo4PtigYtZyxCZ6tTEM1tH1FCQxuyabBwjbSPP2xpnaA+E
rX/7G03DqSXE7y7WvLgkATNpOusK+PzVskSI5diUjBFltrXOiaf9ounBZXirA9NI4+4B5DaeR2g7
k7sztjvRPI0Z8IsrMTfMIt4dsKWgDgN1aQHV5hYyO3WUOhtEBo4zxnRO3uJGiDJ8f6NNL0K0Q4WV
FPmVEBHTbIplVCecym+2cy8F7SV/j6PExlM9H7x9wCBKJ9myVQGMZCbGEOp1uMhYJkIDJLVqH8NW
QVpJi218V7D+tGwC8vBTOFs58uTtQkhSLw+5C6vhMawh6AF8q8rpXt5gnO1aw/VmCkJA4Df9HlIL
voomiA7YEcXppS0iuQ5XZGIYzCcqGbXVRpLS779cajLAkGZKX82D+ejkxSabMjMSUQANgL5UWwn3
jRbsWK2cC6yy6aZqwP1mwy7nmOVBkmYdul7KpZCPf4caj0dJzdSpx9me3EvQYJuT2NtfH33wI94s
jDtrFg9v7jSIYeKwci9N/GmN07HVJne6bzaQuDxa3hMAqon++uLnZOZLOUMnXVh6n60enjvS36Lz
dvUIlw0YLvRsTLP+GiZTiU3iJXdzXAED7oxFzhJzvLPv46frLJvmmTlWthpfcj0gQYNw/S86IJMB
QKnr6HnOxbZOzxlO9Km6lun8Kv0p+jKHM202Ku/O7d2npe7A/4lmNEVXoUcvix0SGYlSWVWCIGIy
4zLzUr7Oe4TWDCY2CE+0l5mEOntETs7vvkM9Jr0kggcrS2W74Lr3rUIjg+XSiH+WJqcgwauBPAlD
wz6NwR2slNlo9KqSF0ubOxIXKZ060e66nR9qnTGMNnXhQyukTw7ve/x7KMBkY7HDb4hFW6PQfZd0
0RWJKadIwBSvTY6Egf2QrkGoCVcWaGnknv51GZyP+i8yqlx0hCn364MO0wWxNIR/gdRmJURsWsyg
lCrPjBPsiL0VK8U6BKtEE1RNn0AKR2w1hL6c67QMyf20L/fMmSo0SF7UcTqPNNvafSXRqZdG7OB9
HRQtT3baFCNgLuy8YOJbGPru21buMke3D+Qszt90Rv6nVyANVOgbMWXStx6FZEgO1BBwnsf2qp8L
8Zp2ee77flJ8ZGj3qLAwvGhS39DSuuusX3R9oI6ua7m7ihLc+IpogvRWzLi9uW1ZBOAlMeGsN3BS
zHFQgkHlwrmvnoQIZ+c5Hnr11G8ZlcU60/cEzWr+smRTF1KsbxPYFLdfGMU0L38AiE2u6D8xV0T9
WBtS0+wWT1PjHTL3d9+DqDbWQbp1f07fCTZAsQiZrf/uq+nUvgKdZITQG5MdqFgKOngTQlC5naHI
jI5HiF+hjzQhf8FK+IYJSfvZPCsWcEoLpk/lFA+HJDsuO5PniAlucZFuH5f5+kGpbmbO1xBBxcJc
NQPMqk71xuKygjGq52rqQv4Oeav6p3P6keyO/xdicn+cWNF6A48Gb2EIzAc4yTmaWxofH6176L7O
vMPN5sG+q2zjy3Sdx6RjtXUCeNmJeHVtz8fKWaolgaCiYz0tnCTKhmJHqi54Ewdw1p+oc/VGWMcr
vQzHueXW4JKm4r/fAJUBoIGW2h0HC9xB/PcY69k9TMaaLDZdYAK+2O+gMP9Sshgz4cG9alZoJTnK
5bIbNndf3fng5HlxDAKqdNsm6pyVf0hbHsTSzdOBkVL2YTPWdR8cJEY+8xKJdrkuM5zWxUiMLKUw
+GJBUtk8uwya9EuOnBDoMU0MRbfwusYbtDnrTb/4pWYU6deiLYw/dj9OQXFF5hGVL9EE78qn5i/C
tsX3GBonkQfrFvjCM7Lqfnrm9heXRo2eDwLn+ZnCUKewtneT/j1C1upMGDc1lqyADy6P06j0CATs
rFOUmhnw8IUdegRQE7d+02/5qomYdXgu5ceDQa7PKWAHk1wbCsn4wmtW9UWRlhAst5aHnPJPpT9r
PFWEfXGpGRI5pdHzQMV+CBphymcpNkli6tx3gzFdWPI0pV0mSL1xPyma9RFJKWlLFBasYOLzS31W
WyomquN6Ssl6J86fb4IbugGQerPE591KuimqpPzxwuS2TxlM1pW3Sdp0+uK0i3eCeoQjS2v5Kb7x
FggEmZGSFVYB77fVFFyAYsED1DiwTXipNvgoPvQ4CWhQ2xc9roxEcbLjGdzOt/djGLib48zBu/xN
jmPc6pfRX8BxFv5xuBOw7pMzX6SOlTW2Y0nj+/9kPONspRy6vUGfLfohbAkZDPmlGPwI+4MQcoJy
p5QmrolDPWt5zL35H0hgAQYZUp6ocyKtDEXVuOsifVQmZLql5vnxNV+sK6b0X20FBK4JQ3b2Tntt
mW+Ueh5tJCvuYb2lYSHybm58MA+AlQpT9uoog17KvwzHg+ERTwAAHeMcRBBYs2rcfDsCT4Q75b7w
GgQl/btUSnpzi0Wk94Aite/nAKOqcYQW2yAZlJziNuHubH7naT8SdFmk5II4Ds0mav2vHHd9PlWy
Z/pBzdmRnZgg6FLR25KHecRy6dvplH95jEKwfjPY9j6j6MkVfpGay7oI2GAUNkXfOUG5FQ5iUa9T
mUhYDG89Pf93ezy1m0sk+ChZ7HJbQbDL0wwasRIcDbI8PNAI8NcXgzLbp/7UY+94+lAmZRJ7dzRo
QzTBs/fGgaFqX+mZfyqcpO92xB1AeowwJ1ToSBh9ECXvmIiNWfG2JFItx8KBSU/pYadJH4ECCsxh
fmRqTNzWvA8SVnYo4cfOVeIyfwVK/5cf4OTHL5rGKF98yFdKl3PIFE/CjyMnBnVjHrCanH71LhNS
5aVnkqd6s8i5Re031Juyhiujhrj59UhUwb//ltw1G0NZ9743iuPilToGZh6CAnhu46+kkxo36k/W
eV7MmQoBN537cG70k8U/l+W0Mx6lUJzdcnZj3xaRYLh4QC9czUhmBSsKhc2IA6oXX24UJTC4AGJN
af5AwfcyVh6h/stRyb1lC3RNl1UBmHUggNLy6tn+vPHQdQh7rQLYwRzI6qB5e7fNWrmUuM5cS16D
SmqhoxbdzkMN9ppH8EmtZUXknp39a6JTR/JU2JdWkoo4kesM2rENC5JzaNWggUWtOmrx5FgEhfLR
OUKYmvj6CCJzNYghtPqkT4uyZlpQFbG1lEirISanLMcRGfOZ8vYjZ4pAJ2kYMugxOnGyd8yXABfE
yKSLr+/i0AOt6OUGlI0VVPJxtU/AUGSom5LXI8Uh7zZdt3dvS9xBtPKq4dK+VnZWTbPs/QfQ5Z4b
W2j8OyZR1BbZMPTWpw+hzvY/nnMp047MchjKjAZnPcXz4QFbvInm383JZc2x+Ix418AhbHATc1h5
QDGb3NIW4Mxu69rHiGRBPImZsglmdvOV5TexSWxO8uVPtnC1nwBaaj7WLd+muAqgdu/fyIOySnmc
Ts3SFaazFejT+T4dItd/8ETVdiq/PBInRkBC9wh1QyLWsSeTfwmj85it1mHcqAyvRbF1hCywCgcc
dP5brARRnC9Ix064bFAdckExOxFeiaRRQ3pygRMrAcA+m6oXol/5PH7VKqXI3oLc/W1l4Sjdw3+3
xkssx9WAsDM+vtspMCDbWcDfrvJgi1hqDSVRpF06uBaW+/fpdrI2SaP78V0WhWOKEdMr8MWMkAW7
vHoa+nkuhGd+TRWmK4t8rKYdhprr2kALtDnRoODVday/2jK28nKML7jT1J5OTJxS27zYTTH9MZNi
cdCFPyAP20uSuZlYP2zzYQhZT8NgFqJ7rHbhD1k3fntZ/qyzBqmvwZimA/K/I4CcxQs+CnmhhKCR
xEriy8E9k+37XiyXRmlZjH1sOxfE5nbEIQX+DYn1xD/wEXboZlTRVE0s0qqDo6Xp3TNbTfprq6D9
2SDY02grvtPK6+bGAQHIaJnVfqEFZuCzm7gp4LsVwfH+5eP+H1RYpW4sIk3hGgNYGNomvg+a5BKT
NXOQJF/bRu3N0tKbMYzODyZz9bve84zf8AZ/mgLA5OclGRm4EEmdDo6g5XUt1ZUbaeg85OdmPRiq
5a6mG3fkliNuTWmn3L6Z0OA47kkrxmDPR1K25KqxO1Z5+3qDwV2N4urEHUny7EkFJo4LsD8G9pIB
MirFb6+2eIQwkqWbbpwGXgOexej2Q0iSqJj3qPhp2vAO/q2NBmtHa+pj7CGtFwt4xIx0T8JxIyoN
RNKrMrCkBenOjRdAYQPTTSEQl/ChlYtd7Zns8pxKVnp6kNMgGWKJW4pyG3jKN1Jb9nibfdAPk+sl
scgwMXp+I+QjNo6s/BKFqx7a18FHZptR85nm4gqyp0ynMkFP6/cvVYwzskFH1lAAvwj629YbQHMD
JALlgQE5D3cIbmThv2URopta9wJcHDN3D4WkGv25gYCKYqFbIkdOxNzRx4PxH8NuhCAaQRXyPphC
FpuTeJvpagueQwvly1zLAPki9j84AuCGq8zWqCrBR302Ooe5d/w870Mf4TBNsA+AwxlHG7+WiHq6
n6pHoOgtfDtBwxwHj+Ei6dlcIRq7lV3hGMMACwj+deV+OPqJiJL5gpetFsZ301kuLnwr1s8/u8X6
RTWICy4C0Fr71uYyw6jU8E396fhR25Dc4F255ZmvdszxtnGDi9Hr92r6qwm9NvN5+s0llIXkBR0g
p79e0ZHieJKFo2XRg9ZJFxWU1hq3V0mVXZIUPhwOQz4MoiPC67mxZHbv2I1wFZVA2KySD75BdlXE
7GTiyOxoEfKuFzQ1AqNq9xrASAZJkq4jyjeDi6MPyXfohCqSWYyEKQSQuCHgkUWeAQEYh/qOwoIl
0oDcsxtCy42Hi17dxFliCRk6srxb8QguGQMVbZxDFWTKt5/cbDxEV1jKWxJjziaWuHsqETOwglai
LY8DIc5HXoyM4Zwc290LE4ZzxYFNAsZFWqPB0utBn8uoA0NfoCZSuraiVzq/hUUXT3ClbBiGasf4
0gdLPiVJOlXGbj5372AX5C7NrIUjQu04nkGcBeKpDTtSh0UYCwnhJjRS+tDTv8W8ZYbm5Pyh+ISC
+eGjXlMDsMidk5foIyhOgT3EIEQunfxysfZa77JicwZhlX/BpZpFIf2aYc0YdCoHLAA4iwfCp4kH
y91SnpnD9OGbu/kYS+H0zOEs3Dpe2ZY4N1M463xGT4iXyjagSOHVQE4TwLefK3AE5d11vKbK+FKQ
D2dnOrOidv3RdmQ9vgJg8JSm98jU6MJAuGNHFpKJLVRDKEbX3RQqPe16xVPSDNdCV54pDAWoqi0u
VDK25BOxZhq0D+6rotvOhShkBnSREwY2e7dmPEDr0xB5TGvXGDa8mUailM7KJ+0lPdjlDFcTorYg
LWMT0y/7JTi+FY4oHXpjJKcdIKNxnK0QD60yxCDKU+Wc5jcEhior2Et4PnDZMVq5bXgcNXF9jlLy
pws1K10JPOiGW/7dmDgTgJzLoM2usysC48FFy0btleL7g2780Yq0KjZgyO39QJ5QWPEJroKFP4Np
yv8g/eHtM2u/cGNUQ+6rotN3HupwGIHTJHb856KxBvF6AT/+oKPjVPlkc2ecDCwRYp0Q0i8cq35d
Vh7JRB/StMsBdeEXiNUh/nsRvQH7P2sR9pGyKeh5KSw6YYwfO34F1H8XlKxUMiC2ZXfagMQEBmZq
onuDqu0TSgZytyojBRY8kX17rFilCGWr1nhcZCTjx5a5Uk4Re9pUlmZ8tJdmCTQ11RXVGDzBOKQk
zI4MGNkG/cR+hS3OOoy3MuuuIXVSwhGAu1ID2aHODMAbowW9w+NvWxsJz+ihcrw9Sa9jHx4bIW+c
CbRXXnJgBWMpcmJ2f0y21GrA6cDPnCYmReWhE6n02T5r3vLkIecr2io3OQDZtZU6hLPkk7BRT6BX
G5LI7HbPlJD8LSP8lovDUYkdth6jpeukVLXHMOeGx7mmqZQMrENu4qaM08brUFaOKJbYrkaDVP5C
sgsrBMIVs05MJUUmk8K164awgJnOrzlmUC56hMtFoxuY7pCqB7LVUeWq8iy19ND5Nz7luIvLpfHH
qxaw1mStdKVbWQqhj4YP3DODSC8M419ObEBRsXYfFlb+tuwY5rZ/sbVEE/yN4gzEcJCWkgxamVY8
ZDjaNPiWve6GnGhKs6ELYzwajhPWuYRJxfhdtDhkWIFxqYRA9LCpTt1FYcZtI3WHYUfCCb8OiMyM
8b0iGRcVOQ5Y3zP2l3N57jz+s3veT4IC/WDxoqiZKn2TdFI5wBf74ap2gs+7WsnnWNhbRAl7wzzb
30yojYPxwzNGiPcOUy+f5O3mejOnQsmlnred1WkEA68gAEvCg6wsVI/9aKbUXdCemzN9vWrKXPFm
UgdWyRfzO6IiXVbrYjCkvO5QKjsMOSOPnrODzXlETK4Qufx/Ii5jx7luiQWG2L63SIcWBsXycLLn
anobq+5eoS32doU//4DbmzchIcyVjtDt1RA2ptx+fNl++9dC/IeF/fFNlFJIFdxUWodPb5/Oew4y
C1vFtBVU1YJHAZzaGh5otDzrtQ/rIwO1k4TDe7Nu+K7KVT1z+3vVLlsvZuj+SHuUKWaKqPYA1qJP
UMUec841/fXx4OmyzvZ2aT/Nk+HmmLLMZ4Eevb7EXPNCfHvnmofrLnUjbKQIwnqPZSCcHQCchsfG
WipWJHJ5W1YVAVVy2IBN9pUdLmA58EqhZRgliAMqxl/w7D9NLRXhUTFizntf08m6A0OuMpjwAWJ7
XB/Rtd6k1BL6yUc8R3xWFSNhnqrsbRVBUKvrfWoaSEbMqb7dPMLQWRraicfNJpKpNUv+6703FWRx
oWrvQoYXSm2cEhzRiEvip4ilHxrRy64DtyoZOhNzOkV8lfeUq8Ijkj8+5/WV7Odm5Fx78bic/rW+
DgjLmCXQLep09uOBcqVVMF8LcTV7p0qIRSqkxhGA9e07jtxRNptbTLVF6x++T+XcwxShtd//KkNi
W2qVBySWcKFXStCaW2vWBFtiV9rwt6nJnOsa/cPzFJWAkc6OlViFkBV4lhZSrjHWmWtgX9h/JpyW
EIg55gKV+sGPzq4cNeaHI6UC+mkNMSkAUz8Lk9EVKf1mZWYCtbGMX95YWBNWzF8oPEL+Ocv8TH9T
C48tabYrHlSR4ZZRW/plVOFap8cUTqI2+Xh5aOAvTnvoR+ZEvrBmOB/wcmDgyXru4PzULb6UsoxJ
fTkzxEHSLRnOI2nuyklg+NgjmnfMVNtPv+hpXzMmFdY/JAXtH+x6egdzU2mwdC5jvLGOrJiJKTEQ
MEIyhebdKKzCZ0FqRQQroH4YU1JiUeSu9XlhNncUUpe4bLJNiV/rcgTpoODRWdmaZS81AWE9eMmJ
xH96iNjAaYlVomWSD7cRVdCu/bUiSsJpARHmSEOMjUgUq17TDA+12SJFuAFHfR+plt1FnOh99m+K
xyb82C+nhMmAhsHsrJ0qtULpubZ3LQqwrdvMz2QhsCbicHsGnEg1bsR1Bqzb4B6hf0xk74oWLhIm
PA5Uy5I8gXXe/H/oS3YFF12ySg0CXgfKRGwCgxxRcQ/ZCIHXKqBrjK9fWAnLjF+xdw6pvdrLm/ZQ
hDQG+prW+BM3uIj6JdqKcgYtqqIuBKkWIYP/io9oQr+U3qtmHXaObA5ATuKdvHofhX0xx2U6KhPv
Ff0fXxOP+PIn0yB6KQE4jJRJUzsWUMN5agX6+KDdJA65pMFALjrh0b+75auVrdDUVMahgU0Zpvcq
Puk0wcAH2as9mSCMgFX3xkcLt4oVDuo5iE5YXnZ9/dcdVII2g45aEvAB1dGcXD1qKeMa+QPmc3jk
019JFKlE0hvIjh26my64JrB19blRr7U1qyJ9GhUARK3YfY6pTUpMYml7kr+4xOdZB5CtMJYzj+4w
4m1jBw0MVsijjA4akRm3ZEO3gG6fhHkEmNIrXKL4t1EGSqkYK7ItssdEAHCds5wf0tyUVzizQyCA
acTZJY8o8mXZG6oqVDl+RLYITLr8vPEFpKiBx49gTUoZG9TGEd/f586xYQJ/XjsIE9G3RudoGfiq
cyemBrPJ57MBUhdZX97MVJj2ebpaNGTenAjafYF+fgrTS5cXyowy5yHTC9SWKv8citTekrN6BuLa
JGYGa2f/pZL1gvUKbWjMrRF1dA1pugtbDSuGNJMUllD93egwEYhB7wq7juFVhBVhBsP48AhPRMxh
XzlbRyiEkaIVHwxzSm8w4adVn7Qmqb/eMvQbLObcj/R94boMchAJG4hyBXmyJ1ku6YCuadLuBx8t
1gZEVM7L7LQ4pc9bwGUWlxgo7kFh9i45HRd7wJAWaTDacskY272z+16txsa0bjgXs5ek5gBzwGSL
3PKaEjmqAk3kCl8GCJLvgkXbK+H9Uz4EAg+s+fiXSaoO3ZD2UaK9Urqb6c9TlgB2ZstrshJVRONX
0gYaUE2zjGC516UL6Qw6nBPvHtlKF6bL4xXhMO2DRSfGNRZu0qUHaCU4F8ecLNo9HeTl2kwPjaqN
kYnOXXNUl4mMILhwlpKWecYBvtUexDoh9aEqK+zcYvSs8yKGIIfKl7oAsYAGFY1fzhQrv4oZdtSE
zRgYO53A15SekxseUJZpddudYkt1bIQqh4cA3bYNX3Y7xdato0FNk+moQAS2Npgq6cnQa5kpNEHv
E+S32e2MMmqR1JXNqZx1sXxnpXtgBoL2zlOALvCk01SfxTBw9J4rbmv3gt4EhpDcwbDquuKvGarn
MwpeLd4646xf1NQEoNFyuLcmKAWk61lls49XMz0BBCgeU/AszhNV2o/eiRalPgW4zH/2b6kD5DAe
ji5YzfFYC0i6MCVQl+ps0Hcty2ODxTZNIGfzALg8tDmR/6ojynpQUiXLjw93k5HWyieV60+Q1VSt
5wXeJhTyH7gnu5kXbNiLHKWAgbmLHp4O2u53v9mN3wEDkgtLYYdtOz3fCaMhwNSf318PhvDRrokn
16V7FODLp3qLKmfPZlC6mRw+RKJ0AqyQtzYMPX0NkwVC75wqACIppZHOYTjcwKDrvMEVbZ69J63q
jf60XA92CWdONO1kbe/RVJ4V7acwbAspr83ZOFduSAK1ZUs2Csr/DOfqq5Gg2WznXk0QH6EylqO6
fvTcze2kIKOcq3C1hkehW2weK2mW5ommXuSMzfyklloddWGkzX/QeigNyr6nI82aEzyH8po5BBJx
aeJFa29FvAZh8ZOFzuXNAfKiMxljobrJJ7AoFD6/vEjh1ceoYLT8VBTTmXeG6ohX+wtLYkRe5vgt
WBC0LrAsiaJa/P7+OQ9JLBimkzwsJOvpUikt/SAdV0OvxxwxAqFL+JFEaX4fYc5/DVg7W6BNRKCO
6VX7kvyx3gkRmRhgBbsU/6Xg8c/ysFaIAVFae+10uVbY32jcvPbagpEOczu1XRNb6OwD1I4oQNwj
+0AhQut0ukfGqyevkLroFJ4MLfb3k7AytwKuUAVDvfoAM1hpgk09rKcCNFbOWKhc8QI0Xz/4NLYq
PWWot6bAaaLmz3RyjzjTUbAlVSdMbQ+G4fmVC9XQ+NvJ+PJBHD4qpGwzEVvIM8oO8l6Jyj1XH00x
g+RzzZPtaLrzaP6Ac7oROBbk1yooiOEywP3gL4D+zlzxaykCW3lH+y01D/CK1nv/svHgYQ/Jxbmp
eBWdJNtVr8OXjUPhPKzonoQqq3i5GYBu5wT0C8X5tDjLxCZqnmNXDRNTsWzvdMqR7p8yALWFHezH
7m/05cYoB1Tz9FJVaLKO35gP1dT9Xd2IAKGh5qlxAQguyAeatk+YHu9ul/lWM8TwHHRLP17YPbVx
uX3SZgviu8ZGAurupdX/k+024od1ayDoHcrSFZWC7k0m1w8InopQZ90m/yid1EY0MqaszC02DCe4
GNSfmEgXSotzsR4H/tSlvvyk5d+9xfUi6numiZ9FeVNXH1dpQKC6Gsv3ZtQnr0hqFPbH4nzpgdST
NCvWEMOOpmlnh2qcuAWCb1VNXAGZlPCyXG/uH1eG4+vYXTOC2ht24ifeZtd41DvZXgEYprtBbJIW
coD1JFgfa0U9V8nlz7ILLn6CNjW39CM1zwOIIO69Yb1LeFxliPjRwOFkfkCuTLBbJSoEN192UD7F
22222RnR8CkMPzkVD8FrRLJFALCCG7uGGNYuTWcg5rxF6qP9tQz27zcFVW0Orzx2KSuihhBtaXf9
KskcOvTQ2q7mRYJAn1fDCc9QpJHxDhYit9EtpK4YZZUeyd08tWNiB+eRflcRGzfvumpRcy7DN3ds
f7yWC7W43fXAY1toxzvWj7O4hDip2GszDjWKUVTxWsfz3fBOXsLdQZRXmH6+V6AdrGtbk322+DPU
9OTqDhXclBXIRp53GvXp7yvn1zL28FTlnboP9gw7F4FV91ZzUIP8tcBJk6zvk0Xq1lMqw3bItEQc
BO9V8YN8gQqTo0/7UkypVV7+1nvl4H6prEWjucY7SF4GYXQVX7ZeGdSDqEQ8zIQiCNv9vWVkUlq4
GYOxmYk4dGpNJOKR+LW5exHpbVht1JZoHjblWZtWkdZUsM9MI8MQr6n+T0KtzgYA5lXALsa5Dptf
yLw1r9+BybMVGAaEHblYx8VHOSZvUMiZACj+hfo96tuFNZZgTcr4se4N5SZ32aqfopBf1kodVVS7
dhQMHVyb7eN9nPuSKBFVVM6DWS/EwCsMceB17IXnsI12//pZV9DleBcMDl0PEUBZJFgtnjoHS/X9
z7Avx5Kkrs7xqyym7Eb8sG/wLR3IUFvweEBCvNIsNzw66lRvFcENsLIA3YW5SCJO28P7DOxjCjSS
nmZc1iypeOieOl5uK7yPQ8/ou7ek4pLuCerp0XePkB+6sWXGlOojHdS8QdA8JaXP6VcFSGPpQy2S
+zdr3oN6qnn6q7a0lm+3rkNtU06pg1guSbZnIhXTJUopxHERqE0tB6AU9OCTslIim/WHVYwq/JTf
ciaZO6vQrQ/SUz1fmE2NDLFn6PonCoOx6pYTNPbDsaBqy7RUwU8az8cAxZP8j9OwSLUvvOh+vuWt
+g8CAROGOfbAR6cSqZVkKmincoDFpS+S9EzxIbN3a+xlnIjFOVwZ3Br2f/IGaJOdyk0Q0Vh7jezP
S3Sf3c7k8pf/dZciufMGGkEoOOuhfC7CC9rUXdXxvFwer3ISIuOtyqelZDQP96/0D5iTj6OsUofO
QDhU0533Q52u6YbtJlZciHzEer0OORXKCZtpf5jyD3xSKZM8TlLGqA6VKeU+hBaIdiMzilXSz4uM
PeToniP8N7barEv5rVd/N+rVgesp83leXt04ZLSjC3BozG+5EVN9CKNctb7g97K2fEP4D+vXnTF/
34h9gSVxzoTmFgpHKLftrkaSRcsBh8izsPuhnvSr1JYqIPpqRN2VUA0lNZKFmX9RggDvAbTwyfAm
zxAibUSVazSRvM4FJBlkzc0xI8vZrNGmeAEyOzRSvSM3aWR+lmICrCeEzp/J0i2LLYjhKB29V/Ob
+RgXXgVdPZl3bW43yMM9Z5x3ZpNmHf+5CVK2d2lewXbFJ7ovkDvKao5fc4QjLgbbFLLd9e71Lt5Z
EjxtdBUOMRrlSOa/sesI1S5iVfpfLobTQJaN7MMBtkz6cxmS0fvaX8VtnVpfSGWQi9OvWT+DYxVA
0xLx+YTgktAFrstLjbwNXmnzBcLbSSkMq/nkrziQyvFHWBAJbPMsxPs4cme96m/a0ygDX8TXMdEb
kqASWgrsTzCXBf3yfsN6HsVV1hWzRnxpZzH51kNZfh4FLF+iEvCC883AgkVvy44s0XC4n8pc6Y9k
w48NQJJT+VKuvHfk4zZM6Mp9Vv6coINTSHOdyE0t9EuGLzdMX/FGzVXLaKvuqXIeNx8LNhxvQf3K
k1APc01DwAXf0bG/4PtN/4XGDRASkY4Bve4EdkEyicVp6ZAD36+n/gC2pJ9MvsvwN/YT6gA+geYs
1/Tl61SDF51ajowUb2QhdNQxx2/QgSD2i//til14DosKVCMI8IFSe8TLNLfKKRAHNV3u4hMTL1pm
RrZrmmZ/4rzhHs1t/VTKuREjsyd9Hnv/O/KRQwWHHaR/5ee+jIHEHvtSsIAbSkdBW7rPHCro/GHT
d+TaIkgChbjD4PhUub2zqbLMVndCH/OvwVK/zJsyNdobLe0lhGy0S5JZTW8K01nJ8SoieJzQKUMk
97d5NExgBCAXO96icOZVojiRjBYK8Ry279WBOpvI3/VSK1W+X8i9hpMnqH5ck1dbpu70KsJrZUs9
e05hG08OztVsg8V5dUao4dgoxPM1xxZbRfTHOiMVm0OPoX7N95iv+UgvMN3mW9INJFGmIz/I3Zq7
eXHInvVMfQdTqo9zxCfrRR+4HmxlJziYACBs1B0KZDJsaxRC0RXE/Pj0g9X0V80OrwSdp6vYO1bN
obameSCo01g+EyahosGVAhMfcUggYPh5mRL8JeuK39gYMPiFr68hs7uZdEhPnbrr1eu7ZGBKxq0q
I3hIkw5Gj8NIqKTuJ66uq9xipbtrqe/Xlgl2xWNsg8/tzsuSyjJCJPbTXbxT4xn9LvkStC090qxR
lCwGlfN+E+gX0SsGfd2AkDRwHe+SBbkTue0+Hr/ek0C9Zi7beBq20uk3XO9pG3+jLnNjDM4x37U6
WgLtUWjZheZSi+ITR9zn8cPHYK+pfqzH1MCAezZhGA6AIR0KeHWlru1OyKN/VgT+aL7qCdD59h0f
w8CuvALha3ssTs1yNAFxw8SGnEF5cRYxZGAWtUSaOwhJGpwCIFLFtWhxf4nLjMeO/BHlsBwORGbB
JJQFsvWv92LAuk/oh+c5Jhix36pGJr26rxxs8SQ398GtE5v6/EkpudTVuoBvc3O/gUoYTXAwgTZt
Uv4Q02mw9HbyEUhZOXwVjQNzpqnksqijGus7eDnKERaYIfZfjoP1aWLZU3GLqvCKLdWTDBDkqv/X
uOpm6w4dScDCQBZJzYsUZ0lPvHnoQtQz1B5D1X3mg5atpOFcQ82jd5WTf0hoLs48QqEEX5h++Vet
AxS4kUNqYlmKsPcn/znrs9JHWm8zTOW4m4qF765cQe0fvhJzrdy2ta9mreMdyuYPYWioFj82YbnU
XaeUD8I/OhTf3MtqPY7D2oq0D8HPZDfKOn8Ds7pNIogSBQVX1ZDnUY7BPZyb0BQbme8A9kj93rOu
ZMPRdH0U81N57VTc0u9TKLwkPdZnGslHALwPPovGHkdrhASQ9T/sPXuxYBY9hmhmszEX2mLEPhuH
DuCuZLlEj0XYDaHhypa7qFJxgZU4MxqsoQKJ0lbVh+v5YWwxolELXoykB10/5ETrbgE9Yxp+Xux9
2J4+E+SSgoONN/5U3POb3hRejogP3oZi1zBwMWDQBcwrbyUTM8shXJdWOB8gRPMXgaJWmZA6H3Y6
HYGpmRu1HiXnE3RWBrsDLFWVAKmuFrNcRDEXQAwmZNYN5NvNY/FA5JSpkVXafNb+a6LpOJoqfixc
q9SOYm+0+UvMTyc9o3WPpFVZ3JH0k3lcT2gagS/pG79ia5iAtqGRh6qPo6meTkoJuTkq94nWH7t2
KVcQxkfP1gwzH1b6UyZLnttoXudx2dr2BxU0W3v99I9MVykLn6RRi+h64pUIO8XbgZv9zuRkaYUT
Dog2WMdPx3fJYPuyD/R+mO9Z0rZdP9B/6S2Qubg8661N3kSiBB8wD2YnSgdjBsICMHHQE0FxMXP3
Fi9TfGC1BR4tBgqKtHQU2gm9b8kly1L4KiN0wJHYRZybWO9EUMzRVwHSF8A1RB1XP+ArffGNlexn
7n0+HCq8dmaAcv7JBFcD065effzpGsrGtgBFDw4AdDUSGtVQHMP7Q/njHmwW0CUYoXb26/VRcx/D
3vOt6VMlTkD3OrPERgqPpWXn1CdHgNv85ojpIksjxpYL6kWh4a8qIllw7/B49OVVTa3bJ6n6dqdm
U7NkwKhBvz6AqHqhy2lGvIWmuSRDl52D1+dIvnb8ZjUEZNuFrpg2bFfIXB6X7ax5bfaoX6x0tMZn
XN8P9p5Ql7qMTk7BF576iDPsfT6yOWvv7Qxfdr3zfMrAtZLU/kXfAbkYm6ln6rqIPcHb9JaaCZkL
1UbtbTJLCDgCvAQ0OHBZiQ5lfnb19LBq+V9qdc7rI7t8JTk3n1sESuoB4qYIS0rd1Kc5PpH8t9nq
9If5XZUQfftiqtd3DbbeFeRa4spFiJB4OqTiFHTibcUiyfUm+oQsWqTTgt+2TgO7wxwdXM5g0XYF
MyQ3l4a67KucNjKVHEO2CtTFnmT0EU20XsCGto+ntmEgz/HEaro4A/Ul0mwTGOd7cCXkl3IbSx9u
fO4v5OfMUB7gOvsGTYBu87z4W0E1cZcqAzeAaFPx9Fx/vf3Ddqzo//5asx+AStvG0Z+Ut6fZ1GxI
HGBhE8Hz0tCU1eV9KXJlwopmSlzbEpHfuxInQDuQTrZESHJr3IKI1OoCADrqdakAps2lIVsyXKC1
I5/Z3dY4bRA103DBaj9vqUI+nR9azQmRcxbewkBSdImkH2QohOc09ILCWpmjLnFhWgDCNrT/eoXA
s+relsQxFmKLN7ydunKc3msTWX9+HbNF769F4nETfP+dV8aA8729VMRo4WqxeExKBbFbxRGa+4uL
fnUnL4SZsHcnpyNf97xtRfc0q1WACIFrkT7IsgCtvMZow/VCLh5Rn6aBmlFZEzBmkuGHUV3ivEdO
HT3LII1pk2V6BVglb5eMg+XqVlKYufri9zBXtPNVf/Bgs9UtZCokVVN/VkqHH5jWvFDyTWbOwNnI
//aqQN0EaIc6KjngfnfKWz7Us7zlkas00OfBODr406FpN196+16I/+hRy1nrCd/qJypEMzQwdMhD
rxVahs+HZjlHlz6wDOEQiWynzGuFV6xRuJx6+Zeb8qiFZzGAKbh253jaiNg6ViqCibh9j4LgzFXz
dlErmvK6AnOdpCGoTb0PVKXEFkZYEAu+Z/QIYrW7mEDwCK+zD2/c7J+U3kSY6veP8fSLOWCtDbF5
5lKz0o9n1XBZ+i+DJ3lrCbPXsvhAhUZ4Jf948SR1iwF/DEuBfXBy28ejb2V7z2zzVuPNl0h+7VZu
hDREp/4VxwHcQP4S4wHw3WPYRz6jnDF8aGaEcvWcKH7bZR/h84TvFp8rzO3wnugq3NDhEjDlmYRl
2iDbKuhWVZvC5QWI20iU4GOjguyn5SitHDH4zAlbqEz9D4Vv88vd9yoil2zBKT6d/p273MqrHL9n
ZwjeM+4kLMwGErkbh7/wjm4KuxsUUAXNYf43dI1C/eJZ/MCAR/41NcKOz31pWZW7PPy2N8++fG9e
pFK3Hmdpq7XhAg/xQDAhMe/I/XhErk+4ouFROaSamaMT9XlAfsgzR+wxjLXK2axTAMrMjIfHVlWT
g02PpMyvNb+PoFmwchuV94jzZ6uChX6M+KYj2Hy1xu7EE3UjU68IreGtO9fML8DbBpjsPASeYUuh
IcjfcQAuRiK5hEe8jeceDDoLsiN3YzpcHTVyszi6JWzFss/pi5Mlqv7A94tLIO3FAJKCqXGfx1k4
gxQjQXONWCfsVaqHUHElVHWoJQoJuodcggZcIUFsmjqHrX0wdZSqzwhBlmaHg+wt58riLZF0Ry0F
Uq60Lh3UBrUPzS64srq6WQxrVc167KdW2U8R0SHz73egQC4dVquxeHDCVEu2cwS6JCJ608Z9FXAo
SbQzk4z5xkEki8+BsDGvkK2iSHMvJbF705Jw6E/QBveVbhBjS+ZMjnrk1GJpxdryDSLVr281N5MW
72R2+r/3z7GV/Dn+pa5HdW1BRD89wzqgEI0PPTrnf0Jp3na1RPyN7Y/0X+eaq8a6Cex3hQzya2aA
+8rZX9idsXd2H35ANxfrvPKbq/zhZ6K0AYm0Ttrpgpn7jQO4MPYVX3xRA+XCAYHTfjGjYmGtx/iE
yHdI9vbrujGDXDXP25Smugn7BetmM0YWwAD7kQunx5qlyrHShJXzizW17y70UdsgCqAV8qm1gnbk
mFNRFdxRjepzfRel76Ezg3CiDcLV1EfH257tRw08Nl4+WBAxNCAh4JgIKYlBbZ1bkw3f2jibh7qU
p4PZz7KhW+CWmw0sXlHgk+u8uxQ8qGpKOI92GTItrjHHMe3WaLf1Izk+gDwTsFWGVKcDIphJ6e86
KVpyiuWYJV5R6/l8+hZ9KhQVbI3Pz4Pp5uHCJrADSv27CDi+oEp7tEHXg4b4WtL0ng+uCLLa1mnp
tG2MOB4jhtDwyMDCihlecvv2+Zcz7Q12IMD6yAoYXBVRQa9pdvS1usM+6+1PLCOQAqQ91GaagBbH
oqYh0nkq500CZBidkJaqUxW6Dypnq1Oq1lTf4mR2f00j6b7U8aZDTYacH73st7FHg0L72D7mtSga
EIib6CD6kwNRiddb0pjvJWnMiWADt/C43zseT4GH+qNByd/oOnRyMbmCNyRvJvEIjhl7haQ34R6X
Nt/A/HoEa7MQ8tPuM+M3GkO+I1IqOBZ7FqfijYRfiD5iEnUB+UHE01jvisPjJuwRlUw0PStgoH7O
TiOcr3pX0tutNafNqsiNSero/0/MbLxelWigM8XgknnTV8n8kPcOrOcJ2/3Muj14eTmVUbqlmlT4
CCjF/hq5QBxY1nkfp3J7qXb5zkXmzhBtmCFsoRDVijwco2vMVLC41uFT71MXLKNT+fn3olLWrdZv
oYOTrg+hB9hip5CQ9KE3kh9ZeKt2QMDhwgORPutxXV5CSU5DSP0gpIWL3+rYUtg/4ZZX8PZ9PwZI
jpv874rUf/WDGpuy87gYLRK384gai+iyei6Nv7LQeqjFLnEhuhZeYkHWZQc7oBKiQb1HLE8A+H9K
HO/h+OBr837J3+php0t3vt3rZy7NvhtRncMNFb3NTlVWAYUWazJBGWf/L+oIqk+uRJ8jhkrejle9
HctEt64rFcqYRDTytVYxwNnn+TmUhBgz0BoFHzaF7V09ZhQs+xHUOYmZJcEv8thkY8oTJ8RlLfgP
VHBkkq7TFhSFft4lpKyBdQfP8Y7NIrrosq1RUVnLWw+5KruLY/VIQ5Yrtncm+HkHvGwIr+lxWwQv
pnnQGn6LYrlRkGklqtRvJ0P85jLay5zrwC9VmfLvK3eyPxvloONvwqA2sj4Hbsrzn9wHyk/49syv
H66WSKQjycFUrZtddHmpISqjq4/wHlW7kbvKw2V3SY8nMsoH7V56xCoqJoZxt4TGi9hVtomcRc+I
hFDKU3a9u7kUqCVrWWgLssCuY9nrpU3XsOEKVzFOYouZYEvKVgvu0OO3kcslmmnNRjYs1ZJvS+DT
s3QySrWaVsz/KweNPvDOJzkmxJR8jtcQFoKYBnRwT7KVK7C/r/1332UE9aHuj07/6AWBo43Uo2MJ
nsiGwCtX+2BK6T9l+1VzU1u90F3C0b1hn8ZD3yQrYIE8VFoAuXdrrdI3gq6YSOFg7k9FwGbJPBb/
hZhPLRsG66gsLt+hdEeQKJdpkV1O8MrL/LpWvjXUOwbsDQqu318y9sUdJ70vrCWqaAxod+nhbAq4
h6NWg0uXTwuYlHm4XXIzfAvu1JEKpGXfCpMx+BUOIeTK+gHuj3FyLoyFXE8VDn0u1lrvF6Oru/Zs
c55MWMR38gJAwkwYkRPbpcGjyEPYEEo+QfNIvik3lg4sqvxZP0elLLIb0Ybrha3UBLH+YS0x/l9W
Dt2nLkFDz7SLxFm8ixkK+xyAHJsjdWjBO8i6gJX59JN2Lbo6gcajSDHTupooa+bvb1lGfdvENJio
n0EDjVpifBZo83KQUUzzdtO/u+xCzk6qQ7ZEX5HeHll3jyyAWci6puXe6EgqKl5ZgMVpztMd3Ye5
yJLWD95Jh8va+/H7NmnWXvAimH5wsTN4AD7R6L034nMc8P5yeOeaWIiyYHxhJ7Iv3e+D4qS/Kmft
TRdjNTpMpElUb87l5wmpuxM+ilEJsDATA+JP3Xik8Y2ZE07mHCRBq/DzQq3yTyt6cZSatXm4XbsH
as7E3/oK3DN9a2bh+4cadcEH/+XuGYKCYZczIb3Plyk2hQLd3vU6X7gHfyn3NHd/2FuWLI7fF7MI
kNI/YA9hIzBJtizuHRjcMx5z6+aFU4fTKKGyTaBgdTP8uA80ynkILBUFesyXl4y2dW0RugsB8u5y
nahrl4NQLP8mlFr6GB29R1cgi2FU7Ar0KjQ51BHjLaWk7/zqzzsjtnUMQgieW9sROkmOE0Stasjw
Qg//f2LbpGSC4+cU40KX6AvyYNgWprDhHUsufk4fpygX8CBNSLqydklEdX5LIL8ct2isfEAgNM2a
H1AUS/lTHipx5ojB8PDfyQJdbr87+Itj5j5iCmKlLkPnZ9tByOzvzMZscUx3/m+gQH6Jx3nTJ3hb
gxHismwW5PpmLJBohBKG8KA+k+dAneqLUoredNU4+XWiw/iYWj1VwxfSQP4YvgB22B30rUKzOvBC
a3lW2BMu/NLEVNz+DoMruNUYrqQkEWtkcB17t6KgaSGhaB4zKlbwrw3i284eizk40QiJIQ5EhzJj
r0gc/p8WZSn4ShOqn69FwqcePDHlEsyFoQLGfi2m4NZzN7GRqBpZy7q0OHbzx6wKgpyo4fuRVM9J
+vygTGKGpZCEjkqYalRjYekHIUsbRJ32t18KYU/NTJcxr8CrXlaTy6zjUSwsG46pxhq8yoyUF8Cm
sXeOg1/ETHm8e3AzB6YvXyPgupZ5ldNjnDAm5jYCChJvhS1VNDzdcapYsUcL0zrVYfMkrb5nX6l3
JhvJNA4Q3GXJDOq/ttETFel5gcMyCeBH4P1lJnBlwRTm6DRkg0KXLM38ReqLVK8RNkI3o1tc+fCZ
/7LPpRGIshsqah0PgBTvn5WE1ZRQ+fAOYnd+QcgGpST3i1BvRnJYnIXIshLMhFRwcBJK1xFrlbvI
55ggOSWsGG3pVqACcLBFEgg19fUld2/9pOm3EuPbTCN5lxMRdFdg++SN7s17FZ4NrshYa96aFrq7
04cI+JPuCqHIs/K5v/LMuTmw8uBMzg2lI6sEhRB3bYKEPTDGNYFCQymNs2Sr6jTB1sA39MRxbTFK
XgHa9XFlp52ixscuGaUse9M+iOwsu7+3pvbo80MIknJBklP0amC9kliuLVr85CMoVfW1AXDfgaFx
Oi++PK3mClfyhCWkjOOtwXBUPnzdZQrj+rZYLbrZLrE2i5lFd0lluJ2/YdI9VJ5CF2FnCc383TI0
bcRcPDMR5kCfidjKi/4wlTBAehzEzEJp6saI1Z5XwuvCBhDQ5HMB3od0Zk2FimQAlV6x58fBqvyX
O8TrkrOYt7qNXc/Oaog0N5QkUX3sMQ+3qTn4VV2OanHm1dn8Mxgnbw8LWILSl+ARBKXTrmX3++Ad
PkXYdcgvlrNyZAUyqaIwxQoI4eSlztDL0+a4krANIirz6HPfctjdtfK4jrgerSpF+wu5TxEeMq3y
Q/fOV0tySLVRqUU+dqR6gOjR55UguJ6gB6HdDN89gS/00/MbWy0ghsro4BzxmlXGFG5/n8C+eNaF
PVbuxZkv5mc29toCXpzsadfwL/2BYHNDth6wsAg5qYuEEh3Q+ZdJUe6MjI608M7gY8dST6RX01dR
LLVYRYkjsCVtdVpkg6PBxammeurf60aLPhTfdzLj7p7cGxcbzD7YMiucLMloWWobO+kxzSkOQtlY
33kqRfmfzvd71K075GTRpki4YPdL6XELg4KpcgwGFl/nTMsJ3kyoG0yjQw3yBZkuIh/+djiWqHkK
30PM8EUU30S4whH1dbLZqEd0A8cgTeeIzOylfUIprw2rQlRojilKVEffxkp9Ndy2hRjs6Wb0bW14
whqmB/7DdNbDgp85A4emFqd/eIMR9+D10cvpGhXPjeBsKy3c2h4IWsXT/sQ2D7EoBts2cL7IS3Oa
xKzGJX1w+D+NofQChLzoj+43sXOsPAjcGUEl6L3xbesMj3PYAPr+Fc00uC4fJjTU5wTeXccHmqQ9
APeQ6kZXIOLTtfEpFjPCQ05tLEvVs673hljD/fLIuwQ7hLtrxkSZvvWy3uhdc+CT9Cft0XnAb15b
v7ONAa8TAfYWUTQX3gBHpFyBFxB7D6DSJTMBg7hbsdlEIBWV1QEGBUZVgsq4RhepriLzYMlHwj0p
fp/6JqGPhXe2ttANPSrm5AhprNmZ7+zMQ6ehdf7EFnBDal2fMGe8tkS9XxhzUxTF1m/9rojDUl4a
jqu02mtFA14TpFOM6A3ClPZ5LJoQWJSFHPWWgObmctBA1p7HH6weF4FhgETWreueQOJmkaWk452q
BaQSKLJZ8/GTpLgCPMarVk9bPxM+Qb1EnBPZ88rb3FZQP/UNfaij4CAafwj/0ucJ5+XjES9fTDcm
E03m7LnUqdeQ07C5zl9MaVAweVzw0gfFTBKgPcYrE7j2mjbDxFMCUNARq8+hFvUuL3g9hRmHbIgk
j1u4nuAtaEBEWWgKWOQZej13XBh1D5/t6hhqgsrkDpSDw4KAhl2UBhVN8MGjWknI9QNMQ1VVTR1G
4y1VdMLCOGX5ukDm1eK7mJQ/3QiyVeJbOaW38uPdf2mMgA3zQLL53KjEYyfhTYEg9heWZW+TYzrK
JFJLKltSsHPE54Bx7tAemdcRKRjEAuYy9tAhUtRHeWGSLCpvgMVgocotOJh2lrq+2t8zpK9TJX6f
w0Dtvw2wALar76s9f6sOPY21TSW6Bez2wNV3C2nRik/HTNlcml0G1nhArqHz1k7lFWefNrNc4w6p
dfqKPSNN1s3tHVfVmvAAzx9d303VliP8AcrOdxPxmdqaJfReHW/muA0cJl8GglDtja1F0gZpk1UY
RC4BQH1nqJ4icn7ynB2epUaCKDlOLo+zd7QfR5lqofwcGVldvmr6WOR3UvIGni1B9MVoNRbsklzT
Z+qz8jI7/uFNtCm9IcQpFTsMyVT0eEJVv+eRm+pPe7D5/VtHVcE3Ta1c/JL8f+kcpSy6nX+DuK4z
WUbtiWzlhiF0IL4UoQdU2TF4o31wN2yJ+won3mibgcrOfaFte7uVS4rKUToCcuqz1jL6hhRSTwd6
KMdSoVltcatFDXF+ju3+zRkhHovRgPnJdptcXAbioR8F6G09KPb1zY6adjJaEvZnYuuF8HiDVH85
I39WSli1uAE9oplenOaawoH+1BN/Rk/rPbI6qc1zqO+gP/3gOZCPvu3RSepd6DLCvo94BMYNKiuL
EHs6sfAkbbCHJ4C5cMBeE6UtTojhKxW9ALhtnAtkHg6ouyxT/zL/v4EJezlpTkMOYb3Wg2D1d65T
DFIPrXs6lbM07Ggk9K7MBE0yY5OTwjpj5bGDQBND6ZiGgpans2Vv1am5YUjl4fcLMYOFyfKFTmT9
qkJgcdFtFeGOCevLa7Ky5FVlbxa001UtON4qiJ1TtG+QZVhufO7LkXeS/AjsYkWhyHPz0NI5QdB7
49Wl/p4oJisX1kAkwgtO1YPGwfB7i/U78nAZSC7Fo5CsTK8kd2lc+XlHs84uDyFQyQFETx6uCdGQ
WWjHTaDhKxfJpx5+TCjFr4jAJrAxAAN2apSe6y5hUeW8FK3T9IevqRsXoGyqZzvMJyYSmsd3UV4r
YUQIOMx8NT9psV3q9w5x1TRITl1p3HsXrHYuhtLfzaE/VQNZNvkur0nOKBElRqkYMzrrnBiCE08l
CsGSQBI4wUGjUOaa1R0hWudsm11UAUTwwcaTZy3Axz3tmtVHim3SYNOpeCATy2mOpXLAeEkXdE+Z
3/zZfvs/pHO46ZlcanufGczJQ9LVsv23vDqUYk7HjxrFi3uGmQtb3h7f6Wk5qxdJDWv8oiFKz2ud
ovSjRYeOLimnp+9jJazC8jiCggYeT7HlyszQx/Hw8nTqao3sCdwWq9cpg41n+As3szE3viaDzsOS
Z5FscYPLobhxKPgddHGFYLpRqxGuoSbGFvxHURmOJeyUBUh0nGsTeid2u1E9HPasI2inP1zA2MnB
Dc8F5/OfQZvBnVqXKkDLQb+OLZ0UseyTsC/XUWb5RdDNSSPWnTB5U/FQeWD90vU9Ngkql7MupfB6
fYdSZgp3KW8q7rBvPIblCCikoCAi7bU6Tv4B/VhcbV8hRnc27TjqjnHYrg7OIatn2kxJDEWhm9gB
EI0qKg0cvK4cZtsaflnJBMgYj4cG7eAZtFNmK7ED+GN9w8LUmPOZVvcnFD99bcSrff8RXEtqB+ly
LOTep6RtIioSBwMCqIoHB4EHbeYjjkov0hqxBsAq0jgJIGYOu9izOCj6op9IdeZf+szu7gxGlOWr
FhVO7T8jaKMWVmsUIL4EdGuvbddnHxG6kM5CuuKpeJlsROIFW+psdAGA65qd/w3WNUR8rphCYZBG
fimHN1Zn0mYLycQcv2MKYo/2mHcoCvfepUrGV9QcGxbM55fO9Dlu8lbT7cOQ/lKhoigHWPXOgJWp
ysplhG+BzKvfSStYeYzQx2H4D6461ZDzbeeCuuPOOy+uDg+zL8X27dsmuVzeobo491UpspbvvgW/
+wF6graMeiQ3teNJCa8d9SWZ+/3g3Uh+1XPcriSmoZPMB8lAiXj7wqsoEMH1Iw9pxBusuSiEguut
pa82EgWtHx7IxLKcE5R32ir0zFLMnwBFmvqhndlg6BoUnO7lSh9HmGI4RwFOOAGhFjSLbTzgi6ic
Ln5DT+vp7annYg8eUkzvnFbY+HZ+1n8KMtQBaJ0JClTmjOeQymnMDybJN0APJtEqFg2L/lq4SM/h
4gnAGuwOUtzZmPytvVqy2UU5er0v7njBsKPNkkSj3pYOmqBv+eUOH4w0gThEx6KXutP6UvLVWeRc
U2VCTX8esuxTy9WQd1W/GZ00KCoKaW7AhTjgclVM0CvRyvFi5fdyPuClzHl2+nZP5spyt9CAjXo1
SEmRnOKZMdpDZymibLw3LjiggmXUylOqa/Su2Tr44j4iPQ3Nnj8FRlxJWq0+1+1qpBSs0UsbrPkr
Im2K5jPW1OmTdA8xhR5qpvlAjakTPi7r7hIlXVkzkMHLeWSxeusG6dozZnn3YtNdKr86120xlD7J
ZYbn+XKh1Se1MCnlO1AeezseayXXZ18n0Lotm9nXes1WMj8NN6vOdSeaaCcdDYG0am6B1VtsvAh7
N/n8xJIB+TcNkgCX0togvUi0JBDq4b/SGIPYhT3ODYP1tMRoqI+aQaS/dUIAgEGZipObEJT1k+2y
2NvU+DT1yQ1PGn32BJTMwIZAvERlztzN4ShacHTL16fDS0Gwnc5sXGWZvb84v3bmVnUC95/CgC7A
m1qunNYSWTQO0NeEREEcInXGAcP7GCIe2IgjAROJ+xDhOTXJW579/eU5hGBr1zchD6nCcUE86Jo8
eaGfmLYuDyyKxRpcZXgcEkKWAnYAupT03hTe4nbHRs+VQfs3AP84yoABP/JdPOuRongqnYDs2oq7
MZRihiprDv+PcaXJa58H/4GqxUOO/yqX/tsIJ36zd1PrHrCiB0wj1GDkNt78CelcSgaKk6ndIglJ
g0oW7f8FGRCwjUthXl4p1vAek8piaQcqJI2ibdCPzOqhkLZlGhAtlEdjhG82pngRqBGFs+leC1uk
psWwL3h5ro88kRsQxCHOqipJ5tE4tH/EdzW3ue0JDsFK86hd7SLFyGOXau37YoSgDQbdxlj195fd
2sI/gJ89aIrcy5Y5AGbs5To2AzTkzFfHrClKY9fXRU4h0H78MiUOvmzTd0N6pNbRtq/OOUkBN+eg
B4XPc4nQUbDOKmTSiu7c3kYnurK6Hqn3A/9eq+osf2o6QB7kuyX0zPa9wSV+K0SK5WNw8fU+kwvS
9FylpHsy1p1LSrJSOGXggIWoRc45jrL4d+z/qrI0NxaPwDw0ZLx9rIT493VKGeTR8XA9Fs5OVfFl
z4xuADJS1TeStq+XmMbGN/K8OqQeyeBxEsQrGiwsH5z2d4czEN51+HGS2V6/ZZimVVKMrouDvISA
/1Zg95YsXTlb4l6483ZV5R+E9RHf9D+KVWDn7fv5zRmtnE+G1RmyUFopbI+Q0PepAJCuDutUufSq
NVMIiBLbhLM/Jv6Tgg6iIxcH9WePMIOWiHMcXQytLijxy0zNL3e+Y7nE7p+dfNQSuoyS1llVUyGe
1jX2fXhmP1i9Q1cuyjdRj86UO1O2cqqFnZgRqs5WMxZ7GfjCepclzEftd1cyLL2asLENgVDy1e3t
qwyljHpu94RI2kyjRv0kCjK2z41j0kNODVx9o4Qmli+IC3UxmQ3cnvsqdRS36T536V5ClDxPmzl0
4BnWaTRpcYjpGsqhYYCx7//M4exify0gFqDsOJWF/aMHNpbmm17jQ4/5bMY/YjnNzYol7NI0B7LL
0KDF9zbGc5xsEwfFQdu0UVXrHjY65p3UxMNdjnDfBemJEnE76glN1bGehgnGQS6R87IhLWBoPRaL
jdvCdU7MwzifCpBHa1zWQh0bVrwPL6e0vC4CQFckyMZXaPtew9SP5Q4i+h58b3Rhl3ZXEFAR67PD
kVVac8nhPPjGv2/NWp08r8KUWW7BM1OIlPXQrbmdo0EbkNxzFfIiozo4VU+wNp0moMNhy2f+MGhs
Lwr7TXLbdMAUFBlo7bbWkT672tzS5D/y3b5uEpv/CXMOmfYybHFmTQQ5IVtDchYZ91La4zKTwF2/
De59e/RObUDYsxLqCappABvi6/Oq1RLs+STNpx4vFeWEgg/0TER1eOob7kcqjgtMyKry1lgsA6nH
m0v0Kl88LABmx5gbrYJe+nuAN6qhFXQ/7PT6V7cblhyQYeYlsyuWmLm4Xt2ZpjdBYqA2FAzyrZD+
qD4Rkj5RIzmVKf4sahqi0LLpnVdSArPunAq0xonWtpwyLWPFBWIw3msxEvJlf/2iKceDzQs7w1wk
RxNxKwVuVBYT401U3FgC78VHM01KgkQOeLey1sTwGAbJsFu4UNr439h22qhl/jHsGvoT58O2QX3j
lL0ETudHaWJjL6G6uXYKnrq6H8OCmCHtElNX/n7HO7Qelf0p1k25ExgVtgpL22ALS1DeET3mW07L
RgT/J7VKr90wE5HlU4fHGR3+STvKc0BBXfS2XBBuQPSOv2RNVutqXY3ojPo38xNdaatthCFsEODv
bkUuP8OAqmcLAW/nU38pwELdukp72dDk9NfhNOogxIEAhIxOzKvGNhBGL/EXBPD9bnAL48M2Jgpn
9od5bon074mbTrN+HPk9y/7u9SHVZYLmDNYT9/9VkXwc0dWntawuR0ePfzkavLvNyPraHBlkdnc9
gNa9KKnB3Vrz/uWqqlmuMvLn2Z3oSIpA/6PRlLs1mzD/NlcC7GZpB48FvRacDcAwCkFjkq8Ae251
veko//WZr5CuEbWyv0xq9fuWOTRCr3eiEwS5alMnWB4Ck06/6zLcOOCwXLnkGAY2JOIl5kvp9x0g
RwvScz4FVC9Kt2RgYUZ/mVXtuLeNlILjelezxvthC0O/cg5c1k1LnQQOSLOAyoaFgl+KdG1TgF6U
oD/Z5TFog3pMj+QtnQWL7fWNMCLdVCyYnVeg32sU7fJbZkRz9Nkc2pFqABlCCO35KsdQT3FstL5Q
QxAM+u4V/wUwZNvlRK66RSDjn+aurN8CR+VcymdjJ0vN6pf+nYt3UApDroQDw6sTIzyCYH/+G2Qr
07lfgPXuqDnRlETTi6GNXH7q5aMA2YNq9wn/l3cR0YqzcP4F31yIrt2kmgGw4M+iTKhl/Hp2mTO4
I5bZaJlFmRGXPymJDlcr70DiPmYToZsv6p7mj3q5zRElKG5z7VGhgFhRYBHSDMJOQbTe4rfaneoN
WHER6e1Eg+DbM22xmM5p6jwGyAIs5nmxZmaMxiStk+JAFIKStil4SPP0HeREE5XCurOvETRggSM0
gmUqMn0qlvbalJpvtpR5IUgTIUcboA5hNMZYQofDKqWVNkWaheelzReqQdvSjFJfTv9S3HUWu2ZC
Ruvcy9+FWT5dFNgBWi11HChuintYzEnO6cArQMmN3S2ZIzBwNCcepAQW3Do8L01hmy1cqnjH5APx
fpad9OklZEsaMlWRopTL7AiGaslo9CnoQJBWpeYb7wWVwsOO2sVmQz4jHzueYXze6TNZhz7oBwEj
dxMPdYKU6ZNdN8zwfYEQE2jSVK31GBh1EdoO1rivVu0WZm/ndSs+1Ht/RSccLy5mVc5bM/+b2kWs
uSNMDymBm9jG1jthJyF05a2xoT4vGPntVBlEpZf+oV+a03jpnRbhjWHT5EfApsbKdQ7HSPZqdICa
2VTEpq++l9W2OI0GarXhYZ7ZLkaQ7SOF+ZFC+Rc/1PEaL/0G/+QLO6V0nPV+oBXg5PaqK8Y0VTuy
ERMB1759eKZYLUvRxvLgIsQArjpvJ4UURqP5HQ2FlktGFfsSZyCASaHLSnqr99qiDgNBsmJBCWJ5
DH+A5DgEg0rjyB4r3KcZQfNbPEnUkxgmz0YMFv4MLpROZcPfXWi8XZLzD9U6aJoFS19s/PDzikeX
wUHKyeqZMg2DsCGDvimKy/Rk0Xv4kHIulpAuHzYzMs/As0Ztr2XA1Op5WnxhyXnQ++Mz2HpN6k2r
msVtu7jHtpbPJ2IegkcDjqgpFqg0EH3vxXU61RgumzBtkQB/GAQ6IPDB5fDQGD4kwRzA0470MK3R
PxdHEAqJ0gnwL4yDe2SeCbUVHA5plF7EeeCQOK3APHRkd+h/6ta6awEjVcVZJ8P3w3Uwl0RnLI00
rXAk1+rZxAiUiVFmbb+OJmk31iMYbbUlXRkqzPbFavDInr68S4PTq2qJuezNt4L/aBM/rcK9Yf3P
sQ5FBbLUzVI3GpGODED6Jd217qo/ng4x7UEZNycCt0oxFzYQeAXdSCKCtIDhDt2ZZZOuwwCGsGCz
7JSA5BfTK8xWHwtTW89H8g7NyMUdR7L6r2wPN7K7BjsA5W5fB56x6oJC6/fJ4DWD2WeiazDmP/dZ
NSRbmsTe4lhXVEjG3bNkTZ5+XLBASJ3SB1xNi69tUQSNiGT8oBT37fN9u7rYPvLXwfNPwHCppyqz
CBoiXhdIc3p0YXj8Za+aPq3EhR3y/+MPhOW5ropU98e+GtwOGbD3Ht6KRbmW/DothE3hWBfoJseP
qVwal0qkV85Odi141PWZPlfdBjNGpTcTL0rWi0+gPxvyMth56rfyblbR3JF1N+kPIA3As9UzDDOg
cxDZr/U6ohCPsjD9Qei7zz4VdGJFZDQf+f+A2CwOUTVD2NgJ35Eet8pFxPKLKPGjwNKBhhw1GyJw
uggin9dWV8WWHc/AVCs9CjMof2BbXKfvBu/GZXvtYbtgHRP648gYeOoIH15MA3RQ+5sQfKoKBkMw
Tuwf4QNjTYqujCmJk0iUqrpaOL2Bw+4aJhcx9Uj+oRAVju49AOQrmNYJo2gf3exA14s/lRFy02dL
UBA3/0Dko9WbES21NQ1ZnnfDACO+47sku3NblYvMnaNwm7wxWOv8PsiNnEGBOzQcGKd1qp+OP5pd
V+s12hCoeeMt9aX6nSd8IJEYknR9e7qMVeQ4t+9tLFMfnzWDkjeTQVnMGDCnU6wAuhl6IpQCt9z5
604aQKUcZoBUBDRXfGbvegupwMvHPCApAgqKspHuH8pVHIec24gMR8kIUF3oAAKEEn3WzTnRVvVM
v6Jum6/5kq6qUwDqE2uJA9Xe3ZwSYao5Ke4AhHcgIE6Iweh1NC4KgDkEvN8gtAdI0mCWWzX1yoE0
3hYXrW3iAhc0srhMhrejTGEeWVQyjvoqDKuJcihxeGkoQrBnepkBqFriNDfeA29Hz+B72DkcGtXC
sdu0FvuvwVwFKazo7F6IRyw54bQbblj31VKs7z0W6x7aAC6+9ETZqu01L+PTatQnEDE6tXhFSM3X
GkVeA989HNzJLsdWDaBW0ZWd1XlcUG1KcO/4nwdGkyHWoN7hWbmGVH86DCWM0CYD8JH8BGbfrjt6
9/bbhoSeVq5avmjsD9T8tbFI/3gSXobtSVQq0LuWYGtEkPEl6wG2xLB3iXg7nCqW60rxe8bKtulO
c/r5HXAuoEnleS6GtOGVcfYMvgzxuVA5HfUH/0FanAhzYPMEcEVx/hyFWOVPo1i1lXLCF8gx70Jh
AsRh/EJpwkzgRRDfuJbaekS7kWz0ggAmmqTyarB95ruyh3RfRGmYXq52tlax51WIKg1dNt805Ntl
twEdHgNNaLwcIXKSq/fMTkcgqdM8hYkgO95Uo6BnN0Q+DUEq9cgDqZS5cTfuLZPRN4ZGUryHnSFh
EViJYJdjuXl7mSUzM/mzL4KQK5oZgdzcYD5GFTQNtZzPDhC0ZYENRgXmlxsK8Ffi7fEMmoSddrUI
67bmH0hLa/9PLwyKoaVyuvOzr1f8vgtYW9DGHGLPEiQQbtYJd60eYY3uwwJ3WTSmjZnBDc8mbOcc
4PJgIyNjXXXsl9AqztkuRro7v+s2En6+qXFBqEftWpQcPHkhyADB/obA4emDO7V99jFbfCqqLXM4
QPdFLo/12uTPWlocA7os+sJ8VS9CfyXGJsBPaPxIIs9v97B71FvDLnaFxm+LvVi7nSyFaCV+UbDD
TubZMAHEhfGwmqgZeplMYkf05x9cQRZUDfeYA/K71/u48fmGywP4p5BHH6SXn6JznUU1aOFSE1+y
UXqE0NaUxA5NsVCzDYxCm0NM1wIL5cRAIkdGzPXJy8chNmQzI7eoI4Z2oADH3VSP5RE6ojhyeXgA
O0luJb6wv5Jau1/ZB63/9LlvOZET1U9ah9qMy7GTO7GV4mvSOrv0bef6dpfJRO/0tUIs5TZuYL4z
kLdrRobPYw9l5K0WbXPlRvsv4NRgKrT2f6CrwenY+bY5xTMz48yDnpCJFclEomTn73arCZbkgpKs
cVbgsIpTO0rui5LO68yFxFc+O/dHu8UH8JjwJJN+/HcUhVKfu2LHBHM7EBCLwjX87PJwCdKkW4V7
gQr6WOlq0I4PY/lVDaz/NBe9K/WzqvzJTfH3GiUX/ilU7dEKywgd5KDxo4CJKlyAf71OYSkwP+Oj
SgZmypN4OMZQwmY6WLaDHONTWkNG8M7YWzbVp9DVmT/FjJzfQYUiAnNpnZ+J6lAoiJ1s2AC+kI6g
hXqYBwRgy5I8olPSwA1n2pgLcX5zWDeDOsgRrFRbmI1mmtOYXpaoTgfZLfXd3HpOqFeFjKwzN5R7
nfhM+r6Iy5sqI05hmq+nm5SH9Hi2iNYVqUVd2AlQp5SwHeWvFYux8VrZTzeQDxDQxvRJ7hOcSnuH
cDJ80o2lW0pwWeZFxYAUYyRjKJdP0nY57kpyyRGiMZZCdsQ4cv9k2ni7Mr8FuVc5C1gizGTRTc75
h48SDLxBodaFeLxckPx0JIamX/Y38iyQYrP6mHT65dktxlmXUxlngxk0t3qCv6sMCOgSfOlYmKs2
CASuiafXF02JRqrMFKwLkKPEjR3AP0TppRUTa/HVDrGGRCmh3/Ic+UMm9x0vGKlU/Qh8+QOeb679
Aum8ASZxkCW4MZRpefidPAujXuGpNa8wUPYsxke+5EwiaZEvrYOTVmf8k8wrgASKj8TQFYXpVuBe
RwL290JiotcFz9Pl1m0DNWqcoCgGdiwu9HKcGAqsEG6DykT6s4RSbpa4/s/8e5rsm+vLjoP1nqhs
osrgGOuietkTDtBWSkLprCjqDpSXxR2sfDLuuThFqkCcXujL+AbjZiFXnMwGI0rcBhQ53dgpy6ll
GxIEUivgFuYnWRV8VM6hfMutnYRfQSP0GWLrUqeguP+3YnGzuyd+wKZRYRHUmuGbzcNA/Q19La5b
nEs87uKEJD6GaJBgK9p0PtcLqF6nusp2JYKDKSi8yI7MvW0X06XlRTWWJzG6oRtLG4vgX7BikkJO
jMv9TU2+o0dKy/7h8TJRhOJ/EmDCiundMuPGYmX7q4KJDKawibaM2Hfoa7PEo1imd1VxJNOBzk17
LKUTZ8ODq6fFZFMYKRLsw4V8ieWnD1A7iOZHvgcfYk134RPmLOK/k1CLkYyLeexTgdWOhCgvs4tL
SUXUdNOAmOUaN+BSKSaI3/95FCViMLhcS6/uuKaFGf/zJkLFfP+ln6NqNBjnAp6UrjZo7uD2VvQe
QZ3DS0PvFaPhTDhhYkOhGlbEtnaz/SRDp9sOgP6eS2PdczpGO6WOR5iZmBku3uwkxzZGMKc8wwWi
5zUbbWllwXpTZPswh8+x5uAhsgTCAfalFE/GgYO7GVDrGd5WfZsencuS3XxuZo64QYsUfCqgXjUL
XLZhZT/v6QCiycgFt8QN1Z5cPtSzkJQkZ4Rb7pTOOeKDtL1ufEM2QUpoWgV1MwBW+NChdeoZVwvf
tUowD/Bcxn2pdj0pjP0xD9llMNcvwqgOhlsRo8f23HWgsruHLrimP2m486hzAvgcvx31syLvW6HZ
BM0x1WWjzZXb67IPTp6BX5E3weiELINvxbXhUAZP7hdy7jM/zIrkQ3aykowQGUVFKO4eho4AvbSS
AsNWOXnNo0xQ5D20eRNkkFh31Ej0wRv5gOQCGrS36BLEgtuTTNV0kO/E/ZC3LKoHdayFOk+EgcEU
+LPx2qEXS5Ei1ObTBXqv/0v0zNHgKyvzz7rEF1qDSTHO3eKczvLd4+kqI/SeQmKFlXzQbCg7i1AT
EI6W4r3XBsKiXpcKVu4XZLOfBUi4rnVhe0VfEWE6ihJfp+RVaaaEK5HmEcl3C8kf2heU+TMSHoBC
8G/ym+fEmAuVUYS0PHOgG+PebTiWg6JNAUscFsUl8QEzQMo5lWP1kpeewBXe80Gxk4VIbJ7YCW9B
ZnwfaeJOEZX3daJ14h3n3a+0wqz7mTk0TMtmW92jQ8uV8IBGf9CzpOKcRzHj89YrPhVUxTkJvHeL
FWGBobSPHps6k3qRHLq8ekiQZ5iZYij2ww5bmzc2G9euW2kT/kuYYtp5CGxSEe5C+iDzrxHF7L58
27k2gcBtqK5eCeW8lnwOQGsB49+O7AqN6jwpzS54ANEGqmRofwP242D5CWhwSKtdtgaGn6sOpWb3
NAcehCDBvt3DshJi4wI/+xvW5ScGkWthqRDfGdCPUJX8vvzg3y1BIla99iyOMGK6uOtu9TKFS0UI
CEvsJhnRHOP3rDK+j3Fau28YWrVRIgb9IVTVsQAw3xlPsqUUnxaWVCQB5UsfvLGUAFVOIh+B7nnj
TIlsIFM4EDWalST2IapkXg06dYvSi75wmPQ3eTIGIyGBx+ZGFDM21PAk9LKeACWucUOTgPhxjNhH
b8wXN12FXKpod+xtTJ67nBElgTpVU3fU+ugjXDKsb4hU48nCnj3pFeb81ADH5lVWUl+A2WRdNBk1
5kXs2kyv5EFJ3JipEkvjFW43q+bOw603l3QXRHhMtPDvp0WkLM5Toxkrw/zOeMNMUskLsSkgsEpL
oqyD//9wNLuOXOsSct+a/WWjoZSB3qhWNEBPGyrw0UgKntekpb6voky8mDLNEU+MYQLQ27K8ppJs
ekIvkdGWOFmzxb7CrnodrUb4n7K8SW/MEmCFmdhtU9q90DirnsSkv0JoCikVi20GuNyDuSDIXItl
JqJJoMW+ea1mG4QCIyLGZ0W46pZuE0kDE9HJRjV3X5pW7nMBKjHfHKEhVBW+jFOiGKwo/sg2T4Yf
MYrV0RymN9H5oGZ7WGm3u4WGF495N860DdchGv5nXHx3Ok5WO7x1C96AABso//k/g9dP/cyWYG87
P3+WB49S0+7CRy/pZY7/Syc8e46aE+4hX02dkX0lIm3JS0af2RZSce2TnFUfmLpQMVr2MX/WO8me
1y8sVqKOwO/Kz0zEzPvIz9ujAx0ap7eVv+0msXmuPN7UoKI4zqXDUdPuO0wbTFWsdASn81DwLwqh
Z+GZBJYVUa8eI9VhUH33/A8SINgdb+MOAyEdaonqPDaEVl6yVxtYC3VCAd+8lZ2Uw7xMMtV32Xrs
DcOwNCZE2cEhcaEtBzJNCJwNxGbOoncrEjx7tAPH1cMBWWIU43UwMfLlfQ4pt73Ht9xFxG/NuRkb
KamcQ3DR7mB7j4t06P5zLmzC44rEhgSiVtFc+SpEY/LJ5DZWxdqEoCfxGktLvIrL1PRc++cm7PyJ
NXpk79HkWOfV/5xSxQH5Au1nlvGkic8ScCPMMtk9PUdqFlcL81eG55lazQSnJFbYFTfxBuib2VZa
gWulOnefLXbyGML26hnOh4YG2p/G1Ohk2xjXiuG7W7arbV9fUPnKHXjIA9TMhESl9LXohTY99lu8
BV1w2U0VsaP0K8JuKyR4NMuLjC3OJ/ftTu+PhbgrGL0xGWRExA3Yj2z9PcBeR903qOuWwD6GtDUa
OGDE9auLITT4iIbQRPz5VYPBwrJ+E6+oZYzBVV9bOnGvbDVUOkI/Z/Yil9hxpT5v84CVzpDF1HG/
7gWCeRQnsUwQuvZBIJWypVTGaO2sJncRAgSeNP2+zIdIkozfSlAKDF8Y84HlO619eXMc3Z+E5koO
+mQT02cAW1wzEYX1aLuBTHsEvUEusF8obzLkgCz9ozr0iPXhwiEh8feEo79Y6IUfZHWrOgZxshUj
6nbDM39fhfcROKqW8/1l0PlxBHv77nHTXXF4uieRLb/g96M+dQe6rj/60of70lTe9+1awtG/Pnii
JIvsiwfewLpIwicGvZHx+M/EIz6GR0Lq8R6OvI+go7Jm0GKtnQugg0QwdEF/3Ideroj42/qFmaEt
7R52aVG5JPfDrc0hC0SqDee9jzXJUl999czIy//BrpqJzHEkU7S8M/MD034yOpZfn3rSmwJjRmBh
ogYtfHjddZDlOOGw1s5z8Ferw2CsebbWYp5hRhCR5lhTJ15N+Na/ihA4rpLJE9aEif5dBj3/JNyR
Dc3JisK2fM7oHv7iXJ4coqkrdSqGmn+/IM7QICH4yvv6XJ2BlK5FX3vFl36K6qkEpGoFvr+r1c3l
A4eUXotvjwAzHfo6G3mYuNBb65DlvvVK8DoJLg037/r776b47/e5z/cX6+pb8au739v6Pto3ffq/
La1LFNINa1xXmj0lWdgShInniZnx+BZwNaU4KnuI1HGgJQ15QOka3XMUl0iLfWbykNDRrxg+S4Jz
1x+iLcZG53P+zSZ10tN81UNGh/T3O2s8krlDqmvnyvcARhTQ8Xqyqw7OjG4Lb9bqBRAvlGgWNkRh
9RvWRHcDk1weQHLt/ch7qvtQqoa9gDTKTl3nJgjlIgg7u9Y94W4v9CLrnPRyyoGJjoyPPtZauA1k
2zjIY5pv2fBCb4B7Nw73W0ZlwLwJgewQgRZGkgOlJSCLir9zJnrMrrbKG5x/5eO5up/pRAYIh6Ab
qLnIyK0Gx2oFn0Hce5864lbmrxkd/UM1CxfKU+qGAt74v7fHwpbAdGyVf287TGnixThy8D9cTXCs
tKUQOotIR8VpLkArA7oMnYMDlW2tXiG3GSzLPlf5jeCYIOilq9lgiOnJMGXwWZRlGil49Ywz8tGI
yoTW0eSpyBk6ivJkYWEwTEMxDqXJwQ8F8SbZ+8v+CwFrySoidq/zD5FsRVupVcNIO19mCLYDYIM7
BX8RISZ96fIYTNXVf1uR1EwZKaOd0Ih7/tsnXxxVHEKKemKGY1WkCcdT8DqQSdfT2Rh+wlUB2g7M
uvWf0/K/n/fuwhA5jQSKSEINKftuPxAZZ1U4euQs+BMNcxaod1budpKR0RZmms9NeQjMN3xyzM8s
tbm+I+f3J/nndNkQRuMnxY5PfDJdCkNHz/t/tXZVlJtfAg0csbLBPAM+G/yzoMEonbKUSEF/sGe5
ftEZXXMZ7G+txawLTL1sRW3EXlca3O4IXmhsaOQ85v8JJC7eJYsuN56vGH90xrRhnS5dAdkn3pT+
UBlLpirxVpTHhSaUXrRMGwIlrqBzI51TJ5NWHLdFIYT+OmB6KqbRlghQrhUZD4bJ9CsdHogaFJY1
PCNVpz2RaORR2Uukj6sbkpELc6gn+tmaXhNq/jTw5VeW3lREF4X1ySrgDnbNNldOMflxzgNy98Kg
BudoS5qn7lC8GREY+dPGp/Q5sRuP/GFpvmtfm+kHOwDiPJ/THIZdN9ROZxkyu0xqO2uKiqLUrsYD
MMaNe1ncfD266VLOs5p+PkJw6q418qIdKMIPkP7uiP3aKCR3WxKnPCy0wYVYdF13sxLaBgMSRRhL
3AIP/N2szmX3mzLM5QGW3vjTPt2uT5lPeAKfJhU8RKIbnqpv5nTMDsKLDdobiNLrOGlMB/uxqdST
/UTmQKiEt6UgF5FFrZPZ2FsfyzQwDsmyptxmUs66KPi/nGIpBeAhbLbw9U5oXXm434DEWwcMswFw
7Xh1x+tApkBPk7J6EWE40URy3psHtF++KLu2G6ibWBkq6XV2xiwopOwgzLT6mRx61wDWaB5tuApx
BhLyHZnoUDwBdEam9CJPQHu2j6mHf+ZWk2MTwlq4AJgAfL06Ys/61HO3DgWtzKe82n2GaNDye2Tw
0lqxZPYGqiKpR6v8MwITRutYp8hiIxvPMNv2mHW7FBePfhGor5H5+o9QEZdVLbiJhQTQYY1eavBF
ubd7ZDO9/RqQQNViuBMnq3LiShyaDkzhMrxDVC+hmJVcmm8boRqgrP2RfiasZJ4CmQPEyx+ikIiv
4fbK9w0m075RPw0kMywih5pgM090mn9i4e2hi1PGaQDlOyBnU+fUbNXfoiKgR34sldYgX55YitZh
C0dKhTDeL3wJDqRWDvAkey132U2ZxAvvk55vITfcfQd6+vIU8AMiLmyX2Tq1Hz9S1v/pb9o9flId
MVNVsQcio+D7Fnj+XaFi3bKpz9umyJh9d2bMwpo9Mi/7BusvkMjdJrr9/eckpvITsAOq5LLcKXeb
3p6i8Cr0wad50yTPaSPlI7hgZossHu0dwYAY6rVxCA08TVLTm4Pjdzuk0ojYXXaHCXsvyTauAcXI
hAr86lglpG0WXTpunXiZX+tpsFewIuelJfi/eJzEIn5ZD8xyo2iQ6qsnj4dnSQEIy6wBKQTNSF9I
tL34P7g25KRQTAuFXyVT8T5e3at6NNtWe0Jly+Fy+mAv4wnDDl/ExIM/qIFgPbdQbMWoqnSu6kcc
WK2EnNRHzRsp1DGFCnKfIGZ0Xqc5/oiJNUYyRuRRBK9/g3O5r4oYtESctves6JZqkLpKfK+/KuRe
Z26nWm8aq9z1BGoQnCtDr3kYi3Np+oE0L4e4vPTjtUV6zhgELKz/zw4i+SVcrm/pgKnnGUBONgrg
7v0Ja3WIJK0QFT628Q3LFU2OnC8kGZTN2SZ9NGMg+vf2j76Tkuq7+mlsDA75qYStLYPPOy4c++2Q
SJefp62kG0JlVNgjvwY7LRvEtLvDZJtECHpIG9IeJst7CXoRdN9YZaJSuZ5FwquHaV2QU61sJVP5
C2NIVrzjzdgLyN6jpA0PSIFubXP414ScErufFJR/haTHksfqbgtWayPIA5MTJodZhvbDmcbmgLoY
/ved95nGGtAJ0LnZbep0LKZptf198ULDsnCzpb4HaGqXch0vvzu/NHz3VDL4cljHzUZ+MALokDcf
d1B7T/fkk546d0MZ2FnCWU+Y09sMVp2Orzig/pGWNFP/wHbimOGmNn0Q3gxsEM+FqhO0A+puNzHf
ZbV4lIdYy1ROXF8Ot1UT2cQRdiVymDQcDnaZIA676STtbDc4w9NBlnfrL3FuDt0y0yVkNSqmuttk
o+URDTVdDU7UhuMJ7Aq2NgU7O7zJ085Yzkne65sod3o2DQtkaJCKIYYXBnHKmrtq4sR6jtDjfQkq
5lQvT76ByNqROj11M2NiPi5I5X8RS94IrwiCQJsWRHDTT+cCbzvUghRelSpF/EOwJHosqTJ70UL1
RED47bU6t6w0Oe4dAIXCzefhUOQzTjMEjhaNNkz6k8gpRslcPTkAiPS5kFnx8NQUAOKGv5XcuMwx
fUKAiIMkRa8W71FKoKeZvrwvQe2ophYKj3FIo1Zs6K6/gD6tIFoYGDlupuzJDE8zuwwNElfOrkQ4
nSwOdpQdje/YMdgx69X/C1IFLWC6b37Ah8rjaBf2btzvP6K0kC3p0Wc7s+B92J/vYWtErXpiZSXm
9/OvZUiPnPL/9PpinMeFqZH5Ycm9ClHDLOEuQsXlvcKRsaG7usShGAYNWAj+kYWPItYyZRlyLCyf
ZtpV3NRRu/06x2TeVyc09vLlFxXevCndMmTpXhSUo1tvtzUUq3ayUuWVUpqLaX7AI4sBqm/nUTkx
GIXYV+p5Osfj8p6qB6IclZgfRr9S9V3iBOReBXiUvG4L4YjRwqh9lTebgkXWPFJupakMMKypIN+P
2muDoPMx8iO2xqc5pNdxfuWVIfgR/Z0WCqK7EYBsrcVIn1aXQm2kbK8PlnB0Fmfk0bZI92FmSMEO
pFIeaVBW0YpMxBmN0LkewTbFlGXWAycr0q9uplMHYFnjvyxTNeNpr4U2aqH6XHDILihK19KwqZO4
UkdBQRtC1JbB23tuwuZxW7IvvKySeftU29gfCucis5v8yU3NEwF8NJmnXbHQ27jBeGvtnMWUyCv6
PsDENuc/FZ6BpSuUPkszsyrQViDaS8kR53eKXQ657LCWiz65SwrSgTBX+WEWq5oKbwCuk27mRdYm
TcpUR/idO/fzv6uu2LSuXrqJw/bfD6LFklJoc9IPG8H2CU9D+ILSAtBNgupqOFIfUmCCVU1ODCDd
yWssFM7Rv4HuDzhAFNBvCanDK/xmEQt2pFu4ebIVX/lSdTT+vp3fAvZAtP/Vyke2UJVj/owSNC+L
0nZ3lvFRTT3E1r8amNQKzRsyIUbayeoeJWLRt6/Dcji73vzGB9DE4eUs/mA7wQXP8j5V/Ws6AyBc
UWsA9qRvzF8fw2ubVYFOMvxSNtoLUYEAAsVxZ2gktt87WG08rvY7BXt70GR4PfBjTfS6SVqynHgk
iPS+ksRqG8zvASbUNlWwXHGU4av/zM8j15Pmli3r7FufToDuYNyxmF1rVA/0W5oHar9nvzcDR0TG
HLpZIn5jdXhD3PKlKPSS2QWOMYeQCVzETFc6Gp1TIsd3NKtLAqmc8T1D5+8eP7UiTnm904c1jSok
69ayEiPVl3QPTys1RHTvDITWCSAtyeMTrHQIs+vClFfQLSdIxRn/MdwTdGnrwrdHoSPzLCuMih0t
Pg9hAF4pZnMhkyKn4MOn5ay46cypf9eTCJaqnaDxgJhpyY6e9RaUBPdrk7r0l53rnpBMC0CWYP5V
r1LX9teIQBIYz3ApoYEELaeLY8VgtEt/MbpmNj9hZEiXrhmQfcIBLBh6izKtCjwDDI8pS76YbuAL
cb+uIb7yX7H9nKzoe+xGLkUrbLxMZKveA19AwzAKGnBjbp/fACXxMCBc+jN4AtGSygMgBKN5FAmq
hvwgbij8I30uJcSb95MQwBL+TVtPuIwF8a6wk3w1IxiIEV2n9sW6S1qZLyTHIMLxm/9/fyAXTD9l
p0yRNxm1LDzJuE0bDDJq46cTyomTJ14i+6zJEJlib0mCBazgSQ4CgC6HUmiU8mMCNCpMYw8FRNuS
pV2wOC/ZJO4DJLbEoIolVMiz9YxcsEG6t6XpLt8CRDhOC8Yp/KUMvmcMSO1HPV7Hc9dntz4052iN
K9CTRu4YYAH1RXfv6i6cxe7rgEnt3VqFuz+vUgsb5fy47JScK2+VOsx4xYCquVN7vd1ZB0uoEuJJ
6Re4e2Q4iZq0qfmt0nuCrLghsWeNhOk1YLAJRkzTcTPfK+zXUlUY4+eQ2+pwkcSba/RCrgmcuOKO
BP10X5MBoEYFbHmiDIi5fIRfSlmKxBoT4mTWNNihg7x65VMuWWi2bfbNJkfiWVDR4JbYZGImUQCt
7UahQ1zjbKBTtiIi5y/ddA6OiD684NwbBmqMGPZADAAS+lIxyXoXphJT0Well/yCIanFdRTl+h7E
+ZD8RRfa5KTFeBNer7NyUig77KdvtCWD6UGeOYRr8x9ELBC2CVj8/Y0yTrZ+Dn8OU6buyuUhDvtW
upPc3XSv/qBosQWJwiDlg62f5QhpPLuY2kpCXqacIgjcfdnz6C4zVSEFmKjKDuHejzXP9+DsdCgC
+vg90gVYzUyQr2U6i3f4YOWb3EmbwuMpSjtHhwam3XM8i4aofKN+q6ff8HwdIwo+bHBtWVgu+40l
XHnuWLnEUrbwqxGvqqCJmNIuUeOV9MKNECcvJS0TrsGYpfyxE+4KD03Kk4UeL6NEPHbdiq7wILEe
0dM1Lryc/ZV0Qpn2FZ4n65fJyJ59iB2YbHDpzgMElM3f6/8Ol5ZhyILZvMxKgiQHvf3JCdcBT3e2
mnqg8Y2uQZLnYOMdYhHe+HObrnqYVi5T2x2aBYP0wUcZhEpb3q78XgaMfuiQ1Il0iyDZ4EC+BWEv
vAS8+1sB/hQYh2L6DV4dvUYq+M6LHKGJsM+elvmM5cYR+fuxr4u91GZcXocUHBPULCn6X3CTVniM
s4W4KbXg8mNgnB4NNEi6U/UUjsu2vCxy5ZdGUtVA3XjrgXmqMbCEmShHeZb/WHeQ9JyzZe2ENTkA
Ad4fUz8D0p66bqNFc5rbXkgLzqMNSbMezvZn6fWVJ9jf8NBy013xKhORKkTChlpedDB19t4RRx78
T3qVZprSUooy43+bcT89fLARIefTL5kUZO+zTCdDxPYVFS8FQPs1vwD+m0vKrEIBjeOPsbjzRGxB
tZPTMT7IuYBIUGWBJEeBZmbH8i3j70gSFruxZC16S7qYLsWAv7A93RE6rC059YysHEYpL/uZq3Oy
hYce1qMeQ4uEjbvOwA6jYI+r384CoMt/M1YQYBAbuHRkfHDb1NwNwNzdL/US7N5BIYcLzeBCrN1K
lcj7I/NLGUyqcdwbV6nVp/8nsxXANji8puHBTbJiDXIq5jZLBIyaNLRld6YrJgAeOYr+3kGozEPJ
U9MH+zK6mM/g1ZB3FwIMPY1SuYlCSTU5GeMjSbiFhsAkcFz08dSU4v4Q2R3JL5sI0BDPIuhhijhG
Js4hyltnwMCldwA//5n/LeESGRli0ISOnw4IPy+W9BUfRzD7gBAQ/aUI331xY7e4XJ7Nrpor+PFU
L2OScSiQvNvlquNx0BMi1rBRc4gbyjZLZyNCwTVpMW18BOdevhF35i4OoMcn7HGbWqFo165v8h9g
MEu9I5LQw0KpnMyK6oCgjJKK5jGIu1txdJxejpjC9E+3gZoZeuOV3R5X9JLCt0ziuQ6qgxZp88Om
MORKO02wBsa94XRsosuM3UfcltZQ774aj0Bxxc7+V50/CLiUkkNNmAYwZNQK/NiR+u8keKC3VSha
2nJ+JjHOR21Ys5QghJIvB2bc7TqeVhcilCIyd4zbPXr+SGcubX1Siy40js6xVWFEwiyNeP+hpO4h
rPQpb+NglkDB7b/jlD3s8hbLPKHmyIn4EuSaCp9HC/12GiYTIGhM7qLKpRGGwqfYCc09YXOfUXQx
rs8tZ0+AryGiIXTkxg1UqHlwJPl80idKqveeLy+RZV7zAiIdwBbf2CPkPL7xMz1BX2JDPcNmO4V0
k+0dJ5l7fZeAHKy1ruYCTuYRUoMQxryQNvchOEI4bKWCmFR8zljQjII0yJAlRViG1aWl8hDwdFo5
dC/qkv7fjbBfQcpBE4+m5rin8XbVfbds9xpogWa5g95Z1SRw7VEtsLCqnHKR+z3VNa9liuDvu2YL
RGaRp6n+yH3kGB2Rfquf2qgBOxNXVztex5MhE/pt55dKtG2gu4aICv2DbP7dRhM8b9C313EZU8ng
LZ05wUw/DjgiihKNu2TslG4HWlYY7Y9IUneJIqxBJP0zcS9Lqo/f9tMJktCwbJK3smPyYm2KHVng
iQJgJYnJeG3no/sbS51IDfbueQgIZZ7ZqWIiXhcxa+KQVLjJ2vIRj5AEEyQNDaPt03/mbfXtQBgK
jfGPXNgEs2jGX/Y4QmaDbO7AogUPn8kLneM1KvCQjEPNtcl6Jija3F+6sjdp9VSVbYZ3rJIFKE9h
BHyWoDIBni5702mfXGdV4AJZ8cOTmthTmEfb1oV+/XWUcCJuZqLkaPanzXZShq2KM54spuDEdhjE
3ShE+4AZDQoIq9Flk9zXF2li46bnmpsNYouj/4qYwC0dtgVdeFur3rVLE5hLTyaiDtnb4aKNUOu+
zpqwJWOcl4z+K7dbanAX+pfz0pp+cvjG4SMFIds+gPBxnrZnlUe8CYM9OKVHX6SQ3lP6I0Au40B6
4CmHFa5XrfGC+2DH4dfwMfeBN9zl6xr2lCgImdBVTOG2VPQZF5Scy4f9M9RJ2+mf5G7/brlI54jJ
EXw/PUdwmy/jYJ93ta7zznTVfiSh9A9ewT5/GKV/2AVhSaBQLfiQmNuGIkOiNQhBZvUfQLwkGSnH
xYvTxud3ImyimZUwKp1lzriY2TUrBkMPS2LGMLJyw1Fkd8t0F01bDtZs3ngbWEfEel2e71jJAERb
aHjvd1WjQC9JwZBbyuyjJwf7/XN3MNg6AU4eh3+4NCnHzED6ZB228Puyc6ufrS0bT5ohH8f6NaTi
yEakx/mcJQAlhmlvLWUURpuGfksPTU4CDeR/vl2SVU5KFwVtgM/XrNYueYr6OqeJq0Q3uxeLgQQp
A83kWGUGZOtS3YSgsuK4vcI2rMMkAzxaPd3ziK4xtywBEfDFGpAauv8DJqkn4x5+c5WASJwX+ec6
e5BHcUgwcGzatH6OdAwg7Gkz1BqJ8TgwzJkOF6YzfXcuzyqdw6dREPKW+Zvdgp7nP6FESCa1SRp+
Dp5K3x4lRmTADSIEmum2sn/LNEjc2/4tS39ScCKUJd33Oy6CwpwDH7+ImkbnyxrXQZnHojk++PK8
XR9+YER/ZIoAyOYIJgWB2NBqCW5p/iFeeJcmjvWUwgA+cV6ctrNASY5jkW7uBpHN5/Q3IVuWKyvo
XvtfFBmppBDHK39+m+cxdWv3orzwIUZefZQ/QvR7bVi1ngpXKg3FJskzb+uUf6i/l8IXbdxvnk7Y
vWAg+5ndQpgFq3anDsibZUDRGI9VcXRD4XsdjO8INNsRRMIwOgBkPJsfDYupTYC15Fzh5/zWHlKc
1Ld/qoCWRZWDJVpMSxA86wcOtEUCGbyZiqs/CQXKXh+iiY6OZ1VdZJvUt0as7+x9w7+fd7xmsfOK
SdyoqfYYv7f6R/buwilwxp1hWTG62oyXUbmEaPVWSmKpY8VdYhKkMpw+lUAuxRqIdrqilnVvFh0C
WF6r4FeRiZ2koVVRlzWfRQijOQCOHNYN7Z4Sn2uZVGuN/rEkqqF8q7CWQJx5aAs1bPgK75uZsPL4
07tBQkhJKEQeLUTQirxlx4ig9GwzSpGP20NOjtp22y3XKOG+XVUdZKtwV50WqUsm1qmiKxZNo8GF
tDJ0i48a2lfGYWUU1i4DHuV26/vEYTmlFA==
`protect end_protected

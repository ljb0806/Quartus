��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y���U� ��i;�N�|��.D\2�kx`k��j"*s������N5�`�ծ�`I
%)yT<2�����W��{*���c��wjA.��<۱�����Nci��9��nӼ�Z%����7�s`7����*ْW�퟿&^>�5�K��C+(���`���jy�ɏ���Y��E��s�t�j&��M�9jh9���7X�+M�3�h����:^\�����X�� }�od��r�@е�N-n^��#-��;*�B�k�}�3���h+��z~�̣3t�]�"%!P"��Z��%�`��%��Gb߈��S�p��I���4�����	 G�	~���Hq�L
��83�b�2�_D�J0Q0�_���?���������Z)ݩ��)x�K�R@*�XdR�������sV�|c�i�T�f� 8@�'�Ă���^�P����+H=y#�;��0�{���<�(��9���t7�^�H�!|��s�e�\sS� w�`���髕�͒����]M�6Y�O��5Q.�-3�
������޾�N�X''/\od A�GLoF��Nw�sq��1Y�/���?A ৥�
;D?�'y�����e��}�j ^��\$�j���@�޼�����>r�@.�D���[�����PY��H�I��������#�߂�T��卓EL�Nġ�t�����{J��>�W]j4g�9҃�W�j�>��ѕ#Fθ����T���}H l��d#�t<'3����n5��H����S�΢�C}*�n�\VY�����d���J���I����Q��z��=��r�+5n�ו���$ӿ�S��R����a�4HR+PU��樍�|�cf'ފ�h+�ۏ4 ͏��T�GK0���nN$"p�.�=[��î����vyb�p����hN�W�璊]r�I�X=:����v
b:��9a��O��k�:_������Ov�}�X��LT�9�
�Jb���:6�X)��,�x���$걧\#��8�.	g���n��@�����z����~��̃6����u��Ou���r�-v����s���q�Y��AO2�W/*���O���@�tK��]��C���@/U�*����sRX�S(V�U�߸��ӍsZ�s~/�M �(��[�E;';�
����:p�|�0�k@�3A�Pa��/o���hs��N��C%�mC(�B�u��������{��~��K�!�#��2�<����v^�P���+]X�2�#��U�#�]��HS�iF���d��`�W�Q�>]>���6����r{�t6Ϝ�";Q�|�V��� 떭���u���G��HS	h�XO�+@�D>�7mJu��9�|�T/X��ڕ����;���׮��Q���v��g	�@8Àb7Ʉ�	��2~�'��R0�kdu�ؖ6A�6�=��s�v1Y巐Olߐ���v�XY���MHh������ /���g�0$ԒnU�Q�{�E�HbVWw���	l1�pD��2�*nHf1�vr��n�#���7w�zyw��un*eedY�A��5���A�k�w2|���GUQp6��Q�fJ��E��*H�]6Bs	bV�o�p�����>U�:�(j*x9d˞35���X�|�=p+���9������c}��HC� ���<R����DG؇Tt�.\��Gl�l��z�Y"��)GhwL�s6=l�L?s&�V�C_L���^�!��܁��k_3�x�}�I��,x���SZ#���%�D9�g��U�_��W} �����Xe丵�]�w�ޖV��B����%������V˩[S��;�r:�2r��� ���'��e�_&�D�?-/|��I�]��'R�P���<YC� �� v�T�	>=��Yz�B\M<MQS	D��]����䢘A� �
�0F|AC�Y^�����lo���������\I3R=#h�yN��S�J://�Q�D�Y�D�ʤ�%>	R�	����8�\�V�M�o�BG�����/�N�X7ʣ��8^[���h����bآ/����h?�?�=ݣY�| GY��®Yڨ.t�g��S����N]]��y=��[l�*aMX�S,<��藰��S��gX�Lm�����D%d��	�-���:zlH8?yg&��`.�	�O��ӫ֦��#�`�ѯ�U��l�D���A�ޗ1KC�	�O7���w���i�*����N��q�u�I03�x�|k��8����b8|4³a��W?��:�HP ��n�1�1|�;S��=wnA�68E��Uc���eR��޷͍����Y쐑�g^x�AI���ݑ�`�&e�_4��ʎ1�`�p�%-\s\
:�����H����[�9YÙ��v��a�������t��o�������B�NS�f��5�12]a�֝�O�m�cL��b����U��^�K�-�� �}0�.	Ms�:��H�@��	;�X_�|2���i"W��2�-z���<����+7�BDPK��oGM��"��,��� �鼦k�ў(����B��ƿR�oW'��Yc"b�[xf�S�G�g����%sY���kt�6l��^��ɦ�"n��y\(����v�8�&��ZzH���ʂ��ht��x	����܄��`\�U�|�+7�#eˈj'� �/��)	D:LT��V���:`�V�9LWtm�l0��̕B�k���f�'Qf{v�l�Z����m����v��;s��*��˜��7�9F�z�����ޣo��Q���VX������^���MT����<�jZ.�]E�&�#���h[���Q��0D�����X��}or;�e��֯bS�}���3S]�����>�e���<�H4N���=����hzc�Q�643�0!_l_!�ix⏫�	S��8�8��
�t�+E���;*��.(*(+�1�.##;U�F9J#���ݤ�`�|/*���ڻdu.�MbʘP@ʇ���n�ܹ���a]�ﴼ�mCaW69�X���Pɉ����C=����n�h
j�Ő�2�
���`��'�Ǳz�َq7:҈6��I���)��g"Ì/I�*DT�co��o���UwF��:�!�⶷������X��끡��֟���=K#?/���\�`=��������9f���r���B����K'��U�ED5�ڰ�ɧ��X?�������{`��.��f@�J���Z����]�A�N�-�wO%�4nk*�DP�I
�,��XG�<�R8��Z?d9�8��VN���ik]%	ce!�X���,�4>m|1Pi��MV����$H:��<؊Eb���9���GD1�#{o�4wY�J�������rY�����˰�HQ��`{���.h�Ж�m��Xel�B2~d���IT�!T1>=⸕�
j.Q���	jR��྽�ڨ�鬂�����v]6$H.�J��_�պe�N��{�	ێ ܈�al=IW����q�J��㟠��l���%}c�����dRQ�P�x��d{�T׻Ug�ⷔ�d&w��$����:�q����7d��9��3D���?I��2 ��/��$����1BQ0���ڈ�[�x����It�T�1c-�1�����A�Z�:��_�j�/4�IF�A�׊�4+�\�8����'�h;Z:<J���>��ڢ�Wh(�!�=�+�VOmi����		���K\�3R���,`}��& �5�A;�? � p�� �A���^/�:���+@G}��)>��a(�D�E�S!E0��+�$jNo��V��=/�+� �{��g�b`�v�e��t'�=��Å��ϭ��{g]���v�֒�B�&;m#(#Y�Q�k3oQ�nw&�+%X�7-LH>"�)�I�[�A����S�a ��lHF���!�	,����3^qK�b�"��}k �TE�S'�G.�־'Yz*i2ú?ߛ~o	��]rAP���4��/ܽx�Y3���U��=�M9L.�˥�����ݬ�������xýyr�8� ���|9F�j�=��i����	�Ą	�Z�С+h�,u��0%@�c=f���J���{����u~ZL&�[�މ5�補[{	�u$0_��ѥ:��`g��He/Ŭ)<x��ἰ�dO���ﴄ�f�C���s���s�����-���]��; �ђ����C$��&�!qЧr_�M��%H +���H�㣪� ��Z"���Kv�L����D#߮D��la��ÁփJ(� �o
�Dow��Ur5��'�UMdM�-P\�0.����y���M�$BS�u_b;;�
�.�0WL-��D��dݢ��(׬�H��= .�,��\aX���ud�`we�a(�:�\: w; w`����'p��a�X����bg-~T�!�7G��N�����Z�s� u�<��BD��%��q}��9tՂ>��n#��j@�+������S�.)0�����6�q5Hv�4sN�{�d��ZZ �X�^��a�'����	��G3������h����gC=be���9٥?�X���U>d)�W(�9��[%���@/�����_�*߷�Hz�Ý-�4|��f���jt��!S��de���^�Z�cۃe��������IW*�$A`���aq��[(`�jd�`j��C���M����jƊ�����-k��\t�#V�Lg3�bCX��g����Rj`ϴ��20xR��	�Ԉ9��0��.F��[�)�k��ߥ�J~Ǝ�U�����C�i��&�49*զa����������"���bV�+><I��He"�y�h�� �,����g��q,���f�������0�E�q��:���Aݡz�:�w�4�d�q
t���;���}m��a�&�(X�(�)]q����_[Y��Yn�rˏ~� �t`�.{�>�l��<�c:�L8)�6��쪖9n�-&��7͚|&W���B�$;3V7m����$��R�h[_�9e����th�MY	Ub��z��S������2_��a���OH��OB���oEiUW�4С����-/��>P�)Z�S�.�4\w�w�{CFFqKK��D��뮲EK��K�����3��7Ζ��M�2����3��J0k��է�W5�>+���8�[���h]����D.A݄�@R�oD�f��y>X7�;�rFy��V�P\��_@�!��l���ԇF�:=�r""4fl�iƈ�@^�+P�T�!��{�����	�I���y�$�'���e�
���p�'A�ۇ�	(�7ȷ��kb,mq� ��3k� ��sI�<YO�*�P!Լ�ePJ���n��˔<�
�Ԗ#p׋�`.0JյG��ױ``I�ˉ��qȆ��ME%\N:���f���g�}���D$�H r�l?~���
��rS�of���!^C3V'�����o�+�9]�A;���NB�d�iᱮ�*����B{�Z�庯Mr�8� Wi�_,���D��8!��0����F�*���(�E����IT��n��Q�j��Մ���s���rٯ4i4������Ū�"���F��
���Y#���k֋"����E�+����נ&�E�������?xSͬ���SY����7ûa�y�h�1I�3쓈z�>�\����rf)!dTP�޲M��q����A�'١,�S,��h���z�Ͳ?�&r��_��BQ���-N�?q�u�]���\�4���p���g��J��!�jjI���,��U�����"i<���2�T#�"0�s��~�-�N��p�������Y��#���m86I@:��W��Zz�3�:�c�1#" �H�?�,�YD�=�I����iP��-�@�j��z}��7;�/�\_�^�DC�UkK��EAiS,��S���Y�.����Iq��?�
��:��O�J��S��������K<�=� U��8@vTt��M���G>��*�l�������?�_	����g��L����c<���$�UC�i䂎�?+8I�9_JS7Ѕ��H���p���&/,؉�o�]�j�2���|���gl�C1�/x��1���֫��U��t�Q�`l����y ��-Ä�ořp,Z�v�t1B����do���
��
��� F�5׶?2#�
1��^<��t��u\T�k>���Aԅ�����4�00�ܘ�$�X���n/%A�k��Иޑ���j�G�#r��ᓯtd:��i��o�f�S
�B�-l9X�xg.Ȝ�k�j��;�Р�J�vi���~���=�A�~x� .zaO}'��V��Xy��	ZS�o!|%���gW�g�?���kuf`m� 'h��:��T�%��U������_��3)j�� �ZS��͢��l���r3O[?��l.�[�{>���D��1��J����E�M�d
��|��rSD Ъ;&�DZ���@.����8S2�����;-���{��R���/x^��K� ��񞔓q$�f�J��:C���Yd�-��3-�����uxi�e�j!u�������_�K���*�Ml�N�ތ�ǫ�vY>A����m2�/%\^�".S�2j���r�+E�h�9&z�)֧�S����j���uIK̷@�ok+c��Z�d�0ВD��2%���@q��
̲ĕ�U"�qh�9�%H}>�N�ҩ]fհE>\p�q����7h�8Tz���B�йDʶ��1'gS%��`�5J��d��Ռ{tAWV�wf~��Gc��JgS|.��Sy���8 ;5VQ�[�����(2d�jPw8�� �@,�'uG���H���Te���:o �U��v��a��Y+!{x�t{Q4PXf=b��1���u_�pi@�#����N���pˌ^w*���#`�w��p�z&��2[x����K ίob*s��B�-��ay�'r�hA��}��$���-ɡS2͏[q>��4�����5����[�դ��*��'��c���y�%��i�rFk�+�$vޒ`�o���'�j�!'�d-�Yt��y�F����mE�2G�~ל�y��a�Ǘ���;�
�f�ڎ}]�!����w�a.��W�ZL��?vߗxn�[��5$t�uM�m5��`7���t|4�H,�e��v.�9��7��i�O/i~0z��I:BTs�<-f�y�X)I�V�3�>��8W[�S!�x�:,�|.4�$�5@�)�Kt��+�J��v��&�_yc}��@���Ֆ���P�Ä���e[��F��3�s��noLF����c��P	5��!w�����ҚI�H�̕��$�ZHh2�zn$KO�ۙŢS�ɤ)s�c-��,���r9�=���S�����] N!7��S����N�5����9����uؤ�&@~�k��mx*��m�6���y�u���#��tӟ]�AT��8y�
�")W I�*m(8^�ۦ�����a��P�;��cE"ǵ�!�
%B$S��������9q�0/�t��K
(Z�o$�yM��Q�+��W��N�bD�H�����#ɒ^-gJ�њa���C�.|'�`ICe���4�Ōg��S�)���⊟O�r!H��z���?j�����sk%���k��]+4�=6
T�J�Dk�����3p�#����V洔o]��*-h��``�����p���c�m��v������̩���zn�?�� �
�k5�?�P��bw��}슴SDyA�n��/�J���J����~H�BE�^�?d�go�U�3�STl��K���>����Ѱ� 2}_O������1`C���K��=�t(nVa��b#�F�NN_�S��\g������Z|���S~;�9�烴6���c�܏mON1%�Zõ��"
+��d��q�}5{�@�M)�a}� �uY4�D��ZƑ��EH� %$��l
�`?�cڊ��R*�F�V@>����8�281u�u�v2ߎ���T �M^�,�pE�@�7rY���oH��]d���I��f�z:��qh;�
$�GrԢ����F�&�-А�B̬��d{���S�-~[�����5/w����/���N����=y�������E�,l|:��
����(y�[��!�ɷ�1����]]j�v���OҪҭp���4�k�c۲}�uﾢ�eA�vd�ԁ�K�`9�=e�M�<�i�〷0M���׼#����YuU�
�ϳ�H7u��
@:� �{�ȀN�t�.��uS�T��rȁ�5z�<+=#oL��%�z�賹��
&k�3�P�ۭ_e0	�:4#\Z�e�zTW%i]�w<iy�\�i�y���T���cz&|S����2�_}��J�R�B!�1��&�4��G�O�A���o5I"����� ч�%���i+��lG)���ۿA���[Z�S_� �Us�?���}���G��yB�Ϧէ97q^,���~�&+�E�DX�D�S�/�Y�ƚ�!ǽ�
 I^���g��&����>;�9�9��l�����dt�)��,ܼ�5��@K�
z?��`�3��O�;�I��L#��%Z1W���J�`\b}�{L`iU�4��"v&����k��:B����WF3�ݍz�$�rOv��i%��A����K��1���1�"�kh"� Q�	��I5?V@f�C�w��^V�o�{F�׿Lu��'�m��M=�G�jo�S��!G��q��S~A�\���a�Q��PE���hk�*�ehnc����RM�Kz�A�U�	�0�qK��8�8z=y
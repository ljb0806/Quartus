-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MffnXLPHOuVM7MY2cyZ01eHtKoyN6o/V7Z+kdx1IpusbN6fgL38MedL+K81o7/lRf09Ie+TbhEro
LxxbgwPS5koo1t4A59oo2vwd82a4D5d9wnklwk/dgQAEmcw9azwSVhZno1ZrFe3TuzMWci+0bbie
rACE+CYUSSELNR8YlLkoGrUaCSpbHq3Bg7M+sAy0IUvj7mMeVVWdfOF3YEY2ALVf4IajvkHVPZ/2
5sMSY7Z2OW9XE9Tq0JHuwdwu5WrMnppZi/8Iim8k31NdEkkyRO5s6TYGWwRNT5CD7IEj0JBTpQGQ
FRraWkvItYnpIV0QUjolPpmMxP/Z1EqvGK3+QA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 194096)
`protect data_block
sYIEpYmMluupSdWs9u8wCvUPz7pL35TFuAY0Y43oVChqw48BoEKs3VJNEhq7j8I1lEzH0X3i0XY2
JfpqHLm3DXerXj6nx3twue6UqtNa+zsxR5DEcZqex0bHwmsVkLD0HePrUrva0BuKZAM0vb17DW8q
wmfxOUq9QxdclDC2WGes5qKTRK5QaLe92KH2qgZKk/uQxQ2umALnGYxkXtCiKXZJhcAYZDgkYENX
cbY7UnneVn2vASupr9HtVdeXHjjcTU9FXZZuGBrybfZR29ZeSZK+CquEchaEWHNCV1tKKuZ1b3qo
ik7kQtUY2PThi1xXdi8uFLMyckEHKUdzu8JvVXCm6MiBu4xtCmxPXX+zzIoUiUBejqfcGMtX1EUD
VD6ulcRk/MxVXTK9HI0qIKMb0kkxZnWllG73e7Q3+AAdBUXEFSNHYtHXpgAuMXTw4NysEgos77ER
mc5pAZ4J8vFiPO1dqRqtPN1s32a1mwPr/IUWvsuw/FzeYzsrwLDz/53PflTWHVVON5a69gH84+qn
shKnRi20IUCP9o2SjjO9zqWnuYl+UEIqE0QvmbQaSuOzlQ5APeLwsTlFc1Zhq0QM/Xq+m3KzwRgR
dfnHshWnECoU7wHbuOq93Aj7JOOS7IQuTMFDNKN9So8CuUbLAqfDMj6M26+urKP1SdZRJIK3+OA0
uVX8Yizm/6krj2F45PsCLRqNx9fXt09QjmYNWijXfUxkp0wEj+u/EX4MQERyHEOrcq0OcTgfEQrG
uCOGs3shxoQPFAGDx1X9KKbjrGp0CeewpXOw0/WovjrOgcm7GTrRQokutzlEzBSlEJ28DWYRv/7f
nYOiVNU0ccYCLeuhiCOvSw01AC2p4DIacFfW3wEps000izpfglq3rj0BcX6aX01ULCYZNerPP7r/
Y4gD1EAImPKYTt4kvPfo5PCoO929bgX8w/IvoHqzQqbPErBQ/eJjbdq/WHS3yXI3tZBb8x6kjvKl
GD+cOXP9jx0hPbKhi90H69UiwkbSm/+qHHHBTJwOu4Txzy6XMa8B49Xx3b6bh9bcX7qlxaf1Yrtx
nK3Tl/pszVkEp4wYm+lXl8hub99UML0HZowpoAKKkjlqyEWQ7gqUmEnb10cQqFQ3YcDThpSENtRs
+pwg9fvqA0vqz9RfWMmh8Ec03FAuF02EjR9VJqAAPG0wmWJimVOlHvm0QrgUjGIye99Rq2R3kNji
iLziX2JCgGQ6HOyy/5eTuFbpqJxORiPLeb3/iYq+2guYVC+0JEUo+kNh/w0e8X7BcnW71AGeAB+I
9lYX9RMV9oC9HZd2pGgLPYYUZcO2Ub3ddAeS5HQW1f9xefg6QcVjhhgCj/ETR+XCvRApWbOCIy+I
js59at4U8asVNCMfUXSVpKWzPIrMopU64GC5xKqJui04CW03FV4vOc8bUQVjm83V7TEIoZKUDoqR
gRCLHZLSH9V/2G9brgfyyrh8HxEyfl750z7BGLmtzXlr5v4xSzRc6EkYO5QS/gRpYMZI9WqBCigr
Iyy04Y/eubi0h9TrVJT9AYZazvogmA5VRVsg2YM9m0KXSzXjeD1Up8BC2aPC4GQpMJmcJeTfiBLQ
7/AApGRlErVDYuSmE8xWlTCJR2EgbRCN1PjRjthpzn5YdE7nmyETjkF815cgVuP+lPWjjP2YCnTu
r4yBK7sd4oA9CyMDOo9atW20WXaj6SoORxuFDyno8CrJ5qzXC5CHgc68yZldjuKbvVBWpNINV2DR
JPxIuqNk3g1hIKJT92WUfoWBk7pz8Gc8dOalMmSWi/V7Y8OduiydzF7SFW3yDSTcE5dJwdX7mLyC
/fiWlV5RHYyZPCJuafWDMH54RGQZ78l4vazc3N7P5jtxnyU9eIxJOjEO1EfJYsZDugxJYt5dVpjJ
xi2HStdQ4+nU6X1PBSzj9H8rijH+gVrpw3nihByt8cHgA8bFPKZ4lxVEg1PecBLtJFeNhX7dzCVa
2ZhRrHZUAy1Wp3Jwr55OxuZLdRGKBO1Tq+7UtMEIxdVhVdlGrki/6cI3LzVRV1i8jrGjbze4DqWk
zrTu/awFPlkmr2iUFRAf8m1TOLZvVzZr6pZe3bU10m2lNhviu/iWact2EWjjn9SChjv9wJA3PnOn
fCRiIGGUOpeGKMT0LNzSC25Y2i2wP9wnUamZq1HZbCdXFC35PZM7ZT5KPyfIU7936Neiuq5xEmA5
rAaQciahcCsD2jnbMaaA/uLv7CZ0tEAVES4L9PElM1AUm7Fg5mawPSFwRCqHEphXegcD4i69dqwr
rpIDtlHKTS1xDdSry2T6TumVSOUeP0oNINIpc9QZ70hCJb81wGhDXIcnfnHoCvtK0U4UiVwrQ2mY
x8d9UA3jkcFhb5CgMehOqckH0V4Tx1ADNp8tiKwQy8iuYnNAdLMdNQ3lx9S1chXN8D/OH5Is9rLu
h84HQkOw7BD67KAbwGGETMHeaYe9IDxpTzMMY21FMzZbNRyQAdfULEOGIHw715NSpkUFTmN0KOcp
mxWlEk0fjbrpjFr2XWGszp2I9ilujFn/9+TJn+VpDFocqHG/lCMPbnheOaAHE85IAe6L4f1NdCbX
ZpWRs+fWoLEUuRTPOMPNS27q0B2ujET0UjWeMfhWL8EIWffvCKAD4SXeQg4PqLISYNQQDUF7iTL+
67AYgRmyOUqA5bMkzz0DK+1XGyL7W+C4HGyVkCRrnuTYsALuW4Ce/3FMb5BoFzoLnqipR6UAGd8+
RymJ+/w3D4WOGhAHLhvO8mdaRH6G6KE4zZuRm1SbS7oSNXPPA20k1GXbqr9HM+VqfL3UI11oBEAz
yqbqyoU1A/+rP/CHylGF1tJuzejHgvzWn+8IKw48bM1bdUXOidH62hZKJuDfyV5Zmn+cUX4jycOg
BuMFMKec6MC/2bD8Q9cS2Vp3qm4jOBW1Dm9siEQ5kjtMLOE6M6LAVzyO9MuuUnEGve0NFGjgsFJy
InLQY/Hlm6SxBC6Bu0nezlAmv10sNQylJXFLmpKZpsJ6dnRaoC2nu2dIhn3z08MWJx0yMTDnDZm/
CCWWIluaQNs8Ix4bdMfMd9GeQkfe3oET6N3y8O1EbMQLxAvnz0UjgxmHoiAdcaWCzW0oxDICUkm5
U6uyx8Buo6B05GYH4IFO/d8Wf0cTDXqwgpMC74a+fVBfGWlrzplUAAoJelEOOH9hOUqIvSAJh8gU
LVMLgS96Dm6Ucoo49S1SgpPO3K1QOUgWZwUDkOuqnFPPlKf1w6cYOF87jVoQ5/MDltnd/WwlR78Y
ud8oDBQpF6SOepEATdZPJ6HJSAhpL4ra0pNuCfawWpGsR2/AafBpyj4zIr+gXp9uEla3vmkbzStl
oD/BEYy1+7dSJWFWW1yVQWGdwFLREaQSIoOzE9LIyo259MT5n5Gr1dfngg7EW9Hz5101a2AiUpKR
AcXu4d6S0KcYDMhE/TJJhJ6IDy/IpD4+M4PHcfjxxnqzmQScASNRiP7QSZHMmKAPTa4t7gqaGg6X
YsNeNE8LCkPfyKqcayF2mQ5gn+aS+uYLdh2Wi/7CNCXHHkONWxsYUsUbU0rkIefCUrn82nWbcTe0
o/SsC/Iv7v7FTQngJQ/y9v9Ntz7cs6AmA/stSlJCkyGQn8wFTtlxi/K4RcTvvORiL3EQaTSfDZaD
l5SzSEf5KI0h2ccs8CtDhFppOZs92JB/Urq7fjVcWByOwZ2D8BNSfLznnWHReoIVKLoHZyLHggno
gZFi0gg+QuoDgeyVr1bc28noU4+DW4sKxUmyGzKNEW7tO291N6cWDhAg4V+dsXTkhwTHfuXLCU+g
cINi7h+7UhZU2Rk5VjE6JooBnlPnoH4hmq0fTd2Ji+1AIhrNJ2vnnApFyenKL+rIbC0JGj3IvdI1
jhoQn9YYIjroUevjUJuNiT6/MDB266etaVaDnogvvWurwSziyOqGf7pzlmWJOrx1PALUVp50JO9A
tXXl+Q7YAkkCWX56I/80NAN/EMsdtgkV+FrUuxkZFFYg2ZgiBrbccO+y/pP9djz3BIYcLKlOXjqh
0xwaGk127Bunve/PKqGfHSqpFLF40xMaJ3h7qLi0Uu4q4bwHXURnclBG+iffjPEbEP6FM8g4eJmh
BmnGSgZfFbDoiXRYpVZXZmx0o2VCm0sVJ8pynMUJRMeQB9YxATvXKSx5zAkLsEvZuI6Aw4y+pt5e
VeLna1BDz7qjj0HpCPQpyc9irSiZAoH6X+c0fDIdO14Y2COGpSzcqwN9Gyv3SZ2XS8to3GItg54U
AzG6shpeATugk9NQ9Gxn76Sk2G7bNVSF1VRFZD+lC4A68MSsBOeo9KUMd6K9utdHLVsbUQhX81LL
erxaGhTic3IAiFr4YOsrexq2U5oQiFLAZ5eKi1hCHHl9KqjENRoGn/1A9e4tB6jFDYA7fTjeZIpW
bPKdZBmFikZK4XVYeZX4VhtLOdjvAxyGL2KAQ0lZJo3tmXEUYPTY0H4zNv/+FUOyHoZOq1P2c4UE
ItPeOcjAPoE7bCzgUhIKAXY9GvnOiEtIj4jYkVV/Hu3OsrLoBrinvu7Dudl3NGgEEhQOB2/vKO6a
RXMW9lzNlVoHpG7hu8Cvr1ooKr5GkdJpC7NncQRxe+4j/c264HnbhBhhV2onmtDKqv3xfFyu95pw
oEvGyPmOsgoiHyBBHqFklOn+jle1AwCjME6PhfOgiNjT+u1OLhLn7WYwV4woBo29Csueqop4fMPn
NCj2PDa0eHsviX0vRVZwcIXOJZ59Y7F72t71yrY9WJKZI1utBr3MwqpSj438FSNi84jpHHLvFsch
vqVNcXHWCVfC9SSN/H+p5kPDmenWEqoPmhx5SPKZJBXBCRl0PZE6ctwhrYac9MNfJRi52yYR5dVU
SUGVVht+CthvnjmMeXyvvojDGLTYLLwggy+zS/n990mrriO8eaFGyFBIuRP2TwLlannGcHZg4wHH
0HTvacunzABHd6aCy/XHRsqSPySzc70PhAXyiMPe8YhjnmEeCnuVu/ThqFaM6iYv0nKP8sxUPeP1
PgH4EDsGnmstJE6wKsRD6usAllhZGeafdWI8VAfWsiNo7HK6I7nnEhtm4PqBUJPaECjOTmst9jEs
pKDDK7+ZadKJjuG4btmWZgE25/+8oZEBkOHLbgXS7GcS9Mg//DB84Oy3pbUSLam9MY16FrhVCBhQ
vrNG7iMLFYW4g7WfOMsi4r62g6/zZoYV2vbXQhtrCGmKbYJdEO6T1LMNvAxtIoGS30Q3sCb91av7
QMB4pnfDs76WK8ISJwglHlwsBZYNPyngGxiFf2y7dSfall6j7iQTgfdmumK/RgD0cBDvaQmMpsGB
SrXbflE1K1eQmL38tiZafc/JmlvxlL+ZHW0sOdr5MvPoDLkWP3T737eDm7XcFzIAaWU9HzXDEyD3
AyN8z8ilYaHQT34lJM/jE/gamGaTnzP+asBSUkkUZFZK3IqhWgd5inC9nZ5Hccg+ub9c+y1Dem9z
qYAcUfMvqXBjhCR31WA7fQThizaxe1/qrSl9euqTnfNWGMrgs9Sw9iz2QpcmrFBeKosQu94XYs0A
cYZ9YVf6QWqO+NzdPi8V+ElZ0f+E6RuAYXe2hwtO2yKevKz8db9UzIFceiNaQEyBH9hZTQ9ovqOl
AXdlBpQs4fgQAPZb2mh4uL3mpSqCIVe8QdCCxlcE+CY8xqk9twt5luB3+1XqAXf+GrpotYy9NJR6
EZAEvN8ynK5faEFfSXkRUwHNQLBlSP06lW8wxlNJaoGsN5zJ+7k/lurt4XlsOC7fc9ec8V6vKSpW
kKhKDcD8OjH5j9wSx59KAHH9A7okyYxHT1WMtIxl/kNvn1Gz3JxQrz6iIxco7D1obN5YSpzoWZLs
IsmiVQFd0mhZEFQtTbWp/4CFidATKHJ+gqNUnTtJqhC5QuroU3JGa9aSFYDxJYWF2mwXOjk7rogP
4j/2xliZk3lok33mTeOqD8iAEy4RIVuMyM7ZS5bbXyX1HusUfrhI2e4ptFddcEIrQadHDwciqQ0f
clwlrRl8mzJiF9579aOSRv/9K3zQHka8q8Vjund8IUDif+Z3qQqFA7Mbvb/rFoZPtJZSmQAjjAOk
jZM0R+M5rdr7ksEeaZDKAw9uok3BAJRq4ZdKGagjcVLG/Qp8r5ic71ryPS9NaQh0J00ABKQTQyFW
Vls+ooqI7OVnY74qCZ5hLkLV1i3pkzAMP3VDvKNhLShF2EuyKg7rvkwdEDczqu91twDEKG3iFXnw
Hnro2gmzG5fQLFneG/J8adnqBUqbs9HEPF4S5MGdxLqqqqOcfnP7VGdziHFYfvgLTKyxxZJPu5WG
63jP8xLBGVI78hqQn+5Z82CdXZ+9coNeA8kFmyYyKwenFonEttEQ4Iu7xLXWjE0FbQJ+JEgcXIO2
EjGOshfiVWUM1wJo1y72BXRu7107XQzPuVwO5oohMtHDaqVlvbIn4cmSBJb8XzQDBJ13kj01oIZS
+AhUvejnSrZ0j5E5z15Xor22XUgB0ytA6rWSuZuG3GwVo3UxFA8cJIwgptxCtDm01vQFS24qWz3Z
uLEE6v7Lk/buiXI4C6025VNIaEavyJ3MzPx+fKLBMzIhMx9iGAplppZ4knl7kJVS4JtXr5XOb1Np
tc/YUSswFIwX4nCd0IOVHPJvgeL+sty+3QlwbGxEvikSWx1aLIMgn6Awwied1T6vq68SfD/xf6EM
wW/wkab2e6YCaUP1grC+WDaAx1NoMuW7icSWUswskV8pg1qqiJAOAOGXSuGzrM0GzdmifUU4Fo6F
dMGvOo7/ZYds9YNwJSw/n7bTIvQoqOg3ZEd/ncmyWFN37qTuKxo3BhlfgC8DsmBsYN9NN0bFM1e1
XiB4dQpme8QT7RayhLQNKiokPnr46Es83XZggmsvpQasyNrHqP526dfqjGvrHWFdtA1kvW+2KCJV
E0XM/Bd7hwXXVy0uMdm8KIWs45dKTbgTAP2s6Ze/zb8jRJEiIrPrY3mUqOZNogclgdEbbAVfE9jD
dFgT4nHszV92AcbXyqEhdsnT6PQerotSl9tBZBJgCS7PU6eJc+OTQtQYzVuV94zKoGbtZ4zyq5E4
rvREHMVPruPXlVGBFbnH8ss/OcQwl5xWq2V3Pagb/JKj0kvFJ2GfcOFcW31tz5CFDJvi1RtzPTRR
ZFIo7bhd1Ns4M1J/JXVpC1GHV60pKdLlSuzutmHW92xI9boxePlEJNV95jTeOL/8csKuZmgpzwZh
h7BO2KXgsH7kOcCsDwQUP40xh39ugwS4btegrNQ0q/gfuOCXYrmPu0Mblov9KKd4EN/T180O2sMt
/NrOI6vLtzg0ASFL29xJ2Ik4YGcpJaO+WbQv37ia/iFthh1bs6tTTxWkf4E8dE6uflYLDgJA2xmu
+MhT7whcKPoywoFCyGQXAbjdzKcP6QVDQRIV/xufYXo0l1Qy4FKNsTHiEQTnACbWml1FuGzYwENl
VTtEyVLNi69r1jJEhR4UhdgBvuhIeVHJ4d82gUyWTBR8vhmS8HQrmvvbyXSns2tsOTbwPws5fhHd
Hu82ZTisJxtA0ztMpov4Mz74cS6EAbowiqo8Y0axvSWvfsD8sxoabiZR8Y5/gdu3A5Kb5SOPI7RC
ksS/cNBpQM2DJMHv4WqUiBqody+4AZcnWGMTbt9GuvMVi4pN/9nE2l66CkAFIDWqQpmzE5EQKHH7
e0IjBvuUIOqijv/DwzpYh5mDAogpT8RKliPqmfH3iUOFpOpIB2NQJDGag+Ih79OE+pccnKuqodBV
67qoOE/XAFn1bAPSASmD8gPuM1GKuZ+APjXOZFS7pp3IfpbyLFF1rIj8iR8Qt20uzo3Cq+0CWh/7
KHv3wgh7OPcyEUELXsCn40iw62lvT1gCYMQK4uxgEw+xR+HWE3ob45LiUdAVZ58icklpF67G8iiO
h4RURXCMXG7hA2miDW86NTO9Q+ujvJ3h9dwdmuhAcnFt+jQ6pU2NDmadH2Je+WG2plD8PVtgWcWM
UdIvQ6nDwdC3EploQGFQMnpZCioSRPYGD0DvBKOlTNyxqqaqW7mwBNvYkBWoKkMqOZbdICSyhRUL
3JUNRmk2dt5UQrLIP/x3sOMNejggfTpTwt5+aqmnin8pgf5t1xDN9o1tafhWFOU9UkPhtEVzeHpJ
k/80r6lFiwtAJshovRsd10ARxJDAzpr60/+gK43ddpck/Qw6fODNsGfZCVHYgGAXD1gPq3TDGRVh
mmNqLt0tKsyXdWI0a/GDvRevv7G31elccfE49bMU+czS1zM9WRobR7o0eOCLKvOJGwhf524zvlzf
yE2j3/yXbzEuMsJQhdeCRwgu5JoV8Ba+xcdFxRlZEss6S9Jalct3BocrUaVIdEl1DrW+HhA3mFAN
t6GF7JoNpBdtVRwAThlF0l9f6hMKQ2pDrUGaGLJ3guM/3I8xinZdt+/Q4sKhlqe+CjtQUbaPAnGg
mfNY8NzTWyVBt17b4eTvDQYCvx88diM5erJAlWHy5lGdnLEeeDgj3iTUrNheVHq6zk4iaXkfEz6N
x19OoCrcUkg3grbEQKvtOQKR82EMLR/RgwM+MlKuZHTjW37RWv+u7wRWs27Fr+zaIsibC+55G7Mb
OfJH+D1w77iLimqO6qUX93KJWyFZOis3G3EAckNGClUlIhcLUGVkALn/qCdk53+K4M77psKChQsQ
XIa37fCfk9AJsXm7WubuIG02xZYBiyqLvJu5IsCmBvBRL/s9Q4ZKadGGEEH39j4tU8fa0ojq0ltT
td62d0m7wT2i5/++lDt0wGNjjmwnG7dM+vUUl6CfWmmyHpiBexUY7LrFATaJUqjiZUyUkRHe4NVC
Wl0MvLywNETav2ck1O90SsJVqoqeoi/4Ob69WUIQn2f04XTiXFXMqsaM6sljwlcZ0qRPHSg43LO+
qz4rp14pUAixUOkq1wZj6U8DeM2QXF6zz04lBIKs/S7Ev4NgnQdpLYQdQ9oLwU08nVBBA/2RNaq0
4hpJH3U/IGBhri/LeuHTGAeEk1FlhO7X/u9tIFnhCpdGqk3RRh2xpHuW/6RLigFR/YwojYb/jh7b
wM10c+NbqG8ISdZ2+P1ga9uqk85IkuJFD2rWCRX7ICJrvQSud0D0vYso0+BEMmXeUIoGchghSOR8
A9Vztwwe8ArnSG3Zt8exNwt8uajPPOgUwJYsAXBQYettPIfB9R6pNmuTNkcJmxEXBklX39ocm5kX
xYbKOhM3cyVHhq8cNQcd2cIRXRRaiuNCCzn7jRgfbGZ0/LFTcZhDyvDUu/MaM4ECBUZ5xIPGRcuY
U7uAspROfSqQKQQk58CBk76S7u5qZbzsvQzw/DnXW7/e4IY+M+HgCD/j54MTDthaZJFqwIMhyhHD
1eSPOrqSPsb165qpatoxvBgQZx5saxv9uX6DNWgKWrj1u179Ywr+1/t3tO3MP42YOf3YDJhye2++
YG3D+x4JQpkkIhHaTgpjqIHh/Li4ABrnJL1OlX+iAyKIJy5iT0O2V16PlG+c8qlSgRFp8eg02Mb3
26sKbtA32wZs5oYp3BNaOTPUtYFdyZZWoAJYIqfPzEvTtv0YmpQPmWCBSti4WwrEO+fs3KFwJdmw
RHzwU1F7rqYNN1I3wKX8tYw0n1A0dIx8AQf176kpI1VbUaG95N4M99sJcVQ/AH/lJgDY2Ho1mAyc
b9vRTto/TMl4xNeBJ/laIbVQO0TAMWIkcGpCHwUBhY6GelwZT+OOj9kbJ55yFlvMgP0CU6/bKjTv
+6Gj+m1cUwJ+Ae9DVlWpKrT4GmFnDk9kyps95UCsPSipmIKdGN1a8DLGoZrUUZowZE5EwbFgF+xc
vN7JBjT7JtVqmpW3HbQaYJFyJl2fqNrDW9AXkfZvI2WuZUJaQlbCD4kPItCod/llSi0btEWgKhqM
y2LMI0lzJkvuTij8sNyugamVBaMI9Hz5MlYCrf59XFRVXxo/InuP6hegq7SU9pPsrMraihF+VZbP
KxZHoZI9ys/DJBaYcW63wIQnJ07ZeAme92DsX/ui826ZH6nI9mcTtf8rGaukW9Z5YT1zqFtI2Afb
Ri5hfgjiDjKKXodDN0ECR5wWrsJAe1q7QhvOHQq19hWaIVUEbE+leDOHvPzq6CD/KKY7VTs6oR/K
xcquqs+p/mSTdvyhhBMAsrkmClXM29IZOJ7hVKCO6rodWAIpOO9gmfjNAkRH8cUcmPlv6gNfKsS4
WxB6ACapFo+1NOS+c98vBNG91uqvquilTrnrBidP0kvr35Qto4h8Tk3M9tjsPm06yuy/7yQpeHJl
evpJUaejBu1WYxKkLP8LV/OQ7k5+2Dmas/Ma/+N6gLvfL/pzx91IgxlnG69f9Id80jXB3wk14bpP
4WLxwJ0KPzHkj9eecUkGwY35SK7oeR9S9b1Bt7Z8q2cFUvj0Dg1m8n+Utib83vGa2KFxOjG9QIWs
n2regIXxpWR3KBe2SsvKQXyMUTQC/dAqdUkwut3rm+Yc6RfsHK0DSxF1hrMwey/U6NGVm1zchX9H
kwOtRANSHTmRI17RCJvkLGk2pa56/f7Jc1j/tO2RXVZVKrN0/oV9vgtvtJJ9Dczr0Xg2XhN3pKV8
otpXzGOOn2S8NnlkREMz6OUApBcXnb8X29pIvSCWxiKaeW4JKxqod2nnZJojRhx/vjvsC3rhsZX5
78VUvQ2OxK1FUXR9SRG7tHfJIBqAV1ysG4chhvRykuoWYOtSDyaGD6v4zJl6eafBqUxvKGizozjB
IJblaeZ9FgvIO+iNIVhBLxDgddrDlvKktv3HOXYvGrfMTWTy7iq93yEUEW5wSyLXXuoqmPh+q9ss
iJyQcz9YlBI/Jke4fNvNn0cgZQ78rLD/JX8Sj6ltD87aIbL2ZUNFKOduBKqyjHzs5jq6fVnNUii4
wFeazc8PYpJIS3zOT+tijCVyduuPZHSU7/JBQCTXr6XqbMu8g9BVlMOBeEC7+ryh1t26dQWKfk7H
Mv8A14I7WEwdK8ZhyKF2CNCU+DyWLDTm7p8fNKpxyWmnmVa8YuEk7r/KtqHdraK73NIiDD18O1Sf
OHfZKgH0onNyHbCP4p0CpKaoxsWtgqCjUo9o+hKj44X5bSfgFBAAciyEutl6hQXbxivcOMQdg6T7
pEosMwoUaPFhLGxKCPtvtGCicKPieUzqj7Cr71zm0MAowqTfxcaonKuMe2iPLRVLX7xfXEcj4Igh
MJjsKlvhRWXkYFPTvUrN0qPe9iXOLwjL0gAncZnGBpc9Mc0CY91biwhYYS2CdkxcvhgdFln4GnhT
J67kgeduW02sJJ6HIkT11id/m+MhxHB1P+oqWj8PLY0G8uh4O8WPTcY/NxF5TmAOJUqoploFYUla
D3mxhyDRzRT0XcToAM2l/azUnDPcnPHVl+0mFDorlvnahvoUfgcCvF4UgheoLiWFcBsX3h6bVIMb
rANbHb/bKJ34VH06kNHmNVHbsUfYSAfazSx4QLOUzY6IcT2KTdIJfH9B+IbIrAMc03XgbxTsltFC
FIgOJpAtWGbeaYM1wSkz9cdVfSM8HKeyw4EITSVkd9ovp4AjLEamlI70m9uD+6fftb3pDaMztkZA
TRjceIWilrzJBoClaVPgMtKacwFUKmYHUfG3qwPjS9MbKKC3tK5r805VPXDORlurJWy8AaufDLA1
Y6F2WW5ore9QgIQetP/Pf8A4p+OhO50bh8CrHFCMU1Jcbebd3FFe0MF5+RpRsBF9f4GJv/id1P7f
yl68n3VXf/uMAV+Pg/73ghFB5FddauKs6CZm/bQnVWhuRbBRUKrezCYyKL3V2MOCuwOki/+xPRTu
/zd+QayJ1bXQeJkqvgmy1nMUi9a1zLkA+J053Jpk/3kCTBboyrw6OJQC0cFPGR73xFC4nuWe8/kQ
YN6mrAsGNP6K0IvUval0infSsPpRnBgMEQ15TKsF5LttEQz2388XpttrEx2dqDe+ooXT/bOcvig7
0dQbYopjzYYOHgNORN55Z26k99mWwwx+Bx4avAZSJ2ZgJn3IA2GoyURqTtzdYflhEkZsHl+l+7q5
mFqq+BIt09hd/MGeCqxJDXJ3tkzJViderWwKduEoy3P720FiT8U01W9ifOXON0fmY10lHYvPW0mt
VREyTVNdwpO55RexA3560EWkI4oqPHm4GCTtmtmSBTu99g6BSuDFse7sOsV2jef3S/XZ5bicYfXG
P3sYS/RZclHZDPDTGaQGlOQqogS5vkCQ3a0JOZER+QxcEb91j4pqyKFM+u0fbqcKH4fGjnyhSpsC
Q7jvPaP+de7HWVwgQi3ry2shzIRQr7Bvc6QGu78nVtKveGCDm/Zq9J+RJ2vKLLkU2JSl3HhOngOM
LIORnUQcZshUcfs2/oyDJhGZe6gw1u+TFXlU98P2N/QG9+7FzZt0J/JOMLYS3XmyrukiQa9aoGDk
PFneqp/4CyEtIfZ2bHHNFip4plkm835Bys9nqjlADXN2m9+tJiPLwRGTgJmMmkjVc2qo6t+pHNXs
0O3V+RDfF2gB9RWe6ePmoiwndxFahTHzXI/RdQJ7o1efsr71xLMByXwt5KIcpkx4lwqt7e64XE9y
OsWMJ6Vin409mfz2GgxG/UNw0FUl1zM6yFXfFeZloG77QiWWQdFDq/E0F8CZsDfNmSKsmbdnEm/n
IvCwVAYQ8i0VN2zM6OI3Y6fvzinKijYw8ZcBynRaJnrqWLUXCuGXMTOIj66f/G0lYRiwRo5exmuX
cqgkzLC0cDr8zk4YhSr2ePfE7ggeWgFudkNxvw/adWJjj6nxlrO1qcO4Z0Q3ZTvw1Bq7U1JCAAxA
roEWSqwfnaHU3JWCCsD/gfysAATWbDVOd6EwGDHupccFVRTbDujw0T5U5tV7wSyqkgnKmLFnZWR+
3sUjyGrTiFIDQeiiWFnDNm2komA7dpjAL2X7eq17FIrtRs1JoMdqrEmEfHrySdXWT9WVdMWKM6sv
HnnTXapIwpTptqLoSSYEWehf1puMkG23x05wIKyMSrGX1Zd+AHlHMpkVaDIIobStHAkWf7XksfGo
xyRCu4B/FU1LAniAtktAC2ghOChOxUzwxr7AKbueKDRnggccrpPiqR5ec7b0Gt+0BSWfmcVz3PIx
NOr4t22nHoylBCdkJbvFzxXEDf2hJKKtHiRx1A10PkqnUNBTbzK5Owkx4+s6mcexq2OFhhQKtyk2
SATIERWHntfSJ5fcc/zs4DYEUfIXMEhGoXLiQrqgDx19Zyc+Xmv6EP/wj5m8buSwMkc51zATPKVj
qO6j6sQxugRbXynQmRsFJ238BgziIna7qja+BjVPpSuDujCOxuL9NXWZBD3eWLkfmLGldx2OJbc1
rLe+zx/1K6mWE9vAExxtdzwwUa6ST0mz1oWoJVWmqAOSj8R7YGYOfMjGFh/DgaFPDTRYOm8EAaOD
wYmTWNWS846E1pt7qIMkfE+Y01+XjEpu0/3B5F/AeGw5L8dCdNvpfrhcrgLbu0Os+CHpac4c92K6
ChZwBTsDp9QpT3cg2RN7LVrA/E4yA+g1290Znv8Braq+s8wKckKM7vxMl3YM1uHkcp/kHvjc/4Hn
4fDr+FPIAZgA4ON3x0kpyy1ZzjMXi0vlttsUPUVUa07MRAvC48PZ5MYA1SouYBQA6GEEm2ws+TqY
NHgv8CGVF88e7gslQm9OtJFx6btiU0jQMxeYSo1A4XCw9FZxhZi25VtSbjw2dyk92MWmRJE+i2nW
+dbio3wzPJGyJUWo6M4p22oqCV6LMlGkMEoRyfnkmzk9HllOxKrv5IE06Qp9shT1wcvb4ScGVC8D
K2icFHaROHftDMaToByKHyyZ4GTufRlfMxKpmN/vtgUcWd7i7G1Uw4PBXq8kDbnLoCsqE1fKkefS
OCZD0A1chQukZCpsOFsW2sEiA1h0CecRiooveSqWMLsHrHcaMr5rzpztKnERYNhsBwlpK4LBPRkA
Df3iLT/EJOnBGenPLMpD+I5RC4D8QDJK2KdoaM6c99YZs9l4syRfLrRwPJJ8qG6NxXfSQF6gZGfs
jY8tQQRN+BfjkRpTiAnSNlyEjKbJPxBBkF/BCWZM/XanJxA8YgaeVmop0ZkRL4yn/wOuuJ40DbN2
j53l5l5ksU15Enl7T3IMluMdX9mKE6t0K8KrWkbIUFOWFwxNtD/VK/s2sI/i2mCyQp25fWeccGqi
OvoZGys43BAz9JU8jtom2XOVfA2CZtMBBTgjTJWHZq7tVeR1SnX7oAn6tISITcwznUIIrD5mzuKM
ElAwWF1aJ1B17u0KTnZtquX4SuHIpzJ2dRWeHhLkbbsTP5C9eJQ/PZZ/k1qK3oilCyg+m08Opvti
ENoICEO+wMGEs7FDa8gWQa8I9JRRwcBF3LdyxWN8TEUduEmPAfWyMr8NqCIUBxZocJEUBQsJKiPO
sJP03OfKr3ltiTjAsTL24fPwLNxqM9cfytoKZ9gsVPq3AhJZPGfr1p6j56BHjJmywZcGCCEQgxR7
CHCTI1BqTTcbEUp+5dJ7/C8vg5Ip0S4XD4Nxnxs6GG4aUD3Nqq0ZtwwOX07yYPRZMThlIiS0UprP
6oBZ+jeFAoYU2eUx/nzeJzibLWujquqnoK7cD4+e2CmpZJkvdZ7ZHKhPOp6AdBsc9u4TOMLSWSsQ
hBQyYTsdB3X3RICVuDLt1QfoHChuQUyti+PpLKWScd8dW8iL1y8g9ULJCIN5HTt16KiCBtDPy1vR
3W4T4n+Yup24/MwSiTiiB/L0/813HbUxCalkJ8w9rNJ8wKwET2wkEEMTEml5G/LSnEhwfpttfav/
SYlHTbmAQ1rSc7QMYdE2C55ns3hfBtI3+9ysYoOq9BF6lQ9u2szUyK2sP8ZlGFL5Kum728WwZq1A
mh4fGNao0OnRJ6tZhX0f6HrB/pnYG+Ea4/upmyhHDKWcdrTMBZm9jITtogjjyTie8YXm9j5CE7q6
aXGs2GoirNvr2jSwvqSXCV2nfix8QkJwF6dka9BfRdh82FP9KtI9R27SFaloSABpMmGnxp39Q/6v
bqVscR1sm6Ruwu5FLgF8xgIlsM6LygYNPDFMGWZHMBzOR0qiR4KFurDcMjrvOjByQUChER5kRlIe
NhRWA9QKk70+kJzygdAXNr9W4X6Y9BApTc97NR48Avzqp3c7YfFwX7OMzf9M1MAZRkSeRbTQQXlb
nCYUzQCZ+WzndSsLrCJfgFCLFaaGPA/BjlmrFdKfwdeTBaG2g3H7PF0h9i9axBD0aGTjzB1KsrPU
797+Ut7Tv9Y8fGFMIJUBQkuZwz39yp1dWhAuL8a0zDj4GRuNTMuWkFoOllmJGmq+/CoKBIOz3JBr
nGH/1+aG6cBFjIR3a2JZfQWIiDoLyNBQh1wVfXKAl7bAOJGJl9Qze2DuFYE8dbwnqtEoTq+KbXMw
UKc8D78NeQkFq8ZQQqcPAblKazlvKhkvATxFhu96XlJfqtIfiL6GMKokLaZy1LBlpeCg/gyNBZtt
j0lSva5v2au3MRLo1uiIP96RPPbwIz0ycnPqMeJJmveRyCMiEjErOrthuTTyNfJmGuUJxeU5EOGi
TreV3n0dIA5ZxXWSDqrjLdMqP+FrBcbF394D3GgVBxhvWr/C2Kj58yOLxNrYJ4sYbTH+d29LPXqN
0iL+zuYn23l0q+4uwdPwyfDtPGdotL6JydCO2ljcLviV3fY6gVp61ogA/CNgGmA22Rp5I5C8Hn71
k5mfDk7HKGFTVoTZhZNChzuULgqLBvPPQN4rs8Tb4JWWUPsdTSXsAFeMW5ks0qimiYNibPZJO012
s1omSH9ScFOfZjL+rEGo3awLPoB/k7pkMfh+2CuANAxj4nc0wGTSMNoW7lQP9rVOSYCs+eSJl2rm
O2xMF17GQYUQ0g6YFBybXzocuHaLjrgTd1fXYpXs5Znx4tfed6WYrmhODi9V9DAxLNcGz+O96aKl
2tYmrv5H8mwbjV4EeQVnJvjJZHC6C8hI1Q9MW4MRxhZFSKLCDZqVVaMzFgOGovRzUym8Fo5BF+D1
YPPXr5B5mWYm+XYqUq6iYA6/wxUsx7VsZ2aIcp8V3A5rxS/4FQdGVRGZ7b2gOQqVvZnZ2sLbUiKp
1SJWzVt1Qsh8QnNo5OCTRvB07rFuILQ5cVrfMphznROtwmj9ws4b5Pp4mvDbWAF20dz/Yx6IIfKg
AqWfTXngaCBSV+uQUJKWkcvn5PDauDARH/KFIaus3jXzD3kMj3i4QiKAYJiidl7XEQqXTh8jOUHd
XcBwSSI5OzOaVkxyXKSuumxkex6hqu3NLdQMaH3Bq6jrM1cZdy3at8aK72IwP3iAVgFUuMzy2p5i
X7ORP9lItPhh/ktrzQ9LUX3bXqgpqCImUnTYNKRlzfk1NEHr4uM2PTT+6bgKgm+Wc7fbn+SSRcX4
pcf5tL5roFHT84PZFS0LRaM6WUAwxpB9MctPLyTPznYopeE18/5hmauZqdwcEY/F2gPutREB3Yaa
e0wS3o8+SXHxxNxffGDz6ymThsaSyTO52XIU2OcJYGMe9ELD42qOLjsUvO0lPEIZpuz+Lk7T9mv9
5hRl33BuuNjcXFsqNFD1nSlBSniNM0SIodkUbvZWlxp4luDif+cJ5QaVRdMFmgyxwnYw2/H5i+Be
X878MPsMhoGg9dsddzcNCqyxP4RLZaB8NSPdWrPyo5EKLSZILX+8zLev51lGcHrIg8wq5zKZqXLI
2q+PoioFsji4pE2UtIfDGGGrYrhCZPv3qEJCS4nS91kftsxZj8oE94iamPqIhGVslmuN4kHdEctz
J+St/eufCVoUhSkTn+pJfuwYiEILIhfxM+oBBTsgol0yP/GQO0j6U0pAlvWLR7T5vRKWEvg3Y/Ic
iT2glHfmI4dAyeIoptxnYKDZnjwIT67AUacDljvPzJAgFxJg2qLvxWdzNuqLSVoMJw2kst3BMFSJ
ULw4KOhMFKtt4dPDHr1RZ2EZTiDcik1BYLFAIdxe99VZOJ8KcZRCvjY0AN7hUAtgT7ZqNPiak3ms
BMK7loHOWkIcVB6ATjf+em9vhWWhE3Y3cKakcs8Z8wry5RSOZ3Vpk3KK1Wl1Z6G8L/6wa8HT2cWX
PO9KRaG/Rdvhqo8ieQlKhCPYcGdb2o7TqXMePdG/6Az3kHN7+o18scgwQ64MdUJk/0DdN+qydrLd
tBlAzBfGpwh8mK3IIJ+wg0XZtMAWp5X8ozOx12O47hUyvWT3qap1/tlyEuQ4nylkxGuEBi+Vw3zT
kz+lLNUdt7vgCdCsZAyTeIXmMeutWQEIP/hVP+4GCsjNvPpCO66iswnC2JCZke0TX3LBL6oRTHRM
N25RS3d2MaiSncj8T8UD7R08ZFHoROmvKGta+E4xam0ehOgerudy+e0Wkex2X24idKHV24LOSULG
NeOqy2YxuY1bStXfvX9iNLLyoxd0DICelooE0+caLre1p0ldVIHX70MuUBbwwnw+mWHUvvrrP+RV
Bc14f2/c6v+PcPR0L68hKWX06GvPg/JFzugG2qcGdbQe5PzyGW6b6kXkfNRoW2FVwSL75KfEUfGd
Xdk/Xrr7LZYRJpmFBfwTRXuqlzH5tHsPP8NCHAUV0ebhmnsFPu7dKW5F2hJlJIl1FuHsSTp/Am5V
dUK4gJNes+XOlbj59Y3CVFPFfke9/KAU+AggTnytNyNT0PwJM+7cAiheIirsgbXpCpUZulr8s41S
gMBpxXA4AJtoK+vZsxPMaqGLviP80wYvEB6/OnFl/Lmrq1Yw5/zBTLQwE3htGjaeVa4WdVXTxxeE
frNAHiimjfFy56whTKZ9XxztCCb5IE7Cdj+C5Gmj2bCw3AZSxQTqSz9qXx1G2ZETKlLJ5Sa+ChDY
bTbj7mTlL4qcpwS1n6XwCKCH+rWA6BOZrYnFZpYxrU/KQhIExF04N2fQT578X9tDi7FXTll6SFUU
a599umO5uGEvcIy0JeoM8CvK9HhQJC99IUlA9FAVFCzqzRR7l7W+yWWIanOpKywBUs7bWl5nx1F6
yK2Do7sIY1JiSLHdt3/r+q5629JVww94i5XTaTsSmZ2Yykh7w9OZ5oGzgQG12iFf6OyORnDR9ZK4
p+I3aKzqvP7ay75pl5ZjW7bUgUxfZb4JNwqT+KAM9gs1swP6ZbP/Sfa86jgp4JJH6izdEW2df1ux
uCczAHJGOigZ/zOjqZm0DTsPbJNkNy/WuSuYMq27YXSa2mhUirl2+UyfqfYpAcMOAs50LHWcm/kt
vhIDcyyqhMIhWD1xwsgBUaHQxgV27N19AOM4C8wa2u0kMU6KoP3kwbrYfQ//58VgB9lHzpSeQZ+B
sfXwMTVFUEr0kOLVvHX7+Rd6tAYMTIRt3uCXfr/6CArwn8bFhDdJB4fk2kjWEj2ubYAlfLnmP9Fe
ux5O7o6OfbVxkjhs2GAPmPPE+iRQKUsvu3gvhXa/rtOl0Cf7JJC9iYN0K7hWrQBJwIjrNR4faN4B
0yUE0rYPH+eJJiXNS2qS9XbINY44eB/tFezQN7aJx5JM9aDFLLHq9GwTVSqXI0AWRAZoEClWErB3
IZ2CxzqWynfXflTFRWE1m0yPRklOs20YbJw+BP8aGbiVYuujSsT2thnLz9+v0+iZcFsA3jw7P4wB
a9hzVPIEnvrhLQUjbq1N5XVO6ALngtHrdeaSuSvGEHsHT+9rCf8B52CQ0dS7KGjISF+t6aqNOwZU
YGxYu7yxGQxomLP0za2Aiyon6H+uBG078y3teSDcLmUIasyzL3miz8gXhmN6VKuoU6zkklSEEWan
WdcFhCVqA2zl8Usu/gdCZ2fir2e4Fun5x8F0bTASP/fu9f7U/ju8vtb9085u86DIVUsEhGb+QqPM
/c4wab7j784wCDNu9B6Sr4vOzZZC9UrEontC22agk+A3mBSM+9S3NI4V6r6YF4A49IrZIdZj7Igs
zSATjajKBOOw88oXcayB+EOPLZtzAAHKlq8DpO34GvIl2Ww7CH+q7YKWqdZQccHL+Oo4qHLZDSrT
29ouUb9/Rp2SYID9ymya21O6sC7w5dxtNqAGrjuP3xrWk6P9iXH/ZT1UQ0Uwtnd5gQm7l9VQ00Py
RPF+vsQnZNazxe3bxtVxRrMlSbPL5i9RZdpqRVFTK9m1WYLoi++Kp6NI0Za3CDY+zsXxX1wIBBMF
hY7cBqLB3u7NUR2hI5OEDJ5Uy9rJLsOaq/ChE7nO7FXH/568wI+o5wD+3F1TtXe3oyVSH9uP8ZXg
o+LmK84sbNipAlAafeXgCwW0SPhXl6fMK8gajXb7YGp/rxTpJcvQiH+Q37Lx6RHKiwLhIeZs5xhF
qAapTNh29A9vXHMiVFqLm429cOxJEE6B2syPEG+m00IhMAyC0sofv9x0YVA5SmIDuFDxu7lutOdI
9gV+mh98hMhKmiOPOCFPxdItQ9kos9kKPvWl5KMJeJ3thMZcIS9R1As8Atfyr5Fa4gzSMjlGy8+5
F6PntaDvFhgjWcxH1trntbIfatwDbWQixeQ1EFTFy15Tc7oalVFANL34QMSHXItZUX7IvkrNONxv
ZLNa80WUcKsfDPG2VW0nfUWhyeZf6e0Yl4WNcCDw/NYAcyIx6ABkVKl7815Bp44G98RYgEDmon7Q
3inWcAPEsP6GvQMJc6r4XFed14iDqeE1L0srVJK8Jpf1C43UUZgTo39fpvD6LUg7Fh97cdKRLFpt
hG5WwI2yCiNEU7fj470z+X91UmbEmCGLWIXN+dD4gZ/L2YvOwYPs2taIhaRQlxGYvAF5OEfJbumg
PxZ/QIbOlTYrkF7GyLsi5pBBuzyJNoYF/4N7/bFxX9rSnWsIezVpA5vN6bLpdpdF0QgJcPYU+Y13
je63mATYBwx55LpIK6lZX6UU5fKDee6u9mwmXZ5dYhMqbYjejH/CdCnaB2PZB/5T6wwiS2j0acBm
dGLc5KItFvriNGsUT7kLsjsOOkITJHBdzZiWyhc0EuQHJiTP6kV/N+JxExwejtYZ0GvAxU6sTglw
Lxq3bv6KmSYX23YZkL5lQnNg4pun+9JhOLv/XI4Ybgf2/xbmsDWGRCe9eYluzmrFiLBXxxo2nnx2
KDxb6r/U7IaGXnk0mRN6+93fmb6dmoz74wqv2EZ2xswjVVpp4gUSyOs6euAvW+v7dEwKWWz+ViiT
xUaPNycNiS6E0GcsUXO4gTFkpooOuDHfAUgOGje0j3UsiiGwHGl7WhM5qPrNM+U19lRHWafIqv+U
FzUo6hqQ6vrvrGTkljeCvYxHx+yXA+NqQyhJdNMQSfT7NsTpCGB6R4A/k5ZO3DN6MbVCRWdYpNP5
TNSeb9l6+dfnzXS4Uc4OADlMSps4enc/43t97KrQPdJ9lJhgyFFXUDEmPWaXO+rCNffrhwd2mcMy
DwKlIy7gH0nvkeSQj30wWdGQ7TqQfmAmvoWJLE/c1CnYtQZDVJsTVSUuLP+vapzg3DvdkKeKTHcq
WjXDPjyYImE7ItnE8aL8WkN9of2Ra1/ks7mNwREzD5V8BxZbusAV2XJheTXs+0KjCx/nh/daCA+9
lMHzF/Rya6tlPTcon6J23WOhSf6AJjmiecsXUb/p0vKOvmvrBGYLuMtuOOCP1QUHxC+/guJmY5yK
NPb8jwz1BtKibtNqBTZwWK+Zf8pLhn0O4iUTw1LhCMdYTI++V5ajta8MkDMrmtECqlBCQxjQIcOx
Zepqdov0i3luhcwzt+KbObkrU433S8poX4h1RQWxStHaRjfD0ANZpj/kyX6jtSM1/m/KE17tvdDp
c0nDesrh+p94ZYHkHu1sZoylxXQlk3AmS7Ruhd3YZEAhioLYJqHXTSybRlOOLXADLlaNWtIP7H6Q
Xr5L2EWp7O8kA1JNNs325kSQDVLc8UEzIko3FHF2ubXcDutFMh08zBRGO+B8pGZOYQdH59Y0wuEj
Bzju5mqzFcqeU9OpT7Nj/FzUALSP8cDJ3t3zEvpGoohLcXNQaZNRJvehVQREeecBXQpPcArwq+6u
q/+Jn9Lxz1KTNFwbmXoWdpqa3VBb8zeRgbs2y72jPmb3MaKDJRKvUvJ0Nxj2Cg6xk32PI0eYe5YT
z+cepCjehdONivIc8FNR+xQLwSG+rLfBcTl7DrDKfGTHWN1HfFMEbJjsn2EzcU+9UswYo3TGyolx
WyWLOVrAyotmyAEPj4LqU47w5DKukX9oXYD+gMU83ovm+gPF40zWyWA8f7GcX7zBdyONxc+Ga16t
4nBzALokScWE58SgBx5tVwc5Dy4PItSHnUWg1ll9rgVjZP17iWk3UqELeEw3obQCIHMvF22EWDLr
ardjBTfDIO4w3JkRcq7QstMejzYJNvmVqLMua8p8ueOmYj/BPABoM+b4nYHbVaz7x6qb8/US/WaQ
g+Mupi5QrlKHbAp41l7hITFDi9sBpmtH2q8/0gJDQugrytpyXnh5kTNjdAXfDPLiYdoLfIKypH/L
UrDHZARQuXiZN8VxtXgmSbIYeLioyvN0LIFXhjbcb9qS3y8eoJbKwnLCHWnSJO9pH2B6NQmxFrmB
Gbaed0/xKhRAI4baWGMBj4MhdyQEJ6kaV9siOPC2svAHx7kkxXbcPRQh8A6c602VOXZdH0rDxCz9
GyIPE23I/NgArow9U6iiQpOopC9ewQ3g1vMOAIMBzsjb09/hRmOtWwXOE3HhehehdYHFbPM//iHU
dHRMbTSDB+S9Tib/2zEBQ2Nsz3Pka57ZwUARx/PzFlB66XHXinB8Rcmk0EAsHPc7nxeQlJOHliSp
t5B1P79HFCeLSQgpXCf6pjqOtvayzxPQ+bHvwJxbHJxtAYuRiF+6OxSFqbsBCQPDtQiYsicDncly
FxXuBFWKA0nGb3oLRNJVynOUgvxkGU9MCZA93idPe45GFoo5i9fBphFolWVLP5X/GEqCpwdEF4Or
oFSDrVsdceNP63244Eis+V2I7qJRB7frV1IKtGN3XgGkX2T1e2KF0h6CcTnrSw1Zix44njbCfnEM
pzLS5o/izncLRv/zF5vlZ5dNBnqGJa5xc9CU1WntBs5SJYfD1hSd6XpF0RYK8sl+uj2S7WZyiopx
1Cuixv6mRlVlFgZ25lNwWFgCdPLXbofI1cNQvcJLEBktH0fBLGDBwDmgtB+l83HliXPfWCyi4EXs
LkXIMfTCVl9XI7uRu/Jm+GatcTUopaHaYhjeopb752jmmrA2QbgohQygg9u39ucLU5eBF0I6skhB
NnM4UcdeBnmjuvJrmYHj1pNgjXkYLJi0PgPhiexpa5tRahQUwD09RaUMp8DxS7rPykXK/1aMh7O5
R6t2LlThNrWuROcSXoS9tbTr/ePlpTqOtrD2390M8OycwOZioneoLRSqdKSiAJoF7crw6iZV+7Qe
0frdbf48uuv2+WRKwgDN8ldcPU61izmgd8Vdmw2Ph7vFVJe6xLVshkQs+fySnNbA44vK5quHqf6f
efydN6/lMnZKEfK7tjKF+7h74lRymktMjxbzdYwsRe+gv8JaGI1j/+++777mU2kjNX3ymXbNkVx6
FO6HgAVYGR3/32xiNbLJBZqYacweWSaAKFtei7FJlnCHS1u3APhjkQLPcxUpKxkk13ntSpTKrUxd
l9niv9JsxX2U/132U/KBkqX53MpOHn0A0PsKKItWgQ5w3J6L0BGIKmuZW+2ChB+Z+p2DTR83/XC7
QgOK9n2T/XoepVUmMewNQIV+cCecv9uThkud+df87+d1p4xVh5zgTUZlq2FEMa9F6/W3+3Wt+X76
F+y6xQQBt9glMH55rNSpIvy6tPSPj4NFC1/Hk9sshvYaVT45caUfJe9I4v01RmODDGlLvgTgH1AI
Dt1JHUMsdKZYkKZExIsDdis4NrwiLV4ROHhYD1FK0RhmVKo5cw5VVb6k9/tGmHl6p1SDsMWRAsPP
vtd1fPP9VTbBGZOweg9bPtp2bealdm1ji6WDo6XTeqSO4eUmA26e3cgWgeoBGm91dUw91xxc9E5N
SxKK8exufwB29/G3Ec98bo52/ABG9Narks6Ouarff3cuLv3i1DMXazZog75dP0LSHe0dUCgujPtt
ASVMktkH80x03w973qsV0mMuYYSQ7O7bw5YjjASIV32FBY9lt031oTnq9s7ZMEHJpwWv3Mm4riVP
9CVWoeDb5uJ/hIfb71pUsoTPdPlFK+FKNAhAJnnlucCg2bxcS+IFY4VDtozdd6tfrazs9QXrdHTe
LvR0Cbk6LdDzLkeVasv0jS8f5pGdTt+Q/tuKWMCjBSd3w1jEbJWuZDlnCTkZHLbFWAkGhb1gPn92
GtImMtB1dstJl7/yStNLt4rd5GokLjrG+SCVUnLvN2+eHWAjHzHhrtoq7pH5+H+FGBkNCM+u9f8e
NCX4W7RO0I49yHqn33MbkP4YY4GFSeE+ABJPfPwdwrxKtlO/Yv9yXcImFZqUwoCtLs5HUROOMYcG
3lIck8khsnVovtz7R3YZJP1CVoUypTR5LKrsXGQ1ohULNx9i4UsTSj+Niwox/hNC8GsGjcf3+jA5
YR5puWFrMv6XCyfE2yeGGRTmAGSVeIdP1sYiThikcSAXZqSH1KZiU6GZ/PnrJzfKV+VEwM9uArPt
mS+/K0sQG+4iV+1xiDc8A2ikvQMIwBcybrDYMUKgStGFcVU7R+VSG7qLN0XfkSVWkT2h6bL8dot0
L/vK5UFhRDkv+BC5o+4/rDaib32KiVStLDU5VgyTSEkgdCR8+n7NeXb7SYw7e5GyJBaEW+8edTd6
rkN7yFOUoplfQuDHHDUaIaRCYI3f89nJ8tqeex3ulv5MgWcIvBjDEAFIFrefrRYkiZAw+98RY2eE
MsTQkJCevfXv1LajzFUVjIEhUBmn1Nc5ylafb7xnPQzmAsBMztqIJ0jMxzRP1yVBNVrVDrklbjlF
xcjwitwhIS8DUAROvzMSGmHz+XkS8h6ZMoYF/RTzcR6iAGyfJTw+KhxCQOmqdmFX2dp8wLG2iaEe
WgTZkZ//5UaQMAqBtVKpx6feqLjH0RBaC/ehQ0edbqKd8MxlV/FMAJv03kLwnIw+krJKoAOn2W9O
JkTtKNS8xXCSQPFptL2mxxwhq2FOgWbc6DeBY+MbtuDn1UI++r+3fItG9kBq+co9akXEiIseLtzx
3VyoBT02rgHeYmQKrmHWzimu+NLV6i6a2Tiw+vsSUueXHsNyG84PjAhwzmhG6W9JWFEaVBjzOQxO
DR7h2Ph/cG1kpV80ld9YhRFK8zmSIpfpx8pwlXn7JLncPYUBIY/+9luQJG92xRBTQaDSNzFvvd9g
397/h4nJW4IDqBW4Xb2SxL60c7C46Y9dxajx7qTMQRJ568MdESfrZJxbfEf++kooWkyOM19PTcTB
2TdnN9yGFZ1u+N0CvZSNVeNB+S2fwGI5Y3c7X+6qnID11ylVrLpH4M49QiXBJYKNwewIirmwVXM8
Dem0gL1CARNSeMRAOUw6tK2c9s481k/kXdhjWADIjnWDoBq4FKi1qC6PbE/+9fTSLIzW8sBpt1ft
jaC8hVUawtzKNhQQEYDzUBl+DiZ7l60vX4UDKE3TV2GgY+fu5zhve5ceKAdwV3N2rLGt0TqqxTlL
B9URrkV4CO12IkxCeLDvlZ8+vFAsxbCM1ZPOWrVpcMSgMxuHHRCUmfcMCJsULDHsDz75Dxuu2if/
7+jXD0yrs94h6eg1IVoQ5vXVpv8yWX+jZ/EE2ZbkrGQB9tpH7pLdof8cbktoYD6DAKHpQGF5TSRj
sSYOmXx0J+FAi+l++QbsI4eA065rewLT9pH0w/KmItLqLzQrB1DKwecJdyeuWtore7THiKIYUOr+
Zoml6p9D7mMnAhRUjXoFlTLF3ILWRnz8DuYzyD7MruUY1sny9DpQyaauaCsu+ytLIUv9hp/6sDcD
ubd+sKjswzIuBaCobm2qQQkP3h9wKxSyie3Vdm8qOqEFTPV6tKMXe98cZCj1HI1zGgBFVwO3cuwn
GU+WFl82cmrLS0gX/COk3+Avuo/TeXGaGeQI1Z3d6S4WNu+nMVf3w7HjnkTeVtl1XFOoB06zo5eg
UGA/O76aq2Cl595Se5UEyF4dRVLGLps5YxMnNRIVaUwiG/VGjjhEMsxMg8lpmptBt3SjWSinVAf/
uKrHXrxOufRBbwwtkSXSiksSCCZQss3Gt4RVHGVXAqTuJi/f8CZ+sxpv2dnZeoWFOMukGVNAkEuJ
EcGE9EB6s89CmUPSsp5A3eD/8WFji7ZBiH9lZcA0PMFI6Xw+JQLDwhJOdlRPERruLHTeIKFhPuPH
kyvGkncyxQphoMnEPQVVJgR0o8eW+qxtnw+DjC/Ii0uRcl0UIOYgDi+jXgzPzXqbH/9gJ7tTozNS
bGtVHERm8gyXIwKoQCe0bRlg2CBlttHAThNNQIPVxWGtqFECQFtDjcMd7k1RYrK9NNuHz1OCEiUQ
FUTnQSIz5rnKqzvIZiOd34zNYv0vHfkhVUKPDHWjEaBBOVskwdE8p4Ki0xINWqPvbIiqTcQtIcsm
aNib89cU9U2F4dCRlj6eBl0Av1FcJPMnbBHtuQzK9EzV48Z1xsG9T9Cidb3uzK1KrxkeMIk/IpsP
ozkcSy7CL0z6WzZv9hC3skEs7kB2DOHRREp9jwy6OYaoVH3/T7TO0UZLs/i3Mvsze5ZqGT1mBbAX
YrO1UmsPgKQJ79Oxewb6bY0kkQi2w2ybE0bsdcCWn1Eymz3dMzeUjB5YKh9l1P6xYG+Yqavt/8q2
5fPZdf29bZW7j4voed4mWX/lw+PO5ueBlCMVCtbyTtu32fDf1wV1aadwTf9LfFEa7yng8CgIfFss
lmIGb5Qb4940nuLJZKw1K1z9A68nDbXEtmFHelJnc9PW9J30D6T/Ag4uOOsf+GhCg/cL4RWBIAbM
ITslQA4sMJgJ/eqW3tZcgKm3Pt9iEfkqwFkPf90Ye7YeaG+tlnnPemC5UflPi3Pqqw1AOzvsT/4A
Vi3e4KcGLpPWjQhjsxdwTjX3hIVgWMBKQFfD5TFQm3rM+9R4A5PUVYbOslWH0NDdYX5UXciT6sal
Wjlq4dxFU+72LMDXYzh9RperwJXvcmjUVD3AdcpXJwYIxcN/573mr0G4e705NecfqdNLU0idhl5l
GalrKrYzrzNtcu8mH40m9Grlu5m2KQsLQOnujn9AXL46tmhBXKBaQ+Jw6nxs/+E9FcjV5TQj+XFX
w/08wHiTtF4IyouNu6RJxDwQFVtaCgUsqDF8vGPx2+TjdvVgRiuJwO6rbWIzGt31wsz2SDqygyEC
0YxA9gPjrkfE6M0pxU+wGbFDvg5TtlJSViFQhJRGN0coYULNx//fklcH7lADEfsQgha1xTSeuMLJ
MBcihEg8Z/xQKoWsZb7sbYon/MMSae3GIoQ97D/cEzt9yr0zlj0J09dje4psKZaxZQR6pEBWtpU/
cToYpEEHcmHYYVL/LA2plzTW5VkjUVw8r20ntdhJqgOKRtrVdunp5WlZ1ZjHx9nXqh4cVQZxBael
KEBgQw55B8TqP4RJeYX0HBM3RvfhuZbS/eOa1gGcrximN9O0Di1e84h3E67YzTo+liCgmKVO0Q+T
Nn2BvcIT2Th5of06XO0JugeJsdcqa1/8Nqb1t9PXuTvxB+SjSmnaPNfZcJPfLYBBB6fJ4bwGlUzX
QO7MM66dyCbgQy00JHHFRnAsh5HE4+FRfoMEbM/dF3eRmrVGJXDTASXxBw8GY+nDhkGGKvUlh1L0
ct/lInYJHYXKzKCRtEo5Pq0RwQ1mPEuEgy2YjJ3HEXbVyNBY/JJDzODRCFG7xCr9e3RMxW+JXoNd
Ix+NttfHBN0hEN9CcPy/ZUuF29zNASfKzNAAUkuXQvwUd8Apfi4wnV0AynZ3vCBjKFQvHoGMnNZJ
z+KywEa3OfPibl1Uzu05Xe86uspsJSWwM6mZbhHtj+rbPWXbxnwNCbOdCVcovFaDm+FVwqz8APfF
4bP9aeo3Hw0XOn2Y9AlvZvcGl9fXLHUE8F03NugeO0wrrJZ6f/hCuzZXgvQCEnrbPt0ds124E5YB
niuPQ/sEyDbsQnHSv1vxklrcCZ1DVqYOq5tfJCMvkfXSexytNbAGGGcHEXb4lzeos0m3ijo9eSfk
Jz7EwUL2KN9d1Y5okYRVkGyO0Q+nDsun+bqUG7gNwbtOw1aNlRcMXe5SEBPsjLmkXB8n2MGzMqhO
rjcohRUNu9QPXzC0ZdkgzUtuW8MgCquYzJ5pKaGA1mTEA16wd1vBEfTRWHkrReiYWCYPMIKzLJBH
5/0m5RqttTr4ynt3d05ARRF7qn99uCWUUtdVAoutJkL8R+jma3H3Wj6+uWk+E9tdZkwp9EXTESDn
HuCaAemy7zWjhsdA5Grs7hLW1T5cacJRn/v3lrG7sS2XMBoGotu8jBomGWQm5tne5jxKLjFZDZZF
ZYddonnLFG7jbAQux0+FIh2xSwVlNFJsDdR4Z4UB+/V4PXBPOMuJ5f6w/Bw57RXNqnzKGzZwWj8g
VdrbATL2Vh/7KfKVcIPVZucpeKTswwnLTXBwjwMhpTZ6n859sY5wT+EEmwjnNWg988MR3DPO9Zz1
MzP2FPyUyooOvGc17S+Wtq2Rn57hW3RBOtqSbkHvKmQ+k8DyEdiXiDrZQyWfG5d3rdYnbJWIRYLN
okfFK3mhRM4eWRmhlZU5ukyKjraAluVLQs+niPhVC64/IneXJcsVknK0QjOLHeknV9YGlihMgWo8
md1Z2YVwchsrYgzaw8E+hLW2i8obZqG+6WUylfSC/bWtgHydfC4B9qrhkP8uTY779+KgK42fA4Ls
a59VWHf/iheu1ZOfSluNC2MamK1BWcKwVp6dIPGG4hbUnHDM7ptNs8l9ePGN2F9jx5lHldMUFSpp
j3nJW4V5aDyVn7+2H3eWRCUCQrpLPc3Cj2qFXLzEHuKg+qtkjj1xhVLFHWJ9tyDuUA/j9lnLtAr8
LLPWajQ6a0pqm2dnwJI2Mv2qboPNeY9Nvmm/81f5NUz2Uzwa+SO5G3/6Z56QhijLQ460c4jHDwj0
ewvDlpGWaBuQKdgA+N6G68y1Z6mNbKhG24cMeA4rr+CdGXTnppZWC/BtIw+MoJ26tgktXut7itUm
fYK6lbqkFcDb+TYQuOWO7QoqiyxKHWRWhPKZcMbtEN/MnWJC/OEFGhUsQ3QHXy5u6408q++QltOG
epxMuZp4rz7yEy0kfyH3vAhve+kZFfBfubEPifJGC5OIiDS+E5HT6X0/7J/wcF9LaTDus+dQY42H
grGKYleWXS1TdM5vveAibdpQg/qK4GFNgBj3M5onF5yfdgbylXGZvDC2ad9JBSsGKZtk2wYCRlzc
LtzzbngVb9gCmaxRd16OpE9qJuOPEADtcAzxb1GJxlzkp4e5UPmerO1YBZzCr7ISUyxp7gSijveq
s3YPDwRcvv/f2wha8rwkIWu0Pwj3QaSKFxuung+rCMJDthsWpFHO9/FmCak/KmU3oBe1GUft/76K
qi15kMrdaYcCJSogYhPgZuybM+p/hyffJXqePAOEba6p00ObppEyhgjMGlV+F61WgLyUtpvs08e5
ybr/LGclmVrlk/+4hteQwg/K9uCBeV9BBnut6oFlTFH7AlPjaGF5WFXyBXhXurJjTRSpJ40Hjbk+
o33S+kIkau8dGXEOTM/2/xv1bvXuSVX3B/5cmtoIzV0ihWL06fwdbcoboi0IsYXN027rrIAW6i9D
jdQXL0aMXbYXWaUrmzOjdtFZE2X+IsiFhTzVB+lCn0SosVkQQlEs2pooERALCmwhqcP8K5RHJV2o
nt80rrW4sEYB3fBB/Y/6UOSzirl+p0bXuuLoj97Ksnv7yYRx3dav2e4GJrh+P/De4qhSrPXHpHY4
+QJvLLmwIi5IJhPE+CDiuQIgkMNn8ZPvCbeVXGUgN2l3DMhAlAXAUjUzRhl7D2r4yfGHQuSUyBgt
mq1bu+MtSbKY4vdr7QsBkJER6w/Qw9mvjdEzssm/N4ysq9H35a3R0Semu0tVsjUXUsp0apHtHBZm
ijeSmWd+wgcJIds5ki6vqgT1xnziq6pJ7qrDDhtdiX9sQCH9ghjtqpyv5PILIZqnFbDcThyl97Tl
JVP6ZTn1A09xaFUtw3YYZyOTTEf2HKKN2A/mfgrgh2HZDU9nYmgAjUhFo6ZjEbRgZfSIGqOlSurY
aUcP5B3ZsCTMK857nJV2fziUNEc8gwZETOsYmouN8gmTEAfikJv+CoSfmeBaVJXBg+chfTTn+meH
jZ9EgLzEhzGqv9BAUGOjVAnGEihF6iufm1gM/x472NgT7xrmWHsTnscNq71mGQyKigX0n1iBCmui
IzBAmoOYHgtCjurQ4Yj7CQroybKkgtkOMI6ZJVJmNYWhG1Zy/unPhaNWpnuOTwmhAzQ7kGpk24mO
Ic13FjAO+XaC2kT5vsyL8VmASpgaXLIxpmK1M7gBNGyS7sXJ3WSuHN88a92K9or1NX+Qv4Y/JD94
2SCzjGneTnOuML8KWlsIAtka+BHCGRLNERP+pSvmFqAfm/VOF32pit/UlGZ0n3r2Pjq3BZ5i4V7r
0kPGhimv6aX2+klNuFoGgtg4iMImxQehy2Rh5tCoigTSV6wtxpmijtEtuQRyjgcMnBZSXDp9MBCc
H+hhT/aWoXFFPx3VPCaPXcu/jS66iJ834PcXVTRGCNt16/X5ai7W74tRFrQXi6dUeqSnIDRCub2h
CxO+8db6Gbgq5ccGDgL7GArExppDCmDUzwFHdVatLh8cFwpwhq7QxU9E4EY/7wqcyFXgEjoQB2HE
BWEZFBIG9G4SlLPkpZlw7YrF55X05bJzsov521LCiWU5Gatb52j6t+bZJrcDmW+HBIooWqgi+sXV
oFjCozb5qFxUwL2AKhSFUYMvOo+zmRo7dm4H7cC4H+kntXwda7K1WJrPAz4Hl+yRP5yJECT8g3nl
CVey29nqYbpO7rH+irSx0/H80VYUg+7JweO0T0jfbv0y69RDO4UZ0NBVrVHXYc23Ge/7afPH0Wn9
hQYlDJpKFSUuvNwIEXnHGNifZ12A/rR9kbJ4FvwHYYxAO9vgYTKrXngp5dbGWYwYqYxSXSRDl78C
/e2CViGnKZpW8u/eI+Jq0xWKsLPPKHT+acpIxEhHMbI3usWZxRbhC8L7RnNS5YgpM4VuD0JkzpvB
G7nrJKUF39aWYwukwqGcUYbGokW9WdwyQCpVhVCSCJOT3eUsqTb1BTaklJddklA2w5Kbs5mBddxX
Ymkk2I08gDv6WqJchsXcFUSkiBglXbXLExh/AQcnLSuZPNzEV/OKsasJyi16W2p3Vr0Iz/7jRKC8
aLozOkiPTfKqXIb8udsD6YYpYtsrEjGThQrQGmoxoHMq29jZARMZ0QrfY6k1RBnRqnClSBNLyqUH
oOmsCj7REbCXeZpSZ9paCC6NGqoAiiq12ojxiOoHZZJFuvQBPLWFGcHlCqKr2bdEsivcQEe45qkl
tDBlGIPhJ0MDKNZ/I8lpOMyYnHiaT5aGwC+UcL+JXvPgTrcALoMNq1r/vEEEjIZOwg2Fz3SvPs98
LBoDwxPSwyVIoKgfH5gDXdgV8cN1HwfpnJRg+Hs9hgh9stGeIZ0HSYxP4U/WZ5d34yFEQnDPyTEc
nSXajUmuJzpp19BZX/V0iPFVDrTyW9HLHN2di353ZZ54YZCELSyYlr+4Sdd1wBKlFLOkHy0T8wnT
UrfKbG+Td1LyhqoIGjnBfx8quJB18RnCJRS4qFL4oFGg8AbfTwG25Pje58AhGedimxg0AYrkIN6c
XOh4b1v04VwBBr084UGEH2z9YKeYk6UwPCuNWWIgqUW08ETklsu+NVQjUv208tbCWO49fqLDvFVo
o/NyBDRxWmmAZa2T6wfMvDhXHqSJ/5msdx8gpSn3n2neYBOdfHvHUl+KHO0jIm2SOD+ljQP5k3lC
/LiU7VcZFghVIUxoJcEg1BTDX2cHRs48Al84eI8euTI3H0mRqbR/16n8GGw0Owf6tEbXG30y71ed
WIR6Epuxok1MFUoQkIopgkiVK0LtaarrghW36ErK/oKI6L2ppNG/N/nN9j1g8/VmWeL5eu4UenO0
GaJBj9v8fl6pILTH7QZATIKpD+e3VO3DCECdCrZvvFPX1Qi0jsxAHfC8kLN3PY+CpHc7lsqIrsl7
NpgthNf9Hsx0mCvTkrf+cv97ZT2p+UVDsSdIiDIPg6AEop8+MaE1unwe1Y6vhOijFSBiQopVnUZe
h5nSvT9k3TCQrzLql7ZOGhNPQYMF3ywnowxIeukzN0FJPlVBRy2NkMxEUkvhbyHMTcUvgq4SY0Xn
vtV3DOwx440LtzLm8001jXF6lHS8D1FW6p7yZWOQ8ANKckZo6gKhovA6ULzLIOhD8qxwY5wotGPQ
1AdTPcrXxoi1E0g5XfEtCsdM6kC2SQ0RhVnZG2X0FpCN5oyRgjcCrVRgFAJ4p6cYS9DfLhm/FmI9
V2QHqtxMdn2IPI16M0zOp5SiHgIy7xXjLuiQWXgdx/gSkAHd9eQS2TPmu94cRBzItUcYGUdlgYQZ
e5PrBITXmzs99vwtkROrZg4Dw9LwY2w4lAAYQgrJu+8EsWEJaCnZ0EatNn0Ljh0N67xFmpMB1W+b
9H87bGKikbeVzA+NUZ8eE5nItfiXiken8UQLXT8n7B+F1QwOedPYmnnEcKCvLBfg+lgvWIxi9Y7t
qgMM9tCkhLmxBofahbPAWq0Y7xAxFpUZ+fISOMiJnBeDUWgvCkxaN5WHJZKFWet3Nni5Hs1lIt2t
vN7hOonRfitfi59ACAfONHT84c7QUSz5fPXeiZzZ5Hd+jqHoRhSVPqWO4r6NDou+u4suZMIpOXHK
s7yROBsndivwCw46V12w0QJ7p7gZ557qwjmwFb5Y0jYjmg9eEN8Tysmd0wr5EZML0+BQ82sj8Yig
TgDj6W9mJCM+weeDU6sOMbOAIqesdoG2FFEe1bnRhWNISsT/gSFBNFcYI/5fZmRzKLv5LGl1+SmP
Zqy356WwEPqhJFpGvfdLv48XPVJlqQj8nOVXh2fNouYypu1v7+UeFFy4kF5IRFRoZoQT6uSTUYxu
FnnheKXRMwUiI+2ewSQ68J2B4VVZ3T9odvdC9r02RnFkkYMwihVsk6nUIxWAmpyj9dtk7nBJSTpM
5J50EmDUUDFcHdVXWap+3DQLuEjAfKTT7j43BE6X96Td7Na4cBIgopjVIr4TzEAvv9s2oJ2G6s4/
T475AB5lVJg0jJmEKK+3Xz5DsnNCmY6D0FY+s8f245c3augaFE2ICFFpF4senRk8C5+K0i/Lr1Vp
NVTVVsoQ5Rk+a/RLhsFJ9QKGGZJi9As/esTYFuOxvXGBBS6BItyi2pNsPhUitG3WvomVGg7FAOCQ
K6GUhTRGqY623bAjiFBisSYnOctT4Lh3Csw8pVuxDWXeKY2/Hq7pqNih4hztftVB+Aah/goEhedf
vgZKt29J4JCPBc3P9vE2ozWAV+QsfrZEg8ke/WqPs4dGEXHEqnLzTGQjMEgpYvcB2yYAGs2fKsEn
Logk65Gawjjl23CvW+aQNO4fs67qIX5wKJ8FCU8Q1/7B4/Ynu6xNf2aZw+UU5bFTP2/iiJ0b7CN3
0Vl5mphKF9LIcPta9+13S2+t3vPhNHGbGLild684ldgHac/ffvJWQu0IEkFyBmEmgHvrXtBePJQN
Qsz31RFMr1/47Y2mSqwxnmcJ6U5EtHLb9Yn+8vS54e77gHGAbB8Nj7hsGwhtsA0HbJviOqZlqtUl
Xz++HDdB2rPiYS79PdlOv6OIxV37uH08ORI4SzYkkIMgpMXHV/4M6hIYw4H0z5fb14MgjKqY41Yq
Hi01CDsirDIpmic7ZVpSKPJAwCpXp5wrnhgaq8GkTyiJVuqWjPrCbJtxZD6NhAb3idgQbMI69jA6
kyTcO4wuD+kn7d3pqmxMO3ReblzQLrmCIY6z6xtqt0ABz2mAxDJHCWqnKIT0rjeGCpJDNCDhcz9p
PNRjX+fMCzRRRhILE5/EURgyJbAURGvfV9OOIJSkx2jNqSapz2pnj18hVptKfawp96nQi169XH8u
S8d7FfBg+cLaKNHRz7uScUYzIO7D3By0BDR/KQ88cqMr2THCLW6kWO3MmBmThomfWRQK7CpHnlVB
eUGz23dzjG5ILHF6Svam3ZlK2fRWjsxPjwUWUqtgIFvzZe/mimBDRGjsPWaDkPHJ/qXUxQDTSB5c
F7vfG8XmDOyHSbyr2M7+BkOnjFtYERrDoRIoncHquE5cbBMLXfsjzChrRByU8iyhxX/KimF05SjE
v/oje2pw3WvsyTYpzEh8cfBPt5Z6KKACNBWdkGLSLZ8y2g6LOLLlM6a1MdOova+L+AIoQYWgnhX5
JYG5daqh2uaDbRrqCurcrVqzdOahuqhj5His8ZgBjwBlBP9wDe/+FFtK/lQEEklozVChjmBuBD0x
0A96DHKOlHZAOsJs8Cfcb8pilzJQWcK5xyQm6zjH22lFxz6CfaEtTCpdn+kzv8l04l9kkFE1Gn07
CP1B9h/4BMTe7Y2D0XMHLCwZVE9W++qKmosdmkI3mDGWBz/xZd1z61N3u5PsxFhaMKiySCNy+WNa
Nu3THwEmX+jueYDFr8XbtUZE6CGDkK0XL8m2dlDcWWFVgLmTeIlfZQHhFyho4ibbItC9CZuK52QA
NhOjwJn1blgxsUzdlsNnKZtblenWTr/DYDdUh8YT842dR2M4zsfZDwmx5LebHeAWkNwhGAqW0DQH
0AVS7M8LYieNRYDtjuYlXEGXcHEkXJUG0ohNYUnGlS370F+XXFEHuHV55U43vXn89JI/Fd6erV2a
LFMcWk/U2Z1AyiR4AU/VbdASkqC/XW3oQR4vbJdkVfM75RXgftIXVA6XdTA26hmKrrOh4jGNTLBO
1M1LCEIhD9lnjoXf5HlOjM4iwEXF/AaMzDsp6w14UF2epfYWU4WuF1lGBg7imrlsCGHdNxkatPuC
ydFPmL1BY09om64R6nfRJuzF/DmAi5ddkhY/JNmIY0hYFwfbk1RJF4lvmI3hkPudjZbqgXoFNIJ2
E+L/zP++oHSowsPgA89VTmSynewwbK6eOLG8EHSUs3XGR20167huHeHeedzd9QxiCAu41pOrMqUn
cU0CGkb4kheNICqPIJObg9fefPCd5p86hrT6BFLZB0jwX3IxVzuJBot9T1XU4AYXFpkrz7MY+xtt
kpwJHgxhOM+UnXR0xkSu0HW2e/+kOLVPWD3HsAZtPY0AmspZcpbE1CO90gtzyVaJa9NffY8fHY7M
Ovw4VhED0xS89x9H/InbmaDc1B48xk/MERZZepFWXXWF4w+L5iO0tp7ITZrEjqoN0xDcHDV4C4P7
2LYoEn5Cm/YdZdqe8o50+OooNMgWIksnp3E6ZYYGgcSsqPHl/G4zbj2XZDYaigACY4aZ9hWsV78v
2ZP4UXirfp9tOoGRSAPTUDmBNSwxeHWPrqL7lh0cNUMyrBz+lV7G4XrkQwPiJcJz7dp1k3nqIUVC
TXf+HSWB3UBxA1NjKXJjtS/aaTM4Y+ZRlSOZCYNjAUZYAdJbonp2MwDyH8wHRLh4sNQYPK6EwBsd
ADGq4MImb/xXSiGMRNtNsGGSIpourXWEqYyJUig6V9VWJmz6M9SdIsonKpT7qPyYApugUIoEcRx9
WmpZ43DkjKoZ4amvtkFziGNE+2vBCkVxVCB4x3D7plz9sM86G11iMlAD+gfUKiwe4WPpRcdMRwTS
CEJtAUWFenVqd0Nc6hAK2WDTcBeN01j8+6b8wkHoiR6mqejsd0TtLSwCBhmUihG8aaUZpux+ua/t
JcgXa9cvXQaHzFMK4j41J3P9uQnI8uy0EDYE5xiObbiJr0hwiMQFH2TpxNvi74Mts53F4bm+KRoB
EY+7F2vEVkA0YEFmk3Ep5KhL/Q2UApgs/NiHrbT2AyGj/mUH05GVla0mzAIKEHkTplNlYMT1XkJ+
nbkY42YFuca7joevdWiH7TC5HZaP0ONbvy1RnhRLVpKiNVcgVwRbKB5S6rY8eEc77Fk72EOEK8Wv
JiLFtyJviO5yLUaCNzdMcEyM0jAfDqLaYc+0oO//yNVv4LWSKDmnRw402Qtrecw7//f6gL4eCxyC
zL+ULeBpg1hogaFP+k8h1Ex5fDRvYod7lMW8pICB7hdRQL2DY7j4vwln8hj2BX30X3watMfc8lbB
CjFH875uis7bmW40sYVBzTNm7EgZ4ZiUUlYGETnk/i0HzTZ3zM7Nq1y+WP5v/OIVgu/vzGLphhXY
zV5+8DARccsG7WHjEoiQfistGNsMoy//6mHLsXhQjfE5iLbPJQxdk306kGpkn5QS8ThPRe5p2Ere
uN6D4WwTflBjh30lQzpW/jIvY1YQPXSPaHLMRQH7XZmuGQueKtMpj0skd6igOLZ2Vl/7Kj8T3jMV
LKgc4oka0Os6wg0VZ+avvFU5AZzmICcsF+gGonIOPGMO9qsQ8R/C2aVQyENxGWws0C6OM+lpWms9
LxOsQRO7XTyGYPfP/OyPWR8ksIwYbXynVW5AhkU0aLO3gxCgZsyAw7A4B3Z9XnPy8fspqfAV1bly
JjJL07rJcJpvcNcwPLuZBUEZOfT+Vag0vk7+NbCLcdB+2Y/jDtaxKxmK6cb5ASne1wDmHhhkBKjP
ERH+KfcJZ7AmbDUeMwGe7UkaYuYONtkj+mvNZCDwb7FijTeXalFPWqA3M4+qYPw3EEb/8Im3hUrg
hNramvWGHbncMiktoYFajuTpgh9plXQZNTBZ+pfFxGGSQmf3Nds4q6QBNGUKnU4IywvyHUc6OAv+
yDhoU/HCAh/6Ry49eM4adP4Pcj3KmLHZ3ByfUhnlkV5SksYD9d7vqlA0duUQUHL+P93SwUFLYUjD
cVIXIEs6YG3iBpnfYbbr0XyuxYQCPdKMB/jiNOFqTFfzB2eNzbKzvi5VVVHDifyqLSXcY0Z89ekU
2mMih9jhZaQJIekmbdPajcTdl6FZSVh910ii2Xt1syuNVl5Pwh269pJDkZyrKYq3m6/KjAtpwGnT
yecEbJz1BbsZqfNJ/T2emoY3j5WA7XQzFNcETkif1H2bO3tpTckydT9em4B4jwFl8ArinY46fRcY
vE/veYegVNQioQPPJInVdzmf2lVLg524JUjoV+x/ebCxI0nazG1DLHI10IaJ6Xxm+5GFMZoIHvsJ
JK0VTQZ0znHLhyhWGRttVo9rxMGDoGe45a8+HheljGtXllGerpT90LZHIP1DEp/A3DRXEmn0uiDp
SQ6WwjXGUs6wb/QVgcLALFqtjhxgXpJ43cbQXR8y7gNi8l0bOJvAVdfl1cWIPsSA9KJa1PSIsADY
DeuM/8wa371ZijLvIEO5uLgFrP2tibCksWHX5YYjrxpRt/l4EoQA5Z1E7rhulsAtlTl8KuyKO7Ey
FlPmxq9ay2RvR3+4rioQbPM36VhYXHNrGsZ6lxGRXYxbJPzDhyofz4tpvr1v0rrG4icfllhn96QZ
9XtU4zfaawsVWEnfHU4Yj+bt/laurA+mcGgxJ4cSqnUUwJvmg6yfuXA9WGP9jWQtyl+0q/cSiSc2
FH2KaBacQPixm38DjESAOSKRrbxFpcwLSMVOF+c11EOQZ8UF+66PwqEsrL0LHWE9q62n69f63n07
XLk51H5jQibUWm4H2R2LCLMFnY/NsMrG3Mu68EXcpVzR9tbFNs3ePJjFAjX4UN5Q8u4Je66DA/OI
YV20euFtbRuP8Qvvc+b8jRMqQRtMixzyFDAt3/3LvKXLStmbkGERm+KxvrUPgsCHkJsm33bSxXb4
VCOXp29bWHGLVb0kNuYNYjVbhHUW6sYjOnkUWiTb75ldt5G8FnxGQaN18oNK/P4lAQJ5jQk1LLtk
l+4ib/KwQQyEwydqt/iS8hTFwonOXEg6Rf9hpy6RpUcyte6D3gqSMsX7bKYY6JOUJt0w5NIx1l8g
w6fiotaBP1Uyez9peyi7I5VpvyvarDRCEBzGLMySO84vlLMEw70zTeovIl8kccBBCOHZxijXXjuP
hPCx1e+hTdHqwGhATnmDfeTzLihnrDdBiFiuM/kT0z/p4aPby75ROcLyckFJV0pq34jNE/J5uZQq
5PljpnN6+suqzw3f7wXTCI1+m11eUrl5GETwJkFz3aBqp2xPb5HVkTZKOOnWx8CxZk/GnHE8okDI
F1o8xg8VkuOmltyyKGG8loY3A371wwJPJwM87zlXiQ9VHpfUx8hjKHWhzkwNTY/it8ddCb3orZad
NqZtxpzIBWsoofhmy5jGTxJHUWQveflpIc1CAGjVnJ2irKsYOqJEn55MRoV6uZItmKYLqWlzBFSH
8D2MAakkWcyxF1YsbqvnuQCRiFyv2lPgsh2few3mfUmcDWj5NvVkLUinHuv17bKaG1MTGdgfqucy
wEGFsk6iytGzqENoNhC1fqjds3QG0GizSYM0E1zLfL/8yTH4/YNQyWt++yJfolDy6jN/pPdnwXRG
1LM/4VJHEWv8kuzteQkV6L/NUGvidT2xPRLZhEaI7tTYEMcbKvuyZullHkDA+5XCFuiOwFOt3gNf
9fD9p82otIL42IKO8m5NP/shYe7GdBFeWyvrVgIKgJgvvGeep/zPx/DCwU3SPWG3PPI6BTDS5Np2
MjlG7wW4w7k8nGtxKJZeRmWkdxQFrZv2zULbjKhm6vH1Qcj3rlh7kPuagdB4gvpYRKpd8tkI7FCK
qE6DYdpDlgBcUVtsXBLc592SYrNH0QvbVJi9oS0ju1VTTb6VCVhR1cHpcsIhsF3YgvUmV0Ky3+dC
YkG9zEFMEJKuuNe3qoNd9kiWeHxDccr/x+hSKBL9151Pqq9veUoWH7ksaTnNrYWl5BCkBRiNNyhU
ARbucLMr3vHHTf2XWNsUVzfb1YvWbyfesTH4JW9TE121HR9esCkBBIy6Y+Hw0CiIqierN3AKKSwd
caYvLmQg9PKBoVlYzQa9gHU3+qce9GVR1FCBWQHlLYH4GR116X7VgqHO8Bs0XxxllhV14etDFBrJ
TfGTCCL9Bh4GFcG6xNd7qijcRMqJ7YSlRncbV5CuUdZVJ4V+eWWVvcK8YplfrEwXK1+2481/fWvr
e5PE0Oha9XvbEnPjeaqmMlZPFP1frXc9nE6nEo0hszz+mEteef4rewwq7fIiRt+LaGyW87Wo/hb3
6IiWgYAX/S7gfyMM38LRwUkKXTmtWUW/I1EOA3hvzYcsNrtdUkwaDMqY/QfZhKxoiT2AdLzs8wYG
uvHF0+/I6GT9xjRnhQ045bYG4KY1DWAjSfAa9OA0Ec5RXEMoq/vd1F8kb7qgGbHhBWoWsUEYADPD
C4JCFAHocFYrGnJ7UbxtZ1Yc4jF51gkvVegp+KaKVCuaOK5tTJaulNsDw2KgXGxGSnOvX0+HgQRX
NOtKGtKbxCSoet4+sLePWL3oSB3Qdanupb9GgCxTk2JI4K9o12wo2ZEpo2J2BdWs/g4F/cJXSdEe
dgzPEP4/0Y5tC3vHHMJ/pd+2gglGv86MqO7Jjen1dOuZz0coFOsCXXCY2ib+O2n/qcjpBjITTP7t
JC0ftlT3GoJg3Xn/s8NIKUR/6n12L17P6t9uXTNKpHN/BSM3tHkoetek8Jekgx7fJsTU/wua6UVG
JAsx2eWiAdbl111VlrSj8A2b9a7yyHb51QzwAM/GdOHK9dEOdsgfwIaIj30UnpnC5fApZGX1IE3A
vsh+2DSI7aZ9XedHEuUyHDuyf3mpEcO5c0oyLmlVmGuGpFb082wXjjBeGjVWc3+PxRmmoiVciOkI
0ZD7HGTjzO3nYdDroBP2HYef5Yz2YnzIYHfqt7rz9sIxUMK+Gi4bHnDrOsEBdALBYrqNHoc9nSt2
tqpwvRue9py7vdK8/GkTl7mvvOyfV3rc5gV9YLgSCllE1Y8twpEHjRizuj9irWxWmw8ZqE4kZmyf
HgG3OpxTBip+podYHEY0kDEhPFxnhXdDCEImM+SJxhLtYACZCxg3h5hyUtbc7CT16Izt8EuaBJEk
JVI6pTf60HGZEXn8y2dufSAO11KRLRiOQDjy80WWcLVuK0yUG713+tulIkU1AWWn+pLAU4QecYiN
dBxJbgPdyVsADIKl6BiaNLO2UVS7wpBXegbK3kPBJGNM4qVpg+T1W3qNOYCy0aMsJLXmjMogu10E
hGO9M7Be28zPxGOKH4bkqVOu+NLuyXaXTN9T1hl5ziMixcmfLuqvmu94Zs11uiBUdwzaGi0v3d2e
je/eVlQsnFyVAYhGDSu89kUFHuDhywaGpUpOfexXRNnLsxmqahX1Vs/EfmweRGrgLPammeOHR0Ry
uqDf9LASbPLvYgflmUZP4NtwA2zD80FVWPCE3FMWrbXX+y6tZ4AnMzRA8FnalXusha3nCrMigBIk
RoBggin1+ny7QYREpi/1bD20nmqS9jxYJgzYh3Nx2woW9/ulRNmJFuLVF9IZJuEsMm3wnMgzC6Nd
gvo7tPXvhGgaQC7uwBoR/54GBCd6PDvVtgEx+qFHwG9Hna7eH1tU+JhE0KH70/nIvP61Ic2XIUBR
3R5GeVJ7P/YgJI09Q195tTsnE4yyhhAPtMkx1vADtGyWykWGRGCejNwnnKBUBQ5uDCv2s+EGG8FR
TraOWUKAw91eOfivql6pmQYWP+fzYOCDA+EZnhiQQFYKGW4dAxdViBeKVGcBjJMGBOZ0m0AvzZYz
teMIJE2R2s6sY9FEaSPlTmX7q+GhdW3f13E3mo7z2sxztVSd/gUxTWb07vd1qvJhUvA6Lqf982DB
kcsS6wTAU876kQGLCavQDI/D2vXtHSsQXwQmIVupxitnq35QDSFWDMZt3HJRQ3Sj4ySWt4q5kVAO
JkajvhO0wAwQ/51HeGyng+9jhr81FAb07p28EOw3dMwQLHM4dX1wB56AAG2SsqmkXBeqsINterP2
uez+j26JOn3sVmcv/bz5UB+zlnPbAJkkANp0D4GraQeb62gV3l3AJOJj0EcKhMEV6pddKJoLFxQo
DEWiaejJHoes1nl62AqmekIBvRigureLvgJy3kdLZW1aKDs5G5ARBMnznxGXDyiAlcYxjDj/OrVJ
mt1LsxbrD5UFYHbuA8DWSG1pDVCFExy/cxAR8DQvNTTXewe4/v8jwG7GadIBc5u4TwPVdnEzAlAt
NjmQqfsS1l/9abOW2LDyfdUKmTMmX3ZVhYvuO3fe42qbVL8akUXVfavRoHhaqd+me+XJcc2+r6hj
UIsasoJLGd/UmfkH5LAS+Vgk9tZPLsYlB/5DjSyrvFQlk7F1jbOdN5f9HQqL3/Lg3sBRz7QcQzFe
2i6Y2XavvXKEqUDGKsTBEj94EW7SfGtc5m0iTDZ0B5gZ9SpKMcIovQIptGEgB1o2HzEHpC34KDMF
xBKog4O8n/O8fVh54ZmRdLXC+/+FE5SOqZosub6fM0IYh9sLEEfNZN2Bq3G0BM4xjpCVgQTElOr1
skmDuPfsWx3ArWlEURZTmcxqdrVdxq6a7TBYiHtao/lqoO/OUVumk3s1wsiNULFcW5S+JZIYq6e1
Gh1Sk3LA3hzhXplf2bhJM3BmcEIZMjKYyhVjIgrrRFevR7laFvH8G8e7eQT2uUQVOR6Py3nb/ECf
Z4NlUGpW93kxFOSCdMMWBl60sfLVOVHWOqKIOd/MeTv7D9NjKETSAZGDCkF9V6Uc70xOLcrmyaQM
+sh942s6HvasD5Itdx0yy4B4VYdpuT3c6OQlsIowwqdftjN89YbancTloHVBJ+u3uF9YaCoiA+6y
CGGNZPJ0xkkySonjw/U6qoeThLGu1ppRl+mR4VXAF7NFMffam5JSVgebyVhw9IE9wrtqfk4zCrkB
T96v4ZAvpK026cTTi+9K86Guz0hnq3axxcdJRXyMKPdZ6rp8M7audV2NtdjxZf5BNlq8JvKvoBEv
+J6xX2aSwcuNJvvg/xO26UCrS1ZszUzhrhj/QqMnKDmvAQfbPtryU4tQAoTsem1clfEctOoJ+tYO
kquR2d66Qpj6ZfDES10x6kr4yuRmLoiko2t5aJWaWJI4yCaz5TH25W/MvD7ahBC8PqRkm+fxEdUb
YYH+0VXT93OOfoTtJ5L1dd0j3+BhQ1Q0xOwnfEeUPOVNb1IcInJRZlULHQd9LycZDg77JVcBswZw
ep8bUtv3xC6U9Oik79DnlNnmo39Ve49Mu/iY+2EIKtqpySjm2X3LyfGMS0h9u7tm3SuG47nAJtjB
LryPy07MR/Fx996QzYob/jOPc2mDEkOsjsZ/9C8f6l4pDhHA6gHth1fpeOq0kOj0ilb9u+NbjuWT
4YBTxp8Vg/o0Rx7+clOc/Wra7WSH9tFR04+0iaw+q5BgKooNJOQNoteZ0qOle/4pd0hPpuo2u5Ve
HCVR7iFxDvT954uilNhSHfDTBRPKTEURo+azqP9n7c5lY4GWhH52HOJwEGIOhNeDeAms+BQ/BaCa
zSvN4jLuVPnHrc9xg2P8INpBTEwHM9SLvaOrMEfAn7UEYfgQBive9zaySJ2vMASKssqzd23IVKfG
qMVxtxifOJlZQkCYdZBVn5l/AQNM8edSxXWMxBfkLFlQa+OK3K7Mvw4K2bqdaitVtqqb2Vmb9XQ1
pvv9UMKoT9I2U6GbnhQ5KLAyBe+2pbUNZvNW4pOPlFDCRqyHiHGW6BeGTG4sNO43S7yLGt67qqwG
mXcIuHWf0WWhqN1ZFY/I382vCNWp9UWspI2FEbs35nmE1eXZc0ZxgN17EWlrT4p9xLIyv7rD83se
XjR5GKQrJg82ryMfGQO6D2F9WoyqqGRjS4YEi2BuwrE/kUO9Enyk8JXMpMwOUYlL5dFoKjzAuwWT
dPIKckp297FCxtTSTSfOf2kpoyXEMN0o5egfGRAsV7ZRID2AD4rDrpc8pTt6B79UsyrIOHSdkQYK
Luif/+lx4BiZTo4CAylXWcx0WndJUDn1K8sz04YJw/D0ZVZrDeqoSr29uVUaoDd10Ud8ofLrXWC0
BVccoYhPUk38b3lA+qyyv6DH5dviboathVz4z0YhMgIA72Kb3dTomBaz9P2NtsRAWeyzgIxi6TDs
Ac5j32KejVdwwOtAGvjuDGVB4RuFCG7EcnTAAECc5oR8ruoBrYA1+8wruWOFYMYUlPSR/OJ1BvMN
7BMBix/rf5hsKRHAMyn4LrCnmVEZ9JwZ6B7p0LeOGmhKRCliyiHUcIrfjDDMpdO76os1JKry98ro
9dUNl6EEG0MxBj05S+6eX77PH6BrMJG3CnE3cqTo2XEUiX56dca4OSNGIEuLQEjvH83UU9y7djo1
MomU/wE7iDWgYw/Uxp5gLOxwyjwBJY42rHZ0iaRCEpngZcFwM6rtZRr12xh3lE6/oc2li3HRxvzZ
pjrVBgc1OBQtlAeTasvqkP74j7+sN6iKCoLU9HCdS/89KIac+80haPJwKZMjE+8f5CtOzM1lZraH
lU9xw9mnEpEiy10qrPB2CwCxLaG1WuPnvaGf+vG3ZMwNkDIaI7DvuRX0IQ9aJujmQ63it2jnzp/m
fJp49p69kTP3Jha1CK1I/3xUnqcTqqHcMkXzrv8ChYWOMYDyQrzA80eR39yquQRgE2TeC4eqMr1R
+GQkpg7JPG+npspWlJmdV2qRVM4Gl9IpGtjVyoh+PvlWcPzsYpVsfx1sup3rtiH2qddn3nzg7tfO
YGiOie2D/NnQ6GHlnvZAqNYlcmLzUaswxhFyLWeMVZDDRWgVrDjaWSqTynNPf9xYgc9T21Yt60HY
gS+ljZuAwrBhqHLDQSnmNeIbgMnIYV/OmOBbPZ1XRklCveJa8BS3sNlpsCH7m18q8R97YitEIP/p
KYYwy6x9v85nc5j6HJiVZei8GuMqra4DplmTiVZXBKolru8E421maz4+C3EQqmaefR9t2ffS0Pfw
aeI6Qx5aFzlpRzgiIm+qtPZepu+aAgZShq2940GNzfkvszETZrukwdsPjAWE4M1zu+o5T+z5kNpV
TSkVEwCHtQo45rd3yWHB05Nna8YmEU1NnNfQrUAgQ9zone3f7hl+Yf0N0ivQkq/5hpBDaMjZ9Rjc
3m6XLjTKmnk+0HJmcNjRj6t6exVyaB38EnnJUgmnnO85IsU+FH6K0QjvaF66zXfEZ+j8E1dozghv
rTpYXIJla35fnFzw56SP3efpypkL6/R/xPpL0XCAoUZpySJ3Ld9YwVRn0iYywwps7dTyLqTcB/4l
onRl9p+a+mWahSzd8VRwzWomBK90d+f/QvD1eFazXmXrSNQCd0fl3KAAvQvj9OCncOb0EvN9qzOI
AR67AeoCpdEYurJrNdvKDZE+1KeYxmiZ1kdm1nWDsc8uDbCmo38QkYN2vNQaSSZCbY06JgmthOMS
UJkuSbs97mzb76hfTzatlaEPO3qbUYHU84gz1TH+vliCkI3C1Mo8BzClpvhP0TBBtm45Cj5q+0nn
LEZ0Z3Uq665PtbKSChnio6HuRNao2W83f5qtg+UMwv9NxNjGEs+KfYNAF/DTvh78GqofLkK29fcq
JGN9ZawoihBLKvIUuKH0Lw9W6e0S2FQny0scdx3hmkL9joxUE+6oPdlbCY3KSvofMVTjaPAykyL2
dbm9HaW8X1s24nxupIbZ/qgkyqqabkX05yQtL9q6lmZXgmgH++TweWoVuiwTfg8qqMOHNNmPxe4k
UwCAcX8zvtl30SdCZrQt74eUNNPuYaiYBtPAPTCiPghmd9uy7G1cQYljGl8garACeDAriOssKtNM
Q1e5JOq/AwXdCpkceY2RA2CUOXk6eXIhyWlaGo+nq0sjoz8Obk10da2KFKHo40wFSNIhQEnYQden
y/xGjUb6xKAk5EWhuKc71NgzhnmupO+9I5rfwCeOkwhGEStENPvD9D9iSCN+pF35wb3NIRbcFXeD
4lrj5FyiozI0eGMvXO7ySseTskW0tpttLqJ7Wo6i+NoEE0ovcP28/qEorc6bUIYe/DMwonjNdwBm
pXFEDU4NWc1hHRDvWuA/MjBgCRNOc/gb7QGGat7vrg5sIUrbrzesP1pPQDYZCiqok+Y5piQ+sqQj
Dlrll6IcgpD0FubqxWD17eSb7Cln4nLPb2pTStgE/J/O0481MjJgL3ps6peRRpjYgO6eZtVqge1S
0lVvS9LhsPMaLFwQCS09r7BdO2wveuB1wQ3mxlChoCJmk8eqYPO1FYZWDg+2NRBuDN/lbalL0YAX
oVsnY3Xa1m+iOeE9Ozx1tgpPRGVBgfB40C3I4OKbfHQFiK48NEW7cazCE2M21hcxrF+/LfiQzU3v
A4NaKY18v5c42NL19pIMd2IG1rfztiCidNS+IK9fZaI3bpG1KAv+thkJtsaUINp+PMvIflwHib/J
CHJj/0uW4s/sGqvPWh0rsYRX/mqB4kuB2YfSzHiHYOC05fM40Q8jdkFIyXaR/YeWWx2j01ExJStV
DC5uyGu8MRzoUdJ3po1H7NTBnXlzEbhHoHc0TdTgsICXFMhiVOkqBTZT80RNTnjLyA5oXL5u9B4N
5EyHSl6GtdP5fDSqkm2ha6rEuiwPsK23Bw7tHesMd7GolxOsFym6OqYyPRdle0gXGXlEEfO2V9+V
ad8e5K9fckZOCdPy3cWr0P98zonuHrM1fNuwZ3C0Cvyo64wRs6AuA3/zcVoPac+2Ki1WyUFp17/c
+t3qWeuok9tzCmCmy0/0j9bf1+EC7EJ8QCceQku1HnRwhmtOpoOL9yXLoplXPbpbxmP+6nANw8aN
ADPH7nIgpjljqhzDn0FBIpkaS5ytFFQYB1Il4F7Jqjh5kGC3AZD8/vvrcfp4iB84pVljBVzwljfR
iTks7RkmgUochVEYothCZHTYCErM45gTqQYG01uKFkPsY4XazDJgPZkDuhDGB9bkCsnHbZdTnUJM
BlaY2srV6XCjQhCFVViPSVbDVyaFXn6Xg/4KiYmKvrjWNlWcWZYVxdKCINWAl+sefGrze/DbHREb
2riI/ja2SeIRI/ck/wiYQud5l16U+zhIIIMb0O/nxfbGoFXo9U5ceOtQp2SDUhQDLU7Um2lNrpwP
lm0bWx2SmWM7l5Ew8HLtXu9peMsoZ8uIxiZKwpW2JZICqN5VWibx0zf8lLcm/Ey+4GjeyvlNWbBy
shGQVFYszKoZYapqG/JhbSh8pe4hboTJUTmv4HVRRdmVQbctmJFbvmARz9lKkxvrC723vL11uM0T
1v7DGZ894PznG1ITwNV8IDXDPZLxDJv/lwDXISIv1Dav24dTp7/OgGhdSUZJ1hQtFVhOg3gZ962o
CHgODCqXdvmDSZ0JbrxyMbTTPJm6+H3XrbdkBJniZGVtkfvRvEG8kJrGQh4yPPV9ACMLjY6oCLFD
sYVu5enaa36VTmTGD6aKvqBOk4+6y420OKpuxvv810GYMkWlOSN1j68PA6EECnIyuuN+6tNfTryR
dxGnM9p29gFjq/8iHSQEjNBWyQalmeZNMjopjGcPnyRxry/Ztu0cCeHDE62C9MiUU52PhcBuzIF7
U6Ftvn0M1P6ctGlOlMakByAeol5cyYGoR4/Ao7MP292mu0kx4GX5QVHMn2DhotOMAh0Wxx1DskLA
mJEKvZVCS3umd6mKLMAaSk4RhXzP2hjAzCejx1mPfZncHpdSEA9iXPpMoj2W3pV2cPmNkTm1BYh3
aIUiQl5GE8nROfPnu9/ppWtKryLvn2apziQFxTnO5UKv2xr4Ug9mMqALn088rTrkaKcDWnLiFa7U
Qbn3NOn3sfX8whgO0n3ZSjkBzOeS5ZAF4Iy6RxanzwX/zA3wdDhQvKdbhtc/LPBOp1c8OwvFu9Fb
tX6WE6eZM82n4KmbI+eT/UtxImronD1rSjg+r/eQ3swxY66dyIaWqFcx0J/GlZZX2BmrjNqbvYNP
luWcCQCmqCLfh0yUMjaKxo2tFyKTlzi87GEF1skUy+IO3aGpRDyPunKcR19jhCBC5tRm/RL1zaZS
zNURweZkkxSdwpDbU7kNCG2jPlsBHsVxBEN1FmxtSWGb07iD7wwrEeTbSsurg6NAYF1rgUJrx6pk
N2HDX//4aPGI7cTAv1SxJ6pZ9wQt/H7OenwVUGwSXLsykDRwFAtB04SvT8rijLfQRDTSl6bjnWY3
h0ViYRAvV1l1qsVPK6Hn8l+Oo7DxgthmDisojBwsj3G15SfswjYvwWkPRqKjFl63gcOqiq9mDiAa
SJS6YYlttHZUqPkYErc7sgcsV+YZ7Tk5mxKrIACV/w+mTF20pvNCsCQSnrWQyKWoR0Lq6bvTQs+D
WfyncH3dXA8pXcy3hNMc4uYEMv6JVJcf435oWymlHSrmju7bdYAJMm4sPsqFxNRFZtpgBHyNbBpD
y90anDc1oTMhJz58N8Eguug0uEWwCU7edEwyQWfP7x2wCYdIwaPL7v+sQe8Ro53lx/SJiX88uXPF
k54zMnGWxB3lql4ryuwNod+M07gNmmTdulf75kmkbFECoe6TYGuHGSQWI3t9WrPhY9Kcdzcn7P2F
c61fwqgiVqpNh43s9sxJVIu1HfsrjEQSwIwV0JHIYuFa35F6Ovomt+WwWnHPykpfonJURIMIg+cO
UzvWA1lJIeFxQn6ozDpa8I03rKhZsYqMKPL2ppsRZ1naYKc6yaUCcBmka0iFVCq0e5ynn/sE+CiW
qVwH/AFuPBo8zG1dVUdbj64CNyZ8mMlLQkG5ddtNwn/tQqj6/165YJypL8VxkbJ9QNI/NTTC77uZ
N9yB0MwpIYt1iyD3NGbgMcRQUf8kTCsGLbRrZUH+TBDXbFS5djTOINJwqtMWfChq3Qj+Z7Y1sgXJ
DCtbKKPudTMBgnXbg6es2j4/Bj0JEVfwHzeBP9tEJ8D9d0ABc1KcLYEuHcVo25vcuESHWXAfDSmA
2XKXV9vdPHFCusaA4QcmqSWoHEu6SGVKnaqqlh2hgDxCrVg85UJCN6fkYxXuKxnWkTeUg1zJbX9s
Aku0vzM5A5jVY8FmE4U24cyk50LVFocwS6QTb2ilv8YeHjHkl8oXCuYTqPlSYz2HjtjeV3Edvjnt
P1oe9u/yKX5weCH7hBP9ZnNKYoCXoGgnMS4/HqO8aOH5rsQ5wtLxE3PvHq4LfZ1YRDVjUz8jwW4R
izoZf7gSU1p45X98GR6Xl1A8zfG5Pl0lsCB7IcGrOyMyUUg/YOAfatx7q9XjBt6eCKG/FQm1vUEr
578zEpbX0eI/rRIf1fNiKyJy1RAGZmbjmx97TOYXKkCAj3D1czMJwenaXN87QsNLluel/LHVFXyj
yGhAonbJNaimARVR9kqfWjUHQzAbJf9r5cyleLAUVBNBEwyk9Peszf5kt6lblWIyTrtWApSwfV9b
6jHF+5rfB4dpxbtqP8Qa6PKi7N4byLG/+pcspdgZ9h8Zwz//bu7uQFcQb1FvTAhBmS4dSMJcVERD
+ULohvLMrhDrbieFQYtjWzzTl6BGNss2XlN/eTqHafLrulrwwAQqfHf1ZNDJd6wgpk2u5+KwSxZZ
212+x9g9R/al8PJzT03USyn32/rR/IpZWoJ8zAC08aAMgbl1b6/oHrB8nHKRCyTMn5CB9ZgubT42
ZHtEBHYHa2vjXIgEPmlsABwVI6HJS90mKK56Eni0AlawkIKQaGOK0o11Ofpx38L1q6yd5b7Rhr9I
OE7poUc1rb7/eg/gmmJwm+BJpm7saKH1nFjxBPMAyUEqQ35CdsNOwNOm4GFQBhVjFwL+1MO2eqZN
3tTSAM3XziC/fTEsQDJuONUkAheTcyIwIAKKCXAS11sVC9XDKUz2psxp2Stii3usebQvnxJVVZjX
DFZfapcTZtfIawdisEJDxeWHR6Or2dajDmyzHBFyDlWGPT0rjw5ysOJI3Nwdosy0xX8Sg/IKNRcz
AKmp0YlWR9MQcbEWjqFig8ELIdTZVTzwaYKJflgHsZ/GxOq0mXNFjgNbEbBy35zVpoQngqxbrHVY
eGklqdTsO/CmMTX9vl8/UJsne5HqiDMwzRHLp1OHzbaIQFkljai3QYvKclSgylwYRWNm+mA7HGkF
DaYRp7LX5sgwMwHQkyE2rwhoqemkycPO+o97zHVXLJnKmZTdOxXmk0EqEitJivz4FfFMMElAm7l5
V5sTrrd9o2QFXaDl2TLSF+R83KIMZ6ASee7hTQnaiTJoZYQIy8t5y4x3sHFs15AyYTu4S33o4wKF
sI+Z70X1sOjM+FEp0g8mPnnPGaKLGA9UfkKyFxVBI/gvL5Pcxa4MOGBga42EiDbeo/2zMm5fRhNJ
Rf74ua1kYhYPtc3TO1WurBthd0RObcXn3PORpiRbALICzI4gn/viNNVoN5u7/5v6XtViQbsJnsAY
r/xFIfABo7z/VsNvyBKhZ2uQJReke2i7p3/5CY87NvtevGNCClGcUxdZZeNAXH55XhfqHtUF2yD7
5P/SLG9ECEd14EPA6fuVUeha24DUlmIhr4UzdbKQO/TmvozjZYR8ZiAUtVIFsEAalsf9H2/A958f
1lavFEkHTvu3gMV8ZMhXh1l4C+Z2Huq99gg6D3um08lfm9L7y/Z8VRis4Z20mjPYT6gyu95CaaiR
XUtjKS7mRDOI9XaVa0D8xC/i5q9d2jsqgOx+pS0EAlPz3uS25OOb3oQBCQjnk5xixjEjyX2QshMl
L+4SB9RTOuDO4h4M2gVmuK9pI+xyONwLNdc5QujiShMpkTo0hVeoQ3frzbkvm9IR4E9pJeG6QaQI
gt2BUqmZcSFqUaQzSN6aByYHmJhEl/qeoqKUh7n++o14MwZPjsGo8nF3HhJwUfVmG2dTEfS0DvUj
4+zcS5ud3UixBjBuAwOdlWW/OideedgeNyDuNlg4Rnp+EYIKslvQ+sgdv9I6IE8pcaJ/LTTJGl7n
WzSIsVpCvUi2aKIDfiXO93IHxDlQi59eHtnTbCDqIM78ZHUc1TfnLqhu8kYMI08sq4zxLvXCj42Q
fOS0Z4Fdmk+bSgejymNnB26PKbvi0dkmRJZgiyKjMt0RBNi2NFdQY+CVbo0OxmmfuiiebhZFQyVv
+ZKEA4mH/Hfzk7gk5TuZPQ2IS0nIHOgATeVSsk2Lp5RPRq+56Tz2ef8NsG4IKW1rMTe9PlHHbu8G
2lwCTbm3cZO4xG6X8SQMJiMydnrVfg952+TeTyXkji49i+SrsEgtfAg3NPJp5LxGaxJNK8YTeIrw
IpzbEPP9bu6a8cvFNrM1bEfwDotQhTS6yObwYcIkAcETvhJxkQEnDXjJ4gmUj2T5sltk8eA/tSCb
pRdUgtBqNqNb7lv844UImiRd3aMaajt3WhpPbj5vMCPseRNXKGgWPNQ9+H700AcoXOSOZlWQ9V+H
rL719L+OHIrPz7M0aO7mVcURKM1/U1FSDmhcB/TKPIRN/+a5a3djfz6pWeRKzq3fbG5WLaVDY5cy
0dVK5q2Dpb7ZrGCxvsoN+HQ8hNiJHj5JzGDv4C62mges/Vbyx6sNDPNs5oEe/iEe1/oCMsJwWIKU
VOOixLBzlwCljxZmsw/flrEwDL6WTGsO82fIe4IKkhQoK6X1L08+yar6d8pC9iGhlELPT60vUzym
33rwJ5JyGJWz3ozxcTKGaIn+LfgfDPy14xJQM96kh1STLcbqOvAUqLsmd6PzEGp/oenWpvNMewbk
hVeJs0LhYKu2vjBgstRsp8AHbwWHh72n/N4nMfZoMrkEKiFL1aykSiJ7Lxkq9dW/9p1SKM79WQBf
NyzPfI6bv/Ly7Y2M/pOQI/T1jFMGnEZD44nPOxXKFMW8lIqdIL9nVCGIcxk8Pn+jqILjy0ff53hs
fFGJ7sVIVCNs4Fx7C+uNpb5BQIOPIYHZQMC+l11CAB2e2WqK4YmwU1wLCv1g8by0WvfQ/Dn200W2
sMhmhw3Ktuy4LsMzELy3qAAez2JuQeHyKXRkrb+91MxfkFZIen0GTfOCVIwxDLgq0xKuo63+Tv70
bhVp87jAlmnkNYrXuTpZmEqMzAKmB4qsnZNOoVGMg9O9DbXHuZ0e/rGB6YRM/5SFGudPmkAYgEu3
8/JtPHRGnBiZEEpf83DNcXvRIMCRTAHnxG4Qi6T5NwbJYG9cQuz1JVLkcuddad/y9z8H+W2BjtHm
s57LC6Qj/0f4Xd5BSUxRmYpuy1D41+kKDgoE36L/gJ1XgGbDigeQn5prR3y26REFHbD0vMM4I5Zp
Y2lzTAK/L7qYklwjhl7gXdklJBhVavUVwCjXgtzU8UAJLDge4XnPx7yXLb2MWAcHJPs6K+NeTbaR
sWGPCoZvSMp3L++m18CIWarpDtvkP3zS74zUmqaUbAIQO6uxvjQWMFamLmCt0EZ9tJO6DBlkvrpg
RH5Qw43QxLbY0uoRqWqChEeYAHViXJfg1IkRi94xtr8/OjiA1oEhZ/1yb2CAqDzfW2WSOvLTjwt0
4H76gxsfmiriaZ11OYDP7qr1bkz0rPDa8c6Aj/XkTfQFzlDB2X6pfdN9olRFq+QgxdRg5iDp3Eda
kF0AKdnIKmNCk1U9CSeTv4liavAso1kXSwI5G33ArmMCWQC3uotIkbdR45uya5vFkbWFqBj4/WEX
s926nT7FlIoZiS+wMgJ+fnIW9cPtVUzKolZPsUVR5ibr13QvJXOPOZdckCQIhUyDCH+GsRgC6+et
kx43KD8hr3mVc1ZrVsWQQ7ZeBb/15KoLbq7trIzR3sNX0g3XjGIPo3O/zRv3TxSPXSf0L63mJq/I
VPeaf10Kiv1mC7rgxbcTC9IxbqaDJQZrWUvVJqdgc2Ow/PjyCBBgA22eL2k3kTcf9SIQX8f76nSz
70M0XtTBGqNV0x4XqNUcNnplDUCg+PR2kMPadakiPxfn8+c3IgJOtKi0h42DRmMm8WUwcDNGyLB6
MtlFLwY/glJrc0Kp5w7+hQEA7nk0CznDUy+LjS7MF9DfKiMEeo91Swz59VHdMeWAng6SBxx8Iq10
93L3vuhK3DYWvd8I4GTQQcfsIF6NlV9+bNIVcTQ5EcZTVvTX+vqs9SjM+2hH2gnK1W48LcuQ2qY5
M395YU9847V8lcCSwIIANfKOkGxQJgbaB5at+da8V6I0/6OT3+suS3RTgz12eMbUNxpT+xlqXUBM
kGCzDMSASPXSSjhX+k32UsQlMly3rJ867Ta/oCJtpL5it6DKkojBGCJUZzhl4gC5Dg8hV1YYhuh/
GzzVPrZP6POazJ36QBv+CVfTXdgOUYpRG7k1fKWvUMS3TLJNswhj31VP99y4SlhEhtZjooPAVB4s
5PQxu6Q7t5wEtNERoP2oOgzBfVujj6l2gjEy2W0/f7CnFE7DpBt8v0/Gfr/jYIqEERBjanedeNCe
VLHdUY2vLE/6JZ59T5jz0KuhiVUrKSlxSukTQlosgth6aALOB6t1qYAXgldAjQwE3/y7lBnqy5iJ
K7/Th1BS3Sge4hX8uztI+T/VqO+N4h7b7iuC0gx/NN0Wc9pStUBHf9NaOpDHq2kCiVI74PEhyyuq
o5sKvuXiN/1z3/v+GQh38PAj4tuY5lHD2B6nRjHwRStuXLfKwN8YpQHKZGp112RidtLSvR4TsRtN
eKa7vnnN3zU2hD9wdt4xyvcA7XehvHFWq1qCkBnCLdubJ81jKZGsPDNKMnz7d2ITANr+JkGCrt57
TerVQ2oYQ603w5ivFMeUyoeURIDUV1CYpEMl/pPoLoO7MQgrATxTZiBe9HhVJBoWeaSsK2tiAjSY
iTNlmhrCwKnEIYHm2Kb6otuKJ7n3knLaXJMkh0XJQVOmETme7td2uQOMdC2kpx0eUTqB/s3+SsjR
AIji9JrBZtqZ+5zqLeAF94pcHlUN0TlhDko0c0FoO0/08RTJp8yAxTjLYWuRUDKBBPVzpmVmL94M
DSBq/TFcisch1rNVfJYk8WOCVTeG2KxMTGHdjkY36tNrl45SmyzFl3R+tI+s//lkR8HGFzDuvmmB
DY2Zk/EI4sswPYFsJqPGkenqYZ1PdMsBsZufqof0PcMQiMNV4iUHoASGSb9hrNIVc1NHrtS9MBP8
cMGikyjL8nJsB9I2V0VEwoEidnNsi0tCYVmvBMf/X8I/PmHSciaSAnWPuWCri2JYqeepNVdYTAmU
YIKwWBBkk/Eryk0LrQZB7md1L1vwPZNhImOf8k2Snm6/LXJ6CdfhIydoqB4Z0aKMVMRk9FqlDtoi
1wbiWTDrTCPGqy119D7+qZjkxESQ67g7piy530H72XtbhunvVJNBCykE6XJkam5+xbZSG2PfCyCl
nJ/gaemoXYt/SYR7FjP5rexFaB9SbqMDAJstNDWz5HY/I+3QRe3cnAfLwy+PqUUtiI7+mFM7Levs
vRBt/Xx+DxBxT3iLtv+RruseJN49TrsSnykflAY9rvk+rv1I5W9+T5pyxvJPZoDHrWy2uEC6qt0I
XAQfbcq8XSGF/mGEYDoW/whvIX8JCxXac9ImluqbuHkg7+WJnKhsyG2dxuITHt+MWkjtqYfF6grW
5WWqOOkNoYiRmkm/hDzTFjuAsXDsniuROuRvmUUZb+wjlgaIgD3z5rW9wgOralHoAy49WH3oYpzh
+U4iHBYGcpiUXBm6a/wfH1LeDWnGpH9B6sR0bH4y6WvqgLbvJdxGrSy0bi3+n51TSIwqQlpfT7B4
QXexVq2Sq9CTQLCw+fzVEJwAcCjEBDZh4XUlKh+/r2JQZ9mLJzkZ02zdSql0hQ+6o3+8OiFrUDdL
9AS6iSVg++8JdJCTfkO6gb/79BLXrNukC1awnP9mLoPN2eDPho/gO0pfTjb/7SDNV8k11xz6uQiv
KALhPHOGoGF4+OO5t9Fsr+y0zA0wyZ+62jmlAxPXGEVDOd/0H/ECrHN3hat366ztkB+6viREFLIF
x/olEts0/ZGISdBXYeId/7RQH2dEUEyZUUCX8dRZIVKunYRH10nOcocmaIUVrtiteTi1IJ0lQX9K
QhE9HN6m4GHrjRjo4DkIpNV8QIQLXEfchgE+VJCKDDTm4gM8UxNsWvyssQiVSR5YgOEnETCmTj2k
XAGmVAJup0UIfQldDKd0hRoA1rqtMc+CZD1xsGdq9+iOm7AcpBnVrp7QfEBJ1ukki5bQ5Yv9gKiQ
5Ewgjp/ZjDvJEY+Z9DyrPWjPXqkXLsAjarI6Lq9RVAtUf4FQzQYei3R3y74oUCxIdxkaUwyDUZ/k
s8+zh0/zS5nUskk8dJ77A3AVaKD/Zth0p6TVhctjz4SVGUUbPM69GQfPr2AsZw4FSxXQxLmOoD5S
FpGnTAvmZTlPHlF6C4Q8GN9xN2R5kN2X11w9inop8QDA/KDjlOTkXpEVx9qVGi/iFcm9M2jWa73a
vn6siFlH2PNF6GtSf43yS/yTIMcIU35B3YEOdzA6ZGp16EkFkEo1ek5imCSEjPcZ5ZC/LBtuXOZU
DeXgiKLdPMiHL0DMVNut8Q4QI9grugtHIPjcnvK+4G4I5hXL4IJashJWykUEnEGd1NLvfY3T608k
FfId1H20pao3/RH+tABwmQMrZdGK0nzUiwhF6zwhZluG1wqUdn+oHGszNfEBJaQJIpwRIZ1TrOq6
FK44TcJfJob5ovAvGd5Zk5ia8zmKvYqUBvH36QG/TXfeVWtT/EYZfXmroJLJNzUBWulAAMLuH5Ak
tzk65at0XhDExMgwO0BYwa71E4RDyEHN1ZK2V/70sTNK2qJdqUvUKgTF8dnHzVfJoY1bzk7HupDo
xPhOJ934dpJrDsSCTygI0Q0NuiWfrBuSyD9nYdvpVqkdnxjifu2lLn4JT2tIjwZ4mHj4Xmt+eb/K
NwcbxrQfgs/0NlVj1sqOaai4pP0xRk0kFYtR9B7+Fiocs/xGm6je/jZOezfzvLaNOAQ0sKJpAB8c
Z0fsWA0rcev+rJR+3I1K3gdfB7YUuuVd/xn3DCz+h3JafezwEBFYCGQdpw7jaQRMGCiLLKbQtb/V
DPHRIeC4jtV6+KtJ+OOZJN3/H9u+pAK841hzHW7eCjmEOwMe9Lw81Jp2fCV17ICy4xu2EfAcF5Zg
o9Ovs9tRYuoBdKaUbCfKJQpgqyo0IE9nMbQ9ziq1zOW7sJVeyjaryXxG397qkE6lARhHsPZBRS9B
X4J3C6GHPc5Lh6lp9MxXJfnEsOLZ8i0AS8fb592qgtD8o0uZWl049I685ul5AxqZwRBFivKPsEej
3YbeK4kDkzKPjCHWQINCN4adJW11OYQc8rwePiQumxgE0Q93AitfdJTRIlZ20nduuhdn3Mu6CYwW
kZTAIt9x0YXkT4B2pNN1Us0o2Wq/3FJ37Mrb35HGev1AdDx8viO685jBhBoqg/eyF7zZ+qNVpnxH
9YUk0i+PcsnmIA2NfkdkY+6WrWyni6oPY642YXjKowTQuoP+3JT7hUhZ/bJG4P4iN8ZHYwBqJzrD
1U8SU1pgZ/hDkIPIvSZ7qNmCMj62sSxxXBMPyA8QSjiAVyww8AFlnGoxzgioxL9aI/hzY3Qej4aY
TQuFOO9+Vtsn37iua/1UrOXbpgS2Acm+0jy/+q+JuNs5Ya6R4Auc6Nt1WrQneqykM84CfOcXIMIO
KCNaG9TE38y8NC6Mf8qTHwIqbu4QIqdXQB2txE4TnkvLb/SgTcnHvRSG5CYME+NfsxRy5p3FEYml
lL6knfJHL1ht/12DJ1Me3w11gDRtp/GOtawVad8Y28uTo7IrhONJVZEVAWAUfcbkwJ0aLnI+hA/O
SraAZVHKdI8hgQCZaTKyd08BozSKu0Z9XeDvz5m5B0xphgD/QGgFLSCJzOGtfJRrrEHGMnQFIZYc
BtchVLOHbJJrRvYCkhI6ojq9OulHjXvI4/eRCQIb4IDk8pCuK0JhCr4Xyp/jwDoBqe/vLrgsqiP7
Hg+a3SnMqy0WC66BU0W6f1bP3FfDJeIyC7NzbjEJzt6qYySxaAMUy6oS8yEoa9LfG/3jHd0Pi3cc
OxLf/il2MDnjA69gWAMu8NI9ArmjdPGp+J6awO5fT/ZeImRH83P6R7wDH4xsT1/di/EuIYIBYqpi
oGPtA0vWDUv1BXAWGGv2GMKEpzcGYgQBvD6gBBTZSupAJEAmLUcjE0/dUzT72reB4yHODOv++pxN
ywC/REFEOluFftd9fLH6mlyzvf1Z/Q0Pu/hTSvHhfSvszaZbIMAalBc0Z5+9ioV2SLKy5c7ST4s3
VLQ5dw5YBs8akm5VThS2qzlqbqGvqK98UvVVjEd4mtQY8J4BDRxOwzC1mB2pMh0Cn8JjJSxzxCJz
RADs0Zl5MM6KMjpMlClMD19ri5xA9Z7g1wt4dd9TZE86q4DvyiSctpVrSvD+vP6uiERNJO3pVFPb
4P649w8gujUvMWAZD0K5lTMbzx+UA5xuIKbj4xZqjWhfdTNsNV8EaNJskGizkZpfWVnSKiJ56PiR
KtjIYYCbVhTGJQzOQdGJgOAUgxHlNVSFD54NzRZoQYATOkyG0ieIPipcMpg0+y1e0KteXuPR9GK0
xdq9H0ze3LO3PboAvpNTgod5qIZGGDtboorR0CQEJWZLSyt1gOB+tLM/IA4SS7q0+EqY9KKyoUt2
ZO2g5Jp5irFKS0IcLZpfDMSUPTOiKQFB326wSbiNdpV7MLth4IVc8mHb2/hG+rXiGQN79fm/Gojc
MRvOpivyStT6UTLXxsn9YPDEnPlSxT4nI/caPgApQQm1pKe7e0MyOlHEgz0Jal2lLS/AJpEAzxCD
Pp+AA4t9BHQ1gpSkkxjBedSjdv3c+NwrjwMA33nLz5Mok2aQH5yr5xJ9fv4OTyYYvus4a5C57xsj
6k44Spd5Fe8VNepChSj7LjmPNOazbwYy12ayvNySMfGXN67hNkP/ZHTEmFa4Mx+wPvLX4FLVSCAi
wulAscEjyYwOQjf3XWfCafgKHEPSySQxAOUVI2HNMm9w4Emuls2QxrhsC4ThMdKp/vRJFqasGRFL
Gj0XSukLalkRdmipKcVZr/ueCXgjDZjyXzK+TpCsOj04lmnmow5szj3HugP66YvTrbpx6jxWb2HM
IaEfQ9DpNFmY3j+hgdbDEo7iVgdqVv+uv5HHMfLGn01O78AvjTosAehsFrMSMTPUeihbJI+YvVrt
G42dtPhwBrywYwmKJGmq2FtJIEksr+XiNVTmJrAxTUbcdEKgwtkVJwlM4PcZmvlA2n78pWiWnslD
5+EUXkuIiN8pfl2g9zfrS2YAKGVCsZ2mi49HlzbDYg/d9M3v9UtqYpYr/ceuUL7tUvk+CbAlNasf
vw3eML2CtoVZmRsiAvIMOs3oT7zTkVoEMYs8fZ5TUbsuVMABxnJgB5z70Nm3Q2IbNol7x0IjcnKZ
KMwnvAEZysn6P16acB3w9GhV8MCHBQ0rHqhtF0kF8Oj1wf3QtsgwVsUCIC/aSr0nuQdgLWTUO56Q
WRas2Vq0gfnl2mHBW3sQPKmPIFdT+hyAsznO2mUfscM6vlv6VvStGLMh02+aggP3WEdhz2ZtbfFv
a5OEnLOauky3g29c/Cd1S8y6zCiVUWyXf5pvijn69ntBfOYho2VdGhyAK9ASnSQ0dHqO8Nf50agK
CJxY/kHOg86RKKbhHwnFEvKGBsnQwITWCS5Q+/Z8LQQ9LbQSjavtfbk9WWFQ79aeCA6H8o56GZ+M
wgZhHAIDR7Q/Ig8ocHjDFoHk5p/HimITGDTfQrdO+3ORGyf9zuWCDDKoemH+sgmjklI1teQIbuNm
efs6ZAhttwcI2+CPQN5X28uVKn0T8p6v0POtMdAdgySmiVMNU4ZSr4iumQCBqWa/XAeroT32zPOJ
t2b0T//Q+N4ycQJdTsjk/B2AIfIypnHn/Tbv8flRwH1BNe1Yp1woJjEIZCo5Dzz8PGQyjoQ9o+zN
YN+/z2Zj4suK9XjyP0pgdXUg8V4kKiUYnbhTz/yRFPenF8A3U2Jw24BNGCu9VV2DSg1XWt9khSsY
of5NUElgUhknDtwOdsaY6VXVVEobNtlCmr1I5jgo1Wun9T8UuAYhwZggFmNF2J20PzWXBP5d0nRs
l6Dm63UZtdYdCMpDgrSkewsmb8U7ztH7V3UJIQhxFwFxoI1h7JxMwytgCvnzkFHfBd7ZhM/2lymt
WjZLK7W9fnl9YOn7P47N0EtvVszFZYic8SjO8hrjsjXQ/m6i6AA4cFJDT8xWJ6cIEyiVBrFcFzYd
s5hv0MzT1YyOTPvHHmlXy0UxOdrxNa2jF7EEQ8CYh6qB9yQGwR8uoKSpXC4MXO9KbWm6rkHGG7UQ
RuoCUmxnA20BfS3oOqmqhYqwrjphF9klv+QfIPRMc52hAu5wX2ddvQGq53Bk7sE9DjdHtaUjmvoF
VGDE1s4bZW5K6uxheGnnc4r5UIPjgkP3bWeQYp3FXLxM5ery7ZrUlDTK+96LNIxPNPr93u2DcGe5
UfHr7J3I4cg7XQ74ia+9tJmXCu/1YN9bSTGuIaLdrgZ7GU6C5/m23O5t0YQxBDCXSJovGGgZyj5E
eGS7rUwzFB+DEa2uhNvc1OB3htzqyaYjulGVKUcUkV5mYuXPzdIIaZrOBrk8IvE94sbhti0bQ/jH
LbJoAcqOuvc/qSbqMtTlXYk1IH9vdmvMB6FAlNMy2MRJzSK96qQfPIysbc+1qRuF2wQjmKaPW5Gk
hcogdKSCxhl063K3pv2nMMgeF5JT03nvEunf0g3g5FtPtc6TvfLEY5ZUt7XBvfQhIg48XQJEe24+
h2ScB/a6vHeaT6+veZ3FH9x063QVDcnLnsUCcQuhhDvm/OFxz2kNkPLntaBq271qZvluraa4ONdq
2QGV8rGYwc2K7SrmeSFzUOnfYz0S+usOPdnjQCn08FtXBceM34w1tvZ81+k9Fd7nhDxS6dsuYCXL
8WPGUaHDTBo5FGLMX6SYO0HWisgbMKc/2nWoOstb125TvRhAk5c/OqxnqDhjhM4nT8b62wfDw8o4
x9nVLOarkcyABAhkY6x+f6SmeS4u6KaYETmEF253N+4NWuJZyHyPCrM9nf1GigdN6jzTi0cP3SwT
PpXDNM9m3MrXQoC3GDyOSimRvB02vZS4LRpLhxXRQk9I8YThUw917ENbHCNDrTUG86mH8fP7u1Xs
NiwMbFmVOqitxpDaAnblt8wmLhTFfINxoLkIp/SEhotWstyDbFrbO1ErkNztroXJPRew3VwSH8Z1
bW4+ewhqbEQyjvFfsrxSQ/8QYklxqNpKX//PqhVYvMwYT2vonaQV4D1yV30+NUPAvC+u508rxT0G
03ituSn0IEKNgsrz/GjCBjGmbWT8vE8SBiLBdBOJ6uOYHOZNRZnzd+/uDj4/Ht77ygE0i3gFcCvB
NjysERUQs9SEHGtlpcsQR/tgYK476stlPKPxNKUNj3QQiXL2YPMWLUyDD1a/Ug3c6l5chZoKlwgL
+xILMjySaTZhYWCW4C7svnB7JB5LURK8Y/h1QgOvrDEZCbARvU20fO+yOidICtgS/Z9wjo61hGmN
23eycXOaX5Ng/N3NhrWepWkOCppNax7F6XRXkPc737X8mgDgRIc0uhv/Y+6fvC8j7BDcl69zC/sb
Qg7KzfUrJCqOukT0upovAF1VrHJe0AyEmmfbYMorLEIvjXKDKaajnJYdQ2OhNp0vi/JrpCvs4gn9
u7yfdjGWC3bdWTfmKSedtQGH0DRSv3FokGm5mZ/4ltHKinm1Jm0GsXOcNbrv1u2kJbfLv3LsTeqz
r5j/xgug4k2b0QJkOOqs4yTvqncBNT6L0qkjwfUtzq4zpHFfEqUEdu0bMuuBDmflIlGnFMmzLEUY
3uR/M86SQnioUCetWX7ZRSFjCfsjA6GIkpnljgjHeGW+QGXTMrKKNdRGaOu47mPlJm+huQmM3Z0u
+55k6cTQTWsNb6Cb5plLYTuT/00PYLH/x7gBMv0Y4YFqZ/PdTsVQmubfSQ1nZ6r3Pfa03/A55bxw
+jQFtArOvJrlOoG/VrVAO4FcdNoPSg9nZ33lBK6+z0FnW8lTgcqoEmD+l+JqVpHKr4KttQF3p8p6
ynh6OSfLm7rJSwn/zMuls5boFHA8uWcWnvTAnlZL9bvxm5zZ9x2s4yTB5QVSBLR8D4qYzpCQGSC9
L0CW9AEUxjoKZdRdrCEjwtzw8Ds0sCgeouzFO0wwKLPR7noeNmnnOghL1dRxRxgqUTwBzAZ4FXFL
dilvXPije0wHs6fX31DANOSZpUua5yD2Kklr1683/K+sWRd+DR/gyzSdlmhMXXJe28n5O+lVicwA
yR40fVO0XbPMt21LMaAvyEoyryVTVyA5351GBV9NHv+JsR4KpcmNf2Ax9QDkJkOY/adAbCWPtoh3
jgc7oSryUOQqLkabSPZrY7cCJ6iLC1e71AwarWdcrgaKnSYuG0aZOIWFMC95RbeQBM1WrZawHItM
T0O//fEF1L75FTzBqBvkum1fO4MzPY7f0JBWIfL0G0d4+Abz2BuD/2trtieSvsUUByfVmhYATcD9
+VHTPVcWcP8dAco87ihDFBccrw0troRFyeCG2a9Tx7dEUWO6/7yGOyAaMh/kdTYvzjQA2SQtZoJ1
RqNXl7YyHCEYEmYmxH+KYRRovIdVccLBLn1ZpJCjLtO7vafxMLUjpf67qD8Mjc0BxGLmysIbL24m
sY5j4go5TrcKd58u2oyeW+SO7YpWBdup1ai++V82cnfYELJ8BZ4AF+OtyDrLF6k9iy7mh3mHa3q/
xE6fXuRXhc1GUbmeUTlyRwyQY37F4VL5kQOKdlqTnaNEfnm5DdCrqWcim2JekyBUIwqMp1QXkDho
t7kdXnvFT5aLD17uD0jQOa7BOHkGdbvTjRP4ROzBIt0of4/AylRyBCMHbcg6k4ReyIWZU1r76pkx
PMel5VpVYoHIMhhTPpFAG78rnEddFdYLvYdBTpAx6gYMoGA0yNkuayWeVVDk58nf4HUXCjZLhwVl
VtF77MchyjO4vDHnvk6FEKLDAfofEfPq+72kmxrN9jVvxjm1LFBKanwYmqQEBXGKAg7ee2U8II+J
K63xxo0SI3AbsNiENB5GwnD9j6E4PQuT+qajqWAcJM60zFfWcTDjE5zsstv85+befRaD7iaIcQJe
S24kMK+Ps4XDF7nOhej5VuQObNL1xqsPQB6Vj2GRcQ+zANDBR233bhg6TV+ZxO1/QtMb+YW+Erie
RytsS+DWopLymLkPfrLDirEtgCWXm3QaXFRQDb3v7CCvynB69M2SgIR4f1BcJaandP6w1i9iobkG
PHF9UaTGVwgbhFncnwmrC/RrBEreE7G57lyxEZicS9NNkNOGx5ifwL5ZMOGwf2BQy+WYaAMXQNby
liK+d2wjmxlOSsSUen+2v0Y43ta2jbCCUPO9dnA1Wz6pDf8XpyyMEeXEElFn/9e9YSDD9O7KcGL+
kPWaA4thwQuEdFe+iM7sENunLwXkibXuf5xU+yFFD15iWtyYauFwEeDvLhu26hi1p+bwd1ISpckG
zu/g9RSSbrnsRFzyIa5owz8Ha8oBQh3PWCUDmHkAKHIFwqiASythaRde52buBjL1QOCBdnXaFs6Q
Cf4DPcCPYR3LP2yJnz5uRSj3PFAfFHadbCIZ8jJKxU85/WVdTVodIt0/l/EN8tcQHQY1GXG5cskH
ADcr6gx6Z4G3bdEJg0Q0CphhFl5hDwaJZembQ9jWtXmGW2xLwMuYiMNIoLniBKs39xN2u147tcyO
gLIkXnMspqTna9o+tJ4exF4uiaiwpvL53erOMjSutmf/XNWOWffSWGQv3tJUswNYsLydetYwcVNh
ftytnbTnoqmjWHgmV4I1wo5QaVAVkFjBCETpz/UXKWLqe1ZUPxTh5hqeEKh0IBf8a6q9uPDkqAS+
qRcf62dA7Ldh2a4VJ08nCEbVI+MnsGaXU9+J8I8AiRAhkxyWm0twleE+rsLKDXS88SyW/Wx/F8jd
Qmqf9vEt0Q9jcrbjEJevTmYC1nUdZM5YxXOUtuRiDp9RroP0lhSq6pfMs/3/FE88LZYOSmYXTNJZ
ZgsoESXg9Okh7xEQj+QsajkHW+49OBLt55Bprd+EsFxD/Dvm40T5XAM6iU8wHWZIX9xeZSwwQkQB
IZsCgLnXXopdxzQnEC3H/UGUL1ECd6Hj7nlD740NVrcR5oRNh4g9c/VLAuTGsAfKlspEK5gLh9cS
oV0tj3Us88OO25oWnTM+NZxUhT6+unQ0BAlOKnt2TUYt6XiRrzPX34im0G8JE5/x07GR3liPYqyj
Uj9tcvbSpYppie1LghkxrCCtQ0rRoVIComxKPCrgkpKDTUZR2DbMxN4femVk6gAN5Am50IkZ+y6y
DUHeOoeNmMBodcoDstlR4q6yziDi6E7VvNpX6FFok9RHeo160YU3o8o8aIVjRfCr6ZOL6QgrBieX
IGx00uQ6yfcFExdX4Tk/B+f7ZBMGQQ+o30gm6Tqea2HPLfINszlDDafOhQfNG9vm8nPCmGWcic43
XwsN0+JMD8+GfDcMMUHY0yGBKwcVD99WPeKLDnibfYCR6cKpGwzr75AM8VW8HoS1J9Fc5s79I674
StWwpRLgd5xWdnc8pR09tcrUG+evsyBxx+Vq2gT6uO3O6yQkwjUjOkVoEqDW4rya4tu0S2Mc2z+J
1bMHSjRjWrCQWcCa+RaQ9eJLl6z+hk/ECX4QwfmQhyOOXyGQiOXYbMvrLPHba7IzXM6SxSr76nai
0BKVww+o6Fw0i5grEyUnohR0W/oz5jYYtZ/GZmXZGmL8atTVbJPTNjt71uqOKsF5mMVFlobvozSO
6sxMfcegIy18lrOioEyxUjjucg0x5SzK+yDBjYdk/sJoGGy/XQGuFwdpJnh+zgQRaTmMuGNXNc9L
lj61xYfrrRzRZmKzgetMzdng3Z+AVY0WTcmF5md9WSrUhtwU8RsBeSUslkMOkYXKeXJ9XfpDO8Ga
5I9ptUuiEN+kdSXu4EmwlbqV8gcU624sG4ekG/9w/jPdjsMlOfsXHjX2wfJBKrVLW5rknIsEGN/U
kBYoGURRTYtDH0FWLdYvwzncw+G4Lhp4N4KtD4y+YOfzfzE+xGd9rr6WRyulCAsrn0mA6varVt03
+X29le9WcUaPuw74b1r9/AP8Jn8GqJ2bWMupWUiM3GWJrACetYsfRb1HOghwdGzQS6H9AyLpedXQ
Yu4RQ9nkiclk33t73bbQAJ+yVSadCXJuNoaRBuTfqYE2LxgZLDE4ctGuSL5A6fbCTRdE7an7JW6t
f5ge6wYDqsJ0m09DizHK2kpoYhs9JGItXFjWELmGtdhpBf4trRKnfE06+zPi/VtzVYdIVPPQWZPF
KsjRIli8MJZ28nCfDj2ZKROtf1ogbjdqLVAjOGhdDj2vjrwhJFn6OWUTYrozMesx6mGL3Jd2bMU/
uuIDpvf4zedIxFm7qjzVCarVejMdJyYQK+w+e1JdLoSK3LpklK2/57/bnB8QuO7+kiq+bfh+hdga
8ZvI6I91O17qzSIM8VzX5HohDB68b2tPnnidZW61V8rk+u62mBHdL8DIHHde1Ok90j4BSXJNpJAH
bSQEgRZ/otw3+2/si234+TekNR0YFyfrpz0mD409RNIocoPOg7xFRWMxsFh6z0OITcAlqBWE9H5m
Jm3Pl8hGNmcXbZ7bthO9kDqlNoFjigKlWWk7eaGMTLz4U3mJqZSOALf3sCVpfc8UPGuKFR+FjZYp
YD/OzzpCiy/GVxxINmEIJu1NGfXxjYNg5cNz0JFNzR7QPHNbkaetP0KoGf9ouKTm5apV3HXJpEGg
zEvZEEATSGR6gJZsiXlRZknsiNlIVLOVaI4pp5H8/dcKW8d4Az8f91/S9bABHvNVP9GZ3l9vMkZk
B2FK5kgQ5U0BhYWvsTVIdmDtfmkFn3wtIqS1R1iNlsY7Ax1XsIPSGMJ3MJg5otSn6dILL0UmpTk/
PF3GIODjRfYKjTUC0HnfLx3yP5uRCrJ3/93BknA9uovwyblVPZoI6qG/tTjHSIc0ERbyn3srw3dD
Z8nYEZC7LuPAK6Q5LD6Nd85ncPgYMKTfZ9afU8ROoLZu5HP2kUjQBz02vRrg1zjdBFuY7mdMOqtJ
NbRoPTJNujrdkfJyY0Urvow1ydJnmzVGQRXjCsCmu1pWwAjEKwYhleKXLY619tSa8iB40s9RJ6+I
CZcCdwEuT0yW5e8MaLFJhmgsyb4T3a7ol7SdXGDfJKk8R50ecKXBKUG3oVJCinnNgVdxrXM/c5Q8
u+e9LB8y2nClFcDL3mzAaCJ16+T9SC62Itk1XrWepXgw0qu9uXoWLsP9fv/At/sAneRoowARhOJT
K9XgLQA8ImoUV/ee/QWU/OGm23OGivtkaeOWs/hoKphj+L7ooEMyUoiDArFggB9uQ6hEi1Tqh4QO
F1fpLjs1K4fnXbBdmvkF/EBopLT+lbLgVR690OBBnhJlSgmCJhcr92Xj8YreaMDCss0NPxm1EV5C
B3DbOLnffjK26bfrRWofdhQZk15+KbPHPECddK4wUWC9RBt5ILjP90xbCG0ZtKShBM47VAh3pyuI
EjnKW4Ywx6n3qOTlRTGCUgdGXZmxFReLCmSwD+Ed1Wxpd9Lv0aof3QupAosYeQgzQJREwafNflp5
lvVfWE9B1NLuB3CDQB9RN81AOa7tbRvmcvGHV/VXXt9D9SP5S7VtwLIOFhADYPRVoc+tr+TeM1Mx
JeSdloBvMJ6YFwMAXoIFz7IRQuM/abOpU3ve04LdwkZENAG9/qv/W7Nkld+WDF+hrNEkWJUI4fjw
n5BKKI0Gt0bwszRhTETHP10JYqVbjNd3TizCWr1RBVPkmYuSeGD8GGJtMKWLR/YyZDzj1t7uAVZ5
CD3hd72KyySDiFTQMk7lQs7eDilVLLZaAQSMSzqsTw6mbO5OAC2VqsxrmsHJPcdUmMqL3sK/GQLd
Uw5rPTtejkBFk0q+PsESVBF05SHL4xtzGtZX/3CcAFOYqFDAMROJ4kdf65xkILzZOeaGwIyMMjE3
OjlYfOKq2dU9OS4yJC1rBWrWq3j1pBdVm70Fuv0oUMck9EIBdlsYMN/G1FEgDxERQzskbrwm2wev
IzPXVG0B+YpFdM8YjHgW+dOl/5iBVOr5WErVteKeLglZhfwpbkcwIXmcYDv6jSjsl2+0P5hzIRpq
QyUlzehnFF+RWFoBtdm72MN4FRjjgYejrwCauiE1N1UubwWRQwrLj94okEC3887fNfRsmH9cbSRU
bGEa/pG5NRuSWQAeiEIIvnfGTgjHO5v5pJdNzKfLqSJw5kcyxu1SGOwN4g5QiPyx/5jpRZGzvQqY
QJsUrsyJxLkRjaTG5d65DgMvCzZf4uRdDxncvs0+LW7o/NNNG+JVj022biFZuT/i12MdqO4EyurY
IEz+PThgXvy+yDGL2iRF6TtnYPwpvHhmFz9GOu4Y2sBsLn1IuXm3gMjiALaHIVGkXGiMj22AqcMq
ILFOa0w/PYWQbQRasumEK7iPbkmhONgrAf2AETVRG4j42ecJ8IM1zYMEVPM87329G7jnx2rBvasZ
bamjSu1xB7kOaw/m0wQhBB3XCDxfvW6lvKAod9D9DiU264qoY33BL9Mz/60j0+RPUOjKcWEkgbTq
sr8X83lpoyg7Kd5ylY0cjvcy/sazqdTAMIGKiJFik9fZXDfd95lgL7KiL0+Wrp4wqns69jMf/nm/
6RE5MB8IofxlXoVFz0abjdPEmkKOghrjolkM5q8UkUAa+EYK8N5UU0XfELlu0k2gC9WbguR1dUMv
C8+gCTbuvllT4kH2l/GGmy8iFT6LXRpDhkSufBCnU/dMzU7xxU7m5gAYxHveXDIlpXmivMq//jhF
dmpU45zOIHccolLsyMSTRDmUJckUq6QYONofY+e676E40gPsiWYujJB9POZOikcLCD5KQ+eZ9W40
YfOFg1VZqm2ieW8H1EYwiJ3X7OGObid1jlCZqHvILZb1VxT+L9s7yKrkEWrK1XxRQwAP/Sr+KSuK
aUNFKQacLo51C5wtPhYUSt27Oqnj+MHaDeOkXkR2GxLiQTMKW577iRiR1Erc1K0vjfh6CDdgvLDf
w74RlD+lKbeM0ZLgQ0JDmXkh65m7BvbMMifoqI+HiNXUQpS0+Sayjvt2bx3TwkZLiLQIgVeK5Yta
S2kt8YZeYFdeHwmpd7J6CgxV7Vajov6FhSF3E5F1+poUx2XoZ833oIrguGqHP4JpzaslFK2NnGVb
Fsqm5JoGdHaGTe0uqqcxXXrloH04oeXjXUJf3TZbNgL50QaJH52rrwwDTZ2SvDejNTrTTmX1HANL
bSkZSx+RB0HrPydv1nFu6qVgnF96QKDtPzw16WOZ878jNXk4z810oVYXKaTQ8C31cPebJAt/a1U+
G9p2XF/1PVX0+mQS4CosB97uJOX2W44TOotrqgsXXxEu1e5o3Dus7hlJKnhl1IBaG5UC0aGHR8TV
JSmFmaNk3SdZh5EOcLG2WFfUPPf/SHrGPh3gM92rN97W/3h2K6P5pEhorCAYzJ7NvYFVpM80E+5o
IkumeLGHfU9qLRKmKCAP2LV5GqvlQMjLJMH3myjIYer1DggtB9V3KU4CZOHXyQ3An+XhkzQggAiJ
1ObPcA93y3q0i84Zu4pGWKcidbR83zIhHL8X5CtSGowcgneErOQkLAtVbWD96L4+9AI+WRF9DBcF
01E/OxJ9r0Rz9cwsivQuzQjUVJSjOXAEyG2N81gEJ68nERTwRAQKo4BWS5vA8brEK3NC54snUXHe
6Qp0eUZ0UsxQsGBYKLRDAjX/YMmcVnLuG+p2ZFT01spjExLbIHaB3Zaw5pJp7U+m2fqcAEvk1DaI
egesEOAjmnsx/L912BkvngkYjP/BcIph7xON3pRdOu5lXJit2St70HezUzbgj/RJasCKD8tufn+m
tAWP0vxFcwqRxG7rmJ0DcuprHne7qLgW7qKq5e9oJXT9wREqw/G7ZXTjgQN8LtnempXG8VnPnygO
0sykuFO9mzH9ve48ta6VQqD8L+Jebkow7hAbBlbkE3S1f4kEoMdUrG30WQPiGi8YEEz+Sx1eJO8x
cU9c97Lw6fDqLZzNxxJ3a011xRg8Hb6LZPcZPBwiVC5KIVUXi+T+PH2NV76Z8eJuEG4MafDQ4IOa
aLq0J4mT00CEACQZ6IPAJcTJ+XUjeljQkzdMoGTIozGtXlUyBgqBPMudEfQGiom3FSmHQus7FfsM
ydsV5keEQ4DUqN8WbVT6UQ6vkxcBrpAky4hek90c92jf68xolWz9Ff0EB7WuC74uE2d549Ut64lB
v2DA7I3+aPVftn6StiOlk96vsgwDN+oTJHubtQ06c+Xeu6yGYu2m65hzDp5HNziaqzGakr6crHI5
/RxiyJQOGnaHQJzLja3q0Wit0UyHwuFlRvqrogBAVBJmjZ+A0j9zdsZYNK79t46gHGTHeUceghof
XVePT5emWJLzUNo+8GiMex4sUvPxRxwy7Ul4ylTJ7eZYpoOrhWz/SKWnJzGgGB+sSRtPzidqGmxq
PTcPr7QnypXW9nMgdd68uby9GJjizcAjJmwTZswVHyHVQ81XtpWX4RMmGsRu5Cpwe5QE9pvS/ala
S28IK34kJO1HbknJp9+ENtjQJFqWAdZpmdhE9mEdQr/GijHXRgZw8TEmwCIpCkBZ/gEOdraeKiIw
hbttKvITSfVNl8uEdzLsmrf1nGqT7SaADKjp3SxO56niw7nMjEOS8e8SOtL1szW8BALrjM7j4vw/
VBBctmN+mSXWh0YOAcg+ffTV+ydQz/PNzBqfdNpEKX4V3Zg2MCPZjGhqiStBD5cECv2ASFb86bcN
Jd8B98b9BJ+Og7zZCRZPy/kCR9U6fRMR24F9189eEwffRv6Kp6FZSD1TbMCz3PkZM515GSOdlMFN
5PTo/dXl9Edorr1ShUEb8BNlKCVFmEe7c0X+gX5Po9g89NhzO2h/FSPEgK2WVNJWaDJfkdoFQqZC
INqOsESCrCFK7B4VyiRMYMUs5bjQUrpv5ACsHtDpJzo4BPJQXE+em5VQnkHA/VZpZIqxlJLBFwrU
pUaMH8cyEy2wJULXdRzHs+W5kCIZUZ4xA+FX66fhhzNNgNU0HT4u9xHJzyyRCiMliB7U8KXEwpW2
s5+JLv6xj7pJBkWYypz0PDarX1UZ6/idh/LfD1TESfsMPu59No12LVyZRpihzjdCcArOACrYkder
XD3szpExAE8ZW/6eUZ8cZVbm/2/7S/scLVfGn2+Yp868s6knBbEaSxuH93AUBr6zuvZCc7ZTsfei
BOmavUT709tG0+x2aEzh56ScqPW5kKzE8CGYcUy20Isvlk0InWElyKymuiBqZ0sDlsF8BqFT+d9C
NqDuxxJWBqVWdQFKKXhHkNACVdEg+pvm4MZbOb4mRjpBtq49nnjk80n6PZuHIwDijAxHc8lUWMQJ
cUvDxTLQk9acsK/ESQNcwjZhprN5IRvd1k9JnSkSXrwkNiMCi5mt9xt4ljc2gVXeKZHaNOfr7/bk
wh/qFtN+bu3tUgbC8br5mTu1hbMAQmSWU+yEJ61l++I6JPSa3wIN2y50aplh1y4KrMIz3iYJ7jyC
qo0WrZHwncIf4zn6kL7V8EdmDaKSkkFfwcx7PkQmAa6bRETBtas6Sbpz6zcqoNrJREPFGW87zPKT
GDBVckDiZbdToC9anq+REqvv7teiWjwQO566Vf832ctMfn4RzJ0EJ6YSSQYhXakzGfkuNbGHEMSl
PEMI2sm5KM9OFUg/yPJIem0TcjpYnvjZdA2r6NUgsXNRBGeQdedzU1uiUHwD2w4jeNcLHvMs922/
QWbEjCinA8of6vhAtfqu9IoIHLuxW05GVj9Eg4WvavJWqUCkD0jUfvewfiyeDQeJbcAdfQTcsoGy
9Xc1psYhj2nBMv8TYRx2gtaTSm6XBkI6rO2F5ohvR2zcSQAuSxECE8UWTewqVZ4xPJUAtDYWhNDw
Z7ip3GTrVxjsbT06OChK3rDBHHT5y+h/wEgPdGMudTBnTO/IfiXzzOcJHjY8BiZ8oDWbeTLjtj9S
hkKLG0fMD06Q6lzgUcfwcDbv2+JByTqdhEzStMEBS6ZNQ/7dl7WPPzfuzyGV3ClZQ8GqvyAhCTty
USl32BgVbXQW4v2jxZfewFOmDMl9zcc3NgzvyvnLux+hR0fAB21DVcdsJU6IaIpPyozI4XHCfG9F
oMNxKzcObbVW+KJLe6nuUz+Xzx1F9cXDKchzj3TkQmGIRBBIgpJywbTUqQIuSJJKUTnuDGomdfSW
s70sEM1kFgZzHkgN/kG/DsTl6IB4Ql5cqF8as7LQDEkdyr22FuHRf50w3zq+ibNRYlKKppiJoHQF
+Cy/4rOBjrSvYKj78HAHIVOuS/UKPdsETROOBESinC1IYi9W0daTqICwDGbqOBlUXv0GGobQBAKD
rs5KYTaYTLx+nC+ggxPdVBeQ2NLQFhXTmo+d0RKGBMoPsCwNovpjvMQi7812rQnwU1DhaDDemm4O
rxObyihffo2ZnhTWtwpn0LlJZ63LLouwfQheAMIOZyXwSYKDnVBFeFCYbmPAdC9LeSQRlfNWeF4o
ukX8BG4+EezDQy5FGWnMcNeucR5999b9Ch57v32bS5+afhqEoNC/R3tw+GkBOTlggOJZSen22d8o
01Ut3aRn2HS+yGVhsranUQa17fnw15l1agjJIr/Nwr7Ry+VsNYFIoFw3SCfrHBzuTn3B8v4mdMyj
nHDrubq0Gs3gGJg6nJIGj4wyO2wdjAILTkhaqvNHfR3MIa7lmvYHQILObXnDuSt5brYsjL8CVy0v
3Z7Xs2V6P2yF48aUWVS2gpw19hTOQWNxmrnbkCvckrIfSf5hwHg93fJRW/XNV6KQ5G7EWEqeRhOF
TAXnDPLkxNhu4xDqL/SHPfSCosGcwR/TjSfO7c/2rz5BvKgp8h7UkAQkq0PvPSSlonfL1g+dX6jV
vV6nUJI39A9i9oj5EYnOQcetCXz/FIZfd+3Qub4Mqzc633/1jopTuHt35gYU4kIudarb2ekdFeZf
OBdRxPyI0HbTUs65X75alL/nhpgbaQHpe9fQVq+Av5joWow4kXFS/wMkjkg4NJu96LXLQ1gcpQx/
Y5BYozzLZIz0a518FBzfamnXmDH6H9Fq/AQQiU6LWkC8XnHCDtNFGX69iYdbeANPL6/64FJ2dGMX
ovuOY7jNmPJiUCp+OsdH6j8cuSju+xai7F3pfsjQiXsRzGBrhjTalXdQjpjmVYXL3RyNeopd3cQ3
kcBBPnWY5LfOrEAOWdBG8Ur70ISwJtcvkAeYDlnHPi+hOlh0h08dQEa+i9J+AxLWdJWLH8enMe/E
c4GL1bbSRCf/bA0y7D5FUu4mspcKsE0qaC4rCnchPM/3PKMRmW0nT3F6ojUdZtOAkPnMKkdmr2cy
DPPnp3hTu6j/ARvDQazT5TTJUejlKb1VTO1KquYRVWJxlugdwUx5WEh4pJysDv6M5eM0F2GfSMtc
9QCwYu2llbNXodLWkdafrrrLKV5Sz9njhtkuZgkF8QyvCkIZVr2GTTC+0H59kBHw24UR9lqC1aZh
EggXP90zNB5dN9MT5RP+FeOGq7OwNGgJfesMQBWzkdstupKMVXQMcFxZBgJ/BlGJhrRTTILNVb7e
UR6HidQN4ESkNVix7HzwiurEPC3YIBc8aQ8OfVHybH6kBaxqPrzmd8iFiK+V+mTp8bFQVO4vOhW8
WBpMjduIf+ydWftFr1v4XMa7ZPJGmgJfTKiolSnWVbqRCdzTnkJrfyhOu0GmvjGQmH6irNC+5xSb
xdb+gxvnxHH+M/m2b3hawSatin3UPeR70smbfjPl2MQzOVuE//WEcrsDWAF9Ef8pxLmNfT6euiAv
UlXoA2tnB7QiTnV34f6E1p0tHPhyd4II6leB5P/bv+z5E6KYqVzR97Z8x4DdtwCEh5m0uBrYkID8
6mGesW9FkI3bTVmwQqBHBaoz2eI6xyLgDL+TzGGgbAee00ft1mvX5iGwYF33OugNyknJe0JSZqS1
gFCew6kwtpIBHR6gQ5F8AoRADbv5VM/RVBqscRB3LOSAhzJSGbIDowNnZ9gnEtqdB4qaU614PNwl
s1Mv4fUPX1YQRJYxisMQZVvv5MR6f8sdtZJqPX6U79bM1Enole0rfpcIIDdYhGi53pFKz5KB49Po
jK/JJhRL6yhTpfi3Yi1Wen7uHqKtm/2ZPKGGGlb+Kzz8lEiD18sIXXpI++AKZYlf6RxJUr3CdK2n
la/eDzsfIkxhAlEQ++Mrif+QGhW1ZV8yzV3bbvjMSn6uZl38p0oQw741rDEIGUMCnTFXtFf1Y/uM
p7uRfKTnwCOs/TcIwn51pZqAFGU5DpB4NOHlxwkXvLhVoqpKO06aXCA8lKIhRyxPnE0L5pf7pwby
+MnFLAuL85bdUrWy/AVPxmvL30rd3iu/U3ay/v2Yp12sjfx20npEtsUtYSFiiweHdL2rLlz1Cnwv
X7I83pK8x5W+y4lCHyXfNzAXdbD4Xba26beArNcnEZ8gfX5vRFruvpuC13XPPp5YFsOPWerH5kFR
4ZSpVsJkTULX/qN6ux7Qke+42JZUOo2f4tSfnurm3Rf1JaPttIoi1V45/+QZ88b1RBcfSNQ7sbpo
Q+sBsdd/SKI6u5oy8ugWWhXKqiVTPfOhRsFdnynxssJxPpsBYyPFhp3VySVuhyUzw9T3szufDV9N
WPa/c/GdJU6o+jD6kmEzkvqAQF02v57o7JlCwYnurGVuNU5d+mzmPEd7hPPvjYF4LsHUCRDlQ996
pb5vX9VphvCkwXwNI3CRYKKYnipZQqe4IEl3PqVCL7WM20EQPrU21Odh7UAQpiWXL72faEnrPkkG
fhWaz5e4Mj40twz5sgydc8bgPb/CMZSqRVIgBwAJ+a/i8xJhwF/KWMvlxeLElp2ny677HwyGx8Ko
PDgBTc2sHMPxN8nL6JXvibxKXmBYHnYxxGvVoc7gAx8o3aAFlTK1SEcATBdf24kg3UYG+8/YsiL2
DpMmG5DhrrvvBjF3D8GOfhhe+n9BEgi/94F9xbehLYtWFW5rJVS+Iy7PBfp7xy9jr5reLbXHvxji
Fci+gIMwtwfwmrza3p3Tl0FdyYAN4d7VdoWqsSTSe8igtt2twTNJYn6V2KQyRui3ZFJa2JLbji/z
pNAQ4fDDu8Ysp95i9qxA3mH12vkkus5kFjIccDKd46+M/L4bzT79JX2UUv+SKahBV/DbWdEx+X/V
qMZxJ2la7AxUNz5NX9O+snCA7Yw51rP0Fxt6LLw6JBHnj5WpLxZOc2e0fbsvEMlW01W8RoLJJFoQ
bTG3ssNPs/uCBmCVI6YPWsP/wu+V8ivs8v4RAVGUDBIOOz0+TzTYxAR49lkNwx6P8jMfrMuL0XiT
Y6xUqPtaTnhuMkQxlFrn1lawqZ1WDEm4WoGYHUonIJZWnHuwPEchqsnFQQlT+Z9WEpZinAEG0iI2
7wnyiv9LitG2Nigddy1EzGX5dbtjb8epsqRs2UI158ND7NfAPTtV4DF5eR6UGeEZ9wyOUNEWknT9
uVXnEj7pR5m+kOJOLv233Zp00vX9WhrgKq2GdGaHn1sZ4xWTK2mT/HOMaKv1KzQ3FSQjurTiShe4
2FQAqmN8lZ4cV/I61VEw98/sR6t1C5MSNonjNUCc3/3dUNmy/meX70Er30oKckXbBJTwg3iMJfvD
RUzMGL5Ox/onKakIZhPBrj+N0x4yBBzLh1HuGZtHX29kskekWvbDNU001tkoav4xJnC1AvZpRJqe
/ziM9BXV90en1O3YMvxo/5uVvYIjMe4QKJr5vRqE+XAaN9UYuA1k+i6VOtCD2D/ZM7GLzNQSVc6j
IuIJ+YmhgCzr4yUvyajGc1Wub/9WiRkLJN9oRRUD/kUtXvxzuaU6ZApkJZsJGmRw9NfcQKcFiG6K
4RKr8PKg4dSihVffqWttMJ7P9kVISzgDys5H3l9VUn/qvX2SQjOATC6wEBu8S9tnJDerA9xckVao
iJgAwVr+Sx1K43nN/wEM0CvqRHOzAeqIoqtN3fAGNUR41ZLUiWoHX9GOuDI5pMQK/77zQhZQyFuX
+cYM4XNXNBgn7PLem095popOEiaLLmtacO30LXgQZl69fWEw/S2pizmWbJJoHcNhyNBPymjdzrOb
TWrEzc7iEAg/kh8NXm46/6aoNAxDgC6Kj2vg49lBICcBNCbRIXuIoQfHT8EIUuNzyFyKyfPTC8Tc
jJKpfSDmBjGVCuNypXb4pLz0FLUpMJQpCW32BbjvXRSGYT86iPkwLsMzL/89fBcB68a+GOiSCTCP
neX6suT10Hq/yvoaf5okwecx9hx4poYv6O13VTMnHtrAm5eepdepZRq+E+oXavusxV/mEdC+l9cm
gSEpDT8GN0GjCKrfnA5S5BdJjFIcISI93JCUet9Qxo38SpY4NThvJ0cLLg1lmQ/g82RgVUMTkykU
nbi0JlF6lspa9bN/wSyf8Djl9TI033nV9t12yYrxDDv1HnzbWFTGIfMs2/ZP/cPgn8nF9HGboNvY
NSN/VflOmGp3aiXacU/KbVmF/AuVVA76ayav7pgGoA8AjlOpkup5GO1ju4iSeKreDmQLy6H3NqNh
N2hWEn361+PlbCiuy+1zjxSWyAb2i996LERNY8gLwxHLRdLIRUxdDJEfgibysiW+NK6CWrxBzC1X
4p0J7rCo6k4gabjmeOI0BgnNKT0gdUuxMXw32n+ubwbF/19QGlp+kZ42QDdK5L5hIbGTSkUBLbeG
KoNMGSfxbDDSZBE5wzAYl9xB0G6+RcovL8diLXfnjrvN1d3xQum57NKEGZkPNMtGQmR0nzbK7ufL
RZNA5e0/kcWLZzyS0NGZqKb8Tr8xv185Mj3qhKWlYsoJW1hOH/peQoQBT30enqkVRpp2dnhHLvvT
rfJHpIIbsxj3AUsIMVijq//Z8cfUh6ywnGGZ+V0RghV3T3ZS6PnYfxUkz3PonYvgaldVCB99yS30
ZXvKh0H9R3Lz6yaan+TkXrFJjgodUGZp/ndWqtuisT7EL8Exk5ANlthvvIMwuQFhvK4SWPr9ZLFi
qO9ja0yh8jqUbX4ysLuWGaXAYnL9HCmm/nt1VyRHYfIrtNaKCZAWM6bTpp/P1mZCpF+wEW0mKbKV
g57pSvNnOIyeR/Q4nUBbQgiBdbELDktpZwfG452xEmveVJfZY2oBe/4xGDuYhK7CSfnnUP6XUBWW
ZPpRk1NRmfNdoTESf9bAvoIEKCYpVA94opFV4AGUGZmZwsiIFoJoW9HzmuDhczpIxhhxfzDuhoZS
4bnal+miuHLjZ2i8zpIxUSkow/RLZLVkWkX4r1/0hBzkAIAjD0Ov8YKs/MER351HbnGoN86uoYMD
Ao2lf2Tv69ehocNtCpTD2UgRKJCuMG10VxztX5z7V/3hMdZKDNDuFFAkZiSMjLngFaaw0pHXO9IF
HBSCx8rWby/5LzF0XeUHGIPXXjkS3Tq+O62TfHe/O+5vi0/f0Kv7HbeadcWAyBa0E48Hhrpla6lB
8LirokzmvG1WF14AyS4cY/e9BfLhggDLxKszCYa4Ya+O3X/RXF1Jbm7zQuCInFsoSeBqU99gDfSK
0IY9JstVOsKxeGagMxAlERq5sP+xA5mZxmT3DJKbFeTmTU7xkNCaagw6xpeNv4/VSYFPyFC//+47
dRi+zWSwpZRvk+9HDky1DghEM/oHgyz7UDeeliI/pl2P4o2TtHlJYuFQ4lZldrKXQpQHze7E5sOk
kZM2KVEiMEWJhpCUHTdPHm3oC1+5jLSOkO5gkMKqdMcBFRybr8lUTK5+otXuck3T3cgdkbtMDY4C
rECHy4WFId6XmYf0pf06Bb62pFbGd6iVE2pczSETe7TcDpPDBArMtpaPgYxdYYDtBMfhtvrJq+oY
6ckRdQGbTDC6wwOEvX395axsDykvEad0H6TonhGSfMkF1uFZVMIjJLY/wDt/93w2onpiaBnPoBQ2
8rP37WI+kASZcMRzoXs0F/bdzcncMgQqaRW+cPKCKtoyJ4YK9saHG2Pi8BXFmEiTtN7BeoxMnwAx
QMzm1HM3Fk1q4ih5CW2IhlgDmlhDtK6wQeA+Q3cs5HX+Wz7jrtWSlsvZPMmOOH9A6f1V+3Eklx84
6yHZsHWGTqcbg2U+PN+d+OY4mHDwirt3yAlG6V1jUEHdd1sANg3pLIg9M+vpxkt0lLMLEBtIMvRk
gAysEJYLPRQ33NseJwHdxFPWzebamYbATg3Og3PVZCHABQ93BmDH299ASLcCtskkyeCQzxPBorZC
U8ryh6/P7q9oC4i9M3T8O4G1OJTc8Mg5mIKe9CrHgkJ4X+2x2vU0axyJMPRVanr7GqQBtXXiXWCS
JGmPDf8aFDhbT0zYazrAl5Jkvx7E5OjuK86A7/GBYlHngkEcjRRQufyY8CM0PsAjj3KxFrMTHB/u
K1U+RkYBwNQAYKhsNBGtR0ZUw8hzc5rKV4wq/TsuSgztM0feO4ezsQcSdOtZcP2gAVAYCQShPhup
XpyHdj4qSHg3Y9xF86MKIkHsXVOfqqJ5+sdTn/ytGfMdmzIllO7HauF9Tb8mnhmpy2EvSBHWSWOZ
VqIarVS5S0oPJR3l5sjXrZo1izkjmK1GrPlefSaEyxKVRkJb1ehO4yvuAPIEwxTCEhgdl2WFS0n2
+fOfQnQ5KV30kCri/XMQ9Mx5xuq6wjbYbS0eRsYZXAajp1Kurh9WhYKqnjDAL8Wjle343KxpyeMV
CsBujVjDgsrb6C/zz/zGfq5ukQx7ysfUI9cuVmxAgSAXHVycYMayzyb47BNYzbTmkuRhCxA8yhwS
WY8bEge9Lc70YxGlBkwwyDuT1xwnKBYnKtsftHRMhYSUd3ETiCRJ4oyV8mD7AfgQrb6u9fhEohmb
gcnKohw7X2E/nryb6IzvD18+GspavFes1CsZKxUMfDJG7GkdJkBrikUW7VFzph3stBpIiUGqjJ02
9zjVYNR5Pd+NbpVSndubHuySoSjeWUNfJMwwPAxr3gmVwEJuAjAZ8nFPzqIgiLCprg2zxpiH0qpz
P4fLH62KXbppl27OqJ/tn3kJ8BlEDy/XrTvZarzR3gLKU4OCLQm8ag/MUQZIIHT8oD9Ji+2f8lY1
JioZ5Pb00et7MMLT1upbnvIXZd97rAbZz2i/qYqCF1XtboV/6n8FvOnr+HPdmrAg8oMjY5LWkgKx
+/OVM819DDSHW1g1lQf71Od2mXplEjW6iRxiKYmIMOQSiFTZs61cCXylcCIhIlueAmEQist/PhLr
hDd+YyEyDuWOgTO98xLEqqwQKxyv9yMNDUU0DuhJb6th1nipj8ElUCuF/xVzZipo6mfcqR52xVA9
OZwlQvXdRKnm6LXz+hoPgxxqOaawn9mY6+Q2Fr2gUt0HCbEFH9u2PkGTfrYwu/7pX6xXjSdAxMHw
RKWsXKCAYHPRuBz0yvazkDqz1sqbsxOdDdW3oqjfMLbpjWCR3fD/qeJMSQ2nnmvC7S2ruxI2BrL3
O7vBVx0UFG8OQZJwww70ZfkhYE5hpeh6g0fd1Bl7TyWX9SJ8aEwPQ/qvx2IMkza/IACG9yvj3DuV
amd6CfWftoCb0NH+/1af+eAPYXwxvtAmC43FuGNnbq+C11QzHTf4uWjXZVgb9b+/TM7ov22EviRo
fdHXPSrsAm3x1kVxyvJgYjd8G7tVMpb2a3ArxQWjpAmrv3QT+gWa/DiIqjAE+lYWh/ULEwZXyC5X
F0bGzPRjfMwYPWdHR4nJVnrleNlgk7rkmjLuNuJmYsMkHdIhrGNkm8gouKp1yOk1/I5mky2NzUYI
Eawc8xmlMJ+XSkB3rBcZqdnAiaijx1MVCNqagL6ojNbNd4p5FCDjEr/zd8q93O/dd3YMUfk9AsHU
eGIaDRQ59026blvjrEOQKJiaI9BedYQ9z7hK+fJim0ZCf8ihoRCJleYh/5Depy1jzKGT3fbEmGiC
+BwDmnDn6e8oDgoYXK30BHxnS/8Kh+WYwcIpBpE4bz37ESi15N0WQnck4dRCabP6UW6Oagc2ZHNn
Nt+K0XfoCFCEy7otpuDcqks5hLTJ85LsQswdpOWWP1mJtZgQ6BqyfHX/Aaw1twP9Yur0rTHFok7a
WEKLmso0C+GmFOcb4NRY2whJCWtlY4KPUYVECSShazm6AZzpZN1MsSt0eTgQTHjS7NOsUFFuqpMH
dGS1dKx10bPtZilotbpKsHbNVQr8Z/rUjwBnhYlFMAbDSODtvIkJ85q0oYQxL6hGmC+QOApQVGdF
vCnMbuhUtM0Xtpo4uzyfXatvsxfvyyCeb14si6aWTdYa+YbXh043gvgGy5QX9lyyb0pef1g+z3nA
ThlyHW7yFlxkZn+d2Y+i8qfdh2fZoi+MxM0KRx4P0dQfIAhdi98zDig62VsmdDAARlhRq6QoVGNF
kMAtnMi4/Aal7dfFVipTodd3IZerMKU29kFHxKjBt7swd/j9/t3QixoQW20EDAH99c3loeYV8gKx
OmNsvcXyMevSvHxMMzlgseZudVJgwcFHozfMQXTy1sXPCJmb6/mO1GjuBcJN47V+AKC+Vwpx+Ub5
1OHweLs81G3+i8N6ZQckqrerW2EIt5eqbQdRfdbmmgUlKOa75yU+0P6G5yxicLsjLiElVGjXXpnP
OlSPUw3jW9BYx3+Ro9J5I0CPZUa5QjS7Epc/AMvNxmxzkfUO9Xftky8exYb7v/zO5hOouFSmqfnb
x9vv6fPIPaupQLM6INmnjybG2/o1lB0SXUQTAdjemWUynRyeCb99A9elC3MopkHdYdRdzP9eghEV
THYx9W3ERGWi90n9Wf/EaX2DMbPnZrfOTRGFRQjebB6F3Jbgylz6PLqaujcjZVP+/xstjJ6l9OjP
rxRpUM4kFP3Kq3C2VXhLSkFMltq8keClTIcJngYOkJjK+JZ1nIjnonYTve/DYQRkhO+8+bxQXHbi
H6fI4LdlqIgDOxE7oCG7iH4PBHinObLFoPLg+TKMTl/bsJ63dj3tYmofjVCnvjFmj2bAbXg//oMR
5IqTmhT2+vJ/6cAoc1aseZOkFzzqjuUYoGiNDn7MMdeg7AcvME+us65+Lv0kENz/98joOwujQXw/
ctN6tr/0sHa3giga+u6riVYN5UKY3aYcfFbMEVizpovT2J8HTiE24MzVL5C7vmGnuD7JeCCR5DVJ
eYU6wXth33jpmpv/yHRfI/UM57CM7e11BmCWB+y1nwgIZGGnCpp5XyDHaGW1oVk192vy6uTexKSh
yABsrMF9BJODlm0OtVbrs9mjk6FEdwHE/L2Yk3llXXtsUbxaZbGYqESd9kVOMgykL1lgIiSwK+JC
uWn2ALGFypkD/2r8OnccrzF1IuoSiKjItyoQ4LXX/331o0BjFFqTK1H0PtEIP9Zfvpf/RnzEAAJd
nGZ37v/FzxgHk/cpwdQtaOaIGCP0QPVlNt2+60p359ggFLu7pMhruUBDp+fW5B+xg3DWh2o9ey+8
4gN83oP6INNa29wHpSghbzJRlbTWr5BGTyTDUoYVKobKs9SzJlMv1GL0zB3M2mk36kJxxTdnRJdK
FCIE1JVaoSL/IPdL6beKeukOPyAhNvzBtn6LKfJnSjhsPHyjrjOZ1regor/+d9BSdzhv88QTCDQS
MTLsfAFcrmaUMUEzfbhiN72QaeCv5XGNDkfZoK1Gg8BOjTHD+7dnmaka8nJuAN3BDNSN4oRHl0TA
03JQ4hz7+TkrwZR6KmjVDTYhubYAfbWqamoImo+/z8e71wRXKIiRDgVLrYD6ISfQHw4gBx0SmtRP
qtY2ugQP1BxiX23oVNhi8eViBz5G1s45oFqax+h6PUDJtbMnpr/8c/2k5NEezKTij7XbhtCJtP9H
/oN1pxo77IPLLHyi67SfsCW4ItZoD+JRzgXiqwgSpliyz9pnpcWt+gZBk9vyMTfWMwiQ3dYsr/O7
Q7xumgs+vUPlaElfzgiNLqy/SSeA4LIYsLxQVd0hR3D0Q39YQlxxXUCfVQHUVIPoPf7AXBUMz2rS
upOnOng4577yfv1L+49R79IEJmqrsR1zVpnK8jLiqE4Dgo+dZq36ywbImO6hDFSm20bGlC+U8fg8
zt+dOhjQG8hrAKXvFr6R1ZTBTWwE0Dx+t57NcprcPsRCO0Dhr+tN/PzQry/2SNjwoBfJzYb27tJW
p/9mEpAEUabh3O4JV1yTaGGVCzCTaubO5eYkJwudH/Y6fODE+saEIy7q8hH737dcuGoMltPNhHXT
0XqvKL0ZfiqgVI2A8nQ77CyPkbfed/U4t6Ecop/DozL/xyU7h3k5V4YrcqV1apDLOIN2kIMyNZN1
PHemqJgCzwWQpBr8/5kUSdl4WaYxwa7RN8L0mnXwwO2ocXpUxPTTZAwyNgLSDn3+Gj5HyXYRST4V
tXS205YDQeqcLysjrbEY3aWTbPXQ+bBrC3b3Sh5Lhdg68q+F3vVPeVFaogHduAP4slZj+s+nDPk3
5diJdMcTKiFe71D/pDulnKDW2jMR+OFA8jgeg7+ozOMH20IbdVhlBDVAwaeSdXB1XAsN5r5ZPIrL
hAj/HPX7v7tPIMqKFiyxbQskFvQ4umRG2kSki3XxP1rq3fA3Qee21kmfYOFeJhk7yPdx3rRtZkZr
7fRE8iWW02nWywdpZWgOlp4+IBHN6w2BF7Bg0/QQ2eFYEmbUy7qWfh3yiG2eJt/6cVNKfmP615Td
06fQV7EQIT+Ank+4WhKdHBNYF76JFoZs+zqGE6G/wZJLJ2IgBN7U6XuB/pLBHqTgCfiOl1+fz0Np
PV2cGjBqFZ4pqw4HuVtRAJpGwQrngw219BBmUBpoW+TJ8QlKYiF6uRyXOHSKNymvLi0wLDTYAlo0
/+Anrom2ZNW3uoRxrXxOytOQ4VEk6gbcUmrBAip492GEMecEtRgniNRluRpqaaOsZgyq50Qvv9D3
PUewlp4Fxg+Sc2yvqotXqH6oIdhDvPAC2NjsFiXzZqDE8QRYK4Fw0B3T7DywI9tkmF6dOqn80pLB
VqNiPVkwgmD2rxe79nLPnZ7GpLDv8FtAhDK9906Na1k8etxleBQ3CogCQQjfkodAx5xKTkgvV33o
oQfGG9F963+jfnuoNf5E7OAO1ihEOBmYKJQ7g0NlaJZbTtFx9nHMA+kSn6DThByxSSgqoXap/xZv
/ZJHA2KVKZhZMGXGZYrIEQ5GvbbNVRL+oKMu2txdq4CB1Dc1I7iQ42byMxubB/obc65/xgNerIiR
u1ihhWtjaWSQ1LYNxdvIXdJ4TQ5mzmVvU4mvzGW3r/lf7FleNJ5R/LdFmmqO4lkpuAX+RPOhDczQ
f84r/V54Ur4MU/PzOYztBaMz12mmtejuWRH7h4h79D7PMei8ci6bliusrsBKEe8aUsuqPIjbxeeO
a1dE2LvmT3dQSZYVi7sxh0NkW4AutudzCK/U1B0LKzJ81SW1Cg2wk+kgf4NMtbtCkuMaPgfGGwU2
EeNpUhjXtodXobFMPQJ0EIs9CYG9Gh4VC/nkNiWyct968OCyaBeDck0QBiyD5bX6t/aM2gsjfCQP
mT1FpETvwX8km+JiTkJ3hdYh27Oe6wdq9J/qLyu14X4r1rxle3pvT0jyQmnQ/AieD0QWinuZunMo
N9UdanzdMx9VVohdnJQ0NfklZhDqaRmKggZGcq7xyfqn0ucb//tdSPoJjjuYhBw1U7NcluvLvCFi
b5gE9Ki7CXuW5Z3VojUqmXtw3syah6UqQSaRlR/+IeWW7uQdi/98Yc6r64GLeUQ0PF3Zq72Qn77E
5Tcj7C6njeQWry959WD7zFbRXz3LfgT8y4j3LZ6aotWP2wCiI8fRLF94s76+o8/9LO7KBvdV8HzK
53TgLnhs8d2Jlxkyu6yDa+cwcwlFbPFl8ZlOE8Vnlo11Kb7woaIuM8MdpTg7sikzWYoX76vw5xiz
9EgOP07F14X7O4KKNc4eDb4N1PKhMCFecESQAuNYRxgxhLfoMcES6+Te6EqJG5TkVACPXrFb9zi2
jNr17d2JbSkltQr3V0SILzKsTu+7iJ5kNIJlanf/mfWtYkOuFkvc/jI90lWobX8GiCNsfOxp4ZE0
agSuRHgkjMgwYUPopJhDOhOaJ+P0fWazb84rjDvmo9lxREEGZyL+9xOxY1zzmTcFMtFMuX/ytWmG
w/IQIbBE4PhfYIZoYBorpvotoW84LxYSwh3Uip05uIEOC+u6EcOqIUrTLPsns5RWhQ+LYwNz1eV4
UUw9Te7zU3iyyjNeHb5DrGOpZjqtok5Jt/OjpCM58PzpgZZ0bvH34raqR7EtZTUIrxNKxH4Kjmzg
AvObXeXkvWAKhvCvUNf5bCfwgG7pYY8QcSmemmF3ExFemWyTDDdoqYUMptqrAOqzOTGIcJelnXvV
UNOzTpnOZ7HMHseg27M/qYVSTrTx9BUzD2L4BxVueFvCisnsvgIP5eEnk3OJ4k37tnx3CyIHkXW2
9lKGL7SW9rq0mgAHMnf/7ewuz+UR2//MqfdEpT5EaTsFlj2ezsL39zrdxdo7PNwb9lVy71dW2sGI
HIEiEwMau4wPUNDKvvzWdQYuOumJM0SDOnQx52ywq91sHt16gWprhIyvez45s4e6c1r3Vqrl2XpY
LRALPT2V68P4BRP/UydMkrxy8N9JJbQE+9Vnaf23n9Evyfd88/C3X1IHShctr3PJ8tFO6rHv+JbG
7EQWI9PD10GEjx76qB/UPW6GN5zYZueAjaerUJf9Zh+09hhq34z74RlM7H3KolEiZIA9Idf17pQp
9ElH3L2oG6TGfOTZb28u2E3QgD7gaWiBDIlS5sCL2Rl7TJaxs+QDMJ6kO5kj2swp4D3AyPAJ3nGX
Hfzr3dIRQ8qNBH1VRW+FS1q0E55Uf9yQBGSUhImGe7W8aWb6Eupg0PF5ApGOCBtDDkiHx+a7C8dc
wAmQCFxCZKEstUn5j9urn+8ezD4C4y+VZek7egUlozuyixkN+fLnfU4TVtFzPpQQzXUcHP916FBf
ONibNuJS7feI80lQzJKbsJLzR1+4bXwZ63XDHjXgw+VDYHrFCEAHTlVmooOoHyz2uNM6uaCZa9sl
0J9YirFGvJPaqSCjY7fCvjrpy38g9Wz4jY1NehJ+dsTVKo3+i71q6kMFT+HnPNWvw6fKaJMWRXuD
4iEgtoBlXp1RzhV12etWClxU+ziJuCu/ALiBGehGmD7olKsczUiV2DJDD/UHrHkX2M92OSSxLTIi
dCqGGjTkZyKj0+ABpWD5Z12x7LNPvxEuQIGsH2vngZWoks/eQ/3rueUwEwdVqJnYjxfyIiUXkkcC
CKZQi9ksl/6vJRG4d+Fwy6J3BwEyECaTbaOjff2rlPHPAbfK5U8au3f/xgqGLhyCL0KtPwJSVfxf
2lgCNvyBdylDjCvAYZAVMxn4i6hDS/sTZdRugEx7k98GtUF9wzpsh/fLsEp3Xh0h228FOpWrYUNf
qt6zLXCRa6tsFU5k0fjxCMkr1d8POysdat+dAKHfmGjZmSyjLDkBT0psOJtLYdQM+wNW8LJKFLUs
tPLwtEXML42EIOI1di7St43hdHlItAsDoetobthz8luYdAx69NxQT+MRFDJ92somNfpYEB7lg2KX
mZK7g8oMj8rxsYQZ8/G9UeMegpmZp2CBg50vs8wdh3R9N2qFufdHnIj+RQFBuhxKslrkScpxwVhV
caMPXKl/HREt493YymYQn4ND4AWH39SISGiLPrnBe8h2siEbZ/slnpla5G6eRUbdidAriEYr1Dki
2bxYD7d6Rksm7KGLEAVpjRSsjEAQK+wmAMI8ObTfxlsYp8FoksCQUV3TaCSM5QfVBWDig9frpULp
YrLug9g+R/TVyvSktG9AwojLGAbqFEi9jis5lcoCfwkZX2l3dEMnGhSwXnlvEX6chxtCyl+6kPK9
ockuv12+QiwkAgpI5wqX6THwXMV6ZVEprktb+zRtSFMpur7QGrQHicsBrLlPZ0wLygZYfe833PqR
F/lqvD5xmz1WiL8wqr8hLwOceyD3HQ+wx3oquphYrUg0UmnlB7PwvEc6hoEBb+13ZBAS6d2xiP/j
510XIpZFmLnmmLAZrxQ1PuUnXwxEWCIjMv+T3rJl9GdKRuKnpVjo8OASkMrQCEhR6SuwuUpSJ8T7
3gJtOGMG7wS6EJx0/BcTtHFNEtk/1Nhv3K5aTnI3l8aQPIZZwVSrubHZ3YpiYyuExgsGDFiFqxMW
zXG1AhPjzHfFB9iFVPwK7HeRQclHFarrGNrzWKJPu0yq7GNbbflYneb5i0NxGPPnZsHkccmfTLss
1n27VmpPF/IEeSprfvhQCEYlL6ukNsG4cONuHTm0CCPxwEup/rVUTBbB+SVaJsEKSNkixb6h9srl
42HNKVOOOceIPF3EMFlZTFJPAfnEUzJRJJB6RnC+HEpdxIj4QeJwipI7hXxYqtIlHUo6Q3bMxWMO
pWE7uMcfq7ffXS5VVx1y9THxN0n3VUqcfoHeqrjcARLfIt+KboJ+dD9QO2VCMFpAq3mVmk3b9kSd
zDqs23KsHL+uRbQyLErQTog4DF2dNezX0W4KQY+Y5I7NEAvjMw9T0XcGcXOjYjN44edoWGKA9p+z
rkHfmtru5Vu2fDBtn0Eor+daqSjOeZrbZU155MyQdXYmznXfMVI/VwiQ79QEou+8Wfim6qkN5IyE
ptVM8ZfaspPb93Cqs4rDhZWT90+lUyD0SfDUbiTcY4tCniBxnGe6PpTTSufRPoTQ1JkAuamXk/8F
YwN8FcMPijjSvlpe+DK3cWI4lvJV4WIcxjl/OBWZSHKjjD4vUfEvaHr12RvtcdUdSsZg/oK6xw5S
eCGV7YGG1+0mzY9PcP9omvEIuwg/7wGOcHNkiXttle/3xlNA+CB2BGGwPA5mx0Tp1r0CHa832oRN
O4xpYRuknddcuSJRNaVt5BG+Kc+OlaBYt/u+RQNpTCeDs6BMcUz//5Vhk/ZC1skfBKXZWtEWE48a
xXx7fZFG9R4HjLENYA1VVVszM+jqsQDkGO6kNTgQ4GrU4+kObtUb9eICNNi5gvi9+gkGWFXtkdZi
oR6IfoXs+Z9hNT249mA4gW3PPnYTCadckxhgM0He2xZuY2YFuZ6G837gYPcEkCMBugQG357TFbl4
Vx0w9eKPdp3K+y64RZiLVQkSrGcKAA+fY6hONYVk2kdVgf2Pf5JnEDqTMy1+VnIj6ag3M6OEeJ3U
LJBhNYtBSOkm4XzL/cC63ZDOXNjrZAIKRhvn5Ld8wjlndkqAY7MDwJV/feQLYaO7ShPXyH4HKPzz
q5ejtYaxzHkXBAr09Q2YlYrMRF8o0rhqkmSl7aNTZsA8eWrzWEtDELStbhioU/G7r7qL6jasohV4
yK46a0duS2aShvZADbGD6eykbvIXqMqwQu5EeSzPkZNVNfSUFOX/cCj1hui1FaRPiWhNSvtYXQ69
w9z/icWur4e9xQRLm2aYrGl3GvR+4RgLQpr+S5eXz3OyV2VCbL1gPZydPlcc6ZFQGRERg+LIDj7U
4A9qqAdleuSnahtzSYESKFxpa8UTLWshbOg23GLB52u0O3yGKCwNwSGmcCU7wgJqZTFPTTJRSR5A
tsEaLf5DdmPTVkBI0gyIha+p2C7c7dHR5rr5q97djwN1Ly0h7j2w/Gb46PmCtDWXj0QuDLaiDkKn
WvXu73v6Fuu3KZ1FePYAv1GjUccVlfIvVUWvE0R2stO9mCWZvrR529XswNVNvP3J0h4ZQ16JjE4d
mZSvkJgHvgwJSIywDH/kJjzd6hu0K4NWM69VpwTjxgeE6sbpEvyqacnwS5tjd3OOoQ5it3Cmt+6R
F5n/CpMmJ5eW4YefrXnFr6UOHWNpdTrFYxFAwiDGYRqx394Lw/es6K1b987jAhxshsfLpUofh936
eKCVKbJ8gyqeIxirKYAzscV8yg5LPb7j2I2BtrAxVyadGSWXS/KxwF1VGfUlfaejOpd7af/s+PLt
4W/c3RmmaqRvZZaUH2dsFOy2w6EA1MdeCi0o8B9no3cnhCuVjzTCKFoBkO5eOA7XNwydzUWsEMk2
wqsYN115SX/wA8rRQScHFGY86lGeQuJtnvDlGURJgJBd2XgypT3MLURvbMba8MXWecM2IyaPvAI2
AMjR3ulwBn/v9BOP5fcuxj6DclI18JJ5RwHgVZMSBP76D7jCOfPvnl7i8SgJGD8gXor7Dt1BckwU
flwQ1GUcOzBU5FzS+xSgg7uHtCZ4XV0At6eq2UN1nddPWa1hWYrsbBNsQnl7LA2abD1cawRglKji
tXYqPFWtSChtrCWPJzoERgfszrP3A046A1fiILA1rtjp2fur9C9LlCjAZM82L1p8z9QO56IYtR3Y
iiCXyowu0qNl9Jf/CvJZrhAkVJnwxhs+h0SAAHwZVpEW/VmQpgvNvlQL+AKoRtF5vXEi1lAhR2p7
XFNXczSkRO6oLG+lEyvE2kUNXL4UPtw3lrJtyrbPwxUKbAF7p65BdTdkZFGZkDYzl6Y98OnRm4Vm
joNQRbw3Ytm1D3EuIKnw1oKEqyhrNdZdpJ3ZT+DmmpbtNC+ymo8mXVzOy8m8E3Q1ZPVk9E61RBMR
WxO1FAR0ZLcnIE5NTmdaKaHqu/Y+nikrV7SM3B8ukYJCV+W0r+GG3PjCrcCWrEn+3qCEUXDTRT8y
7Tq0GY5rkRG2JuaxwU5VPoj6qzr7SwbUs9DI3rp+bIVHr5r5cFhxqJcVhaLuX24D3hwvjWpxoGNg
5D71fPnnO4J1oT4UEpDMsKbartHs8sqs1QzW/CILMh7Pi4WroqJbwIfoyaOQ0Lq1ynQNVb4knWwT
4f1e2+pvkRKBbDTB/d1C7/ZYgqyNfEF9/d9rDSHelB0FqqN+VYa6BAhCpgqdZRRaHQli9kfFW+3f
DYqmRUKLGhn8kmM+ZEPUmzrDifLXY90Td+kFTLpJr6yYOhET7J2rKm+IYyHDCY6wSmJqPOA0Ha4V
ZHLEsfDmNxcbM/epe3qRHWT882J88aNKdLfa9wQlGaCwRTeCFbT0zLKgM8MQS71X5hymUtg7vULA
tj4NULzHTZvozbpeKTUqyp/j2rK6IYG5lI61LjZuLVq79TpqqyUNrPRheF3zL1SNJQTUfrD43+Hf
zrf1/4HyDz3/OpPxxTPrc62sn2jxtRY68HXiM+6YaPqdgShD+kQ3bncK0uAef3RKAE2fu9KrwEr+
Cvv+QMuygQzJSKuhdcwIQt6XGeIbwGxEEjAMjbdF2W+KbM4AxddmASHiDRD6w/unCwO6BFI1nnlI
yjF3VR88X4Dgwe3i8EYc7UfeHxaB63acj1BEPWFapAF3YpabztnQu4mvqZWlOXsDJSp8yxfeSLPC
VacrOm26LV5/jmLnsnADpK1vgMWNxoEG9BHBjQOPgEX8xn4rN/talRohV6/TraJYJLYdviLu2JBz
cpe0uInfOD0ELbvFRugMpmjCatXgdhNe3pEmpi0ByBVEu9HbCbfZSpt5rcQQYagAtEyMe7v1hMMD
6cV9f6knF1eSoI2poeE5aUA8PucghSo5aWXCbKBpe9yqEpeTf2Xi0OR+p9P5vQd7dGu7Q6MXeW1v
LvCljCjQEopetxPCoPstQVD2YZvHb4DJ1AVv9xvms374lsWxrB04h9qZ6M4uPs3jWK721zRM98px
j/iWvAdunisdTfgF54DYGGYz5guOC6J/tqfNdyAV29A7IF586uNL+DwxPxNTyKtR2SaXwzHTXNxq
KQDSxPHEiDEMwcr1VN4ASCQyWoSNE6AwWnyRT4lijpFuyRnxcG2zZ0FkRC8NgbihhFEob8nDetPn
BKN41Q/QHKvvwajIjiUOEX8/wj/NR1mLqboO1HQDhXXnPEX25TUYhIuXPSO8LJKUZqle9PEC+M5R
tBuUMyeULh9hQNpzDJ0byCrgMXi+kF9UHNoF4jHKyKfUzb4+3S7uEft8Ns6WcVS2hy87ZAiBEnpk
P6dJEsvctakWcC+Uxzp8EGyGe2q+EL5pURq27iiw3qZtBwu/H2anhFXXiaNR8rHQlijuFV45+8Ax
YOnew4d4Wp5hRZUiYE7fTxkldyAgN9RyQU8SuySlG4kqI6BIdU7H7I6id33wkTKG+w/01HqGjj02
XO423peke8caDRF6tkCEfrCtxJrGLHD5+A1+Ngt8SQPvkzzSdcHZUyQoQsVezXw9VPBr2hPa9NVJ
4UkSb4Dq9ANFzaqjAAlimhi2GRgK4Dd1KeiLJLyj1LIY5IL6aiutx4zWlCzZZMW7cuXp4Fmlh2tu
hC7bKWQQWKZTxs1FtSGnJwLEQDry4SvJK3QV5CwLcO3/1uSElejIUcpnsPmor/4fyQg8y6ksFPQT
KtPLnfCv8MJE+ema4+0vwtK3+tDKoKnpCqYden6xm1dKwROOxwUU55ZVAj+BoUicKG+rrNNyrDJK
md5lQjoNXfUNuEryk/Bg2tPzMJEVmfiRIE3KHpfavvfsRlwDOkKcDAxJIsRL+sh4FuYbYIXdloYH
qO1WwoETSOoQkdQdVDCvDIHnNxol2t7HgRmRPumpJRZHRoQPQv0xCreNj9b9RJgiWJi42jYVVhE/
nAaSifQMoxVWJ/2ExCsHRcj3KP5HepC1RDDGgKXHnrlvb/Sr7024d5y3XVxw2DslDSJHOhJeK6TT
04Pxre2U4GHVqMmj+S662ACu6yuttMxQGxeZE4BnDR0PwlULZ27WqrsYTC58ENEjnmgv2GOujvvf
46CNfP+e86neQUQCoOq77xOz8kua51kcp4Qonq8n6hokDaLxDB97cXIDYcq1R7Jl1uCs+EIAJiZp
5CPRJF0tCMHUV9PMkHGcQm+Mn6512InPki46SymfGZ7Ip7A4O1mKUbMyj6CvxzzVPcxV3B669kZN
1DfWLef7n25DoUHAxGT0XlGIzRDZoaUGEk3CmMKG80yOIb+uIYJiSGPtWTsGDN4S6Yn2aAPDTr16
mZMmbBuq4W2yHRm0ovS8Rh0+8PEzTaG1Ck58leZqN0ZPuT4vaL2RTfrb+rtO5YJPurRnxoR0FReH
MEVMbBGzSGZcbSGEnlKGgUQTNjYUA97mguRcVdbtryiYAIN4q6XeW6b/v4EiQg1udhj88Px6rL1P
m+ylAHN96MAkGI+zfc/6xH/h5MOvnS7Gu8OkvvXIWyNZZ1OH4E24qUOJo4d5UsJDmDHtkQEgePWF
RqLcjlo3bSolHhJQmx+6hwHmuEUQtzKpD9qy4yLMT8NZ19oJjrWBNHIjGk8Kc/qzLnhLrLDaTy7u
r7KG8k5sHJ8Plc1U92hIZrSMvyDnhxfXIobIX5s3SdyuUo0lL11UdkE+J3TAkRP7YbNQBFl7vcgk
aLBsowzSnodNxOBOsUTbzyUERqcMPFKPPH4YV+NVlnq/VK8c6LpkNwxhJd4NR4f6UKU3XymCcHQA
aZHGF23CNCW3n19Ss65JSvOqqf7R4wNVH0PHbZzZT3KYMzTUvZq1swCFTtaADGk8DGrymU/jsffl
a9TvEVHPCytkfG4hxMsUdu/+KXKvdhEVjyVsc4G9DqLCA0Z7CcA8jUAJiogCol77F8AZq5DvSVfJ
s4JIIa1/roo2ocXmcxoJG5BDRdc3Q/ZYfKtPGLJUbpVdkKPqLOAtINOJlNzAzc/P9kmb3xt8tFxU
kNzv8WTwhYacftz325yKuPxeqiRME1A9+CqFW0wdVOflBGg5W6Rd1BMosiC93WRmZIolQi/Wko63
aphcfkFpYqpOiFfJUj6qXsW6519FOJKg+wvlUoI8VvLQXznBkgE2FrF9pVpesOUBtyMmTehn5NE2
S0i4FaJLJCioBANlUSRwIWdCFVu0NPIybCNUgKweSLr9YNqVdJuc4R/AarKi/e78mCa/EatWu3ZK
v1LqaWS7gHlI4QUYav8Z20Sr0gvu1JOwzn9WYlXR9mB0XQc2eiq26dj1XAQzcxk71st3LmoAYVwx
hAa7QwbWmH542uF319/ampUqw49vdWW+wodtOSX+WofgV3jrhk5qF9Y5xHr6KB24NwZL3CmEyH4d
5YTQ/IlVVr4UOBQ9M6J2Z5Jz6qPwf3EAmHn90Kr6/NglBW6bcatgPRTTqvmykzOIQVBaTtOqSA2r
E1mdByUwBLnnjYkI25tYdfIh1fpc+/K3DdVSR7RYZRulHjm9tCHMiFOlG/KD+U9YFkc6D8yVsCP9
rwDR02R5gF4nhSDy7+XeW0ZpLca75KpoeGb6abNWlzh0u2KADhzwrNdDToWMVPLT/0sy+XQ5sEnj
QhMKog241sTs96B04lzKvnD26QF3MJ2ufNym4PejcWSnsaUPcJZWMJ9dkupiTDo3bQQzf9RIqhy+
8c871r08PKj1Yteab6zrc+lR18nm5E0anjwTPbI+IQcYQsn/dDR5ycxkvFzOUe9QbUDe5xXrpp4f
CqQS8+T/oOqHd4sUjST98Ng9lOP838tNjqDvANXCO2+v7S5omfaXFWfaX3cAgQgnKTqvIFAIb5pM
Rc07EY0EiEBdqEyvtXPYpPiHIvzsNXz4fdc4HQsi9LpNaI6vhnpxc0sFCqNYxN+hpXUTubs42o5a
L+QBHCpqlbL/Er/B9gFMIIE7yZ2maWk7I/fRl5W7MqP0pUhqlEkAdzCouz1M3+YrPlr5AchdaadK
4UM1yI8NBmyTP6vMdIxVOLVX4U78NbUrrwrJA0Ci7u2o7XJlrwBcYLEA62oX595WWPUsmiaijArV
PKKEUXVBni9IZeCCIE3UeX9Pg99aE0/FlbZtKkF9+Sh/s1jy22957cNFx614BstsBoX7YIC15xHg
Nzq8JncDiGqtEpQ+jOuiQ/alLR87hA27I8AuKVykm3TNMP6UG7BVIBQFkYrPk4svD4iducDaW4AG
lB6HpzLwMX3dWQpldGmW9C3XAcRe1LFs85W2UsL+I1YaXFsrWhw4OjdsZz94dFhA9L1gmepgzTDk
O6ZZUvK9qqpeKJoeqelr/iPePz2Iz9M2QTqDAhwHs9n/FuYzKGnBu3Ku8JqbzJ+6WYskDsDYyPAl
FJfDE5ooXXpQzAK7lvRWyme4Zp/l+3cROocy1FcdXyzyjm7CwEMg/Ykhz/GyfBGX6Q5UwekdguL1
EmTGDj/2Weq/ntn/SOm9Gz2fbqlLcL+924mYVQuDJw0NkKgTC12EXnEZtPmSgCpt7Bp16v8IloQQ
XV7NwBpttYcyNaK2jiXuuM0nOFR/d0HrNKIVurpChx2yzonVIZCk7uAPIGPWOvjMfCNJFki9yjqe
AuDmx+0vqGNH/064hCBxaw/m6RIEdJx2c1L9fT9mXXy8MbY6bfwe0n/ekInBi35tUlhxMoC5I+nA
CFx7Xhvie6DyY1Bd9gn4bJfg1D2NTte99aGssnnZV/s8TJ/OvCW4QnxIv6D5pHu4+/609wa+ydTB
7n6ycf0Hh6DoocGzXrXnI2ZdQBmGWgRHfYrckySiSsXVzrKKTY5zcGYm9hTMEFIPi9gaFfQDQFV8
TApoSzTWyxcjtz/vVOSnvRNKYeJEg92KC1xBwN4N5oqgNzRoSiAgjlfv+u9Ogw4ppY8ioSiZisJ2
E1w+zZTx6CQDyPc2AzxoX0jpzwfsKASPt977eMblhBFvjh32Ig3ldyYaYaHA60jLlEAm7CKMYBS4
GSAndoDlUJp7A4OxFczwwnkMi4CGzvJlnrUxLZBL9X8GQpqZ4caOFxHlYwHAa77rzS+tItXnRiLq
srQ6NftPghnIDb6xZ8zrerr9OKSTCqCzN/jtUAC7TPs1LyHXVRsyb52mJwrNEkAr+ncWl84/rtJE
J45xhCyNgI/dz5WEVHNLBrGl04I+mRjYhZNFguNjiLaRySCWoTmYwdL6woedZVM3KAYbX3anLMIF
Us/YtqvjFuxSn7Ya5kGv5O6mAtTCPCghi8s26CVS02seTprNP58FcsN8osY8m8wG42M86HOAN1zA
02gAfhvLNUGhQMPBY2C9K1y+cwHD0bJy0pzNsXiYNadlRoEmMYPCUUZigTIfae+m7UP8nKg+nACq
yUWml1Abv0A2tQUpY8SvRAd7f0N7USnWfKj6UzALiK9CwzcfPvtekWYRJPTrFuEw4h5L95UPh4+b
LElZ7Nq3Hiewq4Mcnyfw2of77BxOIug7CUi0ad5aXOFhhdX8d0/Pwh9qjI8Eib4nBNLYPWrhAZJR
Hhs4yi8uyK7xiU5hlSbCUQeFSeZliYi+ALU+r+VxzPME7aMrAhrDu2MsRr6tlOHyRePh0iHUnu6v
mh2AUhBeteDyWTaGTEvqExBnUg9K/qT9Xq5OJY2OH5jC4MWEXr6Qmqy2aRtTj2DJv7/5/lZOeBHi
os6GTjbIAPXYV/VjCQ/GKQ6QrMC8P/7qdQZjLclEba54z14qlJ0LUPSINHbsQlwB0aFUj/10Auyd
DxE/aNNSacPRbwT8NgqkCQk5IMehN25Kv+3NGryeHWhi+cZSwuZrmbMxwSTbi3XXrytUWP0YokHm
pQ0kHRpoNDqhwpszULMAj34LJfmP1ntCFvPKiypCoW+xI5LIzFs4Nw5P0BG+eTUoszdUmR8TDlEK
EC0bH9/Nm7Ozkoc6sNplAzkKFfbY05eHyeEe62I/0LWntmxyM8Gk7h7G+YmjTLAu/bvHxLXW5nTI
Y5wX8VhrrS0vo+PcMAG7F8vK3iohlTu7z9Be/JXOPcYAJtEfLV6D+rvWLbZr6iW+wURu7w1oMN1Y
FFtmB+nbu2jta8hbvtihcKZMa1gzIHr2vMV23JOSJ+4gCsrtXsx1n9JDnKCMBAlMNQoRjMjCvRKy
nHjptODZ1jT2aoZ77IpXlFsi+s8OxFQFy6kOHslC1NYPI2cqJnNeMj64ukDT0Yej1PMdDDEJCKfy
/MMzlDB6XfSeA7JlJR78p0lu/YoZ7TUHLGoZh9YAZF/BvXH9RT3GFzP/Q41mcSPB3s27c8LXuEr5
fdVSIG2vOQ24EoX8ZOzMHr8+RTtoED8noXvPSdjvmpK92SwwvF1Hdjuu67h65RrwLkCcWvwG2afs
FAQmy0Dh8u0Wjeq92AYS1BlpTMoSWWsCCOTPNBcdt20Ulu77VR3sYEywJRAMEwyWn29fkJE+GP0t
ezJOvV9F/xzkkWFAgSsPq51TJQf8M//38aqTg/hrR8qIaeI2LShtJFln6WLnYvfihC/gg64ude6a
rnQEpQDPBifXRcsPa6Tfl7M71+LI3fnwJSO6Pb8RDUOhsa5LGRfKpDzuj+MR3s4bmMUFsicofZ1L
ZZWxH9p8J9f09lsCl7U2CUjD4p4mRCkcnSg7Bl9+FYQCjTIeZjvXGxfTeJTU88lxNmHGu8Zvvshg
e/ggha/2X366chMTx88AREc1PjirHkwcoRXFmqSUQd3cVtU6zv3WXSOGQeQHLJxIH4QwhskLd4EC
LNEfrYHtRlIa5y/lgLKEsO9TN8Tv8nJD18BPq6F49d0dfh3aOkCuKV1OjlrdD+z5HhdznrAHF1QH
4/JLDEueSgtg88D352AkgRk9MOhSin8kBaxPMSOx2dHatWQoy4b1+PZRmRTVReJvbmBJ4+QHOz+S
zy+ARrvANPhT9jliqzDKUSXxu0zdmOCRkYXx6jXaDKLChCBs3vRPqGz4CWXOUGmqn4ix+j9LH3iP
d9EIKCCGY6fDLrLTMe6ckHEvSF4lUPo5abJrhSl6aVItlq6kY0UJOlPds1r5Oema6AsASQK75QHD
MufdeXKPBi+Z35oHAf4tY/eD5I3SkgXIXLBFIXM5PtGOdUCaK74MpBi/7UgjzLPmk1rPVWlwaAYd
WtaAUC8KYhI1J5M22aFOCJXmYAGHh+YaGJ+tAn4HJ6L9yZlkDjQNpQgWF3S0mX2VOa2SpoifQ82V
BuJzXlkPFUtu6LFh9V+a7z9gUe/mSHPjShn5af6ScrRL9pvtrN9SNIS1iB8zGzZhgLJTXv4V0DTG
Cfi8YN/9qGSPvEsT7D8FFTgHf0CgdX6+A0Ty9B0iwpYxYt3cba1WqSe6uli4F5DQVHq55uamfH4O
tl58dosOk+IvCXZtrEjDljgcI6oyAG2iCge46pgks7JdzwGt1II5qxkZmZofKYpefVjov8ohBzct
4cSXqHml9XDsuAPs/dzQ0dnp0S9sKuDdhgoh+vzvTm/t6vd9jdoJdWN8ls+Lv+BrBbFBCioD5rWX
PklsziMpcIR7IJbcLX0Osb+7gyJgR5sxhP8M/7+ztfsB6hGn8b0YQzZbmaeFagj/e9PpyH32pYdH
kyOMC4JczhQjarjMcGekIzjQCADtPKRPSTttpHSZ6hp7gBU0oUEuRR0ugrcj78VqctawrqIaouJB
WE2j7oNeJ1CoMouiV7qw94Eel9eKbzyTZuTooSqVu7JI4YmXX7GNPvweojdc+lkqbfcDMEejcup2
UaPmGTLWqr02RVdOYfJWVgXOOoXnjbB1szKzpwRCPJxVali4LO3rU7fuuS2gJbVp6g40KpCOTvRQ
YtWMRHxyDHqJCGuPGlnXtefcYRemizKdmY9pnO39VqZE+eg9c1H+Rcy9ChcOSBzVzXDgM4f4NAzE
2GQq7m+f2TJzpH0D6f6jSCZv5yX3R60G3KaqrYxfy7OFDJflzQzX9wkKalF43v1/3yYm2iFC9sIc
pFtlImC32djNfm8yPXKfdS2jPHNRv6I1tv2Bh50pl85EIPxg6EuHFw+X+kUYVGYiT00x2023b3d+
tpVPLQxgNk6SU5XhfoGLUC7P5B7VGDbjKRtzjrTswv3BKU9HEoFDicilxn9uElwEx9hvHVBVC8MQ
DCr+vuUmIsdrHbevYW0LIzc/Zr7QS2eyCK7pJPPd4HR7yD4iT/i+2wcFycESOVx9FfGL4Dbo0KnD
wRNaul4QqFXybo+y6XrmadEDPeVtIbwh8zh+y5xKhTMRgjMPPMlV2Tmew0FH6l6HOxtFUa0C3Cnt
wwVqTimoa/pBEc7ux2k40ghwhs0v1trIFaCo/tbSLuLazgXgwNCipvLiIrNiVJsSsUxIyLlJ/AgQ
IoPzOGUEtFeMN0cpDfaZlL9N/f9ESND+hugkALb0N2b1WyLUqzdc+Ly/x6Si3KXG8leMN9aVqy7T
rPertfPIVCIQnIfoF027hKA6DyT9TUstmMexGXZ8zxDS4lyhibxoSz9HFexjMU6bJ20doSoP5MwE
eQYRu4qI1C1OWZF5RiMQUDqdt3GteQTXUZWm5DDt5Qp3jva3e/61S7L69MJhEMH90A4p5p/x6oXX
CcdInMeK7tHG4mmPWr+sO56pAgAAxmmyQbURTrw1KJDYDbWgiZk21d5szu+xVn8tn+3npIAhLa33
KNLC0Pwm+BGEpZYJsT70z1mFCxAZab5nLAqj5PDCUPc/OZiuP0sSie/BUS1PdQjDMyVrxdbAzlW1
2XA0vAOjRpXvWN69jTwwMtrmbPdjRr4ZLZx0gfZdaC2pawTd2AmGvs4EXiI0DbNBJ90em0NMZswI
jLPOY5rTyCVgfyFNIqrsDeMVorOERevZysuwEz5estPlOhrCh78JKMGt5om/LNLrANsZiG5I1CEe
H3QZcPQubg6z6trlbyjyTCvBKnwEluxZr00bt5mqh4SNeGhJ/hPiBG3gsjWTteCEUv3VBNR5Z1YP
JPzL+ammlIz9HdOKQ4N8/Bx2wEN2mY1clHQhAipNxgZ1Jj9hd5Aq1WMYg8RLkOggHz5LKWDWW2d4
QC8EEJjc25wXk99oK/Nis8e6TXB7vamhJ3iBxQ57Gj9VnXG3YXnv227skuQhvtlMA8T+n8afuveQ
3kLXJcIcvZ1Ec0DTfv2uZW2e2XOrSd6nsRw96taDzQotXwENjRxpdnFKhntlAC1gmb56pBXbU1Mg
8jOHMVIN57Op0NhZlQfMokFOM8Kc/+VK5q5WE4JnLRqXdjcxGDuVWVpXxH2v5NonySMkwPdBFS7W
gQ9mKEjIC00yXV4qtu/JmUMCiDk2mzy298hn/76oOI+46FVWfIcGXQWVaok8GI3aDRBEuOcZXa3n
uZFzGY3wpFPC6dTnm73i9aI5jdip/nyXDO3rQdP+ZNd1BtSMqxpZ6RbNdicIpTGbmAuyzgkaclnl
WbHGq/j3PrVrNAEUVqUJccNxpOxp0IC+YOdIje+OuZgS5v0Kxuxt1lFBL0n05Miewk0OnhLAGI7l
n7DNZ2gfl/bGVCMKA725ZwlJwROcJVjhqcRc1VskqAIgWoni6iiviSGEij4eV/Lp+fEiplDc+/OD
ZiS6Yhk4P/G1hEP2p3vijpI/QcCpvmtUvZaL8K27r84OgQWHHw6i7w3hTQtiqMdJLLFiC3PnC3pY
lfiFJQD1U22WiPQuwPaZGu8vJLhB0QYlRKR4Ypx/Gx9viTxY+qaLYwj7nWORLkaUFKvWgJ86Dr8Q
omUnwjLqfz7MdGhnvYtueQuv5AeLQXFX7T9wzdNX1knNYLdccMIfapQ2x2DyQ87nlHO8UyrZoW8q
UO9gRQc8Ha6BYYMDmLDhWvCoQ05tIETfHeGESKyAUt+ci3QkC692CRq9JqW774U0vRg9MD1yJinZ
Zb/igV3KsSAKBz2uHV0OXDrzMIeZAdD0Mnny0nvWKmGIz5LRc8314k90vYXYlXiwAf8g2y5tznKL
6/yPtGeVCt0zBZNdwHjhmtLNbCHLad3Na6KP3BIGwGARqBnsWPvvOavnD1JbQ4PhHYldgChdrOJZ
U9TYSG0WF8PU84FCxfSzM3kZBLigLWHNahL/ahAwXM7VyyvKtW91zccSbz+WaZPbkmszTzKaYfzH
G4DC0TRnNUbcXGNTX/E3SkX5fXYhm5LOP2wTwABXPsC8KASVeztu/o6JX8dWMdJw2r0168v5l64f
cmfXmALxEjj/PxXS/xxeAh5+hVsx4SJxaID30hIR1pyv4Fafah2AUsSDElrFAtqWr+p+gy9FQ4RV
8PK7rllN0/L6JWWv48+Zc/4erHknKGZe9o5nZerZtG63BTk6PmR0otEnOOHmLnz5MVY4Uaf6FkTx
A/fsuW1AU3vYIJbsWVNU3dn9oNSYnKpcILN5U6kGcMa8q6Zsa5YgHJoYFHCGvArWj3UuS43kRHiO
7gR2CJgOM3vD0G8AZKN1mHvx2dM3AT/UytWAJM1yB/fZwb55W+5sADtUXzFMyBLTgrUdCybLkW4R
H3AqAQHmceG4DDGkevEa+tIzxEy2jR2ev0xXRRxy/QSZq0u5k0Y7bBGDHwXZwzPMyrudTtIVTLO+
zUO6FY95f/7V67IHUP2y25bREjbV71zKaJyStPMAs/GGpGdlMjygfOzqLgUsfKJXegghFOnl2Wjt
0FUjuIiAx8dqLPILILxm8c5dH9R+8xQMvUKDddD+mnkWOgTGHg6cLc/03s+FdMSBT/RAIDxIjEh/
sH1Xbn1PaQF2BLgT8gJXSTgYGQmWGrBLrBdFTF4LpbpkRze5Ei/HNSXQdtLOx7BTqzuezrAZxw9g
ypyg0rHonLseRRLeyZXbwf9S2yquSuwe3dK1DWHL8AL56rzzTDUBtPJ29USScVSAeKcnG8m7SYsI
fwnzv7Pzj0ZNVMG8RuUEWE0PqTangPYkRZiorTyENQySIpCB5ijoBQTrZ7ZAMK14CdFrXD1lRujN
8rjoLMsRsXsdG4yl1PxLRYoSdMXCR6vjx3WF1PXdVCTD3OlHdqIplTSAq0ONoiHzNev+2RVjkEDq
/Vx5RtQTQmXklOiZkhpJr9Tq6Hr6pFm25likieqrdbqT3OitTFAj7FU3irTHdktPXkv6Vmt2Bsqc
yNnGmiPW5CfatyTKj6mDhugqPCejnO4oy88GEg6i0NVLLEWG45Wdy9TJwyIqq1ncRiq1QCxjgROt
8e8ttTAtQR48L7Z+aA+eI0xYyJjr40JcAKhBB6Wq1+2W1c9fMbhGcxwkkDzAJHL7oJgX8/sN8cst
P7/hGABms9dV7hRcTCv2MD307CkHKklJtab6JR6KL6rb38xxBJpfsZ5t8h+RBYQqGk/rMF9Ceuau
fV2MwCwWybFUu3K+zwRmLaRUfLSDbyxuLVmDxAXe60/8tEvGHgwfQ9Dqdc6zHeNRKS9qDl8mcKmh
nCwS3ttUpyB9Bpd+byzt8Canye5AdcrCMw6C+H3thQxBr4zt80tlLkmYt1QZH1TGpIq6IxHGw4op
SyYdB0nAG5Y9+x2+oR2Sq86CS755yCznCJ8a2jW7dJkNAE15cW6hOw6oZewePtCBnLnKuIPC0wRK
1ZvOeAA9+WH0HbAWJ4F8JYSgzbuU4R3O76MB9cQ5YaquW6xvkKECQarHiAGTkQjyDPY8JtXzY1cZ
DsRHmNX4YBiMiiMvmsbvrpqmL84nawAKgSolr6VUVb5fEcAtc1hpUXjsuneykytMB6WsrzZDTTGN
qjyzUe8kXJVwn6YfRrUlKG4R40cJ9gLGUIyQ/H9/g6jIUzXcIsfAxdRXbZ7nvS076RJDw9XbEmNj
VIAWOAD8b+fwX9gxy4f8ByF1zVmaw5UpkEGQgfnLIoAlpAgNs5zqotBAZYo/7YGLiLjgAdzCSMdy
a/KbEIMY+qoe8+bTepM09NRS9sG4NFMaXhzqCibS5amoEygPy+OFiruLZzAU87G9/30gKhcF0QN4
4P9La8Grmd0ZL0OGwlf6mK3RpoQW4pA/5jqDzNtOlDdzcDpaTfzDj7HTSFeEIjnWHiOwpiBvwsAd
Jy1C6IvE/adyxIHC4D6sM/Nj59q5z60BVtwByfmdFlkVNOvoRpZW4ic0RW8VEVG31fv5RAgwpoBv
qFkOxo4Y6DgaDls+SFr9S9AdU2U98p8sEE3l9d/ev3ud99Hxt3I+MG+B0ZImAEZYv2+bKskvATmz
c+VIMi7huP12uNKTVeD/HGcDPB+W9tu19Byr3MhZnDDIaf24Yt2OQ1SO102WrA7X03hiR4bkEf4v
qqBwSVo90GkOuWteayIs48ItVnhMOc2Rtu4hAFnqO2BnNSjSsmHSG9HFKhO3PIP4usBwJXwGomBi
P5ucWMqCjsej0iNjbT/RtrKkMWG+vns1H2l4uAux0Y+gvYaxpiR4pPVSEzZeJEhG8hNj+hCSd+6t
ujq48KfFiRVUsjwUkZjfDYsPjJcJ2gwZi1XpZ80tnlZjP1JCGsGqhIYpVhKc+k1bNgznyC+YMbuI
3A4qAvcZz84B910oVyDB+Zs+Szp/zmP93wiiJzC7xUKa4NollSmuNY+sLh/f8tl+TtuaJdPPxlI8
PnCg/t6ahLGQqzEc600vY0RYykAkTy3hQnoysQrnYxV+F04zWEdp8bJYKOJ0I5O5RZLrbaETdToD
Th8lUcUZ0yiIBJWLCWw028vd7SUEpl9TVh2Ius1cQulH+FM8SedqNEkCGXPDnL+do6y5WtcIgROf
qMW0Fm3ta73BRqfivsuKVT5UyR8Ludrzr6YhkWQjepjdG6RI6vp9QeRmplue+FGJU8Jn5KGqb0kN
7keIBNiULOdjYqSDc8ud4WqwvVngQdNZM5mCVaLQJUTVW6i98/erRTDxFh4aYtWcOuS+2m+HPpDD
+4m5RbxWULlOWukVQvEOU6G70/LrUkXtj8pwlPilMWsLGwvN+v0Du060mwHapso9BVIDkrTliXqp
XArPLr1kFIujJO+d+o0MirOgPvpInD5lHmZj6NEVFdRCNbMDjdbq4+c7Kv4xwBrunzDvfdNFcp/P
vyrQfreN6IbkrJKGGvaAhiG3ortPVdRVS5oYK8qvO1DaiQraO/QbJ62TANbBTQIYs+Tr4QI2gZ8h
AaXJGobXPhEvx+EQyVpgH3ZaIV5SBjy7mEJSK98kAIS/wLaQXFXpufKsTjX+gC0tHB+bco96mOzh
O+IekhIDGr2l+2QNDhxH4APQJNtemE7bAQNC8iot62o8C9J9lBLdFaYjOFD0buKyG4l3PWNfhYZM
+YhYvsN9XYPjDbdAAjgX2qRWay9iEDh9ggCHO3T1R1JDV/UyunmN29+MiCSIgQsWK36GNVYLjFPk
m1YtYvrua8OnPmF/DTNTM8iy+4pfuIG6CuJT4JSD0QHb9uhQFcWOkXy6WZo+PmrOpWMdAGOeQD9S
ljiKhNv1C9ua5YEGY0W6v7jw8KK3ynTeaX52rBsBcDOWBwwCpADFJsWmJpaJuZyLosfrLUQczX8B
YwDvmVjCbp3bCyxnr00zRbhRiLuM1Hhu/5lklLK1Z8Sn66TqkJBlx/unUi+YLU983wKFgzS/N/N5
yuwhyi/tLIitwEB2X7swQfD8KW0NsIVp7zJDqhOkS+gzchpYeMwiUgHAm4t/qdGC9Mp3VvdRRIRg
cUeHd5HY1GbsWsLRHQo9tnv7CqBEBGVBOzWe8pcqLDb0eu2mqaUXv1egT+NH5D7oyRKPe5zjGdeG
jcR03FpsupaPLyC8Fj0I4t1DX7otjOonAbxNUKXL8shmxorM0ZnlzNqW/X5IH3+TVMhtp38TDrah
5Bn8upuLTNvzcdGQC7TlERGqqRmjwc+fM7+YkTgDoGPALXHkOB/QyWzSfAlRXgyixXoV6TN+Y7hP
jKvOzI2YXq6Ulol3VcUWJiJFCa/ng+QzTkdvQvQE5lddmwQVPgMYY6og1ycrcPrI48QaqXsqRsYr
nXxHwInZPwrNH8bQgUHudLpZVWEOPIItPUDOikhJpTwg2bm34aSsblkP5fCfEj7sELUkgY70o3hy
UCKxBenEePEV14iZAWRd3xU/rM/1lwlIf2skw7xn4oV6EQLPYaLlVMFYEPV0NGV95wOlNuBMJz6u
F9lHHzuZDiECdQMog6vNROsgoNcFQadMhNNsmaI4KUxk1fPiAaQ6iFyHdQVGAGaCkDzBqqw1QPtD
fsiLcDizMQoRLTm5cC0KQJ6XOcsUwBK5fCYi48jvmNsXOFYsT4c8bAhHFh2MemQn6WgPvUon8N1I
2ukqsjaJamrpyxw2pj6LgTmJsPlwR0dVqi6a6DDDFHX5U6SH6lTBahDthjGgSxCAM1Z2r2KLj6vO
EmeYQz8FtjOskOH+VkxahbklOgg+nlrju9vcNoPfozaSkAP+0XPwrlSwk5fNItldE40CXbbFtq99
M1EPrF+JLXED4EICqlM55tYsbJ1zZrStcY58/4sSi3TUXV6w/r/ib+e2FGsRf8iVttRkJgeLXNiK
+VlRF/IJ+rDwfMpSoijbzMJKcwmV2I1crnPAdxlaK8bmqADuFP9WXLvtydlQD1zClDH09w66Gz64
/xgWpsEH/00XBxNuyJLe2KGQJnKKLXs3aKbi+MfOt4X0Cxl5jBLZvI4YKcksHgiJQxGob2B7qfV6
5KPd3JQfTZcrlFxCAzxaU1ObfjgPH5yQps2jc6aEBSwPIA7EmUzNGNs1Gjk7O8euHH7Y2JQIbkxK
rbnszkMF1DjhkYlhE4NricEise1HgnYkzsuAGlFthX0/Kekxu6agLmi0rP3xGrad8birjMy0hlin
WwjUXJOEOMNQjKhQcEtZ7QO7sl23S2Hr//ujYe+Sa1vtLqXULYNfWNt+Vf3ljFQg43uPcKBK02sJ
LhxvzKY9M0fu3ZB1DzBwzkyzco16eAu6hwaUV68F/6MmHGnaYtJ4OdpyNstDEYmTGLQrWDBeuLJB
O5f6eYGJ0B2h08mKdkU7li0Ij0ft9UmNIlG42lyik+Dew+uuCfesqmahpCHFKH7mzVRsZ29FnYtS
Wb5fF2Mr9BJF2zkAfzpD3t0kX17OS1bNPosKNkqSGMfOciCCeh5GH3RUHygKiSxgo9nQyei441Qu
g3QNJMAX8g4oZfqayIoYSgxgRv8AoD/+J+RMBzOSpQfACahRTTRQT9Ehjq9n3qgVPeQiWGjKv2cI
VBitp7J/TpVHrUzhd3C5nA0ns1wMRGXX+Drzgyecb9nJ1HZwVhQ5vlJGs/6Nkq1NE2zMRE5th/ZD
KhdxNGJUnp31ri/IRDHoziHW6uJ6Dc+DaRVtvO5UH1S1lpO31s/UeWxBW8d+BLqE84LL5+oMwknQ
Xz6W3vk1bIWoKY0Pj835Iwg+gE8zOu6tTNdm/fwBlFMIbqtD9Rf5D6IcjqUVjdR6LVUHEehplcVT
53+CtIJY1bMY5CpB7ZdqDlg0ePhQBSCFYR8cnSWjW/eOkylnChj80pxrUc75jPNmdb+sPxnalilG
o1IMNCVAApzl48EFcqe85gxsseMoh4eS2NhI/RTW2bwKr7YuIMEp/65qSHWBDWE+E3t60hl6P45e
KL/vB8Cmm7fD7k0XTSi2QjX2yuPjj9PV/x+lbKSxQKw+cTKLGdbs8iRVOKbvZzKD4BA9N2r0A8TT
c8VhXIBJCUNJ77kzOtWLl7Kg4zoqMTIfTjHyjByHUZitobQOdcpj5cjymeBVMT9Gp9LVvoARKguw
G/KUzWS8Qo0ml31zG7iccOB6QqQpa8EiDUUJsXw5W4ATK6fsFeuYuK33zsgVfcSNsz01sRTQr+gK
2tZtI5stC4xGr963Ye7yHL7WcB2VVu8BiImLvAVWfNcaNgDHsTFKoeywoReBhzLV6nBk1uUleVQO
SslUsKN8FOAPMvyOXnxD4HHINAWQVdGMfNj9lErKXIw2Za2qdKJy0lyagmVlV8HPtUB1eZ7CcsbG
QaXp5x+M7JQZac/y8rWUyDUTibXpTsq5SKN/L8urWB58O+0Pz3qqr9yyroWufzq356Vkr19sJzdN
Jnl7oK/3e+qLkeSOBOJ/KQojcQqGrAMQckiYC7JO3Vj+5BF9qQWmBD6UPPbCwJBWzQGP4/LkxGxW
zmRRSaXNfimHqwFirvjUgj//jI4f5mEVswnVtheExjayadkWKKaIphIXGck1OhMnK+R2j3Y4WvmV
iz3MI6/gk4YmDPG3meevKxcLatjujjUxtqZI4kyB7Bhvv/3M48QnzFQTnGq8a3Ym7UKb38jRtrZE
BGuabOGzW/9fVIZj7G/3lJdkhvt9X8wTswJAiWeVABi8Un7REqGy9nVyzfosAlVng8UPW58+jMiG
Gy0KJnDg8pCYNEwY0XOvfv1U8p26JHprGzUklIXpEfAjt5SKD/mEfmxD0be/mNmRQP4a47EGsapW
sfx4vbYn9X64mWXd4Z+T6JD0Vc7+yfqM8NXg1qPkuDkiqLxD4FAfKTRCnTCFwWH9FryH0N8pyyqk
gnopWsKBGAlkJfLy0mY7UL5zQb51LVNJoBEjIntqWBkES+kfvz/ZmrqLA+Y0CtF+mtv3/Q/YnC6t
uJ0s/c9Eka06+ZTS42Suoj/dPBCXMJ0EUekrs7arUaPVN2esKY69vjECpfGmPodujVQABZ1yavMF
D6fMsm9QqniHkbkAf50hyANUb4a5psjmWOMgd0z0zM1hKuRzreIhNN6RDYDmSWxIxJKBMitFLkEI
0HpNrO/wj0irZ32ziCUi3aRT1y7L9aQx4XvtwWkJMC/jVCKFg0eZJGvhXox2iOH6KL0XvQt19Anl
QyIanSOQI3ixHk2lnqH4clMTsD6nLFdIDakTnP8weqbZsFZ7ZDp7TEl8oSC+F4+QqV5BoHCFWpdm
wmfiXXBL4nAJ6Z/lJCbP7lYnMYqaKbpg2FTfn5Etn5QKGV9RbE1MFpk4bnvN+PCIgVa+0sfpBojE
qKsdf3q/OQ6cQnyTLytSZ63XwkxXz553taf9w07fwrV5d++BbvhkZaH+AhV2aLdDA7Tb48nb9Kkk
Utjoy8AdWuaRgfqS1UdCQY7KjERw86PWE/4CBGC6rqwxnFPuabUztOJM5y/neqTGD/6Os7rNMAwi
8BZbYJD+nHVjEM6w1f0z0xRYdaFx76ZL+XdY+grDfVBKfRHRsbK15r4DibR0pvCo7Lj/l6FSv0q1
DHGoenHo3Gx5FEvkshqWXvrhm9rVh0bopXiHsQWmqR5/FhXtRYtxXQnpPB+TydxIPtSPVGlYaNaL
kBhpVTs9j01fv7ZCnDxai9Wut3FCx2cqh6RF+qh6KjOHcJ3p1sPNxzBHt+THFgyzO85NxKZWyj6C
0AJ22nO2011MmxNArbSOJiNBEv6HGQK7E9BHg5MnvhLLrY02Elf1p96h8faGtTJX2dPVpOPagWf8
Hcvs007gBpbZziyxkiLPnd8mrRBOc1EzPysPOHMsYBshA5CHcG/cZFqoM5+g2vfQ56kDKB7JdMvk
Ws2MhoWSkeyUkPgzFBkSvUV9aSSZpcfNDklpg26QR1/80hOo6eimf7xIm/U+LiM02Yzi2fU+QMnc
VrXxgUissieIvFTOgrNqheRUSlUtElaEI2P5J9O1u9mNWxKXWEKJeV19l0sVGUvfKls1hsBncNY5
HvT9SqlDnov5m8QmerQzMCWUG9CAp29svkthtQZ7es+jW+87/g5M3Ak1Uzkp74pvx3KxsZaDJaqN
ntspo/hBSRkmi0U18g7DEPSzhblvcC7xcIfTgMKULCcOPKyIE0HYT+YbT3JE799zhVcib6aKO1F2
izMgqfD3TpiRl+7N8E+5kWbvwKeA3yMCqLkT9y/ddTnBAMB3WRDTVxVl9vwHvLpIM+Zq9dy55Hzu
omCg1Gej40sv9RD4oLN2VQ86Lhm3uGfcIaMyvhBDgrfJjQgtRHuab7UkfHgCQjIxxxwoWlnrz1Lr
TgPCPv7pKumI+PGxuPkWIUKzbkzGZ2m8EBDrJeXKWweO6HDJIvPDG69X2u3P6HkyL+vKmo1iI8ed
k3vtE4QOCXLrUyAcEOQ2cWBS3HlbONrRQdmp91nF7K5W7VUfxvVf99cEG7mt4MuwxxnALXrI9swr
lnUie9hQrIEiK2/yMXXVvTfuKUvqgljUq/9mwavRqQ+jN+h4ZbRVoCKF2vD29S7Ke82Lc3as7dad
FzNUlptG71jc+yQTbL0mVyiUfc/ScjkpGBAsmIt+L9KZr1dSkIWn1KM9X8hn0FleGUugyW01LeA/
+PfX3IdqPBv0BBBEgUjM/rypdDB4ULBp9eyg71jds4zN+58JIEHlMdtdqF+oDYKHGy/lk5JQUJ0o
RN7PtDBnS1afmExuII8byFT6jVlWDsjMe2rze4oEPD4uB5InpL0wWJO73GsqoKF6eEPn7OU/vZcv
IPipBgn1v7RqdspkczuFfgwvVFO2H6uRIGUcpAuPNpIprLd9EciSslZWBbVs3gcyL9WsL0Wmu3Cy
+s8GcR5sRvGMBShvNDDBEtFL1rpSeYSCU+ION7Z9gZNcbbQpS/pz2ewGSEEGuSXnbTU7U4jIlxTC
sfFy9F42wEJtyyHDMTwRH/m4dsrM2cElit4Cw2DML5N6Tuq1h4uJKO3FI5DCEapAuLNjisBdyfhg
+rdB7MAtn4yDruiHjDPGr9Dg4NCedSFJGgC6ESc7UfZXIi1S5cK3PIQZniBjZRb9WWw4c7LECeIs
c6ESUpQef9aw9vwMHop7J8ZtoERY2lcs8r41EJJxJUWcXtyF8TTvMDCMsQ17gik56RAvyjiIfo+r
9smLxy1Pvve241kiTVetS+4ALxPvaMV+wUs/LUMXFqoBX3+c4j+gP43v3NKbkIuqVagWm0xSQSjF
JpnxK7Sq9oGnMmLEZtgFx5hXxTFlWbCRfFsJ7YDcSHeWPKlQAtQtGQnbrdMn53ccs1s2JrGAKS4H
UeGY8/ya80xXnMiwiWP6AmyP0H9qe3Vfpn0ZqwugphYXZP8IgwQzR90KcCQTk9PAPL6eBMxlN1wB
eGZKN1qqhqWy51X0BB5c2Dn4HgpmOSE/cVQhAOn0GsC2Vsxwi2rlAePe2iYGh9DN7m47grKdiMGf
VzbL4LjAbx6d2IYXnafIT1+V7ODnN6Z/NRiin3g8W2OlECF3bj14ZBetXeiYBWNLW4VXBIAVcq67
Ud9yGfxF7RL1ULiv0oCflRGFUJAbXaLBGzpcK2EsV1a1ezbMsOZxmd0XUsXU4nEIN4A7s4S2zRSy
uVQiiItSYtUF5D8KUgHJbObjb9U2JWK5/6armO20mviZ4MVstO6h+VFVOYAlcW75hgySxXfnx0NE
9Gxz8ysjNaE2TBr0PdQDABGxoWjpfiRku23n20qckFGlzJasUfU9TYvkuWdRgqJKVEUj2X19CHst
yIj6Qz5uz+oQgd7fA+eGkpbGJO8zUvp0HInqXqhPNPHit4cvnL+gCBwCqGhJjolv6XPawHYwR6T3
rA10pF0VsEKpaiAyvdQrGIOFx1rw2YEX59o1xcZriSYIPsJuqtLilyFbZpUDsOEhmq1MgcgT+U7O
5N6JueiGf9i3+ldg84wW9JjqVRSCTZdgbNu2E5peCdVa+qL3yBbpM+O5nGeUMmV7RcKOetTVgfCG
rjvrTs3l05ARAMrLXLMNOc9+AGgMhr/CMsbk3tt2aC01WMOtp2DB1BoE/yfXJLDuej5tsZoOUCyS
yE6EixVf0W/URXFxKQLVr4oRNJHNCyaqSm2I5DHFL5DSTC3n/CXSkknSN1NhhxirJh7d67hE3Hay
E3V2FxoWME1NB4oH/J5yWfsr0mZ8gbYnrQZgo1N5KwVsjAjpQcwax1l4g8I3Zv3zKh4ZSOanRq6b
WGgjl0LqAsAYQsFX0DVXq0Ww0CB1Iu7nqVnmN9eqXy3XogbR26AcPQHMscrPnsgcwPcUitbb0CHd
P3MflF/H2bdsmMomyrTynEmXYiKFmehIjBHptLKsHWrfJSfBOWJcYrvLh9TBaVfHdhkljIXZxciw
peGYVNGFU4wW0zkaajJ9c82w5FHqLWVyWgrb5d0ODp3n2R5i7gZcTEumApjRsE6aVOm92yWIXkjn
wVfUVeFHAfv26JmJKSNWTYV96Z7jNss7WKBTgScxyY66aeCzBWLzKDJlI6Zpd9+Q+3gaWlmvVsS8
mfr1yauYOgYULivrlXty2ekNN9l1GSHRjx4e1h/EaQLsdgj64NFMELMigk5NqdIYTJzJxN8WLB/v
ZXiX4xFi83JDRoApWjHE7STPLbU2ScK+zraRYfzWrNvP12vV40unBzujd4kkFWxDDMLuLjq6yw26
sZhZF0h3TMJefis51fJ1iSibRj/eK/uSR2U1VVcQihbN71jKc4FAfh391RO3xsDJeG4QL8eoKkNe
ulTsjv3A8Nhfzbs01AQE9Hgr3Jkja64hSRXbfQc5C+tG/KonDz2cvyd1Gb7DOclJlU6W1yxC4vDq
du1SXS2PlAKkELdJQCCtWk29H04abckgzofXf8xFkadVacgywhAwLYw6saPBJXEB3kHA2357xtRT
wCjCWTCmIQnEjZ73Vc0iEdCJc33URvqgckXp536/RDd5cvCRNk5PaMS7ZUh/9kCa7c7ltr2j5oy8
7C4L9SAq09LKdUt9QRUT9PdgMsdOjs1Y8bxmiDTDukSkoEdL7La60mWiy+5qWZmJ5+ljTP0GgfUE
ug4X7W/gC9CrAeJMGoOn3o5K3glvYzOG7VoK0dO9tOoYUMwXjELsSkPzHqd0CpuduJXG76WBYGaI
vsawISy1JdKT6iGVqg++iOmYytK0+Cl1T9+QS0h2BJgf6+XFUwnlH2SGbf4YvnZYXqzaffTXg9RF
9u6UwM0YPcnXenKVSFXbPo1wGTG8Esc2Gf2qjDVUgLUFPpN9upxo4V1nPwriCeNTUVImh+FSWeJs
fwkG3po5j5UHDGLoFSpzfAP3Rp12ZW3jCOfr/tA8UNiJtT0g4FZlHX3Of4zXHqezhFehD0V3BeT3
0W2kVG4EkzI5SE24kXeRIXzEkd6SXDlX7xAyT+UPYLVL2rbqFxv9l4w9D5wyk/kisufe7+DyHQV7
XVQtQ+iiz9nFrP2DofygjBmPFmVIImH/01cn6NoZQdtX8o77SjqqBAfEBcbircJ6OJ4Nhbj8yFc9
/LaQhHR5qWkj/G6x5l1rqq3IUcoLngjGZeobCdfdXfxFZzAlP7rxZUwe9OTKKmHfHTiY1WPc+pIz
IVRKw525jlD5dn/Y8+aOFW8Xe1kO5g6mo/HW286dO2zIxZItPv293zcZVyCQ7zFhj0ibRniTS915
avjeYk3a+qH/Ztw/MlDoXKKHaHpcLZRMXow+I6gbicKIXCEFp8nFcAeiow6mbahXm7tZxQRx8o74
UYjs/c9YGOCV6p3T85m/L10gm+QYVmKUmGuuK6aHCVYnSRmIL+8ZbAxPkd/+OCwNkJgOgRXCOnFD
mSJOAfet3JRzqYHV1Ak6kKbMQdb+Im56/91O8er+0ICquwbiCwkDvz2k4N8YR4MGNPzlUqZgypf5
PSebTQfoa3fZcx5mDAf+u0XAY3yGVaMaD7VQj5lpblKrrGDf3ZKi0xspU351u8YRpDgdtS4WfRF+
IBzhCVuhWj9i2hjr/3H2BnuobRbJxTEJFrBw6a/y6ma9QwOihZNKR0FiwVV0VAuEsOI/aS4BlXyp
2xMQJppCeVA1qBsUiVunm2e8OPxa7MOo0DRZnupXyKr+yF/jP4Vat9mbWb99oDgKPeA7NnD7wrWY
Nr4I+ZohHsWXWCx8zM+KEb6uVr2RvW5E27Qtpg5r4h2TDEXV16TwIPCaXIgNuXCNON9Smgu8j1Lx
2QvMscvJl56ONVbhkry2UlJyXC1nThWi5J/gO0aeFESL4ZH67ow55KN2nnvnxROuf4R7cuKblYRl
nbNDpk4XQhLlnfaCqhZeHto4hVVjGS5Ix9u7uD7GVevZ15/LwXWU4YWDaNhL8CyyzzsUZiNNTPvC
opYB7izNlHSPIVfFgfrB77vEKrYQXVxn7sK6z74bDeQLYbvH76YWcrGQcZXBfjszIIIBmYCvxmMe
RlVJRdPvY8BOeELLLRycBHAzO/i75IyFuMS3aC4b9ly76ceIGUfqWJYpiqiYlq+HMNlHEcTd4AHM
rz+hT2LnCP+iZ5osg1E4wBiMSiDTKozItmeaxIFjgQoAr7VCSuiRZBte69InGgLqHcK6f1PlBQl3
PHllrjksdZkY6YM1+m7ic1lF00xDNgbVPYG4PTvtYhG+ohNRn6BudwzLyjwajRRLJQpmsXtQ95hi
fxAP+nKacTrg1HRsKFmoreQknQvhhOT24KdhY7AJPD4GT5w+H9hlLvgbqYZoUJdc+PsG5rIRZeFa
xR9eCQl5t8GoTuS6XWAyTw51FrA10MPeYUAMwe5M/iofHAtr/0rUJ5JL7Dv7X8MB0rVFuvdiofc9
Bq1fVpE1Kk1q0+ygBHPoZJioaDRcXlFvIpeaCJWYRy+cMe98sQHpz5gNt319KkLoMDl8+o5eMy3N
9EWmwObv2ycokdla9rl6bRAwoPSTEAxpIO+q9Xje1KTc4jD1F2BWgsfXtRaKEfsKp95tTfRZBQF3
r1NdgVQcRCZb+/KX/uDvGr2de75q4oflIJUnZNdjTpUyW8XWm2LIMJlUOj6v19AaASEa5gwVuTBI
8uvBP2gWgAjxiZ6DeCq2i2J9M+aXWJDhKeyko1j1o/q8F1MWqCUzjm6sO8PWbbdS3MQL+Tk/1M0p
3zrLUCrM8sUybLor1EhnknbagDXZCQZ1DdGYfre4fkLGa7/8CBw4O0jYHGuiBqSaF/Jq5plsNXPK
P7eP4RpiWTo7hwaRtnGvihx7DmJjJlIcdYDwA7+CtBG4m8CdMnpLzkSuseIjJ0HFkH1786421oTr
w0XFCCRneTPNqI/aruO2WvXFIXHP5PMD6oj95WjduENJVGdEkoCQGDGXr3LW1AcXVumAnnzGu5EK
3T5NZbg0JzEvpfVqmNPfzbgwtv4cRgizGrp12S1eSmD/957eA2g9p2KVMSTWyp39c5ePwMUZBigY
Q4svuUi2TyqvTYjcPcIcpzv+hewFJ0Il6TJKyZPgWz9chwVztEUAS4iTwuod4JprbdywNAhrCwVW
QmiqZ/XMNaqBs0PzHJ90M2CBqrQCjnZ5xQt5Z720JFXa1BOWCDQfqx1bdJfAz9Ppdod0LdYthVSl
CuEx0RSZH4TGfUN6M+jdmqMv0FhX2r7m91VhigydzJghGwAsLIzN5hEPINPDJoyqFi5HJ91AOAUs
r4sv7QZCiHH91zdxCuf27P/dzPrjRusS0kt3inx6LyVWiEvxUc9H3bQYfDrKZiia/sQ/EvJO413u
uRGYEshhtJYQBHzaNT8qIhvJALQLhIkTGLeVk85EN4WemaXSeKm+bxjQibxUjL46vfUQSdW6SRmA
rFDZ02ls5QT0A85em64M1LJjIgSemGKpHj3QU4cTUjIO7HKYQ5nhzU1a1fsW8GI0K0ApS+aQf2pv
Ro2uKuBRkkcdJ9SF/HgCO1ltz7w/CoZp9vty6V8n+onNgRjJMLziXXLB5zqJpOXFiESEcq1BsDnM
OT+zvLrRIZFgQbZqmqFnDuxEpu5XZ9F52o+OjMoPM+ma583cOWuIy3C5IHhs2amuOiXL64c37/fP
3R1ip4rrdWtqrzg5sFuCBs5iuyPpJnsdqJmS2orUuzwysdMYZUAtmp2Q977biJli9D8h2HRogMle
bKJJhpy7bdq5egvbFY+oHVUTcJTjrwWfmlwJsLMLxzyeAkmulOaUcBa6YH+doTfvSvUJYbHzyao5
qIkc4Ud3R3dgiNvTFGUgP8R/XR4XcPOHctKb3FqEIQwkOR2fvygLlKIrXHMfWH+b548LuqXgpsJ6
G6OwDwv5WLwnbEDYbnhIHZnuV1/KqU2PgWZo9S3PbsmE+b+2G76Wx92YWaveaJns08E5CJSeO6yG
xyzpcPSQ3BUF+Wo/a6wpSTwaDk4id9iyJCPOQNgVLSg3iKmFLMpGS/dntjiCiDEs+RT4IvDjGO/E
WcfAxrcC9B8qTug6pMG18U8hhqwAx6KlOF4DaaY6gd/7wY7xH2dutGVqFBWLJIFwHoSijp/KCrRH
EURfiQ4d0TlbCFvPGoX6GYelGxrOYD7huaqXJFlFm82g5327qio5IdV7/DwhqqSfy51wF3wFmbxY
NXedcKw5Y3Q5uc3kFfOyliyONllYhUa3ENgHd4BLg6z//alJvzN33MNwGTc0nn01ulK6ad8WSNmR
fBbtGh8zn126pUU1y7/POIONU5McKzRR+ebi7ybsjeQJt7OtH6hGQovLPNUqWBu8M3+0YH/M1q3w
P32IA60gtOs3cAje8UXJb4OmzGs7wVtfUY6A0ylZSUeEg3JRXMxqFpOx/b8q/YeBqHhiRCXWmX/3
CC8YFJ6uan6jizZKnYuOKGm/us8QLeYMau8ib9QtvqM7t3rM9VyJ9zCeO7RIJqRqN+7LCszsGEba
sCDMLJKrOuf3boHbhggxv0TiZRI5xSsWWNz7e+Xkv9RP0crvo3bLqO01c2LXhvvU4+6b0aIssKwA
N3sWerS16Zw0bz5OvWvlGbKZceJ/KWHq4Pc0FhNDxZSCZoribRGRU3a8j0h17TAwkBYgeBN49m81
LMJC5rsFdb79lVzxOHedVDJ5fK8smTob+SqjqQxgK5aPNSu62wIw/2l1H4LZ/DHCIeHdEk86Fuq4
pDQb9kVLpmxBOBxPCnjbOduEBs9l+Pa6i6XuK8wWjHCx8P35dATr0Dn8EY2gNPU1v7SMbu+J3j3+
L26N4s0HGh2L9gUsD0o/9kQPEWRxKszwZEUBHmxra3U8bJBfLHAVhLhz7LtaE/9iaoYCkr/SnbT2
KoH+sAz8lvTJI4QdSmWMRK1J3Mg5in3yaqH/afjL1OHG9a9e3/CdgRWzM8FFVUbmqWOxS3m+4fB5
3ttJj8RUdekg0xhIqUEdQ16PuPIchJPUoPJsV6+kamuxftG40mc1uYWe3l34K6tOprpycbU1v8sj
2gKg2ViRoqtGSiBsDIwcOQ3Zn9Rog3cjtCJM52Jai/AiO+e5Lpq9Up+Opf1hJ1LBkgoSJxuxrIIp
ENtaW5D1bedlHv2cou0aNO8ewAc88r4chkVSr3+LbLKCKGhLQlEcMpSWj6jnToAZSRmloDrTBvAL
6TyOBPA4ILj/UfJehwMyNEuIgs52LJADBIfnbLyTi33SaRpJ2mP2L/WQfMp0HXe+MjEHoGlMFptD
a2RuMk0Dfc5LTlLc/6v5h59wbG1NxU8Lfi2gw2SZUFjMbDbCl4aDxOstwOfXrAmK5h/9hDKsfBLs
tuiAt23TfqMiCP4Ys8xC5WTo+tjsCsvB2RELVZhhrY/KeP2pIroMcQTerYiBDxDYjJdFAO42/bks
aHLuettzKrsP5zgJ6+1YhRfeiOL/P5HZmIbJSo36QTVZ/uW8oVJ6hZpv5xabb47FRKToObaH45G0
c10g8W8hH4CU2Vx2KlKtJekOHMI6qjJ3CX/mdsB6ZinAiu2b+2nAP6ObDPDVTscdcYwetlAxVWML
PdkO4iE+wxmhXAj/cyqSP2I0a9lv3Mh7T8IT6xrfahEQu77yOq9MrQ+kxe0DKQercOSSJqen2t2/
2qgZD//bNk+YCTn1R+VHJOhBpBADTQUQHrstF5apoyjpddxrUQg1nE1/FyEHj5ZLQ6TzYomIcbiM
r83BUPllDQVK7BT/NI26FXZSw/LEeXBPujIa5TAi02Q5oJNejeJ4Vui7JCG2O2j2vYgWky0HvUaE
rsrJK2efeKWH8SDKC/g15h0oSoI6meF5RJPJvZwwsE/ab0Qj+g1U9K+tMfe7rAO1Cxla08xMyF12
7lr7Dzdn7DYfnXttBEZXTQA+F/jBUMkp9JWH5Vuns9ZJIFr13LEdebvdO0opUI/9P0i4jujRvVBH
vgv18Ftq8DriS1cr/ZCUG3IH6WXQmF/qwv1QqSJjilUwvR01/wnOYBNJnaYLubMZWrtyZvM6Eit8
V0MdNVgODDinfiGR5YH/PxJG31OJC5ANiGEtP7jgblmWqTU0gQiQbe5BDhfpo7rq+9d1cqCjKF+M
fG1OTT8RxklUlekHJsqZqnP26u6bUyzbYAAYwiIsKe3pXUPeHKlcUWNK+Php0GLljyv3G0e7YBY7
GHPrIh3CkTAc1gHr6IT1bvyA+U2noGz38B7bBU/j0Ii0L0KyTXlVbR8+gpAaQDg9Yv1Y2XWmcRXw
DeXxG7AgcZ3N8ySI0iCTXHXHrkmMTMTC0xl8UM1FAwK4TNGepriXFLsu2z8DIAfTh2yQUv+xnsfF
o9t7v7WI6yUy49TiFVUIoJ4WJ7GhvU6FGNAfMuQJkx+ilpk1C+Pl7GrGpILV6BTcURsbS2y1MP30
jVBSZY5wRCffI/Qsm25bIC5vas++8/J6g5bJBn1q+pVkiELIYykfUZia93vT6ss4IAjGMHM2KtkL
UQibCoknA+Bc6qwU5FsvAsyk5qqvFG6eM4JrDfCE2XybMLjM6UNzy5oKiSn2G7ZXY+2qOc65n+d9
b9BK3cO7q6/x9flJrGHklDplY95JJw+ND1kOukxNlmd8pfp1KNJNZU6Y5Lez8TCZOtvn2/aeJJX/
U5uz+YSE9n1qKTFMdwtYn6KHa034Qio5Za6b3yBLbC2mZOtZrY8afytMFwWuRJDQ1GX6YGvXeSiT
xeHv8C3RZ5uRQDodm9W4hZCxURllhZ7FBIoKykwxzepx7utSFZTBmrmdszZlxlb9xDhKVcsYB0sE
zgltCSaaAjuLuS05rMZouQtBphglRlu0ev5ZF6v1lDbBPcDxLaP9YSBWY9++iV+qJ/OHnM3P8FSp
APEDPxT8yzZqQU/hEs0gsOu8CwBflg0RDdbcUadr6Z/fahog3QVkXuFHFTvatrY+teLIZAewFW52
dYtZmTgEK3/l1AxHYuyW+QjONVEph8uaRfQetT5TNKfYPEkK7HNkcjOuMM4l7R3MbVeR+wkF5QMq
ZnIk1zZEQKIXt6uPii3/9bk9jIdReA33KzKL0CJ0pCYUtFJaewBkZ+TOFW34+9OQNxx9Q+PzMj7B
2obaMkkLWuAq5zxdgTsuv+5zk4IsT7Edy+pHd8c5voIjFxxS43EgAOoIQereHR1ac1RtXOvQQDiZ
sf6G1YiR7kw03B4m/bioUzHK11ZKwfkObk1fLcnbKSuAnYGlir0Zr75R0vi4T629HsMD0JNIPbit
mE+PON+ybGBLEVEgzbHl04e2lsE+X/D+x02RIPhfIOOjMS3PEuvGQbm1uFikQpH1Ola+ACOHjhIA
GmejyVeUWMAZUIpUqhQsuUslQ44tq6Z+Z0QguAwK6hJHShFFIDo2Zsp1k6u777PXou4YTbdTtDNx
rmAG6J4Uoo14TRbgw1XYBfWD5+3rKDzQjtw/E+LJtj4Y06XC6iHjPK2k/Q6vxHYrnntk9KjNu9bs
rdef5i9vov8CWWct0zmmao0Q7gcscmd9lVAUiWibIfjx4QTedmH0e/rqh1PUsQgzX79QXwRaauhP
BFFuJ3Nbg97C8BiZUmcFiSUzxTBKyUIrhM6K5tNdgBIFvrLswVRRV3H2K7Q7OhZbOc9WBfyK93BJ
ke521uK7QvsN6K0wmwfQnkDYz1dMj3UV86TgRS4tIZhg2d9+xAq1IX89xRXhBIOYyQBI2599CIlg
KewFBRZfWZhj/uvi/NFYKA1HPbC0qDrNheGrb2A5ss0vmxXI50aFc6WbKHs6QhWlERxeAgyL8vRj
M4bupuOmFFCS1z8vRmsLrJ1RpU3dHC6dEmzygrttQ/X/YhrBNW/nXg83ySacISvNOMp9PYWxR+NH
n4RYuvOlcH6DhNIt4X2zOv3MxcgHyDNqRXQEvLyTDMa7Q6VbNTVlBBHsGQ6U0Rkh+B11r1XEFayT
eCjcL0tD82NjZCmVQk3LOu8O3YerI1RjDhRx5naUi1KVRnRvWSPUGeUrP86dpC9fY9Gsmv31El/Z
KDWZkH5IrWm2SuJp9NdOqtBv0zi9nCkTKlXRJdWJUAnfvgAUx1aSVpY4vyZ9D/07GlA2g6q2Vp+Z
GgAgI6ckxE6qJI5yfij4I1y7ADVGSX30uLCT8nAx4V63JjbqDjjKnF5iRcc8h+vzxZbYF6qY3J5c
AcTjFqDJNjhQ0yCnGAVbm/YY1eX9wAd9Ra7bTwRXeLivIRdMxTLbH3ACPgb/+4FGWaZHbl2dwRjl
zZsutF80ll+1ielLCjGEEygS9fYAJwJfgeRDduZWVCe9JZ0Slcl98ooVh0NO8Smch9hfAuCi7vn0
abtahRFKTso33zpQ0/1XnpFMc5t53P7E0WD1qf8niuZ6MCmhAdhmE0HBWtY3WpsK4XinM/ET8iiE
IMgywQqu7cXB3b0PUCDI8h2lKRP4Jh38Vwrs1bxMaWd6mFPGiW1JVDUhA1udA4X11/oU7/rKG003
xvJ4KbTjEo56GPD0J6FnnD0ecHLm7U/aZlWXlL1Xyf0DGL/zXGh6xE/v6Na/bo64GWEDtZgO10CM
eS9mqA5ndrkV87e81wjrNfD+iaUfiYEMPNVanZciStnlcAdqy0wtkJS16MiTBNDqPWbP2l5ONdQ+
96epaW3Nl0sT5TLeR5taMCU919wOMguFPDpathxrTLJ6CD5ahSIsvf1nUdtPSjCQo4dw/bz266ZI
VvBkVDsumsURYbWZcK+d87rMt19PYk8UjZg67aoYw+lRMGBzAiVIlZuHf6YvFqwD+l9QjvO7f7SX
vf33ux9xweIyNyY+wL4hX4X5S+SlL1wpDmWC4trx+55scHWYsv6hTaDzxji+lg1vdshPUxZmtjyu
OPV8b07/UmrDMWfH8srAvdlwTUbAzG3H+UVFPVlll78Wkd5/V30ydmlDNSk24A2lCy0AdVsPagNI
DwNQmO/BD+nwjjfYgQYJMxm8ti/5bTd+CwL1fzN6Rw11Fb6rV9Ex+s9y0eu8PBeMfGWFzeJdzOIv
cRZW3QoHDDEoJEXC+suwryTPHkDPB00J7/hbu73ILtsKL7Bz8RIPPYaRZGc9+oEiCVSr7xz3k3pO
yrrw0xP6yi2988wn4es7ZDylWEqTg8MjdNeTfqqJ/bq1s3DwHxXx4N/9myRxHlpQS7dtNO4peSj/
URZJKfSq2oQ99Msm7rIRUPz99/X0FRVY8lPkQ+KkcTVjRouQwFTc7yzj69x/c49UaNLwifY29AOy
80eNyb2wvt7UB95V2vCHoLce1sj92vVXRKr3GcfH9w3PFZ/Dl4tLt6hH+Wtd6r4SG/DbzyIrNE6i
wIHa0yu8I6ohs0eRY77CIelmPE59WN06cSN7wC9leMFORR2yMpmSFQcL+I/ymv2I8pd3v75D27lk
X9N9jl1r32WX+TXCVPpbeWYHUPpUK9tZTQFd8MTRIAMXbNrDglI2bTjf4miYL7lTnzC44taBUaWb
6YKhidNuMgmLZ813dLWVEjNqxyPD42LOC+5/Ovym8J4Jw1TJDxbABC3fePsBQEpCR5CMNYI2zsGc
6Q8CTrsyQgpF+opCxjejk/lnRp/heADC1xYoe898Hz/chLKJm6Wc8Mj7w4xOkq/jlrAVymw4X+j0
hkbT5f+lbZEMCP6lfB5JR5aPZYjRrTDDDxj6Fz+8wjxOfp4aVcX7cRc3TBiu2dwkcsqIeRnYHD5s
Qo80ZWTtQXKU+fCeRMN0F7NHnZTqyKInXvhYih0HayzmMQIssYrVeB8YarfnWXLJuYSY3VwsZppv
JVWznD34rS4YrcyJNKQd2pVTgQgTneIF4wI37Fm7MoqY/ct+zPFPIHt6x6zkfAteNGCQGU671SL0
USSAdIIkRDhtXcWJ/66dggZX7BLFgUlhQFv9A/0WAfEIXR1GwD4YIC2sdyrXGVo2Dzs2gsO7tPRE
D3kmxxOSgZvR0q0OpRZct2vIYLKI3qRrr7dPSI+RRvg2yAXrPWPuu0JNa4j2V/Hmebo8HJFnAALh
PAOpz2vwpKyB9WuD385gUEz1MeTLnqcuLbbKqIgIGum1I2BU45vHrz1FzqTavMm43llta96fD340
9EHp1IXpi+4cEhFfO4IHLVMqIlQ4G3C2JHPqd2SdERFdBxD1q6uTEmuV2+a25FmWNQsujzbXH/g8
mheg/7LM27AljY1tPMG7HE/5Aryj4ZpvpsdRX9usqBsTrmsFh1K22LN0zJ36uLeG+/bHAluzQzsX
J70XJriJxkpJuRRNxrkPQJFZQb830TFQirY5Kpy+BPpa9hf9YE4PZLC2eZ2v5Al3lkpsFwfiUPte
XXn4bLLAGDJBpLRhHQoarDlTKP3r32Gj1X8xAwKa5I9q/MS8hnmxOAwfBnbIIabyPik4k5iGZhCz
W782pYMrwkooMMn9tAqd8vu8lUq7LNNAmwk3diJWKherJzLqzuqY6TanDUiMdcr8aNGobk+BQzcz
dfuy31ihjeiHRWvldhPPTkgAGnd+xIZDEujTixnRdO/5BGV5U12pC1uqeUKjKKdzRaDaLcuojin0
EIYVliSr5dfJD2KDBDn8bDg3jwrBaKY2KTPCtkKXFG/VQy+1Cqyw/hTv0dEj1f8PAQPzWRhl2Dyu
2LAAn9EgeSucHWnESsIhCV9KFGc6DDTWrPqzTUx1nyZMWZcHEKO+MK7bjLrEE4rkJNB3X4rTDTx4
W65+c9dXDe4fE8M1nnJuuFhOdyhpiatVAYtdnu5LEOzaI2cci5ea53crVWtOL0ECMdNe4P6JiICK
F36KZOn788tGges7u4uyuynxRRxL96ErEkyvapQvytYHAV8RFBm+/nt63lytKAD6LxyV7Mm/fAIp
K6glbv3BEJeAY4H8DmQhtkJw+SdRByvmxnEQxsTWyUnSpBD2PdUONLTQOwRgV9+ccL7IcC6cOd6D
hClVW4bvmtp3XOP68IrMMUfpLhjUkUujHxui0S/8UCZQmjdv108eW2wvRzv+bY5P94XVA2Z4B+fj
aTQQ/YJM3+m36tC+r2pmfUSCkXMYE1xvZQ23k3qM2C0s5/q90xTu1FKVTG4o5hXjdMKlDg3S2FWj
SPAlYNwVY79RfWu9GcWgI/MMOaccdwVBK3pgXBJvMfAKeIaHyd82uuJ/wrT4gkBfyHF2heMhKMDQ
DxRzaYvFPJ3PZ8V8RSTx7EnMw9RqDjcyI1qJTeeqg4fvfjlvf82npKdsf39Uvcip8addGz5Ov0ZZ
MBBkOwR8urQvihq8AlwTt20XTdzIKvRRl+vqht26FLUUPXdBOuUwaEeFAwZbWHnfMEp/QYRmok+Y
E92D1tD3tGng4qjX6RcTyewNlaKlDpyB/f0Lgmh6yOeKfdnfPd7iqcI663Yg9Fx3NAiWACSrhPs9
EY9IBB6vczQrhQlaGSAjEKCl9iFrX58hSwjiWlunSNnf67xZINyOBmoSl8n57zh0GWcahwUfOxbk
Rg6ygJaUqrTMpsERPBAS2yvng9Tom3aBRGpcCZaAbbeVP2oJffILfVL33jYTCX64wHqEsBzUtO+3
2kReTX+1oT/wXvOwppf4kRoubqnM5ZGm6x88YFbH8Gef+XrAZHwob8BbrgUk6RT679LyP0fGlO0y
RHs5tWKxIf5F+KJT76B+AMNov0uvXY7XayznC9KljqMiVmxtReLX8uk61rAXd6KATWQv6cmJkQW0
6T1pYk61x2IRlXV93Eg9gt5Xx7qBudbztYUAKlJsZ6WtGrg9353zuY97X0+vG9QsVo00UOHVewVq
qiZE5bNwwVZFodLSF7W7b9Y/mHMo0K4JJQYazh60zbeOsAnm3PsGB+59c5TDjN6IR23lLeDbaPV4
knX0AMuDSNqaUAfnY/zpUp3k1nJQTqTjDj5jmtJcSotGnMp8k9akn4wKFA628UvXk5wnzWTOxn78
iE492cXXKeS/CFb1+AjIv6KpTXBYYIc3mbWt6SWhQiCqcl13tYfJUMmyJ8Qwrd18+ulbPusUAyn/
D0Nm/08bF2Z2Jx0XawqsXikcVBuhqWYmGmgunkXmnYskRtMye5KzGtD3icB4UOAnTzfhBo4NSd+l
eosM89qsp17xZOQyYwQ8C/GuRac5F6kFgGrIzNVuLMJFwdmOBvYQE6uQpVr2rpRKde2FARxao3n8
wmtJyAs5zAPF5F2ovyzNOfS+5nao+FvWC6WEW50e8wYNsWKSTjYbqyg12LTAR+Z9USeboeIR44Ax
ahjkk4ukOuWP3IpOF9/CJZWqBdgxemeCmfeoEgRQDOHoCCmHY5FoiId2zxf9XoLwkg+R9u6FCZW9
SooJt3A82dJevLdGn5zXtIg5YBCKHymRj4WnZIg8ql20/r2sePIJZakyq2rIhP+Glce04dseEZOI
/FR1zbcqlAS/0fEiA6T0IkuoDdicr+MnQVlXBPaBWyjSyxymAIyho0POtLCwGi0M+T61yhAKabsw
VX0VV+y9xijGCMO/GgxL4bZ5wu7WLSi73o4HJ7CtKQRdTZHkXJ9npi0JM1sMQ22KWLtKQHEs9PTG
Czo/Uy65cGAUFaCLmUG6tojUHtvQDoWd00y6w5sePPXZ0Nz4QONCCo+jeQ/WXl0+7imWn0LpTWZF
+1aCg+HrK9Np+kl3GJtUZVbWlhwOemw/vlDOttr/xaeBJ5o/d544SU2VCMLcmXIgVipztbJ9Jkn+
tDZzB55XavgRhN76cLfnsMvzpgBgz5HbnhXM1JAM/KgnlnQQXE1nJRzi9huU47yFltj3QTxdj300
+5pYFbOexLQtbNgAtkCwohlOZMmtJqaE1/GI7bSvFHjRpAwHe5d+yexb9reg1DXbwIlyOOzszwgO
MVLEZQdqQHAphyTQ9LFcW1zMwLs1+a5qU5Q8Pg8IsSETqHaTgNA7U2EXG0DZpq2O+UTxtfqkDdCm
AQlE8r/hGmYbSjeuKYh61VkkEXGWZWTMs8CuJSjQIoCzmch8Jx23Wpj5mXmNIC2KCjIkPW6WuU4/
F+6XSY3xtey8CV9tfFqRC4NTa3NTMdKH9UyknlR8iQaSfaA1IwoaUpEddv7wYgGbHylrPKoau+j4
vs86sl8x8++6j8Uic8dxfoZth5SQwxmtpIjZkfxPVv+2I/XHwO1lK0alAo4nP0G1RinaR4XsMuwR
S+hhytJclLDVRBJPvyVhEqGHc333DiwmlMsZmVDCP1sKVx0sljw6ONMUGZzKKekcRi9BpYisld4k
9Hy6KSa3E2mx2x8Q6iHWXxX5AoaHWb8FAIP2C4r/f3FsqOTFiJnxsyqyg5XEtxhxsLlvFxch543F
AnVkIKtZGWZWn5r3MhbPax5D8UNlmzX4w4x6RRA7IU8D2tSQNdA6+5SYPZ24Kvt6qXq+7Zo80L8e
qe/LMAtcbGqlnLT11dONnNCEj1R3t5HJFVvdQ8viPGih5Lvy8iiRwb6mXSfjHolJYKH/Hq4Y4yfe
J7G2xKOFqDeTBFHeJARr/agHULob7kk6uHFf3wla9f4GlRxJiu6yPUSXpAF7x5qKGxIJVAvRwoOW
HzHK2WJvgZkH0hU8dWV8sYBGlk0LT4NJpu4e3L2IBKdU7FlHTb5RMPdNKuB2NjXxlrseb22nvEwf
fEng6lAvnSud//TtauzgeztEdtheq7hwtU0dGGhfpya8vNJsjij+JD4CQs8XoGMT4Et9A/A3S1bZ
OvNrx0nRciUfCVXeo9gLjJbMUfrZQ+pB/HTDD88ZWVXnavLsDax2+hoOsdE5dFYMswyn1QwN4eer
hIaM09mB+rD8VSBMdan7HzZHD1dbCZt3MObohIN6CeSdC5prElmkx35BCMiEuMeutwtryVVux3CP
GrAVD8j04lZjh31oZ6q6d5vAtt4TBpzgdTr/9gGmpJbvp1fPso+L5tkebuUoQNC5yQnaJuCnu+q6
yXeB07Kay06TUQU7q+BprH9B1trHPHUAjluJDyrQc8W6ONh9BjuxPW2pJdq4MwkQ2w2P2X03iVbl
AxXf9kOwQMUTUDdF1q0sXuoVe/bGNOijlaCf79aPwY0qtjQqGEc99etB3xstmx6aeaD95pafEBE2
0ekgMQVuAq8fKzxaFopgar3pZkgIH4YDFc3OPuLI6H64Cp+7/aKSNTz+tggZcSYSFhnE6SUsM9gt
bvRIq56SjURWj8czZf0pnGIdHkb9j+r3DR4+TAtBKKPZXZR2x95SfuVE/asZWBNI5gLPIiwbgDzr
5tr26VWdVZkjlANnOo+7WKgAYOcAj4gAr0eCTeFLOf+SSene8qaZl8JEHfcYEZ95YunK8FkxyMFu
CR5lA99/c4DZnZz1hWMa6N+JezY1IBj3FN16jqwcXu+RVPH65+T+bRkG8sc8wDwyid+scfKAwmOW
mcGknmAZiDMC8z7RooMvHv/hF/ed4b9iVygX04WOzWgfj00vu5xGBaPM4hM9bgHfoC7AirdcOnCs
ThX6mH6HeoLf33oZYZ1Aein5fF596Khi/3AcIGuEK6LmFWap5llVvXK2AjOGLo2rJTB7ViUW9qfJ
MPj6tIiz/DDJ2lIJ/N+FhklRZCptrk1AyEOwS4NlWoAHZi8k+0KbkWYqZkuNrU4fvmSDdK9F2s9I
zgmuP/Rkrc7NRQ6l5gT9H1TgQke1CPsanjD68G0L4ARpYRsI1l6euiWUx13V/TC2Lh4oMRqQL2ze
hy1SSDHmUBiaeu8j1x2Aolm9okxGweZZvZxkMgP/rMRCVAsNG85nfKfAavcyCTUGwswbfzYF9RBU
KgYOwQVlyZ474BgRnByj/HPqu8pC2ChW7Rd3WUOwMqPm/bQOlic0sbmQUzlR8Cl9ImHWzTGcrB7i
L1C0m5mkJhSxwv+/p1hEZHT2rzLL/vSBNGBeDLOb4kmf8MGTDWNY/46jpmb4XbBK00UqAHzLbt94
HREZD/9afER7sCcjJubO8T6Vgdzdkr/1wsELBD32oPQBbu4FDZr6G1cS10yFTerA7UZE5au+huuk
KZSpmZ0V/Zc35Jk8HQ8/zOYQ5op3U39z/j4HQoENM2POjUh0fDbqCSSZ3Lhe7OQRMyMdWCCYonl7
UE/GmtfaTkp26B8SuSa3nQeBOBpZzSg4a3avWxKlPrRYIW8fPwSoYQ/AakA5zU4ZHRXzfH9L+JQ4
GaG643CLJjJ7/h7Y63V5fpOPUut5P5/7ZDTfqX6xsk8If6K4I3BcSGiSQn2cZYMBkOPBoBjrnvj3
aXmXpUQYBe3ITb6V9YaAENE5/uAKV/olcEMsDTk9xFN318tSpCgvvYhERDAxkjjsfvrb09MpJq6m
N1gLOwpiL193Wq9jMpypsVLTd2tYfbzYaswSWUBLpTRjr+v6vYR3kYehgnz57U/LAtxZgyh7Ygms
d/VX/kQDewVfwwrf6n0N3MumCyYWZZaizn0BKB7KPRQVASFabgAL8nEVjW3FdEYQiGcLwchIBSfg
hqSUk8oRsLqqj6BOXWkTNmWSQU2c3AJf3SSG3ruDPKlbvuz2y6LEWnN6Na67YUNuZcsiZHQPEl2j
MmJcPPmiIiZ0r3fmHmWz+vfZJH1l1zjDqwkkv/c28y25xFWR+Afj8XiAnwt3RxUfJ/2deOkDv6RO
VeFP68wsp29L8VW2hGO7AqGI7UwuU6+4EHfEuDUOQsbHi3qte99SJ9JyPwZQBQcwebI9yi+kqIeJ
qm6OyQJXZL6Vg+19/3r+dyukr63Z9ShwJtvRRSn0WPISquIAhWfmILWHEvxXkn/l9b55T0Hy4UIh
1dsZN158DYHLKosOF9hcbcSoZgSY8zD+8lZVRy9mJgz053lchgtbRUvfpHSC2DY/2VU7fhWmUcPI
18nNfT/lLmZClhSDl7k2Ut6W5ASC4NG6a0D1BCfAK8DhZlUuxHx/2Xu3jQK7Nnhh2VxPA49PPf5k
xqHdF/bvVV6yTixNIwP3EAsxosxmbD+bML9P0yIHJNP6a/WnDVDU442lQaRa1w5/WVS8axoOuSDn
gKAB7IetlihtuGUpQF4a2HfBGYAld60XrUFewhS+eVtzrX4x+unt0VyCWWd5chmOsukH+XfUfkLC
HUwQDWlbjSs+EGxtjH/2vkSgL6kaY65pmlW6R5Amvif9W/v2xb+eDAfjsqucvSP0FnprAypsGsu7
F/jIjy4QEKJ0GfsfYvtaIwMNf1FUDs38jzsaDfaW4lAVPJ8jt6NzaXJjKKJXSFKxa9at/M/tWnZm
lmK7ETsSk1eVGEIACvB29tULQmY99n3Dgwj4OZXoa7xfyr/523GPAgP4kEUZRdRPmYs9WzW2d/lm
nd4kJ6sbUIPf3yJRqv6nb50xhecjkRnfPUwG3s//alkmBXDEj5NIqYvdJRDj5p09FsLL7MOodWsf
3VFnMPCF8pXPrjs1wPUqb5EJ+bzxhUzqK0K6n9hjTHsNmn1pFF0fSkUt0ZTKyBUlv+EBnjPr5e8G
fyFlI6dWCUaEyBtvoYtM159tu7L4/7z4efs/KsHYhSjVhI2RKYhpQTBNOE5YxpcC805vifYX6Kmn
mi75pLgpdc7GEiInugdmT4SkCMAhLojeeSBZHBzebnMXhekQcT40q49erwkp/Z8czGY4+MWg5BU3
5Svhr5ONNwnK/onmXGEhoa37fS2x5q/2ZU6ahfqaqejZ6R+6A4s9jOoXw0uKnwg+clOT+ncft5gd
CDnlkIbP4su7vatUq9pV8pb/u/7ex4hntNhIDVZkY0AcPNOim3KjWfSQi/VKvFWarZ30D8k9uDzn
K+XXS9RdPzWJs+ZJvUrX4Xq+9PlnoDU8VECbsisYrqUkk7Q06QZAgKxL3w2Lv0fBI36w4d96eXsg
Klf4BW5fA4xSKpWVpRO0BwqEqqHCWjRKWuZLZHBQEKZDjMcCIdKvrPgolGhVDS39FenRvvNoz5Yz
1dgBxXtpnOnQ9N2A5UNvJf2hhEUGESUsPFIW+hixvFiThFH/9swQKqWb/Gv+dAP6RzLYxEeMFeoe
E95aLCIe0z9VhhCTK88Yu/jGl0ruHHfl/8iR1YSf3hL5YuSUeN+hsh7h7nvSmp9Z5+URInYwzYYE
MNAzMe5/9Q7ze/ShE9tyy1TMh88g/N7iuoFnaEc/tw9RNWqWv0dtyAtPGR2tZ+tgu0ORLyU8dJfk
rf4gwu63ghOf/2YnEuh3pd1qXBLq/kKG5xwQQfXl1Y38mjVpF81r5cAkwFG7ORys1Ae2bwunr5Pc
K6ZsVnOjDNtgws5wWQJ83HL2JZ7LfkMbx3fc/sgFlx7eSGzouiJiNnz9rgo0jPez4OyLK5bzA8D6
myBiwts/2TpvuopqAttkdFdMGS0bfYHu5JgtzYgwTQP3KQwpbnE8ZF877C0yBC0WDwMKApqTtNum
TNz+l8wNcsqbW2ScZvHCXhHPSw3MBY6baq7rTjBEZGEPZ75F3s4YtGzgt0nBshhRAR+Xn5uUXGBk
bfFcQbKds8wU/eNtXzSRRs+BR6SPNR3b3zSahr80csbteJ2sQJOXi+NMfFj/ixKN0vnu8+I4NsQU
0MjxOG9EFtEzwqtu5SjIjH7vUTzg2OBbCGUhPdvH3SpV536k7wdLiVIu3iOJWUaKsQEEt/EUt+3+
Una/OEnSwcWaBC8WnZjCIc6ofzCGfUWRwCBWGjwr9/jL0ILo2pz//vPZcW0EDZLos0ss/aO4GvgO
jJQfV74Kn8Urd2RhG13I/achwugP02/ZKaLLIGjNUtllOwY8sl9hJai4foexQU1WQPPc3+6wMdLz
WEZPMMl599A8QRt8bYGZgAEqlfQfwLnC6JlsXrSRy55JfY66nZ4P7FLqA0StSg+rg11KQr8m3TAm
fGvzed872vUKw6JtM/jq1qu/3en/446xtAdd677/D0tZ9ToVryYaXqK18fz7ECPMzJsuL5rkvLc4
TWAoPgymeYXGCZAhFO0EAi/HeFPP6pWQ3I84wkXWEDYG72p25EJfTaKwMBXgC/7Q9/OTjmXBRXnl
nj9/vIJ8jAL5ZVU06XEHXLAeg0MUGLOrTzQia+6J0oUPO5SMQDrVayNxqSQa4Dky0ZVbY66xOE4/
7OWo0FCb3evzj7qgYIKp/xOe8R0//DeLlG+ACBiyB418FpwrG5sqcILH6bggHZTYZvMohYNCh9dQ
UDHvaH/NBMJ2AKx/yEGiN1U07lCja5KkZ2hiBothJwP1VEFLKUge3YOiU/OUQXSLsLBAavtH18E9
EZ3HMo+Dh/LLX4DQiNhARb+7B5iXmJgRVXXcGID4kG+Ni+zYiGRONPBs//8mcEkQIoOuW3ZjwEYJ
AMJk6y5asXSyUkjMrhU2/PCU3rtihmmzckLN+n6du8uD8xdtOwO1qc/dOLN7NPKFLTXQogIv6vcj
4CcMNKw94iGAFDTo7QDj3l9aJX8dnfho60eQJblIft/1QeAg9xk9gwCOGUBANjM46firVDaa+8wE
3GF2kFhcSx5gtB9f/igxGjgy7yT9eaBYra6Rq74Z6WcLgAtEHo9E+O2wVB2FWVfH+Lfcwb7FcmX3
kLId1CQ2XrC0VEmVS73vK18J7IiaikfHLn8Ii+wZnEj5T0UEtyiP08zhzeWiEteMmzfItIKMCiOG
yEcPD5qtlLXEvKnbUqVvG3L6VjoMWm4ZlsEm0f0NX4gpEkb1ETKePikbc1GS312knYfEngf8r+Sp
MoIqEHK3ZDcTXqUgxJIYfp3F/1GCAFn5zFUbxYzfTr36euiuDp063bHql8X3nS4XxSaMM68+EucA
Okqz0D6NT7FDsuiewAZcc/2mhiEYWSQUQPHbWUK7euLEHSfPEVXRTK0dlP4F4wYIiheblKrMysxm
k9UeK2J+AYJ69vFR3iShMKjZ8iI/2RGcl0GZzJFCQB+STHTdNwfzmR0NZyQAKbEpoX/COFLzvmeg
oOQGDELB15X+2EWsaGkxEDabqf/tlFcI+tay1UoxrH/1MjZbwTDkzcNYovp1lKx8wi/sDMi7vzQD
ntA+xmaBx7cTJE2/b1zxaHwBJ4IEEIze7mDYvzL5d9TRnXtWKoCcBvmI28G0N8rQ9GUrIBqGQodX
4+98Xn9VAMgWf6KB8r8eFauHSax7cGsIezUAbYxhepkviHnfPnOx8VnWYWikFB57v4aqNAgfc9jQ
ZMI2QtoPHD+ioc8N5Y/Xi46hXhMAIxu77IX5tg3ZALfpxBkt1U7Dp3SI1/DLy1Ep48OXH7r+Bn0p
+bPes/lGP+hudB9Fw3dq+8IdxtSaB5k/Fwofy1T89L9oIAr4xCQ2KgXxQJa1np+J31VAVCUMZKG4
XJxqU2ZgS23JK5To0q3wi99oDFnOEsJXyyvb+g3yJw9NmD6WASd6ypK4LPj3AlJmvRZ9cOjspPNx
wnAd0ZWpwJcMD4LPV77zpveCF2r156OZFxkevLZZuMnmv7kVFVd9nY6UBUARZH/VEg/WtlxhZZqN
/PR7zR2YfuC6AF1WO7SCifi1ynYC8spgRQwyeKh6oU3r1PLSwBhUV+9H2RySMECThataLc/Nvdes
5cMNhdxsIkOGP7mittl+2iU8VbvJVgB6flZwGso91HDL6aT1TSHQgg+fz+bkx5OG46rBCl8hyZQm
TEdlb5LGXpbVeMOaoljpUvEc6IpBLVbKGSd+NpZ1wBQxvSTTOkdCzPadU0to3VRBeKdS47sp7QLb
5jEvWNVW24Mn2SF+XDii4oCKC4Hptj/W4t3J/2jHLvIo5zE+9c1u/XYXUarzf+Zooe4ew9HSjPx1
IC6oT1H7aAFaoo6OLel0OKG44En/bva+woceXLbs/qyjNvDrAxBIBRm9uU+L8RxR0WjMz7xbsW2z
DbbIYElFlmik4lz2gyX/TtQKR3cagKJYuNkxGlY1I4CFlCOhcQ2JJsslcaG5+ZVX+LhhU8NiJeyI
n1S+DLFxjfKuHRTFr1dXUOtqH5n6jbG9enbVSVYQmzwXZmsmIWk/nnibvCO0nyUspQaSp3NN9Czw
2soa2O0i/vXnz4TzBCCuosls3zFwttUg6ERymg07clc6+rihoE34w/yLJ0pRThUCQmb/QLp1NZwM
Ig+gYcMYx7EMTJXNSJtdCtoGPqSeVHAM/idYbQV3Q9F57PmMH5XdlJrloe3iFoTnNrytLJM2cCyU
g4lGY7Avws9Y+2x1CCNTKXsEyXUaqB/hu+OI2kX7Y0QN0U2UIbQWzKzLPE2Px9WLG4rOj0k2JjYD
w2YuR7e268wqPO1sLQeug6vqYLmawP2es2LWEWsKyFzIZFEFebgP0iOHItr5gI5Jx28le0S781nd
nuqiWBANIBcTGGHJW18Q8diCiSHh1Yza/EC3BJ3RF6YjG3nY+P5cmedO4+waWz5ENjrZtBE/BH3R
l8Ypv/uar3Ono3nd5a+8k7njCwIS2ZFTcmnOzhDv8oWN8u1c/AFQz15WsBbUB7udg5UFUNMViIvQ
PZxklgOLkhXt+nAnqCIyt0wPFQdhZwyghcr0+MBC9UdphjA/C7u4X6pQcF4vGrWhP/jPRF6YVcXw
ewkK6DUnT+1cXs2uvpYvZxdgu8K/zmz9q4L6GadRdoSniWM0LsISw/s+nLuMM2ZCcsbBkEckv73p
b29m5eZP+sSWK1aMs5mut4wYLrIrb7DBi6GxtgbUbzbRhRk3zm2VOQ8rDKZgqj1K7abeboHWaFZ1
r3nDL9PkcGCh22XpQlAkuUjrV5H/3e7lUok+0X6RINpZrunDjwCCIrQnMd68Rs9i03T9AbCQQZ79
IDfSCjPKBR4kXTkQPuTL6N43pUKcI6BSVu6WWzz5WKUj5WTj0Ndsxq3Y3jrumGW/hMXHcZrLl7SD
ky+gG/GFC/e9JosTwQPUN8rBI5f5SAVTuQCrSZVQH909D4cPPlzlpN5U+fgLpE69FIEpPtZZepsM
ZSgMP8Fl/Dy71wOWf2uKvFJM6YZVMI6hLxREfhlAEnNZTg8DxuiZ6ULKshqcbFNDh4W+kyjn/tG/
aJylV5hdaGR34dz2lUeOEP4LGz7skgBM7HFBP+9j4rsvrzTux9CX6yz6JA7WVc/uIhe58KsRTtNp
NvnWci8MyC3LWhNGn/1uwwna6RdO/ZTfE4SJkvAiMMbihSIur9RfoTM1lJQUsLhFZOgg5mfDpLCZ
o7CTrCZyDi6NoWdscSp0uPWG3nt0lrJAqUD35uQ8mKvlZTgO8hwLTBCewOnWoDgDsVZUmIyyGwEH
4eucwKAz0CrAvKzYovtyzRw64ILME4BwMogm+PjJ/AkVP2GUf9f/QYAM3KNMMTthEZfPNP4/C9bW
UGM7DWlMEL4+OJsM4Ah4x9OOu7AtpSCZOIOhvBPT4smDGIyzeZyHmR9ZlqsiACk5UTzOcM3GC1yX
LJGY3O+QMw8TghbmIqD+CKONijmaJN2ClsLq+VQy67ChdXUopOyxzairxjQ8GbRA9jqcGru/z1Ku
F0aE4UmobX8+3UhZCH6Qbbw7HPrcm4reMZxxqlryM+n5O1/BnCHT+HlFb18umpBfb5q7VX+4OGIn
0dXBCcHzMZvohA1nBMGNV9r01v1CzE3xAx2I5wRHpLGrskp+hrwvItQDgwcsE2hYAWqDrv2jexHi
2G3jxQf0mpPWTAq8SXiCZTIRxnl1ZMlmMcSorvl6RxtvnEaklg0wn61NEPaqbKVFKYzUaaK0a+qY
zo+Euu2q8lHYxZcbnewrYFtVFNngBVhbwC0jIZaCIV8ecWAfbvdDqPwDw9Ou7hgS1pWKgR2XOvNy
21Y3bFag78Q2jVpZzqZdtJLJpDXhqI3TY1erW2YXi4QhfGx+/PIGtALFatY0V5BwyE0sdtRK1MU2
eDMrkU3Y2rhqo9FX4yiUURvBU8RBPX0SpdDGnmNqz5vMBhP0Kpl1p7I7WMqfC8AhrNjV06IkXf3+
QCeouHAbbq3fpqAuKqZAPgCMrUmoERGn8dZfK2Tz36DCsJbYDQdHcNRxiYqxX1kMqQzRE27ylJcq
QgEPv2ojp/IC4P3Yl70U1lm99ZPv9Nc8gTXRe2fK+IXyhQf2KUuejWHabG9VtfvHK4yZVuogaHEy
VrbpEWbtUqUfk9KTbE6N/KDU9GvRV3Mfl+R8cFNhyxfxPDo0AlIIlcPE6c+Ac9/5J+SJTiKMNWjE
aaC1luTpnKk21/161SfY8nVLbGhfdUi2UG05XRRMQrgmcbvVCODRpWFoh+/aCH9vJ4gk5YpnY+dg
/UMO52i6hRqjRwzUVigkToo3BbzPFZb8GLCVe5Z1HkojJGvcN8GURzW53vSMQ5BgkUgFCsSqgGHo
9jCtAuJTQdgIusjNnFBjPgGswkUeOsMTfkuka6WbJ7Qc3m1BqwNIzQBbZ94td/HOUoaJZ/hv42Ia
88XefSyCl8Ovy1f1hASnD/+iYrIjLDX+prM9ethmiKLWf0/+6yktlMg8t9FLTiwTxTJcetiNT+tS
dQIuNjNWUelOd0EjRq2FL1Ee4PN7Prgj426zxSlSrnoV1TBSQAdwjyVZea4mBqWYJrz7b9TxmTI+
8LE6u87GC6w4Lymvv+IwkuXd3vFmG11HYfeXUfgjBLukr1eGJ2S6z2RGJ2xFnOJfV5LJgc0BGDY3
me3pcxeqq4MMQPWTVpQpMSJfOgpAALjK0TdDp6B1Gg9H7Nh3WH4fNun1omTiBP1tv1/tsB6kDmUp
OlG9d0RJNIJYoqiZWDK2S/RTUr9Ku53CkJKMPW7FF+tkZvdqLHG2Q0cpqGOlZZGnQ8nf8GIdqufv
KgLPldZZ3JVAAH5ndu+yPCmpJaVpwmbapDO67xZ6veTGHmuNM/FjF8s28ibgN6TWtPpl7mBw80H9
w/disaN3RUebkPqU8fLxPrqr4Zuc1m7sJbx1tPENHmwcGVn3dobA7jXhS8PueLvrAwI+uPeYDcBP
R+IbrsnzMkPAipzrI6ml8GZzxYFnlUmyRA7Y4dgnJqSvvpb9qybDC8l3IqSektLoYg/CLWHNzzlQ
Dsy157hCVQDiO3/LAH6RJz/mMbHhROTtgNL4DlNey4JXk0RL8KWGVF6HnassD1fy2p5//MZb9EHc
z29oiSoeyb/OFqNFuIC9bglDrOsWUZhF3XkM1UX9jqEYsl2WSF8j3N/lHpR4zw0Q4P4TISfRJq41
fntcwqYA2zLiEB7vKvR24aGRdqfVUgQ2SAhXpJMxigbiI4RNkxVyUp5SrJhgYEDN1FrQL1dn4dIb
7zuqoCdzDedK01IVp4LuYiWOjgnFi6ExBtUzeNobXr+9ZkdykN8MDPnGK8fb/y/wJgwNhQyZ2nxE
YWxUgOTYJBRLm4cQBz1ypM9SJLdbGnhy0CQbpCL0dDCKN+d8rGrcyWumvh4NcvyBQYq2jRK4lAHA
VE3d20suFkIHB3dWiZL+qY+jGWG1aUYfUDRPQlu51oqIhdvmuBASKpvDQadTfgL1udAG/8Wwq5Rg
IBLUMMtYfpK6lkR0VqwN62yXKpmCEsCRspmtvGgWVl4YSol3hK4WHIRIzqEy5Dj10dIGnJpv6uyg
SlkhGuE0rEceaOGVFYRswqDuvDp2HGzVjtC/eU6fy+2e6zxQmLPVJy6MuePdUHWhD2TVMspIrRmP
AoHvRZu62HnTx9L2dqoOrOkkFpjZoo+4gtjyGfWf7hFHiR95k7wA3Ob9gwEvgsJ5Af6VrdP8EEQ9
+vZQsLwo7Rw1/8bbv8AblFtOxkDpJXK+roHLPy8sWl19DO05l0yRRr4B8bzCCSVdISIS2TbL7UTh
14MwSkKyAxXMflU7BH6GM27+rVC3yLGSKNe0/qM6v2fdRXMlM34ns6RCdcSYW2vYWXbGzrrYmQhk
dLRvbosy6Ib4b2u8Wvmxb/PUcl1Z7FsRQpaso7WwxGHq37+NyqaeWqFXo8iTgFIL8Z2kfV/W/Ysc
VgjHiPynrC0V5W4/KinX1hIM9yMdTH4blipmUA6gRBDMe8cj+QlzITqpqXqHxGWZp/PRyhNxrkFn
20lC4tBOPPVWcZE8U30n6r+1ulGkRsktwAknVcQCE5IrBX1A4Nx5g9vO6fHfQ9mKw7ih5/mixLOW
I9VBn7l+R8EK/tGP+mdIwDhXx01bu4uE4echJiQEV0IW4AZmdxFZApY/R6qlem5yOXAIYvgNDVv9
2Uvzu0MDnMyImUpJiKhbtrN6r7aQpFPM7AK044w5jQh0aEp6Bh47GFqP1ttUMGegUPTQm/dZ4T7Z
ETGHquWP5l1Ci0FimpCCyZy+XkOogonlrG+NFGZBdGTf10PourXxZXXC+AcWFNopVzAokHoK58Ek
BiBkWoveDdhJwGTY8eLCDm951crg/BfRVugaBPLTExKXLg8aJwYAAEzLQ7i2IrVctmHixKCYbf6i
trGthP+6FOE1HRhNzkOif322BXN4RVIu5fv5PT2Kg8q+MRAWWEEd8hH9y8qlaFg76qC5O8zE4R1n
Tiw8aCdwNsOK7++MuoeXgs/0CwQ1T4cWoNK/XTsUKKQVFhTqKXSbpwQFWkgdmngNEeHxfH4QT+wT
PoYAyiiiZtIaD0prE29fIJynP9jYZXFjiWz8KMkSnKCN6CenFmNU9jgjmt+2fQHDvxEyxhcSGcrn
6MFZeylbLjVPDViLk+O7r36BiPdnDuaEP1RYUv/xed/F2sxtuGN70C3EDk9Qe0nJerfubMtei6Xo
4XZRDIBi41DXbMdy/vqPyZ6HoN+R+q2wUSkTX2pG6zwKaC90GEPsRznlT3co2SyyRl5bb+eLlQIx
zijFC7q/F7m9/CaMOF8nO91ezdD39/LoCaNBFbwEyuAHSl2/XhMQZZ8KVZzOgUdiqoKv2P4SSB4h
6kpg5AyPQORitP8hbPmoKoruQtb/K/TpssX+j18adYPW+JXPYBhSqhIZDoRhQEuraDaqNjLdcInA
qDHaiclKbwa4MZiaquYyw8aenCJoqgEO4RWClkwF70e0UhpAtFNr0H2R8YHaTJ1j1V0vj0QfMoa1
RUWITKCzk0QSv8IJCQlY8Jgy55RfrssQD45KY77Zq9XX8PGWc57MnV229yjTILps/UAtzUDjUbXf
BrQ8cuAJzrKxv76ILwFlylGcPCMqjrShMZ3sYeKoAMvF0KvejZcC/Lhsza+0J+vuT1bzMc3z9tNN
V26jlAxRZB/V9rcCb0Ruv7b0kuUhUv3XCaab8saYNZg1KnhRmH0ATo8wHxtw9mGK8zNan+5xHtXl
CXRR4MhztIs2YhYMqjZP1yBk8YPUVe1GMyKTjLElwgc7BXS3jf31A25e+JxUkuBOaFlJZlWv+9Kp
ejcIkBwSEsay28QUVGZOhSnMRVmyOOdZlzLEG9dh6W9V/f+7rXrZQye6u3wy7td1HpolFiVoUrAZ
k/peX2mJndcWbTHEKzlOlSxMvlyXYQqkLbdoXrrYltLAQeIxj9lqkj8SQ2H1dTmncp/QuJUVKZDI
UXCSq39tXktVqQU/dXni/UIPfB7K4pf+VS4sq+CHRSGyzmBf5uOwkF1lSAvPzYSdDCWnapDmrLqR
AkqamOBW0+eyeyPt3Cx6ak3jGqNCSwnvkX75+DJaxoAzDrlnB+Bn89YWiJmazdr+IEE7ajS3pVHt
/9D8qGFEYk6TcbbrW9IL3RZ9PI/vNFQr6mXkXfiRsu2wyx8TSHfakETY+fPLW4U/DiTALcvpcyLc
qOAJwhmJXX7ZCZndScVI7QTyKE1ZufV2A9G/qo6QpOllj8G4V9ypCrSsPF4Afien6CiVYejP8FCB
82iFFMeGcSyxluIGmbAJkNbCXuWirvXnfGRiTkNU1FnjkHHngr2VPz5KbogP2d1NifWuIixb+A/q
k7KmJl//w3GdE9QECL5Y/oZ6Zbw7gaw9glQUDV4JEWKTieauk0VWPcGUetu9UcTqM2fPzRi05DHI
HzWM9Mt8sxfSK03CMtBP/mFyRsoLnxLo+E5fpzOciQv/xGnJDJilJyT9mQlCxMQkeAYE2Mxp2y0Y
uMRqd5n+23oFUKSj/cvoLAQjLqChNj92sxdq65nVvbtP24o15ZwWjRr1BRIaF7TZwLgMYZDwCTZh
+qzrcLWbqhASNTZLutd1D5FhqW0y0pKjPMHSQVESlHsi75oPZIer++dRrVQOL7wiP42xX32vruRj
H9WqPGWRE24lKz9GCOn6oNOHN+1RR19SOMEQ8FlXBk+sGbQXs++q8Jxu7fmb2si/IdgtockxP1wy
MyBuQ2F80VJh3pt+GMZ+uj4B7diQzuWFhntzRzha3q+JjyimnpoaxIxTPGFJnOOd/qF43lyKCNde
FkRAlZCGnlFIS6JF72jr+mUGWE7LO83hCAsIXVjaic0QMgli3P9ckKgUA7vUBoi4Jm4qlnDwhc/T
BrJz8FOzoQq/vb/zA4EAtwjRiA9VHoaEr6jO5K361R5nG4iRZ0r0zs9QbqpYUdiHV5hdCSxAcye0
5DTuWLnMYxWrF2+fv5jAhBFEOZdtut8Ah1qtufILnvkbq8jt+kn9S/I161GAN46YzC63BAFl5LIp
5Ogwt/30atyVt0/13ePqlb7SbE/T2PkyfeJeioHFQ66CI+KdkbibcVvoOwsaPN/nnLSq69J5f8Io
k1OkUGKerboWBTlaS7R5weBI3/gCA+j/WA+OQrG6xhWALOWKgPi1WM4f8yJw0twknf9yD+zPgkMV
axAA9hZEprNykEWmBLSyYf0nDtBq6mq94nEGpfahVRdQacvl5nKU9V6TjEUXscYkQrwVex62HxlL
latki4WllUXNDttDRBeDfZNP+PDbeQe8GzZY91CEhudDw2Zwc1Vvt+s0XmELd8LeP9/yoktBEGbC
pEt/C/lL7OywnobzyUedjphk6AUGJ7LfDJSxUNZmski1QacLKq7aGRtNu0eafEzZAeScAl0jhwoC
3QEpm2Ji0TKzN0+JcB6DEo0OBux0T8ReOU5julKgl8NYyYuyf/Wg17AFMjX1WI/hXnV8VFNIAZer
7zQDMAXQH/JljRc/lSAfCXjZea84hp5Nq6t0sb+4xDuJpvIGlhrBn3qpf2am0hliwVsY5Yj7qqLS
HtcWGE46+DbqxPvPh/BDz8nNWzzuONoJp1RvD18f4b67AVkvIaUsU0/xknpieiBgEdLF2oL+hPUA
HVoH4cOiRbm8TSb143ENf6At7usXnjpFgDYahqY5Xe0XRPCLytmTDIeT+YPm64Tpas4xiH6/ix8C
Irs4hh9rxMdUxS6z+XoazSXghG+zgiTo5ryZjkrRrCM5BtkwFXJEHfoDW16PdhptWaCldad5kW4m
kFovTjiNre/SWuO5CcZUpawFN5F7DTVeXexci6LrKMpe4l6cP2lxj+zSOephQIQX3nFYeFrOoJ+w
ymA17uxeqPWyHbSrefCDgzKz0UgZ6Mx5s0XTH7wIZzLKFM5gAi11aVvgESmFmRvHZ+ONGthvi7Un
TUxuGJLa5B4+DlreLT1YkGHiNN0mTwM9W57il11SdGWPIzktO6xp6l+YWqGofZrfLxpM3UDnGy7b
ML+7aSXUC2Qh8STPjEXv9A/y5us3oimndrFXL2mtGFzwlwP/d5aOWhnNCO8377HHmWtpUqa4M8aN
qjrxYxDe2IVl7IGrCS93J1hqQ1O3RidlKLUVo7Jw6yaDiAf/tbpEF/xJ095jRb+KaA+0Xlv8rVo+
edPPFaSwDkAxlFHVReJechq3Tm6RExffwsiP/G8iudtbCXO40YslRa7D2ZItFZ9045Xxt5ZQ4Hb3
1F5uPhWP5bS+hDiy8LthLhWdEIXTlt5B+SLXno6jcZK2FeAeRDNb7GQqTBHMnYqUIIi6+1pNsM/l
r4d6bqisVkJWABoPDpwdR/NPCG7H+OedXwoV0kuebsxqTZ359tj0OkV5i6PobgS65Xe8E0L1SZCF
y8LdAC7CzqFrAN/Q+GI806plsiOSRvFXB+qSgpRKqIMBHwSy1ER9zICZPqrmNoCTLZ6qxbGCL8Ub
gL6ciHHVWx1jc3ILhWHWkgdrPceT2YssxDLSw1DgJVEyoD9n7mep6ppNUgkwF6yMBsUzX39TyGUs
ihjf1eTfB2iV2WtGCUyx3HUYPFcBCapJywcLUlHbdxtTx0v/FFaLZRcmo4VhcZAhAVExRwovN9+X
weIbmtKwjhQBikcJyEGM8UrIfP/RR9BPbCutbinDvM7FnSC1wN3A+diuRctXVciEUDFABVOn/2mc
ygGYAzKbG4eEmdCpaD5i1SN71I/kIAoxpKwON0QtWZ+FYteu34uZf7jIkbLkYxgdlyBnlm0ehIVe
vlsWhesfdxyeYe+vthqIW/qxjMe3uOOmOliliMYqw2ugxgACUr7Ir/K2g8uYttV+8ud/97PsAt9H
H6dInIp84jQuXAn+k4M1Yv+0yEP9UFqVY+XpKeE1n+pGQjzSOzeVTzBKAkHC32ftlCmxnNTGcnUA
gcjohrj5fS44VoBFhmV5dDxCaQaEFzDCiaDBz7doHKf2rjsRzK67qHbHpaeUjT1mIfi6NDQOpvXL
rvKJ7HsDPUAiFQvolxXemqNQo5Zv/VATQxW/S5NOU75ANW3bSE1e1m6WghdV2bScs8eAnfs7/gHJ
v9tVVRX7viwKG/XTgP3AFklyT1bvMGCYRysII/hX0FhAsyRMx+w116Io6r6n4f+1ZTdGwjBFHTD6
wK19YXFiA6lhj61Oo78Sb3W296SjSYNtGeUYAGX4FMuaqCO5zc3/XP4eZv3wsPWdMlvaKsb9O07I
b3xf2WGtvK0q6yVi+JZVJTq4wyoG7XbJyP1GQXf1aCr1Pm/lEq9iWdToJYtgRbOm2cusowiDusWR
Vnd76k0EpPJKW3xGTCZ93NlUXyqsjNnkN223DtOnJwlepuMefE3HxuCtNtgjgyzU7XAT2fpB7R+3
JFiLAaBPvNKo0FoZ95tNhzr3sa5BZBjFs7IrPPaiO5lmML1NKPGSaejt4eHU5SYCUrg/MJB2/O+F
OQAnz68s4LYv0qUlIU+P+5DNNKNz3/1mZTUJRmVAq4JXEe1dhp6Mjuy1Y/Ojw8aIUJupKh3nXW0I
LDd7OE2NcgcXQIPND/5Go/xg/W11PqhUo3i8C/vW8suo5ZTjVh248BuHoDQlLNIBKajPoU5zmyP0
fObnF1luaTN4l1cN00NA8L6fi6bk5fCxjDi/yO/5+aRekIO6+AKFkYDynRZEil0H7xOUS/J3rEkA
syLeEFAKouYFDQJ3wWAdeolamHoYT/3TAJ3NSMPFZz+teMlOT91dMZowpYhOrWnzzvYhn6o/agXJ
uukU3kyVNj1L+NDaRt+E9A3tiH+TOlBzMiE8hdZYHzRtSkheWFirZXUzIU5Arx39Lubp4172V1W2
himkO8wz6ajcovmhs3gXT598oRb2/e4wMKT1J9vjamgPuG//op8cJnXNDWqsa4922eMqe3gvxiGd
kGa0oeSeJ2DBPaXmxBXdwJ+9MSqrTICCM0l5H93tat4VABvF9C5Y2pY3UOEKacgi0f4o9lLae3T4
aqsfxmBxfxgIZrGCncJGYGgnpGFxbwaq25hLtHXTH/9awu+A852F1kPTPmVVb8qUJYSO09XcNvmK
KFwIgSrvWpbBQZgG4ILgykmARsHTkX9Eo2oTelT0vny39MRCSoN2lSzLpRTlGsBB1xOcZ587KZLA
2iXXhwu/oCDOlAzuHalInTn/A3I0tyASQydy6d0QqD7zoGUGqNNH0J4NCcw2IpFjMBNGuJfkM7jI
nwKG/NnLhi15ctmOVLRumVY6jay53zJYc73VWg6j/8avueHKIvU68YEGLEs734+S4RiXK9h6arXx
DqYTU43/mb3QGDalKsQ06w+y4kgYVx7Zct33J7mrRCa0YwArc5lsM6rzasUptuLrh3pQc3ywGTr8
vnzeiAtgNolTWwpJmUCGaoh/tBlfiYUafI/xSEx+9iVhDdv0jMg4U0TZEjm+UOjdAWv6EKFsp4aH
r++UDQ6bBqE2olZfTv1ZzIUKyiOgu/kfi2mUutrBn+4/fL/v97a/1ykAPfx6HTCpHvCSK6kWshTV
Inxdvesm6uGN6lhln1SGLe1ccKevqAFBdE5Lf0ogQ7v9SM6Y3R/vkftY6v3f5d1whLJ6pyXvLecD
psFdiMdOUrkfmobo+fNJa4sMQROnQn8z1TJZzyjLHgNvOySl92vy68nZl8d0iK45UbI8S04jx0qj
NAqS1yre1UCfWG6ZuwIygNgmWwuOTE/WmU6TPntyqc3bBy2vR+usI79JLAcio459nQpf1pfzjbCn
C0QqXBzP/zBfhA4F68Xy1zlfwuKCHjVBlnPUuMRrwF+b9PmH29WSANjgOqMjkfu2dBCBTQBlVpJt
6FKJ4zrdNBh4va7oYKpf2gtLc5JhXD34thdHF81I3VtaUv+cItGOugCZM3Y8EA8n1GnT0nEPzkQI
pyaFcs201OZxA3Ghjp7pBpXlE1dqHAHVljKBtki5wPW3HKMA1HM9VzbchyNq84Rd7cT4nvDf6Fon
Ecq3f8ZU83GlSnhPJQtmpGRPZsYK2yatLKYcJTmERCCY+WRNZWLU6GVVej8ffMDP3zkMp+SGDVfg
CkEaB8KK2JBUmfouT3nttBG6OGEv0GNMyfQXs4zopf1XiElYO3xsbm9csGWf09+W0Z72azE2AsLY
Sa4lTLor1fgkOfYaesP8T03ALeXgZl/1Vr2jK0JMQut+ovBQmIEc5BvCK0qtb+XYHggppalWpsfL
d3PBQocHzbJ1OEsmiIxNqCnqFE7KMi/Lhldlyj9ZUgCb5YOEYYq/NkX0i/ST5i0FFmvqZeoYP21d
ZVvWnQzZnCNDj6pZJqga8xo+7ioptg6Y+q1m99GSpO++nMoTXouhy/rFeVijUoMkDtEUZTUatY4+
aLzm+8J8hSE3vBQy4rveo8z5FybC95x/YfSGEQoTKPFZuItSaB9UjP2oOJqNFdD9l437gv9wLZuO
q1c/BNKJgdoLTQHy/wbWv03P6jy/Nc10yNypplTnPFYlukV5zU2ni+lJ45llnenjJnZp1x7+oI5o
la8OdFR1HX10VMGIimg9daAohHX0IBf2micW2bwef8WrDhRDqbgmR+XNrONg78LADnTsNdvIt806
ENiYxKgEMBSZnc6F0Kfdcn3oNatXL696tnr54jI9bEyQ+s8CzWVmnOMgGFIEWRQwzrTKLUcfmkSd
a8OjitLCDZd2BJmIO/b4TFFZW6JHIniDvO+dSzf0JeIglHT46OMBli1ZFBrATCp1RIkjn7IuGlAp
jT0aeoOWAZ8i6xJs1VUMexqtMqOwghlm/LooghZesWhGS2EHBjksGXiGRYWM4z5GRSlauETExd3Y
+byRayxZkM8aiy4AIab02G7S3cF9QAHlPr80RxfD8O3/r55gN1sFwd9KVYHg+h3/fsz3ZvBxS7k7
VVuHVbFJSln576g6cZxDwipeXoBWrkB4sPP+26DS7rn6O8FemAUy3S6sKtnACyjeTT68yY5KJbQ7
lec9LIfo5T+W/iIAzDSLBFJAQMjtT7Pc+NWRSU53keqmtCgJQ306rETxKOel/ps67a1looRQHa0V
98QRudzJ/HDNbLCAahZQhIh2Svj0gTYQ5oInHX0I7raCocISjK/atT3Cbmj7HiduKYmvwZ/S/nJg
AwVfIj8e5XK7IImdDjUdt2hLBLt94rake+f2Tz4eRdTugK0LaoyqacR8K++JYOPT8Gz2TmzyWtJS
7x481FXAv79/JyttFYkVDvT5d/1eHw8T72CXtrVpVDf+wgDoxM79RMIvZyGM0K14vuWZ2zTSRPzG
PctV/iRPlcqAAZp8k95UVLhYwDZ117zGpj7Y5cCiINpKOVSzwKAtq1eBJPkdfJ2Wm18LJmdMoWxU
dppBkK7syq5lYsK8iCS07KDtDvJ5CyyAvit6nitVGDzMoWPsVDAJoRK4o+KfCc52KkZ2Anh2jpPm
IJeoSJ8M0MYrjDSOwx6u1E43zX5/9/gZ210SbjVOfjqfzeyRUiFa/piNX/m5od8qs4m2PO4U1NDm
eLxPgvcucB2lrDrWFg2OTjBRscLKSQQxg0Tq2QVi5PaKFOAXsdf493p+EfYor8/7KCKc/CsgxX8g
cK95B0p0BtRk26O/hxIn3NS6wXK0G2I4SAPhOUhz2995EUPIUTH3FhP5jnefJYuNfsKbX4/VD/PQ
CSy7uPEyLUIATUZmuKlYNRCXU786EXJqtrAZMkqhSHXD+PSkt/16UCjbiag46sVg0dmG/2OnyA8A
habsMARypHfWiYOEWaaSLAqe1XqWH9e9PINo9o51jmXuuWHGG3vOMzkn6kxavbRcYsEDQjDhJ5+H
R8whr2KNnA0oA1rOQ7Yc5d9QHyOEcZa4WYF90fDc8T5ISr+FnXypfuGchRzYBKLsgtqIGy9FLEA7
3/IYdLvJ78OEr0Ah4QAhSwOofB52zdsGirpnP/6wb6MAvmwYceHedq/ZhiDK4BKknTaBDDxl7R9L
uJyedDMaxCgy4Z8usyBgz3mK8Tv2ZssyrTwxCo21Yps4CTqOLmP68viNhbS2XLohyo0iuMwCM78i
ZvIsuSxgsofqwVu7k7vt7z9O0af2lEdhuAckVZzEcCmpQ8Pwp1zbLPy0sxn6TV1gkh4+5MqVUFWk
NmHiBLTWdBIQfZ23YShoHyoGx+4bJ2AAG51bleRJn/oHX62/ee1ZqpFbs5jffx8eaI1PSlXhqmmc
dDTV8HApcE3EFJmTLdufE4OiTywI3qmQwsguu2BeY4Y6X0/ZxeLpGcJ8/C1daWYnnf1PIYD0/1ZN
f/5SUYrnHtCSaXxwKxBzJS/MkGxS1/uLDW7Ph8hieiq4R45GV1MT5AL+HbRPBALhB7BQJGbqLX4c
EXOmHHp/K3N9uHhIQNsh1HbrcpenlCSrDQd/F0XGqvW1b9skM8mwgsu+cjtqNrivptfyHOd9gRkQ
V8NuOlJP8wQa64zDEKGYtKYIriR6Tt+pYUvdBlwKhi/GELfTue+XWgc3Xm+UfpyYFfyWN81CNxUI
yrYo5DhIuqKdpG0lLqSXukEzql5HCfcqOUaM3ZgqBYB2zMR39AZuCxGXFPXxqGb1sS7U/2hNYTIV
87ymuYZPnnwzWFtNSH2jSYL6jFF6+98F0HtpHk7CSZlWv/XY1+8kHyzO+IsG+xyt1g3qrpv6vUis
PMuqJjZt9kR4RoZX9yE26Tojpq7Q6JHWBVyFREG8QRS7dj8k1NQfMfn9wh957oWE7CQJsBwMC++a
NmJjpjsCWB47P7IWBjjW459+HYl1jpRzg+xWeee/ZAvmeHcolkWmBnu50HweO743LXhzq19S87Z2
QxfmAnF3ePigeajxsQnLCsmlOehv4J20VQ4LIpvVqxtGtngQuCFGl8lsu+S2Qr4RPI85r0mObJi+
1UPmNzq3oKFk7zQYBvhRlai6018jDKLRYgCZsMsgYDxO7RjUFiMnBw6ul7YO09dIjMhxYBaRTyiG
II5I4zJyJghWTTo5u9DHiERaepugT3YAlWiIZufpiQ/3J+uMiRuEj/OBjvWUUoC2E6mssBqeHeoO
WBel6gcbHTD7DzQ+rNfb0R0sGgmQYQ1Bg0m3QXLwQ22tT+eaTV4r/bq3Yj7K9mieW7tL2/+CsJPO
AzJ7H6Ju3b+hqc8Ep0hsqYwO5+EhdRjRq8I/kBJM+Vepw+EzJermaw8IGIiNVXl1egiHgGcakKrH
JE2Fb7HgHgO7uIlOlL/DE7f31JGNl3uAIiUEv4NUb/s3rzTA225WKgXAxkAnWTk44zOgwsm0d7E0
lAoMuVSxeXY2rmppRzIecPTiwXjGpcdIDQ23/p8DhyPjm/fM0AOE3Ibx9lsqhq5as2Jr3220WRW7
m/9kfGsI8AmmXij+dJ/MO87JV7hM6NciytVQfPPlVDZlLwZqd4q05afChTrSpvoh1EaQFsFtA5TC
FQQY09HksjZLwTeVWrcPuioqfDfkKdynX0ccRVTBENIRPuQ/e6Wu5mBibY8anhy6J1yD2P1pW4r9
B77hlLq5PUvKm8X5BP7CiE6J2DeNmOj66DmMtRoJm7ytXbdd0R19fKXy5ChjoMuR2puHeT/Y5gE2
Xueu9LnHYP50WzXFFhhU/h2FPjdeU9Pd+gDEFErU5HFIZRwba+UeVBfaD2W+Okae3D0i8o2bRBBT
fzuZAojrC0J9ASYcbuUkY+tzGyJJJ68PrOuYquWPCac9ey6PvjLNbPW0H2pF7YXnT1YeSlX87Jdj
iVBf9EOBXqXTropN8ifc2GiVRoUmjdHGgIDXv9KmhffPsisvRleiaBWTZmTAttFWXhNn8XBqcz2u
CnUVkXKoO5ixiqmS7WglxZ2pt0/+0AQq1M3KP+hdXaYf+IPd4LwIWVfGGPWiQ/ZA3wymOreAvImf
g6MgS3sHOIJm52CsREiyp+3WD1wWUVNoInJ3qbqedUEbty9Ih98b5kzyaapUix713uyiwQRrxFvN
45cgL9wwdrqgO5waRyrKclvy4dUM5sz8F1Ttc9e7hxnVe++lQ9B1Zsy8UtLrR7MduAPdmjcE4sSv
3LTgSIcpu5wSuDcSF9U04Q3kKn6SjaMQ2/ksozYgxZUeKzQWL/YD/22dMWwklNmuWGv1u9Zq6bQv
b/S5BMoMi7yvr5Ql897YdVHy0DJZriM6B67kAGA9YU2kCZihw3aUNwfCZ10f6TWopLy0qewSFwXt
DW6s/ieSF85XU8nryallgD/Orkn84EnDDlh00tfgYqInXZQF/ghPLytQfqnXQm/OQG9abbvJCod4
7Uu07yrxeQCFl3mErfqqs3YjNQSaa/t0zYrcnsnsUL7421E6OCmILApcmzVWrtdNBnbw2tAyxKYJ
FpccIx232EN2ycQARoY7l+sLoEgyu1s1TgeYSq6Q3IwxL6eh0XrkOmraTM14ITFMWUDDt6IB4CdP
uW0oGn+L5DGCQBEDliGKCfBwbgBy+E8ahC0yvS/x7R62rnDdQJBxpajYXJGTmrh2dCEkcb8eANH2
KA1T7jL/c3HX5cqWS9RuMHtGS0EZV2pCjDWjWsg90tbLvJ+TyxQJlN6fcSllnPjrzpNQjvBpL9MU
0ReFOEjUbq/aPzCccQ5/LiuGaWpD+yJ8GK7K919AcoZzS50PyJV0dq9O60eNWSdSpx2gYbxa5DnV
IfMtvt8alVqjK/r3IjEZClA8YKPrWDTcW1Hkal3XHAxGMzeQjnu0EY+XDkVbN/+ujQTQMejdsbaV
8QaUTmNIcUJopMTkx4UcE+pmYkORygn6JRkDSOIcsRWWsOsNLJc9bpUDwpCRIh9PQbtVE+P02YOk
eoR4+Sehs0h99KX2wmOm0npHs48lric3l1SphNmKfAXlfVgmXL8rqGcc4vZ3lBvZ0NbxxP+cepXi
4pf+NzCg5Fr15rLvT++WcHBQn0tekqISKnxIFTLCYaDBw+UUbb3PQBB05AMLHi9Bq3V0zyuXN6HZ
pjo0HDCLXqLyVsqb73sgH4njMl8dcGR8wICcyuuSuLV2sf5mTJjyPquXjyK52pxHHJiNfE+FILet
2Fg6slGsc5DRL9MJ8C6oKPuNT4eGEtz0r672ZQfUubwA6J3xQY8J3GBq0OSRrLwx+AKO7tvUMtPU
VpPzSftHaRakz4O9lnWEqlCC2Whr6eEXjzSMs+d8JjljgoLpB1uoTZGPvK/UnsFg2CQq1Ub3+joh
PZw+IZzRvSu5LXl7WMcNUEPEmyTermQG9mhlpdZuMweZYMMm+1w3NqFAkF9uM6U5y/Yvpl00hi9B
gVKZ9cN5Nm11glNUpFkBIB+6jonpUAKiQevsn0vMyi4aTI96194xeuzXr2rF0s0pIyvi0oNRNWmR
7aHlCsm4JD8X1VK+4Tg5JyFPa5votMGkjqyMEeSSGtUFnqYn2sz6fRkzZYPQbGyuUzHbaDvOqrWo
jpfN4iwXg84WcRU9bFzggr2QH8e/Pgg4iN/DGT9YXWgV9iWsNDS2kF6OUl5cuMczbrIo7+4WDrvk
T6uswFbX3nXnDjpPOdmO9DTiAZF+Fih8KWhWFVmtZcNXNx5TAfBZYxtpfdg+9Ii/vN2mWMoyA/XX
ohoNT0awuzWtGK2j/doVY37zB3r31VniAE1YIMPLHxuhauLu0lGR635sBZyyBjRQWnQR74NC4GYM
PvIcXo8nyZvaR3efu20Fa+dbTec2E0DB8SsAxOtUaFEgQP5cMExOXn6+iPCkR/VBN6xM+utRn23Y
9RRdnr3++MwDup3EIfKaljEbBXzF56AAgD5kKBdttDoA4HPHcy5Jreu0HLK9n3WShuJ6/SXlKUFQ
SP2VfzdPOYAaLWDjlhrIW7zEX2Co9/1lE2beb+fGbJhqwnBOzKPBUYI4rbEUGaWL/+Fqn0GLocLo
MD4rEuCcd2VR008CsgsNJ+jaKquJGqAiCT9hFWD1CTEyijF16j3NnvxneI4ElZn6tdvdJ08s5BS1
hcCoS9scqYxVxSVzLliw76cKB+i0P8zFCd1zSMPjAbR0GVfOXoVKI+Kv0XBAm9rneeUstmdYcHMa
MEaKI49KRZ9XW1Q5EvT/uCJ7G185logFrJTjuU0K9ciztHF80X9kNfKQCT+6+5sG0pCKjIN8xyas
/uztBYLTfAWquKF908QNjxONbhLJidQx4mklY95TNhRudERvAs+NHhx7Hnt1BPx4u6dYqXxlfIFU
uY5PY8YTeMpF9H/mUIo4HnUvyL/ZzDxeldq09efvgI/LaI5OUSrBEuvlTm1cZ32w0hC3WmGS9qyu
ax1KUl7oeo/wjzKz8+Ij21C6lPDtWEOcfDlgrgTSrZRFE8sedaZc4o4gtkMGXLQpgZigiwaf6DfH
eFk7fZZuzZEEedj9WE2yH6kD/U3rKpEbD8ZvRWCJb3XlQDoi+C2LltYoLV5vWCGcHZwM7Tnj5dIU
u8CIGeh3D+iuBfWYqVfOiW8zjspiBo8srRl9drEMgnsXfk7l0H49gRyxYuuG8A2ij133sn26Rcv6
OnrcNmrItQcOIJfVgDuRc1olZ2bVFxKPt+G6VSwv2R0dygwA1dHROxsCTP7EL0VBYVwVC+mt7r4e
/ngJpuFr8rkGksWAJ74gbq6uGPqJhbDAQC1/FCy2jGdDKFcawz/9nEwAqsEfX3xy7HLpflxyvdzY
wHTFjG3rRdZpXib4Kln4ljC7aZcGH8cIyGV2tUTcukP6v249yMwKO504aMn7QBI8kgvZumHtQYHF
JP9tjc0T243JsDzAnyYntHuGrJqFl8IOeFnUU4T3QYFU0VGqJ2pFV6xDhzm23HdNk/04Zoj3LhP1
IwgEr9BBy05KbpBltRW0rd+BzQmWWAYxxnseDa4rSqgHE+WcYG8k5jhNrlaeM1Dj+yCNKUXAzmQ4
/TN28qi+/rJk77opDGKHGbSBYWgFJogDTNh9PFHfWaJt6VwIKYWRwKrwN/Y9eqyD4v9FHZdvzw6Y
m0xZm1gdBcL1MMyEcQrxe2+PlRBaRH5uVnyRL8Mppxet2m1q4/RYx0TS0m5n1Q7n/Q9qrJp1V46R
whOZEPX/Hpww90p6h1RROyflsIdWrrQssEKRaDhMKvh7jfIHShR3hiLDid2QbnHqQUGeaib70ma3
+i5uIcEmcF/TZbJQEFSkY13COyuhG8wHEw4nOxdacR8m+BmoE79TR3Q4fYQSzOoZ3OP3u0TcTCNX
m4gZS3LQVCx5hzq2Vk26BwlnzTjWE9o1Ls1dvHc7EbktnKRr+3WoiTXtJ/nQUIZwMw9nfFoGx1By
qTlmtg9aNfKdYe/NV+hTXOPf4w2nhOxA/LGjnjCYYNuJWOq0hNpQF2TL1kUyluxvcnkTHrECJlXq
QZyo8Fx//VEKPq671On30630WWdT8LPvLLBIHKrI0uPUS6/ECyqQ1HF20Kogs4QKnmr+F1xox/LB
U6XngNA20ldkdeXmW4myAdXw4NuNclF8Qc8XdTvLV5R03fMlC+/JMe04QbrQaXQ/tiPJWIFjU9Zm
6G8oc1Z4XQYdSgEw7BLknaFtQicQliKA8IYrWRbdNaZRlytedl7Krwh0lM/eVgCFRcs80z7E6d6Z
Ctt0vSc16wfg3vlLedhC0IUyCBbnDNbNIqfRkXjhoqOzP1T8uX8nA5HqOJjfHbqL5FLPSjtrsS3N
TF7tW4pmtp88xmCUjPyQaEaT/G6LDVPeCYKImlv2MGUZxiZJnu0PldbCQa+Lbt/v3mj/to36Pn3N
oet3MeAG6djMBm9MQSAhIS40BCkaw9A1grheSdWBkmsZYkx+2wrLL7KlAeHC+A5QKhlyrgBajlFp
Q5aDgpyCzNFBHzh0tjIpuTDmVOw8kYTLguNxLWMOluwcS1+P7LVxM3jckF/2bUWxMaZPeQhjNSoe
2wN+RqkngDlQDpe7NWkVR/90vph0PtecR/wX3BOn89D+leUkf1lSX7EoCnEimoeK0HUUBaumDnoM
QodoM+EA9ajhhbbMF4OVhUAMHZTGe/XB5oWAUg2k0RzoA5+6SeG7T0whPavPv47Lyl2TiHJ2XwFG
LM7enACxiC2Y5/ABmhit3gvY4iL5dtPfXXHNrYPDA9N+qLiT6fuRemUQtF6A0qwfHTM1RX2OyRwr
zlJGR7vp4+joxKSX08lANXJ0GU+4gR/j5Q7w6BVmQeDe6y2RkOwdpXfU+rV7o/uwAjAKt1E0lIRa
L3EEvIjWZIiTPp7Jy+32/5468zmlK7kZbRBK0oj54Egma4E7YiNB/SoSzJrnZCjKgXpd+B/F2RGJ
/ZokrJPv7AZhLLxWbPjcKJ3kwoEsXYl3x2jiQK7drIixQAQDYYdfQ6Qkm5paZ1qo69jXzEWR4OvS
Ev2Ng3QwjmtvliXPIiXxDL28LmlTctbJFCN5eOkwR8XX0NvfR4fTQF0b9UyYkX7E3isKPgVz3Tbo
MrXV4MZz7Y1IzE6UrcZmtuooWtZyeD0mPnYKTvy+WK4cPkCTrocYK2uYpzLWTQtZHHpinuts6S4z
TDg19oCuBnjk/8IQOPc0rI0PPjgakliP++WB2HN8SAqt8ocXrsTSAHb9VBfLPiXN7nwFcvRNMlYd
RYO3/q6n3oA6tdhPMX2oAV+g0rgwH3YG8+trEZcxRAVaQHvgm9l/xC4r+Yp/bkTej4r6+5qcyuzx
a+rg8h4NgAteYW4xK7DiOT2Xw/cGZDYf/aRa29EBUMCeH0o0Y0Jecr+6VR419KayiHJ9F+UJw+bG
x8bjVMKocnr9GUiK4XY+JjFJ4YfnvORz5XfThEnqLqsiRrJxbQklrCdArj8Nmq6xq+9udhL35CRe
xA1WGQCPljGa2VzKEcEqqS68nBjylxdrQ7D0JtYV+QURjXlh0dChgiJ6CRKt1QFMsW5F1qs8YZaI
M1lwo4tEA/yy3sBqFYjM7J6fnysPlCytqiXccRJ7RYrjoHW7Gan6CuQyRny+5z7+xTzc/GUk7B92
yXwxKau4kT9E482kP9fognorwOEOFd9+D5fYQNR2NE72p18ahCWB9NXBsXnZ01LFUu0662XjBU0i
Ol56zO12rnRvEnQJ2ADdJvBA/YP2ChwX2bayb2SvLporXx+1BIyf/HvO9ejOX5Fx7eyvRbnmvfzw
+PUJHUb9hs5GGLj5Fkm5xtYrBFuqc3ECprT6JX4ADMcfaK36DDfFuOltUbBxUUwW/DvIzn48bViY
fLjYDOTHWp+N1nGVqhw1xl7M5HyRb/JaiIO1UI1UiI/vd42Vorgs8oltZjhXQJTSYXmd3zpIUFm1
s59/IM6ERQcw86Bha3b/NFKE4LzItigyn/aEN5WxTiBDVZuzKGEeZmo4QSkVlkDbXUP+60+62sle
Si19xXPA7DMEvChVWHsVZi4KMCzfaun6D4NcvAfFmCsHxhq+EAmlIXTtYTtBfHQq9Uuo2YsatwO0
0mWVuoiakDJg+G3HoMtRytPaJSQckltMZWwhQo7ROTJCMr2xa8i/neRtZGSPDLaovN7tAJ89vSSH
j5BAQxlHX26lRFWmpYizxkUXCegTU8RXaQuXblw8mPZM1Zw1iI7jH7Q/dcrLzabmhpY1kaEMfC00
oJheXzQumqrYiabc/c4vVSHJMycZlrFy3gY5Da2ZYXARUVDPzfV0MyHf4tsRBJrzYS7YNqgkDY8B
X2JKDLCr0k6R8+5NQjvQf8ama0JWx8MmRbsBiYLaacUTlZZGbEs6eTKNFrrkEWf/9I6Ivoad4owh
jFK2qjpkVeH8OFGnHwMOWjdPti2MOs+p+FVwDqoixbBB7CgSHasqfJM8Non+i+iAF/EW8mzHXqZC
cgMdBkG1birKdC0bxQT7I2/F7mtmnVhHCFXa84JcJt0GgI+COLTo1W4rruMIFgf/hW8GCwZZPCoZ
bpVEfD0PdY3jp4yL8mc/dg75rKzofzwJmVA9qweYoQmx2xw1MGKNibiNZHrTxJ7TRBr2Z45IlRPy
pjXZ7hc8CpxaQaBUEUUduuFCDMHeFF2U+br68eZuXWIan3+39EK+NeOTbwVyT9mSulYA+THqki6A
V0C8Aui612srJymg2Emhjd4td1JUw/vJGy4YQAukqkM3yr3qSVOMMujqLmHlVEYAbEbnaTEiZEJd
ql4eaLdL7fuHx7H0w9NsCIXKX7MbGLDPEMPhTXKLZ7Ez85QiI49OqpcTlI7Mr7tS0kTKULtHlqX+
yND2eFvdz/a7YlS/KSwuvQ1RpgQLzVUrj6F11CEcQCznUF5l6TCO/mUrjSP+ru2W7VK7LaqgkAaH
b1XiN8A5rGeX05Sp6mZCu2J7D4sxgvwKDpMTkH+/DE979+hl/0CXg6pQk7W3ryZtoSbBYIH444wY
IJUO1Bp+yDDq4p6zkbjhV7QcFXX+B0FXQj/KNkcT2gxKD3z3EefLmUUGHoZKh95kaV84rM7yeelu
tO1sMw3yMQgcWAcvWfnANec+t53UB+4xYeY0AdQMFLIjCuztpOuBsX8s7PLSukfdkB4EH0oUX85H
7HqkvTEqtHMwkGngLXgSejI4iV4BXNfg54jsIOOg6faH5iUbLawKqgoVgCXA5zdzobJnsFLCavVq
0lEEY645NgBri+GTfogjlMoVLEXnrVGxt7X4wifDDX/ghp3D4Ym04nxBEl7RdwYl1bJ+GapJ+Kl/
xVr1bVJgGcB4VXNal/feONsd05Ik6FJ/S9/tfsiCe6D4WAWlKXv68tjes1cbOmk61F2NwyQ7k1Zi
WIrYYK2KO8gl813jRNU8+wUinxlt54KP/CMaNoJqMVm5/JYr0YLdexe002ZwfSUOFAaCE0qNtS0x
DMY8neSPq26bgKL639SMN4WIEYesVtxYiW1SZSw80GrDu5RBiIrUnbxHzYJqWJR5GMja4WqrdouI
FQCOraC/s7ssi9PgplnpdhOgjv1nHnzPmzambEsHUYG1IIdeh+TggNCT07iodleXx63xvA8xZ/ki
4mdlogQCRZHMNxz8mbGjwiln++ByZbaCj+KLXlIVDcj4ps0u6iR+hZOzBBCERhwBOSEr1By4yQec
llb7vfXu/ksP3pZCcXapKkRp4fQC0ZOQneAuO66f/0F769qxnKjK2gDU5iIHiYQAdqkN41uJkDtp
hAvCOCKuMlFDzoDnXq+6XVggKT9FLsTSea6PPyeg1JPsv2Z/eIHwWoN7pvStWKtT8wuqScgpBTN3
Jo3i4HoiUHp/9XKUlYaAG3Iy+FuZt9Ik8x31ufocC2p0dPrwX/216dKdwGhNxEvSOFL9HzdPWogb
HozFeAFecs8cyEy/btCRUR3bUJOipvRxcdR171gtFJr4J/GSrvWaCEi6/eMWNaIs4QQb4x7mrGUc
cQrHOdf/ByliNZfkWVRAwojuzzk2gm0mpoMVe/2S4rX8satQuMCQtuBBU+XRISkWKZVpNJKZlm8a
5xkneYCQZhmalAzu4r4hrF4fgQqB6kSLw8HczdkzO1OcbNJ8FWHAxtOoIIRd4gUHjEZp23Qzvc/n
mxag5oiqHNO4bmiRz1Gmn7cIq8e1/C16yfgt2zvvM9lFvrfRf2FppsxHS2PCQiH3PiJ3EEvfByOj
sQmrddVUCn9X8w200uWLKFQm2N6XwxsFmSh/gFA6VEw9KGbCboOqbG+mFNhjZgdt/0RlV3xTH6DM
rAyBdDz+laadqw50K+mxylcRBwgVpOv1wMlTLZ8IkRV52WCoKtpLfvyH0eyV50W9ezJspkdcxHSB
ZpRvEip/OHzIhlsVtVuZyzs7+w2Sx9JFmcIQgXy2arfqqoQ+fBQH1pRsA6BD2SMmy4O8T8RIIcbO
y3Y9B3Jkm8acLul/DhH22LOvwPoDkqjnGAZYZIq69MrGFJw+Y3EIY43XpzmkAttUA255calKC2lG
pnRhUMpLkT5n4JTkkazuWvOsDDCj8rQ7VSiZ9bufIPhg0o8Jw3NAkHUfAPfcgJI8IBxrx3Fdkk+k
g6cW8+ftwkUfO3KMZvUfUN+M1+LDFM/r1R23vGTB1OxDWvi+BecJ4FSKjGinHgJvo/BrUaP/YptL
hB76ebrAPpP/fLLijwlTGWyfB+KPlW8Vv6L4+qs57r/3JgzY2Rk0HFIBTmsMewL2Dm2bQyRBYIs+
y+SBfGlLUAwTm3mmzyGA9k6RdynOnMFm2VRKMaNb6q9/G0S9tnobEct2z7rtbmOyFOet/JBw/J47
ARnfWxhSOZqBKo5ZSteXDlkJCodu3HvAQMekTPJ3StlgXfZdDmQdotSdE/Yry8R890+vn9xx4Xxq
ib6/g2fCjQua0k0SaiumjbEc1mR3JH3LsukBGTE7/u/CGq1V0qNByHNYCximozF6GewA4DykScQa
pxoARdWXHLJZaq1DcjIUCsVgM0cGVSaKwo0H4RSL0bzXjjsJ09reME1DpJZmFXi2+Tk0K+c8r/5E
rccbCe1mvyl6p7pVdtKewC2iDEET4v4ohXfIxxvdUJDZ1fmaLNE+flhYRQBW6fKKrCI6WFigJ7n9
eY1T/LmHWXbFXq5WY4ehpR9hBIFDtjiufxf/+zRP/nByf2d8tYnZEDi6mfpbk7yGA4SS72A2cgEf
hIJ92QA3IL8kjcQf+OqTQ0TfGDJlb8GgRKYSDDgG1IBnc6Hf7NBBBdkkZBH6af+T0fEsqTotZV87
klvOaXFjIVuf3u/DkXaSLBQWqG2byClOgQQK8lfecTdlO4N4AYunteK3GowrVRc5088QVtkAEQpH
OqDHTbmcF2vOGIsOQqymqE5v4Nc6yOOJdL/OPpt9h3Jgz9RpwZnw1uejoiqzxDmy9q3mPvmMKtph
V1uDF0TXWsOGHFylRjMEDvk/DidAKBx1aD3ZAswPMJbNBAu+bpDqh1Ha+gFDeusTxKigQo2hs/KQ
tsGOtnbdPW0geczeH5PFpYKKplo4o4wdV6RlPjDwe2ImKHjjCT8tMM9mZd6zdlExc0cjPeIKBUCM
H45HlZULADVs+tFa3VJ2z+2Uk8Ez6oJ3yOcw3QjfsDfTGJ8Y9nfPJBSEjBiLwmeGwl5UTeG0/055
8F+74G6hDfYTQkU9XA+TLNzHZDwTku+NZiL0f3DBpR+yfQJ0gUUCAx3PdKYrz1tVOu93/WzbYRJk
2Sl70nT9YnKhSYGlxoBjT/nmp3yrBpB2vcCEUumoWCiCIMUXFFjHYeKK+hLy1qmAsuHCAfZXibiZ
fEX6gafocgCWIiHjfuF5CoHFZ29ky96/CHXa4bU9K0EDudTUTNgnIMJy+OWjxR3+Axe1i3UIVyNC
FrpJt8SaNHD0UqZzzqDQQDoC8esFYxOwve0H83FuVP35uaTcVPKFtUktMuEwpANAvVhfvUqCOa3s
Xp6fWyE35m+6NHxP5q6TNh6X92dHbTcP7WhVYFiFJPUrPTaBWDGOFzXnw5qfC9kNSS0ZiFxW+aQT
i95YtwzfqSP7J9RDIQVjykIzPBpv+vFjBdGriiu0SjK5rHRD/A6p48CpnfstyAw0UyUeA7iiCeQf
8mhUikjbDhGjKUl/4XygEGy2jjiEuFgUmT6YOPWQ5gzKIMYZ+OiwyVnEOzetbwYRLJJLV7cDPdOm
GKgHz3giMuvL7ErlMKQNYN42PW8sgWnp+SibcMO/KQlOL6NE1eOtH9+JmeMk3vaBjMG4PzFR6kEx
BMzhpH+7V7krRq0ajOd/S4DqG7d7Io4GLPZPo5QpjanZO499hEtNuwv5A/K1nvt2DCpq51O0niEa
J9qAlPBsD3YuJellx+Jlust7wYcuAQq0lQBOGy/GB6xrK6qw2wqjYIHEYLEggsZDgobSiVBWHR7E
fCzt9TBJQDAVlrkAGiiB4xzJnMP7xmK4O2FOPccsU6Ag8Gfy5nXCw13qP7LBhPIZLIH88vo9henc
hB3hPGuDbA5o0NC6SUnufOo44R/OdIKvcSQV88arWRFKGhbeBWC20+3zB8NaCq5ZJTdJuCfQr+il
mqpiHSUq2Zq4BXxy1yVJyOxRBEngXi78dDEYcja0CO7xCpgAfNoq1rj6TedBSTGJzk3z9DdPQcob
O1lmKd4/Rp6xTRTxX2nyv4tKXvXWlMzC5DI2QilEeSR0rv51U/vM0Wh290ybh5SiSCSxz6ZcbOlb
6V4t+RB/nD+4ce1jB1nH1B5rkuN24VXM6hS1uJITbGh78JJXwhbkdyIH4MqxBVCSyaI5/qch2PnI
WtcIlwTCyXY1YBK8OHmkCPGod/nWPgUaC4WgdfvbBmR71nRPOgO+IYgkzGfPDvZ89AV1WURfmuY6
vAiMLXM8SQ/hk3DHDrzDV3RkBlYNtKy4o4vZBCdCTbH2CH/5rFy+5vpVwHgtaTzfaCiretNW96x+
x7K5sf3KA6YtWyhs2UUEqvxXDZx4qgolM7FsoEPe40fO2RntU2zKbKcJU91ZAkHpLhvxg9kXGRjf
ScmWmFarFofTD08gTlPc9OQgDD+F6Ll5QlgBvCHWIe4SUsEZD1NWq9kraZOulUTQ1mjBH5iisiN4
/UhEolxHi0JLZyWgVMvsmPv+3MKuJJWJSkDHrbijKQVSqK8AiSO3jkEt7v3xxcwWrnJ8ebesU4vF
+CkqYjNRGpQxR1K+xozCTB0PDrqJUiAzoUOxYGPUHZOLaG5KsTxRKNsDMllvQc61fzy5J2KYYUKd
q0viB6gZLoZ4+uM11eJQf6/FSGUvOFk06TfOuoKnYnpetCSwiCei0wc0tZTiF1eQZ/85Zcw6DdV2
x6mN1/CHrNw5dmrxUxMzGFfKITYNSsrm+vjsXIZOU10ttGQOBxujKSyY2zfnk0qMGqiP2MQ+ud5v
PjMu0yD99nRBUXvTl+BAD3bOYwfW4RrhUsfH+A5d0QPDCM0JI+hvYuctgE9lOYiF0HSDpLl/Ge22
S0WZH1AuOJVZVAQ2xRpW4Me6GZXBBVrggsYpTDMXOb0TrXoKv+HYImIfIncYq38Ehve7ek4vdO7z
/k1iNwa93p3Tb/KsfigZsjCXwDZU3W4G4tP5D/lHMKlHhPkoWJswyGycMqwcAeiDQPndkp8VmZTj
pIh2bEJ7DbilCYihowLK65U4XTC4g47YTVCfnSi3ahe2NyXIxPZBJHf7v264YEDzGOUxMf9MJ5Ni
FWg/i2nYGN6Xu8tqL9IP+OgL0kOLDTjQohP3UrSNaxAlqvwX1C9CbOoRIE7myyHlY9On29ELyMBm
dt2AA5IvkVjfHdraXoGJbCW9zwd9WpfIQn7QCtemsWU2aMksArt1mnIcXfFnPnsGheAjM0kfI+uG
4sYUQKMQqyeWpNn0jU/loowC1R5uMRZ+lJZsu8spGOC2DwRewWjVweDpOmO86FkBOK0ZZPP8rFGU
FMbe7P/3VJ3/CP0s13dKrrPjqZHWEIcdIZ+9XLBQGL3PvvEJqsM7aww++fCFgiCzLcP20TJe4qqE
7XdD0Dy6J7d7MXuDjSPx0wau1ZID2Z91Tvq+XdiKtQTuNlpOUV4yTE7rv/ttF+DovDrv79f9Enyl
UlFTdyzvQxVfjYz27f1o7TUOozp1NHpdemJ1YlqI6lOibkPE8cXOO1HoSNGX3w0RIF0NilPKuFnR
J3UsbFoovxN2f9pWHY0/9PJZIrZ1+mpreiaK8b1bRvyEEpqQsfu5KOn/SpyJOFBj2bfcJBqLOTBH
1fHUM2JVJbkyLWyDWYApwxKtV0JMUpgFBPDoflaTnInOpNn4gUAV0PdYm0PPe8OLYug9tL8dEtcn
KKr33IQPm6bLm/GFESxVICjiZbMWYP9YWFYVMdd8/9wUlX744rKx2oEzhSDeOex5DHua9SDz1fjv
KVxXqEjt7w5PXlNfjAvHuldZSQqQF0QshQ2fPMvRNQlpulFNRKEzaL7HbUG7tC8XJgNsrhyQk1tQ
kNI3GNFCShT5S91UmvdOL6yaGVXZ9HEQo8sfv4uTPAUmY5lkNgnuUyuPJ6nFUOYUKruX3jIXS3bQ
rrBtLDKmk8wKzbxKleWm8dUxImg8sUFaBAhHzcNvXzCkSgYp83AHWs3LpuarFv1/7sKPGPwwjxB3
vGRAnn6POZQi+6gcmNxsfLiQ/B8Ma8psO/jb30URH04KmNiIWD4qcaQ7uw6eI3/tuv7ogLLlin/q
u0NTyhCq3WAvRtSzOlKai2JC6qBaiYncI0uy4rwTB7G0XF9JKz1QESHQUYF0XzTrrIRkdhyOWsHo
/txof/ufaezCAwoAwZeVHeklIuXsc4YpwpxFmqjjoqZizPOCX+DYZJPIewRsOo1nGZENuh61j37l
mAAbBDHmSU8JlY5frhTVyKumw9jJ9jej6+l2PTkvTsooDjH+mJ0jSfe8LL8zJAJb6+Q9DzMT5wRj
YxvBYHWsgFehg2A2K+E2yF7vPW489dTSpBD01tZwq+Rl2Ypl2Gdk051xd8MFMHDXK1ls7FkpF+8A
kC+HhVKB5vGxOyidxTIWx2n7p4X1rdJ9co1PmIog7dPJmDvGttfFY85JoVhblMIajnmgRXlsOOdY
4Fe+Rr2EAWIPr6rkodAv4fZUlZLnTPPQ+Zk1TwNQye5hn8UoGAehMEEt3s7ztvpbXt6xzNLQqpTr
fyzXWMfCxP2gAPx2v0mtXx8PuzVaZdRtb8AJMU8xwTw2pWlg962HFEkdvTTsN4CE6C+3fiTIw3Zk
9GsAnDrCPSlRPM9nBsvRyg5gh8jq3BPA1Jo9k03Y2bAd11L6g2WDhEkejLAkVuxgzpdmP/yFDHGs
W5NS+VGUILRzUZ2tOntc6UJ31tNvriFx7wsTNmEf5D6iGie7Zqhiw7YdqrMXmNwx8qPyZBBzXRDO
lsLGJv8KJLV8LErot3ODzjZZRwyUEzkirg7O0DYzaFnQEYBu3vnbAUDSK1YXH+0Bg7Zz1+RQo/TX
Xw4aUCKab5UjPZO1pi18ddugb1pdYtNLzEJnXqOU5cjyEYXmpN+2ffE5GO1dbM5BGgX9yzvHg+PY
zDlL5gYvRwxr2g/7duf+ivl9lEt/krJ/0xkcNey6BaBFuYlZ91udgwKwivesuwiwq3HKAkIwiOAb
uMvOBoIvJW61cg2zcxgvp0GiTT4NB7JYzpXlYUSArSN6pbEpgJnVp95t7XakpmRScB2bt9qO0oj2
CcP10nFeTdfPIHf2VumejYysLEC5RzC5LRmWOIGucHGPMXlMiAOWXkXY9wQE1o/MXAax0pPjPuit
HB/gptaQ+xU/rtAnX9BpNWnd/cRhCIcE0K0s4EafBGXe/jeP12k8E68OyQQ+5J00kgOs/xtcIr20
XCUdT6wa3TaXwjHP19bzheezXrxSACODLMdO/6UlQOl5vLSR3HQ0sc0Q44DgqWozPmEQu7RAF/Vz
hAif4FifV1ep2hFGe+qBCRUJ+TDSWl6q72BOXojirViJ3EqKfhaI46ai2qjVv4JLYHjoLyKXtsQm
2PSPqcIGtlcBMyleFj9ZP8cr0woBESANB0JgxNoKXU+hgU1bVbaSpBMg2na+eDHvdz2CMefdcdMD
8vya1sndBT6Lzhzv9ez62k6ETJgQCfjeoMzWCJ7VScGSIjwaUXn9qyksQtpmjlsLICWtF0pjohId
YSFFVmSnjqXMUcjQZDuvmOU3H3o+DKDmSZAK0lsxxOlDmLaQ7kNOW/UXr4ePJywLIMo9UfqiVcvV
doZ2aEuOjo7Ya/G4gw8Zc6zFqxSmkkzyR5YfeLvVccz47fYMwXHywi4hvJxxywpuA3UuxpzmZOER
/+1i38+Owm9rPqUg5axahrcMBTMdbUvZZX9tqL5gYxiubuu3xeT565hUlHcJR8B4BVe/payjXS6Z
U0hp5JMd/0dW4VptChsK5091twBznTlf1FJS2ilKQb0tVrGlJW276reJHDaBAw6NfZsaqKz77txq
zncZ2wf94mRA3fcHlytS/30PkY/pm2NpMrg8RZcd7NLze2gDYUfxsI10qspsTVE30Cu2zT0Kn9yl
GMUseoqYag1hhjwaXGUwXtm6SC3JSmrqiYSp9kkiEW063rp9bXp/97lRM6yrTXrCu2r+f4vUvGFj
ibtaWihl3V7y+N7Y5Gc8fDGLBmkLZDGY8bvlBRD8XRFGB13H5kxzgFynsMt7F8rKcofhsaprwfsr
Vi5zqxPZZ5CuPXd5fmIdhi2LWKfFR7TakbXX8qIptMgTMzG4kSm7zdwzDyPH2iF532/oAZKinH9p
DMmYUGV0Txtk7cMbtqhguKTLAXCqo+Lgo4jRVFXVhhanFyYxTcA9y84w7O4xAqZ8LA5u/yw/Bo83
Ac2bWfhO58W9cjdopXeYEi1VgDXRDWd5D0iDb1OuPcYEgxeSMQrfJ2dkEujvHVlh0zk9gwcC6bFj
W84JjBjOaEmlk5wYMF7eUv52nDxkR2xHEZXyDKJTEFR0jIbSc6ZFtSGEjgpWJVvVKThoADK3wez0
fOSjoWnH3wRX8PmGEEiVz7siqfPv3OwXtBt5PYaLiSV6IpmNAFk7XVen6xngTY1s2su4qSHh3RNZ
64VoW8uFO1FeVvn6IF7uDTZr/mY1anQ10rR8jpBs9nmkPqe6OX+QWsS+5h37vRbkM/E2bcFuRgEG
S1mYdOfm5neRipjsCMhgCYdAtsC077M+IaG0cz4CmJ99eIuOyO2qJP+d40clA5/ybVKlg/19Klf4
ucYzWi/b9AUklhxqEMAnPq6iMStu8+cVVADJjWUXQZa18aORuf9sPg0V4sBVr0eE52Q+/jiQ+3E/
i9XxNTTUUaxMxhZpKeFT1RbmoGok/H8p9IsX2663FAMUbX69B1KK5BBusGspxs8AUkCoacH6DEXQ
3fGcOem+7/mPkP/O1Z+/vE+7UVsGX37Il7gXL905kqZ/040yzihrNoCH2zLTjGSc//DEIzXRB+u+
1EHb0fQjRPogtHvVLj9AZQRWj79VsKtH2iZLGg/PbdyG0Lb4kvuiPTt4hszckSyjZSP469An12PU
bWHZ0v9j2CuA735IHrZudlBo6KyF9KiQbhyiAkrtXdNNMulxGbkxtXZTn2S9uZjcrtVv+1WXoeTs
D8CGBKtZKY2M1tsro4sPBnSMgYFto3bjmJ3ZINT3i5uajdKUfpuIIypvXqTLBgnv5z4IQ76aqzTH
i/+Kl3jQVln14BWMJ+ka9Oep0H3r4JJsqKqx28BvkqSwMKO9vPhW7bWXwVE8oXMFATzZ+mfBnq/v
3w6UwyTXyznrTiyoscScx3QxoqdwqPcZa1gJNqHh5JglPE2OB7oslwcBHIp/TZMyUQJKyVASFbV1
xvT/GEcsa5dfXx0L6Bpaz2MvzpbVyH4dgbjM4BqQ5+MmnXoYZVy64qGpAXR4pb32T9ogupcenxNR
/JngqU+INr1NAC4nr1AC+KTJK2htYLUW2emcAMMXeuqMYadEqVb6wrLCe0dezQPTLv+lMVLR1PaL
5y7vk/E1NdFOryQf8ZtJYZKd/UpkpMe5qdCht15JYNQhaDX2MTGmOTpIimGLnAUdf0Dk2dKBbd7L
EiSo7CW3QS37xgCcFzEy8yJn6ivRG9pF2F71gNjpp6zwqZOFc6MOKspkOPmIQyfU9yqKduFZuxYa
qfE1mW5CC/gZK99QFCwc/kfmlorA+OaKzXB/NSoy7Y97bb7j82QjCtbah7iILyndw8aq/MI+3w7j
4FDcp/evoFy2lLCGMv5cOt6FZ5xMpAscM7aQ70IcNNBO9JpG3HmJTPYw8/eggN0dB5WTyuamqL2Y
9FtU2C3KUwuj//8HGDRv6s9JbUgh6jODkzJCUP/a7Dc3g8wvxP3WNRfJ2qwgsI3O7QCsLP9MvA9r
WI6rfWd2Mdfzr6+MZZw6wnk2klWcD95sk7dWoKqeInNKPinMixwBjeNImqVRekSZcr7FBXx3gEls
VGAH9clItEZ9NXh7TvhymheZy9Gc5n3vSA+euObwpZZo7PPzZ6TPhucrFRTTAD8NgZlWz98c8MX9
Nqx3iMRTq99l54qIn8DCz1ipxdKZPa8wXgfntFFYNhJ3ykrbJ6FtrOJ8TJtROgfLNkQRKlhYs4ft
z4V9eUd5jHHXXKwg+gWvOKXa79fJNY5NbzwPfaoQ3tmORGkdeZLDDHeNARSXwoZjj+kW3w5RiD0r
nyI1HeQrS+X/e/Ttu/72CP7DjjVBGFtnhErrMyHjO26+F/PQHZMS9HZbmtrbIb9XrlvxrmpMLMBF
qJT8HhGsVEFuAQsc9vxa+hfxW+u6A1Hb2l1bHK+oAVoMY8Y/YVO1flvBVjzrH8Jedeq4FIeyEDdN
JMwwWa95AStifJJbzdoTG+wRI0g8Lj4hauVC9mMabu5sOpHFK+c3xAbmoyNYNxN/8dFhVGhUH/9l
oWT5lMqBX4Ej8Kx2VbnijEa/WBobObiaFdj8rNTedcSAWFryPQztBjgxSPPSk7fMTv18RBKukC3X
QVBKcVdVDeidP5OniSBxqvgGZWt//X/FwbOSljvNX6oJa1+/KN6TJF75spmVpPbR4lZ79FCM9n1L
x28TvE1hIb8NAvQzSh7zJqxxNCHOcy4S6bunQvZtyijjXLxGEdNnV6dvMwL6T1tnjuEvfAZPDU77
qlAFLF0p1Xb2EFkEjubq8kumFCB7to6YhTBdqA+hx3kom91Myy0JxtKkzCOfZSaEUZKjbYC7yD99
5EVkTPdc75nR8nHSVYYlxs29efeO1kFFVaFhxql+gpNLESBtfjhJnh6IH+y89aY69AdRmjX1xnlC
HhfIBks7ozBHBAfSHuOWXAE0uPEiW+ZJC+gkK3V3Tr8S3scaiBXsLbChwbJyAGEe7z6UrpBRev6S
QGoZdpjosC5qKTyU+ruI+gbyjIzULa+2MAJ4Ox85uATuMAHYnQxh/ipwH0ph/DPvnmmnZdKBHNdL
WB3TgUbEFek0QK+AvIzsR0zGjYZCCPdT0r4J6nGaO1afbAyZ7+ZbJUjfB8uTHItQrYroXKgvyjsp
R+4szS1BI/PGFa1cc1/Ul3EBwLcaK804PJlYfRhaGGPCesL+SJflWWDUsFeZHcyschIixFfsO6C8
uBCBh7ADDf2YBuEM5j0ZTddRqNWI23V9CHpO7hPBQak89tWoPtmmhKEBEjvxO/7l9SzVVdw4QKyv
9PdJ6lyNmjt+WMVtWJrvfunY3xqVqe4ogz3Bpc/gpFSiNHibm/hy8daK1oqgtu4ARCS9W/BVVXIZ
ZYTc9a8gjlDD4b2dD8r996XwE4biw3aOSuz5LBh+oNgEIwjF9shG1RziWS3TC3IMXu97vxg0GSX0
abFhDDUURK3xEQmmc+H5zdGa1HC7bjFRQQm2Gbhm5Ds4k9+Gxt4A4Aw/Bww0yVVFmg6lCAEX6SSv
7hzAD5YLZJskUdKsFyNudMPPVlWTC28OD62ojyYngyval7qOvgwPA1g6y0/jY+96FCYrHOaDjM7z
ecLMqXvSQO9ACvCLuoQcp8AvW34U/3dXkJa7mWfrhcBhQ/v0f4Vl7YjVLzMe9kIc4xRE5N+6peVG
eQg0tzYKXU4IRvUlNmnERWZWS1DTqGnOrcYcXvqnSj+BUtziThmksJQtl1GaJoF5gn/LH+l7hL5F
1MazWEMFVzTclT+CE7mn8WxhnXjtAmpa7wk1Rh3UtbEagKXWoCwMFvreVW9xjd9Bh1UucKMk0gpf
DABPKAJ7aM7cHxkYUMG58ysquwn1XMn4BnExmu4Z4dFiAvCQq2Ro/jKrCKFcAq/0UvVHdP0AfcL7
D9VFH4oh5s/PWkAk1ZPtXXyMZAvmFQF3V4jJmFsYhyTyn5uTslOSgXTKwu9j0gvieMJigF7YgosU
a2YzTawPfMT8cCc8HhRJBJSypPCJWpjVMNFi0BR/n2Gz7rfcz02+/J4tLXU+a8n2d34ubl3dsTUl
dFzBCuwC3S3/M2Jqqprpd4T0PqgnkRoUnIK4VIVaHKZX/qXR6Du3xuml8IgrRQJpPj4svlQ3wDd4
PDp3+7si802bWaYiM4b3qp8F7QH8DeaJuYHF24oiRvKEPUFLjP8x6vEYJ/pY+wGp5wbnemus8gCs
d31RRVEnXUOnixyRKvuAjYjl37naLUk5pZOX3HGRVl3k5sYguzd82ruj4WIuJi8GA+aimjOU4heZ
MLQtxHIO386lLZysJdbfUkhYz4eLNz7rkqoVdIT+TLT6p3Sn125ty/qR+JdKNkQQ3X0LxR5HBdAV
ANgXa10Sxf2fJPnklmWlTvJsl4g0kjVBnDf9lih0dyfAhkVV2CEPyrgfruSUsBUiaOSxGmSuCzLG
rrbh+A3IQR0wFzSKKEgH4gMsQihCIUOSMEYSapj1YqJsPXTchFUloax4ENnNn9wIpXpv0eK+oILR
ce02C9N0wc4cnf/RZ40h8i/9ftrT3Y+ptokfO/T11GHOtI9KHzrjbT4ZnjHewUJvhXlAkbqDUOCW
wUSyfMylwApWreKNOHlybjQCuciQ8bvmd7x0H021Edf8DDKGVLeKeQzIBSytYQVgtkEDljBIvEyg
kHjpLr9kyR/cqQ+gqB0S7N0BStBf8aeY+um3u7LPFk4rpAn44smez9dJof6xbtqAjOdutN120uer
ONLtRf8T5baeB8ypCXo5MteHL7Ex8CXwF+s8M8b8ubNlyVlgw24UAf1YuEzVE1lzYhhem83Mi8BV
N/7i3i+ix/rt5YmR8ctseEJcCJ3gpFvDmLxpSP028MXcrh1vwsMvZFv4gEW4HLP8o9VbbJpv+JPx
YDakTBLZIqCq4NOkUgYMjrsD8Y8CxsZj2LuCc/nohymIC/THvBBg1DrbnsEvftZmnx8ULe41zEJ7
853web4bz9nUqo/aRZjTRTRtUloPTt61thAMZd6+Ms2w9tnb41JxMtImja2thvxNkgdKmBAvV/1t
fq3FwBTFYKG8F15Qt5WQ24NhHFjuAijL3oQWjyJ+FBAifkaWodaP9TBo3gLFXl1AU39uBA8+jEHL
4evfL+LzzQXZEE4TANejH5KLqMrjz5d02NptxXUe1rl64RKNtajjIOn3faxEHGxX+dqNvfPspf5S
wH58U/bhZng6HjPxn7enpeTDVoL9iRBgW9jbiw+rmAThmIS/LuwHNm1tcuAyWmfNu3cPw/11NwB3
r+z9KJySlEmCHLcV4PQo3vVfK/qarvZ0idzWE0ZYVwYUBAJrv5h7Y9wrg5gAvbRkzFjLyo9ttW17
t4nkDbb4fAvmz9HlYCCRXZ+0S/c/X+cpSBVjQv5NRAUav0axKXTVOObr2ohHTN4nWYUCMnsvvQUh
ui4Cn0CFlytpjHmktNO4kRUVNLBIoR72I9IaBbkQ9O7m7MPweqlPG0M04fHwIfWVa6NX9HlXkLez
flQ3k3g05OIEe5pr9QIxgz8afeTgA7dZV7byhr3Lr97zfmzcfwkn7V2Aw9FExvCtRNGJ+YSX6Iqz
nAyi4udWpMJqQSvUD3vbRyVv1CRAxrx6Ixj9V1fxaBghvkNbRbySiVUg2T3rXPr/fah14D/FjoPa
Qy2o6hU+FpwUn1ldIAf4vAig+vUGrCxRD1EeRmq9fD9MSAh6kN+SnIJLFQemLaPncqD7eKfRYvOm
GPb2GAXud+m7CA9wOeXiG5yVWcSAvcfiV1b0gupaWmlPh2Akg6ljy9n+3yxp4slxhu8G36cASzRo
fO2E1YMXG9+2LQbzAWZRdHXBZL2WUVNGhLCZMhBGyw/YzuFmv1VXUFSF0nBW9l5IaP5Dk3Zv+YHf
NSxnNr0k8thXPPCcodG1ZptT+8yHIYzOwCIt18gQCoI96ZC1PYZm+x2x62bi+HnUevqBbYxiswyG
qgJ1uf/zps7neO+YlGn5djU4262+wvogji9mUBmLWNWEhwkDXKah3LJdwicPkE45s1CVkmQ5hFVO
N46X0SfAOhWVMZDDiUrcksJeDCDWzMehCrwrddpzHxUVm2FCHsV2DTFmroUVh2OF/x0QAkKv+xqP
c+r+TXjJM6vb8Es1JkPx+CkeZQVGwd435B7Ps8aZq6F5NxmYUnu4qHXUL06l25LubuMZWtt3MxfX
6I/1QngeYSAf6tWNgA/nv6RnsAWpWk/BoRQhZE0og228MZaOVvTnNzPK2A01AOebdc+wmRgmN8Rf
gDLqTc9aB/Dffw1Ls2J5OgUzUsnhsYalKyKcApOH9gSToaLBQSVCoqRd4GY37+w2VUKaXrdNw1Cv
N+dgrjRojgmI2rqMLkup00bC8uYw7z85VCvmVt2XIJ/BcZIfdRpHPHypA7GrwA/0pzajKoA7hKUE
+0UDyLcSaSaUWgOF3pWsDYRG0sBdcra3sXJsMcnHkpaFG4ZGPuSlmjyoIHlYPEuADXmKjn4GfRLj
hlvFWb6iud6a4fpF6BqGaw2rMOB93D+doE0KAPcdV0At/s8gBmOur4F/Y9ODRS5PiYO5wz3rFRDC
6RuZUzPUKlt8T4CTtEIruYT/BGx16pLKh+a4W1wH/jvEhWynAkr3ERYpJVzzy7tWoUb8mK0hxkw6
plIlHMlTNnOGS/5CuiBqvZpReOy5dRkM06h1P0Z1l/TUeZV1NpD3Fn7niVHSoVIgQD7wOIQIapFx
AHgdVQu6J8N3MOu2PufhYeAoOoasP3pmTX44L1UrTnV8xgXaD6wklLguotwMGhR8Pd562NxMzl6y
IDa1h2iuMui9FBqIC72CB9jkjKaZaHDhgNGXiGTY8RhxYPgZPWp+vkTvHhaNgegocLTJwqD/EQ+L
7wsP7UsPBjWiq1IvogRMLAXIltEaNhXJEpWgfnbVuETgah1CfFsSU9m0Ari1h9LExClM/NEE8Gs8
7EIREQtH6VTSMQrmJGg4v2DAs7cVWryAJ0Lr+limHAtvux3HgmuaJ/qN4nR8XptegVoGL5poRPwt
wS03StyuMXP9x3j6SDpSZnmrJcgiv8Q/F+1Az028IJ7kp9CM9HCNmEXeAKOp2qOvr0hikaxKTFqE
tVnuFa6x3ptsHD7D9kOX5TxkQ4mXAhdau9CtsDLFRvAta4cjcth5YH91pE8s9h1sG5iqgLh7bJzg
PIcch3tElnryL/rOoVbAyzIA2FT6dostTjUNfCL6uPDs5tlsfG7w2b4L2+DoFTxp5ihhscFamdnH
bCqwLD6/bcEhvn1crE+wMi/txsi32cYsLDiaUu+a4xPc+zdUYnbbanHBrqoJ5az5j0m47/jLYTYV
hQwc/EkoWgiL9RDnzU7BdZdaVhVOZ94T9Y4nhAnSbsyG51kfivvE3RQjQT86FrhJzA1lVmqQyoBT
BBtZapx9jlCNZBnI0sd1jwn1Z73aUi2KVuCC0J586CmwBou8coQpKxTtwxhuJ0dMUL6fRRXJpKXo
iBjt9A7x/TQYWGVk6Pnr35aHypFwi4OLOZh7AVHhyYD3iZCzAKvVasd1Hq1VsAx4TdL9BHCAe8Fn
6LKxp5hetYwsE0vVvF+ADvs+9JmbrItjp4NI13B/ldi7DgA/YQh+0LRW2AOm24+XZ65cNxqnlnoB
228gqPT7DpiZar15aMVJarDri6QR+3GuAXkWavhhVzlP3rZgZXXhqzf9M6T4ciFLG8fbt2YilhnP
1dJeJDYIvlVNRMueZbnsON9F0A3eCdvEM6lazilmjfxY1mtjyvcCUiJqanPTkvIPpksHtWve3Pa4
g5PqQUGX7EN9xO2CmwxnaszVXNMAk7HcQUYbHEN0PQbt9bKfjzcMIHqPIfrKK24H47P1KinbmB+6
P0HovNoTrvLiUgy+oQmQd6s5kLrAXhRc3TylZkn86Nn//J1mBSK0o2htOSsSM2YBIyyd2vf0r5o1
WxQ/SSOxfvGRJc8UqaraMvnjAZ6b/cnpqUZzJsv2jD+KcPzBHYRkbv+ScjlpxHEznnWfW1EwSk1C
MLn9NQFR0XlPQfLmZoaX8d5ILi7mIs6V5QDg7mtfaTFw//WasezAWJEVHmN7sLpVs0kafMjOcwfL
ubfzlYAcPaXNVFjeeZozsAHUnDgGAa+ODJV4YYg1ZOFebqQqdPNw3PJp/iG+1ln6JX0p1PQWS0wd
jFI4SGL56dWTYTLycEZJSyfqOYncd7Oy71kXTf3zRtuvsm58ZdSQO9CkuTw+MEfViO6ZiPRn6jbS
jiWIlaWdK/8aeoXUj3Dax5Wh0FvqHtvf6ae5l+mt6WzNQx1Sx1WCNO26boWrubXVu+tcqhrEbCGA
/mVMsVZGyWFEHsKLu7efA6wRUF74VhY3wXgvGfb0ZAG88NiTaCTB8Kf5lUtJAlDzHyAzRhZa+rI1
ubaZv1cZCn2hv9WCcBb8SrXDeOMmpRvPavDPMCHOlLAK9hWNmjad5a6/U4F+1BKoZ3KOBjAFaQju
zuMXp/eLcaUcM0VQ5kiA3KtOapaNwygud6BJRz+q7dOmoAd4F7xBAfJjYkvFtBhFpfTJWa1goktG
VUBm9TXdtWdb7Tz+2T0wfV3KcGgiQhAW94W9u3iWVrflbRJoAI8cMWaSSEEjhqkDdHLsPvO3DxF8
kHR/Y4RhBYbMrr2Wk63vL56FF35WQUhsWzfHkzzkhTC5OJtHUpTQdUZ5a9w2lWtFyNximx3/nXy7
BADKO00GsdnFzDX8+cwifChvMSH/fL401z0tkX0NTQlNviIy2wTpMQoFZ79o1p6JIy159acz37Ua
u5h5Mqzfn7ecgAc3UdAUFaEI85EgedkEDz+WBXI4ruohblkBgHkZfZ/QWmDM16Po3Y4w+mdBTzuG
WoJB2o6UxvPJA2PIQDIYLcOdWHA50jKfZH7681xedT33xC9vc56p4IkDkjNxpiqVErBZfNxQq7Bm
1J0uPKWsDnUscrZSy4JhrfxHikx/h8Fu5PU/HB4w8wJpt0Z+w7sgpbC/bzrOc7f3D+wGpxH6dfPS
0YjldqpG7mlgl4BtQ/5tHOaNgvrRolV/sS5dMQUtxjopnm8GUdqMthcTJXKAF5u85CRvceDXLMHa
S7j9v0nxeJuC+yLTF/OVT/JA/EisIaT1iFhm/vtCSE6vUtIqHQqlYDTUOwBbvsDOGHT4sOGsfcDB
bxEAUteWKAfXy3vxiKI0+HOEp4U/zVHN08VyWd+I/lvdIxyAsRuglmSoyrrqRpSzYunAioqIxuDG
nr6oVj2pv9CfOrWSTgKFYZMf6weK+PA8aZWT2zwCMEqD2oRbGo8zlKqJNji4TM1FkoGTkLmblosZ
ZIY4TF6TyLYCZOLDwPeVFvRdn5BeKDbbxOxxZ9ZAG2oQ5xC/T3bnnb/ogR2QRFA8ofeA0CvVgTAm
ZyKZLQNHrGlI/hdJtTOZkDUT0CNxQMFVt7PNANVhJIQ1LdUaqhbNgHfHfRvLNFzpjWJBx7nGBRRu
arzjAGnVkxU+h4S3Tr5JHQ+HQxwWEdr/IxonX9Vea8iEpu6Jt8Gqtw+mt8CtuPEywUyOgYJf7fhU
/XusBk3dSxKh/ga8YpBb6GIJRZ5VU/nCK3+ckwyyNEixwv+G8CYB9j746iYQmpvY+yfmw/Y9RFmm
oQE4dVqcsBw0BCfSiHX9Ly065yZFZ8VXoNILNr1gvNgn3Qdyzdg0V0wA/fSZGQIX/CcAmX8ZtpxW
0V8l01hHCNa0W54I0DZ+1x14EmRYQKjCSZyNafwWtanFoG2tZcl313al8XVhuQJ5KiO4nkag3TEP
LMxQK4+xY5Lbg51L8UDOCYRgFobQMrPCEPMH+34yHT2D/0PtMwwX228yUdMqRhxsUqj3UJp9gzAg
Yyyi4XNUZ2sX6rcuYwTVqn4kvHyCELHTEUdsGVK9M3Ha4DK3CI2nP2wX5drHMtemapdQ4E6xQ6Ie
JaUjecAtWn9FagMwu4wfEbzno/sXn7VR5wiFmrjCYKuRMH/g6WTV4+NIF+8Pa0+1Ic6AGMjhUGu+
X5D6k+gIEzdw6PlieTS01e9T/hI8JMtx5+Eg8fSzx8Ymil5HUTzP2d9Pnv7xMuOWV2AFjphgL+bA
ucKzF7C6FsatNfejQHCLkib029pPzep9m5EdQhGk+IPrKRII/U1wJavue0zokjafhZOUzBmwnsMy
Tn6Rpi+4QjhDZ1vOIIvW+pcBmDMdZvLvDMJ8SHOEOkopFw+6jcrVqk29AxSqGxqw6Y78X2L5m96c
NgR2dnMVyRx7RPVkECZIkykev/nBHJAkFaCj3P9JzTJesS044nbdOthuayZW5pff+hvnVkn9w0Y1
ZF8RxY03shbLiKAar2RpqRG3/ptMp1HY6anwY45ZlDbFfUHV6u5b5XPnR1AJ4iVUIEPK8lQTODjX
F4+OOVIJ+JrVhVKeLOeHaPTLt4Md1KjTwl3wT5GXkbkRISS2GTGTxuu8zvjODE+kwoAfeya1Usbr
d7JvWkzIwX1Vc2lYCW6jEatwUo9oBPln7OOH4kt6ZnNl2E+2vKzpzoI8f/Pb1x/dYGPm1WI+g9+B
wMK/Fz06oC81TbkAQiLDEx18fNeFyr4CbfLe64uCBnB97MW3wjPB5WyenEsSx5wn6wZ5cBeV8XOE
msmCA5n9VBJmTVtMHBINA/9WgUaOq0zd2FYXyzYAKPfwqflc4uq1+GOKCiPHUFfF/K1Gj/nyOHNF
kMXekGzjqBfwMMpCmQBqA8moJeD/3rMLIkSSbphJV6UZaiZ+vcb3eo3xLPkV6Tob95yWStkZYpb6
v0hC+ha77mcoxXJpLbe/S9cKA3gsb324wws74jHc6mcDhz/SQ8OduOBvt7i9KTkhMZWPU4KQBIgT
rXBuyM4AI9Imcmf7IYTvk1SpYWF6xMRnmb3f35W8USQ1/mt8LU+PjEtnJme78oAawT4mLqdEjnhy
jSKZH7fdvpRosm4Z5GEkHcyItWWrOSLYrHli8H0MKGa6vroX0t1VefSFtt7IrZOBoJvhPdje7yJp
gjeXMDeWjKxhUpfDyE/P68CzAo2wS1hbF3c4FX8XknMxGUZPAgLRCVXXVSR/L2Zjs3r/i8FnsHR8
Dq4YuvIWcgd5ZF/DYRmJBp7D6HSXZGZpyJGbjyf63c5ngUiaSFuMovl7I9hTj2KUlsKA39YnEy5Y
Hq29vHcXcvUCVPzXPoaBb/UYlVTtGDibBCQsHNGjoRCHBf1jhjn+CbimV07H1Q/HdfgE13ZcDonj
5mXCKnWBPrmSRUbeBRrImxOKRnK9d84vgDzySHLFkztlnegRJZl9uVf7+VMLnLaolnK9W3a7CgNx
RUCZ6iYoXWo94paQAmUfi2HtqhvijS7R4RHwVF6QnYJMMW6febtfv5OeJ/LNLyZVV38rQAvMUadx
I0U5cAIsuAZCD4JHcr8X4omAqyo7mQ6hzTqjVYPXH3HWCaS4G0SuamneHgNLnGBHJsLKuvv1aNjL
BMiBoULiSotbwblWq5GagqAzDx2aEJwa4TxebDa4Bo486xzIUuyJRjRUJZ/QtU9X7050NVgcpCxH
XoMfvTR0cL5iA/EUJLerjKcY/Mi0HwkaHy1fKhNpuVsPXRvBbZ1nFdYK4fI+GD/PAghE+bZEL3ew
NNF2CWREgVt1JC+5d+6r/E5qhk6bKG1IhYXc0v/bBI7U81sWlK9AT/zfhPpqLW9vmzIKrRadjCLn
NDZSf9ByO7QUHlLfj0eSbcYkf08ySvAczDyHC6d28ovxFC7oPe1q8nvXniL0nqa9iH74T4SIV53N
Pm3iXHmamVyvJ6cEZRpTATQT+6mUOvd1OId9Q6NTVPf9AXF7Xnk0p0RQx99GclIRowYaBPWvdJsF
TzfnjroFEJlee/Q+73jJsLYN2PHVicGdlyOYELMBdp9cBYWCYd0SPtM/M5F+4+sGedGkHdUu6ljG
RNR/fb3Qqr1XG3IvNOkUdaFlQ+55R3MWh9VxwQUpmpo7jTJN5wazPaNOcQ/Xd9xfwJ3T6LVSODCG
MtGf0t0dTkgOQsZid1gNgpH+EnBsLGpyNIL2HoaBnJuLonnddo73wcsPi+f+/UIAISyslJXon/vx
DXJi9Mh1uL7EZbK8dYumLM/tDxK/zHrT7e/pU+XiwO3JOizW0hH0Brq2B+4VQpAGBmd6fDZwoCp9
toK6KytSHnfyHnhtxVcaMihzaphxROnj8PdjsoLw3+pV0QK8YTne2S3e4PFOx+I+xud+q/76tgF3
+5zvmW6mualBXLQF9kPzh1872WYA3XCthgh09xqCE6KEhhw0bDCbvTdxpxZxWEyDuMcB6ofTHs3Q
xW4q2BthSNjxiL8ANxoG24W7KX7Z2acgoyRGoWf30izOQVntgDcbNy4FBOA8GM7vSivSN4XgCMZg
wD4XlMc9C8DB2+EkalF+8l+9g6RmOctwEHPvYQcR7fRUvNCEl7mKKfZc/XKqAdjNGRQJjAYslj1+
ZLGb+MYkEqQk5eoN2b4sN3w5pb6d9PCGiYFd+WsHdlqh3jUe+HSjdTmMWyXrCENrt2kRQCKFVEqi
qIx/yNxH8718S+9alaTLEKiVRG0WgEGsgjZ2Gl2oBvu4Z8KDSfth9ysFOfJ/Jb75THISQEHeErH3
XKSB0QlNARm6dYlJSfcyCp1HYjTeUhLZG3FJOu1VVhrHXXky9ilXDtejuXbcBtt5RMqZbd3T7n7G
dkxX019U3WRtq8TzhvzdYF5ERxdhvM9/LFyeVsb59/SHIFDqikZ/XTXWR5nqPnQrYfkBftfsnTnS
S3qIgXImy/4ITrYMuVTU87BECURNTqwPgsYIUFkbleiQPxlmVUwYMNSoUryysWbFOGI/OycrmYg0
Q2SRXIT5piNOoYu0ShaZQByeLbytfqLOMNPSo5qRbf7fjjr5XEJdjbtH7hm/ufpccMZHypptXcMJ
/HcIyt5g1PI8c2seRxERgMe9lPiK2Bp09pwBqbGTQxoyeJlDOHCJOIFFaffDEI3q+4gPluEZafcz
PiaXajRkM8HZdtNlpi7fHCp/p3FsxtN2K8/Qxd5d0eUmP9n9VgTOCTnaCux0QuGV7hvpCpow4Uol
vrMX4hS7WQwpK+h6XIZoINOLvX77BYvZQJLQwF0HkfFmXfj3F8X9L25J5n1Eh/TDNpfiikgABeG0
xsh4vE+R2M4cCeWu4568LOt2U7TBUUFFzsit/rI/oLdRLri50xFd57wdQkj4a0ZY0wWpcJj+y4V3
+CqYUQXwD32nDuLVFHz3ZgBegKb7ii3DltBGi8pSHF4QXb7JvhzCURQT7Jb1SgNyhNQNGSl7IrP4
syS1fAivXeujsUWxATG4QkO2WqfKPlm13pWqQvXojVgjgEr1GQL17CJTjR0KosruK7nLRi7PCej0
CfgMPyAMWGB5F2Cr0vup7sBc5tp+YpbxHjJhhicUu3bdoOAKYhK/IFKdbHRoQOkLJhv/0EP4JQoJ
iRNZVls64oOlkUurMu2kWeIF89wpHAkEuSMAO4rEg3UMlXA5wWtbXcKnoVX2UMx0gs4Sk5OKnjJv
gtNY6QEQb++sRiDRJsiT5Vsh5LBe2E4X6xznE0zga5kWzrF8p/68BAvYlg1ZJ2zteX+di4fpWjKq
2E4eN8+81WY5vovGSCIoOM148XeXSZZhXEFsT5wBAAWpAzRJ1fWzipqAnE8yHdoUx5hmAMf9uqA0
jLm4GjjTR/slGzNwUvYMYCYJjeXqPnON3zO/Yv81zAHxYWsTjcwqjEZQQoCx44qYZIKbdf3BMWlQ
2UGzkCkT9kd6pGQbN/hTMLxmCs7MpgVlPXKdpUz4OELN736BrA7TdSa7N1Bv0dzc2Q+ivxASoLjG
snL6HcMCXVhXfUITXE+sL4KWnuEI2XoWihfMo0C6rJBshEXkwi+EHvpGhpiIDHQJf+80Zrdk6JOf
fwSp1OOOdudwIi2Egrnty2BLBj3+uj/l7LGRdLM3tzNrS9trAzGQ8+IXvkMQWmSKjQV/8VQ78ZPb
JZ89Z5igfsfyWOacekHfx3I9P8vx+GgD+g7F7iSD5cIAv2sqyVTsUEo+Bl3sKWIdrAyd3kpOCI61
0IUKnyEHO5WHbgZAWcmZOoVnTNdAl4g6rqw+LBzWPtZYla27F7XMYF02Myuy5WLe/Fiy+iqyYD8t
Ay3ZzX3kFv6siRg3uNmXWuJ5il67e2K4bRaBLRg39+FGcL6gSR8rMZN8j+t0Ez+5FbyYtIvDYLq4
YFWOPxMLziZhqpplSdH2JJnMct6cawlptXGP5xeGOXWRGhiGHGDtCPCZa5H7lcI6n1xYwpYzCqlI
rJMeBC2qMTJBUyxCuW9TZmnbUAcEFEsk/pw3eeyQI6481nsbaDxLXKErnxlbJM42Nj7LiwWP127o
f3EPIZT4zpUOF4OpAjLNcLJhk3xnEut6+qATOBwRhlgYCIKwLDWSyd8S1h0K9xMZwqLRSaqhGLYA
Q9T8APcWH/X9bPCoGnhLO88nD5ZRP/ciOiKQegjIaK13+o8B/z93dHBhB4x1r2ov0qVawxkUMru4
nG0w8mIxqhFYpUyEl7cZKI25GuKbt/et/B0aLRNYkWPG144l86DBcA2lLMJnZ5mZdx3OugwuabAk
tq8r8l3pG0nL3dOoaD5QVXsFAupnjy7ch1Yzq8wvfaiwHvUx0gkcwuJzMO1Yq3zxt/gt1g3t+Azm
iCX3/GIzPwGxcUvL9KUm7dBrGe/BJL5vMV91Od19f4PYbLUsx2zWeFt8BbPOMNl8wDTt1Q+UF6a0
dnusmbn3v0iuEI7Cn9x7BlBQNEzs695qafzfmBG0c3uWc9NQi1JbjonaW+9n03ta7iLqvXLbbRNW
cs/rUk9/Hb9o9o2Mb+zywmwYh0ti0TbReVZRBTCYz42APZ9A2RuEzSZ5QYXv5N7h0XXe8sn+/Ziw
bNNoVjY9unsTDtLc6YaeGQmuHAYUK5EyUZwbLSfFqRj1KL35BkaaieCLsWV/C0sPJCL08l5vMtaC
ISeEmR0Ua63bhbKZoN1A3f4xqa6qPXvHXP/O29DvuGq4LxLl9WlJnjxr2obQC0eYp6wqUcUiKHCW
9W4CDUh4oJ14FDUhHoRFrlNxCqbHEuAy93z+fNUa9IsJMxMDnJIwOusUqz9fInoOEOGwteX92m8u
Xs2GB7ObCgs8Vl4/Zq2Iyq9m/7Xa2VDBN8WmclAgq9aKTp3es7+AUOwi6p/6Np7Qoo74QJh97E/v
ZHw8TZaO2ju8BRmVHjsaA+l+mr9IRYXZ1kVgqXZFEOSLFrUhf8HyXdhcfJP8hTTAD8uhfSkGD240
37PLBHo4Nc9IsEhlPmEkWN6kNs32J0a2boXUswCb8cp1v6O7jcrfyPntU3RcEH5ZQUaYwHUQVRHj
K1S0fwYbidzyDg+bEjoPl7qhYil2DSZeSWTXwFzu9OmiaZlCpIYu9Aybl89RHPeaFel7h+7p9wvL
J5WhClmBjlYIs9Y8PFKyII+8Z8c5/XgadpxM575eHjN8k/XUhV030C1ZD0asTsp/WeOSsfSqHf9N
Kp1JErPv9GX2uUPZUuv/1mm4fZ3MHISx/LAz6jS8E96chvyydxGnR224E6xS7jfq/1ZS5VpaMkuR
Ojgl8sr+CvZM197/3Iro8wskHs9rWx0/5V0c/goWJZbBVZ8FVW8lXkRGjdDuPfyurhsd9sWx9jtC
gn9nCiVcJO57oyPCWUwckgsIl34jydS2X7vvRf1VpVsVjAVSk4LrHIr7rPt3CTmq9vSpjSNHRwQb
NPaiE39MJaXxkq2mqReUF6iakPMKW/ldFwUq/F4k4azT2Lh3UGSCCU9VB5iQns0cKmye3ajTx0YD
n4HgsmKtXcO5dJupvK/FvVMmoFVNgeO+1wLD2lnotdUsv9an5PTGc1sHLZPRZa1CJ++oWvaHEx+v
3Pd/vxQRKTF0WJ5XEOCNap8SFAo/DyD0eTQy7vmgV5I6omADUab4ItpfOfVZ9wOvjdpiITfwu+/c
Bza1rvroO+qvEInuuf4Xv1rpXiaDvALDlhIFvH6vvcICVPONPMw9ox1Gskf3kPnpvFoUqK9yI3Ii
7CBxV2E9EIjWvVVo5+pRtYvLAHkbvV/0dGXHZb4YBNftIIgcl8D5O7/1fODm0iA2WkEE5gd6y/8R
QOEyu6ZPt1O8GKLG36aBevIbFsztmQDa4YftWFzhkAcLnIW2st456EaXtpsTcBGa9Wpqru4mSZ3e
3/lc2E/eeaSyO4QlJZjYLThAHeFJ/ZoIDrkWacwYSKQ1S+SIa4KrkNzeI0Y92NAzXcwcTSocrjth
AiEBBAcBd1yFwr5xKzBJNkfqE4ishUrV+kdEtiIy9egHk5VyPa4qyKsf338TeG8CGJCI0MlfG11N
5/vDVVjioMwWiCUnb4cG6otWH4xuY2w3vE9uRby39VB4IDnlJZ9l2x1WzcBU1c7Vpxt+RbTIdZ/P
lNP7f9GMKLrKlpX3oBK1dYmW2ftZ2tKGXTD2rJhYkzOmxmk+nSYE7YzYlOqJp5b//32O74EbKLN7
aUynuGfCs8JWLu2ogu0TreD0A67MrzR+zNWlWSnKW3Pw372DAHGpNl1phEiQvD21vTF5Qv6jCLjq
jWgrWqtDaaHpjDuZo92zSmQ3GhMB2BwmR1wxBsNtQQpTldYO7QOh0HiwptN6hTyKqmDV6Nu+Yj5P
BGWhvlra84W823QSSY76Z+t0rMqn0tith1EvkYDMARg+K7+euhvC3zOS03L42lgGW3kEdeT4ozzx
FqHL+kH7IPB4EDXPw1Fws4ctCqfPLzT33iopTPSK9nYmASiTHC4H8U3Pa4166U3cjbYZ6CkPgFc/
QpB1+TaFarYM755TkvJw5tWCmaBf2U5oD90H7g6sh/jeeNGsgKrIM0jEbYyn4V9J8hVuNDVlPKpQ
bTPCnTFpGuHeHiSzW4RI55qe/dgoQW64OMMtxchhD5YIqEuKNTkDA5qyB7sSmvOTGKntiE0Lhft0
2S33t/xSg5SxV1izwLgE3f145CSFENB8RIDe2F1yhpn9ty7Cn1qTgvJTWmH4s3WwpmNl9Qh8dAPj
klu8brUXcz60WuVPkRIoOEtFVXVcaHX5a5717c8S6ARZ0i+Jj1eVOrhLK+na6QBK4p+qF211MuUv
iWnhjG5YP/s+5t4m2rfomQkT1ixw06zzZoCj1DNL/jN5qrqvn4hytRI7cUMDRkHTWtVG5K9m2tJk
D8uBRHq+Ukz4Q1x/Pl2ZH5vB34FU4BSON8F+g2PsFQTB8VVKAfm84N83hzKOq0grmlhzyMCb53Cf
6RMYftC5V9sDVVGmSF/ntQcWuuV++HFk/NJVVidxpVrmlGGJ4H6YYVp3d/1nQWw/751BZNDYPuHM
zZnfLVMlWAPDrR9C93yBMMBELtuIewTc3f5rDnjLAM48qbVBCJVQ+rvUy7U9FGNwAdHBxhF1ubZo
e2dtO0EXYv3wcxZEv18CgytBYM2t3MGUvHVkVAnTbRd6aUCnuTPISa6XCbx25fvxuuYqZ4a+7ZDk
MqGyoDUVqLVBVyXiOHJvmiZWd/6yTmG2pO476aT+MlCWOhxVBlW5m2MKBldK2i/NkUvDVOyzW9d2
HyXWe6/Y5Mu6DUVUtad1Af50wMsiEGOpLZxfFn6Hsecn4Vu+4bw1wS1WAYdboxTsG/WUQ4asL5b8
e38ABiAG2w7VoKD6gJv6fXqSzQ4nDzQn99DgY0mfSYqv/DUVS4ytTQyboTF5Jkwg6LNIHe1Cl37c
pUHOh3BEhNDIBi7wg/PvfqPvEj6FqTQNdnrJNofHZfdUisZUsd90XwZdcLpcB7CWjm0o2LmcFR26
CLYlPuWelOMrEE49w9dvXyMm/w5znlO/ZOXY2QHB4FbsddDmqvxRdy6GmAXK9svzhfJ8bUEbJ3eD
mkPP8jWjAYOLiOS7xQnQ9lYk8mOw6SQce1O0aUlvpZjGSLPI8l8O2ZeDfdFn3EyL56o5EnCJwndK
cnKTh0xd9+XDE3Q2IKRcS9fQrMWAIEfIYC1fUrR5pDyEhwjYTNtn8oHO0plIzauYeiVzHFfuUcaL
UItFkRmHt7ZAF9jSW5b6l0bu1uGUUf3dS768hf1zqDCWi7RdhI/shkSJ1jvhI9gTt6guLBcD9jnh
DzaxbE5kTHoaj6/XxUjlMJwI6/v7luv+DcedYpYi7jB2Yg/t0er4+yMxneAdjooXKjpl75kKDcDy
I4sh8CPj0K8gWE+cfX8gFDs+8jNOq8jm6ghfXlCotWDB8rHpmddNAUAb8P2rQDNw4FzX8jpBvsiM
MRuSSAleM1ngFZw+H/PHT1p6lCsU0dPCrjJMuZF+oEaFkq3u9LU/okufRwNXhOSrsTZDTo2idn05
fhauxgMw0piSMvmPX3kguNwIfZPfriYM2F2FtCSnbMmr/QsgEqGZ5sl2iG4BzYLMUbYoUo9cTrZM
SNm9QLx5DZFRE7BJgjCjuSRGoby2a9/us7HVlPhmvR0ydfdgLy5E7TriCEx7Ri2vLnrYgoZaKI1S
Lr36odYHDKFyONCIqyI5hpFRwAuVJzMaNQHcamnfFDQxt6Tt6LSW9B8g9bY1nT0EUg6zAGn4YlLA
tMZcejLzJT1l/CO9dSQUgvbpD0+lHbAey7QUYvKduqZUcSQMdXt5jYtNxhA0lOHoojokVrqhi9OW
pXM+QwntOp28TB6Ataqnw/uWlx3ooHrLOmYKGUNsyACAE3PiYDmtdlcgRKt/aXR1NKfBxkz/5bcG
sx8XRro5YAqlbKB3UF0NwK2OKTd0YiyJCAv0nsPRS8v6lXhP7v6Dn829/dri6tVlwMXqckf2rJ3l
ldvzNh+krojH5zVhqb6QMjJOQrYvG1IBupMs4gaqvdSLG3raGKUfqJ8VZBL2fdKKBufIHEYJlmMX
8XKyU7KWJSQvFA8OwrEDZpQ93/n3/hzyZs+/L4wHnDlek39jBcTnrJ8sc8nuhZxaaQ3YNWfQjMJp
Sj0eHv9qYnETYcxoqTOBlH5w7liGMDFGW7+FPz0HkEsUArAQJtET/jieOdvKulyuIJZOGr3ZIMHW
QYTJWcerDZ8Za080JEaWXFySl50/i3WqMibvpp3GGmqDFFQKcX+OuHjdbqHFINGqhPlW+1SqE0zX
3kHykoOb/kj9nASuNjOavhvFFhTh1h2YwvDScBsL3T5o9kce+nA0D1teqS5IrjnUvR9m+cKdrKfS
qpn7tYMnxoWP1uMoVxb4x12sGpaMt7k7vDS1VSAeJMZjLuCE0TWsE+bYlwZYcjUd9oNMFvhYfMYu
eKrA0KIsAQd6ahzsOuBrDN1VngUH7Wp2CQMYdbWqFW7/d/d8P3gF3emaoscbgc6h7D0vnoqOjWXb
P/qDaHpRc+Thkn5HVKHEgGnfsSuNnl/Zx+1WmjOBZCyEaLwy0wQ7jl12fcuZur5Kh8Nf5bSPE05M
W96XOVs76EVMx/OtdfUHm1Lu9vnDEdVEyFKQWaa5JnRiULSjPyBwG90dDfqZY29IsIt9sDHfSJXq
OgVwfPtXSRdlM8Uax2C45G7An0Jfo2lGclouibjuHvOQ0l+UKY5wsazy569s7mUw0TIf2HRFrzM9
x9ZIPNHC2v+cNw/LUOQChSrL4Ja/EPi3XNnGayrgXySo/jaO4WCSyuDUbha7SYec983gkM3oBa8r
IX+cP7SwJpydx9RQbHPBCTCj7ffLDtHyQj7sKhIVFvt3gRaycu1+up2yAml5Ynpa82L8hJV2y9p+
Io++QTyfXg73xUF1kk6QRu/3lFQnNUYaPN4pwhUdIdOEdHCxqcOz2gDcBFuzthfVOF6ScJM51iVV
lnydp8ezoTxme+r7bpO6ebhA/M239QQDBJMRM3a+bvHx/p4X0QRovR9UeLLEIx2pWR6xCNvp7ti6
B5Nfm+44wg0K1CInYJjEbZLUKwtsUhdxgICYzM+8QH+3c9cSrIPAf3wA8Gbl+5sWh50LwCkVaqZ2
GQOdlTFqYtkZ3QAnalBwQAeciKONpFXaBfPYYmTlmbrhDvSukNaHjmdE6Z+HBWQ6qk96O3LPcXPE
6ILTVWvzVyx2gKQgeJw/G1s7WzFsR6P3xaaYUS3K7qzRmEwV4mW21bU/29YLFHIpDn7UwAORzfsh
d7ASVDQCem7FbWWXwx8zBP9Z9laR5N3GoCTBRBLz/4oK9PKQ1IkkB/MK7J9rpOYp2gNTa0+AX9lk
Wj2jMGY2aDtMA4hdrsgVPLDfAKErhuJuXxcUERo+fggt6tfKjSD6aVkl2DLvv+JMnpxGZT5chOE+
zfdTQgyA9dKy7Aebb2GOrp9hSVWzysrk5pfDBO31NiB6VdtpJSNylESaMpLtvxMdGw/ulH8tbGoL
RcQcYc+I1uWXPYOv5K38iAldqyiV52XKOki4ymFC2ifflk1GkrZ6VHJRojIGfSw0nn5k6vGAFOmc
2pfD5sPyIlT1gVGBNXVjZtdjpMSvatPJbWTqyPVod2GW+AaHktNaWvq1rWX8qLEVkwLYWOeIEWrl
uh66GWC16O56UmxI35s6PeW1/iV6PsThS9dn7A1h0qb4zOntIwG0tjxKmoQQfx3Mb4IkMWJss5Fp
bS0okP2ZKUnO7kl805d7xV/INCmkc8dOnNDpKQhs0zfKIKDnzU7g3w6AarRvJTTBAeV4RQ/DJ3BQ
aHDdMtx9+jXQ4Z5gOAzJVrARSqP4Xux9ePN/tepJYe7Ag4i/D+ismv2IoFmX9+REnVXTGizvIn8b
xqSUzWZ5ZaG1PWCJbJ8nquOHuDJw4xUqPKD3Ldc9TC+VwyDu0KLMISUeI30QHtCxDPj1mXkfvNDb
FeRNFZsZI6PEbH23clNEWyCSLq488/74czH9VlPNqHTA+0KDjQZm+dqRJiGQECaAK5/yGsEMPf8u
OKXbEIaDgExi9U0BRQ4RGSXSuwCJGT7CJbJYuV6b69to5jx2/t/ZqqGiYUaOUjzrKbb+ae8mkp0r
7QuDipaLwr+6495qwv3ez3e0RmnhC2zLv2ntbUwHc8bprWpjZF+tEOk56W51crLfCYau0ryzYBGx
8OhJtrEBrDU10xzvuFOlbfDztMEIxC6n+zKr6/fx/kCCJmJiJA7Q27Ur70psTc/JeXD8G/z6XccU
ld5ccG5ZBBsIQb/m1+b3T1vMbrMr4mubKP0hVa2z7JxqLwjPnxHsKzelqG4ob9MriwrUHhu9ffed
OgYKS6it2Mv2mRL+DuthzuhWMoIhn6j5fjqmbZVIBGGj6qIJRQD/LQ4DLCy5HYKiU7LTW1nn2Aza
k3la/D1DTx5Ge6Ke7fE7/MAgqo4ELXp7RpHp4w7C3pVdEy7+UAdHH0ckMheh3CTjbo6FYWosbCl7
c3uROsXXVAtIVJNrGkMcUkTx/Y+rmYL5/J7bawJ6EejcP4GrVH9HsHsnB32HPmLbekhsVrKrr4j/
bvsSx+k8Wh70bgEiz/yjJkmjwB2VRZ5714ftbZSyhx+iODfnggccSfmtiSHYaT5wv4gxyAiBVIdO
QyTqpfdcrf3Wwn4OpQKDfq13cHrnCZPIE/wT07LwMe4zL/tS7trAi3vSEfaDJEW89v5ZekoNaKYn
4cmn9iNrQvcVw1SCbBq7zwwLhUDk5LkR8tvpnG33WtkMylewkB27eYWTkyct1zUf0VsJrr0hTAGP
ebkJrCs3vu7t1NYUIda5tuG1tugkkxsGWWQpM95zz9SAa74IpD4yx2SUyrVo6ez0OcazrjRyyMF9
6fMGH1635wYdKHLEK7r4iiG7eNkOjZjlm9/grWDrgRew1R1qZQMKQg58j/SYd7B49OwdLdYAE6ab
dpGkYv5A3gH0gL5ngEY+7IuwTY9+NvjOkXvlrPk4PM8QxlQW81Lep/1tdP+lOgn8ABcjdK8ut1b6
we3pWpF5bdr4mN8lb9GumrdH+OL2Nf58r4Irda8PSMaJmvGfZ99O4kjTK8yhxLb1UUatAE4NC1pO
MVj0+IZlDyXmI/+wssdSikXat+DJ4cRmmUbnci37Q6s6kqUdF86m+/Bz9JYdBUSk84qx3flhpy2h
uA4CYUtEuQNLKT2swnExgJzL9qPBK+cwt49dU+KkglW/V24MotxCbip3+05by/X5/w4KHO6OFJMX
87NgB78+it6IW7fu9vpDcfUn+kIyTJ8SXcErpby3+43yXGmiHfhte6SOFpBTqHfuRVchR4fIXmwq
8FdNmlfx2QxFt6YyVch2GjzHi52vXpH4vPgp4Na6pSJ1UGdMFrcBGfxyeuoO1g0imL5Fg6vebacj
+2irce3eJPP+yKQYeAuHJ5ZzEec4xzSZvxjTMkODfV2CqqKtcIbuOtkWST+vXJykEgb+Ov3NlUS9
18XF9dC56o7/Gk4+Rd5XKAzLhHDSAWPK0729KDSr/kwA4I9ZDS3FrxSdt2GEDbyd9/WqLs0ohDcM
pttU/H8I2Ip7sfl1rDK944RbZfHRrBxb9/kadv44Wh1Ru6FNZR/ayFCTBYBH5yg7lanwprdues3P
yQM5u5irduQrECXFTOo6Um+TVWKI56Et6a6RRERteqY/cMDRzVEpf2OkIw180rqUWMYND/mzCPyq
+5J9jByiwWMgZrifAModvwfNDakXOoZgrDW1L//3V/h1sXRtI2Px4Yyyb9ufVU+qllCQx70E4XRw
FuA1pWc3AC2qvLdA6EP+iHrvT7hlyksTJ6VoWn8oV+6NYKh6wZiRqGmN6JPmf+W72XGxJ7E3AWVd
3iWg8vs8BTBOevcjT0ey/n6wVSCWVXVT7A7em1so0dqQzgCZhSoySKEMKIEasBuOoHLTBOThS7As
g9x4L4ylcQGwVqRqRUSTbhM1Cdeopzd88KgPYPkBM0qzQJ9GLbyODLDmfh5gbXeFFwfl6wlJPZnq
FbMi/LynLcPQL3h9GzUUlYsGEp5DLiDjXcbIlh+8Wss8dytIkfpCOf9qH5Fgm2Ttlssbm0Na18dH
jGebv807qn0FGi9EQYAhm488tHjl9/lWiSXUhOuBhkL9k+JaVhLjiamaOBDoGr/SdmQfGgcW0e8/
QqEneaPcHqo+TL5anFig5C7LqVrZFL98zPg2KSFJzsP06C11R/MOpJqITWSGwEX+YltmTwYbFMM1
z1F9IP/YFjSBC8md6h+uDeLDfob56b7HT4BNRNYk/iXTEkxJuiGq+PcDJ/kdVwKSg787AoiJHb7R
zXuoe99FKtNyy8nQJjnG7YLFYkAUsXR6j0oU8pDCtVRCrR6PR7i7zMBg7Jt+36h3UCNFrr0cBh81
Lu4toQio1wwuCen4QsK5IuIA8QYjGDKLhgSqvP7MuazBElD5w+03kLbmC31decA5uAtwRMSUauhB
FmqMCfOOxXapA1W7HS/L7JlNPiJ4WZatDmeGkMUy0bvYorLqvZt5KSdc1t0WMDnJTYqkqmxf32jo
mbDwnZKl1j7wZO6qUkiWmzlVMW0faUzkstA7dM93pYUK4LyIbsACoVvKggWaNj68LHcdFQKdYpnR
MGDlThBfJLbUJYmmHeV9tWh1mX5dJBWJVlE/a1XfFh314kKH0SUQgmTgZIUMNBBsgbpwsPPZdnVp
iMNGrdS/iPDWwP4nmaxlsPR4Tk2NrmFe8V3ov+o68uh2DtiwWtwzzAfy+fy/2b3hNq3p3G7ZiKgD
1UldLa2TkiQ/KlsAvRXknKnultdir2f+v1kMEdHMPTxX4jV198UPDNmk8zQTIT40ibbMX+k+PmJ5
B7Fz+/QlkG+kS3DpsSZsK5LgIjcETtV6ZppPVug3E+mKCnKaj/CVAv32MgIyyxSlNBjW/uar/kR2
fUFgj7+wutWjSUOHlSDlBsq48V7ADn24kdJW/ei1gHWAlGyuMlEO2YiVcksHntap12vBwgWieDUN
jeiCHBEdFPwHqCcIwBybYWA+6uVIArc1Qh11TIjFuY1Q2tUfJ+tErDqeQErsqm2g53A4IsqcfpVm
4AKOduzJ87w6bvmgmmgeZ4WSyH7q+d9lHN21K/qOOUsefC84kuGS5Fh6TXMdNH11ntDqN4b3Q9OR
eGidMSQ8Mqr3V61HsOlIVjXLP3FOap/xYFKmOQLT8EF8RFoK8cckU29D+RETRo6IupUg8lFzQXT6
jpMZL1xUWVjj1yO1tCWts5nXs+uHjdmUlahRQmvm6djibU2UJZyOlQCE3LSpca7DUvH1+Ma0CzWN
TBmTiUVj8SvGVp5T2r44cKKZWGzA+cu52tVPwhdNJl9MXMrmrv8eAtxLiN0Xy81QvdF3e6+JiTfo
0O66WEcGFxf/6d0MjMPrk0oG+WyCJj56l46R3BkJMg+e80riJB7XaxLMn+O2B7LfzlSp2ZSEfCB4
8MDPeD3qcbgvbkuLp/THrdxYduSMrxNtW4U/NB4yw5yWeX6Q90GHGSomCRdSaILK+4rpFBg55w9l
6po/GMS71tRSaKP4VEwZo82AmTezIE3zEYrQ3kHrRyNYa87JT7lnZ30jOMJ5not8bcawPufKigH2
r5DK3Zs7KkDVT/zJNeSvbxU3eDAmvBCpgSYM4TNm3A28wBGnjEgKbNx93e3Yo98NCkxFP8FbxQbb
f4J9Voq5+SRCJbxV35a8lg6o7AhNukOgq4RkXLMLdxpdIs4OpcAkHyrSLHMqKtbLNctOCkszZiBN
4TWfsEv6G2G54JZnGXJlt9HvFHcRGJ119mKx1GHLHxnR78UbXa8pausgAJhuHdBMiC8htRsANuTc
Q0GBiUDgLaNnWqMvzLqW85BY4wZJb5KaH9z0fiGq9hd1Bpew1w/n8Apq/6fYJSkrXv7OmW35Bryc
gj9GMAOPvK0hZ4Ek9Qs5+WSwzJrFJlRfgxOOni7bqzK1B8X3/M1Gt9QiA57TRcQsipO8dZPfpywS
tNJ7InvFjx3EWVhrxU6FXw1cRH3ErAd0XbMNSQpioj/uYKXatq3BOGfqiVsJFBTtpDoPL8DZgs9L
IBLnuUgL3Yir9GakJlNzDVckEjfp6QNOeySNIa0rTT0yeaveu1NZYlgsvC45QPyIInbE0DEJXRqf
FlYiEHGz+0J2Ltuam8NjTQzQUFb7rbm9dRX5lfkwdZrerSqJUIancH2JZh56dXsdDXRyGjZuOr6U
LhTAUBBjQBHEHnT5TelXiEJ0ohR1sczdqRgwQJlAt0yA9CEGnL4lEyos6OoLmxj8qJUTH+Re2PQx
v/mZnBDdHOtPy4Zwg9U3BTBL61GYUu9aOnQmWQFSOMTMW83HB0zIeXkS23LwP9nxAcdLqJ+qAEUp
ANUupxnUY+CaGofPHiySesMAV5TpKHwJ8meGW+0GpHLZ8P5oT9rWimjyAHChLMhWpkwGME3Lf7kD
gx6uT3vMQgXv5PauEjgDDdFZ6cobMuOexDmQONJtaIRr3kA5wNFdyLiCPTKDADueDG60d8NV5odE
RwnVZGO3bKVFKZYn0oA2Bi3TUtwq/aCEnIh2V0rUT8WULTxLJXePE1ySs90lRGn2eQaQhhlxbuNW
eALxdzM8TO1oWOeqs7zoiYOBqz4ChQ8ToiwqgJCFPAx3aRQ4Vx1T/aoa5D7tpDLZYHc/cwYJPXR7
rvTQkkPF1m94CWBhCE29XvOYgkx9quBkxD4k72w87aCeOWHkkT5sH0MP6xZ5X3MgJ/L9d+w0p+Nx
Cxhx07ThFAiKveZuq9o80r1Wxb0SYfhTfCakTMoDGYN70jc5Au6uzYTJ18xhqLY73OmnxNHZgFbV
mCR59txPn2CTAOdN9r8pAz2Mwpx2J5snJfD/7IoISFn7L2udWTN+1holb93tmzOKkYm0CnbD1sAW
e9GN/r9ZpyuqHsNtof7qw9813d4qukMY2TY9ee/VWoIQi50aiYJKxxOECIrlBQwYTBl6gY5CVvJb
kBgKR5zzHo/mbk5Bs3aoWx5KtFWxCViy1JVkS5WIKbt76+Qn3qTRkidYeMfEiXCDjEcfvsMmqT21
3NTEy0WyPk8i/Ea50Rt4CEZpg4YHzdGFzq6I21gVCLtobYYteYW43ld/5/Z3vaB3TmBU6orFzfKD
G+enthO4dYiqzPc89+dmRznEMMkP0WD61r7TyShNa+PSUr5RbBEQ30szbtfyNxQfULYs3vZmG1+E
41q+dZFEroW7aofJebVdVaDdBGeReejH2JFE4X+KCUf7g99ZB+kzXIwIDgB1u010XJOy41CZ3sJ1
XmKUtz5K31VqnMTH/EpsIRl2CM/SbJZxmW8S9CepJp83CQQgUSgHJhO2DtXots9j+q0I8f6H2zB9
R5JmxqIIQiyudOR6qTYgK0jUV0CL3eXuY/4X5kxmBaIymVZqbBKeXMefvpf8kG+RtaP+DC1rdssG
G8Mr/JymtshLnhL6Effh2XosfZVLTQvpcIoIf4BDGj26cFxb3lw1JnpKbSfz2644pMn4oo5gv5+M
PNO+Hvd4QMi25BLYxURCSIAuEyHL9z9gma8KfB3D/U6N+ML1QI+E6pGZI8D2lIf8W25ci1pucv5P
9bRwA9JqOFhx92oTt4SR5Y0QVnM9cLkz8iR98EpOBpElzyJvQqbG9t2/2PO7i4osgTiLxYiqDBas
Iw2ZC/YqF4xqZGo+bGRnt0t6ot7dWhdBIECFn4gSc4gZEC1jR8SpIXOimHq0Yo60EPN5opIBrbjg
balqzwjxfehXONo2fxNWNNeMmFOLgDxeOi25CZnHqB3BAXK14gFTYOZK5tDGF5wxznhAnqkcLRyH
XHaNP+u3VTF4ED8mFYGWJVW97kedVWKuSHzIB9mnKsqg9x2Dg6jeKbiUZ0wFHsSCD0ZsJehFFVhd
Twaw6oSFV4hDBltXjanPvqKGa9jUaSmDc9lfW6gBPjqxGghCQJPL04OCmz/b+V1FQwmikn/m25x7
o3ka0Bk1WnEoUtwQAS54PwejQSBaRzkBbcFjh5oKpqOCXi0/A+s+37PfnhuZ09uR/Akmd4QT96DL
02VrFYrxHQIr4HotykgwnzN+groqYbaCCkHr9/IX1+eH+qy5Gu5wOHuAsSp7yvVlI6n9Q+fdvjmf
Tn1hRdWT7hMEJvsJoUHzfROdt5BEPSIhC8y7hogLJVNQV27ikSjleIOWQYsKf/dYBxe2+lRlLkSf
mitjuBxFt5hHJn28IUV+89rLg1XiF1AnZI7obnCnw2zT5ASteiuTju2EW3YnCzokTbpTnq5y5gCX
Sy7qIb29sF/d/WTYI9RDcV9NfEAE0tIEtzR0EnWHFipdyLXffbiupxDDhLGiryitvSaold7+ypxS
SYjRzOI05D6bJiibQt7AI6ji67YWnHotUZTXhvAKLq9j1/hBThBMOIuaVO25mSkdiaJbkrvupGGZ
YzO4y0XTT9yOWXita/+ukM+XdKoCXr113tkro5r41ExBkfvudOCstD4zbRAYc8LwLL28sjFgUV5R
ou3L5ZQ82yx7N6AUMPoWS2w8NW1r+3F4HUY6dYUjRmP/dtNAW/33GI+meEKCPWEdKqp3plA1brKZ
bhzpC+bzdSVXZ6qgFCvOTpPfPJesT3xm/s0NMK/QCJucRODlXOVkndVbIWQ7pti1q2LhblIiqY2y
CshQlQANv/zjW86d2iennZUK9up2r4oXoqM74AjD5+d1bRLGxB23fKfwPj5euiRuYOwovAiS5dR4
Tmv9AXHde40AAA98jgdpjaWqS2opeBp2UoIxGxK3X/haLZ7nSL3ZhfjhtLgqv5LVfUoaAy2MyEaU
XOiMXr+mC+NIgbLTGqnX3z/i7GUXFcj30OZwdY7CQ+Nr4g6gr2wTUKnGPTr58OXUEBLf9Fd1pohz
myB+XsopDi02j653DfI89s/lv2p2kruNS1BlYJZbuiJnX4qMqpdN3Q3vltcAKohI5zfJtVQ1QKlG
gUXWrMXnVZyUfvGt3HUBKhy58cCw2wdn6iwsXIzC+719yuRMhAAaRXwVKueX3vAKyD1d4HPmCdro
eDFLvF1JC/tnNaWSWnAntTbGSODQ5FX4/KgEQfH+gFzaN2UeCPskRBurSsd+J9HBY/I+AfIWk/jg
iNLZYHZBR6cAlkFSVB+gB5/KWMOSl7kElL+CiqN1GQYHtTLdonNYumgh2BAkgwD8ZKmCuhVpM0F9
w6votwA+tZtMRVcXU6BeAIboD2I7+0ei1on0gqlLLg1hZtG3kO9wZi8NdFhP2/H8J/lF5RCbhw1Y
o+2prClZp2YcvCwRYDU8l85VFwuAdYJ+Wvv8Zc5cOgiETFcPHDbMTlQodGouOL2X+9qfQd5h07AV
Ak1l9kA+BrLOcXDCIfDQt8JukiI4wntN9HsKm/JLCnnm5e5Yu6AhgpAWn1eB4qJtvO55o7ZTeVCO
zmLmdpWoHMZ/4cheK/2Yygr3gG/E1wYfNeZUb78YWo2VOZO76Yu5a3zDQ1t/D54ZctPeBpLXWOGZ
UyRH41Hu75Bsx6y0WKokDA0tQiy7jDa+Dri5bFZjfHaTYoBSoOXmWAY8tVkWKEX/opZhcaGgSGiN
8AUbGShi2kykE+Bl47jEWuFqW74EH+E8Ic8QjVa3mAn5AFigL+EnNERwcOIHIXI8pdROwKYy8vm8
9GYs/EL6CmPmRg+8kF7eOvuNC1QIJkQfWtBEkoVuFonQDlUqpYTzi2yuJMu45mJISX/U/GUl5hOG
zFCLUMT4OtUV0/2nD9Bya8vTRQWDvcaujprt2+nhhrFFN6aPAntfZFcVPYXIHet+vD2ROr6ATfEG
+2bvuxJPnNF2F1KX01q93Bm72+Vf8uWBvrRY5SyqwPa93BNhlIZl4yCxrUl/PWlGbiCbnl6fHXje
oQ7sMBW/5vmR9Ff1uvzIkPYv9ha3Dk/HqAzXosHb/rQ98OmUQ57W9wyRxm+81F5SyCUYTDxxu+0e
doG+b7gHhn+9/GjFMOHRMAVJfJ/7OTToQqaFda2X8vLd+W5SZFP1thaTTM1d5OS/+Q9yCRAb4GhH
Vg4lJzK2VCpKmIlVvjK5tstAskF2DHyIre/yOhzqfQ1EsbCpHMi0YnoNneUZ8AskzsAog9ydRtys
4b976+1YwBvudKAfZ90/8PxsLcT74XirkeLbSMOKNB5bD335MMjex2qocxoEPk9mJuDLSqu9gzav
wOfxhJEmZcmF9/LBeuf4RBbV52ICV+/D7fJQdlvLGfFRCZqwgioqNrZx5Nb26hsVTCRfjH0hl5yj
de6wFeBqiOUx/ZeZWVuUjG/PD3aOu9qLaJBk9w/xrMPLHtCNGohE7LXRssynCJUuZ7OsqLD25uaa
e7CVXw64ps0OTh076bQK4bOIL1rMQMNM7nDKQ8ffZatqvHhxchcAjMoRL/nMioTedWx3n0fhZD+z
5AU+7kbztPJJbiHy56BHDaKeArNAuR7IPfWaILxgZS7yhZ0MSEohiT4wvLfRItxBjZ7kmQaEp2UN
vgUGUyumR5NO1Z5+DOkXd9rlwYd4nV8znOGf/saG0gjwwJ47UrO9uI1UNVLV9I2WkYT0bT1Wjp+O
wwFTSDzAXPQMFLyNpkdLg1KfRztNrR7JGOOFwCuE9OwVtGov4TIfpYZ0SwHekVWmJ9kXrfVPxwMZ
73C3U/W7vv5wAbZAb/jZ+bh53boJHepXVtRW6w2C2sLF0XA2CosC5/BWJTmLXOL5ek+cMTkGj40K
BQ9cI76QTR8EBYV23rrrOeXrbz685Imefj6WMGjmDej5ygmHI+zzeacMf7ucRE/g+a7RAMrXLLrB
1D9cqGA9mY4FnCgXUSCW5YTbXVwFa9QyQ1j1OXaI1PE3g2T4hIlgoXwxLT9Vp9iTLii6MTllo0tJ
ZdocXF1aaO7g32WTcuWODaUqKqj6pktkCD8MjHYshwBg4VTJJ9Bn60tmmfbT1WXzoLN5h2Qi4A0C
3XCScAiV0ejJGy/jtoIJPw9Lhin6dnj6JaUMOYYW6Q6oJdqOD2fYKJb4qCwoCid5+nj4Qzgvu+SV
1VOVOhEv1InU3c/4z5lEjHz12akvSsURbLhAQvMkLwtOtCbmIqo772lXFyk8UPTv3mDPuee9iY4d
CtjrSBXJxi5wIecRpUV9AHaa2dgYyrmKQGBx+BGrJ9Tv7iI+4GMPs5no9BmBfweUlcrKdBjjWusD
VZfJlnEFs9SvS5h4X2Wjw+PoqokQlGPfVHYYmFAyIx2K2GaN4PTw+4Y0XwZyH93hKeikpIqdA16M
23QEXiuSFHqdOFxJ82Jks2pZqxNqw1tvtMNRkTtWhWeMX6d6KGX3gk26JuhcITvSyQt+DbkBTHMa
7BOalR92kwuHt1Jw2moEJXrtyvm6SwI0VUBBipVePXxy8PXXdQiNOqAOZt8dsbWu181OgqEkrb3v
J3jsMMlE2SbExxEGxZ/+nR3Wf1ZmQDuxi3zo3Oe1lEWx0QBf2pjdRHGTB134Tu2t7wqHXB+zOU9G
MwlAUyVcJVNCFBGwZO8pECOPfq2Vj+wfydIO+yItiqF59lPE/32QH2LcKDhKxcaEeoUSuu9+jHhW
SDj0BijLjODRCmPx693/KMFq6+B8NPEZBcY9GCwdyRNwxvqDY0Cit543UzC3K2DweSdMi6V6E2Mr
3yLRfTqPLPqWNYOTq1G5V1s8h95MfqJuoFGsUQ87Bnkx5sMtMi2jVB67d3zUChtvzBLK4QuD4fCp
Od0tJih11MekOmDrIEDcojhtfk5F4cyzLt9EfyIZ5/PSwEJrRoKXbQyJ83M9meBEXk2NH8mAV/dc
dKrwRvGipuC08EEzh7nDFxDrGgFUpPwJOiyN8cOry1u9edlm8RTMeyO/gHHPC0PzY2erWY+F3sD0
2Mayfp0ETcjNX+ey4U7l/xJa+vt1dApu7O4A3wv7CA2ZheTY/UnVrMod0wBAk31+LGKimIeCs2A8
vN60647DY5dquElAiS/bD2fYDS41Xger1YIlQNe6BZcMFFAchjAHtFd+2WdK9IUrks8tPmcIalM0
K9xOm1N0MsrsDY3JO8QbblyQhs/TjuNEJCKFyAQbE7b+Luj3Agi50wvm5JJXJ0RUb3qwuNxwe1Mi
CNzjnKltcVx3//W7DJehg32iJuGK7cwrnT4VPN/xm7MvJ7nIyBIhokDt74My0RDaqVOWy3KQZI7A
Ibz63wnn4VpRzCQX/tT3bxV/KBijJqYEu9CiFZKdoCB5E9gr/g+5i998Fep7uq2CGMVlqZYnWvLR
2Zw+k8wLTUnSyUmqNr9NcMbuSY5RX2UM3zKFfP6i4zxygLW417zGETd1Xr8ljVfXhZFQ8QQ7vtYa
/uqmJIdXku59xVT6POwiWed3xl4dxIxwEmuf4+ycfXet6pp7tw4zV4nZaJumhls6hn0AxthRXwRD
fOUv+Pgha/nLwDt2PfMfEWK4RsOoaWvsG97hTsYMvmIsshUgjvFHaI7tPYSAj52d4tF1SVGW5Wje
hwLyXZJew4efeTExBz4OqCi2yn9fmab06k0juLknHuXTUZk4sQJs5B3u1CMPKV5dySZhz7J7wP4b
F0JNen/nnOHRzWgaaUS5Bky0WfvcQ6CAOzy0fjJ8rFbL09Qbc13kh2b0bHMpEYZr2cTd3cgJjC4d
iqbqowta5tdKfyCZXDvmuoRI7VzUICDnzJzShsbGlYkh7R9ECkM16sAKRfctUTW8BfaFtF/8yKkQ
iosvru6EdylR4gQTnDct4WhMz3Ut39Pz7+8xg6aFGsBprplof28j0rnbcvBkl4TNgJxjdGOoezmj
FscRqsA7ZLrDsRunb+B5u14+68pqkOgPp/vPFWI8YFD81LhGarCnulLBxY+dayvJR2nNzBgwwly+
L/ism90MB/BOkuO++qPsPvR2axW3onuedre3b1LqrifpByZkgBccUn1rvCCd52VmL/f0l4AZVjYb
YUGkZsjDKw/zRLKnRDabcI+vVGk7IpxeJcmuABvwlwJNt4iimZkHIf1y4ue4s7pTRPpZqcvexLi5
AZpttx4VoG4fKT2Kdzt9NElb3/szE3l0h8FKnGSywP/xGO2EfCH4cuAQeA8+nwbqg+Ct/EBEudrY
DbM5AXXvuM8hpmRELIFYrjfeHwBShqKmSAlWSl+s/y9gEB80H43zK+0QwvMEIVaJ7e93Ug8wc7Ju
DhQ9Q5OINLUQm77GIK5kFkw5qTZC1xEiiaLc4j5jjuU0LfLHDUd4SADdkkFWfEj/59het+k0nMkb
L3ejE+tEtAzNL/+r9O6w+M9kNpGMM6E9w5oGjRCkBzJdEyVZaLVWp+5HIPtW+XWy95y1J7fhxX76
mgBdxyZW/VfGjkmjIr+StL1b1VR5AQ3zJwXoalIotsJ5apx3sUdy4JWpsxOcNQodrknHv50Gp2Ts
e9MDBn/neJymNi8GdunjXjp85kQ12Q+6Egu9durzTeepwr11jYHip3huAqGCY26CPKf3gJcPwPrj
rovjZ/vlpGvpJKouIIGrY973y47M7bzUBFSzZa5QSAVAn5Xz56LQ2DxFnJF12yrT5l6JQgIcnhJo
N46Eh3eOKBsGWm9uDnkCIEu6JM3d4xV5+Mjxbp6P/DlPy+yJ+eoOuBlFvj9ejsrQPZUxQI/iY6cC
M46z0ETu1mMDT6lewDzfEl3hMBLlCQ2+1k+mS3AjNEuhyk7yMlY5gqjJyJkUlYoyZWe8YBm3Y9bB
pDb9CnYhpWCSjpPESvk1u/ukk7NGOi+feOU5RvdKl1jLdle/wBnRQb7IY6WY+S3IxG3a9Uy9+GOH
rHaoqlMBFYPDtw3M9iTqJRJpeW152NaTrsD8maDJ+rFaoXTpGlmzY8FW1SO4PL4H6RoW4mLOJiCw
v375cH08lRZKoL1Qa+S4eq0lgdSx3Rddts05i/5HdWAWFkVlh6yJLNMvOZtrxUvHsZgyrnFQRJ2f
cjZjEqcmZBh6P/DvW7ioVkNhgQ5Y7MMveQ/3zxfFR3qxwmFdy/25+Ni8AkUEJNEbppsIA187qJ79
m7M7QWXbuV45+UZ00aBx5sK5n7zd5xFkuSxG68Xl7ax5IzmFDjeZ1NdTB3wsN9N4LY4lGkQyJE1H
WP4UwHgnlp8KQ6rcy8eoJVLtlX376eATyEPTb5bD1xZRxFozG3uFf8X/rNt4+AcCZazFdSdXS5ua
9MJPC6AIpl1/QSzqv91Gf7GfCwFmseJkA7QyUGsI8Ty+ytHjf5EJS2H3aGR2nt3Tny2+UEo0HuLz
JaRKxKURYa0RNc+ayoNBz7uOZYq2XKKYSGXeRjlM03ZBuumKdy8QMAgy7PiKkN8PQZ76flwRzZv+
018demajDf+ThaxpcA5FwHbk0QNFC+Ko2Z/tnhh5Z818Mo6cSCGi8nSalVYSi7u/BqKiIuFidHpC
SHaWA2Qgw+xztvnwXBnX6UB2haOW127SknOOstoHugVKNkpqZdJcawh24tLIvtOJIOTGlU3QMEmA
xZqU5Jm525QagUdSJYW+f6n370/GEB00ydfivFI5ygC6ogYtuWvqIcpEszs9ah/4ZxcOySn7VMjB
IS1KjAtX+FwA8vD8AuOXXaG47KObCg00wNbCnYcSS+ri1INf4vnGbgO+yNW0mlAplr3zWZ9YUaaU
NLeXyWX7CjlATKdY/PRIV56Bn7qXUmwtrN8gn5zHzvdzGyWqdG8vB6MpZ9vuwEM6IRBAkgGI/+qZ
aCS+UFRDsNrGfNK/sCQcV6gjWFCCoMVzYp3qVMhQuZbEfz02G7R1wgNYqpUhi1pAm8tsKMcvI3ch
jdDbyn9xFb813x9c5BcphxWEGxXtnndedrurujJJRdMvTWEDWBBe+8+05iKwSCyMU69MyH3HjRK/
nnu3a7yTcmZTc8AJ71E8HMwKyDdpPSI+T+++o13AGUDS4CZq6cUaOTMPMxEpfLK+MIR5cg5+29Fc
CEa0pDoVbfn5f+Ieeis2zFs5yoAbv0f/Lix8sN9yFXOentzrn9JVDsV+C4V1HVdVlJFfplnVsaXo
+YSDFzfZLR74L4mQZRS4rDylmyEHp6ltTGEzctnkNZVb3JsgpBUxmOTeSQMUMbZMJP42LbWHhF4Q
Z9gPF33HJCauQEwDjzYaTBHwvx+XNMH77qNjcmSG3gwthNyGgFuoqAPbIHbDSeO1/7exP7k1Sny6
8evESFV0+nD+/fLKg1BwuabNV8r8D0x+w73usJwZrQ/owvZPV9e23PzLJCGVwpJ2TVkJCbb6wzSV
+2HDCGa1+1ewjzQHiJq8dedzty+1znvJS/88LfmmtemVkZThL+lhvFSYTm02XmBzYT7JrqJikKSi
QafWngbb5cEiGt5ViSQ1xInQs1upEjmQKNLvmptKW0vzlJCiLYZHjrBEUwq/TcbTDSK4vYcBDcYH
GPkbpmI/JJU5gnzmb20u+xcIxm4YE7Fs6CM1VT3+S3B83oQKZBN+O0NMdFTdCSW7j05WHYYSN5td
ITg7ZER9CHU0kGUlWJxa6nijcRyQtenHgaP/xLagoAxo4WXR5l1/E1Nrvz/oFM7YBmGsFJWYOa51
g1qK2ADaEYP8JW0Ohq2KFH4uD+CxRmMfZZyyT+0F1COLoAvkOdEZFWD8m3OuZ/gZEPRP0JZhi/Rs
6XH4hG/LTeGoBtFdux282kt9dEmp7kT2DOXkI9tAnS8/TpVy2Ef/S+NmZVz2u6rD78hOjO0ZJ36Y
jDD3eg088d5/j82qlkR61BMIe+uCCgtVG+NAZW4gS0D45AdbRqwCoFNmmnfEEh29f0GVrlTbMCwp
XVxFU5EA1RZFczN8n4aB5/PRRcnOkSqFXap9p2DTTk8EO5wz2wxfXn2jF1ue6eb8ZaLvnsBn4kI/
BXto/Rfch7uf3LjysIaQDMFR0J1oQMrjR0Y57/A0jjHZAliN9EXesTKjjpHmG7U8CIAnicTidz55
Mq3/rGzT07ORbSv9uFoIpbCE/zKAbF7YqKRvMyIsBfPTKRoVqa80+CQT4dgOLjRUhzKSExzTKjdq
iathiFM62Q6lb3T5PUhBlO+Zl+Se99lXnfPZJjiABI+AK86G+gFpOUYO8RGUiZAerTnBzIytkiHL
6kJCtb4q46aA3Wxuz1JPqzq2J9ryZI4oDw1zk1mc2Q2LhS5RunpH+KS6mpA/9mpnNvWiKTTP+Qan
aAKudIwYTdn/+Ei6tjbRRU+yYg4dfPK6keQA+TmUosy6nVYhNoLhA/E6IAsccjXQmPTk8Ju9/ixP
IRWWmpH5l2Kx+Firk/x0UQbYTbW0Aa6zU2fr7RoTgeTkcoyrbz+uzb7hIYCuj7f2IpG8SRdL8pOV
IworUdjvUY57rqpxeugibetvq7PonkNmR/vt545K/3DrYdT0XJPfPNa0EbjdF/QPDh9fyNi0GIBh
0gJLcpdEaCQj8Twxc4Kr62dOHxsI538+UZZfxi5Y47nCn4+Cz8i9ikfawM/OgzFqtJRoCRZbUqHu
YxRxlDz9z/c3oNofuD8aX5/3fv4kjZNogfxWVDCq7FDBaM11fN0P9kcqoVJxiAj9Dp+9vQrdATFh
6LnJ2SyWkjCqpU/tIXmEGVcTyPyRnrvXnDTKiRFYDxgYV9KlQ4gI3GOxvQce+/x8yq/iU8NOOz8w
HyB3MrNtZ349dLgaVU0VsUykVqGFZUnTt0gkDSJKsxQ81xOOif8bC6QVsN+5G9oGZ2Ikpj62iaFe
pUYpLWAEdJS54US8khIVmUSFvZuuxhg0SKehSOwt34rbsAcLIDdcyumrRRFjmz7uOoCiYcf3U9YO
RqYkT9mEeVnAAt9oGW0RahIs5UFPygHLlMX/DZCcaJxSdiWQ3ZYB5iM02jRd3oCnlt7BCaCI8lMQ
IE0+MUSXAC9gU7MM41x0R3X9j4kvNoKkP7nP9kAL9rHCeFBaSQStZW8XP6Z8KMDThoVfLvMRPxzX
G2kvSMOCnn80g94drqvYvfjl9NNzHo9dG5alpfMRMsnrQpPY3eP0YtAgwp0rRi/bY3WVGPUJ7oRt
ctlGL9qkaTY1roCTO6/BaThu7gE56zNhzzmaGt4mlK5TVlnhYX5L07o8W6OZP++YM3LjXlFFmCHJ
JU/d4DLueEJvQRSWFnAl2bZeS3mjJTQacH267Iq14RK9UXXJug4uvHpYjqakUVLFcfd+VICXCjdp
k2oiZrxHZUJ2Lq+6raoYcYiSpj/ZfcsSXXDvTPhAvB26N34L8O/zxUqNG/48Tugh/LnAPOVVwiq7
XiAXtsTiw8tIcAfKOMivv0TLfmkoYc+qNKIgpkKLH8zDcSIExcO24d/qeGOLLFIop2bmeVm/ekgk
ide9zQjik9CtTcDoHI1LzKVWzBZb1klXglamRd8kr98PINuYvA6cghl8PHbZX8laXdGju8nthv9q
0Dyo7J2n1uZ66A7UikjxM9n/mrE82NdVs/+FrdrzgqkaAH6SFcI+bICJhcpyf9tY3jmqK3iX4R7c
Ib4c3/uN/XUAQ1usgUF882Md/YXyROja5Z7bXVW411UB2HwNx/YwMCTIbSffJSEUUaQR52rSaK2i
GHuuV4rpC880SYwC/8NfF86iyWXRuckTqeseW+87pC/VlAV156Hx6XcXvuVRm1j5RpzIpfYSjQSZ
v5TRj+mkTUsRuAfxy5anDDkpOly3WkyReH7iRK/zu1A1rYRoCN7bI3VU0lSgJAfgL8aJsS7HdnXI
A4KoQ6XtuKfz75B4EtcuLBdqPYinkeeoUHIYVyMGUhlqb3NBZjgPXolJEOVqSS9V+51BpBbE8zr6
fMoldhTjnyIwtkOoyGuINkX5N4H79SEpTPgOILLHW388do63aAqQp6Td2O0TvOWX6mHzmLM250//
fWz3V6AeZAx2N8Yk5PWLw2TPQoK9KywiA+6BQlSktSiAU8vJT+l/YxitqdLZCtozBb86Kv1O63rQ
eqT13HSdCeBfhitB4i5VyzrumEdMSHfCsVkaYkA3IXY4ZvA2G+gzessUIWAiApyZI06oPBy0aFax
WOk6J2WyzOvpCaHvB3lgFllkGEhDrMQ3z/St17QJrsFD5ayc1SCiG4t4/NNxQhkDXuaCDogky7dM
hUhn2XRQOCVbV8JFq2XfhVako7D8rKcmqN5Rtx3o4T4E/8FkyZkfChpWjotitcgdfEil7aRMaVfY
GIwntB00SYl+1yeGPih59npS1ykkuJOydCr6Gl2S/CjU79oosHJ2D/JaIZngtJGIh9j3PrlSThan
wNZ8FBAjYZgnhSoPo+tu52o3SSDS9VkE6jhFP6NGBe4Leujv29h9dcShr+tFRN93INWGH4YeuN2l
EBR7jNcLmTppcI1s0t6BYuTSxRvAtFgd7tFCG/AuA2yA0bXhBRy88SQyF2aGqFmA27L+2744QnNv
y31hOQc/TZkA70CqPSyxFz+GrvuzCMdpy3DrRnm3tPRTJn1d0HiClTaPnCMm+HlF+e7Y+0e+tGeS
I+o74HiIPLqhtx4vI5vwIhrds9njelCoGVSp1D1zX1ge3mDwM5ciLNJaXv1XpyeZP0G5HT64U1k8
WTeJmDxSE+yKBb0Ozp9fN12GEmtd0Idv8UwBisMx874Yv4T43BFk2StO8PK548izvbIzrZq6lQNV
lJg+5GIYUmVcR9uwX8QHyUF95pVL4YCoLqVRKfy5PKU7djunosfHTpkxr8caUdt3Z+m8O85hLbuk
QRw3PIWFP7goNXx6WnXIXoB4JBqL2+H2bJo03WMosxtJazzG3K8UtMnPQjFnaRX/4CY/dFZL5bz+
HgSMhHRJE6ZkDT+F0xdY0wRr27sRae/2VioANe08rrNVd5VY+D/735XHNAIYlaTMWkTMHTzj6L5u
Z4J7q20+XE3Bwj4e8DbITIv9YufkNA1vkCoy8lZU8HddjJP5ca2G3f3JPJiCVlVcrFikZ9bQfIHt
OzL8ZgDSdj7TdjdudZJgboiXvH9GE93xEoddu4cPU7DgryUlnjkViLPjNK5mDq9lpaPGhHX9RAP0
0UIkZWRz9SxVArYSNZ/ADohGKrvSURRAdc12egXcB+WAP5b/bIRX7FPXYGzYzJ9mgCGRo4TwWGOO
9KjG2O4dGcoBYmHKvcRmZ4Xj/Wu9R7GnOtEG/0b++Cv+8O/2kU/3XHBH6XWhfRPTox9WpnaOCp8a
EIo5PrVgl/A8yDT0WKHR7ErRJ3F2l/XAv1oWyBa+bilRnA/KDhY8/HRLk1xf5qRe440iRrt950YY
ExyDSBc+NjdCRJxdmCuLFMXwzjpdc1LIv29bZhc8Fr0R/eYhSjSIX70kGgy6Gl6tgrfhLRhsCyvy
TCci5wU9Q/2iTnqa+2rs/lnfWYhEupURjaN9D5Xz/RH1Z8iRZFw7osBOCzmhA76J/CBTx5o5ndoS
CMYTvMzwtekPUXeEF5V/ZuI1Fbx7uCH02oW4xNgJDFcHxFDiHm8uSskzLz8gqanQN81R8mH5Hwnz
0KdjsbBlfYTFLpS2zgbm24QyTqxMSIbnjofCiy3fdECDZtVknqQNkDcH+02VWOrkcin02Oi+quG8
hly4+Mifo2at2Db8uKvmaLCjOO5GBk0mIOYad+KPqkoLPYbct8N5Jf6VD4qnmGF+hS8UbqFLtejO
twt1Cbdk9IqJxNdBMDr6gIHBRLbpSFyDhHrLJ1FmOI6PfxUJBbuRZZBBihww4mQdWzGdj11Ty5qC
tOXGc/sF1ufcy0UjWffzRKT3IJ9Qrp2bmilZsRNZFrHkSXBjmQH2/+jnH1WG6e//1nroypWzFPRQ
dQYSrxIks7vtZJ3GmGgAWeUo7LWjBZw2Qls1mXd1e7/l/GtOsSLlFPuyiSMsu5dYlgOW4bbGucOV
yZRhs+f5OVC6eNWw70Dr/6qm5q5IPxjVCCPJvb1APdt30S37FqEkU4cz2B+brn0CT9HnEgTq3398
BKrJslAbSTCVzvdmUMPe4/O6ioNqwuabFXSaXuq9NZsTJ/oAOUrqIGAYR+qYAJVKXWb5r0JLA9YE
jQARreQvRQwDej3evwX5YUFB8bVKgpALZ6nwuZmiyr5LQYFGozmLXDhq69XwRldcaXTPHd9SLM08
Da59ls+rnnHDQBxMTnKmjX5ne2yPk+ryFqJZV1nzMNMzyrFEEaHrGTdzCDPhyouZ7KvJEe0cDx7W
rBuClNRJSGEyc7NoHsGwotrulFsCmkt3j10ftBCqrepDxdMsqwibitxcPME2yerhl4lVKpDMrSN8
C3cnlY6PymypedzzuJgnuiz7wtXj7KbbOreUSBCul4UpLWnPfuN4yIlgdLp4iHVELCfJlqxK75VK
D1SfWuoa9jEkXI+1Q5tik+W6/d2pR0CRccFsKX0CtLc+Mm3+6oX50Mfv4kGw5fQga508XM1yqIEq
iZr8te1Wd4vgCfpFjXCpyRTcEVjtcHfg+1411yIR/oWkap+6WViMI/RlAvF2ewVQgxXMh6cD0C8p
iUVC8qkjgWfVgIxVjz/wKBGom7PwVoU4iTBKkfA5ZmMEau6BgE8B+xrnJDy8AYV6cudH9OR1Av8m
PqsQYvn2gLyPaKZYTq/mAlGFcu8Ad6m++trP/KfRCKF385zEboLRO8u5S2nConyn+6q/8QwzJJFM
zDTWBY/J4keDoNam3ZbLG6FfUQ4eaniRcXjfxDHDE3x/5YZ1YHsQoKB/6fDYP1oJXbb9rIS02kZ5
2K3KQ32BRyAWHv1MMLzjT5IMZxkRucn/aD9r4lLUGMFg1zte6CzC70ur20Nx9jpFF/wtyr24uXvd
s7QqLE4TgLv564lm6KdNhSumyjzIzBAN9BgOAJKI2w/vamd35JrG9F6PWKe9SbhMHay9yBFPGWOI
aEsEsWAJ1S4p9u8Qbnrv4EpGAmzDmNTiyTHVofXKUx4puVdT31aMHqsw5fQR09/z9rjXkP6+uYKy
GMuqRfnlmFUz6MWxTI4gxmui4Wkl5sOm/TW1SYZEW+gYE2vlJ9I7nNOpifYjuBchngvFW6Dy8CtY
84iuhPBw/Jw8TYc6lUuuMZ4jrUDNnuEdCI4ixZcEP3d/nzsQYs2Z44H2TiatfvcXWr4IHRGdnt55
2g31KEWYmdXZSQZdKUr5eq1lHVYa7bT/GfFaSrmc3OR0Rgl9R/zynRaq3YpsZqe4Ce+Zv52jfh6l
WVLMB2BgfQLJaDF18OrJW2I9+qjPsNJdQbgMunzLW+jZ4/j4GhhPMH2FW9CDP3RLJfOMaI5xZ79U
hW0x5LkbgGKrSifv8nmiqlOLlqqMHOoWhll/RW4W7/+m6UCOUZIG3BTwgNKe27VFFrVbanJwk7k+
1DFdVIXHaT7WtBzRWuSfeDbN44qET55sufRVYdmB/dJh+wfPn5uK/Of00axRKTpug0gtleM/RmOs
MtC6PF08LOrfLVYmvIcy5AazUfzXi8qwEy182qpkHdscRx2qaynv24uWbYOxWWbbxjoQ01cFa2M8
A58wD4AbXpwTn/mObrTKfHwxk9xCpcFwjUMu4fT0/1KkWmC1rxm4kyEK+5C0CJFAT9vEnmUl4wuZ
o+gvr69GFdpf9wUJyaTbQpBiQllNcmCP0d7vwaVXuupSnUfOfd21XUd6FcGTlujl31gKY1aLdijE
HEEExHLYUUiRktaR8bDw6JLg3d/rVUfD/iFcIC68kaCEBdDwsSjd06XZIYCV/h0IUDNojNv5uRo1
5esAG/rHIOijxJNi4h7kn3OZICFYPNQyp2DmG76xMUuhlbBerUdn4yWddn8aXe6reKKCaFL5rIfh
04YetgB3txnJvjHRaxMuh4/na0M3F+UJhnI8PlOkc40s/x71wd5/sy3sO0zedmWn9fjMxNXO/WVu
QdCD8H5I1+ttuGk6VGggtRBLvMR0dVHZKlAMt+aymgzj6L00q0YhzkhP3ymky7YModPF5b0bPzRE
Qgydc7evDuTlBMCztIl138VZheHvBoL5QFCxJ8GOKMn0ol1fhdCHQMTsSqFJ7GQFZVSzh3N/zPp5
0FtMxCbpw4dqILKW9K6glfWFaEOb/dm1s2E72NS/fCFIACE+3IhrTJyuKmk8Rf9FxDPpNsi5DZAw
o1sHYIqXKpzlDa2C2m95sdDfSeo5TTmaM7u1Y19zogLP1KtToCg7S2ju53BWw8Qi3rptS4phk5ks
zvK8Zo/2bczpsdZHFidRboSifDPG7eooEoV9Zes2f/8bDUHc8PVZEOxvWRK4rgj7FivRyM6+quUS
eH5qFOBUKJCVN8GEiXIDGd7J1PCRlx52fSLB979t/WqeHagCNTyq4Rmc++kseKSm8IFknh1T6Io+
wdGdN/I2Dv+7VCrouDTw4/s/gL2uC5wNuX45nE4YkIQJSnpGsv7JhA24M/LIRUYj/3EWTnlAOybY
jl+c/jhJhU50OhdIeqmi9jQc62CULQroto8tw1JPo+fn2xiIFEl++REoedhpz78w1N4HPLoArMi/
v22UA88WXas/rMbRmGV2gIc5Vwe7+XEwKgRjdx/zCdsuz5n2nWvt1J7oqY0e5C4E07bdnSReVqFA
xRHYyVKZXkU3kLXQYNC9qnaf6L0eNpYquEIgcOM2cUSKPvj+sR3LVPQZvT0gNTxsl6OndTbEts/i
XJ0dYj6mLZ95kWaKOYLbxBduBiI15cQoqhlXh1wfUCAsofwWgv1+Pqc687Hzb2CtFt1xba6QYokP
Rq0eCoqr9QrgVdnlN50y5LWwYU0fbLDLJssVGgDebG2Dwa49OPlB7/6en836uKki9OmbYQHBhtFw
Tpa6ExXxzYcSIv121A9G5/ri1l85/v5xmQ3f5/9IxoITkyVbG4LGUW2gAa4oNG6ONYHR4PN+eHZR
Hvr1kPgUxfWzFXN3/Nkq3JW5STvqkIQhvGLvcxs2Df9yL1dMHKKvwJRtquiyl5yFtxrEARomXkP4
Yf4vRTH7j1Z3uh3A2Ldc3Cywa+vdh/EPsMwDdS//of7tTnoi7XplXENVMK/EzrOELd1gfCVVQGnX
qSQ6K8NiL6PoZc8VO3n8hrbS5YUIOq9NC1Ipis95oDoa3vicBN8Ar2riMoSSZJbaTKmavvQSZh2q
4pNL0L65ucm7oFBhFKiLprazS7N/aIfInSNNv5/m5Oy6NHiXzIYwXLPj9Vl4fl/GIiCbg2ImCsTc
t6wQv2aaJm/XoImqUo7uBNwyr+hPxdi9HVBJ008jwI4XiSR2xrBfwSoyRSNpMXeQLDa8hs0aqU7I
Smsk/r3MnQF6YkOvC4u2V6X/zfVmD//7HyigskOHt39FFW0guZXEbZyZjg1G0C2TJwJ1RTZjsqNk
vYLL8CVBSH0WILbtqWRIXQHYRvUm97Mm+utxXv+dgA3H10UOyDDow0cqk1GHp7QJKeSM1UrFlMdR
PfJYPJYn01sh0TS4dhVZTgaSEA8lfvLeLYXHjVDBEx/BOcaw0ufe7tHmW3Lp8syNSay39gHfGPgH
KDPgzOICNjgOg5YqRAsM4xfwr/lz92TAj+FqFv+beg+vqiK4MOH1ilqg02GpHnF76jyKD/sxSMdc
NQEpRnqNvZuux/BO8ibfR+bZVxiQDK06Y1O4SMwdHXab7CbonzqMvD1fESVah8CQlhPlM3eOZCls
/mwzpt1HsFxf4F52i1AINVM7jraIRCRmenw2fDCIloFZRS0IhBou/Tja9mTWlf68j/rKShkMrLRi
dYVrt4DDHaVoAmFS52C11NHGvMEDtiZVtBZqtOma+o1dA97TEib5NdgJp70U0Mc0Q3jPae8A7hcj
Kjc0+wL+V8cy5ZMZYEQ+S2cCH3y+KXn0kKmZd/fnijR3XFCb7YdoRBWEY494a/KP0013p9vF2m3a
zhGlX6RwwqUro+d5PrHZpCibx3p7mX8SyuRWnjCNqfuCOtP5WwCpV4QwRR9vJN/y9BngkUJ5j+Wd
qOYckYZe850eVVGqojn939RX2QwaXED9pgc5lsJzsWhRbPe012OszMCAx/1BGRvDKNCAaIJnE1Gb
AZNGGGPujYaE3oi4etqYWZS2esoHV2baIN+/wGeJFX8Jxg+m6JXEvQPJoM1SfzOOYV6P+TDD/6xb
scP3y1R0Yb8q22SElBVIpkNm370fIPnW93kLuyrh+uwl4FbkQMdwQ5o/04Ekn6G1NGqFO7eEGRYD
9Z3nK8UV5AYf69s5XEHTaVe/dm+cO3bPx+g/WDs0VU/t0OIsmefQX0ACJNwrRBgncMPiEkiWqck6
pmx9F609fQF14nRGhJfZZBDEHY/EkpFSx3vwxDNkpExGQsfhwMJnIv2s9cP/n7mpyY0YwLq4xcHV
1SWIugKUMySISamWjaKvadDL1Skv51pTj/stYZbGWEWmxnW9YbbO3WDhMYQNgKXfuB460XaoqIdK
oaDa7XZS1QVg+XFHeVKYjsDjoe+GDzxd9rnEjzC1TBeOPb+h1XOPhl8s+ULgRZdhxqTOkbvwdPYb
SRwa7SxFjhJov0fWZUo8Oei9oDZX2MzOiHcoyhGegcyzBKBMeMq9gCL/3S9ki1ea+okKyeezU27r
8FnGxcajMAZ4wy9opNoXjVtVhLaxl0xWP2mjBmfD8sqGWm+AbfXsIs5DftI7Atxq62qwk0xKiZQu
FdWIqkCOL5jw4eY9DI1eMqaxBuK0boLoS/kNhXtaBeBgEFhpqk9dj9omDWynnji/sgkkD0A34dxv
++6jUZHbLR3iRVDDggLO2BHxO+l45x+Oy6BnarQP1TwKm87SEFRRPRPvLShmasR4CfnVUi/UhpqO
idSCwVDfDfNOFEJk11/ijAlT4QSso6r6+JctMU2G5we0k0ILwrFHLzfBEwJmxN4jcjltSeEGgdOc
9RMXNUZWBFRcCJtqpzMbc2wIXax7oSPu0rRkAa8WPitHRb0wmie7j7UOeBYbuZ1nYfZrlTtiTsyt
BsiFROtSFOAA6/x70Kk7L0PFpwnSXLFVlC43RCRHxJbJkFOihQZKgivx/TtUIu7NDBLw2vqtIms2
C4oNREmpsOoA7NqXVJ/RGJcDf3UhIAa2rcEnWuRhXo+GmSRxYtLaoBhXNK6491g7rrvx0vDz35zo
pD6PY5VrlJNLEs3eOtXiiBUwykFkfZRkw1LTAlVmuvP+vJ7W7PCsNkZU72USQAY9OEZ5NqoJQqWr
pWWBOFTsRI1V1JNGJaBrydzo8usrwK8NxXN+TlWXxZUuDSj2GZncF5pAyoDsZwc7+gjsCogHaXSp
WbWJYWGFRC0wBdnrD+Xow0NQWpvu9uilvTr1t6UxRSr9LXqpeSIu6zFSI+x6VVLEzHX2bS9OApeX
UL6Wcv2S6Bk5zcwvt4mWVmZodwIsuz0f0l1gVEjt5Q/CpS4x/ZNoj7W8Qy3YMsMxQ6+jY+BZJnL4
KnKLOmD527hrKeL4Gy1Ks0ZbZnpC5WIvuT7M9wmsEpmr++N0DUaoV5B1K6Q0bJrp9qUjHAFNaTyC
C/unFrLPAuqlL3g3LHzAkU7D728qs04VNR/GMKwQdtSONPA5+fVT94lHxALSN7uiHN172KGgs+LP
RoY+IDU6v5A/jTY9/xG4UyjFU5nBpYhbtebX1fQRvlmH1HIff1x8XvOthdhk8H19+VMhnt6F1l8W
Y2p3a+Z0C37qPhwZQ7TyR4fSjl9sE+fAeYeq3pf35l62d+z8/YivX8TplWmrD9IogrcMGZl3ZyEw
hQ0J6XKe+mCF1u6MWTVp1JOiiz0oNe7JFzCD93REM5F6NFJwLhWU3OaVTxtF+NUiN6fNUhpIkBR0
8tn7z+6PkheVRRi3icwHYnucYJKhxdrrbO+veI57Ddb/J2C6ihOgSAsVR07s58Ob1Gn277LkhLWc
TDBlbDAefAcij7z1EmG9yG68XfgHXEivSpvz20CUqnaadSrB6UoLzyVJ9wh3gMs0Ek1XMiWnnHnt
QBx21f2G9SpHG24mgDDPWWhgYwzLG8HxjWpN5NP2vHQw/ahJ8sr1ABSfowHO00rUgQzbOPctp+Oc
xx588NZC89UPCr8X6RoMfuhtVm6bIiGg7lTyBmWLWzV19VzwNf8DqPDwzbs5sLpXIzI6KoDjJo0C
tqMOMa/4JXgVmeGhjOO70GmjEUthpjgaBq+0lVKqrkiB2Okiw22Z1WFRZv/VKjQePd0tGQubCs0v
6YdqWRZMn7tDCvAz144qTl43sUDVU26PvBi1loSPnHF2rr5fzzcMaNTBZvDMj/7DiVuoM66FHep3
ZHjwEzalHS+xERc7ZIutIw9URom9Mu+iInDllJL/n7giIcWJXYW4Jz2WDSrZ4AcU+13Fn9Iz5KXX
hUR87OhI9JZyB+t1W8VTr9ModeV9nchB8kOSjcloNr8ESZO2+NJ0QD3/Je7ahknqSnrP/Er0cUcM
33c3ec8j1buzp66vqX19960pCrYIDv8SKjUdn4QMf4EewKgrNfpmFnqjtjtGhgp8oiIIhT+4NIhz
dcLoip2c4WgDSzVL2U0y3Ydjvtv1+W+zrgfENHxBngOAhAp4803r758f0rSswuQ2W8FaHDhRQJkt
k6rrLnrU+igtcgtDdF41XUbsbENHW6AUXqArn1eO1dtkYQxwmQtrha/EsaQdAU/MYpeFsj9dH5hK
opCEiLdEzKWVAlJiM2c2xeBoaPgljkNmhUzaEcf25RfBu1kdsCy52GYQNqhR4j1rk7ah3qFk4u8x
ODaffU9977QJIA8JAKK5IxFNqNSFqfNCuiy7VilaZx5fkkVg1syt7ag3AI5wXO0jlc+76veD5fpN
OecR0m7tK408ZIokluaTgDxZe6flBWaXw78FGcXX31zdfc/6M2t7xkcGuBeEBeM93rnAgbN6Qj2O
XRt8ohT2WsoKfSEQLzi8K0osSjXz0yOTNQg+6I7FkXzlWMikXRmb2khoN1tycaouqC1/XbMiaM6G
uP0ld629D0PRBXEzLysKBQRExu9PG+0DTzR5b7E6Qrnr8wIFN5YIgnN9Kgy9pOg5f78a9Jm6PW6u
ABYuc+xvFdPuW87iaDsSz27EgnhjhswW7fMdFsqqJxmt4QTLpf1wjYeda3xU9Qmafd45Vyg0KSoz
P/az1mBM2vEdEcLKzKO8wUHUs74jj+OMYnQc2kUGnDF8r+G30g3DjDDhX8aUwAEX8JJfFPT8pPeq
yHmpeeRGlKh6OFoNwx4LRndUdbgx5W5V24ze5FeyMfJ/WlRlmg9RbPehcLsAg4B7gzIg9G9igfZK
IuQi/G/P48q4mAFhrinM8Ib2cAxHkaAAGJ8H4wadxhGxfhjT0NGHmXP68FLFhHrQx3e2MJVTBaBn
kDSOLFcFmljcMPXHS1ORtfNR19AV4PKvk/AVkeXtkjJHFUaZ0Gf0yc5OWYxqMM7L8Edbkk/4bTUM
FLw/hIqNS4BbZXlCRnu0MKqavY/JzTV48LpH9Nw6JI+h69xMH2YTjb7eV3caDqlx4/D7VgKBIYNN
xOD3CkvQoz318WTGjoHfLIBcmignPFUnOQypmWHJLkfrGHVgDL5Kx+p8ZyVQPt3XXlDZDE7E48LW
+E/74hfwaHFrHxwQy6mBkML+5gmftdygjLcK2HLwRnyZUA4m61A4ljcCCV6/AwCZ3XOZpbOmtxO3
0CP1TLMRRg0SHshw/zBlywOR1Y+OQqqukd17+uR7y7gZP7LwKW6L5zpjK81UaOe5WTy3bm8KmPZR
CXWFRcKbV7IfVjFFfISYDTsLZ3BwjwPv2WlSjDtkW7PTIBgcMDuZMivtHdLy7K7qXYySxOeFFjTD
OLcXDXQeuEEAzbinutcPfUJjTJBxppOAzOB81XaGs7qigsdjQ6lbjtiAz5sN0w0a6eRBFeUz6GSE
zED1nAAK4S2mwqj97AEyoTZ9QOrw6dKESxhR8RSn/BxW5zLnlbgs4Zl2YNHkvbLv2KC3mysXT9RA
/Pmy9ZWVcp8R3iHuU89myma8DdJ+AdkCe8dQs9CLwLncPVV48nJZCAtNnzFD676ay/eZSP1KGddx
qEJ5T9lWdwlFBHkcr817lcX/tS5Rf//IbAtpAETlATPx5tsNqGix6z7i+w2XeoJCKAhrFufZGwQi
9vkWm7Tvq+VbwnBsw/nXoBVplHe2PtEkHDyrVgvwfYITO6tZ8P3Bd+mlZ+pf74CtJ6NIlbucexBw
PF8aBMnvmJqfEorMLoqjZgZU0UYeQ8nnmfyLTtenw61rs4VaxInKLJaVZWKw53eWE747wFP8I+iK
KiQu6BxcWzx5Z4yff6XWkGT2j7Lz6wm8kyo4JbIOBwDuxAckLfmLSzHP4EvOrPI0PGNtTD9tA7SI
OxHzbRokRJ5fsLNTq/Z5bI8gg+cmUCpETXN3Q0z9BUiIUr0p5ydeDVA5XG963zxb9accPly5rm6N
4p8EPv44JbWjDgDjMR/O5LFZi6JKEk1U+BKrbRaDJdS3atA+dlwMmhAd08GsjdgP5RJwBLHNKEa+
ht9NhtcIjxwOOeuZn+BLJwiusqEtKAbFJs9nQreb4dOB+pnaDXf/zp53Qi4vA20mdxkHewLHk/2O
OvECH2uBiuF2Z4qnuoWX2F9oY9OiOnD0nDaM9f1VzFz1rHYbv0i8amMahW0y7ua3lYiJh43yMoCR
p5+7iODYqebTOAYaCZji0DFoVUj3TyXTwHwjSsKXf1lvPWKmHmowryN/j8+8rRmgWgU6Zea5TuYB
D9Fxl+V+hg/J42u/9YvpY+0Q403nHJzFypqvb6HrqTBhIlduXJxrpmeFMQ8I2WsPjIMRl7DvbC1V
RZlpnKShCdH19ynlbqLwj/CNJDri+YlAQmtSFqDjGGYFZyyq1ncKicy+Hub5WSAh27eNpJbIRawG
SGzqyoNWmxbBioM0Du6yg2NvKeEHGbQw8QZvWx58XrA0WTPhvejUKjNNdY+2CkoMyEap9VzZmtww
dSaOUqbEyaRCaXXtjcgYtyWS9lTIYdMAX4oUHrjJuy9NMk8daJz0xeckyGgt2sKFODtLY7KluCO0
L8aI194g646Vua7wmYwTnQvysRi3kDn21CVgUosnVVoJ1VMwY+6u2I+ZGqljbP/zP418ZRfQjxX4
ozSdDuvt2Xi3oTmR07JVIm4a0pDvPQGUIl3tXoKYkrSeBNovWOJffhZDQgTyyJfAQeyNDesTNPGu
BVWQvPt6azDMEnu8p+CJ8VPgsgXDAwIAXpOoMlmCMsIZYuokth/1Herfg4hVaMG8PzgUVc0Zv+bP
orvwVIeJR0csIVWovW3mZpq+gAMWwFn6ofAZIvJXXIvmxxB7KJFKmY2Wy3S4uAfCcV1UiaDHpjN5
EMsR+g7lwPbL6mRo6DZm4Hx4cpJHgfHHDn70cDbrnOxSN5bR3Iksdoh6pTyABHDuDqUk/7gn8lb/
Uc+oKrkHLp+jHE7B+YoCgkjNz8y4xSDKeE5LPJnChgOXq9R5z3g3r1U1w+HzHhI5LZV0hnLhdbR9
lWmESX2lhOOl4NHZ0VL7pT5BSl3vQAPQOQbd3U4qGXc4WhHxaUPw1zr0ADMQGwDD2i7bYBP2QyHr
BH+AZq0m5pCKyo8zMuDr98X5rgxWuHmCug24OsbktZwIbJVIBXAa2rIeGEKoKUxlJE0VNzbud2jS
lV6bDCuV+eTu2mXSPbgut7DB8uCC0wRpe2lPtKwkFA3cL2BDmF0AQ/deuBUCITL0/WE6eQv4CI72
A4ydnTFBemxWQ12StTi4qCSORtnMs1equ35CwEo0A72hB/uCwDj4S/a5TptSSpZ1bCkba86H6ZLX
cSVLccQdo1GG8ABzUjagDkKdWSVRdTAk4lJfPUYls+O0bxfURr1dq6RW1ibd3xTpYKwVN1iFh86O
AKmaI9Nf2q+Ckpq0SACzXcu8u65YXUXeggGDM/nlhQjSMohSvulC1vJ/4wWjFPz5THU5xc7hNYR6
aPkasD8sFp90TGJHoz2miQvRIlFLMnpBOZasEG4BImj89/Mx9c75DI2UnzQYOKqRCr4m8h6kSklQ
+zSG7tveLxO5eswlmfnxBTBL5Fjbu0PqH99Vzftvmgnxc4rk6biw6pCzjxWzccWV4sSfU7XOo5DH
eNK2RML277C6do2MYpRkUOXtvDDq3WIEAJT135ZK/VvOYdyVCorPbBATttzmHODCuTW4TOpa58rI
BM9ktl8xtaTEp0/BoelHnHWIVdvF6JqCjEYzd5iHIMIBS1Dji3JB3nKYE9+XWpxgqmpEOHP+YLUH
o2Dw8EMk8omqQGhn1VV3kgoPJ+jAD0MmgOAR2TBO5yDe8XZaofs8ijBXjb1ERF1huiqFlyb201xV
8bc7iU1utm7Ll1RUKc9ikbAYp1qOy/cZRFz+WQJDeW2cqidM+lw/f/IkvgHJIQ27hn8nxTgoAczg
f5zKZv/uCvBoa+8Ld3TorTFzyo91tnVOnfqhRIoHyNy/NcZMzJr4EzBq3AqSV5OtF3VQnhfDgfyC
Mp5geK+IdUfsJjJiwSXk7rNWE1nPSf0e54PE9I4IH1+iLIcoyWLik5yQmn4vGQrHCvaQTynZxzXm
jg55LqL3PTHauj7d7Gtye/wF2Plgf0MOWzRyup/bYxjXH45G9khzYBovHdKN9Ss9O5HxqGUBFmGU
1LGZdJaSp8n4byxlyjbXPEsO56lZYaR59pk8Rg9svXB8ho+QIsZnQhOyACaYipY6mO+0i4SpImIW
PAgIZhl4+TpT1HZoi+P7h3GmWd/rImN6cGwVzJaUUIjkVDhQmD47k4u4JfUjMlbwNbhJVtjblQkE
lW+Fpq+06wacmidNh5gzfWMRxaQO56j2hSexfa1/xSTBx8omSUCb1NKJYWIz3ykcu0QmUYTUgBMh
hZS9bJitun3VCbItwHQBhzgXOrBFSa7kzxZDG5VzKM54xi5JebHweZrwU6+lfLbwpw9e21zLQDQv
Whf8cnDi+6wk1rEEdpM2cLS94VvJMVTl2U8ro0pKBpuRsQa0ih7hrYVIbFWwyCkshmZUfZAa65gH
HEql/xASM0LFeWJAxunEz52tSSkOH3s0WErDNGZTo6TgfLNbFobh9MLJSrx3gdQgsgwvrNL94Byi
PXgBOtU6S4D4NkkJP+8FVkD1eIEjSORhGfTGp984XTEXn/NbziYdKu/EJy4bdRsTDClP6Z+vDq9U
IiR/YsUzcQncBbzEKgdapcIylR+LveyDyI/ddyX39r13ESamYVej0aZcxF8xFH9xzx6BhNvplkuO
bPVwbnRs/zqd5/GnB564rzuqjxI9MucqQWZCrTdlYaNpsdioHHJEZzijMb5hxauXEkmwRzn0a2F+
hIMlWd3nAvvODqP1oAEjym6M1l9fUfDZzAl9LGIv7AUi256BPwRvv08uXMP3ufg2k3mMmrP3C8HY
xCF3xA3BVJffyyPu2lmNySQKKiiTZIv+fnTuYr+EiPVGTpbCcA8OXyAXutxatmzipBsHS9j/MHEb
LZNgUbPP+p92m3Aq4PGuNT8mE/EUPPlOvqqEAoXwtxobv18Xqb0INKlOx2UlaZy3id4TictFYEmx
YlLmu0ApWb+myAEJbcfT1W93c1SqvQLkv+21tPkJQ+bvaZKAF/fcyF7iDbv4aHxtIvCmbcXQZOPo
c8SIaLq3OOt/v0NnNkrQeZjqbFy+8tVlEUZRkRCHWMJKWCGLH9ctUmB1uGpsqxIn8jAYhXBAewuA
wliiiuS47eonawWx2j+jED3H/3LDjRS87sM52CZ5LQ6ZSeI7gXWcOSTGjiHPyfxebUkx6XdvDlM9
UoLf3ahlDN8QTeZTpc+4gd2BB6Hev0gImBGsG8v3d8HquWyU2RyUgJHVFHbzXupY7ZFzUGIOPcWZ
7jSBKtg8sHsrPT6T6rFsVY9fnkFNOlOaq1zuDqkvvXsek2uTw+W3KZ1rzh2qWPoK4PJJdRYC0Iar
4LrCLSOfJkCsNogYxqa/MPlJO4Z/DX7ghAMmkGeh/P+qI4s4pA475acfoCg/VAI/0t7fmEtuNFf9
1xwZS0WStDUC25DLhuvWtN6Cx5xYgncI3lwCSGXxbSWFW5UdPrhCBPz4epFsxAG2CJ8JjX8C5mg1
+yWKymkVvIFJ/piO5agXRNbVpUxlZDPMzq1n1LV8dVcxkeosxVPlIXCDF3uWa1jhmYlloYSoX5zS
aTrSF0o82kVfe++oxQZ1NE/u7KQ28YnAQs021zy7QjrCpvNsYdlcaiqQKwEHxq4ieboesFY/Bxhx
e40qVrF+XRIpaVsmgTJXhxe+9e+tVuZs/X+3CkLg7XDKigmR0M7eTQBktA/K99y6QsYOm3tMtWiG
J2Nd28NsvvTl2P1TKz1mRMuKFUBnNEXqkFgL73fZLS7jSGuBgqaSQwMjFrzc6OiHiVShCEWZUZsZ
xAUKX3YzcFWbG5KX639CFGMz2x3CMx+QkYgXcqdQAvv2GcmshIi1zTNIZOaBi2IPnTYIxNx8oHLZ
Ka+ajrcvTB8Xc3RK1OJzVfLXZLvrQ8zAPx9y90URSTwC+OGYnAfFuD8d+pCcmgWM8JSDDue1/xvS
iLEANmwjtnT9RQItP4kPk1yTzR5jLq+Eywcz6ewRhUr62iRwmlB7hzUj1pUsdijPty0JTyv6fR1Z
+JlkmGnKy+fmvKp80GNqkmvBoHwKbiPXqhiUYjm6lUotNxe6vVMtlWTFqiCGoWYAgVLi0avRFCU+
CrSdEhKiTdFZg/3zj774XxOZpf0UslVMq+nIXJgMw8X2gh8jeZ2NbIZS3OQJSLvTbENz8l/iBXgH
9U4mhf1P/tII85DHtokivSyYf9EiIlJDtil3i25iiHOl0ETpIP6EEJhvXUttrnDD5U1MPcOWRxVY
1OTczg2xE6PVO129EDzk9WD4S2ErKQCWtgvEMo6BTL1h0XRPxiOF2DgcTb+X4gxMx5yygwXB5EhJ
1m2ajnoUh0p+0UjqK00W+xCXKf4HMHMPu9npjoUaVvJRjP2eHti1I1vGN+17mx6gNP3hoKydOlhP
ZKneg0f81DBLCAwmBZJfitw1mmcmz37noWGmn7epaIzzZ1MzmEB7C4xp+bOvFV42OODDkEc3sFG1
NtY1GD1YxTlCZLOyBb52ZwP3f+BFpCpTMk9/QZFWp7BJCKR7iYat3bp3IxEHdkfrRYyuzSzR+RFM
Lw59q01ZYhlCp+igMYDEccntxNlGk9GBN6XGNRB4gVylpc0bm/Qv88QrmTregd3FbdQjT1mky+eb
7vyiTxCH3qk2TEomWpDK02IjoLVL7CH/htvV88GWFPqqmIlbgym+hI4VCDGOX3JCc4TUJNOAnmqU
IxTBdiWhWW3WAK0+nEW3v5ws2Zayt38Co021ybXEgnUBD/juJLAQDnfSYG+rvRIeoAfXzOBTgieS
0IVtlSCoWRmFEg4Hp0DpzEXkoV8PKXTla9HdgFLj00CWK0j7HhSqU8XNmZOcHW35oYOl4tRXsy55
5woShRMsAT71+xrNmHKQOB1W/VMztO72YUaOZbuu728mUX6xEjUPhafcasYFYWAjtqrF+1e24Opq
bpaEgtPGiWLxvg2DJNHuX6JjlZdcCbQHHEp1wVCXZLNfi6P4YhrCEpAu5Rt2lSPM/oNKskO3y3h8
r6Rw6DEIa2kK9SgtO4rVj88JLMHgq7BuOzn2KutG9QN6YlhF+o7Jak+pjkTelEk/KnfK28OTtHDf
fUo8wLqzab6+OPXi7XDv10qF9fjocb/vxRLpIEonvkzQT5Ag1Vtgl3kWYockyTm9t+YAZPfyC2xW
ULf3T37GucTWQto+FeZpzcuzCWwzlYPUFSxsPxpY5hMcEQYYRIQzyA6JMThOICTyPBDcWWLeqjgw
+IVLc8jo6GV3gVy30A/dM+hQBPkJ1Cxu5SHKYpbssZ9pArzHI90yv9bZ+96yXjRWRDTzqwdPWflV
mkbo4dKymkD4yxg944adKkHuO/p3NqtivXtIyPN6tQTN5/DLCXfZTLgIQrYv9IzuWu1mwGkWTpzX
hqp84UE0reTgXNSSHQjXa7TxRWzYyJbJeIMZfXoQwU2u0ZGaDDE0zyhArjjfzN27HKtXjuLB8Jaw
F5eqLQe/LArppKYXMtscbHtzsUY/j8gamUeDXu+xjq4H+bh090D509ZMkjY4Mx2AdM5RaI+TmYP3
uh/xWgUyL9yE7WJ6Ju1ZVXLLAiciKEGVhd/dRWq3AcQnJZuAPE1qHoKn7BBMhhZ+iuNF6JfQCfed
/WiSDmvOpKyOyl5ts/pRhskYZ/bZy54CDeuw1kq5oYC2hNCN0T9Zu0D2uGyRHC+TJJwdZFMnb5nk
dO2So1vtmmrryQF/OQH0gHJm+Bt5d3HcAeMw4vtfuuupciLxzkNQqTN7Rn/6JjUDZyHy2KbAoU8m
Gy760Ez2UzzaM7mGd6mJNIvdVC+WoDYmdhE28YsAp6qZaNrV07lWjs9oVbbKqEKHNGO+vjUHlKY7
thlPBH7UPlD9PwPWWgeHNOwgXvjQEZldJT4mR3Oo7+ltlGGgojsoPMu+S8t3gj/DGneHgN0ihkt0
YS9FQEHAYYqfbNxB0GS4YnhFSmlOSjDHBtGzd5uMQV3m+1VHtHaOeZuAM1+LYk8azGCmiDc4eO0d
1D5onjrWLVHmJ+SKREon/vuFp6fahahmyposB19b+9Uk9R0BEtrvSnJkI3CwXm2zFqRDTBCGB0qn
0FtRoYK3tyBt2sGJDCGxaHGos2IV6onIrJ2ofGsk7kC+djjKqBA5kJmWr8wX/R+3o5qSwmpoKjd/
BV0DDC+E5+j6RLGVDMcHtoFBd89NuUFu0gdatu29HaNGSXltgsH8OqrltEccab2G6GDU7rdJpWiF
BG0uHsgmcEi9VHhMu4zF0lFrOERwYYZ0+HKcUUCSqPEFSeyra+YtP/WHra6SNYGIGtRqWzThgdbh
4VkKYklt8GePWF7lnKX8PsVT28bjZhJUWIrvxMim+X7CQPB6hko4gvK66Hj7zuALONnk3j8v/ci3
V1hqsZe7ALSQicabAzNsmvDcIoGEOVCCIosGDzlL95kCsUtudcGMdkbrvDsUuSueN5X4jIjeStpG
SeZDnWLt53ZzJ2McDNw92CH5QMo/TxVSa42h0ClpSvL4aoKu+O6JtVU9JQgchPCrVMUHZ8NMjLV9
98ULYn4UNk8GqRHMK4chCYE7Qn78DRXER2eDfIZOMEYG1HyYFyb+nxtg/MbcikUhRCXYAdQXfmts
9CvZ/iQeEI8VyDIhd14csfGgZlM/aPCabtFGyC6BkEErwetqwAudFzBzmS11Hrpq3kIYsykVoOli
4aD+LiKpfaZ47Dc1iXRJu1Uve7tnl2MF9MG6mk9a3mU8AxEd84h3ThKTNVwOzUwib7XzhzDdgpvU
tCeqjvFI37l4vdzhiuTuTreWpxVu950U1t7TZLLXmi2Nhfhu3LMSnx+HsOGboY3f5aB60FxAXwie
ht8SQ13auL8Gl47k5VaNc6PJAbQShqemLkvEv4wSzT+Lnpj1snddif8Ap8Hr11fzTR5B0VjtHh3p
1XvO88EAwP9zqCldQ/nZPUTW7ucI4Wy6vVcmT8MHavt8MqFXqJI6lxz2TrmueZ71ONCieYtDOtUb
pEXgl4P4w4Ad2nEuTlBMA336t//snX+asN+mSwgCKD7FHGAXME4bJn6ayxqKI3LobUjHMEs6Ed9+
AW9JyF823pWunLG4IvNBX6NUQtg2vbthsMX+CWz0gndjoS/bf+Dv/+Q+qy3nXPwxe1P1d4szAnwa
IGTRb1W+/mswoMzMNAKEVZKPOYh0wJZu6/b6D9+rrsB3dlH52IqgIisb/D38+2h2AfixRkJPu9rE
yOsHfiQxGysSdfh+u1noDW9n17G+e69ZpqYcTEsvhg+4o85IupHLUjTUs5KIA80Ezy5eQpsgmemj
KLVkuL6O8FRN0/h30h5hLajmIHpFZUm9uQ66I9tnZIvRBGQTgLxlNun4ZGqO7wIHHAckIXibqZ7i
/E77EiVoZKuuBdERCk+kISGlls+vgtX33+AphVXc1ppMK/AvI7cpi2ngI5jkVPvPJVnJARSajfLi
Zueq0sJtUH0XAquuHfYKijPVz0MV+XBZV3b0w5jw0pKx71LzGkrxH93oEeABS07DPK7juWXVPAqT
tUDFeRML8XSqRQ90Q52QMbojfLH1NTyhOVssOe+O5DyZ7gErRtwVj+5XRQYiqPZiwoCkzA1eLppV
7ZJVelSADUTY4dAByYwmM38YhyGQXGhoB/NLtC6wRowRdolSphpUdihDXBB0ElQvhnPunnORz4Vx
KpxNFp/qdnAzBDpThMIetOmSG4Foc+hgQSHBbBa1N5m9znDbdpoUXVLKgUj+ii29wNB73DkPmrpz
8lh1mTkfPz+6mYQ+iEAd85guQXdLGP6Mn/aa4f/akwNuCEqB/OPYo6BJIK+y22mjnnOi/S67IuGm
9JIOKdpQimHp11DPXBXZI/z0Er0zEA9db0sPtbJdV9STjzp/+oWirfhQ0cyNp1w4+KEjVacM08NE
v3nplTRd0Z06dwkcXF9681/kUqRUiv6ZN1RLFgAKFKph+4QcrKFPXXeBQFlKaGHVvr2fXchJnA6Q
JBCuv/235xC5nlwFYOsMIkTkgqd5qChmA4tkUdlRofhc+v03q5u/+eoRl4O8rZxASGaKV5NedRBk
7LDzpvLwt8rrWYLMcvK/WRPdbS4K1XrebtMO6/uD16CZfidPdeuVfONk8pSaxRxMiTDOOgjVLOxe
69dXxU+rfp6S3Q6OBr2eTWJjjQCxWsB3iUA8PDeDyYvQmXK1wIBgvCo7O5wsUradYKNmXsWrqa4w
cICPEup4Ry6UxKbfPEhMrYNPRVZjjQp7r6CZ4S7VWAkkPQJUKSPHzQdhaPN04XWp6EK1ZLkuKHkH
RneLMJkZH79KOz1sRqnMrzzUoE5ZsKueWNj/v0sA7S4t1Elo9jaifhdAfTkPb4o2urCf4iexDbzb
8t/IpdUA9Oq4QdFYVycTkeXwQwa8Sg+AZwbLb00598YrRqPGEOrGMO0ITH6iDGeteGxFtG6ngysQ
oFe0ZEPvBtflmQ8Js/qZMwUajioUImpeqxFT3mLaw3cd0K5m1aL0kVY2CDk+3joKVRn5z+rkkXlb
OSxV+5HH7V5BV8ghmpZ78jMSRfTLQ9TBufrfIJicnrCkPSrAvfk2+FzHQlaIv9YNTHif9SKyjO46
N4aFQ1XHsDIjvvj8P5B8tSRTbYLBuiWVU4gozeGv59sLUDyZ/gBDJngPptlbAXRcJxPgRlK6VrD/
zDr2PKks69LrgX3zrDF5uroBoo1LLRd+dfra+c7zFSwGeZwci1wNRpRZKhumIbhATazcURo9WgtM
8J4z+7BOdI7/R25Zc/QQJV4eFvHBO2Y2LwYur5+T9TUwXrHmvRjpdvc1l+Eb4xYK+WGBwe5ghb8M
y+hVO1nzhaS4TAf/MbBHgftOSfHRGDpHRl2XxsHDwRorBLdxYdUcpXrfLStv85Yn+KVxGT1S0WOS
vMFeLGz4f7wDWmlxRw8leEMh6uoxfq/e34AOy11HuhRWwLG+KzZXVC3srj449iaWcv/GbQGVgCzp
+AkuYwU8IyOlvwSdn3lczS7Dsm10a0/aB7IAoLLeW1ssrIzYGHRP78AXksWQNpe9r4qta1xHUxbF
dXjbxtY51AEJV0jR2CJwzf2SSXgzPrmmj8/Ej8Av1vUN79vRSb3rGYQ/34RFGC1nUuu1QMFWbbbU
ldKgDVc+V10g8Lvv1KDhDYAwmG2yb3J0It3P659jUCCJwATyLu+xEHqloi7SOPTNi3LgUBuMYnNK
xa15uJrN4KTaeLYzd8a4jyBVFS9bBevr6czRv1pZb6Iscxfhbzf4hFu6rwf76WBV2KNi98ghgtOc
9r1l79mJ/4SeuqezfWeiaqMw6l7S0jwBcvLH/+PYHZ3I4V5gQrcFFKjrMy1ZlyXrE4geUGzkl5jt
kUHY02bnYRlO03GoWaZfnXShKp3vdRQVvQkIAqtTGbozetpR+1URCHIRzXQWrgSQHb91bCqwUjw8
FtOQGED7b9uClx2U22OH56PCHmCvkTw+JeJNdWx0ORx3FjQv+r9cJXuSNPYX16+KWCwkgOwTo04j
QobcIc4vRTZJW79960U7t1GHENCCUUkAe/Jg0dAKVXgsMf1scTyFnpasSCsqfNWWLqg9kbgeE8OU
77equGUwmj+0N4+y8Xnd3SuAsN/Upun7bQEP4Kr80qN1ziXmDwU6dfMNaLyKJQA/mjKyvOUKWxEg
vcGIumeUomEjRidTeAZdy1lJG/C/fSfzPSJ4fB0cRrPW3M5NQ+hr4214iCVN+pZ2rxvZoyWey1zU
o56KRGoymeUvWSgcUU1e7cCmyNK1NrwzcreppX1G7xBqO2OmX1UOAYKwleUOP0+FnwEMzoZh1ojw
BYwxP0yL1KYecOjs2aSrEOfzqhkE1mhhG3V4xBIc+mU7x4DZ9+UzUnLAb5WwFAiFnbN8Y+WU/1Tv
GxTkX3twLOfTkMLZUSKuszpwxneBlt4ngLM9uis2lrkpnYiwxNCzMPTBbdsLDEpyoBCRseB6dk7b
Dc9deJKOzzA5DWCHNJScoHUHeffYHQR4Qf2hjioVIlrtg1dvODEZ2saqLoSfWKQz0PkNRr1T1dGQ
96oxtPbspZ6JrmcJDEdVrfNwak+XYizXJe5EwwXKgUaaaOSjWV0hKZ7Pqp34K7R2P1pYAuSlEaTZ
4lE9xUvDM1EqOjHT2ArEtUdqyMK/Jw5fq/Z8X928FattGNfDBlq30h0UFc1QPXrEevVhH5aVIlUT
e3jkw3Vd2hoNU77OkifLLt3gf6m9xQVJc6H3oXc7WiOKN+oZZ2APVQ2u8B6RltOf/2OSayjI2//L
8aC9869o8yOI7QaBebwEr9InNgyLR78P+ztgNyoL9FB8FXFVo5VDNgupyraIkdKpZCmndkKc1DFK
1b8W/NZzzK1n+dRFaR7Rz+YkBNyXwmFTSBcmCMvJE8p4jSyb/B90rHkwXp2SBwyqn9wFjMbYyEeT
BdKvBk6du37KevAHYVgrkBn/IoWUF0Dqn2DEmFKIbAoQtxKHu6zCS7+lpUaGZd544AATKTmWDzB7
zHQVt068TZvzaFPKAHJR/F+RiPNZFsUpntOqogiPFJ+QxMU118e9BgJWDff0o26pql1Txz4MgV5D
nNe3c2WWaCsgZSQo/lzZk1tAJM6Dl1W3c1FTwcE3TZA9HAxWn9/gTX2MOpV/3Lk4SW04NmUBVVNs
j9QYNBCaTIG4ctgb4Bvx4lR7CeeBKO6Sqc0+zJhFyYkFuduX36wqIG2i1AMnlcO9r4olyXGKvXZj
uHfzDxeMShmiAFe4hFMbhXigB3kHNuEJxMCKUGgi1kY1F32IENTswz3oqDFVHkekRIKKR9mgXROf
sM80qeFrB3plwyDAD1mVvLu5MqhDTpKcWtrVuTsyHyXTQ47homowminhJQEC3debSabo7xVcmrMU
OjsnKposQy8+tAzrszrCiBjHMrb6eLlWEqXoCDSqQWvsmuRLjbwNCP5PtIgwhmycLAQbOKijxit2
w+ZbIK9J6e+IiRtefApl7MWw2h7uNo4GqdS9eQtgFFdlTt/1/zCzZJqM+gchLOKou4BHoFtzDjwC
08mqWRpShArqC+pW3davINmGEEt6YNRvEObj9wOejfHApU6677sLsqZjOFpDp6PVxCdQ8SJkYbxH
7kpBJAYsghMIOXOKWTyM6qcPNpTYEjP88zqeZ0GPHTFVesfwzxd0NMAhh3Nxlh7SGzDlbHO3hu20
yJM54OpvRfTS50MoJQ4G2asRFpEfcfEzXboLgqlLCE6PwK25s+bzOpcAv1eJGQ1wTRWiAYPHcKJy
KiVbEZoFWdGGz8lSr4n8AXEbmEDUdXwg6MWvJfGWBA8uF117OWC8Tamt3F6TojpkpzI/CJa6WZ1u
J6NvI1ydYBBDrdNA06SKA7dCaRwpMpfqDLAPj2OFIP2V/9w21oigvkTQH/wCD3Hltd8L4i3wP0KN
kveaZKfe+vKz+Upm4xuiE5xNAX2PcNCbhdqMR/agQohvYnUy3PuJJ7qHIkzVowr3zG5CfpvJ9p2W
rYqzvRLxxjuYY/ykNzFOeHvSfzaLqT0sTdWCquwDbTJxNbQT6/ELbY8sgxEhuBaY0XyLIXNMUjaY
BfDbT7N60t7a9rnP8dCsJR7LpU1HVYSdj5Mqs+XevYGYLHNzE2mqNR7sXmUem1s25egrvbHgS1by
fMvEub5EHsdaVKxyvS9jWF2t+fO5K29zvf2OUEF//388iIJKa0Pkk8DXoP14G19FtTE1TALz2uPM
QHQJkW3sldyEWnWLcOJIPI7T85IuYPiCHrmp26ZIS5iQEIJ5tWS9Jc3+qd0hnXwrKhVp6xKFoSYp
NJVcJavOsBLa40GJEc74OiUtzF2l0tOdNMGaVvlumaNq5j/B+dh4CXZb0+IYvoxe/ailU1ThlmZn
8nnGg4Q1vxpeovmx/7SFe6kDcd+dzNPGxFNeS7h1y23pCJFcLdmyxuPHkJm27S3mTbLhmp/yQK28
sOkn2sSZluendJKMI+xzNNcUr6BC01WH7ZKh9I1LAfAkdNYpWsONgmfqOi/jP6xRp5cKtaLoR0bz
Q66yev+mHcBfCDZHKCKVemMWCJe2rYjkuoL7HAk3YAk1dxjJKDE/0N+usM6HkZn9QEeFRdLnWvre
2dWfx0BRoon+oWbfXIGlTdo0cu2+Oi+XXyWbFlhFPm3OO1LzySyZh2mgj1avR44tNrIviKIlRAGG
OIcP32k/0g6LsH5ORqfIoZ6iJ/CpTQce/ofr4kHnxFiKaVvpsmLqVHKnBZEw+Vm7BHoRCpw1AqvJ
QcLY1X+C9e+imQr8drLJs3pcmcRgMhixAfg5bnyQgmY69uZjJgNc/cw26/U2HRPGtN1SatlT+baO
CBwSX3u/CbQryUL8TsphBHAGYJtxFF5VKiX+ONUuqo4ykotWwJtpzIpYKIQJDgTZ8Lxb+a5wk31+
eLw2fzgBNqEZAOZuOOYx4cJuGaIrGpDXQ2giSD9PJZe0L6EipsAdpdpNXmU8DjRTS/fsowlRMJmn
XNoelcY2ig6Y0EBby1cJiBLXBwF9RRC7lUrnDENZlrSvLl1xHjLrBvBhwHgu4s4AgG/21vAwSBUo
W7VR1+4V/nKpwnVZRAiWQlFdqIUDs97DtteCJBg/4ZstQ9V6AcMMpGtkLAd9Tv57tnbAunwYaTFu
CvgDXeoUh/QR5bbTcwCYOtlmuocfnNeJaecAQx3EGCr53xwuWRnoa21598L72Oq77eeWZNMZeM7f
UC1x+eywsLKKH68wKSUhQClVhGUfDM70Yxai92lXUQuHnNlKcPbreEPXtli8ywETohtzG32+c+Bu
TiYYtiqqDBEWCQJcmT2TnhZqghl9IAB0EjV1ijDxKY6U+RydyCu7ERTG15T5Jrk/CraNTW0crezM
E+yphW9FAIuXXyHI7Xn0A6b89c99qP02lBCJkMFoiAhwrbRMi3XL1SwQU21UJY+8x/3s33S0105E
J5QR2ROSMn3stODJrLARaCk9SgUXQ4txztF4EmksxtLEqZnCMWOcTFBzbadUAiA3epDqEoQpmFhn
Clru8DnrBVASbiKp6GMY2obuByBy3T98+q+y+1z+hr3/N4saRZpyBRDjkq9WCvcu3Lu8nb8/cnhD
QDClKPEF+uytuNioQfBH+tha7l6HjoG+O3kx/KsHfVAg7vB6nzryG2gbBvarsOaHZoeSissNtVJY
/LfuXKPJbAHcvNRStcmLubGfHYuF4QwC4lB4jxG8trNzAcaVftjrouuhdb3Oa4sFGkUAkYI2zpwJ
AxDzMBONUz3TzI1vyFYFeREn5HEsF+V+nAho/0MjbZpngCUXDzD3cUmLkpG8AXVyuUkvnx3dObfR
dLaTDF2RMCeMezXLwa4QaiEW9A7TqX3+OBvEiWyzeMeDjlRuJSTwxOFkGMVj/fNy52J9hSBuYikj
xU+0az/2j9eBpiP3D1NgIvG05V/BMLjIvxt1nlY0zfKuhDeXuoneSrov1jbNtT9m2zpe3W9ks3Ic
gBrgh/dD7xGHvkHIXi51xvzO9I/NsPudI2rSX+/WFpTtjkzJz/S0MEfOsfvjYkM189AYOj6FCpee
PZlM9+d/tSY+fCbNp+5WZla5d8PYZ5rdFNqiicRDw0FuCY51V3LK+dGBZE05FJFMxqFQvCClvmDM
Cop+SZqgwVBRjKS0WZiqswiFW2DG129uWlJP79/T/Y40M6XHeqRaoCboto5EJSbpPbv5+7bTJ4V8
gnba2EmlcSpAhfjHyIarH/pRUSoWfdO+x6FnnYj5nFGzdv1lwpbbsQhVrAHOtKmeMJf5AXmtzBBv
s5/WsLetjSOMD0iv9k95UyB9Us5UP8XQY2RbSwyrspoRdKm9zrfde9uBxotWjLekUbCGF+WAZoLA
mbU8sTb5btihZBWYhH6hmay4bNC8mMqoZv7ihnEY0mBkDxnQ7wSYY84v/PjPrboOT7x172sY0Vf1
jdofWSi6pqKllq+mDpevgwO+UYh3mPQKZoQHiykuUwrUiipJu4SR378tCdxzhnBHV73XfVb+2aSs
DVDWXStgv5PTwQb/gcRidVLXVzf9QZxqhS1lZWR6SkIVFnCdkzbQSkCto9SMU1amVtNNuSJ296Mv
c5PshRvJRej3jrg66PxHSGcu8WkKSB93SAWlml+Wltq5SoCNfcjMyHJ8orMH2XNUqQKSXOTOeAR9
NLVvy7F40N5FzbK2d4YzVMQCJfkCx+YgeKViqSOEa2ZIPFvTvOcTP/EyJAFdqwz5JVasC8RaNwbm
5DzIQ7THbhrVFxbQCjWVp6oI68ONrJBEz6Lga4Mb+oyRIcfSHYyXED3g8hLtwwg9/ghIU2rVKkhc
Vhn3R0eKcIhU0D3T3bhDrmVPbY3oW0jhOsSDc+xCcpSSvQZKmfUWKrJNmbhaqrbtUICEV/2xAQpW
u9w+rMweg8b/kAaS/mX0nx9RtLU0Bn1F5M6eSDwcXrujpSUEX8fEW462Ug9A9cy3ZxL4P+Ci839D
hLmA6y9ogiYYXocMhkspbdf2OWR1Thx4ZCsdEhPWMqHeGoVj0cH+6DtYHVZn+Ht9vgNIW1mojK1i
qYLERx0RLyimA+OFdQBcuMsWs9IqN04fCkI25k0OtEopChOy9LjT1CgKHUWvLAZ423kymERV2wkX
knKc0NFoF6kx8SQXSFw0CqokbJ4GecCqWhCqYJUttJJWRmXyoVeU709PndyfttXHYQbXf5lbCUS0
ufl8kzNdJeq0WN/bgRKVuzHq9qVuNOauzGj8exP6ZFwfH+jlyczFisC4su/UH/FziuQpITHlN5Kh
sREPs3HQdKIPnEOH8hc9UUoHxKKyfLlgNgfvhQYQgjbF2fFgIXSsrE4YI7Y0te2b5maG1zWdSjW2
Ldiv7IdHB4Vmxi4ikB0O/ecKlPlZv31fhdKB6Zp95re8PzM0a3rdZA1TZXa/JaOk9MhLFtZpZ/7w
KieXuXlQL1dJzLjcBboKboIytYTbRqvocx4XQmpWU4uCuUuhBRH8vtruBQBHC9vObhY3gl7KjDq/
iKwRwPsWwKtgbSaHOA2S9RrJkGBf1Hf8gh64VIe8uF+reeHYxRNOIrW1quPoS0SIsyxZfIb6oq7/
2Zns/AOTnhYqC+g0DZ7Fu5vYulvWqfZ3iKs3ASoXeD3wBQm9k21XuGclDhTfz04FB7pYoGi/OYJQ
4zjsco1rj9mFTwYvaPJATpW6e6+BSY9oB8vKvlI8eOHZJtSGxffEpBTbN1hXfGtXNWuTvPrRPuYk
mTVBvDhYu/MVsm9pZ0jFySe2QQVjRh88VuSnDcP0Uncuu8koftC1bChzpDYfPkEtxgm7SxMvDhgm
DlDIKY+hgu/y1yBb6KGbv+kUU+FnG76OmQOrlfQklEmCLqOoGM/bIjYjBeYs8zW8EALRPOl6NVmx
xj5PQBYhJsXlNRCFAOXbkJAciY9PizxiVx7Wh2sKXXGvye6PNthEumKm+JKF7nB1fpBZqzY64VRo
kYG7fwKZ4AiibiI8iA/qmc4spZSXeM5/y8w9MREZq14+Jf979XnvMCJuRkcwOi5+iUMr2JmdhoXd
AlBx8Ql+KIMThnX4ULOTGHxAmAd7J1ZX9nFih1dIagdSwWh3I/JYkyOZtkXAV0cqfymV26TR73az
FDN0OufOQsLRx+7y5UvG1NErPRvPSFscxiW1qorTDSnmGcW6CExU2qxscJ8kDH+mIea1H4gTRRX4
FFzf6irT6RTl0wuS2hlt9tn8f9vs2CwaZQ7+IKDSv6oRmnRv0vEfadNbmH7t9ho2hHD47yd65lbw
fdgIu827kEfn9xo3pi9fH/m2IHHHINiRF7OwP2pDP1WXqIPS+zWljvBcV7Mogckt+ulNW+r3iP69
ZpWJw6qgzuacmFGvSojBpqgokBXGNTEYaBtN2MvuSz6AGM2tvXV0aVOpUPdq3VJqbUPhZqIVtOlR
gHuI+MOgBrKLeKes0bym19t9VHgLBg0tYmpxmWYFnBJdTK3CqHPrvLDFs4E4wk0HkGsrxmLUoVxk
0ZEQ9k2e+DQ/3ZuMiF/wJXjAZYd1tKUuFdRaJiGdbVYIw570Zgvle1Ud5lJqkKU0X8ilT1SchlNe
ZDSDYjZXBtcSV0qQgsHHDd0bAlWfCuPAZKrgEbD9fuqVyh4kWXhTnP2hcEIaU28SArQATliVaD2J
yH4GoHJi+dI3g6EqR6l53AGB667K94oZ5tzDhTp/tItcxt9TyGrFQ8iijqv2UfWzsrAEkKl1rzPq
QzNXkvrX9piY3epj6lFsX7GCSTSHkhs2gJ9oFAwOYKr6xr6oXNKMU7ftdig81lp3W+peKcypme/G
MLjv+nlrhKx5pv5fwCOcENy5eb5Y2AbZdq5MZzfcAt2KDu92V26ab7QSekYahHSiaOoMR3dner7U
zajxKqIaOKTaGIcaoUjNOJr9JQPdGv7q/ExrMtwIDwzzoEC0UBqZf14R/dnb1NRB1C9EPjEyFR4w
Caqn5Z5SXvSaMdCVGo9IW8piTqHL1UXwYePW9opU+rrRGsMcScYUKOzd1Ka6E4FITQEiaKofSuMU
1mm6cBzKqVd3xScdMnb4I6vUZ/rTPpVm2uqDk9i/iyT3koEfLINKxRlgpGPShpj2brng+RQDKjGH
x6pLBgsROTXKHwbBPNaOezhBJRbja8VQwK8lcF634CvX/f4cbGKxqDoYzFRMzp0iqWiYzzh12pkT
XMs/LdkMXByq8fxlGosagNTeydOOXRFk8wEXtfrjympVCzm2aWJ2shDX8aiKBEBaN+eSF7jnf/QY
QWM3HP1xFN5m8hdOgRq/sBNKjE0kiVdqK8iYWSp1WQq+7sgPcTIh+x5Ub/1zReGICnTEk1wMFQAS
JANmJdt61I+SOnhojRC5z5GgX3AXaS5U9KUwVg6RoVZ0TLhPpN+MJS2SUGbC2v5txs9xuh/2Y7At
DGpgBBLjO/wCEtAyBcNaQwDgm+QywmXAOuA2mnRA9mSi31pQZaWx7a0hoB9PCBcqk25i9veQIaAQ
WQIPPHYv2agCnIxez9D+6qx2wZg3hyy4s6FgqRVZDj19QtWRViM+IFMoWFO8q7Oeeryk0rwSJjof
0SMCNw4SFVnoz54abGtcp7PANipvNaFGORrMhSuSxDexwwATYlfJyAp5BLcVd1YvJp1kNcMBCQlh
cIzBtb6IYvRgqo77mTmyWAMmY8eS/C/4JbZvJImy3Ex/tRV8w/ntAfqjXCOv9eLVrjSKVUEfR2b2
I7g9sdpYr/q6oC2gy6QLzT/RFVx/tAPmueFJCex63XTae0yX1YAgAKnJl3JjGZ8paj8jQlLuJ2jt
HXVcVxQrlbc4d6TUt9N/lRBe2q4DIZjUYe/b+Z655zHZaecd94RmBIXdUN8fek7qr2qwRCmHFH6L
GisyeTZy+710k5IwounOsPZexQ8mg/yOIoIF6OA1NC3w5lKpQhAVqHtPEbcHR1FvsbLbSRGZU2aV
CoqrpqKYGrflTuFoFdNEdU23W1oPjSA2vm+nqWHBG7aeZ/UCudnJjsOWfvQHBKF/nXVUizMJ9D/B
nGFIhvNrtqneKlmvAEjFKkJz5HtilTGoqf9GeFvAmZMYbzXBR2baQmf5Q74LxYQLlb+AWr7xYKh4
DBaHO+n6quT8whtd5ByWvb8ptO5nbsgWAtVdX3qsI3QDt65VF4Re6EkCAlEwy7qqIFiuyfXGvggs
pD3ke4hejMrd45DCRm8Lhj+3XkMgYjdiENYcmUylOo5RZe8LDrUKJnAU+dCm3JBlCQT+BE2xxors
4yOOPtrZUY6oaxDErb4FXIGypvl/BADhPbdf4twR/xg3BUGKOALk8aqErg+Q1jvgbEShKc8wEPDo
8YAGFO3Z/bwXJl7VcSX9OKNOfDgjCuwLyaNQztueNgyQ9Pe+Cy0qRULRynw3W5yQDe0jDfkvSJLE
ijp3y6zkILusqNvYKvVaWd845YW/i4/MWdywHMM89APw4KqlFWu+YMWlRYYB901NRsmBmR5LB7z0
W+o0vZaNRoiCYZrOzCsnTJH1jBTfrEPv61jw7F4Bk2r2W02I6e54lk6Vf1rUGTHYIVL6T1UvKG7U
6s2q9zWHvEWRO57JBikiZQFVkh+DNRTQViwLha9TwoEGYWNYn4jNOMU364cn6utWp6sucv5gZwBk
8nEA22G8GZRknvxw4o1EV+RpjPB9Qz+ZhTaYNW4U7k/dFUK6cNCUI+i3G7qyFG8cUn1X7k7d6gP7
cEwtVpA5Iezi6Bln+sjDC0cBvFLoxQqabo1EO9hbJE2iIjCiXLR2TxSmavH5HUymZ3PeYEDHLdNb
DNibRP1P9E1F8bzIiF9u/yNb/c14OGn5gixOXqqsT+y6PhPev+D2x4uje9mMu6OHKSdb6QIg04U0
YQH8SfM2+6K/JbfXGr5gHscGEMNCXJDThSoEuXW+5uhppZTF3iTyiXd7psx3EQbelYuY+U+qYq0W
F4qHPofZv6go5g+WOgBQJXAl184lk7/jYtRfe9sp2K87coYvyH++Ia6XeBad7aiW3K7694JtM2GJ
ea6PImWlIqBHhR622XgaX2cFUCXdqgrxhvGI8CbYhRkBn11mSPhInBCnNxve52Q7oE1ax05MVxCN
Eiob8qQM+5Rb8cCEzy159C8jgS/Fr9Ax8cyTOkYwIBmIrrMpFz/kgwxSmhz2Z7zBuhtzO6U/fOxT
q2xKM2S0cpoDGsgyOAHU5Ml6GCnjU7kAGymu93e2v3CbMzBlArl/bt6+u7wNXFgIQhXAMXMmiY+c
cVpWcAzXunjITyi9Gwh7kwlPUvqGj5ksDkpznfS5F8HB+6fAF2zebpiIPrV3J+Z7GYtLHGAzMNvX
yspf2CmSWrnb2B9LLTve9m12H0mgcd/qihUrGTemAEQKzw/dKZbHD4nejRDQ3ddurGfHiovMPC9h
6cVeNiS72lpjxPG000ee5CawFTZvvvANM+GtffvYaceHm5tcGhqfE1b+Q4B+/UJKT04mh/dNdK+L
bkeFGUQJGOroCsA6YW+oYgrsbqPV3ZMRxc3rfmxwUFCkNLzbeSGsMST7jtM/J6mTiXAwndvNul4h
G6A/FD4N4aSS8k3kjGsw4nkH5oOJemXbkrYqy6sI8bJVcM+kObE6JHwtF6ZAjaCz9IRybiRTHXdX
1xMYaFdEoUw/jaeE+NnJkQzq1tKMlGy8uKFXcHNMy/FvRpdAgoOvQMIK8OveokOIADt1KQSrvSez
cusFfloSjKSe2UDdEP31s9MIRt9d6RuQK8QkbQGk++wC5RjwP7P0R7xK3NbAnSu9OOk2XobJqC0K
YKorp9MxcCw8B1TslpUbLw4oOMqZOK27/1EU4wTrr3MPF1WVHaT+z1sTz2gd5QCexZZ1fLV6LhA8
uTykmrmHz+ACpllTo9694cMyhMG9NZObdZeC/fG7Juxuy1BSCLHYOoj23+3tjALdJXxb6V19S1xe
xkcVUZohL7s71/Mh1UdC9Wd1ZSc0Pmhg/SMOM8EG7Bta1hIWjDK+7eVS2kQ1rwfmsKqoR72zhs4G
EeTTIIIAx9LIQuFBArEOgDo80JgMBEJ2faRm28XPaSsGTkRPdWpXZBln38EiwQCKoE87Uxkpdxci
zJ0Xg0wExa5LpO2V0+sSm9aZK6HiUR0La4SbkTCiLYlFjxCOJf8Dd3FK1hu0k3S5o/cxZpcGf+IG
Vo1xQ5ClxEtrf2wJ0upO2xa0WAxQBYdZGXTFlCGybTJ7p1jot5x/fk35jD/ztsRHjAkWL2rsUP6N
5Vl4EUUzYwxYu+Hl7Aw9DueWYYWS17dJSqyv9tlb1qo1JHlNwypy6aPTdSdtYk3MNcVq+/Gkj4yQ
pXPbN769GHh1BKVuQPSLU1RlbHOSuauQpHq6TTvVc5Cr4gJWMY0VZVR6xe1u/YLHshnB8gXRU94h
MKXXOgyk3rtIz5Z+QH9INBfiK4myhY/2lvry2M2urzCeKu7rMapq0Pa5jpqKk4NSj8RjZ/TE3bX1
ws0gl8Jt17l18R4CEBtYhAAozUQvcPN0uCQtpMKSHdsCUNCG2I2hwP26ckhBU2sEdMrrSK39KxFP
g7EJv0U/L3kH3DLNzSxXgw3oKmCHDLP5D+vdaVF6FMZkVVnJF+emtFOQZt5Z3+1pe3ZKh5Da63Ws
LZP40iNEph3INCC5iwg293c04ygnaGuiSEA4DRpzqi+afAeV/rwGeEMXzp0qIkxaMBbNmSd6hqVB
YtPyCVEI7mzIu3nTQhjeX+SDiqMztcyINPWDqYRlpoYLjgWfWW7PvV0CQKkwwo6W6VrhmeBAOzhv
bCgSXKCmJa3uPg1BsbIwX0HNeWDF55psYJyAkJ3eSGchWxXdUnJZNYzTmwGfINr9ytW9LPM2w49q
hPpcgTvOH7i0Rkd4iKnQPELg9tOEKfgYzaCSVZWzzvHkb+xEYv2bQpJoN9HzYrKbNhmNb6J+7OnA
f/k3P/nEdInFehOomBHQtzy/CmNLkAM/UUJfxw+kKL5jdh1tyW0mj5Ef1DECL4YdaoFMmTePqYDE
iJf1VRNdWFWuMqjWLJOriQ1MW02scGdUemZVAbnKqDgJSlTSyA76Rxr9lJQuc+8Qjq9dojQWjYsz
dDFr2X4CYJ7FAhaucGBhfEtXudynkpK8f4hrcmGVvaZIANavbVJib+ESTJCCqGSZyDHuE0K7dGLQ
hphpLhkbBO8KP93b1tIHiMr7HkCDUBBqamjfrYF3Rce6TSL58B5Gqsez3PvebeBD7GppRv7CqiNY
H9IH0M3Nk4PctQRRaYI7EQ/FaYH3jSxtIIQ+FJap8Sx8Q6a4NMaFSVJ0gBgLGVvtqjeFGR5/QIy5
i6ibomrnDwOfe/20vnE5tA8md062cbsQ2LzUUXkbvSv0XGPg8n0f5+hwXdZ4exhQLBNtj0TS/HxV
pDYLqMPZhhseaQCbtz3gyfuvNtUO6ijJICXTOaTMpM52eWyvg3k4GbYC6JpV03BL6an0b0uJhXKi
ydCPPPDmVqXF1wgjk+DErru+Jj5UgnjcSiyd54N72vXugIX3mMv2spsEzRa+/qFMDKd5PhbRkWtA
8AxKnlGRIyA+dJPH3dFgbCR3JIUYOZBxbJ2TbD3H/i1EQ+yGoUArtl47QVLHv4k9GNXSrZ59WAm5
mym3sNmIOA0DoTiypUdOypPuHUFYfcx0bWKJ9CsVZchuar/Ds6cu9CEu3P5nXBBLMKKGe5TZDIcP
mOOhFve5q7BJ2L7cVV5AqNSWzgAPxzWER8ynEATEIjJKXcOHtLwGxrKKs7B+MlSW8mRhfQ/hJ3M8
ovqmIaHSvSN48zfAkzfDhowlyNselLklS8FI/FRNhRaadqDsrCrLur8obh/3ls0EwQLOlavq81bE
Us3gTFKHtjshXUdJrbtKqNaR2NicXA7goEa2qjAR9SoCyiHD4yV9PqDy6/PJcwm72H0QyPxVOQm8
p8EYKMoh+cA6f/7fZ/zcCJJvFaFjbmEkIUuVGr1CBz8g0xpvtrdeZsD1AouV8+scg78yOeEsomLT
lYlbrr03VmaeeKRJyv7lHKUcPvyKYwKaR8GQkv06zJCgrqphTd8ds74N76YWwOYhVd80ToU+4JRg
rIkCdhz/X2o77YYExEMgm4FprwGW7SVGwYYJiNAQBwTSAhUVUFynOQ2jcz9i2fW2RDqpl8z+rZkq
CtwrqOTzE9voz6Gl9XJxkug0tRp9qYR2hhj6i1h6oe4DnkRsjIDiYSqQcIAFaZGhf23Z+bF5O/bt
0lQUeSXE6XtWyNPvuzFjDg3eHSSBB3cLAyy7QoQ0b2Th7v1xCfUaxteQKA/IxPWyHT41sh55JtYe
CIY6qPlivtin+IYCXtczRxW4CnBogS0TjknKKby25hur9lBZYHMi0eaATIhVCt+h/x+5ul0nc6Rg
W/ryjI+tBwOfPSCUyEyO2R94vfgjKL94/hes7DpGhLMtB7Wa516C4V6O6PbbpWu+jixnSkQ86Og4
C+x5X7v7VzxoKhFlYDnHmC5Gfzx3uPN8+00jH9AXEgzpGiGFkJcH0b93AgORnxfdQEykdXOYttXS
g4iylw2MP8tqx35RYATw/6vHcMh4ZeWvgPGgHhrBEWEiCHaV77gfP3/Wj0ISBZnBr7xMEf5a1ig5
Vw5rMfUyFxGO/bOIBDHBqQvUqmtfAXHM00UYBp50rcJdO4kC+XnRpFnQvxiyPTsIrsPyozgzr3hg
P/u/V49/8GwMd38vcnyhGJFoUWlyr/emURIAR1qiS76VnesOdbwS4DwT564bHn/tYX78FYS7lw1m
qmWm0FlYceQHqPl8Xg05iL2hsMc1s6eryZN9PC7hzOdSrraZVfuvdbyDMuxQgMABKcJCrRb31t0z
cirifMKVWk/vbPOq0d0qgTs5Myq7U6jJm7wiR38b5L8yWK1PTIihErJDHBvnb3uKHEk8ubq/2VEM
AptXzCUTRTtL0PwWeyq/vqVm+OIQGfSthJZ2knKCwpQWOPzjkhZGPWZ23S0RnndbOKlv+1s3YRPm
FqFDR3kX2mttFtMzkWXBLLrMIRDCi8I74l2Xi6zQo+IgUQgNODL6cZZxViNh8fSEdR8uCbTGN1YB
tahdDWJrjr6MO4KO074puQXErVYpyc0QClqkElds+8Y/b80yFQKwSgft8aSAaoaIdyRJryZn2Cbf
xOKkvtlTFE1g1IsPjSOuE62XncdjFkxIQuzpCi2qx6gfuuNCzXw7XqjDIONNhTgyLKeU0lfnDfHB
gY4vCeeLrTVIwBcQjeUoJPIdcujBfDxJ+wpu+iJEC9jGnWiJuSMBHY5ZjDTEus5p7RnZnvkRpQSj
SRXevCgb0AlXweIL9fL+RicRNJmDF9IAWNTsLWEbQfs+HGS2LcuFx+lFxD+5Et84s+03ptdXz0a9
MKDPqS1vOT2ZdRTI5zixzi7V+lEAM4nFbMZ29m9zhzV+Az1IE8eouEUT/2KD+V63wS4T4WOSnX0s
vVG5hw6ghpCcR5hAW80Ip7k7sujVA0XBQI8INqY8By/LhUdri0u+omQ44NSLMcxP8tIZ6P7+c8h2
hHLdCjYCQeacl+LuuJMj6asY0qBMYGAjszCde+USkkqmlm3YFsFP76l0z5Ap8uj4zlMl8SABG79e
guWUe1DvT514r9ogGtgtvMpTU4E7M6ljGGF1fifBaB19KuFhVnP8CI3kyeXvPHJ12IPyTUL5hc8j
vauZtdGuBQWbHezoUMjUlrnqXcih3pjswutR2V7CpN+fH45S0/zKSuMqhKq//drcsmPKFEG3r+3e
66nVFA+6gHZtxl4vJZBdMZ/OQ/rrxRw/+jWi7yn0+/yr7rynjypYAf/n0Ra/vW4lpv5/EuYsfDYZ
eXelskbO3nH90/J90ZT4AZBQt9xgyL6lDnQiLErKXx93w9Au6wLT3gbbwFHrRvat57+DlYpVvyQ/
rw2Hrnb/lISe/O7ugjNUJk6mOYGNw0DbVDYvAHG4lE1FOx2TvH1dqMzOLs9j7I9uiCbEIovL7Krr
WqazBuP6xh/CwI0HFVzwsl6kZG+hVf05xqFtwAKNayiRIXN45bnLrxj69CBDDW0vREEbQKKydybb
nzsEJYzuLx9LOCaq/qyYAPRhu9WjySrP9yYrxltIJ8wsYu2OETWIrwjb/mD2wY+BTfkSRj5TOOK4
i/MFHPtJ0K6hFxA6MC9YUwoaMSLpTkvDxWmWojdOApJRvXcyw/N4rjtAFl1BfDoAKcAuPDildkxo
Fyi65L/tDzamb2SJZM3Yhf0SF+UiAqwRVmCXQDxDAznCM1VNwhjRfMHdgfGgjqa1+WEImRm27XNF
fa3fMJtiNLYIjTGfISp53URIGVZVGl6iiqPznfhAvYcng4msbyjrUz7Ggj9xWCKFsf+fvg4iJe2g
s3pIEOq0l746vhEXVO/f/wcuOBkdVsS5CC4so31/P/ZlIfUoRL+9KAnf2DoRYlAIYsfX9Gr9Z0M/
d/3L8XaNVhC6gtAtfSgYXRinZuJDEK+ePeJKWA1vmjdfZ5H8rJycB3xZx+MPWRuGvvgTulxXeE64
KYnfBQGu11qViBjGiPzWNjjTHEp837p6l8BaGB1yZ0hvbshfFxREOgEd/dCYtCYtYnUKHS7FKvuE
pWNdHI7O3z2e4HSf2vW7U8/gSXVfCRzyTbxLX6LDA099iQAyF58IebVu+IU+j2Nj4A3t+gCdanZ/
yp1YK3bQ06m/gEDTw1AE32oLe+Su1IBGGt7GbI7d2XSE+AjFPkdy1LyHHgsfWvz9ii1c9L8WrqGU
fDmcLFN2YlOaO3WgIHQ48G2/gaMcByT6N4wiNpcDHaHRTa8ch07Xw60V0JaKfNQocX+moC+DpfpZ
tc5m6otckCn+27ORIco+OIDT4UVSEWstXCAnUWmkka3sxN0X6tnYWcaQ4C7f65VWDTIapLmFlBIo
ofWSnwRC0q4Ku4VawtmJEaiOr/GQm10tR4de84/lLb1GkEF9ctpiXDURGDWZshqF8abDXinDB0rK
z/FkTTOAymEDK2DfmCI9qjmvXGHXz2Pi+9d4lN77YhwSv7FUD5gNBmYmngJ6zxj1uZZu7dhcskkP
VbHZN/mtPbUlzU4D+L/Jt8g64bsR6A/ndQj4dIgLbRTi2snwTB5Xn4r7a6al5cAFQeBsSMnDu7lZ
PZACkRlX4d4y0HRimotCABxbSB679Ep2xS2AhZ8gE8uxukSV9EgqXqa3NzbG3GkXDCsIMd/cTCa2
j3ZAa/dOFlLRL8tVueEPtX7q6YRD+q+VusLAu9/hVYKymEmTI3BdTbNbd2vrjIplkBhwAVQh0Rjl
jfaXFXZtiqQP8s2VfsfzCtJNYA9PRTyDjix/6p9VZ1V5yf6DEJTtBEf32ZvT40W3/x8NpLjESje8
EzMi8KDHyNtqZMJsTNvLUn0RoquaeAAnznIhxwaSgVRqSd+jAhJCduWN8Ei4IzGvucUG20FMKCP/
u7ax5FSpYY8Fxbved0xc4R0GrC/ZmHpoBCPuKbhQWVwQ79tiAABaZmeBMk3V1rFsg/OsicYKmvDG
qKqGp692y0It5mDJZAam9eogMw/7bXZZ31tDIR23WrnEqG3zchalXtvdKQUUvIPpCp1plm3WDOCn
sx9cghLCtF8CYdxnM6QruQkfpCgBAuntI8jAgTxi7qfSK0I8J3nEYg+obRxmVRkScd/vwCOL1RN0
CyB/qYizWV/7e9/rJojfZhxCGoo3GjCn0v4pLXrudegEU4einehW7tRDUxjvrDCZfz3cPtodFxde
+DCWQayKaHpr2841xp1sijInIqxPzFLgouZ6xum7wfsHELM2ngMbHz0mPnzVV30Z7CjStsvHVL9A
H+RF/HFkY8NZHdGZnszUfj5pSiMN1bcz1dYMmeaxuliPDb/c4QPeKkIEcj/KILjo8ffYNusQblsH
8rvx55oYMQR2SfJewj+GlZXiRlsGmY8dTNv06i+qM4/Z3AyA6BuSKtospHCwEgrKGFdlAtirm52h
L7EFEtfHTsmL60bPb2cvOOCNs2j+fckx4l1BU5kQHMAUyZUzOsOHOagagNuCSF16KrrwgfXMFbWm
cO8DmFpQjw1M+x5c2uSt+WGwbsT4shz+Wj76ZYKVgSIXoHrKiX9pLeqdKgGNyOHUqotQQME0dj9k
yrBCzAYVFQ5z8lfYkGWVw8qd6xxqo46IktKA0fXCQsIRS0X8U7ltiRmHAm1YQLzLlbeWWVG1ghgk
h2XvDpNV+mg+NWLYiyswBF2CNS6LoD9+R9P9E/ekjyTIZiCQgPaSrFW2Nxaq8L4S46+HfV6xcQiN
0yIzoEFt7RdawhRWWMw+cMPTl5ZzAMKZDcZdtzuEf5kG9sBQpsJV1k/iSSi8M+CJcNkQ7IaoAhaO
bbWfY/rp3dONbP6GqKhm4LpBlLp0a+iIfmvzkzjM8l7DK66vCaWR3Ji3g4CKYAklf9YfD0lVtzEP
3+YsDaAaNSiFFiVuZtldQmY81EA8TaY+MfSi3tYYJ33lK2mmrJ9htnGVwGVgdCEB35lraWx6NlQi
jmkC49JkJSpgsXB4Nm8NzFcoWo7cSp1PsQ71s4n1PTyKwC37kUdL1Zx9gMF+WaVSXltyV/CWWapk
C8HUGqA5vO9KX6LF9HuOp0a8RZwtw4EWzWrmmUmxeTHwX7FkyTF3OE3G409k0Ta5XOcYdOuv2n5o
VdMNqBUiLqOJhAnvle4hrAr5t8MO54aGXfmT8CPC9n2rfD8OSc82TvrQFBc1oxNaSPwEhumH9J5c
ULfhKuoRVuv0OgnWGd6tVQ1bOXoZOg7vUBcSBknOJycZSi4RIhIlAwLZjONN2tH+9wAJos109chw
x6jJ7ycG4AGIH/AXzCR8/kmy0Zpw6RW3/ZpDLk+XdFlxrydb+u/bbP8BjlhSazg19mqhNJApslJh
C1LOALaScadf1CUfv03TVR0bpkbbaF0JaWRbdvS1EOL5mnpHBVSQZXVnhnLWLHJ9mJry1w4qZkvz
5l3gMoRsYj8tKc2yh+qZjskv9sh8c6SiPdVif0nAxhYCfx+x0aZNikCM/0KyDz7ZVUzHvVs8C4Ag
i61gibcv4m1DgkctAdhRPk3VAASwpv2qvFhTugkFTnV3EVRbaXFc/OzkM+T6VNJw/QBQ2j58fgcv
i2SF2P0xz44RNhVsrNfnALOZta0jUmfkaHcjbaLD5e2torK52Euo9fNUM7xaf7s31inu4YQkU5bc
47Z2LG0Jq+eKoXhoq1Geonj58HFnQorgMS+8GZIKnM+WIAha+QhRIrBiTt4zxqQGoHnGVDyeB311
R3Ca8BX1m5itZrofRYZpWlSK83cKcZ+9MUOZUveslENHIxMI7prkzub/HyxjZYqlxV04PItecGU/
6N0T1b9zA7Lcy+zLLuHp7GP8FdYpMD1xIgz5mkRrZq1r3YV/+rvrRskwYW20Qkk5WB6MyNLhQWj0
6OssvGaz+9QIc1v4JIiRA9RJqKejfvcjRR0y9ug0qf5YCNv9Qb31b2oN027vYqEa0zW/I3hcOwUz
zX0dj5mDfgzs4M+cZ7Fic1UgD5zfUcn9lHKQokaMKBkSJvw2SHsAKwcQza57wipXpEFqR9kEuR+y
l5G4h9D/TlORNtmeuKGKnG8nyybl2rYFeTe800wNHRkDxlvQTtoHMX69ocsRP4FEVPL/vih+i2WQ
M/3KbdhONQR0/RDQV1WcBaHtk6s3o9CjT0IlGIs+TcYiTuYWVZ1krkVK1VTB1PVEUWgASF4upyaF
Rm7chn16iWEjfY0QjGiQe+zDW3b/aCnY6H9ExJ1iR5kTVnA/H5lMzrXyOapicocofGm54fsuuxi+
rMxUJU0jMsnPhAJQAAQisVDLWiIVdPD/hBt2CAMgmBMk0T3pXcJMhvuPfTr0c7FO+n0uyXRJbjyL
3u5YLrSCv0d1LQ5oPzt3H8cOOwhMIJRSicthPPjTiS3tR86wuQvjutjLGsWkZJPQkzucZhRoqn/R
TJKLwBufuQLYoar9LXbe12m+AV2SwsQTwTxHorK1RKCUStOhAUJRoMALfPpwRaNQ8LSD3hHWg3ij
96rphvHwa5lbEAeqjIlVvsfKV+7ZWQ1iMrJAJud77iTW/HLGRfmH2N2ROttgeLvWWmktQ0DIxObc
9ft7UAa+iXYvbXh6t3/5XKqruzreeug1GhiA8MtEAJoz7NXNtHeuBsh1iq4BU6rTzHUQ4kzwNtxN
CIg78xPjANQpAeDdh7IfLxGhM9zCrWFbLIf+M4/6TWh2a8nLbtx+25L1pZqHtK/rW2IFYOk07xJA
lDW9Hq6vJSCfV6IJLba6BUYcbH9ufiXz0HcEeBmAycMON7uGz0n1A7wsnZmCsBh12zYmApXU7aLN
GtQl6CciGdmgT+X2cCRjKDtFtoYeMM77ya9h04Lsq/MKCB/QYAp3nAVH1doikEpZ8kwI90dWFIs/
P9nZcEryLrTEl1Tkg7rIFa/SIxWdTw9xcmnjI23MVbyGRlsA7o5+cP0/rdi9118eeX50uKrVdeca
o94QCxUPYSAOKXfdvs+xomXwfjKqblb5zkkEPgdF5qD5LbaLTHjUXfQVB8EoSQWiLW2LfqHsDXBJ
VbdIZ5iRHZRoYdv5EuMqOaHu8d8amr6A2v/dpK+c40MnXwRVq61j0lxUkBlqkhBKw6YKuFBga7Iw
f1NkxHuhLIc1WuwxUKnUH+6xmkHbUTzrtZiXWI2DBIekFup1DwYuHzCvTbyZ8vzLVpfBCI42nsK4
bt6Kmdwfu0pR4ZP0d602kheO3RmGeYIPISp9Ykfo7glJOXIYNpCnuPtfQ/1QmYzoOzEsV1ilG501
ZdC7qnPt8kEx44SDmhwqm/4BRYBN6B+p3wbbTruxNKhPYtFYeZMKH03L1CUWwdqiAOrsYZUavYxL
VvlviXDGrB0f+a6XSGdEU4VLOsSxwjnxAw3jIOSRibMMQ1NCibAdLCg1C7aWRaS22vQZrfJG4Apt
6AqZEkFrGjyvR6r9NZ8ndjoTxC0lzjiSL6ZuCI96zzfR6EYYW/c6chxqxJ7SLnvgdgov2cMuc8QJ
VH9LWfi6dU/qHC1/vsKLkF//owk9osdtI6jES6XjxYiDyU+sGPpI+yaMTTNDA3buv5fwUnmkRkRw
IkqyPvPw3V8JS85kaHXNRlN0VAjbtcfoKG9C50rqL6xMoxTJgeTdnA2SMHTa0xLr2luHUupcvtEM
OtS2KDSXRC+bQWHdecFbg+GiSJx6iXPMB7Wmof/UmZC4ZDnBxMC+jI5JMHVIqj+ZZwignB4nmUG8
xIEgHs+X6HOousy3bXrKBh6BeNxtWkPFtNq0sXCKqBKZpxGRuyYliZrpJzTX7OvPvXrLaNc8rcrp
BkYH0TB0fzKGRnHTv7Ssd34JfH86a67zGchJb7vYzOfLkR33z8M/WN82vqRbFOQFw5HQhsOtfpn6
HmvJNLZt/64dO2P2yC6cgNo8zsD0F6EQ7K0UxKKSlPQA3I36ffOJSJMUsz0LN1oBZF8Fm1qI6TZ5
pXCibGCbUdvq8DRaYuOB2S2O2lTIxr+xRx1YtEmRMBESejb5q1aF8xnuzfaOskeUIEIIsfdd56OY
n1+FNifioJoOV0oaPPsDiIA70dokQNKJP1KqdNWEOdSlpYu45d2hOtJ7uIOrRJTzGWvsMiSpXa17
4MS1sSB5KNLJELO1GtbCpq/4CNVL/qVXOowSHliUJXrLhrQKDtT22fSXud8eYxKVk1Zl/ZgAYdag
/4W1rEiy6fTiFCZW6GNLcGDS7/roAGGs2jIotRXCCB8M1LWnzo8yQIYFfflLlytNpv4z6jvhSlaQ
7G5Y5bTTcoa6fvNW0LDvyiMabq5ldyzW2SevvnZQLu9bIsYEgcQ3pdeiGPczCTonvtadiEiuGS2Q
M06ImOhuMJHESZNSTYnE03a7QTocaEU9rwVN6j/4R8V/EWSG9R5wLenMHCUjDLITkyZ3VsREGC9x
85JrBjRmwN9dHJ9xxwN7UktOkH+TBEu+3hU0k2ui0/TmHlo56ACAHWXsnofDFOrNm/yhAcDaTmqo
pTxEvgS6AsLNnKeQKzetBFqdoQjXbCW3H4vkYd1sXzdkmJcjaryH2eC3jgwRy6KUTCWfDx744CJ6
A1gqhdvDF3n0agssRLirK2UtcpyOJkwn4vLmqV3wqpEXD3kEtQJ4/FEITqyZrpBHCdSlZrqNnYj3
f06EMPwwiLA4lrqSB2SbQ5DztTF2ZfyJY/AMy7CM9pu3jsvIQOc1fhJcbP9sFvcu/3E6sKZiuewk
kK1F0EOM1iufVdKqvd1Hk8QStdIbgGTjQGEQnqS+ucKsBwJqFPy0YuSOgZo0pcz3Vr6cg3O0ujrY
+4i6h/GRVStSn3RU1rkXSiSfVV7HNtI4f6GqvXJdlFjzlJTlE1Q/vvCCqECOZVDMN5hirxZxSHcJ
/M6cTNH54vq1wMD+j6ckmN1Uv3ZUSduUclV/hT5m1Bu4ZCW2+bFk8c24RWqPy7E7Cvdn9aO9SB+e
TOmW6DuOoEGX58P+5AJ1pHwGDHH6A7YPG7ElCt3yZ69pfT2BuE2XY0wYNM04QQRZM5IfC5kMLV4E
dPs5NoKoC2n0G5U3cq39DqXAh71vP72GrAMIkSwGPy3akxmdJ+Hn2huzigqUwelLt/dL1ZiydPmz
nWl5Wl1MxqLwIQHTJm5TVvFIao+vhk6BiV2XTQurd/sCzDm39ICZBrfvrha8E7dzXPgyqUKUwvTl
Jj/VzZRYFJ7MSDYqkTOuHfBtve2kyJey8zIqOjKXmGSxW6xg/SgimAqZCQCb1jTnzrJzR4UFgLVK
t+sVPaUvUqj3SQxQRXLpwQ9SKLPadYz4JeE9/IgueYgevSEO5IjIihRUC2s+HJ3Q7VnCF+SwQtIU
VW12FWgXFaS5iIlyufYuzlfdOIvCw9w+KVmUvl20HOvNhJQFyLRF8LM64MCGDl2Mr2PCbD+WXk+A
13NYWssYvTDEIKwT2wSWcAEAIBe+h2kzaAS1RVqLE/ii26px5TpIUHCSWLjBjavcKZklmU1FZAxH
S9+JnonLJZLTg+Lp/pLQeyWMURSanHbQJ1Ptj/i3bluz9A14ZkU7JPLHJEvm7Il4fb0RjpXCoDpX
/mKzMxoldsUlsQVfLVnlR3aSL7J078LJveVp8E5JZrgY7VXbJqjQQebY3w6TIJ1NiR6RT+1txu08
RYYb9/ZPZBdrHkRkYVw9yGm75tCTu3TzPqltLeacTRqkn7DRr1apXoSeoce0eonXqhsR8SfEBXAS
AEp0S/EPuZdgMw5le/LFV9BfoodkM7ypnHWQ+mvicQoztU849WHn43Y+PmQLe8i9rEkDjLRcV8y7
i02JI4yi2lVXzZ+kGx4BCUMJXtt0Vp1o5JadLg1o0a6gdWcVIv121PVOrdEBA3Qbyotw63RHKCPX
3ZXplVQLA0VEsYi4/A0juMs0P4Tp6UysVSutf6IxV3ZGiW0NF0tUT1m55YK46qjQC7TfH98BCon9
0YEkXrh8qOYZ0+qlANmKMaouyWFakHo+g8aF47wrUC8Pejx8bMbfBgkboBswRXd1JgBSlfy9nbY/
UPB4FotC4V3yUO4hdf/1dV61UWLRVPE8j7/PeTLOFqSyW+qYutM+eNGJ7GrA4klpPefuW6ln15uR
kdprCBMA5ueqg6Oc+qeorv1PLBXbYuyhrIFZQQ7HW0kdM1NVmEHuy69+a0zaD5h6u60zT/e0z9Po
CLHR3pW7LPG2IObpotA83wqCoN7trR8Hgw6PXxyaiucX5ox0Rppk4+l+iA/pBa8ytVKqKsxLTz12
gATMXwzSGghjBb3/JslAYvOOOGFRG9L2+2LiIkGenN+YHJeWBcpAKN4MTtYkVcwORwEHchXrAVGA
0JREQloGb8OsL0QD9i8xyUQEMAMpp6F93nmV3jDHBpSwRVdiXpscBVwih7cRmhRPItV4/pijLTKG
aulMBCr2xKwqKZaMBrF3aFmM1I3toJnS+FDcxlIjsE8CttTvW6Oty02uqm8pFoiU3rldPFAcXFBL
n1INWgOj52w4lCfmkp/xz4pzUM/yLTUxlowy+PcFuu3XqCAwhRVRU0hHMq+Ght9Wq4xdzMmNRCqy
ocWP4epmE4dqiO0E7r/rQNvlg0dyAo4pywtf1cMN+F6uyviwX/sXy1lCEDDyKpn9nUUMb/uilpC1
VxQ/Iq33rw8vTlPUAGUIWCHG2icPjIN5ezV9fIsGIv+SyA1cFpB4w++82EWOklvCRinak2IwG3+D
RmrngSd9MgYS0mGwHKUI32H83C0JXpMyksuYHypbxI7Ioor9u9Uq/rb36lBdyt69KwW5c798qcsF
+V73W8iGD4iACgBHdGL1pLTk6+2pWx34Cp97Oc2rEgZiAf7rTRwAqLu30KGBwcEfLc27/CHIINMe
azpMVDAURXR2DLa7+ybQXHwhd7jKjQEUR9YqYAeVGmTR7N86lrrRDyES61JIxZvjPp/RShCWIMaY
muyq5EpE7/32vT8+6GHozzeD0YlPvC/sbNdFMLMZu8lgZ/xoIoIqC/6rV+dsQn63V7/CY90yjH0C
4idWGnkIa8gW6OPYgIA2XW/76fw/pHRCNi36ZysOrU8NVEMI3iBBn4RusAyEiCuxUZ7B/mOFzU2x
n8ZdkjOUs7XUStRsTo5YaBtOeyzlVY6yGYjRJ8+OJQsVyyuUlbL9ivXANfjiJvtSUW5DiNhDjfJk
uXpHc+8I5rC54qmmt4zQyovSSRLhyrE/bBpPpUjHPAjO7NUa+O8tX8ig3kM2jGRL9B8fnvra9e1V
xMdrjDzN6oRhn4y61SJGcoLWa2SWqSnoq2mfgTDuh604CWvJ8i5hPpaw3lSagBX1lNEv4vDI4W94
m/PWAjhdc7V7XAqMxZVuy4nAqX60Mizy6Mn+Bv0l6MF47WR4qtNmy/PinXeQb3dRKVZtqR9zSdL8
9PYIlXPpAmURtoMQilWacKpNQpu5y+MqyyFhTLOWABKde3GypHeF/gGICF4sRogx4KHT5i8TTgnm
KboxOZxzrF2sorH+mR5Q8nUwvDEGcllyki7+JpyDHf9zfiXyCl41vU8tGMICa8GSyp/CBdzW1pJB
AkY1QwrZxKwrClH9WdStSnO6hMQq13Ot2MxGVq7O/ME3NaszbuBMQKPYbu6UY8EMsWoHtGEmJLGr
RQ/yyQmWdgo9YeooPYQ0nNUxYVDhBquxgcxNg0NBiIerOd7D+a7rxCCKsdfIHrmZATzyFGiOz3BJ
FDz3SSjq7tvL8W1RyyMubOWY/p/gDW43AjJ4ZSqqBIACRh/Tu6bVUYJGolEMWpZ3qfhYTpSZnb8o
qYmXu/sRA+mto0vNPrUl91ECq54pH/KULRizN6CMo8V0BdGBsU7r14/CujrN+d9be0uBE2W6Bs3E
D3Q65Kg21WtUSv5F6EoFVOSvoj8Q5bBF/z1T2LU6iu/6xj2UZYaTo19OLwpzS1FgDkcPkyS+QnnZ
2LwlPE0sjzKmt0xBLVU2EK2yiGXn1HJGHVvr0zGNjydZHxgLfjLtypK2wJXzHdy6PXiiuuCTnt1C
pswG2KEpaaV9ASnWAyo0f0PDsHyLa9eE7Hq7ED8hW3Fl0fHgQNkqBcwGxdHxjL9ETGzGbZlpQEKg
4T7WKbKN8k1dl1lPh1SjNIL8+aRpgUOiRvcF22dD1EXn2BUMzIfUYa5uXDSjwlVJEpa0QiOYBLIL
v40jx1Q9DBoRQ/azMErHh+tYdIhc4kp5FkgYLbQgLW/hUVcsEGFrHPfdw/nPdbiwJ8xlbgps9Ht1
s5zi+lXZAheFroHgKQifXlxxDkRrccv9bcw2CC+cBSV9QTO84S6ccrzfxiaJtuv57Sc/UWlA3/9o
sTXhxp/Ho7/QHpD+Kdt9T6u3Hmj/rvQzeNcZB2o4v7GBcFYTa1pi7F9E+zmNjBmzZaXtTqNFtec/
QdcM5A5BBy4TKK9Ho1jc7U4mUANQWY9WGMC+ziefT6NbAFtxer8jOTZwP1tWKy8O0AvsQ8C8Rjni
r2PlPeBtTaXOR6WgoxwVqHMryLyM9yEGdtFTFNDD69n3pOcgqo3ukUAJlPsBPe2ttGF6HT47F6sq
2vktbE0CJEXXtfOgOpt+7q9I7ME4ql4gKtL1Hty8MhyyOACNiV/pFXDptV8p2i6tQiAAa0NnQreO
Ue1bPm5ZN/L9ZSPdeLtZorbrvHYdkfH5EzjOQk43Q33ii0lLyXKSsqCivjcDY4aeJJYGX1J5wQTY
yAk1qi+fAi5l2Eu/w9BIGgU3amNqQv8FageGSlx8QAldzYsAjQ7EjCuFq7ZSWHZCObxdGTjhxvbL
XZG0EmIHgCY+Oa2n14Jmdi/L4XPDesjDHMvcF+VhDXMmGR41BR78NCsMi4KAxf5+0J5yLY7uK0By
7T7YNdJLGzQyfzeNvFpbknSeV6fCeMz6vLX4wRYzEQRmeT4V0451LdeevDRH43FcAK+67CKOTVMh
5UY3GwUBtfHab9oaZPcdu7hMc9FeTxaVTf+SOmMFHg+x92zBjUtPTzbbs+ZiiIj+mDhW8SbAmWaU
UkNpZfgachI6LsfywevFqs34P3AMq9wygbVlyua1kwELTKLy/gwvQQgA6ubXN4gxziRG1LHkr/fG
3I10Ad38Sr3fS4gFAz9TEtFpIZ9jlP8qLMxFeGicgwVcdDR5KEa3P2IKRTr+NBzlu7MsaO/CFOYJ
x5iVvO9zUpaWNqob+v4JLtZJDTcoXgV1upezG1i2NUXsdd7dOpOxsF3AxFrSoVimHOWUOs22n4a9
vSzZLundlzitxUZoFQKSHFBqfaXaoUG6B22kE4pdpycoIF+09CcMGSK8jkOXaluiPHBlD5GRzN5i
vydI3WCNzGF3AtpdUicGd6BaIjd/mAEieonNx1u3OB5jDiO9J7WgGMBI7VydSil/64yQ6ypMpbKL
nOiFxIpX6AsScczW6pqaT/Au4vnhREarq43Oj3ru2zSeGnztYpDiRqT0zdizu4mQTlSz2PCVG8Ik
1jsi7f6GBkWNOQ+3Af5yi7Pz64XkyeaVTzcBzZ37V+JQN2wg0I+pxaaTwUp77oqfDjFh48CUUKVI
oBV3/6aNrKQ9uy7mDJ2aNgo9XtYLHhgoGvR0jLN1zY6HwWL+Qo9sT5BTV6vZTWiiAKPXbtfbjpYZ
459DZOTAkvOONJRWxgjlNZrTJDxAQbrWWhwDj3ALwfhGj/rjmVWWJ1sG0eLscwO0gBNKpFIukjMM
42NJHgJfFiKypQJP8JO2bnyR6F6KXc1CwRwMaUAxWsTtrcCpm/zt4ngY08qZ3iyQQgWQSNYt05sx
29Cd2b10690GqzIJPlCX5dlKindhKLyHp1xfUH2PYGfTBoX9a/u2y/fV5IrhRw9Jn331pVKJFBxo
82Vv/rVbvo/fh7EBuv/WUV5gnzcDLrn9W8QOu154Dt1BQhCVdQ9pJW8Xm8n7cdDoXCAfKyjds5D9
UxLJU2GbnxtNslnIY3qptPyFKq5/QQkT1cf8bif/bYMxYZG0S1o+9qmy4+DBaskWgpNh4TmBvSRZ
Z+uLFGKX22P3o/DCnf61HVPPVHfvMmwRHMqmBS/ADDSMAUUHMRGB0EQHFMs7K8nDnqe2oV8V4WuW
iShJItDZhH4vMHkoGi2NW/BEJvg+a6iKjbcB0IKASmEWotfZMVqIZ/Fyb9XCQ+GBELfOdNDnMEM6
9Yg0WsK5uM/kd4rU2CiArfTw1T09MYZFu11eH0LRdgfSgex/FNrQrpWRtkPGvzu7lwiMh2IZ4DIZ
5cI91PLAIbg4T2X5rw1AdpUoxTDuYXgaDUlnSN9W9XeX9KGZ89LjeH7S/rxyaMLRMOoXy3KZbroV
pc1lAhlbg+H7eQYK3ueqHwXWx2m2retfY3pSV0ljfeZPrZYABeRFFhb2H/t6Hkn0QsqlJOorH02M
XEOiLJWJdvdtw8Ao+xirZjuVYYIdEBohbaUzn9E1piL9pc3r5buf08qMO4pF+0T6UCQxGeihFOXQ
6wQ/NPFWR7MngrZA7/ALrMDTfBEc/vLmqdestE2iRHNvAeYPzme1/YQAt6FZgxKzk/OOBt/MuNsd
1MOm3KlQItGR1ttIhgiz5qWIaNk8IdWPwYPEVpns5cvYPwrNmhdP+/UHRMlpUQn/OdTQ5M1Dn62O
aBDfEp1B7B6z51OWJ64aUSPwO27F7lNwCHkuoLSBlxsllcExuwl7bnMk57OFcdyIoVz1JM05slCF
mO4fblqF5/RrikY7XRsTBOPmrNxW0OJFZtfONwXN4PGF2+EnQB6/cB/ZyKRONxcXu5HFtnk8OFnW
NUUJ5aI/R6bFI4yxjRtPim70gPVdroLO2FZOGckjbOWsPwnHnY/MtudUejygVB6BiDS0Zs4KN2iB
C7cZV4inOQFITq+v1qXgJq4csyAGlWaldZgDrrE9QO7GXTx3r+5a9qXTrrxFLnJvt8jHPCOrV/jO
gS8P7pXCkJFzSuCURuk6vdHHlrYclCJC7xLvHe3cMBZLJYapzf4+RTH0EOPOmcnC+PezzZttik12
SfhYrqnKdTgxb8ewmfJY67on/UK2V519B9CgMrxxicX6XQwqBjpusSqANm9nEB2U7F2wGXD7VbU5
fDTDXCyYGjQ+c4OFLLyS6WLbdNrl4FF8wsQGqQyYX89jYwogI0sArUzuH4xJrmLvIsIPAaVid9zY
4tAb45UJEml65d+trMWtmchXARMFLAOMTXMk6WYpN9NeG5kGmkhtq7auKFpbBh8s5ZVVxi4Qz8Qh
EpIQuHZOjKi3z3vGKTiHod8ux3u39Nv92Wyrx0L/q/qEqDVIkIIIMKaF1vSbp6WOQHYIhMP52zng
MnaUZz2asklnqnMdZW0a0WNhKggLPNal204epeVcr83/ui8SLObI3Y9gfKcjVXY0s+gZadyShWcj
t8o7vYIsgcJZm4/tmxVLvFOHOA5VkcKvTHj3d6UkNnYVcNv0gbOG73fEFlmjRONEFPB+5bRUvToY
rrM4e/omQ6W52tBjOG7kook5ff575kwj9rKcPbeg4Fsq/UXrgvtKdTYr7n4S8WMPU+WuD+UztywH
hxO/kbT9EkCXkL9AwJl+ozC9g5UGMChBHEvJpyUPwYl9zk2+sCUVcw3qo79PrC1DgKL8k7WQoNUS
2ACpjAcH6lFqHxtwmQShFqw6u9JAK72RvRaFP/ICSy0dMkG+ls8Mtlw0eBYxeuhMl9dcgJhs3QwI
ZN+jphNwFYvIfPMmalir3AMKUlaLvtcnDQKlR0FPY9oOl18f9yYdeLGEIUiPMexZnceuTjMbWZqj
xhIccJPZ3JAJK1IuTrnB407It2DXUlsohS8OlA+zqd2k/zl0ayBUEncE2y3lauMbpWyvTWlI8TuE
OhytAZiJF4/JvhM0sKNdmN67u/Iqim8BvdZ47NNh1OY4VCgCrC0F8lXXR39GQpl6SVr+gh89J4qv
YazvvRAayWoMT4hKWwEB7ilhGfCh9acHbT/OD0JeeqBHIL7Akc3VHdkzgmez/BKuBKFP1mjhyb9d
dREfkq/toCcIEPqv3u3lfMuZLDiJov5Bkmtwn8htHdIBB7OLbrrrbjqHHmrFN7z7i5/GkdfNVy8N
eJsjbe4h6wBq6mPiv2kTk+/Nm/UacdHkJ3RaHw5NR3ZS2ufqGRMkwX1xYHthxlddtis+vdmBwslV
VIOG4ebXxh+uK7mcM6Kl6cd378I8Ksu/p6ShlAY21W2wGz+xInvUfJd60dqx0Yo7Fnhfm4mweG0E
BArpblNzJQQz9mewZkLnoL42+YR6vI7ZyJOcEY5ZSOJ02on+NudeVYY++OExS40PmpM49C9VRI1R
91sWpsBylwK2/MnsA0m0HQLKaISQv6Kr6RxKBYirXZXYW55EfN8kj57x3D1tWEFZalIkiAWf8KQy
JXLwoIeEKfC9ubPDxplryZJjJhktrUZ25MwzfkVJDm7G5vA9MBHAATnphDJjESz/FTZBMT5+nMxJ
30GZhFHKmWhS9AiWV6xJYYAECWH8Krs39ToGyrxbEge25g/rhyh0OwyCIYY4yrTlfcNM+kqPfnQl
Y5resRZNLwhdQpPco8MJdlQi1REfFGa/6beOYNepkXMFSG7aySlFFVBdYPQu03Q4qCx89fiOkkqA
f8WL+5hqf6g6RyurESGbcW9dxRinISjbCCUYCbIZZyjMRqaugBGIvq3+asL5BZ1HZZJdk8yo6/b+
fY0AVsixOaRznZJHboqGh4kQd4F5HMh+hVdJpG/kmu7VXI0Xoz8ndy3LRlgfwZiNZ6alQusec2g/
D767Y/z+L88ykYT2OKR1zge+OIRp8Qmf/sbsQvMWT1cUxtq2e1N+dGhZZRKh2Hy2xkMC0j9A40vp
YuJE33+J9DavYoh3/IyBNxoffy/FKvplquZG+ouVqmSQgJysqc0U11hCOA++27PzenoV8Xn7Rfs5
ssJQdOsYAiRYLGjf7YQ5QzWgaEZIHA/nToZSDIE2d17RJlYHFV2LsYygXjLB6XxfGCcxy2+ei8y/
ANZzyFRMbQCeQqS03mKOCejKo2zTq70ZNCadY4J9TQPmm0fRjpv2GoClLz9UiK+kPo59X4B5e58k
BKQDaPd7i8ku2b9q2oiN/UTKA9uof6GJU4K1vuk1uhlp/splcYLuHE7NavtdrKAGuIjT554Vy1mU
mDSD/2C8UbRfUPlwNHawQ5Fgby34zRvhmrbAliLGANRSNO+pUZEo8czDJhK4jQLIRSkCzJIu3Glo
nQutlNlDR9uwUT1onMv+kOYxJOIlLNor09VkSkUhN5dQTn6lWIFChzZyZVwYWVHA2jM+EiJLYcjt
XKLdnH5C4BdGDAGhm/CVHYP69t7FHkln80MW6i1rly00lZzY+IEFJZAp9vGTU3r8xAgJaCeuHDF7
RjzYMyr4OkqeEFocCS1/p3987S1wWrVkFgKj2xOqUuHtuMktWshr1gWMYMjT/C5SSVun2c4C1Qgj
Ery0J5p9Uc7b1I3mkEZ4clPubnTVxMnMBE7bvbODE5qkuTXnNqclEM6W9dRJca4/jvo8V98Sxd0a
BW3InyzHDfkRSkRjx8I070ybqTp5XkaxAE7lLO+VDfynAeEbFrBZ4eZxBrLakubumC/enaLJiw8p
smeQAm2gy2pReuriNelbFyztqVCrspmJuv1XOJ3VYRfMqkpk/b62acKC1s9vS/y8IO5mdjXObk3L
XbNUzK/DJOdU+kcx2DHu0PMI7IFByzK/laIBPMfUumTV4HlARABQH+xvwjOj7+SUOo76VzDWcvAL
e9zA8+13ZCklLiuU8BcQLUNtmdyshQz1ZvLmSXdEs26CNGJNplE7e3YEQBO/1+wbgNEiJaMn++En
lxw3lBC2a/MVyNbNBlhG3CCE5OhwDkQ9w4oDsToVuUhFabTHKKB4ZHBucH5zOYCP6QtGY6ArbNIu
WOn2kQ8n9aNkBMoabUSgDHQvSTCjinPrCIFfQ+onYGxz8yPiK4Mul2lsTw8n7ZqIYhRT6510piTf
+7QLMqnKG/SH4yS12Yj2xMFhxGHoGyvBbAemkYBeUCW1FbuMoXJGrmVgBslPsNEux5EEh0yglyto
/+x92dwEakh5SsLsRY+c2yYjd36AtZ6Y47UqZNRe3ZpoGBohw3d+KJUNQt5vnN11k4lrqt9+OVmC
jKFJtttudZ/jOJiSBwrplcfvagSEFP2ToWEtnyXiHcsMZMGWfPRTgUQj2M2Nv/QsNR/T89d03nlB
BqhKR1BQQJlSRAMyxSPjFvUOvz6zjyw7aLjbexS930bX895Gu4lzkkSjpK4wynff/QLdA04MSO/J
1aRq9O7TyNyTFfmebWYTxO6qY/eFvWMzYeWEI1nvMZ7+0R01F7q4e3gaGYD7Xitzmogrm00f7dMi
MY0VDWISdCscfcBVCak2v9uaxBXigQRUdC710hszQuOsvJw9gZCQ6YFX4Y8jVhVwtYSuQGaQr1FM
++TTteTjXttoHHu614LMqat2WXnscvxt7d9lbUt+XTO4uGPgvFabMnfrd9VFHv8Gg5nXfKpoButW
qgWf8EKQ6Bis+krk2zBVrfJYq6Cbv/qkXIBynnJak+1qd9A2fn+dI8xNXpHsSRh3unfpnl92nnIl
dvmXuVWOpHmIz+uuOct21YTJTaDFk1IyaqmFxT8q3Mf1syF6mmrF2WttSCW9D5ZeDn2SIRXIWPd4
5UI58LH2XECr3RseCweENLPA4s3EKaxv/vGf3+qtmubauN/V3Kdi5AvO54Wl4QE3mXODSqa3zbCv
3V3gcqjAzRU9qocnvd+6WblzaY8VhBs3k6A9/mKxmxROCsLuvF8c4oT5nxsWyzZqLGz26gt9uC+F
Q/sQJlxHVCCh35CaU3H9dh7z/6M2oPkJC7rVsKVhGq9s2rLKhW4qYwIJD8jd0MutVVz+QFPi0gW5
UebbJN0Jab6IqgRmBiJPdrDQGL4h6gvZsjo2n+iuZ7Li7tkKrkql5SWDw0i4ToqLsuWX3U+fp6nV
tCx/vklYjCqXt6hoyslUXaS11XtvFx22jkM5psPofhSwkhxV+WfckQIFMEgsr14Wr+vJPM+zkgL7
HdoDEIV/+CrlY81UR1xTafkzNfeP09fVITcd4hjIlpXvPm4bhcUzuxqVe3QRSF2HOvz9/u5k8/Ap
SyAUCZYKdO7HHDyXYc7WWoADPwZ+zzWfVYYy3H4f+eSpxWzz6tb3oLcYWMpBoBeIRuFwm2yYXwuH
rCVYuQ9rC4M+PnAxoMbXf96Fnhy+ariI2fyaCmKST/Sxer9vttGvCT08eYW9xGzCHN6s7k9EiDin
QKozKIyEVwZKntn7WWdntsNZ5WqGRgDKT2/OZhJXBmpCe0/QRSODUYNlDLdN3vyeN3niELInfdNt
IE6U7fuyb79Ev7N50+aXxyVKxyHJGB9KpREhtpPxY/nL3egXUpebZdjFfsT1DwB3C4LOZAgxQyQP
V3nA6+DeymS0AQuih3xK8hlTtPZYR9A2DDCwVKj0bxEuUFR0VApfvdYIpqSvyWe4ChPsLGVYarW0
aopCAlbG8IgPGqNokKiMw0yf4di2yvVinsKlbgMeX3FFQ+Kq5SfdYEiUkMfTOPoCa8+lUAmiCj0b
boKC6aYD8XPc9WvYbuilFPHaTNpZ0ZgZ9oCnlaeip4BGea+BNyrgZEe7BjoFcfsIQpt/MKAN3MEb
dkWdZ1Fg2Unpq5zutzyB8PUuSfQ2rB68IDj7acDak4Xn4unr/MBExctt949wnKRCgrHvoo4VejeQ
3gdn8kx5ICPXnkffrE3l2abgSqTkr/2ez544B2bhbcPx6hQdwjvqV7JIVXb/SRjySZBiWk8vlwdG
iJjxwepYg5jX6O9pcLFMxqrEwG5tDP8uw+dKnqgDrqCeyWIdbVmLAFNNcF1U8h/2CFqfrY5kkENr
ouqgoCZvYydSypQXSrxPq2XiMH3wmX3cm6yPc7giVSJ/WfszvAVUfCD5qD+xuAIYOUVJpD4hglfk
fZZJ++R/9JWN6vKN/E9ri+4NcTn2roUmGuqOHwmMDgBXf/tIJIKnva/7hagUFRjOGP3c2LIftU4r
y0yir0dfyEx6M7Ud9EhNwW3r+tiV3d/RgMJtGA6XSo8Sac/8NsCfuiWcgqm6ifg9Bp61qyHQQZ1N
ujyQvFHoRmaYwSuDJ9xsBXEgaPnBdiJ3Pat0Iw9MJ4KGvQ2jBcrupmB0DVNZdS2mEdsdUwOjub4+
afriuYGdLsri6XkiGoSD5O8pq7CMRBAkswnzmzecV2pGE2nX0+FYAV5iKg0DvtqWUgzpQVQziNIc
gpLIgLYRxrWMJmlcDCNrlFXgr6vfz5iGg8yEiM9vEWeYT8dOy+aN3nj/YZOkTcaUkn0VWB4TBBFq
1dQClF83WhMGeQWA1mX3oBmAJODrzEYOD9BLRGpW2SMb6VBhT6LJFzePVRPVIDBAYdj48c6ufykm
CwlnS6DZLUereVc8NwEXE/4Mq+BO7TE/s2XvV22iHeqVzSRD7zTvbY77KeAIXt/AAtJUP26ZYYFQ
A/DHHEzthKRLKEipibbw8d829rCQRzALgyNLsHyN8N8rkaT9SRFmmweEXpMUrE9fvSLXM0iXXu9g
2Yc/2rRc+h+12yIjCcMh3ukgCjfSqUgwB2AaOKzrjX8zfUcVcHrnHn+ZgKR4NpQZQ6cW9A0/kRAn
liJYu5YwhS5/l1TvFMm9q5sE1pk7LHdXdwiyPCEHlFcayQLBSt7gw2F96N1TLtCFSG5pT23kplhN
Q4H6DFoVIGanNCGUWyBRmRb2cqnN/3kNOX8ZpV0bK8Q3FFT1QCCdsWYxsPqES6CSMoNjeswILhxK
j7zLGo5qJB6hGeCTm7Szl8xlk8d0Hy5+kkoTHTESZqBHA1v6fGK4xuxjM5f+8JpeQdiCDgOQnGpw
9s4G9gNfbaO5mRJbzp4qjPW5ICGE5/oIDRrj4YlgJld3TuRVYCBQPDhR9PDWY2v8PRCBUrjVzmXV
zZf55piVzHC4WaOem7/zPxxXJ25+7OlKELoZgZgxnQNPpn29K/qyDvWsCFzhUbtWOwLHHtke54zt
PVgTk5jGV2u5q0YmRlPqrEYJs73pGgNq9aBTWxSjKwv/So0mcLcpLR/tdTnpTFcPfSq3B6f6qxD3
LJbbU0qXE750Hj4xGSw6xN8xQarSxatDiN4CffCYpln6ChGiur4sm7WCEvbr0qikWt9gHuH8taMX
jHbizOX/7cmBd5f/fymRtoS1Emc+fZt2tyo6duQt0Y3jllbkqnMMlKCrlx059MbtTKRVa/wiBk6J
1aB46ErmCbQQLL2ixakJDaacc/u8GjaB61xsJOdEANpgDZIZsU2qFSBIbTPgKh2+fmm5gy1Bp490
2QARMBLOuukpvig+2x5RyN0R7mDQWqm02yQNxCrcVkNK9it4CfPBsJnXBQdwgm1f+H7PuLnMRpCm
Y843uMPlXEXt2g0aH4XjkHWlC1GvW8pd6Evkjw+DAIeKGSCjB8jPmvsqnGjUiHjNxel+yTDOkn5L
5A6dNkh/zl0VsFvum9aU6NyjoN6jOqAyYB6e54ihKhFBpjpc4MIRBotXFieEuHZve50VQvaq5wmk
h0Q/AFipk2jMM92eyN7vMOtZc+sZCsbXvrMm6X0lABA1oCAQTPwk+CDbpE6QcE9rZPqmmMDyHGka
gXPDCu5I+BCSmNWAIfEsKhij1QsVN6j0tHNnr2EVUMT4wwQ8V+gNesw47hQo7YrGZ6BGygQ53hm7
HexHtFMUq9K3k8db9b5zs1iTI8LmL50YM6L4um+UogKD3pVVTBTQLCbjYRgJs6zNIA+zhwdmEwQ5
yWVsPYZZlFvEuHXF1zan6x21SkLM6xR05pPhPfGTSQ3g938ACiU0XDW8wKOVCNGhk7G4sUClBvnh
GxRReg51+l1DiwFNZas1uP94qwFZWZfr2qV9dqn0TqeQYFZracbnyuKGz119OCdmljeiyqkJBEiJ
zrQ5IgiE0/bTF4K9FKk+rtXnlkTafm35WqKWuQ1Ip0CPzOPN9KpccuD/3WRSGLfPPG6bG1jTj/qs
AkyQeHaxlvtygoLuf3CvjsUNwwhZmw/vstG6iO31thwh0DQPAeziTRV8UpFzGonyKRhraexgRDw+
9tRFAszOafq5BfeN0rO8fsZkBO6X/flnCmyL98YqgK/TglCBp7LtcHPphfv3n6hUn800arMqYxof
rmoLHoTGj7gYAMVlMSw0MsO7mJUPp0ZQqpshyE8ptBH7ersxJ9TcZ4NZDxhyo/NusY9lqNdKNQ2s
zd+8pH4q2Bl4jodJWPUPyosjALRKpLSQriX8s7+QYt5olE6zWuoU3ootXRYJ+7rFIYJ4lNP1aS8F
Spjq+LXiMAD9uLcQz6oAgU2l0FaxH7p0nlOl2Orqvil+WhbNMu4kjze9s8VL4qF5wP+sAePX99vQ
162Pmyg9fuzMjZpWXYzpkz6zqFuFaUMpJV2slsR7DRbIvFjG5O8QkGMRqPOTfV9v+QSvSHVs0byQ
6IGhCr+570UgNP6Sn8vuzLQFVgCQUDaWFC3Cm1FmWeU1qv1BjMDS7nBE49leSwm6oQLrId4SbY4d
1Pfu44u6dcOkF3tDfpbYh05uEGpPX4SeLBgxrQVpq3+zwJOAHXchIijpmT3jikHu6lUjdtpGGbiC
MlEPNs6/nCMoSHRpWVv4g2oZUETYlvgbBkHmARXHEtD1rR4FrIRIYAdMfaBAUOsF1WPfKp2rawJt
9oPFy/pv4ZBV0Socoj+tSl+ZXGb2D2wLtkmRxZhwwLiFIdFNCpgxCPVU0ludZ+NkEsarZcvilSgd
/6teytfqOnR+znXNju4wXl1o2NS4moTEbK2pgKIk5CIwxz8NiS0QhHcBgsWhTqNIEEF74Zu/t0iH
K41Tv97CStNRuq1kjoqDTHnDUl24Pno/9YvHebZF83Zshp+DeG+CaG3+eVBsvTO34R820ZH9C4NI
IJxZiCpSAJ1ARkWJNJQobGTmTx8PRn3NHNaI9K/Ga1fKnDKqybIS8XTuVWADezR/mIdzT4ADLUOl
9QwTDonzwXItaZ9J0j/j2yCwmLydE07nK4XI52mrBBjPgRTdXCspSWfsCJYs8UuYmtxUd09dAOiX
czMsFF2f4utgiJEp7PIlpzx9nNls84BELW9hQH1ac6zn1uQvr0i7GCUpcYkx8tDyK9zg/nbFn6xK
RJwp5uxoSQnhh0Gqt/M8DwngZvuWHAcFlGHL3Xyv3grsCAn7fFySqqXxvi79EmQbrEYLAzOYLVs7
h5zD8VKEJQdCvqX/VrgGd+dPVxDEzTrpVnQuWOtqzpU9Flz4KD4HR3DapVBdMA1I+kwXSb9sle3s
mfEQfMfbKHEwWelgHJNuijZ94sRV1XdS+TRc4qWDomNoPkVZqg8z8Em0n/BVV0oJnoJ11dcm/2bE
k7qLRFgVdKNKRKgp0YVPUJjHTQSTM12LFzKRBMr3jy3eFz9JVTV4ovphU1iPAFRTFTf84ye56KcO
/KsopVaEShmlyhUrq9Bh99h9yKIV6OvjG8VVAMzdWer0YCuLARU11ABMt/LFd3GeFJ+y+f8SGOTE
QjRDXonNINKo+k93iZp6fvLz4qzbF6Mst9Q7dkzgn3R3N5oj4ECEv54NWAXqjSWiwmz3+w553BdP
iweAu/O5WlDqA7NYLJXI65nwDvQxt4ltDbo09gxOUVqoEGfPLVv/lq+i03n+m0PJy8lsDWxE5P9j
AIXkOxyFjoA//oCArkFw8pZHhYkKVMfXeUVEoJljdce9hngd0JmC+a8tHPTy/q88jXp2aKhZx1xN
RmJEPl2Nm76lwMSygwlT8b0n+CFszaFbw3WjLHq2ybLti4fq46/iKT2Chx0Z5kzamvx+FNz0URg/
HoBJlCpwCPYwykfG5LYnyonOlYNk3/cJkAC2aGvC43G+/AX8G55TDWrHIndHVcZ/TXFrRzK+pUrJ
U6t0J/PMKu8fuU2t+FM+ZBUB/HXrDZ1X0K0ajGLOfrSyRKNytii0VLbmTR9yCqHi+5npPEJVKZUU
j8ug0lCgEyVDQ075+T2Qr91dr8GW065FDGUOM3vffqXw9SkwhD4gvUEfd9zfY2eFCorhgz8l6kRq
O/iEwGwxdV/rUasxHSCijHLtKgX5uYaHQPS/xZhPLB4dqX0fJ0DGAV0Su33uEnar+j/9u1FXb9Hx
18LwZwmFwTxrPH91KVduuAKzoMmgBfPLoHkxMKXbMap//o0cgO+nqj2/+VQDfXiQXSxNior1k0No
hmXBBTZ+pfN+VixcYCVZa+POaTlGg7ONJCgb9S2WEbuvl+6TfU2f5eUX9FJWXecynuDvnphcBTF+
mggDInEXESSqpfgXKi2wmy51pdkYTm1aJk6eq+HT/hImVLupCI3GNsjajY0wJWgskOUfcZ9D9mqL
nMTjKm3MhtIkaiyXO00oeqYFLokzRqyxhtCUf1jlgNjx+D1rgdZMkTiuNyCYxFRAnZ3GeZP1HgV4
vKwvQEDkv3+rfzxbWQHcTGNAwB2ee4LTbTfstzhN4MKfelHHT65O7GrfJjlqUCKBuitFIo+jhf7c
68tbyeSEJ4SxYRJr+5IR7OEgFfS+bZ0hll0Lm/GR5B1XPgMXXqLvI4IPKdmmND08MHyaxHsNLblx
ydXm6LgOwYW/datAHY5vYA3iLXNL7fklUj6zcIwMVYUwxkZJ88PAZLNz4wiz0JTWviDlAq/b/kan
paaAyhq694QkjDhz4EfRtVKd6+drceOJN2XNs4GKZAe2WW0NO5XXctRlq8TyontIe1tC7nQLT0SU
nf8CZue3P7bjyjPmr5GbGkYjpmeBEVeyl/vcrvjaeDPYiauxVrRlp1w3zSTgsPQPMR/MsAI/U5iK
U56BeQMmtmtDCMcderV4e0ySgBVhm1ZabOvMvtHuJifatAo4/X6VgoNHRoDdepJr67mbuuOYT+7t
Wg3d2FZQplP8FuygbFHagmAMhJNeLsbhingfCY7RzIOMzFZGni/9KfBzkmml7HD5rkYPjM8o+Rpp
QEplilEXdOTabU6Ee1dvpmYZS5YvtnVCn4U6aH0PD0bfCayem5oUVZWoxpGgN2MQ1f4Ty3lcp+39
/qxCIrWvrozzMCoYV9ZmIch+SKcuj7ej8ibkg4apqVr5YEfSRjXrxJm2zs6sC9nnDqSmxYC8crsr
oLN1VffiZ5LG+FiXM/h5WQTV6D9jq1QtHCf5RxU+gIPoVgOmFJXQBG4Zql4hj5bOY9uadF1fKPpW
IOAmAcpIXaaHPchDSdp/dsDyLoGcfWdWCHyQZedDpika60MjTA9Ny6u8rxuztYGzKTZuuDl462s6
TnGPzd7wdidmH01vuv1EGa1I4MbMWKC7hLHYY97Kz53Dxut0CjYHUn536qb5Y0t1MzaK5UGQQfgq
ft69XOFMRiyTjezTAkZaFInKC+9ZxwaEI6I4IejmE6gZyfsbd12w99nH3sEnUt9Q3UDshXRV6vZl
9sH2XC8nmwQVziRKIXpwegoN3yBYfe9iRmOyhrLarVAYKBsqrmap8NQVeh7igB34zwYIoZPvY0kX
N86z54myUe46FET8tHvd49QjzT5b/nybQP3sWmdui6Z/PJy1UNEYKDCLamNY3vDBpR+ERNNIT4M3
cNQh3bOqxq+O2NxzDIZ/fxOJaeMUpdbBNvyjF0+VjdqXslT/J+jvVEPHTWOgLri6KdQ3b7f3VN6f
D5oeZ1CH0znNej+5xZ5ZJpM31ZGfHLvpYgtySwdY5Iz6SxsOL9RYWF1A9JzI0qygzEme4nA7eR8D
+nzN9Ut6vx82e58pIdbSxN/9WkesoKP+vEa+E9f3p4DghaHV4QLPmzctj2vjXBPsqVjq5CP9Gdz2
4PtsWcDlshB7VUsW/n9eIYMnSRz+daHgNMsHng7o/4zdkenonEP5NsjZXNeV0vsPtAwvOfUNjrak
4bvP5CTf1fhZQyZMxJRPIRPHOO8YvR1SeMwANB/u0tnkgzXaakr2Vs178eNe5t7hthWKFuZ0iwyJ
+SHk1+hd1IAvlCQalm3afkoW8cBQZsnnzkZz4jPdCrSApTzMt0KeFLPYvw/Yyx75TwyQeE4TQFqj
y9LJsGX/PjIOklUcXlpyklffOaZ2CKYRERvKIW/aE1KPOOwKHgRh7wpSelXbR7bGdTmXeZ+sCuXo
1v9lGrO8OWEfD/lqcpzB0b0N1HH9IT31q4favkT9ZpHXE2gpTlIoCkMOYmg8LJ0XVUfqA5QXo8kk
iQvB8PfDIFuan5v755i3RzQHCjLSa2lAQlX/SZMM45xY7xUyCtiQnb/8ntUAdaws6UQ7vMUV7sOm
Kt6LPsbaHNXRzVlHGpM5bgUt28UKrFSVQFY4I+Lnmpi6wT5extQR+WV82tw81CbVPh1ynk11mi1C
2kE4fn/bq8ldlL7uIrj73a6kN/DygfZn2Vf+8c0ptP3eTMP5z6LheWCL6BGc0Uwk3BuZJswyiDTq
AFEqrQVtFiGob+EsuvT2lfd6UAhHtvVZ38wRb9vwksS0pkJgSE2YER+CRoN47ZbfmSR6E51DBR3O
75SlY6YO7AnG503v2wO7rK4Y1hkGPfAQ4sCV1AZS/fV2P7naedmwakB3p4qv6NvnBbpiFzd/xa/4
7PH0yVKgL8YE5NPiX9ZCR/0vuqM92mVYHbqTHPcGAg4b6bN4mPx4xRf8Va8gO9TXd11SgbU55vqG
dEFDN+nJYkO+iOY0RcOvc01FwsvajCPiY2JXgcQIqznU2IZtMtyTIYqHvnkWS1OV5OuhkDqsFiVo
pKf9OFJq2wRhz9o2Y790YOj1bhnUTbiUjPzTYiTJVIT2w4q4T7Sbb7C/Pi/m0/3mYol7ocfM5Y3x
X+5de/TUEdYNojzdeXHQDmawEpuZSCGFeTs1rw0rAOMgf16L51dM5zSFujdda/9dqYzSa7ZFEKwc
TEW8aLX4pxAvVGr9Z/Fkibeqrkw44tKXonAWWEEg9UmbNMHGiIgsg7wgvzSfyPnbl0uuVntzMzzO
g9CJwVR0R6EHXRGQ0+LrwU6ipiufv8xSSbZWhu2Ub+EwyozZTT9GOotqSDNY2aLS2Kh+6yd1I3wg
KVrrcD96ZydcKD8DKXjAOi6qegmNHcrCldRdsWCEElZNMKWC8AHBvzVIdYtto7m6KXMRM0BKW5i0
TfQAg1OaLYydUc1x1lGILZdGMa5jaZhhhy33/lafX+iWewYeQol3XkxfaLM6Qjd1sKYeXxi4F7Tn
kym1KFKXs2tGzpvENgfuCHmRtkX/Mcst8JKXpfToXvBY6SvzBbDzgA8vdvJ8iDb8+StHRk5UE0AF
+gDHGLjGDzkv48G7XvkaWceY0D40YiyCfL0sDbx2T/ARGkqjmABoXKvKhLneLp2yW+dsDTobrvvp
0IaSndyrfet1nPQ1zXDPRiRylinewnrUg8pBeZmLHIItT6Rcxor7rm3DHxUk4Py13bzQWKhkPUNb
pRI1XvcfABuXVzV9uUjPL1HQ74aqwx1TqQi246Tx9eUMhQHVzKkWI1XV4NQ+IRryM3N412FH4fY4
rGsd4dSZV1bD/fPnwK+Hx+qPpslHrbB2XB7R1Ic0iQp5d8bmMiS1xCKc5FAYTP/iRAkCVXqxXkJp
v0Tsev+d4cdDmRLN7BjejIztlfVt3vEuhoCpiwBY6FclUFvb+XfNLEtVADepqG2AhJ3Z6KLGNEU+
FrKmy5n7AjaZ/Rg5SYV+WRfN+A2+de+j2oz7qKztvCnEUsBoSXpXIEUbAAAX5IFW4E4JS1QJyOFf
AluHCctISLTAdhRBL0fVPv754zXAWXR6XBJ5NezNbmzcRj80kwLu2nJkku0AjsSMxywrP94cUZdZ
NbInYC6QCPBnvba+KiIfd9w66clHsEX6ORNNxaxaBb/EX1LEy/Mdq5iZziqfyRZhhKTMfHC8ELtw
auvXfYxYxDud91RDvLh9TY8BZtvAH53cdI/s374WFHTpvHMcSn/PoYk2ZsSTdIJbhBTwer7Bd5WF
LALolug9WudhamYMgjJzI+n6JnPvQFYT/q8liqjE2imD7kn+xLSol7oTXnCDBztx/ICTQFsN2L8V
PiQ03LcCd+SFYaeio423k6OXGoNEg8uSzktal3PvtDkfJvFxWawVyEUUXeErJcaaSOYr6qnvuWAE
qf9DIqzvWUJfqylkYvg0DNzrMHiDAT/YG8wLQnDQ1lWlc7yKtHcr9K7OpSv5JBplRN5EuHm7vkYe
rWebIWdryVFUGwYyuXI53G8AV6Ojah9os0a6RRlR37rXwrha7jv/IRDLR7iFaqGpN8qdODiJjEKr
UYekzSF8qtwSCRmHoh721I75/RnUgmJc3uVscqTZAduIEV4Ba48FeSOqlb1dahyqkxDkSe4/yiUL
z5p7t7psYeFqg0LJ3deWnugOsVd3TClOQuvpMoX2TnPtIN8xY4spFNFGgn8AsYgFRIt9/VutsETj
ovses0H2jCeQIn8xyv19rACqRDWzavcL9pILmjAHwFRva7IWZH1pAnZEXFjd/iLXXuCNgOtRgipc
Qqe4fI2OfXZpsFzmguPIw4b7TgLAH4vbKWD/ONJ8beaSZxPDSfycdkpEGq1sEjViZuNZ8ICTKh9/
XslI6TfBh7qJS0P1y6Im7R2uG2u5BU1TwEAZGL7Mc0eJrDDopswqqzGMS0vl45HnimjDmPTWaybY
9z4+W62p8U6Y3mQ2BZHBh7bmZvZWsyKcUjqS1VPe/oUtAg9DCy5LkxrjGo1YT/itUm0BaeHPSTJo
1rvBkes5sguEynnYhjyJIToBiEEDICXqkxrZWgwGoPguf1TwCUClOevBef3CbuHsLyIlZg9edbx+
cvCzdkQOMmBqt7O+zxvr+679rTexe4fMvwzUXkHBI+gxN7zhynNl1Su6Xj2Su6/zKoVuSTQupirT
jW1hbS46wp61uS+10n1fU3P91TKYMFNwnxTnFMGGc+Oj6aJXKdr5uNfwZ2WmCt7I3n7QVBI0CNck
WOHPTOIBz05IfqWR1RtjjgaZSzzYGBfgQfPbQBMuCrRgEFTUgCBi7beO5ZUr/MhtyPqLUCFnmn7Z
FyeEKCqOR6W2rxHu+TynUtjFD4FQamh+b0k9DEu7gD6eRc2Dk5JhdqKa+KlF3e3ivSQuSGmNCcvC
KZHYD03mnvH+XWVDcrjljOzDHShLhtNtWYkw77TfWlglR8UMdjAoF8nkZszhoFQS5YG2q/6Cniny
p9fAiDOqEputWibs47iJpoHqBhP1+TIhDVWuxyuk4Ikjrk+uHqgcn0I3lrq/KEHGCSTAl/dUf/WZ
98gcQqzEa3ymT8ZFPo0XwStxk4BUU+Mtl/MlgQv+2vz4zJh4ylqtzZdX0EWOgyWSODZ6IzAIpBh7
Mm17loBDH64+lRbn9zFz+Eeghf3Ewr4Sk5+HugjFHt2TZbDHY0Ll5Xk1dsO5k17bgPaDT2cX6FtM
UPgf/wHpUK5IY7z1B4QRh9yJ+P/J6jViXoyFFDqVOiQukQl2GkKUwveO+VDpPYCd1LRxtaFyYdZj
wiIIKUluXZjTj2RlIiBgDJLLIoblpVtAaUhEB3m5/82m/vuht6BEaXMrd69YNNo1c1xuGpyli79r
6SHsidca5pOjXMq+I23aZKjT5ZkrL6Z22VFQ5LGT1ynrAcAJAfI59EYmrG7n0PuAQqfsDjNY69aA
zlCnSE4ioYQfLHT2bdariZsY6XkhRc4LZ3GOSt2LpjEo4lllH8gx9fNDma2YxrJQ55CbdXVGYrd3
mH+Ci6vfPmV0vpgjeJ0EKcrZrJiTqB8sp9ZSrKObSLHEPQdUFfkjpZqWKexzEDHnVu9KN0H/niJC
gYu9MCRnRqLRWUbTlU+rPCvWxPtALg2/96mkVnayUSveiJR7VbcKrc/3vgJBVAC5gOyDgJiKBEM4
7BXcShFFDkGv/slsfv/NF1SO2S6DmLLov+2yW4OEQxajnOX+Sm3vpmScUOn9H4dzimMDbeOruGts
jjI4aTBd2Q0jXh9cau1eyfTT6yolx52olQRna33xxL4bh1X44xggrn+u0c/dmAJegw668rFWoJc8
o2f2aUpWzlWZbIh+hQy3wbJYMKke75lPBRMJTwuVi/Ieck+yRfbhEX/3YfnRLj5FQq4JI59cTqu3
Ogm8XiubASnCw6LUTJbaENQU3y8BNxHU5uQ7MJfx8USj2Tuk0RW1XcB7e4tZIkRZUsIYc1hVn00o
qNFFETpgXebABOqCJrBkutQ7GaZfzwP2OwXs0c07h2zkKZg3g99PHcEl32FN/30NlSq6/qH2qOfZ
hEv5bnjhDInlTnHzio8j0jTxQImcYmEitsOh4mOD5g3XIUTELuLjSfluYmx4gzadobNW1ra/nWYR
e1kjp2pEr4BF+brY5forvy+NNvlPIe3XEckncJBitqg4vHd56NAGDJJZ4+OSzFlWySY5ZOpHVqjT
IbkDNSZP4eXhvD+hOThVlgKtWGvHV3HQw5kCb/Kt8twJ8+vlbZ5JRKkhRamRl9UV2i/CBxQhQcK0
n9iRU4JLr9+qTjSxGMKdsf7m1coV/5C82oqhTCccHM1ae4EDUSwjiLKSI7exVUzd3nPtfmJESVr6
TRBbnd1Kv8GyBMHY43cYxR/4LuWtK809wvNYc2Y47flvfnLzQdvZVYNHplK7bagz1B/QmEG9RUKI
Xnt5mrzoU86nqNgHHC/fN2sHWFXadohLUjV+Rcwm+J+qwy0t25QPrblqGQIPmMjd9Rrq7NXWUsPx
1VvMoGVIV/TiFDMvz2h+b7FmhXtA0zCEdI6sRHZ7oo4MMVnZhuCUtxoyGiNcrdGUEmeVKRQEU9zt
7H5uwm4s5FwQHCiVO5Qg9i7lADZL+YSeJynQAPXwl7AQkHBLweCvd7oBQnNONZQ7Fr0LUFiDaTSC
CQs24fmEvLsNuQklEJCNWlmRIHOI96HxuLBCHNcAg+Pe4oOWzUUzbhOkJKXEJda/p+b0e9AxiRax
8TyYnr1uYb54b66vm3Pdi3Ko20WkwnOtjIr+pMyXC2AMUVSwNMU0WQLAIJ9B3tnzGQs87fFlr2K8
1Jo+QjxiWoDG36bxq6zkrHmBUpsY/oeNYG0RsZoMB0VtpeTacqwWZfy/DmagM2H0oW7ZGu9FinCT
reMl1b7noHaM3LAyaIQhHR+59gR79z4Wcj6hLoDHXVGjgKnVS66Lt6G4ZVbJ2tOPzTPfIF62G1V4
4CJeyhzV9CkYrjNMycxf6ENWE8TaxpBGm50CzmPoK9BkxgxbZIDvHKHpobbFVxaGyYlUItJ3cR0X
qtRx0yzzw9uhUifQSL7VhX5zT6d67ih+EMzbgsi43PJjbiA9KDfW35oMzfQeFzoArIkgv8o6fZw5
F4NM93uH/q8cu+D2+CeUohlH2muu4CuESJ88dVQX25FKQriv3h1itfAkFMDR73XVL+SvcwpIffIp
4dVBz0yPVkf9K6J0eOoHuFyC0EMkehCw1NolW6An1Gi1t8hjIWai5b/2ECsVM2+0aMXBcgmmpdYJ
9TOMcDifQssjZIasEvE8kj5Hyql4BVhHcYUuogrObTYnOP4iv5uRJtR5i97FzvQ7SzsouXw7Sawl
w9yP6R4Jz8DgLvzhY50iVatDK0m0xJxG4LCh9ojztXxeZu3zPAXJcPdoRPsUqX4dWDx5PiU+rHXu
552iaM0/kemmtYq0+EE3GT69s0erwFmLWBx0FYisauR0gESvKiZ7gQCNVU8WjHNUlNfapMx+z/fK
fJzYkb9aa4HKjEytDbgMC39fc1A+UAIdafv+b3GLQvhPvxiBdjj6te06l8hDjnVNZe8HJlcspc6t
0tlZV4rLGHskd2BFwS33dqqwHZVDTVJj49Sh6PA13Z/776NtdnAZKV0VLpcV5qJ+N/JLRF2RY1lg
vLdnx8U26d5/HGuOq61f2Nhx31p5uPxKreDLK+8b1imrVOKjmmcCK2/uRk3tSTzes8+WO+/LB6k/
GqTtLzogxp3yfP4SX1BBIOMQ/b9k4HXp7AmRA3S4E07cEGW0JK76bO9X/lJnl7+6AWTNHnaMnLBx
3XgGp+l38pK0Kg7e5WBd029izpX0E3xVu7mRp1wdtbI6PGO3ty4gOIcqKJ9QyIe6+nOSgLRHgRs5
dUCTK97clEi0pJOtQ0IW100MLSZJdPVMN656vCNgAdb9wYlbWJrVV8NWFHSlj4pYW2ddJ5FGWCeF
gjfjTMuKzuOva3tmi1UkOQFlG6tVreKb03mCS2silrED7/uFSdvtIJxRGgd93MaVpw5GDskvttMY
55GwmqnDMhcFprsP4m4uN0rxMrwh3WZRfU+lCsXq/blvYf3BFkk+B4EdlkWwlYjg0Ov+vwVNVQJW
QAhUZBpf5O0aTKWEfOavFdo1L+FvD0Uu8VMyaEGQXywXZ4lqProiLU+tIUXUStPWPSYsFOkXBR9A
PLTx6Ec/Oda7nWoJlw7/HdRlkgnYbGbRkZIKIbc3ozNOrYVNe9t65beIZfcq7hp7Vg33kouaq2wc
M+UzYUklVaqulviOqNOueJ7EXsJ8/cwsl6Bu4+mV6LbcMsldsGkOl3Kr2gnNRaSsav5gcct/LsS8
NNv56TEaHkB7xAn5p2Y7Cqx4jNI7uA90aFeQQmM+BlH7xZ+Grr8xGhn2RdSJK8SeHwdpT6A9tOKz
ocRU6mFSZk2+g+lGRwPog1bRwRLwyS7tTNYsEmcEnUy+myfV0M1l/wH0lhU6JY4QwxhBZC0lSZp8
FhegbfUk1QqJnbvcExlEBezsao9077jgV9gt+NWx937AtEDpXGuX0C8rqKcGOSF0wQUxCVdhaXEN
kmopMeHjeRk2knNWkPyIT24tF0+owGVbe6/Ze7Z7fsw9iNEljfGGlENAsGDjdDGN0btxM3aEX9ev
HaYhidznG9HPTEuIW5wBoT5yugiO2IYPOWFCkA7iD4obw3gIHuayrv27MjxT2zLCCUbpAd0xfyoc
+UVdlAg8djQZ9ls2m8NK+/nOwvuYmR4bGTbwUGWKOfjG8BSwNB8KN/W3YfFOH2xxZNy+pwtVysvj
uhdi7KU39b3A8XoSDdRN9VXNPFc9nWOcNi7eLwIsX3QxU6UxqQXrB4+KGSgNJk+xbLyHb6B0BO1O
fOEwRMkZVsL4lYpjJrx8BZv/HiylT/ayujohcaATTB5cpB+LEBwSjZV9OfL0h8I9hM9URVy8TN8u
7BmkbiTWfrLeVpIqs7HhTFv1oIi7C4jtz0jM0VyzXHX7LFWllNjc4EhTJd27wAEiFGH3fm0F9Tn6
nBvj5+Fwf9NeI5bTaGeq+ZNUfZakScVKKAvP/EbYTqqEqDoZlrHLOjyCAcFF4dp0j2Tf6C+ZNOtb
fn4qQFuGo37seQb47UpP6Q0ZscS1KN78T+jZ29oQvFLlmFj8I5GEKc3yifxKrWUvURR9LH4PmoO3
Tt27YAGj4IMEoT+BZmx7lmYE1YPZzYv0Qk/9iOPzT332I0TYiRxFiSs+jsN/lp1pS6Uyxwe5U2v9
v1ZEkQ/TsB+1ezm+asJwUcC+I8cCNsCjYUS5X8fJdewEV4/GjluZXH9OYGl/4MYESR47VWihr7WD
MDIKe/whRFdk/LEku+E9zOatllP48IlXWx8z377QRkvr1n2zt1xENBVPBBZu5qI8al494NygSGYU
JocUz+e/zbo6j1YHsdZ8scC9RKUX+3k1wCM6rdFe3rRM+Ugx54cluH6Zcl/lU0P+uvGLfVyWk4aV
fv+pBfbxL1r6n2/g2abM/k9v4/lnfmLtGhWilyUYWlwUAT6yYVrFuUNP3NLTtv8HJDHFXSfcTlPD
lMk1dryHH+HdDWpsCnygtd0T851EC3o++yJ7rAYcxLQbJD9/Mku1vRLPPoZ6iIRVjio5nEcFQk3O
7Jp+4hpcRjGoC/iVgTBrjy0uBgEYMZFizSx06S+wWEVFWAn59SQflwUhZR7J4bynrILoSwJIjUVe
ZK2jGYdRP5rRZ29qRYdb0uBmMiPlcy8boY4nl62xJJrubd94dG9LO0nl4+DPPeis5rKH0tzFAA4U
eKilY/MLU7fxFvDxE+2m3/237d71yPHAb0wkm4J0Vi07AQAegAfiOwnK8vNlii/c0UgIvG6Hs+H3
xRysiTFSlMoAXG+AF/SuIJ1/3h5RVILkzE3h5KN1Bu7svfRX5xI302/pWa4EahUpEcGqUG3wUBI/
Yv4/lZtD77FYkIPvnjfrkhIAM9Uk/Mv70CDD51TQu6yb3fxlUawV+AoZ3ulc5uVFXeL9ZQuCRzaH
4qTIuw+grlNb7z97bkTOwW9q8XtTKx1JnL65bUalvxtSaziB5pZwY6ILpn4ptTYd94/u6EC0QrCP
SOCkQoelum/evVgogmcpjujJuVJIFIU1YlXTOo4ffy45Khw0fgFVCO6Xbcx4LLIfx4MWP6n1tLmT
Yd0+Zu3i9mIMCL9Mj1ljAtw3g3HpL8BZIyUYrwxr0YeDC6Sx8167bsnm89hoHiLzpY7B9+PstFSZ
o8NqeQ8sziBgDLJCuZJXmhPeI/oBR/aODn76+rbngEX4uHo7Ol9m2Q3iWikeTj2vbg+Z9wLgBhiu
0+fLoarlyKUWAxxKlrQ3KXbWuDUSMiZki7c5EZikiaeiPpVnJTPBsYQBjIkaW9KDbOupWlma+7ts
1hwbQwfe8Jl1aJpLuBNB9729xbbMLiI3NUogm2LKP1YHgDAqGSIuOFw9RNY8Oe6DL9YPUcQiDMHq
iCL6FLtcq2fefJOHS4LanWUX9L06Ms/UfzIgLjk/1LBM13iIzqbAf2rVcm3Uxgx0ulMhzKlOwxUC
l8nth1/UinjSGzMNTJsE0lo7DYq6mH9SCCbrdDamiBauYVb7bGfZ2XMU0w8kZnvabmRub4FIIJJH
4EmNMa8HdBGkoYiWnZ+3S3lMRAGfs44ajZqAaaB4hK1iZ32a67R3m9GZZDAqkbdB2pIqpfNhwu8Y
elWdlCf7HKpGD6d8o3BHti2pWbysBvAPhPwo+Csu3xriPFL6+0qFTSL38YUu0QjKQ/pzWzbZd0V4
fLK9GHoGdJcfFbqRwed3KZsWwHZWySGdjBx4MLSPtKqahZjBq8DyqC/5xP+e4rlQZ0iynV4ipqMu
8XQDgti0/yBFxoOayx2g+uO3MyZPJ0ExR8JFstP/EHdt2t1V/WSMDtycM1QxUDct2qUQ2hUXhrDG
157FHUt4tSJ22i0nBRimbKR/rKsyHeMGlpLpKBT7eg6ytbVBH9ievZGdmXhjMjHnVgskNAUib2yN
d3LLUZrkYm8jwRUomzHPEbs6ChTJNcAv5MhBVJUHLMBWcj9f5wY6OrEc9aWGJN94nW/9gJ6NYzlp
1aZfey+vGa6krEZTp2YEwafWSrrOHjerk3FWNg2IaKy/ph3iYLQD3FZN89tQKFuuuG/i/zCl6QcK
yg8+UET8uJmfiHrFg4Q4Sny2Obhx870e4Mhyt9hmGWHPuaYQcpzjnqldf3RSMu+L01umLA2sRbO2
Gb0+SWf/7mM2YQaWnXfGbP/D2MpX5LHMOpLtFPo2G1XqejC3wp6/oqJ9DDkTztfd5z3bd6TcLyPg
DPUCH8VFjDG42zRC6f99+MauJhE3LYC2aKf53ff4hq1jMDo9Zgz29ZX57meisDszZartq3avcmWO
6iGxWDSy55QBG9+k/KXNfkFtSPbm/nOy9BNQeTSyQoqzJHc6SgIypn1/QcEUMtm2L/x6Wx941iRV
e93maZacGZSostUst6QgSKp0oQi97E+iXZZS7GFjhnN6TjLTNCslX0HCKonY2VcPl2Jt8plfTPhy
8Q9MhTOqV/lvHkmxjsAnw6og4chMP7Y7nhJxP4WDmp1oNEN5lD7oN5HCRyJxb4IOfKFuCHfTtc25
pXjH6s0z6vuXMVj6qLpc+S81YhAMzI/MSmqP7Zf7j3db6CLsr/8SdxhJu2bbslY3ye1KEE+J4grd
iXHWbN+j4V+dx/vr0YqtF/u3RFeasqohWbHtWVsI8G3zfj/gB9HDaehU8AYRNS0UvqfsI6ntcLju
cXKBwgcAJIju6Tr7h46j6QtmYfYqSQwDN8cPO0s5rg50oRMVAMmA4qoYDk0cFsn2mcj2EG7ncsuc
Giy9Jxm+TSAuAbyuQaMbvUf0EB8sFjjveWIyi8Fu7o4vOwqGxiOXz84bOSuE8POd4oRoFkmMqAGB
4+nzICZGC3cF/fhrq3fEVgMqtfTixD41Qnx9qW/TcBhJIeWANSs21lT3VGYqzvBqXIvMuVZ8pdNn
yRB9WXaTY/gMhV0L+oOE8PYiIg14V5ubrDun84A3I2VnB0xrSMHAJds5XitRXQhIdrYIZ9AVtYd+
v6Ez0R4/uSgHED9Y9lV7L/GT5v0el9362uR9DsZ2hA9EYcYBwa6TqjNXTFiQNPYag6PIktcXcAFb
dCEbGZHGD6PEza1fe0h+zW9IZs//jHy7+AtfP0tRgY5R+6heZRn6No/+PFIptswo2sLJ15Rzfb8n
fWlAZOsMuLDdeLyKm8Lr/xyMYZJjR3aBhKmzqA/l1bJdYVqlTvCNXU5ty389g2rA3hAVmik4CudT
9rfbkfZKxIryLfQvmD1z246Br+MPVrGPwjDSHfIjyiKzcO7yzM2pf/Mhf7nXz5vSFh08xE0VO/pO
xQrYrzVfRhBl+UcZN6zns9QqeyKgkpr49EatOPU+z66j6C0CY0zUfCwzzPmdNR5SqKwGbVnEBFox
p+11RFCb7LK0LFx7TC1WaXkjdlAnpf8GrZ80qiCXhMWfrPT0LOll0FWoqT+BBS3+miqh3vn262QL
CV3la6UbOpodbOoyt8rip/YEEIsjgrdlMZ/TxhnghlGbh0l6O2yrusYAnr4qQO9DffRYiWa3x2Ow
LKhnqdy10iZPbl/dmZcjdzOi9sveHWomztGOTJP/qwIjU7/JkMVi2rZPWqOK2Fdqe340q7+LXzly
ztA+8LctvC0mvx5QM6b4Ku0NH364awO7BfRXPufaIJC0r9/THHNN/3I+O9NdxKF7dEMC3VOcZLzC
BGH1Q+LqY/fp8tOtFt8+slaTPa4FCOZrWAopzdN527dGgh07XA+zTHnIrqV0NrBwTjZU+BiaRF95
ctwigwlmvu9X/PKLl7vzZ1mwugzyndz4Ga0YlHbWCrxG3zt8cTTTCWOepfrm+m+pHxi+J64qiztN
38Ea5fcqBWfTEXo8HFPQ1NljpdyUbS2GyeIxvfTQJeAKiK2nwgAhJGJr1AyVYUUfS7Z4yItu9u64
OIESPiQna/8TPqTf9hgrTSNFHVLsUltkuRl5q7Pb2cnW8Ycj0veR2LSMT95AN7ckm6rHIjDgnuL8
+UrGzRsJjuYSxAuJ9M/v7AaAu46xxqXL1sfLINftjHMAAPUI9ENeyF6PAr6wwABCz/hnv9aXbzY/
nZbL0Q63kJxwGKov8+fxmBFDIn/umV8g19DE55YeXCfCUZ3paJFR02wKsueeCIBj02vFD0/aBAY8
TWWeN45hY6k6C+mdI36yP6vxEtL+UjLfKd5g1Re6RsXdf3sGdr1GwVicabJBGbSKp8I5q80fh5zy
M1fU0F32Fbgrcw1BnKxAQriNYmakBUmbM/FWHaGvgYlf9I1zTAb9CfK0VSuKDzEYPn0ON/JhyrPV
QVBSD+tkWIYo/hWMOe2AURXyZFa86isuCK4FWe9A0QgnpCyFVugP1LNiyjHr6UYypxocIYKEstX0
MFvt3OjLGUUiaIYjYCV0DGhgSi7oUra3NXsxF1LbJD1n4ATPd3M2TZtyLaDHyUKSmbbfSvQYExAq
Oj+tWRqTuVLqgM2CCQ0ggnLj6mYcTx6QjK4yfk8lV+d/oWrCzo9RhuBk/QjkSvl4FTtsli+z52I8
y0HhhmT1o7GBzIE6yzJ7eCOphVuRBImb2RIEbidc56/LCBMzV8UIOf9ReLjvQtI0Z1lbBN3aTAAP
mhCI3f+dqO91rlAO2GnzHmHuOkZlNMzRsrDN9WMuXPr5KjSvJ6F7evkB/xSKNxXLqoJ+l3Kltemp
ROG47JRQouEOGglrmQssF7qa8oweZLB2aofm3dp1mYBI3IO73vovAZw3dYdfQnYS3MWF1yowuMg9
nEAxIkW4031AC7Wih9Z6aZyKASFGaHhUYO9DMBcQ0ZQxvgu/KGGkJ8RGk5VrzbtxeKTDkEUJ/kM7
mJLX3fursASQGKrCNnGUkDgIyBaw62NxkTO0iiImwShzVfWRJjCsGX92SzQmLdRINitfJs8JYkQi
a7ybM9s/APD7J+vo3lirVI3nVO3z3jexU+aPy08Wq46DXmAP5pzwMJOPSVS5vfmcMOFhp1C1UzIS
ieIghMQ2UorTmSGWyEY0oQIvocxVQssfpq0e7Q+eTU+bfeur7i8LY0XDPPNJlwwG+YDDn6CmdwTQ
QJ8+OYS3FaYfAMi9V40Y3cxyNHq89Cw5OolFAknFaAZMj6QFQAMz7R0mqPohfoL1gPKQ9wvD5pW2
NsGmbgrAosUXc2lWxpvRE9xUXtoYu2oDjnMwKG/OzQIWG4XdCQLisUeJD8dTbJ8/rjiWVPwDW/d+
8ojA5ENyLKF93GxaOHeOJtEosedoGGJmGLJXgZSqC5DYBdaAArMcKJGMQC1BXVG8cyjJt+HCUoY/
zzVLVZHFpld7qr5BW8V3NI3COXyI4+J/yeBUv8FiljKpLdFMe7PkRLmW9qSH5ODdbFcN53+QRRAU
+upJF6j5rkewmvSCYj4l/mTb76cHYT0s9zBFlObE5SYMMY+lAaf1JMfc9lAN6AvNzShVPPLPWF7A
MmxUZSl9XVaIKa2oTrBxPzO7P/3p11P4Q2h2pQxzUEMWsUhdNRxRUdFckG3HBVfNSI0yjlVXPTaD
4hqc/eJJ6KUNnzLhMbc2dc+NRyT3aJYEzwAbsOWGO/jIxBtKLadvZ9gyyzCT5I+2zT7rzx68XfVJ
8ihEGeFl3uKE2SeIhuzkVtqDL0i7YBQC1ahJgFbyPaRAmepC89DP5RVkH1UbXri1zUViE+2MXbWu
r8As0LeI8mwhtqgneDibS2BsYq+R749KH3HzmX59jBqvRaoExcaEABAjkjxuqVkMFo1KOTzlZARl
w3wA6S/6KMOY66s=
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qWWqp+6u6P8BZZmo/i9PFmAW/+jayTQZFsphhHMGrZunhvPUZYuMe84otTHxZwfonViYryGXZHfV
gU7xIIVlSSO1ryE0qJ0NLhR5UVyc1UE/xBmMXoJ89KNC7pVaBjNhjBnxNZhzzpV4nGMtG7mNKjkD
siyn2lUK4HZzYrdYcGvX8KGarzqR9+3sOChYE3S6EIGlE46oQMBJzzIBtYfX7yNr70tWiO/J+/5z
+MnlHVBeiAe1O+9kaXAIU1ucp9JiLax8xIv0atO/3FuTL34y7NUkovIaGkoT4pTdVUwk8hFhZjiF
Z1aLhozPhIp9ZKwS+FtXK1spa1VmUTX0l/pDQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5824)
`protect data_block
JAhZvHAxewalQ//v3pS16Xl680dVnS0QPzzSODxwqnH3g8SZpFgwoOs4WC9Dt9eFwUYmx79jf5i8
e0XR77kZuMGAOgcSDp+LdcBhjGzUB1uH8NnrHSqbWkSp8hDgOnbnkAUW0Psn97dQfOw7W1ZYc9EQ
5aNZaQG4gGz81lZl0Mdm9LIK1hQ2rxAvBI6piojtPTKIrSSv9TrwvLru4nA0mq2elk0cfdU375PZ
pK2wPiT7M/L0DdxhXH9jUC1ogedrjKIJYo0KbdOLp1gIEgk6pUhohGwzedW0/7hGGDpY7gqW0XRw
aiNAKE7rZugXn6QpdmLhVzuRyaNcdVLqa6FrinA0lKEEXIYPRirLDUCt8Cqsj/fjwlf8NqUkQKgo
ZkqMsXiXG+6xXasUCxwN8B9OMaeieaJhknDWHaoWkWRHo+9eHBfHQ4/fS7QRUSFj8ff/TM9YNWTa
DYwyoIo+G5yOatYgur8yqBjW/HSqXfo6jxzTqYdpVFaoilSHP17B+adEM4dcwl+RM43glhKC0OmW
fXYjpp2M1hCfAYfJwTYavu3DQ1AX2Cl1HYqQDpYPlEl7jrMOwa+y7fVNSm4uKAe/3feJnJ29vAkO
icfsbQ02ad9tdO5ErgCqac4r0EFM/9FvZySE1vWw9o+H4GHLVVlJt/OCVlJ5jUZhw7faPUZcS5Ea
pQavB2SJ2aMBUyk1YJLBMvQHW/9UEASWdp54wUc/Bn3LptUYVbkY1W1vIWXdbRpoOuvwUSVNak17
l7Lz1Sd/fnunAkU7wAZmKs0sGrzyOr5ZROPdbKbIwo8igkMRBmKrmM1XsT/LRnZM5q1YKdbmu0Wg
OqBfTy0hrsuixJYpmEn7NUEA9lU2GhygEgelC29rQ0mQW0/gYgmkQcrCTjrcB6obX+Gqr4/uBfM4
b3oVSAW9M2VRMdge0bk4R7uWzzLNrzStycDSDK68bkd3FzsJYdfu4Z5224g4v2PvwBKXSMaPqS18
cck2QSL0chIP3aUIMLwTzXPW1hnEMrs22OtVXWk1H0qJGegwzOvYtTIUOIEl83DReHAL6MOzFmBR
pyVaa3nCzMFSOtdO9s2n9DnCjlsdQFrXH9VG+hpf1CPzTf1rJxiheWuxkJMSy/o6ipUDyCugs5/E
ruljWdL2LWF6eI8rSedysXw5txeeG8UcoY+Fx+nul/vFceEVWl88cyBAl9ETE5J5TuJU9i7SjTHl
hoYPaFWQZDSETQi/4WAEXzWpP/8F4Ro8Thy/JJWZwNxlbaV52FTtLEOuf3592u7v1w08InqqET3z
3/QTImnRDakN1Ik8pL5+/MTni8+v4eWY9tkc6df+XwREzBD1+SCvUOd1d5xalXylf4o+diZbe9Z+
WW1QA+GPYHQ8cuEpjOyOfDRChj5jOKhdYJF3VDOp5UftM47lKW2uc3PfAMc/dB2yfp8inubxgqpF
V3wb/u6eusxvhpylDh/gcolEITyHrgpT5pMRW6UKBgxmcvGE2/1e2IOBFcwEIrQ2XJkFd60lv6SJ
vXMVdXRg1z2VSAIDD8JmGtPDoByfaqZvRQeV9J5oyN/w8g+Jwk+HGRnkwgF5ESjzsORKtz/t/d0U
WkKT68cQzjIfaktfSffqwTkdflKXg4goPzo4pjFZqIKArsGzkiC/7DekrISMHt6ImpyL4jbe8+9Y
UlYrih+47wj1qC1IYo7JhABJjhrkVtoJxWqyvSOhbNYLQjtA7Nmq7qgFcVq/p5h354CjoyG+wMgm
+Jqph4BUYBAByy0O00Ms1jhFD9AHu9ob3nvrTkrvezmJbS7fNPPFCp7xLGxPF2pZE3rdTQ78TuRR
5biHV5EAGMKI33z4wf6QgdvPEHHbd8EF1//nHovr6qRutUyKebf8ewrf3E4c17ts7tDVy6C3Co6d
Y6qdgojAl3ALDs3LgO3UgRRXYPqePZnLOV3f2Ic00toi77RcPN+mKCQ428+FM302NDQgcaDwMy7A
Rz2yftCktHoj9tF90rP1k6TKyOI4sMYXAzAW4agEmzAec88Qz7ojYJMCdemSCEDMQaQYTCPOlwIT
WLYwbGCkjX6qTNeIF3N9+/lA3cQHbeJh7XdhkAPeZu+MP7Kn3Gj3K10A+5R3bc77LxdRlr65yrWy
nfk0BrfJ6jZOLp7XkkDxW50JIOWCwh9OEScFz+1vTJ1mRiuCPd2lskqsUvjjFGNwGBMJPXeYBIna
8ZyUrUczPTZpNZBx4+MmUNVaMizl07tr5qxCayhdKjFeWF/jcAYSmEgyhvbghU7yz2xWW+G5rtsn
t1tS6hUG42Y6UA4/NmllfZ+ENxyU7o3F5QIDLwH9F2wsHLftAG/z2wtK/UE5sHLKQdRfXXRVCqNn
dPdU0l/UgHsvakEkDLmOWx85sLstk6ksZRQI0dOpG/Hyyc5CntlAAc3IcI8u8GD+KB9JSr7Vjp+e
04qdCkAcjotoc9GyQ1UKxqGSHN+2yyaIXs5lJLhbhbiZSsT+z23YIg+fPvQCxSsrnbMXI3InKZwd
DY8YBnJiXHxQl/2srWNYyF9vUPJJH/0L/akiKkZPx2qq2T91tRcgJaR59VV9z8U+2gpQzmRGifpS
Hgqi4boYMWK0I1ZMFBOIBUs/RkR/XQ87tvMMKtQF81B0O5Rq2hv7hq2wJI50fPwpWm6j7mcV/bE7
sCFHIWeJuR7c+umqwFTEb9hhEggK3113jOrativXscYkGwmJVcKwrXz2U050d1a4Qa4VVhwFF0uV
X0eW9zBViZXAy7HD0RK4G8xisssUPAywQEHuUxGwR+MOU6oE0bhNssDGLni7GxpQv2k8waucRWaA
6MSM+/GLKKIKrm9/xxbSScCsBUNzU6uejBcZEmT0fwkc73akp3Sq6HyMToaf61HI2Tio1FR7rRig
DDfjh3O0MZZs6SXHQkj1YTI6yu8ThO6YqxVL3fj5B8snpA/YN4DkKaSxiaCckyExRnx+eppdEN2W
pOinBQQ4cse+ju2vg5pYuxbpAOP5D3lu81PjkMrqYXgza0jT2egHD75W6hQHB4j/qOVRILJnYbEU
I3wNiYa1OoAS1/aljv0V6c/K0gm4/rEwoW6D0E62kLpQQ2HoEaaY2PVOqWByIgZdzqxmQ/Dzu84s
HIAMweqYcuRv7Y5v2uh2m3avp2PnHWPNxGFygl5O6CBpeIyDTd7KD4PL1auUVmt/bQLYEKioPfuk
pbdGOZwML7iXtzEW3xfm+Rc9jMA6Zo12jAUTodw1B5aEh85/RibAcV5vOMEwJ97OG3CQEGp0sLvK
QlTjuxImYYohPnWBSTLehL8pirJj0bhWhfiTMO/br5tq166rN4Tj3eSheXEB/q8uMb2RlGvQw4bn
Uof7E9KIZAWvQtu9YKF0UUjridbz/s3QRQ4IpdJbLGeJLgVCA6ZHr9m6rRS1ra24qVs4C5tHcxym
RM4TReeb69JHAqfVfPi/ouWO5ebwICqjUEnEkg5RMB9RFRNqunMt3b6AT787zgH9vnaKf6Me7yz4
GI2fGlMJY6pm/XaKPfp+ts106hJ8F7gINmr10ZlCvo90VHDVZh4yGIRQVtkXzvJDdVenXefL9P61
kUcbjau+ZdE/XWCRymWgPrrG4udY9EYuhALWBBa4rwglw+UIobZyhT9z6dhol+gCiQp8QeUTjz1s
GfWpmR+xA+L4DF3yRmBEHdl7TOgrPYm0FLKw4l14ALuKzX7qJv4eSlEH3G5fO9hE97raGLKYo7gU
982SylnLLRmSjyLZqeRuFeDDo5Z2gMRgApQgweklMqm44292KNIanlrFj+SfomH3LEPwYqqdN1dY
L6lgFB9oi6kPZ5XpJ1Y1xcz/LGioERNgPykoKsLadhs8gzM5hpgf39+5CJr0QUh+9RySD7zoI71A
eCusQF7SkP3nMyure6CBYf1vnXQiuqWayJXt+3hFN5VhWYqfzcELE/qGjNGUnrWptV7YsXjqGMds
cGAOpaLH+kVOQONwHuddNU19ZaOuARJgcm1/YtwTsn2nEjTuQupdjffiXJrFqt1p75gzgXglHGvK
hXF0Byjw1FU100Wqri1mhEPLVscL14ysLGx+OIBheZlHa+gMGcarMdxaz6xMxickqWVNToSagvrY
sHdwK+l97z/jxsITN1OVQfPO7CI3aKoQdQgtXkGij/RBKsCnyN54oh5mDI07nb0N5QQuZZCFOwYz
b65a+81J7nKdilgKbuitsRwURrOTKP23VvxNvSlQNxHtYoeUusY0l/iLN1J+9JKRPonMmLzPETJr
6jKh6IthPlMhC7GtCGRngVcNEfPiVuSFVCqhCH/+9Sg67lnuE7PeYj4qgJHU3sUvdPB9L3VboNgw
8PT0H4owfuiHH3cxfZ5U7HX/C5dnvzKw44zQE7VLh+2f4G2Nhk8Bz8Bv7zAxckbFWDbtaGcEg4xU
ET/wTNbaMHOhmFmorZL8pWTcGgGhVeefpHP2bfX1O9JdfQ5xRh3F0NW31APUDcqJeRR9xUUzPsLR
DAWiFany4HCiHqcOzmiy8jgXaesmeEB5Eo417qC99GdBllpONGidDe8WqC1rumSKOO+CaDinwOYJ
QhR+lcG9uhO2qEYYTGW8XNTIDQbEwkhHiF6I5yu7CvHPVuc9LxlMDHKxAA2T9f5OjlKwe5ZcTF4G
MULvo8PE7Rl+0TORuxuyEfaJCXoyJ1wqz+qKr6MrSs132plOH5frE+A3zfO3Qf8ki3F4n7/5ctP6
BeSRafd1HZkP/2qgehOBDShTT9m+a8dY2W+6JmF/IEBkyKHfa8FrD71/00TVoU7AWEnHRVtWnQrL
1THHRgPKdPt/y2q2EbQA8oYjvs49+Nsbbt77i1zEXuF6ng0HvmOFQZpZfIYP8c6EMREMKMuDsoJu
olZResWa8BDl6PFXbnmsS+1JSpKjXJ6H88XBfS38ocFDhT/DnWHcwP2xRFs7e/tan5wPg/PXTwgI
POYy+z/m73Jxx2wPpsczWxafF2y/E65gpqnY/u8jLsniEqQl+8b+SjFJh3Z4GT1+Jb11/nMu4BLa
1nCAzu5i0/eJsgyQnD217rLVvnFhQjL6J4Ak5lH957IegpwjGEEsIETXp097OcoldRx3OFP1NJFL
M4ZOayDZ0OoRt/HoZWG5GuGGRG9Pg+bDlgQ2O6ZG0ZOyOyWrcg3AUz9rDWx6l8WdKJ/PKF1GE/3h
F2eSfKV40QibEC63A8LZdc9XSNwYNpp/evvFx189rAVHDQFg9Yx2eVe1yPG37slnXTPqIUaOUW/B
+sFPHqVu4Ft26EkZ6qLvGjB+joZSqbnf6jIEKHqUFEbFsDoEMnylh8Jr9fu3PuzH/4tYZKrupzN9
rs7+boDb8dUOSpT85dLkmnUTf2a/vMKqFoMoHMJEZ6xD6Vy6zYURKRUHwdnAv5MngV6R/d30rmI1
edqk8k1RiLjAsR7zGgMinqx35OUnMyrbQfe39petw5LH2R1ttVuwkPDmk0zXj4/bCT3wCHRB7Cpr
oEcRo+bmmXU3xtIj/MnfL5uR8oFKG3NoPjG1J3XXyeKevkSfZjDo3frg1ynOWM3uUwNgwehp/Zo4
ImH9HOL+Bw9+o5IWkGtTaJ8A3dmg1ueLUBpA9fnGqVrNVF7IR8/tqQQhZ0ym3sZhFmOoHm7wVU7v
vea2m+qCGhUbWwZg7YZmGo+kIFaFSw7yn28GvvgFUbsU2KS//aCc+w70TVskqVQkRbnx0RTPCrxs
0Mfi3/z8txH/LD0bH/zm7uhZJqa2ZCyXTd0NcLwmm+C9Ryu8MKLeFxWRly7gAwFU41MhQZXxMLnQ
+hEtDgzFr7fhgxO5iBqJ4rjS3VaPYP4NwDNzD/Bl+Fd74g31dfp37UyLGA2Kar9KGHMGU9con52a
hG9ywydt+tb/R59pvNaUmS22DMhsE2nFHTunJFPUX85ovY0gBfEwao/UNpjMecrVXMZCUnbEhJy+
oyd7lPvjL2IPBGCQCwE08BAXWZMj2dhnXpaQTGjwL1/WVGYaTtr65pR/eEiMLspKKZsSQ1VrQSti
HOH3lgZgXo/+/TBzjuiR66cOLzp23Cyk+S3EjYqL5b2hqqJuUt5xHUOw6+IrsEzX6hDJbeFSLU5l
dhqCxVwsRcQAFVv5+LWfxycHYDxHlh0Mi6QL2JMvyVU1ln+v8f/2U0SsPj6+Z5rgnuQz6xghyvsn
JLsfMODVojTY0p2cmTXa81RGSEtxv3sW+TQcYbcDkPf5EwyfORUpaKw1NogRo/BbyZDTFeC7qjdc
Gh9eTbEyNGRkg+XR3xL3SNx/6+boEjY/p9/wAVlANd2KcCLJZXaR5b21eD70RJqnUUzewDq0+lyy
ewYHxKrfx/4I3EzEr+4RmTXZ7+TTRzGL78poZvPSWAwIM28hbgchBIKxinzRgF8pDnLweujfIhkl
s9dzmAhWZ2flc5X6hnm+aw/68CkvVKVsOnp4Fhun/5fRNGCCPSpiKZYw4nbodslxTds6SaoargBm
KUB7ePOKQg9xx8fXksL8BaxYIOpp7MM4hNfeCbOZqcJ4R8m215GBNG6OZUYp4/YaQDzEv3LoPmd8
rzMJZGQG5kCVhD6UnbY7tgukEaOesF9ViVuA6/oaPInpc9eUNh3xGOcXUMvtXm+1f0XBdlVx784g
mQaE+pfq3qOT4EXWkdfs8go6afX8l1vIvXQIuHx6XF013ozpqNQrAxeu0R6W7frv+ZSVHdCooRNu
IQwDjiJ1pFMjIAjMI7LSh3aht+HnpdwXw9vfm4hqw0sQbpSif5HjjtHaCe5MKzyUnoNmhTRet8wi
+pU3aR4DzKgdDGt/K3PaHJWw4P3nGH44Z23yxZ2JcikKKVe0zph5t/YR50ZDeU+Cy7GtwP4ft0Jb
SgefwoPedeKVIvUDTBZFjfM5H+7pcUjCcJifczoefKGjlkZ9gaJ5S2a2JR287zIebmu9SbKPcH3W
M9arUkXTIU1ONzaSHY5dUcUPA0622x9Y848h9BceMMJcZjXAx/qLc0CtYg8c+/eFLNIBxX5EM0N1
SIywF9SsQ2G/i1NJLJVQ/TKesF4TU4uNy3KVSTz4ACJMBzsujbmAPkE8hKmPq2PGv+Hcn4/d7WHK
b/rOp9LYKdwz3jpC0GMFIQ6ZytTdTDgjQbOO7TQ2PUjktkECu1FTcJOG6ywXV6f/M8cHERs68Cqw
yvyqpavU3e2mqm/iXGqfgM8n6WML4lqhnH3FPT22cn/31wJYGa66SC7GLi92d7LTprgF+N84LKfL
JkYgY2qFeTkdfyVFRPFilhpMaxPca3EiTFVW3xUVc4xLc2ghNWCADbcg7X/mHwWwQPwXyg9mVv8O
YKRgImwJQulpEsoWHBMG7hwu4Vi7iMY3uOr3cZID5yFupXOnfXrzs4eseM9jfRVI/CSnFZU0I4GF
ngMponPc2W/pgRyMBcYNUSPz+7ZAgnyFhImHCEmqgkGMYbQHTB8HlmfVbs01foOoXA5+jkwVzOeM
SnaorN0pX2Tu0wPuL/3ia9phyoIdAZpdmh5RCdmWmDOqGeyBxXIvc5ClMDB2c58qNnDbZ/FLB/zz
0L/FsaeUKhnElkJ7dEjZ4SYuG3UWNbVZIMi3mBSRXtSdkLz7JXRXtHB0gmomz/hKyu/SuriUast5
KnfLDWRb9yOWH7wtra/w3ht9DEzaz764Ym4r4ogkI8D0VQznW3TzhbOQJVOQREpQGBD2iloYXuJD
JSyBov1XKWpQ1g/OEPnuONQhonXpgRVOY+r1s1r0PljG04+uXtjdz5PK+qwfQxKComBfiU1c+9CX
QMBNzvDYPTgAXA==
`protect end_protected

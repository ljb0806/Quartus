-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fY7Cq/qD6CKoR8KqYMOvQcnS8JKSou+qXiuHDiTFX+c0aJslYxH9CUf2wE7jEB7dBwfwKY25gY/o
D+4hJplNaYt0AixFnLu4y5Xmlkm3GtifJnBNmlYV+EtSAmlDima5eq+ciHJ3GmxtXCHkIGIjM1lr
XFkYrxTjoQ/fl27KksO66pOAYbixxHlq3sPnnu2JlhBdaXDFlsrbJS7fd742rxsKFOy7sp8jAILm
ofVJpimzemBDySy3VV5Weaxf1WlU6pSgsE+hXwiQuXXdPGrtunoCw7+KJQbTxxB4ViJScKug6Mtc
n1dUwO0Z8X/zcAHZQwarCPjbGT3J+C97/5thFg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3680)
`protect data_block
LO1lHIJ/e+yBQ3VCILC9irN7Pr2RVQPS35knfZAodgkEjVBQfLKtd5HNa3hsnXeJmJoA4qswB/iX
pkYGCfutHEWnm+McUKMEkp58xhhOnXWVvPe3aSzYNLj2V4HYkkx9bFk+DdJzbpTJwHVGYqHwc30B
9z0onF2SXdYJk6v6yCWeztJOQogtxCASLs4Q7+OO011ahzJGkhCKaBsXuM8559SlRZZ6fWlqpE7V
kV3Es0mhsFX0E/VZ2TP958KyHQg7OmwvFNcD1AvGNZmelIP/6c/x21+NTsM0/69ipc9pUaU+LD+u
hIT7o7fu023udavUszVLaqaV5FxHGA/bRQi2EA187LVb+sv16Hz8wvBvCGEMEIMdo3CFndyRDkYl
1x7Wzx76GbHW3MCJrI0DjEMnXX9GD4RPN9RuyeLnIzQOWjtmxnAU3wz6vpmFMZsHp2ET9YuawT7v
DxNB9UP3dOmjqOmsoCfWuS4gKGM/ecke6AvWDQ3ai0jDOX3sB74lZH/V85904ju8XtWYotcviHBU
gLb3F5oRI2D+x9gdljPzMAKL3c4ygKB6teNq2O2Oy5U6SbZdg9bbFelO+902wpSSi5CieuHpguK9
SJs2meC/QA3bfnR193yfJSIssdC6RBVcZHR2cIF1jkezl/5vg3g8oR7Ot3KC555rc/nyTOpL5Tja
Ov3ftPwt7BWk+Dk9HPOdYeYJACZMpcGmD8brX0ykEse2mqtrum5tVKA6H/OdmZpwVI9grNAhNzsI
kq5ua4t2XMedtBDSMkhmOsjnwstOjXOVX7NmGSx7xfrUGhYQCoUIRTyowK/mAsjThIovWg2dAe0x
Z2jojL1pHapRCiO4/PA6QtGQu8Im6SPgyKgbJZVNXNXwkfwJMVsUJI3aOLQvvj/Kdxx1Egloz3WX
R6UsR72gJfq/ocZ3UFLcjXrJp06ncPSAzHfAmoPONwoHsQRH2K3OfYzJhCkan2Hobij9pyR/w6Xo
7EP0OYa5sv24X7KROOHJHyyzKz5TzXTi2imq3rR0VNqyzCZtGxyrGQ3SRJoDEre+Xc2V3fIpnbkQ
V4d3xo0Pxp7Zbri7bTCsrDi4VyIGAfank1yy5OvpAGuz9kPoTXstZG7BCXcAX3K47CG9z1bd0mfc
odmJS5XRlSGffgAQHqkhVn/+IqRYEKa1qlQMvHzR3xX3z05tSLrjLGa914ePXwxecQUbgP/hW7Cq
hkKzATEjfB+/zEbdnE6pzQqudzpyBpD0cDdiyPgIMqX4eo2o54jB1l7i8DtdHwYjuKRqVhrnO0lM
6dqdjOfF7+612VjdHs0FaY0wsMxOJsoZSIu6rKHYD9V3EfPlmlk7b+KFW226UOrVitmh2s6/wW4i
FVuiMyIeIRtumpg159hqPdwlvYFRRTpjBmLduclRBplKi/qzMpXDKVui5rDDMTm8kLkv1K92uMIr
eTslQylM9M0y1JXlKQmZqmUnvKbd8mG+yXOrrF44inU+zdl3UKTJ3MEwZ9HrjQSYioWSlEazAyaa
NzaVPWlfh5yltvjPbOtfwokexkwWOqt3t4+wkK837N5iGA0d9SRa6wI/mDd9DK2KDqcoTifHwitE
Yq+/20acLdq4uF/2jeWRakr6CNxBprfStO12U6kpy6kRixokTbD7SEAgAsHA1mvSJotzJuYFyOSS
NQoPPHcYsEFjUdyb8lJZABKHcslWD/AAekW4f6MNfGQCmeh2kEWDD7mNjKtsTKUDFi7p1LUCKGc2
vLkO0IZoo4vVVw+PdH0qC4Z99MuUlNcL4RMKxbGNS6k+pjyGVR8Mh8TYXHlNlqiSWhfwryCMugVg
EYWZbhKiU7/+61mX32QdBrnrujd3+RjCdqlpzup2LVslrfu9VaYkwxV3FXcMy9sbZfy0TRv8UZBl
PQfyXjCVbzqDQY/A8BAw55WsjuGbmG6vkDLdsfrO+P2FgKFSigx5nqlPa0nlgSbB8QLeeAbz0xth
XFbsHwlbDJVk1GkQ46PgSadp000KWZ66hIyo+K568NMTC7lb0A04vdcaf01KEZVFnv6TPsIMeWev
CH7SEjBULI2RvwTlXaKKDrBzCyVWvwlY680ZrN06oAeKPMNRx53TtrDFNOQBSG0duVyeYbvlUc6g
cYdk6gLqKWxhFPDL4RdmyBxy47Nr3Ckz7hnJsgEscSKOhREonB6BxlWR7hJwBsP87q23xa4q9Lmc
2xCB6LVLiudl69dMAZ1dD3Vvpc+fRp85tbUVbKu445J+GTOq2y0Z/y5MhBujLyLTxeJOQaRypQqd
nD2z0L1/d7u76P6P54IVMULh0prfcmzi7aHC7OQ9K8YEOolf3jZaqEiuEZOEE+lO0aiHi4cyDntA
tQgz5jFTkL8bYOC6RpgzvK7LbZGyWWX4aZpI4334SwkVXQ7Mwxf9MyFzAYTgHVpx03f+2F8i4CIx
j2UdijN94JcpRBcxFhCWyf/ujxBm67kxH9e8pdKw/Gk+BEIqHgzuCHCyIJoR2VniBmU4UY/YJItA
Gy7MzHbkUcKjv1ItmcZv0q4ekMW8T2jzUKWK2Rr0oWm3oyfrGC9+2Gvf+Wn3QvNsKcT2K9eW1qkD
SZ8TQkG04BmBB6QBz1UBSeEKHJ6XxvLNxgAhYhRZcSx4OBpJo309ZogXOE0hjNiiWaI7b+hMQUqr
PnmCcXR4dvyjEqqjKxtU3AnlNyGB9qMlxqgQFBE1ypWRjo7wUOKT8euAXeHXi8xh4e4b3ZqbVKX3
EeLP/pV9rQQ4830gW7ibA36gUPK0LEW6v2ypF3AS72xgw8blQCb6+I79pye+ivkIPj61VuMd8c8s
dZnoWE1PL49RD2eBClu5NPh0zehubo5eSio+K0q7Ux4L45zQPtnS2/hgMTQX0fu/w1OR7jn76cjh
+EFH0CWVbktLFSKKeWPrXvAYOwWX4iVCZ3+b5Uk2SVCmIHdccJyNxZoxk/WXhiO2lOHqiaZ/WqZj
hfwKUEAjbmUZVXsWUSs4hdmHqdLilsvjXRxW7c1FKuCqtvdnHSlJxOq1GvmataQjZ8CRe53Os9Kx
NSKrB4lFt/1wxc1lA+9aEkc02gPmBoPlt1ZXnu1A1DJRHQ1624c568SAQ3pc5FMRFinDjJeubJgF
DqolbBRdEHCy79oggij4oFvFvBZLhQdF6HTbKbV0MCKY3F+7KQubN4ZSRdsmTtgSTDNHc/MySu+u
Oro7451EU7xrvwQHOXNF6R/wt84QaYbFYmb0O2O4cGlbD/EDFbrlmhaYfUOUrdyjk0hci22gTrqY
PwLMkebGPYrmAAa7iK5yZyrFy3p2xmozrCllleVQqzPGodxaf40O2ZpF84z3r2ntj/9P1xu/gtQz
YTXwF0vBaHnRKCXAzfwU7dDumEX+Nk0F6pZu+Qj8y2J+zLcA9CrVDkRq40ZYHpnK+eyp5uCZizBk
3rBHG23y21zB5QwQw+9kqw9bkxFh04Lniq0lVb8vSv1CN/+AdYYEbfxevDPmaL+NSqvBOSHxjuYA
1YmqaeGzl2ZPgcf6+fvGy1k3odvY8GIQCR7QvqeBPbtFeCgVfUZBGvctKKXJ9Mx7itX9ALSu3EdU
pVH3HpH6TEjSEmdvEQMF8bXvvC73Aaxd6L/B/vixPqaWhBwVJV0CYD+MJHxgwppV15MEKL5p1iLu
q6B5PFjT11yXV8VLg28jrG/KFBBJ5LnD0NGPVQPHTxy5xxNKNB0H8ceXDL+hA0RDJGhNLIIGtAeK
B1iq5z52KMUUIjf85IZ4t1XhOSqDnliktJsXd10eMyHAnaOBKeDD2LpeYuszps+N28qSYOIEMM5V
DrOiiGBX0IRX2eVacEpqQbNBUQlciK1lT32dU770ygprXZdJ1KPlVccHIoz7Zot2vZajZjCiJ3Bv
CBK1wcmG8gGuxsCbuCGXVOV3PrNX06emvxkd+cq7547TReOFC0DvmcgZZEiQFWFZpz6Q1iHkjyfe
J/NwCKyc6wHCjeVdtxZGYp3IYAKbNpD0eUVMB3/KpjmuC7w3pYSfS3Xh6U9izXoe2rf6vymhp3+f
AklXlWedF87TtGvDe06XnuUZZH8dAtS0ya4lwDbnGWfTesjpXUsH8HQ0OSVZHaFtQaZNaXjlHstB
/mH7NWSoO6VTBJUceeCe5EfaChnfVtDFYQtVsoWYaHlMfHOW51xADjsz+g8XHlQCOEzg9NddPoxB
kR2fajb9r5av6mqwujPJ+AUiW09aLPd7NWgO1fYFyes53LMnhKVgbWg7rQ+Ho1A81TxzZnHQGQU5
lUQygAfh4sP795lLPVtQQGwe2uTRmqYfCrGGkuXy3CLwBj02jPwVAWyHr0Tt2iRvc7TciYrFwems
arfPmjf+qwD3OvDw1DQKx5Stc89jVXzwpbbkeYFzeYTP/541K81efvA1J74wUYV/bYGUxV8kVEIl
YuvWuDPsR/1SI7HwVor/PENXLqWvT2Lxi+N6uHjjlhVQZ1R+cz272pCeagpxVzROC3jXQ7OKYoOV
KF1/G9Kf6c54v8UXycw9E4oVluFY0QrHTk7i021GmL2mI6WAslJTswJrEmqmqElPgopWq7huxQLe
qGgJl2V+gTsa0/b2+UT4Eigq12nYHrDASDRjFl/7dig5UWBIve6hGVhQnwEFsU5AqGGm/WIuVclI
6j+Hbx/uF619CVGPnW5EIWVr31a0KzziB5FrUgQeO7l21wqMZ+FE8SGuySgkaghvEBb3pKUITtQ/
kICVrkv6+llDbssxXvcFfSpMAPsLw/s10/yAxBtTAdyKItefYSOvlAEmJTdYCVRlJq7Gvn+IgnpE
KhGCBVhhN/7I5CUqrfDwEzVofVfp24xgk3kXTiL+cqBB0eqPmVfklK6VvrDBwrMNryugmn5XTuzC
m8h+OvzZ51PAhzVTuebJx7lmbNQlKr5z1+UusflOagI=
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�BE��C�,W��ܠ�p*�v6��A��"����Kg�����4���YWs�����9���㡳�.���|�p��%�h\'.��,���C�I�,ҤQ���`���>}�ƚ��g�����a����M$ ������Y�O0D��U����l��l�4F#���m�&?�@V�>bIM��֔~z����c=�C �]c�By�W��o��!��*U�L��.t�o�D$~D�BdB��#'s���$���-���Sk	5U�#֩��{��FZ))Ð�˙���leZɜ�`j���ɽ���cr�#ٻ.�x̹�����G�#�`Nۿ�&��_鱻�~����>���n�AɖLim*�LrΟ��[�1��	�C�����|ҕ��������m:�OPoq�G��%�_����y9�uo�[���l��J�a3:O��6�<��K_mst���xaA�؛h�	I5�ۀ��hg�Z��Q[Q�7-�S@���74�Њ��^�����b�x{�ǝ���|�6���\���ɓ��=+_uHK0~ ��홇q��&���r�؀�����}\`��O#��S���Ϯ�|��}�O4�����sRZ�>�O�?W�4t�%;i`v�Q� �ܡ���)��qeXE�U���w��L}J���V긔��ywj�4|������f;H~~l�laN�Ap�(���|avؓ9V>�L��cY}�$O�F�`����z(���aԊ܇�BM
��>�&R犵�z
��EjrB�?�m�_\�j!lʟ�o�5�'j>�?L!��ց���ZpkǙGR쀟���h�i�g��J�
�P���ER��g�߁����Mm쒬�u�2W���rLj�vz'�d�ll8��?͚��Ս�$�h��[���ak��P�rE-����=��nx��)\"�L��[,gvd�R�e�g�gx�C�l'|財����"�ٹ�	n�\-��|)�Kf�+}]N�N4hp�i9��4Y��9�'{�Tly:M�� bu���6<	�bP��׬qb�Y{ЗF��u��b���d���MK2MC��o�cA9�P�v�I�ɐ���G���GZ��z�k|�E/�z�-6�� "�����=�Xm��S�Y�f�ϴ��"�� �.M���=ׯ�qn̏�X�#����H�,�:����y��������u����<���/�j"�]z�n޷��`n�+�S���0�d�7�,a�ő%k�}
�P�<E�+]����ǽ��.*5���R�1BV�p&�tA�Ӌ؇U=�ɴ������)'����������LK��L9$�����j���h,�4�I�A6�>C�t1� �V>���\��͈�$�щDQ�2m^/^K�R�؎�kvkIa��J�TQ�������RXg�6t�Io������������/*Yצ��Gॊ8��|y�1w�ȥ�&��茀�Z�<�b2����˕9in�%�׆�"ji }S�VQv��]�5v�K��_S�|�8! �7y�������Br6݅#��z�Se0��ȧp���^�&�q{`3�!_���]�K�w�F��ѷ:��HÀ�
ݹ��r��z"B���LcBد��p�\R�}}x��;���Ծ�c�L=����f�4�x>W%�c�E�E�����T����q.�'��åm��0'<.~�?�����\-|�X�b�O�#�Bk;�&_�d+�WY4Z���&�5r�.�4wKk�#u�l����y���lf����n��~j$G`�ib�Cs��\��Z��(�K}���ǈpB�[�7�[q�ϴ�d2�&^�IW��v��5��4�4�^}���Û�����e�[�>�|4�3��<L�A#N�iE�0��1���ʙ+��C���F���Wv-�λ��Upi�1�b��u�!�����������@1>[UD]|l�:e�^�b��y�� �W��F�i�.�z�'�t=Xf(��mv���g����4��^�2N�:�J���^��䷵%�����8nQ�a�C���*/������iz���kţ.�jF/-�i���\:Z�M#�{\t�d�2�5ڮj�A�5�M�]���\ �xھ&��"�p��U�}�Q��ñ�4�k����e�����+��:�����n������`[\�d��+�ž����%9�i�}�q��!׀��|
J�oғ��Rģ�<6=٭z��l>�dY�r�X�p|��,Z6�+�WӥG-Hz�-�*>7�e�����Q���J�����z���6n?z��*�y�[��x��s� D@o��Y�*�!$�"^amQ����*������;t,�����(E8��=�s�������iV)���Qz�Z2�[q��n��e$,�`킞BOSab�E�\����
_�����Y��ܷ�%��b�J��ܸl~��
r����ʯ��P6:�2�ʴ�K��s��ۂ��HAjOj8V�կ��HP�?kq�׸3�6/?/E/��i�-.��{��k��k&���U��e%&\�C��.��(?��!�i
��h*N}9I�D�/?���G��l�MS��UFu'*<�<k�;��4L��~�,3W�au)l����(i��`�'���ZJpt�w��P�ʘ��e4��D$`��td���5��jS����8�lȒa�=!7�]�B�����E4�}�?'!1X8�"u����Wi~2:"�wX�`pԛ��j�ˤ'������Է|��H�VH�Gt�V�n'��mXo�u�b�W�����am@*�l�O�}��fw��C���Nq��k�WV192�C �sߤ
uQe�S��B1d�5Z ��U�5w�=������j/6���� �s'���JIA��6q 	�e�G�Rv��7�`�6n����Q{P�����)_mr��D �ΚaQ'��b�,�NE?Q����2�ki3TI�H��\܍�0�����#/���f���\M����]����?�ȨH������Sdm-(Vȷ�"�u��$�d$ط�"]P}����\���^�h�x��6%q����&������8K��(ܩö*+H�Jv��y.7x��d���˖)B�X�i(g��8HrK�	"%d�Oޮtm�#F��}�wq�ҐOs�������m�������6jTۢѾg�1�����w!>*
!��b����z,w�:��:���&������v�@�ְ��z�o��T �#|�Lq��:��Q�'�d����,��b>��@��{�)�Y��s�J�ʮ���ƀ�G��������h���)���&�N�?�a�r���(H��+D1�O��h�u���
a\l��)�0�6DN�����zkGt��8��R�����{���-߃��#踁�)�du����lڑf&jF�����tD����3�8��ֽQ���NM&Z�vٗ���[�m}�>{y�7#`�h۵*f4�G���#�3���Q	DtT�gRzX/�j�n��Ⱦ��&Б��1L������ܙr(�����ք�T�iM��Ǳ���$Dt#��q����N�i��'1�J�����vbmr�r�[�����-Ь1���%ܵA��6]K���?� )�0���l��`"�S3Vm��%2(��?Z�Z8�J1X�j�Sse�Y����S��Hi�e��Q�&I�4�;�7��1S`PK�9�n�P�}y�mɋ �MK���tt���ս)-���kG�����hl\g$
r
\ p�S~��r��6�/1.����iK:�&�o|�d�^��:!9ۿ�	Y�9���I�(�t���3� �n���.�g��[b����_|����~c��l�ţ=�� ��<���4�!�sG�������|*���$�~{�G�/�S�a��h#zZ��u2�Y(2~e���J���D>EG��α���r�b��Q����ހo;U#��w��i�׃]۳>�Ҷj*�gF=J�{̕z�3���\[�3z��F�ȥBb,h��8�:�}�nk�?���}��`�B@5Si�X�
��ĵ��1������W?2e�����ټe1�<  ��[��Bq݌������P����&���6H��v��^�w�?V� ��s���t$A�-���a��r�ӥj�Q:�D�m�R�l�� �s~��5�����G�\0��z�)������doBs(��e�) �Y���9�Eއ7��J�^߉L�5�	u�Ȏs�.�R<s�'+������١�Dюv���
�<����oP��T�J��&�@�r|����(�ĺ��8@�QB���_-�����H'�M��w�t��(Q�g��V�>��8w%�JՇ$$�i�*L���?M�±9Kanb��͸P)�<�F���e�I��חC�<٣���ꑼ.��AV��k%+h89+n~��Y�H�Ƌ���I�ӫ�.�-,u�91YM�O�&x}� ֣S�5���T\$���X����r*ʻ.>; �'½mA��at�x� �I�?º�\����[s���JuƼ_��h� ��s�r��c�$=*z�BRu���O��g���}�װ���I�����_�QL�u�U�h�(�l��Z������������|�L�d����IX����.�#F�f�H�Aڮ(,-9%lE��@"�jh�o���� �qwX�h�B��P���u����<<T˻��R�������?�䓠E�A�꣩��+�:+uCs��ٚ� zs_$d�Л�@a���(�gtZ�k�x�l�V@�)f��]8��U�D�Y7�.�Z8yy��&�B�k���#��r<핱)�%-��M4�2	�����w�"	�a�H`���=����ғ}��c']��"d���K��c�����"i��kj��<��w�z�=��^_�;�8g1��/�%��[[Y<Ћ8��W��P;WV6�+�	(�_y<�Z��P����3��uX�R]�o[V���8���S�U��� ���Hc�EM�z�ۘ�/�ӫ��(�\cEґ��^�;ñ	��	6��jX]D]DN��9�<�M?6wri�85N������\R�T��2Q�m?���1�?����-���:`��H�`ɓZ1��ۮ"����Y흍B�����+�r��A%���5�� �\��6O��}}r�ކ�keCK��g&��0P�q
P�7ʢ_��a�|�$����J�O���*�<ζ�xc@N�o�w���9 �I�.�+3)��4�c���E�+���'~(�1�DB����uL�3.K����cW&�yQ�Ɋ��X�B9duv�\$]�ɴ�;ڈ�e�
G��3Ӟ��9��I��O�oL�T<,KdiG��6�{��oh/u�*u��z��`k1�g
�xE���8�n�2�O�:�Œn�`풯��L
Q�������s�>p||pE$IC�*�2�6��$H/�����/ӤGʰ��E��̋�]�FZo�J�	����T��B��#���헻,����WzAy<L����/
Rd��_�o�`v��ٮ��@1���������j����<���&C�)��n|���RZ<�^a���Ln�U��\\�=���9&�1��URzk͊	�� ���|�
A�Ư���;����L�>۞�,��!(�C��
1b��hv����_�i�0��af���O�Q(
�~f����S��{1Kq؞O�;.���w(�m�|��eڗ���3��ϳ&���U�7f��L-� ��۶lΚ�L�Rnl��-u�6��Z�h(��?�B�K�yK|5�6�¢������?�x �_���&Dpf�e�q��a
 V�ŤH?��A�oX6��\h�X�����7��j��B�G`7y12���@e�<��;.� ?Ci�-r�ՁP�!B�_B!
�32���-o��@[�'b:��O���{F4��Žb�C�����
Nl�q�;�Y�g!�7�`�f�ɀS2;�ٗn���Ğ2���GW�gQ�ˠ�Ԋz%S�~w�q��-z���7.N\��!�w��%L=m�f5����V�>UH�6�.vF�	�~n|�'�Pk���\E>GD�]��"������a��/��'�P�$'�_�)�_a�4�xL��οG�
��no�_.���DLoe��y�S�
���>m������9A��_k|��<�s�'NY���![F
�XK�j����]��|Qn���f)*ǈ�`j����i*����G�D�m�.�A怋x�E6���O�D8.C�'�(B8�فH�j�)��~��&�"n�X���Ps�8Q�žf�ݧvQ��{Li_{ ������э��0��D&cd�7�W��jJ�=��n#�1��9()rl
^ƴ��U��Pg�L+��,|�|D��)�(�f9��������
��D
��ݧ���H+�|"1w�{�	���nt9YP��i5�t+�E�j�E�N���M�w���u����Ԋ�$ͩ����9Ho2��g@�>�&�~����(�b�FY�{�M��0��{_fgT�X0��J�<FD�����=��<M�J�����WP��eI���_�◣UA���6D�wQ��*�nB�T���ߪ�����T���Y�8-<�����A²�{gJ�����9w��:�oD��a�}4&HQ�Ѻ~� ��7}>��JO�+���c�L`9�w�5V����B)Z*���=6n����s;���!� �=��Vd	�K'��������p�����My������-�.blϩ`8`E���e�*D�u��kP�s��2�?��Z���L��T^�Y���KNQ�.$�~^W��!kʗ{ٛΪd9�ӆ���XL}_o���҃��n'R�8J���^>��A��@���[(8E��RG��}A܀F}ԸEA׼Dѐ蹳{���,���u@s�T�II�kh�����1�c�6SK��'(ٻ%������qn�t�)��z�Р��C�����7�T�l�W&ޤ�!]��@������~����B���$��kt� c.<��?�+k���5��:�8^��-ڙT,�ܵ�4^����M��کrE_�^Ckq���ϝܲ�6	c�K�j�+*(���*�Y$�>���F���ت�(
&L���V�R�U����Z)��w˖��w�T��⡙�����b7��D-�ϒ��4X�qbm��A$^��}"걎�ޢ5���4�*"�"�,���틐�>`�EO4��3��#��1��M�ѕ!.m�m=��&}����@+�6˃?�%-�Q��o�愽<�B1a32r�ęm��P��0�^���vt+lMA�}qh�L�ܑ�Ӯ'\��L�{i�OP%�*þ?y�k�]H��<�8�ۺ�f�zj
�oW���N��GP�������Icy��-�����T��Дb��gg�Y)�k���5"ˡ? y%l�f;T��0��0�I�o�z^0U�%[˶$���7���]�ƥbN�P�0'�~9��~
¬c�.�Ia{͌�����5,��Y�M| ��_U�
";F��!�ԣL��oCb��n�N=�w3�cx�b��a:��^̪S3��ء>R{y���4S�*N�z��)⇄2���+[�1!�\2�D)��������oo��,(Cm�,)�Y�������n�>�B۝�48a-�4��8�������qB��������y������g�_Z[�;�p�t���͇5�o��Z����3�%T��ٸJ��ٸ��U>,�-TA|�>�]�����s)8�sp�u$����A�pj��w51Exf�=�"���C��<��\�!�-��T�K���bH��.�7�f��e;`1�Q��!
�MC�Boe�'�jM�)��YB�;Ӵ`by�@x��-U�
|�L�{�p᢬��}�\s��x��ݫ�oY��4�V���x$FJ7sI/�a���8�/_>��y��:Q�h�"��Ã�9௜�l*�V������H"J�ΆlObx�W;Uf|&w�ճ��|Q�(�J�S������FD�x8A�V������j���I8l�8Α�o�i�B��y^��	ɓF-��0ү
��*�F�a��L���O�4]7�i�\�D�֯x�=M����sP��2�B�5|�|/�m������_>��o/� -�� �� H�vG��'��uM��U��N�3O�X ����HqxF%Yy�!8�>O��(�KBz5R^�n�h���t����#��Fc��S=?/]���x�sx���� � ���ruz�"�04]U�
T� �~4�ϰ��E�,r%z�]��s��Rυ?��w-����ֲQ���)lq���$GȺMG���@�,/����RhZQ�:��S$
 uM�ڸ܃S]=� N�XO�AB!�_h�Q���2IX�A��h�'(͚kģ�:��OG�N	��"��fv:�A+���;�J(�G^K�)V'�����M<�r�/������-�a��ܷ��1�,���!D�'Y{�&����ЪD��;?D���ԫN�$^n�.�I��� ?ƹ�8�-��뒪͙Z��Yb�x�R�g5��Ɩ{1��rn̴��a���_����8)!��k�Fo��K�P�'�փN�x�X��wz-�������^��4xY���MyRr&��0aX<�"A�(7	�hbS�5L%����<�,8�GU�k2꽴�͛1Iϖm�a���y4b�7l��g4��2�g �3Y�c�ta ���2uگ���+�K��z���挡G�%%���Q�+�x��z�0D��ECj�v7��#��U��{H�gX`���{r�k�'�(r�f��%V��3�7C�{,�do��kn��#���{���^n⣔ߟ�m ݑz����*_���G^%�?$��!/�sG�յ�E6˦9�V�I��M�}����A�t���!�P�`Ǔ� 1���¿�o1#7g�ĺ%�jņ���,�����:��U6�3�3d��56��Q��\��>���+�AW'��fGXb�eN[� ��'�"�3��ّW�K�N��*�b�WYV�(@��Q8�\�:+{��:���cz��Pe��	{�8p�վ���g��5_�k���~���&+q5��Q�PMS)￞�ل���+���U_A��wkۈ.k<��C�gB���X�A�ᣃ��?.�	AHs�jYP��S�g8���ٟ~�����sD	��4������'���V{#Q����]��L�|WLŊr�DE�PE�=K��uIg�옉��D�Ҹ�dl�SϮ��/��x��R�
6<FOe�v���_�g{��z���Ψ]~m�\��B���b�X��%�69`��Ha�	�	D�	h6��t*�_ ����y/OUY�t@[�m�O8�Ү�(�+�.)�h�6��Q���f�&MhP�r/�5�9-m����7�>9S��#ݲ�B�Y��S<���%n��M}7��^	�(j��I9�4�2���_:=i�ƕ�r��i1�ů|	+य��=�2@D�E�y��0{S���p�E��a� �����U�$ ~j���V(>��@��]�D��-e��ۓ�jD�\�!	�%�^��-�o ����q��O��D(O?���+���WG:���G�����t�-�4zUdCH���� ��K��C��U�ao0mֽ-�z����~j��]F������*NQ�y�ùL����L�?窃�� ��⇏���q�}�)��Κ!�#w����$Ā�=`��1��x�1��Y���A�
��E��x��ۋ7V��_�D;�<!�����4R>ʒ5��+�2%SV3�>�����U]�L�З��تp�@�x�����#�{�K�C��"i�s�E����=�+��vIT��C|��8�V0iJ��F�R�(��Ι�=c�) X���R�1�g�9�&oˁzׯ���'�e_�ڝ�Efp)_BR���Ο��;>�ڛvůJe$2�]L��o�j�����I[���;��7�b* W����OUwK`�h�Ӊn�W/K5!5!�:;/��YB��.���aƯ�*V�F�p��g�7Z�ٹ9�X���S:�/���L�������Rg�)|���θh!��	�fn_��8��Q/[5�=~؅�Bp���p��A����g��}�nM��f�:���8� '2���J@��
���.��r7�>N&=wZ0�-j�f���ytn���ȹ����Z�E&>�g��&3d)�	�T.�F��@���I�g?���`������ �,���H��5s�ٸ}/ ��7Ĭz��;(�^�6���̔�(�؜���i�[ݍHv��m� z�I����	l�M�j���薑�ҼXZ�Is��죱���61���g��ܯ����(��lo+��U� �Z�G�ҒU#�8�{�(��>��!z���, B��n �r��~���p��:�)��n՜y��sm0ͪj�]8_�H����4��@zBrL�gUVڍZ��vfx�&l4�X�6�힓N:k����ј���\����V������s6р�ZV�{�7U4��W`D�xN�0��$���_�*�����X��$�/(��5�: ���e����
��j�2J�,�`]�����L��݀�6Y�|P�ן�ݜGo�����x=,���R]'jO������@��}��9����c����9�R`C���*ʑ;�L�#Pb �0��G��*z��Jy��z+*��Q8G�F_[���G̡VVڜ� �u�ۂv�ȎY�E�b���L��w)�Z�b�\�AGvAKf��7�+7�9nH���eIa��9�g����
B���}P�[o�F��hHiW7��S��������b��� ka�4�Q|���r�O�P���g���F�����0��p�~9�
w���䝍�#��M�^�@��\�@P�_C�`�h�$BQ�* ��C�|�p�.M*Ԗљ����f_��՛{�^谣\��"��H]��*�t�@����ϱ�9���|72qj��a�I��1�+#�V$����t՛.""��l����,w:��fdg,Ѡm��g�H�	��.^W�>����z����Ǫmk��1�.FnĪF�$�HdP����"ن�	������W����
�u����/C�>*�:KB�gp�O	:�� ����@��FI�_�������	�S-�lp%Ր��b�����p�Emh������i`]��B���N��ԣ�b\��!0:�,����_i� o*ڃ� ��N�7u�����!�L$�
U�"H?
�H
��X�L�	Cdǥ:ce3�님u�	aG���7mrm����9��ʇ�T�`���T���#�ۜ���u'^D�?(���a�>o��=W[�Vu��կ>4#�M���4��2�	?���%9� �H!��8�zo�&��m4@d>�_��­2Lx���ȏM���q�<�i?	,v{=��:(h�!�Y�Ԇ���J\ňHّ�{�s��tLQ�6��=BR�5�m^�p����t��_=�L*b49�8�emFQ�_�.� �']�n��@��T�-'� ������xI��y:�����YL��`�,�I���,��)��%���:ɍ���+1��	��&uc��x}���v���<�FX`qN�����j�t�^~#m:#*_֑Ve]��`(�n��W����H��A#q
�TU��������E����^Յ[�t0&펿=�P�k���_[�����;+��|uj�Z��qh-p&t<�|�Em��"��@�Ei�6Pˍ�,;�2 �1���j��Ā�e'�Rf+�߼@P�~6���r�b{8[z�) ٙӂ܈�>���]v��P�d7�+��CdZ����|�T��dޭ�Ė����tBc�P"��&i����=@�?�RЂ���E�0$|��i78-��O���2#<�� ��>��RM�<=π�$�_�uXE�1d��VT�ݳ��@i��}F����Ss#nB5Sc�5I�����o���=XE�vDsM��<+�����6 ˄�>��}[�yO�J�%3)K\�pр�*>=zј�$�x�A�AJ�we{b)7%i�N���é�E��i�\7j\ݠ�;1%��Ӵ�,+ѭ&}J������{@����_W�Ǐ�O�?-�1�W2��'���\6���^�K��c���y���%Ћ����f�Q{�gj4}�I%6<���K�t�G�/I+jF٬6��L�w&�o�ԭ������M_��r6:W�O��)ʂ�e5rn�?;��/�)}@��c�'^��T*��~������v
��:Q�>P�C-6?�C�F� >�b=�L]͇Q{�D3�b�T���G�xǱ��"���9^ԙ����E�n��J�J O��Zo0zއ0js4�])=��5~L[E�`��	���C���]��e�L��P�4�m�pV��~����M�(�^�%������(���̕2�ۓ�C�����x�j�������*M���z>�et���~��9�e�tٱ_A�O���юg4���,8>��Ul��8W�I����m��L�J���܀�jb�ҧ�.����T���:�L3FG�G��r�}x:>?�Ftd$��R�j'ukv��+���3�Q�1��2�̳�P�2.IaHPI�>��v�T#����Ѕ��8���\���!W��� ��5�M��]���1��Û�}{*�y�� ��~���;�K��Ô��k������&�̹v^c+JA!q����b����L����nơZ�NGMۮ�(3��%�Kg���-�u2u�C��m`z#dPF�_�s2�g���C���ަ6�L�>=�j���?���pP:><|�[�X1���ݢ�aU���K܎�����P�
���R����Lk�&�j{Т#OF����+l�b��6B+J��mF� ���G@���O��@P� �$��3	$e���Q��ueg���|7Z[gt��ZM~	�,c])����P�11��g#d�=�ڶ���t^%�[.�7(ʞp�@/ݫ�uP=8�<iK�N���<`n�-B�#΀
����i�j?���=t��6���)W��2y	q⭯��<Ks��L2{qߕ
i�
Ol��Aٴ9(R�����x��\u���ܭ���^����T�1����U?�@�9�� ��Us�I��J��j��;�X�-�8B8F�(�s=9�N�o�Om�SX�P�⶚�>R�zݳM�$"J;��Redj�V���ًDcT����ߧ���=��s6��ּ���{W���4�}�L$�"{O�]]����g��ma�;誠�p7�+�es���O��6�O�t�+�����͉KC�Y��=&�a�Ř�������"CQ��wQ���yA�g���l{q;*��y�fOfcZ�:J����L���c_�S�,k%�F�_���f�Ԅ�H�&�i�VOsǘ�D�u��~3QU�
�]�|�ɍ��[�82,-�vɿd'CF7���P����=(��]�zq�M�}|fEO�cg�f��XE&���2J�8�>�v��S=�\N�;-��tb�k��crE�3L�8�G��u���������'v�����\B�������<m�c~٦��ᬩ"5E�V��Є#���9��0��~��#�����_O�X�Q=tߝ̈}j�)�LK ���q����P[�F�fwz�>c�ߌn��j�*X�(}�-��s2!w�o�GI(�CLۥ���!]�M�JG���f}Pח	\����1.p`��+��\����,(���
bk�BHC�8�ܱ?2̖���1F]����w����޾y��� \y�Vm�Z�΅�sP���)��`�8>	�T�Ð_�-ނp;?Pt�?�/+j����7���|��K<��ԛ7��H���OZCs{���C�����Uq���������hJ��A�Ⱦ��ib� �+��b�x�ytӸ�
肌�:�kkpfs��,|�B8����yb�>�M�=Fg�T��'��!� ����uD�2�u��j
,$��Y��AIX%1�3��ԅc[�`�ʰ~^�x�uq��&�b����"8��L��E;���bx�'�u�$<f(I��u.����{��Q����|�V �Ԁ	w~jX@�$ݧ�n���]x�%���[i���|�r��$��q����� ,>���l5]�G��A�WKK!QZ� 'j+ޘ���ۆ\g�W�.8�~���h����+�#�F��m�>��C|2����+�	�+� �΄�Gy彤\�P�k��<f����g�J���EM�C���'!�MuJ��#�n[*"8��mY�k�����!,$����tN��r�5���z�Ө���+�T�|���j�z�Œ��9��$:����3���M�v$p����YC��x�o6%q3Q=9�ޓ^�.�����іH_u��Z�Yꒆ7gČ�ؑX�8�f����茪� T�P�-�1щ�;i���p�������.�VY0�ȧ�ֽN��^��q�V�1a=����d�p�KJr�I���\g���.�ΐ��H�A�;���
�R�&��U�����y�¢=�V���iv|I֑xZ�
(R|*�@W8[���<.�9�
J�`:���9��G��]�j��@/Y����Ψx��+Ng����4��^�2��OJb���ɮ5���4��D|1��"���Wd�������I_E����ؙnb�o�D�7�O�]F.��U*��N���M��GQ�j\W@;B���;�qV��R�	�+���z|�X:����뀍��s��{P��b�W�ښm�-���Vov,�c���&��gƇi;�V�<�~}�Y��E"kA>	�0���3WW�J\�s�`oJ��vo~���!�P�L���%s\sU�l�`����q\�D ��f���S����,����P�����s��R����u�7WP.�"�q�)8C�1Nk|t?�1g��YBۊ���G Kbk�F���C>�,���-IXG���w��������Zɇ\D�*Ily�	��{˘;EQ'�#��+r�Q����I�X�U��]�^�Q6I��y	<�sd'�D��q�ZdU	6(pT��нs��f���']Q���C�� *�������F��F 51b<)Y�|�J�@L�	����3�Vİ����v����9��`�������f^�f�i��O����P��cH�%R��D:�9�Z��o25�L1�8fL�%��)��M��X�_I���N{��?FK��؞g�k35j˄xR|��� ���!Y�����NRK�
�?KP�������1�hO�ZM���	H����, �:v���HB-�25q�!H�ŵ��P3�w��x"h1��M�����w�Z�e@�� ��3������黿�0%س��(^֓�L�3�������1kS�2cÌ � �`�I��z_�@ ���Z���q�=��� �NP׻Gհ��`�PRM�������Dp��u�hE���jv��	�;��}�O"'S�y���x@!i��Q�ȴ��N�g�������u�j 0�{�"�M*1�h�2�}H���E8_��~����Y��������0as� 9$��bOʉI��t���#��c�-0 �G���4����:����W�^���xcs�v�1�*�q�A#S���L%�E����|��tZH�|�$pz-W�m�ꟲ%cS_W^_��Z��XR��i�/�k�g ���ZT4�dd���扞�9ET��U�/%��v�h��N�Uk�۠�L���2�,5�B
�9���f�D`v����o(�Ջ�;z�[��`����4#�Щ6�P:
���{�a���9���/����c�&�!�����b�p��@����1�č�u�'�ɛIԷ>�:�G�2�6^��<T��Be��.H��YdL.�G�ZQ�wK�6yդ����\t�|#��~	�ר�44����#m��ѶO�}�-�C��ȒS���e��J�z����Qz�.�{eݳ�߿�n��K�0	��@�J�U��݋%�1�K;� y��w���� H�Nq�^j�=��|I1��"C"�hJ\��ըi
cӏVey���[b��)=�Œ�����\����x��S�.8�&�ncK���q�-�m����}K���K`?/�W<�06�qD`��Ç����H���j1�Zx���wh���7�B�]e�zgmj#ʖ��U��t����ϗT,ͪBE�c��#�2�������Ɏ��w��������W3�.�����wiƮ�\@s���45P�*�����\�oR|�0!>h�%����?B�=�I	p� �&:�%��^�,e�L��5O�'!b5�P���+ba�]{-da�u���S��PL���T�ڙ�C26��bV.3�3��Ÿ/�P��i󵀴7
&Ȥ3��O_'�����g�&>NēC�wI�y����I��Bg0���?�ְ+mD-��;�5������?j[z��o���/�!K�GK�Dˋ��s��5T�o���ƺ0-��Xs���Q-�ҷi���i@k�0��O�.�7���~^̅$m&���A�4l���q6��t0M��@;�����򃙬�+�\R#����K�Ӕ'!K-�F���?��%�r�镼�M�����#!�4�i��#�y�j���/�����b�tE�����YI�R�X���A�4�S�H`�s*9������@X����P"�76�r���I��ƹB���Vm2F���c����胛+��=3���n�+EP��Z�>V�b�v^��P�=�/�q� �M%"����6.��ir���Xd�����po��p��e��F(]3d� �<BRmRa�g�bZ�X|dIdT!ٷ�Y�JGQ[{����Ęӱ�4�1�(	�P�y=��T�*���S^�k��U��{��"���X��!�u>����!���QŘ��z4>|せ~A@���F0�g�� �&������([�N�u{�}��6����C#�O��ۄ@Z�H�ߍj��T�H_�s�挛����w�J�=��_�_Y�	Q�k��Ðk�P�%{�N�'�b�P#H�ɜ1��D����� �&CȾs"�'�Z�b��8�3�|��-�>̂A�� R=%垿W-g���1;)��c"Z���[����WKY^ľ�M�l����r�4ATGl���(�(��x��C�����ҧʇ.�UEؗ�7,���*��H���f��`��}Λ�RAh+Q�������F'���<�mGWd���H�p�Y��1�_�*L��S	��$L%	�!��+�E���Q�ږO�@xV*#N��இ0d���F�h�~=}��z��:�,V�o��"�7 �8g���ۈ�E;h���ƈ��rݺ_��#�N���(Zj��z=0�l��=�菄�M�h�dX��'EZ>[&�"|u*��$DN��ic��BD$'�C��������;�m�i�a)��Y�h��?�%��@�����W��qig�q̠5yW�t�a�h{�"���Z���/H�C!r��_����]�d�a��AZܔ�B��$N]+>�(NueY�L��t�_����B��H͋ɠ��+{iv "���D�$�E��`�`�7�񠰦 ��@l}���sl�R �ȍ�i�@ߔ�M������{�Q�Lt��Hb���x
�w�Q�!X4����eB�D����w��\dze	�}��ƏR[z�1͓�eo�0�GE��-��Jޤ�`ϥ�ܒ�&#M"�����,@��cK���ɹ�{T���?G�,-?& U=L�r�:�򈤫��SXLgoؠ���%ȡxY���`G��s$C|JZn�������"L\/x�J����ERH�b���m���T,'�����ƐǍ��L^�ĸ��r�F8�(4/D�Y?%�'Z	���6Nq���v]]�pAF��©і��T����!#�9 e���u�%C�yO4�|ό�)h��}�j����n�A ��aXX�ݳ?�l�wm���)�0�2�m��ޗc⾘��|��Y-�1-@��L���>=jt�3���
�.���eX6�B��f�X�f�^��>޴��8#)���w�}NnU:cϦ�d%���o@.U^�9�d@��4��WU�.4�]��y�pе CEiNդ�E;������$�!�>KN�Y�+X�;5Y���ė,�b����%{,Qws�3�|'ܤ�c̶3K몁�WR�|�ݠ��������L��z�����l�ZX�z	�K��|����sx|��'Ҋ��Ң�!�ݶS2��+�f;%\�� �pi��|&�1�{#t�Jy:V���؄�8�k�7��+���ͺ�F䈥��R�P�-d8�`��&��V����d�u�X&e�R�a����ŕ��ȯ_�^(�!�������xo�OE���b��v�Pߓ��И�9�4o�wa�����m`�a�灪�O��&|�F�cYN�<pZ�k����O��k��뾤l�h�.<�/(�`x-b����G���W��|?vJ�hc����6�nc���l0����g����k
�?�
�&�­����� ��u���up�,Ġ#���F���)ˁ�]>1�Ǵ����2�6ڽG<��G�[�>��E�)�cJ���k Y�qj�}@�*�'�U���|��;l/��E"��=[lڦ�H$AQt����k�� ���m�,Qs]��z�]�{�i�)���ig�;��Y��8�\��p�&�=�^]Ɏ�,�z$��Tp�J��$y+m�7ꖖ`�z��㐯�tnx�o��`C��6j�+U��U(d��R��pp��M���o:�Ĝ���@�8��� JMC���Em�O��.�����8"��'\;=�	[ts�P
Ja�X*(Ƅ����j.�O{
�f��A�e�$_Ѐ���y@0�͌
�ѷ/E��6��~k�-�Ow��9'��Py�#�T�ֱf*���4�TUD���X_ü\E�eY�B������kZ����x$]��9��Vd��V����#�/��Ka`={��bn�	�Ӑ����؅Rj��L����{�VB�V,��X�|���g�{ɆV���'���pˤ����ȭ��~/���/&3�53�%ɬ�H���$���{z�%?Z�v3p�[i�A��y{v�/�4�,g�D}�މ������~W�C�sO��#<�3�er�iZnk2��O<"�Y*^\[#ҵ��H�����0G�\��
ꌌb2��֒Ek^�g��0B�(�wEN�B$�L�����*h!�s�
gƢe ��k�U{�O�ܕ�䝥�je��J@�x3q��V� M�	���&�[�n0�'�F�8V7��/i�
6~�\�f�x������^%�Ks�2����ʼHF�jr����N\x�1��B{�[��Mix��Κ�Dc6Y�s��h8������ұ;�Kx���üM�3��jd��X���c'ٸ�s�l;سZ�QM>R��@t!7Fc�o�dM&c]k�ӠM�;���@��܉}�~��b1�+&%dї�ۻ�����yV���.Ox�l<z�+�&^K��UQt�g��	@���X��VB���k3���$�m&�#��yl����M�j�K�� �ײ�l�<�|f��!�^�;=�7-=8հ��khݭǢP���r�^-���FA�I��c��c}���~��4H��8F���C�b�`���A1�h�>���@� �o�x~�D�f��暀kfD���r��f�*K�m~��:6#��Q���t�Х��N��gÞb=v�*}A�+A�x��O�Y�p2^Z����JB4��p�F������������
:�M����	��kL$�J��ǽ����v��R$?)���w�M��ZcZ�ÝzE	�gR�y�x�/p��T�l��i�M0n��1?�SCeq��	bFܕ�_͡ՖCV����&��+#����8D�}�ۏYQ�8Y��j�7ת;�u}��"���y��s;�'vCM��k�l(�%9�U:;*
U�C������X����S�0��6���b較x�['ű:�������X�`&`��������!��#TӰ� ]��������։ ��V����o����;���lE&�_�Ф-�d�=�r`�f8���+��xM��!�p`�����h���8=�F�ƐS��n�S8uy��È���J���]6���dS(:��W7�Fl;Gd�#��bF��f�2�^�����%�;��t��*s �L��w�ݵ�;q�$�Ο�E)�í�/9hv!��b�f�q��.aqhBB���ۗ�M��K[go�l�EF��O��V���h�^�(�C�ö�`j�H1>lW��sh���W'm�=�y�J�F00mS���Y?�ճ _�v��Ń��\�-%���ܚ�#��,�����z�di�ncf�m �k~��Y�ᘖ\^�~�H�Ϋ3e��<����#!
�S��wg�ww��] ^�k��*fDmSm�=�7�/ng:U�t�v^-"��oS�C��M�$	q�����D{���� ^&�����tƻ))�:�-��Y�h�ꀄ-w��b65��7�| 4�]`��G��z��������<�b�e
9��B2곲��: ^z��(�����L�����c�K����
@�%��Xp��ޔ���P�p��6��?��ۡ#"n�a�H���۸DUW�"��KIs
�;�7D����QP����_gDW�!�_α�\ό��k+�����[+��'�o]�*�_���pO���h�)Ɛ������&Hή~՜S(�iqE<,�Y�3�|Z�|�ah�@JC�P��s �x׿TM���?yAA��l4�[ܱ�=�6>�������ؑ6�#q�t,K��(	ڣ���`��#�J\�w�H��O��JB52����Ά���ƚ��x��'�:O�ZƳI�z������ndq/F�7�\e(oⱽ�7ZO���6��{�L� �?�H��	��؟U���� t�E��I{7�18�o.�(	���R�\{��&�'̛1;��W��p*W�� W��f ��&G�x����L5��yzz�+�U����3����f�vf��\Ë�Ǧ!������g��n�E�ל���1�2����j�&A�G�](o�{���0�ww�{p̍TKNT��΀t<s�(��P��c<��5��S�}p/=�����Pc��o=yɾ,������9��̈́�qr��R�v;���k��j�FK�`�v#�!� _�Q�i
�K��vDDDG1π8^qc��[K��x_�*P��:}Kz��M��U#�#u�����z`yvhq�3��ln��Ѩ]9�-���.�Zqj*�/�)����l	Sm���̤���>!���4o�5�+-.�*Gǥ��1��x:����������J��?�6Y�Z^q��)�`���|���
�U� +d�B�QR��|b_۵�ӆ��JՄ�l̺rR�%hɮUQ�n�`����������cϓ���/yrsV!X_L��L=��u �����B��0�z�F�U<��b�{&�
�W��L��"�I	��	u�n>��-����&m�<�h"����wlq����Y�PO-2n���؝t�ER��$h*+ȅNm���-�e�;��7@�a��gm	������j��[\a�vf�F�5U�:%r���f@Z���[v�e�	�%(8Dh��Y6%��.*��\Q�(��U��#uע�h5xbNA���o�6���i���e�h��1�3���&�UwlV�GU��8I��[�� �}J#�[
z~�vx��X�Љ�T`��r�\j�TV���ΑeQ�f%Daf�
i�+1x_�uQ� �+f���ڳ��q����9��w�M�g�v��i�(���!���b8�}\kfNT��]��d)��"�I�
Z[TO*�W�ç�2ls?F��N	������˛�%��4����X�Yh�p�d$K�$�_j)���$�ɳ��XJWCr$�e�������;�7��Ğ��eia�	���H����{s8��t��7��D�T�N�TAY JL�X��^����7H����9k��J�~��;([��=j]k��},�E���h��j["٧��Z߇%���A��2��f�n� ~%"�Xv�W@D�Z*J�Y_��_���(������;��A�0$���w,��6ן��ŹQg�[W�ĥ�bD����Q·�@��,��U���˨�Fv�'X����w6R*[����S�&�X�g��|�{B�Q�S�q��]�E�l5��z[���Wj�0��»ݯ1�������e�0%�F�j��7��?~Qh6\b�v�q@ذ���m"�N�/�,D�Rحʘ�$���ے�yL��L���~�E���.���b��Z����Spu��BZ��	M�@Ȥ~�^H��sG~?�7��-��M�Q�|~��;���'ݸÒ�P?}�d�v��֋�Vӭ��y�\"<j/�OЀJ�E���F���I��g��ͪY�����HGǕ��.�"��B��%t�b�2�������d���K�԰	�>D�L'�ƞB�Y�pW��Nwh�⮬�54�=L�ʤ-.t��l��ΊF��f�����+W��c��$알t���9.9��i���J/��
P��IrE�س��<�� �u?-/q�!�/�A��}(�#�q����Q��>��fnaC�]Q�Q��^LY�16��toI��#^�p��@W��l�P�HM�n��9=(5B���)�8��R�yhׇe̩�tH�DC���:Z�Ѡ�eg�&�JHxǎD��H����1����Y���zs.���R�[0X�#���@ ��e���Dv���B~8�eq�tS�B~�Jl��!�0
[�����,�tLj�w�Ķ��-#����k��(��uc�����\?��Dj�Z/�j��L��0o��E�!OA���2,^~C6ss˚ۉZD4yBi����{��_#5<V�-J�0�FJ�\GV�I����NL��#�2�k��g��[s�2y-Ԩ��}w�[.x\���L*���H�e��{Yϙ_�eڒ2�����ƓS���袎�s��'��!�|/[��/3l��*��4�4�.H�c6WԪ��h03��#�9C������bM�PB����ـ�W�v�� .Ք��n�k��>��eh��Gi��Ў#N@l���ݧO	-L�Fjƫq���a�����a��O1��p�b��A��qyn8R�p	�B�B��^��II��1�����q�ɜ���n-��h������3D�����ZR�2G)oր�����7���)�X��G
�y�����,Y(3g����Xv�U]c�����۴�i���P� �A"k �e{��"�8�y���/�q�����'��R!]��ךz� :��W�\�Q��!�EL~��������J��D$�ׯW����j�@���w�&�Z��[��ϥ�7+�zᆿkfXH8||��`�����2t����V�������Y~qna�{�>�A@�ɘP�x܂KH�V�#T=X�G��>��J?�&�3�"�d�KP&Z�Kh��y�,��x5{=�K�,��`�
�3�p���8�GA8X-������}|'=��d9d{ Ou�(�{��5,}�p�bXo�� �X
���C�&;��DC�>�=�x�p�Lӿ=	���:�}Ȝ@`[� �O�@!�A��c�krP2�gS;,_��A�=��`�qx�Hͳo�VK�3���� �[("��GѴ��u�7n�.�t�}����z��,������9��|w�w�
��좋'�/�JPR��M>S�X�;�F�NQ��`t{�����n: �'m�Oc�;��@�V�!��Klð��iD �·���]�ҸF5#׵\�沢q�;r��7����[���(đ�����.A�Ų|:�����O�r&�n�L�FG˖�s��#dCNiI��&֋��[��p�T���:���/ 8��!0����J� ���h���mh���+9�q����ĉ�P��"�Pɠ�7��2�k�����K��>�sm=�?�"v��|��_Ǔf�(>'��=�:li������S��?ٱ��RJ�{tDd|r��&�B�X�Q�p kV ����j6,Km#{�^�V�\��ż�U�M�Lj��;K%���GS"u�(�"��ߏx�L}�``8��H+���˞#ޛ�!_DзF�Јd����.��+�VZc�V�9aic��?��=(�jP����?��`?�J%u�Y����7����� <��rv"��.;Xe�QiDz�H�����ֈ�:Ԛ~��b}`$=��;�[Z+~筋O��?����Ys�ޜ�.R������U�rkam���^`�7R�����0�ѼӭS����^=k���U.�3�#ʅ%�fN��[m
`��az~�-H{�8N�"�c��Q����ƍ��+�]�h�#�o	�������(z$�U�N8����B��
=�{�X�����^�C;d���Wn4�w�r5F�O=һ���i&�QYꏣ��Z�gq�7��-�?U}��gb�zBFn�3S�I��љ�f�	y]�,8j����Յ_�t@�7��K�Y��ZvM�
*���l�o ��U��[ws�I�y���2���'`�Ȑ,8mm�a)<�'HY��?a���<["�A�"���i�X����sS&�{k���%y�G?�o"�K��$J��B�z_��ܘD@��-��C���tF
��I+������=0���1�^,��������n�����,b��9d�؏R: ����I��?�ls�##��y�ݲ�b��B2�����*������`����~C�
�N���h���2�W$����O�ty���6���aO")M2	�1�'\Ы��c��a�[}��L�����W�Q9�;����\L⣪�2����s���@�Q� O�%am��Lb��������G\vFpj+{�������m��4%;��V��!���e�~�`���h6fkX�N6��������f�$m�v�UXe��Q�&Ě[�(��R�k9Y��)S@a�b�XJ�A.��T7�:�̩�
�=�\;��Kr��|�u�@HÅ��d��&k���Ϣ�U+�&�?,4�8a2dT�EY/W���jHg-���!��;������A�� /7�Z"zMr\�"a�k2�� Èd�m�c�P��	Ċ��.��;�4�0�;�-�dY�(gY�$�8v��tY;��$),��'6n�A�\`�5�0�na`�7F�^q�⏩��Ꮪ[�r��.mTdM��I^�]������Kj�t��*�,[���2q��\=����v~�z��g���uAy�An�"]���߾Y?��Q�Iބk��}�Eќ�m�����S�ϔZ?�Tr���(��Ր#ɺ�@��y�}�֩<�X~Z@-�x�+�.�5�β"k3�� �.-����T����w(k��h��o+�!�M�whj�5cg�����TF���l�aqo3�������*XƯ|GU@,�gŸ�%���5�J����Z��j� �8��žLJ��_���V2/�/E����iN�#7�� ��A׿Ռl��y�.��:{�-�D�E�����G��q�DYqD�������|Yi��PO˂��Tnz��?�$�xF��~6�g��g9-�J����Fn硨ǡ��p%���>��;����Y��a�����ʯ2��v�D`$>�F3���o�Lע���K�#�$���X��#��(rQF�z��5��,����n��_݄�g������L�m.��t��$-0̼h�U#*\����mR%�f�M5�oq��,h*{G��n�C����9;z��|��O�Dc:0�����-H��2{���*����TG�BFr������s Ա	��6�W�T3�V���)A{]�j7������|�{̭)�)���Ge/]�{J��&����٥`4A#�m	�z����P��Θ����9��������+�Lka���W��u�<Q��k=ݼ�(��>Rc܃�k�s\UYNbλ�Q&,�R�w�ю��g�~	�N;-|3:xY1��o�Kڷ���*��y�"�ӾR��()��-=��:t�&��k�k&,�w���9����ك�~ǳR	�(qcJ��VE�ѯb����+5�AR>v�w��rk�s3jl���,(\s����{4*�z4�l��w�����MQA8l3�� �<�]��	N��9$T�L0��C�/ ��+�Ѩ�΀�4#��H"7QT3i����}�����z��7�����W{~�+�![��N��F�>�;\��3� ��8�������3y�d�F�6;`"�Ǡ<1��e=�4���j&,�* {&xő��%��V�i��fX^�;�QPU�lh����k��(�����S$z�d� �M�5��-;���[@��J�n��U�N�%ϡp~�H��\Z�=��\}E�+�T�`��Z��XW���}�LN�j������7�T?��{�ʫ�������;��F� �����Ba��)Z杴��|���#\�5�|s�Ұ[�8jk>��s��e4(�Y8��a� ݸCؓht�:s,�[N��o��4aAĵ$$(}�������F7���l{�Bٺd�H�Q�a���R~5����|>}�G:"����*2/�,hCz��K�?�A�]e���-7��%�k��sNDk(����򚬀Q�uN�f����VmT0MN?T÷ff��(�&����3��8�@N�C�L����8:Sb���@����|�[<ڑ=G��O���z�7U�~�����v;�Ű��M���ôw�0d��O15�ƌar-���VR���@��Y�ۚ٪ؐ�v�7�j�+�w^�2P����n`�Ϗ�i`� ̀./1��P���Y��H�l����1U�5(��O��^���Z&?��Bv���x+��(C��[�x[�)H�3>�.9��k�,�G\?�]B����X��*$�,�f�z�vH<��ᫍߟ?��P��X><ϣڸ_|����
k�U��N�+�X���Ė���  9D�S��6��X-kE���!xc]S��]�S��:Ē�M�ns����^�nT���1�,'g���o�'*+��H%A��
Bl�);|�(�y��"���'hӡ)7�ro�-b�5��S��KĔ���k	��̸�DW��Du{�i>�4ʣv��;Mgj� ��^�X��ẩp��cN@�$�z_Wh�F��n�8�cs8���|6�C��Q$�Q��5���C�h��B�S�z>�ri��V�S��b���ƥ��`��B;�-�Ԥ��c�h˵
��Id{�(z\m�F����^>_��WF�i���·���T�yRu�m�;������������~�@�}��fj9nZ3��Ge��$Eu�w��õYd@��N�@�y�����a�۱&�J�*�7 �O��#�Tp����6�+)ݜ����\"KuR+b���3g8zZ\�"���.�"����XQf�W����O�Q�.	U�Ʃ'�JMC�#��!Ш�p�5��!�wg��t�6�����Ph�+�/��X���C�� �S�<�Bj�:�ȱ�(��X�� w�����z�U��<��M�(�Q�#��q�Y��oj�^6�ӊ<�Ƌ����%V����aQR,VNa��g�-�
�	�?�4ӊT@��H`�H�j3@�{��|���Kʇ�Ѧ�u�#�=L&�mN�ő�l����p��Ii�w	U�"O����4F1WY�@��KAQsw&��!���}�礓p�L) c�#��<�1aJg�Oř}C+J�0�D,q�����KK���4��>m��~�����_�M"msZ*HY�V��A��h�21&����Ґ�R_	UQS:Z�	Lϖ�eXus�|۵�\ç��6��z�J~D��B�������R�0F8�#uL<��'r�ˏ#��ZϢ$����� b����	��L��]��J��5�7�(���<`���S��H�R�#�{!��x~���<Pmz���j���F��� B^p˂E3|宝��m��C�*z��<>�������ϻ���F�f�0S��m-Ffha�b�5���h�?��m���N�~���m��veU�	�:\U:���T<%�0Y�%�bk�C�/NM��5�؝��H;=�+�Y_�4�K�b�VQs�^���J5;DX�E���Z��J&� ��eQE;C�
�5��I�2�����l�0��u�8T��F���G��[��g�y�\�B�l� �q��<:�qtp�CZ�}rcx��R���ZGI�L���F��%�)�!��I�~W���H��n�X�����^�z�ͮ~��<�B�I�X��X1U	�[��r!vם�6���&v%�g����!�k2�y��%�"5���TU��>��I$�GM�=�^+O>�o?���F=cA�Il�����:K�0b�~����;F��᜿+���^��e~�lܜ��9��T酤<o�!^;��C���¹M֏P;�:��F&S_�l�x�rwe��<����������`!L��DL�B�!Zʟ��р��*w�璐H�Z�ŵ+�W�tϠ�D��$~�}���](�0j�w~��S��� ��Ή|��k3�a�~B�|Ph�P4D<�m�(��Z�Z�Z����]����o��T=�=��~h��ve	<�Q:J�9�@K->:?�F���O�5��*�6�1�,�0*���A����9��_�:���|��O�n��)�L��\��7Zf��Sa`8.1v!/�=	Z�(��C}r�'XNw<� �-�
;��a U)v���l��_���چ]�M��mi��^���^a��-H���lj �Q�+1_�
_A�TLI��r�r�����A����E�6�+U��֬��InAx��Ψ�݉���e�/�+P�A��<ɻd��!��S�nr��v�V}��3e����?9��+1'�[ր^jD����"pbGrW��#Y6̀��g��l���hO�]@XM�?�t�_2h�ږP	������x�Cun"*�@R%=�A����20�VӭnEW�O�`������iv~"(LxJ�}�p(G�>|����5��+e^�]�����A3�ڹ��y/k2'�w1�D�p���a۹m&�s7�&��WxjC;��0�ju�S^>u�|�2+Zw�&U<m.Up-����l��t��rY�r�Q�?=D�����{E.
�f��B��#<�h[)��H�Cgp?YM���i��]�'�m�A.�<��V��0��K6=��� �ZX)��GR���On��DbB���iT�(��o�Rڒ%�'�_���'�"��[�M\��#)�y����DW��c]0�1¾���k��N�9�h�R�^�m�CR[�[��ȉ�����)�<=f�i�N�c^���ֵe#�}���2�s�xq���q�Uΰ���ˈ��c ����CUb�}��f�k�"��7��_sx}�����G��f�\�� úe�M�_�i?�Ex�a\�`6��%�1��h��n�'[_����,%{��v���܆�1�>���B࿫۬�gUR�;�,ƶ�r�O����N�{|}Ѡ_GV|b��K'=�F]�R���Z�Ž1�7Ϊy�Ԛ�*@�]����<��G6yШ?Ǜ�a�4�2I�wa"q�{�7,���x��������n�����d���d�qL�Kg����IY����[�	 �Uu8�7����=�
Z9Y���"�ќ�A^��k�����9��QϜ��0[ۿ���Z��A�PS�c��MO����d^�`3괠wu��܃n�,��[l�X��t��άM�����;��kl���~�0���H@+� �r����_I韣��,p[��Tg����0���q��dSS��I�����B%�{�r#���m+΢s_U;_ Җ\�ֲ? sl�NN�i�����$�$B Pr�E��88�u2ۙ�)��-׽ ����h��0NK�zDQz[rrV<�<
�N%����/�&��8Ĺ�#�x�切{�W��
É>�*-H���PA\6lJ=�~��B��8v(�vPK+ߘ{�Ͻ���ln"[g|jj��e��*����g���gf�̜�+%�f��e��L˰4�J',]��L�\Gv(���w,�-[������g���?N�9��(�#�W��0�/~r�ě��I��"�.|\����s�=b,Zs�ٵ��rz�0�kۓF|�Wtɖ��q0C8�F?J������NG`$�a�B�/�Wj�1HE���	�I�s4�9���ń=h���:�A�Z�:�im� �Y66!�c:�k�O+^��`�q\�)5�j���X�%3?7��02t��"�L�s����%�|w�90�S�U�;$M�X<@.��!iԈ�ߕ�����o��f���Ы��7x<�E��a�o��B�O�N��X�b��1��;ԃ��"��Cw�Ir��J$����]$з��u�碱�N^�Yu"R�	5f-ഷ�D�w�S%[�����*�E��V,���.u臰��)���Ӱ�}�o%�;Q���'&e.��6�Ո�Q�)f;�t��>jB'�1�]f5�ǌW��[�\�,j�)Nz#K�}���C�f`|�A�2�mD�iǿ�Q��x<�m��d�𣴥e4`��J�w(ľ�8`�\>� �Ƀӥ�yk~{;�����S*0��MӟR@�r�ȯ��.��t��5�6֞^�����
C�o�s9h����j�x�z��� !�]y9��f{��a�?��_�~)�p��,JJx�0�_ӄZ�����p̈��K��k\c�(��8z�.oE�!�O�����鄇�g�TX�Q�J�����(a�1�+�|bj���Z�:ީ��-��cCħ�����_7���$��$��r�(�,�)&�Ѡtn��:�N�NȵH��G�N�	!�c��aA��>�6������).7�}e�sɟ�K��֏�/�GIy�q�D��g�2��ғ���ؐ8��J��*�Igl��:�y٬�>�'y�k��X>����뇿Бuf&f��I�Ä*����d��*�")l�tJT&)�3i���%�:̥<� +J�B-6����#߻o��j!f��{JSH�=���B�����y@������w|)��j,�a����dx�A��:�p��;��{
���U�Phn�=^�k
b��:��뫺���[�?����;`F_�� ���RC� q����=�����N-�:��3[�V�.v����i=��)|
�e�!��Bs��B*F�1�_� W'�BW[�'<������,��?�ag�|���c��W����2c������Oyʹ<}%�F��;nU�.�t�%���}�#u���I�M�^܌���#E�׾8Uڐ�'���h�XFB^Mh���i�HN!��a��I�r���CPCHSv$"ꆊQ�6�^b�6�&��>�{�P.B�&%���8��5u4�&pÆ=&�1r><����\~>ܗc-�?_>5��۹M�#�}E��M�����S���M���)�-{1	z���0�T���-�)r�7gprYG1����mA*>��f���
�pX��s`��|;���|��>Y�[٨p��y�ތSg3"E�N���4�F	��|(ڀ<��i�	S*�y�#�7Y�5`Enfqy�7� \b�gT�i�e��4bM=gM���Ma���1xF�g �M�$���嗪䮽��6�r7���J�SM��ꍦ�hOC��n���DzNC���h��:�0�f���]7d�� 8i2������Ū�0o�߯%�1�!�r�s���c���Y�#���<fb5�f3���_`d(�M<�宖0�_[�-NQ���G2���S������|fk�2I.Q.M~
�!I5	��0��ӖL
�����^h�����&U��U��ɸv֖�`B��FGD�?t>]��A�O�!ým�aOc�>�R�S���p��_���+D�)Ӱu�)I�˖�Oea޶Q@�5�y����v�
���&���u��q@��D}0���6f�k�:�^��9�$��h4"A��͗*#B������M� O4��&�c�O��򪂙0�B���;y�Pbj,0}�?�zא�+PǷ��Ż�o�@��%��24s���Xu�K|��3C�v��I$D(�7�n|Y4$�>�'��-dO�2X'�S�."��J�� 9o���OQTYO@�����:��.6�i�܀��'2�n��=�51o9u���Y�����͉	�8ӟ�w��s���85q��AwZ�;�_� z̅Vp%�0�.i-$��� D�t�l"d�wnf~��]��4p6�\/�g��w�
	L��v���^Nx��m^�Y���W[�<��kR=�ɛC K
��r1B�+f-=Bw�9WT�(�4����(�oo�	Z��>�Y��`�r����p����1�2!���b�0u'�4811؞e{��d/��g�-�7�HżgrɍV#�O���"���y໽�E��/o:b
�2X&������(U_e
5��ᆑ�g�ɴQ�\�l>�.o՞�L�Y����2��X#����K��Z�*��Ha-�g!5{���0Mf����+���c���
[�-�G�{zQ���'G����$��Ga�K�Q��N�V���n��"���^�f\	wf�m���q  ��ڟg�Gն&�_e��QC�i�N�[��>!�{�Ӄa��or�dH��@� >:p�*;�m;c���]�xm�r#���V�[Cmן��$��0?Q�����vc��zV-�.liS˻#�@Qy�54�Zj���@��xo��y�ɸ�]�R)1�
�����br�tY�C%q��coJ`�������1(����� *fZޗP��{�h���c��PY�Ϋ�㲶�������'ܞL�ð���-[,坟�?b����
���+/^&���=-�Y���!����iӢ�Bʛ���)��p9s�Ns�XA�mdR�X1��~�}�HE�Ur�{���g@�yT�Qa�Y�1��!p<�ǭ� ���S/>�Z��c�S��s�e�I\a��W��6F�S�����E�9Q�5������j�	$s�� �l�_��z�6���(���w>� �d�S_p�'����#�3i) U�'� e�N6��2��Q) r����R'����'Y�_������j��.��D�5�K������mb��yW/�O/�N�g�?Iq�>`�"��z�����:��sI,��o3v��`��TM;f�ㅛ2�(E^�pQ hmW�J}��L�Ǵe���oߴ����+l�2�������s���Gh�4��r:v��P	't�0k!Q`@�ؐZ���5���zk��w���yvɿ�M�_|�����p��95��~�:h��N˘Ϯ�-�7�ϟΐ���`WIȤB�2�K��S:i�~,s�Y����Lg���rlԄ�y.��g�+Xئi*��1�҂������pߙ0�9� e^ׇ�%
V��s��)��������ơ~�U�	���v���b6�S��ŉ����e��i�Vq��i��Sb	z�*���� �ķ�|B&���Dyd���p5��ӏWw�M�A�Wsm�A��m�A��MPCT,�պt���C����Z�������c˰��L��8���A�᭘�#D�dI|N�̥{�� N�#��"�-	�B��麰Z.XkB35��4�I���=�լM�B^��c���_lR�[ɲh�� 6[���J�:��W+�_�ݡ^��8���-����ZR�Pp�Cf����^��Q��N�C�Q�����sa���s9���։hG�͉�RDr��І~S�_�Vuۨ�It���NnM��؃�"���b֡w귞ӻ���M�st�ՙ
��i��1�#'@ͷ������17�k��\�'}�-6q�j��C'�������n�+��C#�@�ށ�.�>T���) �c�P������	E�zP�;��؁l#�������$�.L�<T9�ɼ����[�ݹ�yˏ~�I.Rz�=���j��4!����K���ʯ�[���kR�R�>R��.}A����c�ܺ@�����4��J`���lb4�MVK8�63Z�qv���)^}"Ż��"4hG��!�+$ "�U��|J����9��M���[.�@��&1�ߓ�/���DH����h���Ip����zA���v\R��a�������@o�Ӷ���X֍�CUGMJ�o�{N�^Q_:Y��}�J�P
r)��G��:T���׬��WF+I���xb���}y�Zf�(+( K�k�|�[���ߝ ������f+@��7��e'}\ط3k��z�e�r�`fY�mʫ|�G�R-�GhR�Z����<��J�T����?�ȴ. ��3�r'_�����
Mp<z�0Շ�y��y���7Y��$�5����K럪`�Y� �MtFj�ho.��D�����lm�Bcd�$�����|�ɪڡ� ������{��;p'��������)����!.߮l,B�5�����<*4M�[L���4<}ȇ����@U�kPn���yRI�r�'4wu-��"�g���ɆZ�GU>�xа�(��%:v!��5&2OйD���8����4�$(�h�B<2��;z񶉌��a�xA��NfJ�21�>���~%��B;��^������NL�]'��*{ϕ$��#ͨ4�j@Nh�/}�R��ۻ�C	y��������N���9��n� Gվq;�t�a���U���p�6��T�W�n<�H�f�Z���y�Ga����A�g�w��B�P�p��qT%c�EJg�E'=8�� �\��罂V{���6��rѿiE����$�z����̧cV��Ԡ�<�^�<*|�(]��8�,�1�[�`q�J%'�;�ץ��k"W�k�P;���b�F_�z�Im3��N$aD�v�u8�k�jy��:�4 Y|K|�=��
x�競�G��<�	�p���I��YSJ�|J瑬V��#~�	Ļ(-�}nĩffL3C�l����b�u���A�C{zK�7��:@�����_6��3�*�xN�/�.��+�7�~�f�����BaY���뜍���H��)[��Ky]�n�6��,B8(�4d��D�wm�������onJ�Q�6� �����k ���t	�*�hFQ����	���pUn�Å�����G�^58k&��(u���<�����2i��CS�3^�j�h<��̎��ˢ��碡i�w���^ٟ���!W�G�5��}9�N2Z���6Q���.�z13�1lV����	�Ͽ]@��߽�U��l��@��eՙ��$��� Z��r��Om����05}�͏=Fq��9md����A�������c��f�����X{K�4\)YD�,�T�E��w���ߞ��*�-p�K��I��ו��A�z@��\B�_�Pj���8��*6�e�E�6�g�}M���U�l��6#2�cEH���x�y�w<8~ISu�o��MK���z�c�����IO����)�Ax�S�VU���+62s�>in�.��*��'!�2�c�M����Z�0�ƥТ%x��>ْ��O�Sa��ٙ)��r��9E��'���m)�NdǾ�~�Ork���(��XV䰠H����� 3�.��[LYG�^S�*&z��w7��E�֭~cQ�����E�,��Þ��2���܁]�; �=EXQ��"&Xp,脇\ar�;�]�rF���F�KjX`�=ļ�أcd:���B$jN���B	�l�<���g(���"!�#�{�t��Զ�>��\(M�)��ME�3[��Xs>H<a@?�+��Q��#����s�hC%C�4Y.�ao� �a�B;�+�uK��1�#��aeS�~��b�����l���	���-u
{{װڢ�����((`�Z�O����[���PT���uG��;e��_�K�McVb*ڞ(�9f΄�)�'S2*�c-��R}c��h�=\���h��b�L�Vі�r]B{�zs����ԉUW���=�F&�@��\���=��6�ThQ^'
�z�����`��)�iL�3�k疗A��ѰP=;w��fa�|ψ�Fzs�}�l���5�T���������u;F\�U8�o�ؚ���Sm�iT��<�-"P%O������5�����J��+Q��~�i��:���_~����"�|g޲�@��c��n"�NZ�X�I��R�@q骟^n~=2?�B��-�~�f��7�~V%[���#>�1޺�BV��e��Ғ��6��{�#�OS��g8{��Ƞ�;�����'��D&�S5���Hv�+�4�(C��	���.^ǧj�VE֏�:Y���}�hV"�(�Y-dmxF�e8�}Q��+$��,z)3d����f��~w�V���hb�Hz�!��g��t()ު���[@�Ep � Kx�FL�ȧ�|�˵�.�b3������F���X�Y�n�H���	��u0L^����KٮI�>��'=�R�X�Q�XV43��A��~D&>��}E �}��Z�vA�vE�F����.��+d��nJk<���[���b�ͤ���E�?L��1q���p��ۙ��X̸�݈GP� �Y	I��p����}< K���O�.W_u���%�Z#����,�xd9��W�aJ�-�f�lP@,Y�+�t*��U�3 <X{@�g��@U{<�0�F�˵�V��X�>	sqd"������_	�5'餐 i�^�a<��&�����o��Q�+��A���ä��o��n�N�e�Ŵ"�&�Z��o��Il����]s��[D�ߐ�k�Ŗ�쁳_ev�#�U��a���S��o/F�j�5���8���0�33�м�AM�*t��V�]0K�"�H�Đ�[�{>>9�Ux���u�3w�$�6ǩ��ۛD���\���wj"�S[��zX���oL�d���-F�J(3>�\k������_Sj�Fc��,gY\
W�X_��pj�s�W�<U!v��h]���R��0-�/�����c�� d�B�}���o�&ǘ�ͪ�O�SO�V��<E͇P�\��{9���wWΑ��4dj�x.�_>�Q���4}~�/���)��B���uv�?�5�fr�+�[!|=���I<�~ǆ�L��̉lc"䰃�5� �)>�^*R)���c�Nb����3����6Q�G}.�L��f��܄�C��� �J���]-��s�u�$���ݣ;����6V[]m#Q�)�?�N��I�+$�].�]�;l�,�C���H��;:ǟu���}-�_���픒��+,�����K)6}E�P�_.eGeP��q}A�X��P� 鴹3����R��?����
]`&���(e��'��Iގ��e>�>t}T�H�o���*���t�Q�M��=VZ��
�;viX��xW	��h�jV���~�.�aW�M;�J�lg��
�?�tT�G�����ҏ)ü�P$m��Q�8��E�����!IG��+��UԐ!CE�kd��!GM��7&���G�)u`�=/NƎD|u6����8�����͕�&�b�����!.��5#<��U�rz��ko�k�JV��?-�8"�!��Fj��WH=i7 `�.����DB9Q��������¾e �{�$?�����Go[AWs�_A�ly��Q�']���y̾%��p�� ��%x�c��ꡝ.�#���EP�-Y }���Y�At���~Q�*-�����x�F7���$,a�Ǧ���0�\j��Ms%�z�CX)U�|�z0^��	Ut�i�Ĕ�}4I�R�g�w��iY�|t�\�4-�)|ޑ��Y�����c�HtHM\�����Hd�#_N�uݗ���|�V��	�"�
E�f��DzI-#�`��ow�-��8��/S����P�n諧>9�C%<)'�:`� 9A�nA%o��O�\lo�0A��kU`�٪���� ��n�	;.K_�<l��B�տC����C�C�e��Ϝh��d�o� ��]���J�&"؛ӂ�+"�C�JB���f�P��P��Z���a���$���}��\������jQ ���z��4�4'����{u�订ns(7��'���휳]oֱN��f������k9	�`��f0%��25������&�ѭ�3)��U���f�G���$���@Jt�ɗx�Xi���6�ÖC�{L���UM嚿����~��7���y�>:s�v����	~9��H��Ǧ���H �e�"�ި�'��7��ՠGT�̀�-Q�#�s.��L}����8�����C��aR:���F��~)��7;��q����l	 �&M�D�NJj}�kB�'�G�]?�
a1��j7�
30X ��\q�5Y�CAOm�$��4�
���׹f���$o���4,[<��w�(�U�:?�R�v{0.@_|�t{�����5��Fg��~�������]R��br%��ܖ���3��%����Hn��%��\�=`�Y����fnҕ��@�Ig�,~��P�]��)
}�Ii,S��ښ������ �kT)��� ?�Z���b��L�mH���1�n�t��ba� ���_�7��P4����,��mʑ��62��� o����m�q�����`6��#H]�l껱E�ƙ˶p��X ����!y�I`OVP��^���tY����nNJS$�Kn��6�H���f怃E%��pֹ��ň,7��J#��p"�^P(�=��ޮ��uC�����t��m�d&k=M�@4�f��j�%�(Ey�r�|5�K(]�Ph������+�'	�܊6��佶�����D�7E�~�#�����x�_�m~�
T`�*-D���1�d�s2Y��+��{�B�u�LH�����i�c]�|�m�ѭn���	�c;��ğ��!Pu���f��g�궒?�O.J8����]0vJ׸�x��C�x�%�`a4!�������Ȼ��>\�~?�wv�S�$j,;� P��(��i2x��8ޡ��v��U����l�kEʱo�3�g%Ih�xj�s0�q]���a���02�G�%Rq<�#s*���	t�F�x�Dlg4e51^Q�p�p�\"�8�c���p�ʪ����e��`ʋ� ��e��o����翣2���5I?��K�0'
M�d��%Pe!0*���%ϔKw�žyW=�bF�p�3sB�Mx�i��/��<#:��U~�p_�*P&վ��{�/�E^_�Vg2ݲf����� G��c�g�y�!c��b/��y�]�Z�D��6<tO�GC�M|i�QT�� �Q^W���k���T��+���_�š
�Q`�!x�=���T)�:F��H��$���XZm��'�G]ݖ3Jl��9k���x�(�:k3�N|��W"A��"��.����z�[оVGb�	S��O�oFF�A��]��0���v�2 �'_Yv_1g��Koչ31�^.�U7�� �8���%�b5A�a1�F�b�B
��s���,q,^�x~�.xQ�sX�k�$8o2���P:������X�_�JƆ��Sv1�Gƕ�ls�Ȇ��v�q~>F|��h- ��. �?Ed��4^-�"�B���i*���ޥ|Y'M1����0�K���.%�S8-$�b�\=�!W���?���Gb��iW����Q��k[�_��!�P�qJ:�{2��N���*v��a�|�>��>l���wz����1���@�=4
&�&���QQ���m��cOM��D��[�Xu�j��ܹn𗞁��Xn�F�.�N0���V��k#ӇR�X�-�-�
���3���y��c+ ��,�\e�!��!O1I!P ~=����Ō��\��zNqKX|g��H�5xG����ߙ���tRА�K&-�?i�5]|�#�e��+1 {��I)A��z� &!Xg~��[m,���U���Y�+���^�{��"İ�符����u����{�����t�|�� ��)t7g#�>��Uȶ݆� 
����J���jh��y�=��@aĻ-8��0"���ؿ���BLM�!��<�`H�Tp��vM��VJ᜞kuhK�i�8��4T��
��UL�3�|Q�y!n��=szγ��+�����?�P���7!.s9��({��"��z�m�ԯm��굔�j�G\����c���ɷ|5�� �Ӕc�_������,-���j��<�ˈ���Y�ֿ�OjcȺX��}��p�!G��Ző�uu��a�hذ�>�s��=�J�gvU�#�S;���:�gj�,�6=?��~�W�M���R�+�2����**aA�������ٵ|�kZ�D��hXhf�u��b1׽�P7����o"9����ʞ��m~�����'s������s��wD�a��[�^�)�õS�|7Q�d������j��/��^�bWϵ^�H�}D��	���m٨���r����X�'��<���i��L�ղ�>4���=s/��I�0����C-�9�W֢���ß6h�V-ѠR��#e�@$����q��N��-^�v�ʹ���P�sY�x�yu�Z5l���Ś'��L�Ked��o���TX����[�+�Ϧ�h:�0�_�΂�a3dt�E7Y�CFl��!%�	4>3�F�drd�N�A����f7�	�ɾ6�g�b�|�>2�^�,y��Q3�"�8���B��]���<���#@no�p��5Af�x������PlQHF�x���>��/9��1���bn��"w(��#X.ԃF�Ds7u-F�ZRܑP������yEҔjw�W@���e��0n��{]q=W�0�\�zK�Ϟ����3��q(y�s�~�8���zw;�)�4�8�w����o�r�,��Q��*o�B��-Ju�-�o��Pgj׶�Me&�!������$k�w��'C/�=ڊ8,�:��`����������e���������~K}#�J�� �'�ǘ�/N��tXG��|����.!5X�c�)idR#�~�Y������C?[��5����T
�E
�j�vŨ�2��)1W办}�Y��!���M�ݶ�_�I��d�	��͈!�mʦ�E\�h6=Z�-�����Z���`d!�Π�;VEd�~8���nZe��
��t7�"9��2�o#��+��Zu<��Dy�Kc�������7��/=�|<L�_�~*U��w`#��  r`TQ������	E��"}x{�C�d��lM��>i|8���'��p�9t*���ISj_�â� ]~4 ��~�H5b���]�����<Y���j{XRu_���N]`<{4���W�u���~�
���@W�E�_0n�by���G@�Ά�mS���L��m_1vME��o�Y�G���|�l(*���8�����!�R��ҽ?71�շ�oZ�L?,|4��K�	�i�8���Z��csxș�����1����L�)�� �TX>���I�V���������H������?/��4l'Q��"�f1�����@����B�w���Ŝ��)�B���!&�\�1�B�G�����0�
s`��
aI����BV2�ӥ(��to��@̯C�y~��'��3�����`�F��Rau\X!h�&	8g�o/�c�<+��"��zZ�<�:�G�Wr���%�W%�nb�UO=>�����h��B�@o>�/�c��ϨfΗ��ڿ�޵�,��������2=�Q��ck1�f)��:8��a�\��8���1�`��$P�<��b3��f�0_�+��9U0��kT6!M��aU����7���^z5�48���UH�=菼�k��ǭ*��y�#��(��?Ó���WH�U�O�+ʎ�0�q�-�����˺��S4`��T�ѻ�3rd4�Bq��㗭�~��ABiR���ۄ��H��Pދ�/�Ĝ�)��"���dWP����5e����8���S�Q%��	7u7�p�96�Ƀ��yo�ED��dZi3G��gF�Ҍ����),�]��x%�įaBv���)�5��/->�u02f���CB+0(nO��pj�'D+F�G:i��š����>��"��ғe5�*��1^�f@�w9ICʔ	;�9��s�SJ@$Eg�,^p��G*������,��ͯ����J&��*��aw�[M�#���|��������N⯔�hgm���'F�E�1�2ѷn��gF��e��m����H>-���{D1�`��J��^]�I�V�pg�^{B$5 ��~(�>��
��h*���q)l�5�W���_�
k���ʝ�ڶ��}0@��j<b��Ѓ�<*��<$���%¾���	�_���&<�F��z����e==Pkt�����{[2�1$������g���>�8�w�Ofy�"o�Rl�6��:H��r���8ۣ�i�G������!���^��[����}�ء[�ΔK��M?-�j��}��Y��u�$l�ek�����=P|�Ye��yo�;����R=~��g[��`�e�t������]����`1s�l�^q���3?�Y&��i*z>�W�|��a%Д���j��oN��?�����P#�I�T� ��޺�sgy��Ÿ�罂�0��߇$�.&���/�_PQ���q�I�Z�@�&���Aƅλ>��Y� ^/8�0q\�[���Q��u����ڰv��'�3浧��Vp?�/౴�ZЊ�.��H3��^Μa���GGb>� hKkt��ZU�ÍϔV��ͻ*��"�a	��)H+#�ڡ����+�zC��',�CzF���Y��9+bR4m2d���p�>����7%g��j�7 Qy�Ma|�F�'���R��G�7a��Rx܄t�Ft�bWF�7F�"���/���M,��\oY���u�A������H��W׵�L���O�'����8dH�C��.���nؗ;��u]1w�M�T��Od�~�.�!�� ��\�<bF�������X�pؤI���m�h 5�Fp|1��)p�x�
:|�v�S�hmS������͓ f��H�w���?�9h�t�E�x}�sۿ�eŬ�q�"��26����t��?�5��~�� �!�]�!l�(@�B��"�1�D��n�҈���X�l��QJ+n'�H$u������`T�?[�����r��� �,v�'������G<k��ա��N��l4ORdM�bj 1��|۲� ;u�/*�I����@��3�������\k���x���O+��w���A�o\����N�����_X�f�35Dհ���2�T��I��%"&���a���RiK�r�m��3�'���#"���RC��LҔU����+60_�ay��ν8�i��Iu�߃�b��3���u��#�zj~(̯��Tw�)�;=3��D�H?V&<���+[��a{�p`2�������a�`2�Tb�Hp�}cV1ݴ�"��F�!�n(Ɵ���un�,+��P�K��_73��3�3����z��iV���~�F �2Â�d.	�{�	���&�⑂:��H�3���2�^�"Y7�?��Yc����9�T��r8�Ź����m�3�AyBU�@i�!�����۠<(jvlAZ�O�� 3�3���)-u�����(�E�����O�v[Om���#�V�]8c:(�[�qC4=�&��g�Tԟi�����E���4�M<�!�;	9��x {b� �� O��_�ˁf8��nP�6_�rH���"�o��Pc[#B�*�����:�>�	��l\r�<���=�D+���ӟ��!���s�B?_~���<+�,�����2Ƶ�1��b_�x0��iu1���ױ&���#K�Si_���6�V�6�=ʷn-����6UE.;sl0w��K-�O�WI���s2�t�r��Q+�0�����1y��'���nODCXy�'t�&�.~xhCd�&d��4	iD����J�4�O�S��3i_�V��NR鶩���l,9L0�c�|�b���YC=7�u�3F��1oG����f&l�K#IW��c�ֽ�3�8�dZ����%��z�<�E*p0���Q�6V������ɿ=���q� ��4�s��ϗ��Z(!��`Md0���{�~���,��4���bC��90�m�����:�zc��{��z0^$>ꢀ_�Ю9�� ���Ӣ�5W&���(��R�z'`lL�U��<����Stt��%y�d`��p�00�'	����iF�EH�7w�T*i��{G���j�w��	��9-�]�K=�]F��66�I/�w2���B͍����@�)����ؾ��B�^v%���Ǟ���0���xT�qx7`��a�`��䊖���;�.��E�#��>s����g��[$��{J��";���%���Y�8!�1�'xEz�h�|m��9d3�O/[�-��	�dA�U��]I)%�"�FR�Rٯ7�:o�����Ð=��\̉�XKO$\/*�{�S��}����v#��X�2�W�J��8iD��R�����LO�1�ǉ6���
Mֲv���8D���9�Z�*n�{�%Yo�mBY���#��Ac'���7`�%�^�}8c�!�j�_���#c�ˁJO V'a0܆)2"�+���ڎf�M���Y��0�6/��N}-<�(�X1k���Ih_�}����)o��~�A��-��:2"6�r��o<[Z#�ҙ@|d���J��ʆ�Β�V;D�Wu��u�꣡���ǻ�c�+@!�)��n�x��R�Q�����M�(d�M����B
���ڼCd��;I�U�N���7U�CǊ��b�����6@�a�31_!��Lq�����j�Ep��N*��
�%�ƇЈ���ԭ����Sڦ��c_X��S	� WBO
������.��=&5�a���0�b* �p��/)S���#��*w˦�7�������?�ϊ���+��e�M�~��<�vll����H��^��c�1a�$4����I�&�7L��{4�s�F�oE�d\b���W�Ӹ"�����p��42�*�4
�]���S��~�n���b>v��?%�8d�|Y����Wg]:0KrE��g��ځ�\,�Ï-���b�;k�ka9҂����F����ʈvh�l��rO!�S��2����ur�#_n��tn��Nk���?b��0A�����#���r�u��s����.����3��z�>��R��٪�߰��	#k��D�֜"������������ҡ�xh�4�,�4���0�$?�S� ���%=P�4�QSj`��B���վ�� ��Pe�`�����e����w-�E	�(��i�
 �>K"�򀌫����RO��2ʢ�ި_+���gP|��!���4ȼ��;d�cH�{$;N�V_]Qw�e�e�m.���u��v���K�b���)K5���P`�Ü	��2j���jy'�3�WW'HO���%[#U;r�R�>���Uݞք�_�l���$��m� 뙹�4�n�x)g���F���:�Pe�}o:�?��z�X'�U7�OŅ/�D'*�,����t�{��^&���޸Un=p��vZ��0�$�Fsn����on�fjْ�~�;Z�G�lT;ף������롂J_�$	��`���v���-��;5��/����<�ȠV<j�4�e��0�|�?��BoW�)��I���i�D���{�4)<m��VyQp���o[��ƹ��+b�1*v��T���0N[攆��==��q~�	V�rm7��]*��H��t�x���{�S܎L���};[^��Yyr��J��"�E::�O�����T_G?�8-X��6�;C�����#��Zdcó7b~��C}��y}2���Y
M`�ptH�r���ϫ1;��w��\nO�f��p2�M\���w�j�b�aW(���65�^�`�J�>���āYw/dR�(l�Y��zl��o�FY�	��"����BA�Q��5c7H^�����d�@dl۫�*'3�lU����_��{��w�扆��󤳑�mY�+Q���$��
 B�}VʷW�1�}Zu�8��fo�z����(�b�T\���v7\��!h|"��M�`EhL"��h8ϫ�\9�Ћ�\w��4(�☧}��	�9o��،B��H����"aSI���:*a�(;��Fi�	�-G���9�_p�)8W�1�"��ɏ��,�<��^d� ��� ��(e&��.j���/Y���-7s~]���͑e鎽�߻N�%_��sƸ�.8�q�<��v4�~��C�Q�p&�U�<R����ѻG?N:U��X=����ۭ#O��X7���\b��$`q�F<r1�M$��Τ�n��6Qf�8 ��|T>�ax?֧�e��R
_�{�c"�t�Ϋ�-�o����dڒ�)y�RR��*O ��6^*>�\3T�#rR+F<|�F>�Ȧ�ИG۩�G=�xQl�K�m�/[����zrS�&4��,��)8�R�#rD�>sm�Bɍ�-"Í6�w�Z������j��Ĩ���F�A��;3�c!��7��B�>-S��m輁�G���Œ;`�`�QW�EB�D�����9,!k�Xӂ�c�H�ңV���q�Y����HfE�,^Տcy����JPRċp��G�0�qc�/�\"�M2��Q:Ԃ�~�c��&y0X)�c!$)�\���me@μ¯{��'�E���e�%y��T�X#e5Kӱ�t����hK���{���6�/�#:��f���kۚ!G%-�X�UA�O$W�w��t���p�4O*��6���Kވ�M�:�|�ۑ�L�2��m��#[�S�&B��"͘�]�`����a��e�l�+��OG��yϘ�)h�7+p@^3��*�`t�>�"9:��?�Dl
�=���)�f�h�[>X껆1&Kȑ~H�Y�^�����L�����6]��N��=�S������Xת�Ͻ4m��sHqD��7��t	�)�Ux9���7bG�̄�&~V���|		�v�ъ�m� ��m�ٝ�@BL�b�°�^L��kc/<`�v�%dt�k�#��^��8U���M���/�-�tu0����]v��E�~� ��SA��Y%�~����p*ó~ϟ�b$�0�Z���	�[�GK/���mw�UΞq����;���:K�pxw�i^�D�2>gjO��n$�xBu�Q&�b��>�Œx�M������
��b��r�� ��=J8��(������yEh�'��N�n��J&�6�+�����ׯ
~�� C&;d��J�=Ŀ]�~(�&�d�d����i���?g&RN��=��(��9��]B��*K6"93QZ(ѧ��#��"�(i(���Ź���A1"1Ł˔Z�P�4�e�4�a�4J�N���y�2�����x�l��)GO��7@yEx�>�%bV�Yz�4�@�%�uۋ�[ �;7�"��5⬅�������m$�cϰr��x�x����6��W8!rqҙ�6`��2��|R�(O����C�5߅���-���y�
��%jE�I�Ù�r��Ф.L� �Ĭk%�á[P��� �s�3n�"8�tѩ%YE �o�� W�®��THQP�fH�9��M"�M�j\��Ε�VL��u󣌰S��V�x^&�%���D-��s�Zp��� �6��px{5�S����P�>='1iq%����]_�%���hG�.�q5	�B�)��6�Z��B{�Z/��x��6�l;���K��w.r��ɰԠaѓ0�ԺbI�r
����6�:ȥ������������v���ۺ]|_nC[�3����HU�W��i�VjX��Ԕ�e�w�(+@�ju@�=�lBx��sX[�H>5�&{�Ԗ�M�=����}<ݡ�ѧ}~*s�e*����W���j�d�1w��\��dK��:8����j�h4���!�f�m�z6�).EC^F��#�g�h��[d�b��y`t�m�va~pP����D.5*w��׀��k�2!�?��u�c�v��o��Gix���f�r�O#�a�����2eC1_udS+:��;|϶�������3O�`���3dp���j�B@fh�Ć �F=�����	D�Zs_�i�j�'��>�?�%�uf�*����)����\�RI�c[��P����g({��N%O�#�eP�O���W���S�])�N����A���ߍ�Y�l��#��G/�~��� ����2/��J�fz�I�%�GK�g�f{�6�=��*��Ys$��L���V�ħ
��$��߂��C�t
�Y7`(�C��W#֟ٲ51�V4��;����-V��Kcϊ��qQ@M����cn���b��1�A�4;xUwF��d���kķ</�x�!"��>��$���qqxґ���� �X�,e�C�uκ tr�&해iPX�dFC�L���$��bV����U(�F!|@՚E��g�Ơ���2DB��P0�9��J��8��
!��s�Zd�~;?Ix��p�k��,&:=�y&5�]�P�>�
%��@Em������E`���|��R=��(Կ�}4K�T��m0c}�͊���t��}u�}�$�B����d�i'�v���8�@�#5�@|�n����$���1�b���?���"ڇYn����.c��{?��\���HŃ���N���6@�S*�4��G"�@����G ��[e�R�=F����<���FdN��Gu�M��WDR<- �;����71���a�'9e9��4�v�nU�ٶ �Gn�X)�������c��L�ټ�-�.��\�񔱡9��)��}w,���>��O��_k��pt�L��)q���'B"���p��4^�,=^שy�Q�R�/��T�y+�F���#n�K����yz��z���k��1�(Z(����8K���Ʈ�@A�C��&�*���#��D��`	i$�Eݦ@ʡGc���y���u�T#)v�E��`p4�/2�h�B�Nk��;08!c�9B=A!S�_�-&T�ĭ�B5��G�Z�n�x�&��~�a����+�xr�bޢ�4)���=,����q�]c��%��x���}S�hZ�|�K@�)���#���H�*7��^�@�܃�3v���W�,��ʭ	��T��EۗZ-�钙����Y`	�~��R��@�<o[#������� �E�a�2W�`:�L.&&O
��v�qtNdP��5\�1>�d~�(�-��s�Mqء6��T�%pl9��xQ�C��`�+�����X"�1U��*c�6ؤ���O�ӊ��D���]��m~m�� ��К��qwA�P��z��\�q������tk�ۖ��x�x�Qᙉ���{n �4E����o@<���Y��'�Qu���`�u��m�ڢ�wk]��9"6�N[�C��T��cM,8�H� ������w���$�D��u�=�D��O�
&��vue����V (�A��oU�H7�ҕ;��ķ%kWbe�]�O�������g�'�����p����yu�5 $]ig;��d����«�Y$��v3���)�{+v�]��[��<[]sɹ���A�e!��o��	齖�a��&{z���y�Y��ni���23��(в����6K��>�ά��Ý�>±.��ҟ$������� ��:m�ܹ��QUɒŝ�僥� �{���{���t��j�ǡ���o(�r�)�n+6�E��TX㞞:=�	�I����(��<g��e3U��C��F4���W$r^3���Y�!!ʇ
�'���|�7O�es_��W�d"�J-�ܹ�P��S,Qp��v��HC��!Tܠ'S֗����b/�T��b�u�y�'�X��P���X�LHê���� �b�Ǚ>QT��Q��B�`�K2�&'�6�w����0;�n�?�g�h�Ԉ���|�b��������{� �h�I���#,V?W�6��'
"�=ܼ��3�:��Aُa�]�^mF�7�K͉�2��Ӓ9Vf�~a�3�;��Y�1 ^:'�P�`߿�\�#��Q��T1�wo�f�w��ơ� :����FF7"���H�W�Tl�O��\�.ͻ�8��/ga��]�tc��{�૏����s�y�5`aTQh��~����Y��۠��3|s�:AѺ�:)���ߩ��g~���9>3�G�&�t�ڍ�[�U N��d3����j�g��"F�����%�lv]�8���^��z�-xjoP����
�5�dRWC�+�w������pn��k �������.�a�p�z��_U�7�%�� �1�8���U1%�Ld��N1�C�,-j ��Xy�����Wj%�*��\
�6V*H2���Cf_��H\CKPc}E��@�U����ܽ����;+�=���f\3�& ?�ѥ�p�3Ń�f�>ŢͪF�0 R:C��@��U`�3֖|a�lh��Bh䇾n$��ۜԕ3v���~���N˜���p�1�cni�iG�~�@0@��asmj���M�+��7;�]��E̞h��w�%�7�y�뺚�V����p�k�4E��J���d!�N�.Szq��r5#�l��a�1�8�:y�h'{��+8a�����P&@V�X
}ޞBpJf���nTd1݃�-�?�:����.�G��Y=l�����W=�	��J�!d\Q�jA�R� �d,���N#+�)W�����Y�ݙ7�P	)��6��-H�b	-	��Ҟ�4"K$��)�g+E�k����{*d�$p��ø ᬛr��Ӹ۬�x2.:�{�����~��i`X���Ұ�>�݃)���b�Y��D�|1YS���Qo�a^��M����SТ�yV[��
��Me/)�iX{�82�X�Ѿ���?��#'5��ݖ�/|���^$)KW���)#՟�S�h�?�[�m��њY��9�;P�Go�z?���uaFg1���y��@p�C�ǎ�W�	Iv�źe~{ А��w,q����aƪBQ(�ŵ��\��?����"��2��E����+Mb��~��>�j&�(��JJUn�tIvP���)�Ss夻ON�n{F��({S�G���z��"�->W<�*q���������/��7&Q6�ﶟ��V��^�tB����
I���mn����1���T�)�O���U���*M���?�� ^٥�  Xy��D2��!���b`A:�?u�G'I�ܓ|��:mT�)O:C���G�e�)hB�&
d�q�~����\�N.�<���tBlƏ��Y}�	P��+n��J�#�ް)cp�"�ה�73D|z���RV|zM9o�G��_�wO��Cg��(�0�="d�-7[���Sm�%�G�DW� j�OI=Wo<�t�[�H7r-�/�vk�S�
�h\r�c�dQ33�Z�b���4�B���tw�@�n���YBT�3��Q�Z�ii���V-@A��w��7X��}��2B-�n�rQ����U-8~���7W�J�i(����|�]�u x[5[�z~�C�z�y�3���u��t�;Ka��ַ�fP�ybo�w�r�U)p�K�PX��R��'�ӹ�B���o��=�IY�Y4�Y�W��k�]���l���5��8�8ƶ&Oy�.�EfЇ�Rظ��!�&S=������v��FnG���}�l�P��%�F����"H҃\_h���Ra��
^���>��r�Dfрk�\���M���x=�.
������*Ƃ��KJJ}\������O7��9ъ��Ñ�����x����?���.vsǘ���`NA�U:�"4T��݊���!��)[���7f{�=x�㭴��Z��2i]���<p"�WO��vZ�t�����������lT��|2
��T�{��<dP[��DQ5��Yo�ٖw�J����h�/	W���T֧�=� ��^��=��V�q5�g���t�Epk����\�TQ.c-S������Mح�l�uss>��@K��X��6�!\�{�L�����=Մw�^��جR9���b~�m��e��JNM����{C\ힸ3iP[�3�x��q<���V����A8�N/��1��l'�"���~��6x�����Y#�����r�ئ�~�<�(��-����G�:���D�4���D�D	A��xǍ�����*�L��4�|�C�]�Mw,�m-�R��W+$m���q����ߐ��f4՝1x^��`�x:��<�u=�I�lPb�)��s%)��ʿ�k�����|P��]�N��\9�z��2�MiX����T�F� 1>Y��"����� �%�w�ċ�F��&^A7([��}aA��B�?O ����nZ�q��Ό�d,�6�;�A�Hϓ�����>[$3]�8�(\�d�T���|��GQ��$�3�%�+���f����nÃN��b5��1T�
�E���V��=�mWdc��U�w'�]�ƾ��t�cҖ�����/�y����e��*?W��I��R{���Y�r���9"���l����m��,Pz�f��UO�R�6��퍒8���@���M](�����[E�|�9"�F3곗WI��ԩH��`�건�Ռ�m��sl�f�_Eu��^}R�_�g+��Ӕ�I�sO���O��B�J:�T�{�A8x����x@h������������#pd�zN������r2A�ζX���y��h/��5�����ʀ��,��n�֩p�M��3�KoL85v_�U-�_c�l��5�\���`ݖ�!XlQ b]V���S�g�����ܕd�Tfլ1E�T�j��C�q	���l�6�3O���M��O_~��3r6(b��g�O��d��Ƽ�C͌�$��W0�M�C��z��Xi�#e�'�_�����ǣ-��H�x��R,�_��Ӌ��r�܂�Q`��w<͌�JL莻���W�U��K/�7��,�,g�Kƀ�u�$^\�f��0AX�"!�N%���l����GN�{*@�����?���"�J�p�F�׶�/���(\��0q�,���Wv��T~����S!P�����X|l�q�j�&����sl�
�y��F����@ͽ��" -� �Eg�������)���l~ �$�N�z���9b�x�>�7�(��EKڴ�����>6��$$.� �`ץGs��Q9���̛�,ɑ�%�ދ�lǲg5쯨����Ό,cS�U���a����ɳo"�
�Yf"c*�~zYcb���B�^��q���7�u�>��L@˺�f��	5p�O�⁽)u�]
��{ \^��3Xv�	އ�b&��1c���OD
��BQ���[1��us�<@&��{P����D�L]����%��d�Y�Y�ZL�$N[�\;�%�RMy�uT��J.�8�-rK���.
���fD�o��QQ�p���ۙ��E�rZ�M���`�B~I���}W��Pv-����ڝ��g�@�o���x�S�|�!{�K�/�^��8>���Oc|x��r����eꡈ(n�e;��H�LU`	<�Q�炌I^
,�/���OU����ّ�i^�%����tT9.��O��V�>�x�d��GR�/�@`��J�.N��}Y�����:$�H��@�P��"���9�\
3�o�T�c��^�$����PI[}����8�%a���B13����&Id4Q��A�$������=,#ӽ�.������վD�h�n\U�G��Q{@9)m"f��F���?ǖ'r���rχ�_�t^�ᤎ�z�MF"@֯���O���-bN�A��l�a�K)6.�H�G�X�J�т�b/9��J�U�Y�jtW~���[������pm�����RRQ(xI���]cGo���q���I��5>���{�����Ot��Bp!А���?:�:�KCp�*�+dwP�� �>�,���'a)TiEx�>vOg[_!l+tՋ��F�_+�zV��5������ʠ���/���G��U�`7�/�ZG�����=B�<IT/��@D����X�KI��]9|G�tA�G���9�����O��[����b�^
Pg �ˇq^���~[5�#
���ٽ��������O�3�x9� _)1��Lȁ�X�s�g�}��3����ƪf�1�O�`��擁)�A�s%ـ���RT�_��OB��A�r�_'1�[�T hE� ��
�&�T�Μ=�g ֞s��+�ӣ��ab
Z�@,R �3�λRs�7Ȝ�ԣ���I1�ęr�@�	��a��7?�mj��0|�8YH��.���Oi�G��#극��Ju։#/ߛݡ\��޷0%�~,I`�+	�H��AH&=0Hϑ��Z�������4�,UI�z$D�Qk9�����^?.���yF54��*��?/t��s�A�-􌥍$�mZ�P~�E�O5HF0`��> )ͭ<p���E�#��:}	ȕ;���r�mAݟ4jP_^y��׵:�~{wͱ�	���Xu�`ac�6sX[*!�c,�#��]��Q�c�o�o�7~�����[M=7b��NE�ސ�x�aɆ��ˬ�d"�h~��~��n�쒜���d��'�zi�ţfn6�����t�U���.��v��V���m���P��'~V��x��������i=���6�W���-MrB��({�s�8�<Nv�WI�I������[C<��:�ΛB�ޣ�8��S�*�Y�v�Xr���;�M0|5D�q���r�B���32�jL녙��+ـWQns
�p'O��*1F2�葥
;�\X=+�(��K��S��_��gze�&s	���S�
̝Ȓ1���#�_�h�(�FSu����^W̏ ��:��e�Ù�y�[À>˾Ԩ��b s��D#�u��A���N���ReQ�E�h�K���%�Zd 9�M���}x�4>=��v=����ᇢ;��_��"/�0�v��@	j�F��j� ����G��ʬ�Q��3~��q����Mp�;�䬜+Z�4��+(�*ަc�N��3���?Z���U�Z����k�1ҋ����V��!y:\��>�Fu]鿌�ګ�W̚�:|��%rykǈW�>\��)���.l���`���%�q�x�r�~b�1�v�Qžn���0w�Z|�����$Jh��R����pADY>�ʆ�yJ&��͞\V��7^��'΢�84��V	�����z�ь�3�Y>*��a/�),&8�]<�fEf��`E��X��l �k�O��OT+[ב�)��&G�苕h� Q�g���h��.���ܜ���B�*cm�@am�^�N��Wܦ	��'%��Z!��?&W8�įHÒ���Ѐʀc�&� 5�
�(��K8i����~������'}���]�xD��3���F�<�h�����06q�83��g]nE�|A(����2���2�
��,���Q� Ω�Z�tS'">8�(��;�ry8~(ppi?�q�\LF�@j�#���)6�M_�!�ײ�ƞi �����Z���r�R�4�Ӊ��n�Z�2�) �yM#����[�ܲRZ��@󶃐�e9�9��g@X?E���1w��bq�`�3Y4�;��c��\tϛ{�����x9�Uˍ}x鈇5�Q���K��w(���vw�p�1���E�8՗#�5s0�b$W�=Q3l�h�9Ne5g"nm���f�܉	��q@��D�s���x�`A�?�������u~�y����������y�BS
x��=8přS=Ƽ�n
���&���4�L{V.�B��pH�b���0yt�VC�0���u(�d �9�)^UFČ�uL4j��SڔT��$��@7;�g}l|r�I�"�0�ya��FIż��ָ��eo�\�b��M��|+Pw��$��vW5~'��pȢ�\�f�������)��',�^���֋&Q֜����V59Tc�s*n������-3�*i+`�Z)�Խ�G�E2�O��ɽˇ�v�I�Y�Å|Uq�^y,+:��p��o�v8f9�[S��U�J%���nQǈg�R" '`(A��uG��x��3�m;�=�8`˯�5��|BG�"դ��p������O�ms$���h��I�2�8��濱ߏR vIV�5 CFIAO�}����?�E��N�)���e*��H��i�~ ,i�:/�F�B�h(ǹ��B�e���>	W�[وx%��5�!����`�R�Z������4T��&�s#hy�x���1�m�h�4"�$sUW���g�"̧��S�=6�/�|]JÙRR=� Y��!9Ѳ�mr�(}1����r�V:�e;��~R�fp˸|³p䅖��D��)]��ԡG�	3[㨂q�E�1� i��cX�9*=��n4ɐ[�ή�zn��b�kȨ��T���!��5i��p uꀩK��� �!��~�{���:n@u�sA�������f��o,��f
oM溴5�t�曊���*wP6��*�F�3���UʤP�u����\<�7�3F�����B3�0f�τZ:s�G�"376�d��̸J�R1֝��������:X	E#).fϪ��0ʘ�V�٬��!Z��4&_W��\#�C=�Ƨ��`�v��B�D����t0b]t�0V��n(�_~"����0�%)K7B3ǔOB ��5�[=F�M]��v�����|����ݦ���:���cJ��,���v!��fR��uY�b�6��IF'O	���m;��2z�.h�>��-��Q��]vI� f��~d�F���;Eu��&�	Q��J����0~5�Bɒ���/&���k�G���A��O|RW�V���V��O{,�X�jYF��ME�F�e�ʍe�S�7)�����^������T����O脄�����I�!_�-�Z�������n��e�!��\'�#�9U[1�,׍�mʛ~�-c5�:krS�S�\,�y~U��bC[88� <��Ϲ���)`~ka`J,q�r1(��쇆�T�����8HY 4S�ՀPr0�����4:�6�-x�,:OȤM�5���[~�8�Ę��F�#��#���m��Fj���.%��Fo�*�
Η��@^]{����fr�#�
�S�&��2OY���Ot�]��޼�n������%��Nex��#"�`@J20��l,��H�U'�Z��������69��}���M�P�ul������t�b��K/���;��挄��j����^�1�x���4)ŏ�D6[]�5��MGP�Z����y"���L�Ζ(#���z��v�(��y��C�%p�C�	`!�aHLV��8T���GXǱ��8E*��ڻ���Wt_��|��K"�qժA��V(�vt#�^�{��:f��Yؼ��J�>z��l�J�=�[�`.~7G]̾��[5��~V���d A�QP)1�V"g��U��(��o&,Y�_:pa��ޮ��[K��:� JIފ���a<n�����P;����M�嘽Q������	�.���I���~kq�3��Oh?4V���"yk'�{��`�_*��^�_�]4^��A�I-ȅ�.$$ᆗ=",�E��@k���&�D��O3�0VTqe�S�aa���<��+&T�Z��**���(YP�*�Y��n����*����8��}y9q�����E*뷟/�%kT;@�?-��nC�y!]{�{_4��o	R�����2�"ZwX�'�	O	|���d����T�v����wa��47�c"������s]`/l�	*�����W�*���1f�k+�BT�\,8�;i�9���������c?�x�u��6;i3A�� c�*�vI}����f��nH�s_�?�6����g�
n@��i�

m�������s�eQ�|��.�����H�ӻ�{s����](b� ?���L^�K��Z��Q�.�P�%8��7��HNN����g  ��<`�?P�y�(�Wn�dS�!�Vyu��ܿ���U��݈7����l{�:�{��A`��F[5�Sg���t�[�׏g<c�L3(���H�2��|}�s-���}&N֕�Ah
25��f7�+~������1袦0�;[����$��JR�c�m���Mc Cʰpb@,ɰc44��c���I�G��ň�_x��w�g���� x�.����e���!�	�E� �9��V�P��1
�7tuo��~9>GEF�y@���"�ۿpK����h�ҩC���dJ H����5�!�����wI=+���}'M	���uO* �(�#m�����YZ�>��-�Iǁ�x:�&�3$.E�P�O������D�����Ʌ�[���DX���5	=:՜T����U�2/��/��������8��aZ$0�?�Z�	����˘xJ�d����y��y��<���ߓ���b};�R�z�{�o�[��$���8�b��'C��@��2c���K ��*P��0�=^�sL�~H���S���6�%la��_�OY�|dY-�夈�=&�=S贀�+�T���#���?�g�k�y<�2��ڄ��9��\tC*'�[$V�S�ɡI��f��v2�H�5��la\ӳ,D����	^E���kK�r��}�k+�Ec�g���x���?�6:���7OBM:8�����;�U��3�v�Z*]�+04��m�O<k����E�)�OXGc��T�9&e�(����M��ظ���볼��(���������e/���m�t,�Jh$��*���%�����[p@�7#���������%�W��N�Xe��	�M�y>9���uV8�
m�L7W��Lv/o�M=OMYe$���hyH�{|��u�����!p[�8Ҡ�TJ5G)x�b\���tH�Vu�0q�X5�D���B��T��\MM�c[J���/G���{�3:�:Aژw�>	�#�4���3^l�=��K���/��S�Pc����"��p�v�]�ڐ?�Q<]��q��lul�i�Ӳ�⠐%:�r��Nl�n9���f��$����N�q�̇`v�����lK<ަ���N��;�$�i�x���2`QRU+��A������+��dY�^U!MT�y�su���l���g��V�'�� �D)f:��uL&*''$?4ƿ���u�ih�"֙����^��c�.pVxeO�[����R)��o�]��e�Q��C2��?�/k��{�G�{2��g�~s9����DK�R�UȲ�d���p>���E�@�v-9�54���2��r��]��XIK^u�/���捎0y�g��*ѾJ�hh-�S}O7�I���?���~Sus��7�Tç�$��)�m,���e�e3����~7U� ;K��cb������ˈG�k��3�����Vt��Z�k�i(��d�hM:�\�(&�?Q��gf=1�1�
���U��}��ؕCp�3B���E��20Z�ɱ�N��zK�Cdr�M��X��=�s$����-���j!,�w���z�{������1�3��8�e{h8���^���9�1�I+n��z�r� ܊ w�,ـ�W��f�3˟QhÖZh��T��}�l��nT����cszYg��op
W�<7��Aܴ~�p�@��?��L�Ţr�>u�B���a�'��@�h�O|��X�(�,�[y<��XW� v�f���@�: �G/�Џkѥ.�p�t��	 �6���rE��Jo컷�t�se���ee�m|�`7�t;k	��#2�X�3ѥO ���#��A�7���?�W�g�����v:d&�Új�#	fY0<��?�����!��; ��4���:�GI�"b�	�4t?�� ތ��O�:
��v���ƀ��@�����m;�~�@�F�8���e�{a���Z]icR��.���ݔ>�P,�w����Rr
��  $%>g����j�DS�Ph�a�ag�\l�����p��O��O����OE�dNߡ�̐b��(�٨���C@4��ٹ�F��?u�,��us�"��^aD�Jc�tL0��ۇ̠�2!�)0}^�OG����{��S!T��)�m/&Ut-����5����W+��V��ş�M��Y�h�4���BU��&��+�4� ����V�������R�½�j� ����-����p�����V�g>��և��6�H�?))�uR��x2�6<n�ɷ���l��XL�f���J���{7V+x�J\��AA^g"ܷ��D��֔�#È sѺh�&qO�Y��h-���d��$�bx���L~K�U���x�W���~�PP�bҽxc
Ml���� �0_�KIo�r�b�R��Y��\�$��f��;`�Rj�yC���ǲ����zM��K���)��|i�%�;Uw�#1%)��AjW4��eq��ʰ8hF8՞�`٩�"O���b�g��?�t�{�R��d|�+�!E���<e΢�8������d:�x���ݳmBM�b�f2 /��?g�j�ԥ���͕zK�oG �<������@�,֒R�b吐ʁ��3�r�j�G8%��C�l٪i���X���;����}�5|}ը�{�� �H?�t*23lbG �)�/�z���r���h�� �` ��IM�唀 w�#�M?�}QR���H$���=7��w��bS+��Ǒ)C�z�0
�v�L��K�"�Y��v'|��=�Z��b�?9{3�qi�g��p,PJ��xP,vy��kk��o���˫d+K�*]�G���߽6���K˽��K|ߒ}5�ku��$��c_���Fإ�w�ST���y��%Fa\��o��IG$gu}%r�)�nG�v��d>c��M�t�̥hØ22�'��<|>��q���X��ΤE�c�|w�~�{C�6��c�r���۞j��ѝ�eʞpwdY�:)I"�ީR�i��J\9s�;|~Z��p�d6}F��ӄ�w+��j�O�9H`Ğ��gK�ĝ�/�cJ\��^ȍ��A]+�q\���;&I��OS���i�+�E�h�{��_%h�c ̪��-6x�#2�(Y�t���exÔ*M�3���6��Yҳ:B��N4D�t�_۱�]`0��g��cZ^�J�S�v Ʃ�;�!��wo�����[/,��&�K��.� ��Q:��Ìz�8ѵv�W�s(%�7��&2n�����}����K���| ��>�A�j�1?��=|/;����h�ڧ�����������e�(���Ի�̞t&88s�H�Cj[����E<�!Jݩ>Kh���7U�q�P.�<.}�a"����g�C��T�#
/��s���ﷅ*)ޟj?o�c��c�o��"B	��6����7y�_׎(Iu��"?���}�����1�~��`���I����`!{|0���Ԗg�R9����ҊtB=�F������~Ӥ=�%-�Go8�^5
����$mzĳ�r���_o4��O�DVO�}����Wr�h`j$����t��U�~Egrڡ3�hD}���Ħ����<OtN��5����Z����>S�c~��+ �O� �8 �H�"�-��!d����}yb�$A�����so��W����%���/g���~X���ȅ˒��"�&�y^R����	�`ס؝�N��l��?`yܼ��!hf`��ל����Xb�����%l#w��ԯ�4Q"�f҈&��
-� �%wɷ=�3v����7!�m�O��l��W��O\s��
�˰��Z���,��`ں��O��-�.��d�˽�O��;>R4�x����d4�:�?j��+;�wp,���:.��@#-r�ZJ+�%u�a�� {= k�M<�LM�	���醴��M!Xd�M�'I{�<���g��d8m�A��5A�E՝�׹/L�f�HuZ�yUz�Q�5y����Y�D트Y;f�O>tQ�a�K���&��͹��뚡���w$�(�} ȿ5�hB�1ob��/^�}L����?ޓĊ���D��v�x���IH�$���h�;�����G0�:'���Ay��5�4��+�I[�3��p�!�~�G�0��P�7̳����_u����.(�Ќ��/�G"2��b'c�C�v!f|�tv.�K�ab^� 7�K*����Èy�y}J�C����ڢ�sb��~MÀ��������Uͺa.���f�1:K�j������qKS��-������!�N �G|
?|/~�D����V�`1}Yk_d �)C��
���99��:�q�Th+�my9�/�5,�ȮݲZt�1�@�N:��E@�Ҋ�<t'�2q�'�>7(�TItjq�K���.,�	����&�{�W[Ip��%�y?@��3|C���1�����r�6���H�i�y�.T�	�V2h[#�DD��iIy˃y�Vn��BS;'��֓6��s�������m bm�*��NT�e�a�����L[L� V���\Hp T9��n�����6>ō��/���Q�H���N� @�e��)�Hğ{��Ѯ���>�>��z�yt�ǔ�ծ����"��+hA҂�SҸ|�����nFq��~�  �?�H������hl��7x3�)���A�Ϸ�	�ٍWl{���zo�  �3���+��3���6"�ퟧe�c��������(w�G���4Ze���'
���d4:�����l$^Ќ�,R�J~��\ԁ��-�=��m���3���A��G6��H��;��x)�vY)��,��5e؁�w�Y����w�Wƾ! �5�RU����^3�j�ܔ���Se��j�x�8�>�nGH���1K�����M��Gs���<	NjUΑ�:����/׋�H���h|M.�r�T�Q��GD�~8���X������R�H� 	��5�an~51��E<~���x�d�ډ0�{^�9���)����;��Nu)��*Ɲ�������v���Tfࠪm��P����M���38�Bu�7+��@���G�1Ț��^�B@x
�'��|��s�hm -LK����8��i�VMM�����\��uIG�=�30������$���/m��!�|�=柠��s"ؾ����=
�M�!���n�-v� �&���)[�pqh�I�p�Ы��%&d�u	����sԨ������J�v�iu��	�P��ouv 5�T��Ĥ�����5@Y���tB���y�-��<ס��ӱ��|��[5�5p�ަ�N�,�̇r�k�R����{	�nd�r��h&$zpt�}�V�'�9�?K�P ,q�0��8Eߝ�S&$�ף+�X�٨�iG�x���~���~��h'N���UE���
�S)����M���l���BD���TK8�_r #!���w�M��}^�q���>���Y���e3!W��%-,�If�LC�m���.�0�^<-�?��X��(9C�R��t���nTS'�%A�G>4Y���'T�r��4��h�yb�1Øj������$��!�ř�)r�?�v�M.�G>R?��f��D�i�#f�z��7�a;�4'�惟�o�`�M���c�g��t����;+��M������/�����#�C�rD�	�t0R�C�aO��.Q�"���/�s�`(��U�l��5�A����L�2���ؔG�:����O�7�1B�0��K�B�nMB�9���ROt�|���:B
w51Ʌ�E�5��.��"ɡ,����Jq�z�8Vo1U�Q�š�� |@<��A?,�lTwF*&�΀���~c��-*}�����#�("�e��
q�j�n�:@�):"�0=ӽ� ΔAG(�e�l��r���q���iP�t��.V�IG�i���(����'J����~�[ ��`�-�J�ȱĤ�Xgtm������O����Ao��^�w��ݺy���6�0خ�n����bqTX�T�ѧIK9L�������9/',v@��'P�����MA�|?n�L��X?�bg��,^�t����mt�Ƅ�~� ~��M,���m�2}�3������:M���O�.\���7���x��D$����%P�� ��Q���R��I$���̏�Bϑ���+fY�k3����'�G����~��OO�rV2K��	[RB���u��@��Ak�'�a�8q�2yr����6�SȨx�T��!������$q%��q�W6��`n�zfɄ�\S�x$DrɅ�p�
b�`H�6�f)^e#��>sAR��%�U�􃩴a�Շ��T�Ɨ��5����y�9ވ�kl|l���P�d�v�&�^e��=3B�~��1A���]���״t_�e��@,��A��,��qv;%�|�bz��9���{�P%l���'�p(ung{�ą�@�)��6���GQ��i�LI�9���0���l�_Z�_h�"jҗa:`���^�х�f�EKk}��+¸�2�cON=�zl���������3�R�Ȕ���E��ػ�+� ;"Z��< �;���1��@;� u��̗�2r͐��%��߿��O�ƣp/l���@*�	�NS<���1�t' �oR���F4
���|e�H�=��eֳ�&fp��,� ���X��m�
�{b��_��r�s䞣�`c!��ϣ���)����xI<�_'�Zҝ�� ��ڦK���ǒ�S��������ճn���p� j%��YT���Q�o��̨K��W/������ރX{�NB�(31��?�����	�>�u���� U �#<hژ-��'�s��L����H��(�����L�N�z�"D�������-���*i��0-y��#����Z��΀5r�V��'>��	 =�96
Ş�h��'nE�i�-��P��S�H�	����j��@�B��{����#X*sX󖖑�����v�y�.M��_�M}#6]��ĕ�mCMj?T����r�v�O��^r�Ή����|B0J�o0\�.۸��މ����K��9}#�p�lͥ���.��4�� ���fX��ڱ1��8NY�=:
 �]��,��
UI~�]���;�E���֟j?˪����L��f�9~����+��r�8_��?DO��9#��)��ښ��<&���>@�2H���w��L�E� ���V��N��#x�12W�07�_c��J��$�_s4�P���	ґ����g@�YJ]^{w�7$���E'> )�H�/.�����n�D3_{:�CuL�^
$�����$醞+2+f�34�A�Q�jɑmi5R)]�Ŝ'� �������>5���E�4h����K%��3G�	��ڛ:#�:J���[45��a{�[���P��^��}ԩ��
���/Z2�~�qvZ3|�.�p��o��f��ʹ��N���U����ovm��$��f3� �x:��`&C�%�-���T�<`nw����WX��0C�	foAX�E�  u�a}���Ue�R�����CL���aթKm��w��x�����W�͟�ހF�o]pM+���O/���㌳�3�Yk�pE�>�7÷Ȝ����Ŭ��q��|��H6�nD:�� X.��0m@��, �%s��`�	�F�Z��XqpC9t7�iKaf/~�Zde�w4K�L�OdMp�sD���2���C�I���jhu�ُ]�\W����!O�M�
�t���ɗ�}F�S����_M=�7��W�5�f�2�:j{��f�^�C����)t^��<��LQm��!���ڱ�����R�e��^�s�hp�o�9�@���|,����0&��Ja���Ԕ �_B�fw�i�A� ��k���&r^��UP��{����J�"|��E#��Fv�Y�i���XR;��a4��ͅ�����W2(��փ�"�Ew��/�$�!>����R�U��<'�����4��A�ٛ��P�,]#�A�����)|�®֑��
�T��d�¦Os|��E����ʲ���������r@c�ͳ�1hS��257bʝ�*Wn�����*[{����YI��|���/��i.��X��JQW ��F��dXT��PfLL/a��碦���K�x�Ը��k��'~u��6�s��b�6&�*��ۅ�*r#��s�F���	P��	k
�iX$���{�<�H�P���?:��˂1yfx��Լ4) =N�.�9����f��W��(�DWh�� :w�d��_uW��g&ZBݡ	9	|��M������刻v���u��mJ������j�Y���v�V����~�\�};���*��)�!u�)���
�S5*�sǡ���He��ؓ�sC���#k&�G_������>����P�.�ÂchY��nn�lߥ�(�c#�>#��'u	o�IM-��G�k[�֍����Y�}��l0�K�G���m���Z؇�N�N����>�5P��Ϟl�^,�z�ZRM;R���C^2�����zzlG(����pwl�mZq+�EY��/	��p��m��S= ����S9FP�.�tXa�o�vmMaE� ��p��|J_�K1�4Q��h���󏤑|7��A��ЮtrX�\�W`��8=�ˆ�p�p�)��S���Ԅ!H�n6*j����6I?z� �!T�˓�E�5�O�H�i'lgK�$�cd0��;n�`݃���(vZL��/�6��P���Aj_2�qss�wQ]�{v~W��|Q�X����m�k��cn[N�4X���ѳ��$�F� ��"aƸ4 �&_��_�ƔKd�p��e���6���Y0�P��N;�r��Ϝ�� ��7���`^�_�Q�0>Ga!)�A��.����%C/=9W#~x7�yA�s�>@Z>TK�%�>Ab.
�s�_7ŀK��W��o$�S0M�����϶{=�A��\7�W8I��y:,���n�c�b�e�Eĕ��r���t��Ǘ���͠�:۟�tE:_�������poX��2r�=ƽ@��;o}[W�l�S�#�SV�/t�N���������˄lc��ਲ਼͗��v��yf[6��
��M�];��[�������zb�\[��ڏË�\'�C�$罙���e�P�u�~��hx��sq��2��9)B
f���ǥ�h��1��w�&;;.��!b��J�H+�o�����AE�Fk��;ZeK%s�m\��}���̜"K}9rǽ\�>fc�pK���9r*P�׌��3a�o������X�X7��F-�t��QWYk�?l`12'��ڻ�	�4���:0�3��Hvވk��Q|�F�2ߓ��7���{��d[�������tb˒g������ oG��rSw��\�Bb� ^H���I�F
N�=�2Z��U��Y�L���+����0�������.w��G6ur�5a��,�mbS�dR�l�j�r�|IX��G�Z��n_�|k�L}Pt��/�d,y�+��ܯ!��%�jB���r�h쐰�:ky��4Ҹk�h�.*��Wk�}<
0H,kCjq�+=>�8�r��O��Z����=�3�"fx�1h ������Z+l7c��ѫ���2f�s��Ka��P~�=�s�J���'����Q�����um%����>�F
Eq�@��?�n�[������(`Z�t�%��I��H:'M�a�8�Og�4�^���f�Fb�`-���\+y�S�_#JU�.�$D�V��/Z��i��+81*�b�?�I#�h���5�~;�n?�4���}�1:M���0y���'�ԸZO����u�q. ?~`�-�]���X���%��Φ)t��xi��J���qb��8�~�z�TM5=6My���$@�r� �i:�@c�EY֘���.�vV�8-������ [2���dd}TO =��)^�:����U�˷�%��ӎ)��ɿt�q#����J��Y�uV��G*�)�W|��׾7��\��:?��b�u�p�NuC��F�i�m��4��;����T^�,��QB���12�oeQ�y������h<2i����Ye8�I��h�DU�GZ 6$hc�5g6Ҙ����]u�U���=\Cr[�Y�j���m��L�9�\�b���/����r���u�A�5t�1���8��U�,Z�A�JwJYI����L��]��	�f�@��
,��a>�K����3~J��������4)�!�9���s�n��5Oʎ���4��*���cL��?##m1J�������x���,6~�L�y�h��7��g�;e�xNZ�%��L%g������%*�R�ϻ�"���,<
@i�R�	[H"}�}݆�P�JFVܢ���'R����~���#E��m�Ά�IbN�[���B���?��,��5�=r��d̑<��C��/�s8����.�t�7	?�J3�S
�u�U�4���缲=��Ǹ�!L�W�,2�����H��k��g+蓈:�aZS���
|E�e/4�	p]�m��|�#�mg��/ƈir3X��;�6C;m��WTǳ�2�,v�G�����ƫ��c��m�H�8'E\^U�W�6�t��-C�j-AF�@i�Z�cJš��r�&��)��q�oCt؁����Y�^p�@)�E]1�P�
Q�@.uC�����C���������m�sb�&g*d=2�R�"���K��,�Sn�ve_�M��b����^̠�®�F�B���#�c����n|T�2#�pG)%\�ς�\�Z�c�g�,j�LH[���ވߢ+��D�NJ	�;�p
�B�	X��}ȥ�W�f�.�wO��H��H�F�@3�&�RxR���|�N�#7ʂ��t����]�/��zo��W�,ّap�!�r8#��.K����BevW��Y��$V{Q@+�[���B~KI��X{�P��;�$vۖ����s�	��b���"d���ll$�|��/��m^�0�e:���}z(
�]{x�̱�T$m2���^�/<�Sq���CݰnzpN��κ#��@,�ƺ��_�6�_Cn�)����o�'��s�C=���06�s�Vb���Vw�*c6�j�J�X�c#��uu���M���nŤ�R6F�h$�8�r����c	]}�����I�Cӱ>����G��x�Bs�͖��p$�<m�Z�R�F�#��?n9�eS�^��Fݸ��-��fi�����V�l�^����;�fP[�D��-2�}��dwF0���[�JU���O�c����u��>���������4��,�r8q��,��h@�<�s*�g�ί�8�`����=:�G���]��Y�i��W}W'��n?>I�W�~g��R�#̅h�"n�M�{Hr�H���tQXy~z��N3��!RX��U\w��v�g�q���8�ʡ�4���-4S@���d���Z�o3���+"��&2դhG��WQ�R<��Ď���@�k�q����ϠB�O�.�d�p��q��𿖬#1?��7��X���VU�G�ם& ��f�#華:Ň�Qg�2Ϛ��R=O�,���x̲�Y5e7*'��0��z�<�2�O�ʃ� �N���^���9���JS����6�=���$U��XC�Yt�Օ����@Ew;[s��� ����k+"i��MB�s�f?P[I�}������i_h�?���Sŭz���k'WN����R��W�4�4�:��cp��OG�
_�/�;&���{��CN�9���B��uΣ2��R��Ck�r4��y"<�D�5����[С���
�ٽs���T5��עz���M��5�!j�2NvX���¦�@�d��7��sY��~��3-�@��U��C<pO:� Wp�V�q��
��$p�VHE`���ǣ��k�sPMQ:ǁ��=3 �������N�d�b���ڤ��
qz�Y7<�YWk��8���s-I�D�B��?"���ކ<��3�,�9Ɛ�w�4�14�L�ߓ�{�Բ���T�����J�⑀jnU��s��U�i���O4�p��W�j�Q�"V�Fb:�j�BM����ED�JBO����w7��T'����3S#%9@��A��[.�V�A@��a�4H9l�$&.p��.!&��VdG��ȳ�¢�'zg���L|�30rbg8H>H�I����G&�r:_��׊�Y샏5b�$��x�$,@%J'TlW����J��.�L��b�ah�߻߅;��R���z����?�d0��Q�O���T^zP7��KVB#q1�6B���rA�3�8��%����������X�+'`g� ���+Zm$7Z��b�܏�j'�K�~࢖�}#H��������y���dT�jw/��� �q�E5��d��Y��?J�;�}�ˬ5��.O�p�����k7+�"Hv(]�Bl�P	�
�F�J�%��K������@�	C �����I�| Y��X�g�}�Lh8-��G�0�Ԁ�>Ց2��!��$������|HK�RW�\��S�ĥ�-��]��l�썁��>$��v�$�ȱ-�l��*
�d��N�X��v�H9��)K۾�g�6��x�m�f��1~��v3@p�\�F6�5`���#�y�R�O@u�
q-0�� �&�椄��5¹��3?�]�kfm�ګ^�w/�����)�8�)�Qo�U�ơ�������v%�JƂ:l/v 24�����lec\��ꗧ������&5p.� ֝s�M " &�݀4ge�e������6�7p�(Ud�����)!p"p��Q)ޅ�����̭��VP_�l<�TMX�'�"{]ށ�#�����(גv;�X�b� �ޔW`��C�Hf`�9Ny|�������9�v�cu=̈�Ǽ��MĂ�T~0�ع�F*�`!�ڦK��~�bA���ߩ,qH���%>�6\����!��*��v��w��Q�����'�4���-� !��%O ;�֚s�5�HUӸ�Tw&QWŇ��+n��a�%҄<�����j����+�A������>G����0{���f~�<�2o�+�'���� 4��r$���}c��]�1A֖�p�S!��zc"��#������~8��l��6�0�tg����e���"�&s�X�4n�[��om��|FGW���x3�媌�(	�ɏ�qZ���j���kN�����K���k �*m��j��4��);u�?��w���ڙH֐��_��j���똫�&5���+�<�X�8�f�`9���0����J�A)��96�9�	�#����X5��h��e�������+n�U��}-���S-���W�P�C_C�5F��m���)�W�T·D�����b}���<��vT��[��5�PB����ඛ�ӕ��T��-M��!��_����
��9+�y��yi�}�,Orm��U*�vM�"�^�*^�]�Yq*���	%p�I��ͪaC��Q�.��➉���ޤ/���w�1;�}r��E�7��/�^\�w��M��皋?j�@#sP��l�!��މ(����?,�.�.�4��u��EڸkiVh�H��rD�V8�o�8 u�܉��4��W�aH<{�,�|��+^.)"H�<�q᫦.��X���hm�^n�-���C�b1E�']I>V�c_GI;���Ow�Yr�n����cΩCd�+�\#��8#��c?s��h�H��˛�����=���4��6�O�^Aل�kz��:�X�D[���\�JW����yӮ$�M��`��ʥސ�>+@�)�^��� �{�L5uF�V�H���$�D�t�bO����i.;]�%���R�������V� ���d���+E�`�1��	�K��3�2j��w+���$�Y�ݭ�������{b���w1[}|�/o��^���h�L���U�`�f�6 ��?%۞i�p�/�m�����*�Z�j`�ۅ���ĕ<8*�yo�98������<J��Ks`�ʣnb�GJ�L�V��՟C��߂���i1�4K�J�ի�����(T?_�q��ծ?��a�T�VN�D��)��$��A�w�����5L[n�N	��B�v�\G}�\E`=�MP���0a�Ry�p?�z=e������Ac����$�,?h0	��o�S4G�}rs����J�$]�r��f��z�!��&]]-L@Uq/��Z>���l����hD�����/��|��,u�C��2qC����'�/`2�ܺ�e������3u3���,B��[�͞Q�>2���%`W���n���dy}]Ȝ�������J������5'�Mu��D�m��_�"&���fz��%F���M6G�ڵ�+!������Cr��<���n�
������U����3zl"-���U��0̶��x
�14�����YSݿ����4\��I�t @���É[�x�i�Y�C��,�Gy�rPi\96�+�� U�>3��h�v�^��m@L[+�ُ�Z8�� ����\�����>���o���),���d�]Wsc?HI�ֲ���N�ڲ�iT?���p���1�����g�݋v�u$������l/��Ƨ�I����LV4�F�� \��z��&gn�����~$�D����;�����M]�VY��)F[�O�F�����\��dy5r����j*��}N:�ͫ��4����zS�%��|>�uiF<�����j��g�3qa.%c���ehC�%�pp/m��c?�{��{^3������1��h���R�`��v�:o8��_J$��+��
���%�G2e�Z� �kE��*a`���Q���Rh|����a��װ�̚|� �Cv҃���A�?tЂ�m	��$쀕	}�����n=Ae�4��r4ӏ��iyЕFkG�Ȫ���.X���!EQ/�=�N�(R����!���_����_
�zU�j$na�[쩁
�� ���r��װ�oD����|��l�2w���h�-���+�Mȅ����~c�H�\�ٺ���i+��MeoG�Y,���m��D�0@on�oj����ɥ�s}q]N�W�	T�`M��B��jh��� �o{�t=*�(��ݵ$�p�BMQE�L>�	a��b�QNz@I՗�f�Q�ٹA�LYz�ڳ�kz�.�ӥ���֑J8G��6��?�|6�1���e]U.�2ȡNlj��f�9q��H�CHҦ�̆�������g��`I��,��:e-��7US� �+�D�HF�,5����G�O�J�R��kBz(�h0��,��1+�Bk�(��*�]�F_jq����K8e�9	���EmC�(8qC��X�'�M�PV�Vy~�� �̔ݸ"M&�6w�l�v7K�2�]}�
�fK�wr·�Lm)��o�P��5�=X%��k7rH�]FVS�{tľ�d���_��e.�<��q���ƀ_����
B��8���=�ﱯ���kO�{9���kڤ���v���Y�d���au21�\��&�,B�4��@p��q������68��2��LN�s��䧻��`N�;��e$�̧�L��VW+�8�W��M��H������V+�W�X7�5j����\N�%%~��g�ԵR8�%�	��N9��=i�p�W��0짌ǘ���wu>	��Ic�P�7��\����#<,�_�D����f�0�j�rL��o�����hV聥l(p��!yR��ջ�{�κ`��]�Q&�:�3էD �\����}����!�GP��1\�9�sdډ�L���o�C�ϼ�6�\�PO�f���H�]t�G8������ �i�n�^��r���L�tyŝhQ���L,n��V��i�|��s����^.�O>�Y昅liT�>sT:�ZL�ˠ©�H���:�Xq�c"U�
ە�|�Ǚ����ogD��brc38Y���P� �k2Qcx��m%�м��
l�ڍ񢻭���PD����\�:�Q������K�a�k�A��׮���������h���ۍ6n�y*Y�fk�ɪ���?��س{�͵���o ���X���ΐI�MޟI����&��<P#p8k zu�`�(�
�å��M�p���]Ӧ��'��i8�|�y�����AX�t���$�UT�Nt�3DՙM���U ��7�:��į�(ph�_ٷ����Y~ӓ�I��\$�^"\y�v%h��9&.=k��@�>83�$�_�]�}ݻ�˳&1;O-�r��b��Z�Ct6�>\(I�x�)\ԍo߃�N�+���=��+���-�U��Q3��#���lߊ�Tu+���
�Xzj��̠�9@����^�ơI&�W���L�e�5�f�D>�,��G6�+�H^_$.�滭K�N ͻ�jF7�a�4����7�}�Q�\�D�*O$#f�e�P��NjL_�s)�G�M�z����c?�_2�b�a.Y9�0�1����8�,8��8��&�5}�����ū>��>�j^i�<w�0�)`�H+�U�c���i��m�xTA��-���W���hM�j_���F�w�'��w��)�ݝ���'��YmmK�5+�*3/X ^�m�j�_���E�����.2�p����x!��-*b`Z�4���'GI���(hAn�����P��!�Xv�s�~�;C� ��xy���g�Df�t���������=Zv�@Vr��4�Ի�
�)kGY��
�s��XW�>����ߘc>�d�P�� ���m6S��ש��^8��:	�`>	�z�t��`�2�csZDoO_�,�.�=l��.Z7oZ$�;q��[���fO�4³�v�7@zh��?7&�Jm��XnWS�����n�0�H e��*��V������w� )�S�\���܎�!ڈ��ئK��ƃZ��3�(:�]�t��)��1���	:�#6�{��h�ϊc���F���6�-������R�_����j"�@���T�D+x�e���׸+��+����X�i� n��(�oE8o��ml�</��?}&\PNc+��s��M�Aj��n �q��^e3�~�.hc��(����Cy:�"�*fx����p4�L���o_�e���^�Ͷ�6��hS֦N��� �A�~�u�J~&$ٴxd��p�Wo����R���Q��X�s>Ke��SO1�V�n��uh�ͭ����13��y� ��g�zK��+.`oj��a�/l�sZ�VlK�9��^�;�@9�ȳxi_Zn �Gm{�a�F �T�ܼ���:�$�vl[�s2}��=�.6g�:����yhV�[�s=Ȼ.-�E�
�^2����9��zW �`H��g��b�ፘ3��yAl�Bc�&ԡ��2���4�+~��J�����q(I�������c	Q����o�"f�%��Ͱ�hXE���p: �{m�����z��@JB�c]�}#��� �K4�Mi	��o�K�޻�W�25Ù)m�-�;Qҵf�����K�r&MEc�& �M���+�B�q������_2c�&��z��ew�s�E��ȷ"(�]�Ua#�H�h��E��(?瞢��Se�%��b�}�a޶/R�"�SX�a�ʩ�Jk�h@���������{��N#���N�zVA�(�q���~D"���{��l�� g��ib�1���V���r�v¦g#����@)��-s��HŨ<�t"v���,�TNAMy�O�P)�iuK:.~��}�;ŀT�.�PF��r4؈��~��&�J����
�n%�(��bW�{!� ��t��{3peo��]�D!��C?Y`C�Q�� �@�d�aٝ�M.z�/�'7m�	[_��~�\�3� m.l�!�O����*�x��?�2����^�[������ʠO����k[���]=x��dtŸ��Xc�m���t���F���I%����{k�<B�b~y��a'@����c�[M����@��E��Tm.�cW��MV���n��7�On^lwc/�"s2[���ڭm,"������xM�޼������8!��eϯ]�S�pb���r��e\:@y�7A=z�wI:�քp���T�wv!��g�(1������d4���5aw(�P���7hqř�{�c� ��r�5�#��N�*��|��b�c3Cy���W�B�rH5ڂN��N��.z�+R6��Z��P.XGǑ%ߌT�цFUl}t���et�LQ��_�2��܎�o9�\=�{f�)Փ�a�T�/�ά�pGK�B�aņ��s�kb�}�q�5������0n��.V���� 7�v1AÕ5aI�u��	�3׀=�G|F���Qv��j�7�Qe� ��qbS�}�$9	�D~ظ���C������`��*�3��L�F}5F<a�Y]$~#߿t�l�\��HQ?��$1:����,��!�[�Q �v��Dߤ�R$�ֻ���� L5�s^z�>=�����A�~A��9V�{?�rE��t��0$��}�l_�Y�>搕�6[�����3�.�Nq����Wٜ��H��*��"ZyĵU�I]U�@��Lo��{��n�]�xrg+�0�>��OQ���&�?P�%.��۾|��k`<XQʿ����8t��z�FB�>��y�.�ܲ؃�,�"��)�Y9��Oh��#s�j��-�x�<�{m;����u+I����8��z��ڻ�$�.w����k��K�_^�׭�b��
s�٦������>��Z}�J�Ӹ_Co~�A����˖�M�Z�Z0�#�,�Ո�nuQٍ�Ze>՟' ����O��ч�uH%�n��@�2�,����A�gA���:�kG���>���
�Z��|�e-�+����ch��[�`D�љ�]�q�Ɠ������j��y����^K��u3��S��=�჈c�FŐa��J�'w'�
���j�h�'5�l`6�̢��/�u|Cؘ0��̑cd����VX�'��.(����տ`?|�ʥZ�(wfkM������c ̓��@����\��v�=9�H�C�DB�`�9��q���:�*ՙ�������U\������z#�щ,�A�\�;�ޯ���o���LV)������m4#�:e��H����Q�x����j�/c�#k�k�1 �h%��~i"�Z������nRfқx�}�
������m>.�l�I5�?��Ù� (=TVq'�(�
���
v��a�h�|�u�x5��＆�%��jtM=��s8��Q{�S]�n�OP���Ńp��G}��ON1�K��c����O�1�wW@�U��,�#�|k��z�-Z��T���7���g�:\G%%��B�=����F��WDzNK�Ȃ�b����zi���&�qx1����}�'|�S�N�k@D���� 	n4��\f�v������6��������D�B(��0�'��x?ȝ��v�w����&Zw�.�&��cٚ�d�߅gRo�̙��;�wɚ��x��py�<�/d�9�0�V�J���K]�y#���ޣֵn�|,Q-%�_����'��*v�^�v+O(�.)�	����r����l��;YR���*GwsDa2^�`M�6�R��L>{ Z(�����F��9�|u�0�m#p	q׷��?:���hܼ��bo���~���q�%���%<��J��j^]��qfTҖ9�V�8c���۳!¡B����t0��v;"0�Q+ٴ'��.{�Ak�ؗ"-:�.�4��J�:m��`��*�`�����
T��lF!'E�i�DM�ig1�T�4�T^b&�}�����l!vG3i���,�ui�= ,�L�1� ��߉�ZI�Ql��܇��&�Z�:F�.	��.��rᾝ�z�+�V�-���ݛy��^w&�>��j��_��u�e��6G,��2��������by�8��r�VN���-�zE�%~�p�>xҗ��뺌J��	~4i�V�&z��i �Z� �5q.���K��ͪuL] e7��B7�`���_�D��R��4~�+�#N8������r�݄M��ZM��v��1���Mkq���ݒ"�����x��οΜeH&�P9��g�j����,vas�/����/0XܡaWU15�K����M�C�p-�����G�X�����>G��wW6����%���[���n��=tr��h^� F�fT�۷?�F�P�Y=b�j��2:�&�<ow9a&�O@D��|��ګ�٥D�s�pF�s�I�*)a���T�'�?Ŭc���^����i��eK�l��䠼�H�����o�@g�7R�pn0LRʝ��K_p�B�:؁���O-��/��J`bAo�
�P��B��	eF�;4��ӵ�C���GH���=�1�V'��G��b���츘	�]FG�"��pxCQ(/W�?@�Jt��e��)P��np�,Dqys��a�.^��뛓וb��S~~Lr��ʀJ��V�*�v􋰪�� u��[ ������ĶD�j�d©Cw�K��Yn5-��&���� +|���pu~��o>~)7�����Owu,{��<;r�d����%����I�[��s��:���
�6w#�(�>�K������b�+:����5�H����ͪ��a�>�	�mAH��� �ʿ(󱥔�q�b;�ڴ=8��c/�UaN��asMJW�3�Q2�곅�,��饠�-�!V�����{jW�>˂z��G�9�jY�Yx�>Q@�}�@(�wp��W%-��,�?:�C�b�\ۑ/MP��by����U8ۦ�|����*��Wrb�����ֿV�s�<���*�8=q��*A�Pmu9�Yڢ����7��P�l��~����W��~���}��x��P�C-�_�� �2����C�<`� @�ja��7�Ǭ��9H��9K'�J�#l��^G�YG����S�R���^��+��6�����,��8�-[쎢Y,!ǉ���IX���V��TG7�v@�q��3�=gY��(�1�u��<�{��Ńe�Ҝ�a�/v��
��]A~�k��M�
��h�5�v�<�Y]G1��a�Qֳ�0�O�q��Տd�UT�3�>`V��#Y̸�K�Up]鱦��� ���"��6f���+z^U� �M���s��̹�D����{��9v���>�r��<�MZhf܍:^l�ݒ:ص���^^ݼ#6�M-��7E��9���sL�LM��M��8<!|
J �����n|tlF˱#;�eI��ka��.}�hw�O�2!y�Ԛݫمjy*lh�=<���������ڝ��#`s���mi�L
k��[�46,v?6O1�Ξ���b:B����c'f�=�m�N.Ր�C�����W�Z+�6-�DB�#�s J��z������y��U���ݣ4q.GD��Tgc6�]Mִ��q�-�`Md}�����U��6�fol����fA��΃x4ګ�(y�6���k6N� ���y[vg �D�_D��,0ۣ�3�"��,B�
�c����p�G|~,�+�j^����W��G�Y���8=Vo@�~'1і��w[�@-���ǘ��z��\������j����[�q�d��Z�u9��L9��yj�W��l�0EZ�� 偘lUɨ��*��E$�Y(j�B4�����X �B�K�ӏ�V��'��19����<�{j�\!�vWa�d�S�l�}���W1a�G�Dk.�;qS8`�W�vnDV"�?~�}��q[��ݬ��k�LI�����CCa�xG?a^��y�����SMR垾L3���ms�'��-皔-'ӻ�Ш�iAx������-U�BR�U�V���~ӓ�Gy���v[�1Fl���)G�H\e&`�@�1+�w�l|������x#����I��u_�����҃1���� 1S��Xղ-D���ٜn�q����FxX��ĝ��hd�Z".fέ���$��흲��y't�ނ����{d^�R�a��� ��Q����I���(x|�ܿ
�U/o\�G�6Y�n6.���S��	��UK{�茛�d'x�O�ۘG�9�G����c�*�;���es��u�-*���6S�����b�f�9��������
8v}s���w�7\W���eH5��dV�o ��*��7
R�f,����0�`�d�0���-hBVU��@��Z`Ql��9�y!�لK&m��S-I���k惯$L��������3�텅����o�!�>M�l��3�]h}�e�u�n#�_L���y8���y#ivZd(���A���Z<�4��U�����Vu�
}�!��g�$������r�M��Fx���W�����T-׫+�!K��w��i@"�pp�O��|k�G���	�)F�5Bu�1�8F\ja�1�J��ES��[��hF̅J٦��xj���	��[ܖ	U�m���Ɛ�Y��M�Jgԧ��[�+=���E���38���
X���
^c�d&���A��u�V��[P�z�X=�f�m��\*`����BF0@�;���@O�&�̏3feG�0��d?���,��xy�q�/uI��ԩ,��3b0���\��HD�/*"S�X�r�J��]&�&�Qq��9�{%�7��ځ�c�(�xp���y�7�4�:~����<@� ���e�M7y��'9G6�<�=���9����:[E'Y��ɚ?��4��e7�7,�������������^M�4�{m9��]K7
��D���)S�ՈnĈ�wE4�d��G��{O��n���#�H2���jN#��#���x�hSV�ݧW7����q���2���ī%�����f�+���g8��l�����N��^g�7>� �n�q��mA��)�?�R5CK�j��Q���S�����v=-��nH�4����e�V;ύو�7�%�"�m9�\���8؊G)Z!��0Yk���_7Z�*,�vs��H�N�] �)�D�j�Ao���e�����=R�� ˬ��ǄM��+�4ۑ�6uUI�t�c�S3�V��ͮ�8GVHހVn�n��Eˬ��L��|�h�,�c�5�rWG�����$�!�i-�����k�Ğ��[h����NS��c|a1<#z�)pn�v�Ү�|6w���x�8\^9�L(7Ĺ�MT�"��QwJ�b0wWU/L5Ap�}�����a(\�0���\�?��0���Qә��q���̖h�� h��_��և�mn]2���9�r�YJ��5�Z}�bk�� �̐��PT貐ME9��3 �L���>�[��2�]N�w�IdŬUu^�e9�L"�Y2�Z�[GB�<üY�.O�X�$����a9t�l�j{b����w���E{Ϯ���/M��X��F
�z���̄���a�[r��>�o�I����'|k�vI��bS�R>,���;������/���'�ȦWG>��5�����:�ԐS��@�UĮ�Dy���·X����y�!F%x���,s8��}���x��W8M3�hpt�Z���Lt:}����-�D���
@>g+i���{�&0FƄ8d�>x��zC�m).��n�/o�S����>Y��CJ
���"�΃)B���~�ub�vS� b+�p���SR�0|��#�~���������dG5ݢ}}3b�.�4��4�@�|��N��e�Ddp��`�����3e��=�V�  ��pu������������5yq�Ԝ������#m/�#�XG�n;ꙬD��F��e�M2	����zC�ܡ%��_`;�i�Ѱ���u}f��9�c��%�7�p.��
�0~��	�9�?T�P�%���^vY�k>>�_A�Tu	��_oRǤ��ƞ9t-.p!�x����2��+`�_��CLuȨ��6�u��)�"���4��GԲk���%l�ΡN��� 4�A�-D��?ʟ�#šEy#,}
��VW3���1�f ��ܹ	�ڎ��WC~���~��_�zv%��/NN�f�ZؘEb�̾��]j����� ]"~��]V͇��@�y�.vRvf�eQo��W�F��J�j�����t���E0���$ey�d�$��j�::���3q`qK�V��8����"�j�&?ƮtL�Z�#����ɷ2���xTX����<^=��V�m|>� O�T�=_�!a�)��FZ^�aG��I�SF�Q?�TI[� V,�yu��k���VB����S����@��09�
Ϡ�K$�qp~�jF�o�Ab8�c�iBr��}����D�;i2�u0�8�4L�b��ٷ�*j�:�R�|6ޤT�R?��aB/ N�a�cU�>Ƣ�G�B?8n^�g�
=ӋB�w����8[�tI��Y�B�nA��� 9U�4��?�ѯ�8#���v�)b�FE�h�L���a@���k�Cw�&NsMw:A��]X�`>Y����i�X��P�����n���˿ަ��t���<u�[I]�'�w��^���)��Ȟ�=�kA����a:�� �呃�| ��~I����g��q�����&C�l�܁(�c��P����.��?D�v��Vj�:��T#�a��#�ؿ�'��ƋBX�'���	�lK,�7L����lǃ��-�#*�S8]�i�(s���s�A7K�]�9�������"�����D7�wJ9��
?�Jy�O-���2x���o���P�ˈ�ž}M�M�ۻ�Ͳ�l��/R�4��Q̶:��!����P"M�c!�-g�q@�A��f}���,��#T]M����<�����^�wK'�P��A
}���O^o{Dt%�)�s�L�v��&�
i�j�WQq�����ӎ�=>Qr��W��U�U9�)O��=%7�]I.mC�~��H_���
����}5Zb%�iq5�8:��	T����ax�3]"-�L�յ/��2vs�z�{"2hw��6q����B	���H��:�^Sr-B�e�9E��d��{U����?����P��F(%hEy�nE�I(��K;�:2@�mgh���B�p�H��w��o=����o��j.��W[��e�O[�D;�'K���!�2�s_��o\�3�nvo�Z݇��4�{���c��:�g[��=�����&�����њ^���^#Z�)� hI\�;fd�
�E�{b8�өK�`e��I��-��̢"��՟0��i~�����UI�<�.ꑵ�ewI�i21�s,GFљb� ^�%?�P�=09�2���B&5���+��C���(�v��L��4���HIk�?�Z��<
��K0�ac�Y����V�(��ۗ�� �U��QF�LSp>�t盶א�-�m�-��f��&��FHK���r�C|���"����|H���*��=��4�t�`؃=����t�>�1��3��EWf��N`<䈾7�������~]~��͋M��gka�*�	�����v�n�c{�f-ב�8Ғ/.\��i�=eH��ǷX���S���,V��Q��5K�����׼c�b���})P:_��w	����z�qܧ�axx��>�g�r�1�$cU�0+�u��$�hT�S�JE�!��OU�K�l�*�%C���gΊ��I�f�I8�(gr�y ϝ�Q����o�g�FsW���r<���C}���tt��B�X�+rv�KQx�ˆ����n�ٚ�}�:�֎���x8*��\���n_g֟7]�ߝ���B�D�r��H5Qd�^҇�����:A�o�dť��C+���K�{Ĉ��&[��H��kD4��jg0�Ҕg���~T����-N�|	Up�TlyM��[�1!���ϒ��/V���`�s�T���r��uJ�i&Xko�x��j,�?��K�To@��^����k��3�L�a� �C�Ni�c��d=+�r�=�������[K�z��:*ߟi ���v7�!r,e6P&�Γ��75�RN������j��7D�K�)խ�a�>"�!0Š�B�3&9�c�>������;���bMh�HΧu�H�$�>A2��o�����c�q���*���%�������Ϟ�_��KŨx?�m g��%�}큀~;��sL�r^dT��j�6C�@3���;v�' b�?Y�����GC��'F"Ȟ6v�`�n1X�4ˏ�7��X7��10��\�!Tʤ8�&L:	�,�_�,fl��W=�\�JF滠0(f���% 1��$2f����!�\_]�f�#�)�۷O۠Cp_��Y���ʕ�YR�:Rm��+��>�� ��ѫJ�!�[��xq�}�w:1��*�Z��IkҦ�����{gݺ^9s(j?���@ԋ|�H���J�".P=G��QE�*�p���ܥ����s]�Je�\7d�.�|��|��@�*���7m`�y��xy������P�7��n���̚x���J�>��[���,�{���R�R�Br��Rolj�x~���b;�g��J�Ȟ�[2m�!� �423��`f��ɳ���W3]��L_q�v��F�PM�W�WS�p$X��٧ʳV{��!S��rqN��!I�yӀ0qh�2�B�=H�WhJ�2�9Jk�ٯ�0$"�I��WbB�(I�:�/�θ��4�D�AAh�E����!���[h�\�si��q\Iq?��Y;at�!���ɟ��7��Q��D�6ХbNb>��
��i�+a}a.(�C}��߬^%�K�����RAr���2��2o8�ۃ`�kա�q��H@$��qQum� <.z;vV�� ����da�PW8�mIך�Ch��ǝ�ޤ���2j��V���+5���}��o/�d��8[�"�C���7�W	�1��U�w�8�9���!�<�p|�?�痚�4�� K�J�����؝4��7��hS������l�ja���+K��"���p�^C,F|�ܯJ��>29�	F�����@����$%�.�'1Cp�)��\x㰴���$P�0�Rw��|��S'V�d}���e�w��Z�b���h�v�%Ne+��)1���.�Q�E�}{D�%����*De>�<�}8�f�\4}�l!_�59�H1H���ԤtQ��F��^����M=�8�D�40���Q�ZH4OS9��H��G��:%�>)�'�?���J�6:����p�>��|��BG�Rx��<�������0�4��q��Wy2�綈��\ڌ[��#����m��!H���˓EmZ��I_x�m���޴��]ng��A������u��i_̍Z~z��䚔���<x\Qd�𡓁1�(�i5�lp�wtn˓e��(F��fVHCN��I��;�%�a�kW�#������aل`;���G��):F��U�z|�B]h��C�w m+�(`c�j��qzw�KÉ,���"/PU���}�l|�tY<0!-�UV�[˗�EaA���mFRT7��\s�_�\�:�i���쿌�6
�ee�r=��{5�h��ADV���2�½�;�\A�G6V��O{��8�c0���W	�2����1aXf oW�V�1���l�򫤐�6+��~���p/ڦ\o>���c/N�`5.Y���$����Ǔ1� ��Sx���D��/�ǂ`{z�T�����G�4?pY��^��8��-X�(�>�K�1��A�5!�x0�:gR���Jt��2%�H��̆��k"M,H�R�������G��e*�����) ^Q�{)�CK�����=a��S`�4nXjp���)e��1]W9l�h� �y����D-�@��Pv�īǑ��(=-3���a=4rٚ�0��>J��!�75���{�{=s ɫ7!�f�U^������(Yp�}`n4]`&��(þU�����T���ͬQR�2#F�I���1���+�/\�j	��T�����Ɏē�c)B��=�}�~�	��o�<ϗ�F��e��ϓ��Q��so I�h��+�Du����,���4�F�3R���.	v��tN�D&<�=���ER�q���Z�\Y51�r��9]n��<��b0!��KR���ZT��KV�;�LF#�|��Y
�G�;�5r�ѡD�A�p<�<
�R�^w�F(!;iBH=-l9R��KH%r��.Z�sǫdQT��OgE��Ms&,7�F#�r��v;z�|$��<�
I��n�M�_nu#�!�~Z�K��Q��4����9�W�3P�R&�?�l��X�"/�ޙ�h������:>���	�R�&�w�о*[*[)��yG�لq�a�wQ��Ϲv�� ��S/�b�}~e}���Lo- �8	a��*�j@Vۅ�!����%5������12C>�K�H�\���0��&:C�_�y����=�S���Y��
Q��Y�7�@+y�P*��ŉ=��|a�#f�M)sj��ܽ6�k�U��x{c�	�g�Ԝ��B�\�2��v��*�,��G�u�>�J~m�l�G��܋��!�ͥb��a����Z�5�^�!.F��>y1hj[f�l	H���U��3�<�]���BA6,����<�g^�=M�m�J)�B��.)���qb�o�s�&h�hc+|�T��T��#�#]s.3FC��3�bWi��@6Ɉ���Ɩ͗Y�t���hN�| s�J�إ|>�]��F�s�$�\���XM{����,��Bl�m+ʛt�����Y(D�	���H�]`L���8FV�N�qYϢ��-"Ch��+��E0:YR&�]��;�����7�iV �|p�5Z^%�uv1
J}���D�]���L�Xu�?y����W�����E���G���{8evH�Z�=�)�6&��2����NU�ə��;{8�����}#A��怀P*��:"a�hܱ�}�[c��ɗ��W�G,��Hyz�|L�"P�-/f6=��X����nځ�"���)dޥ+F>�ɿ'�D1{�ב�ĝM]ṭf]�
�8]�=2P(\�b�}a<.�qY.^w��S�F�ͽ����� �̮�ܖ�Z��c|���\�r�r���ݽ>���b@�a�����e���^�;1E��v��\��\ :�T��=�m��[�F�P���GW����_>u�8�{�#
a�I��y��Y:���\>MXk�e��{������(�������_�����z���:G�  8�k��<�/�	jxk�-~ςܤw��9�PPL1��e�p�DY�ݐ��`�8�{�A�֋�t6�5���X1��Ѹ�j\���Ux�;�^�r�s��.�G��ZKb�V�ǝ�Y{���Q.B��3��z��	P�d_ȃ����K��,�U?��*,D���]�V��&E����q���}a��9.F�)	:�ֵ���,����#��O 	l/�Kŉ��y�SuF���3v��e(X������Rģ��B��0}*�SQ��Q	-�Agg��f�S��?}|�ob�,������^�:�Z|Ӧ7�	��Tkf3���B+���g�M�3�贘Z��s���ӗ��LdF�#3��tߗ��K_�3��8�e\Xg[��׉�ޞ5��͙���J��x�^�Y���ǠX���"�>?v1*�����Ov�AF�n^� 
�U��tXae⽎K� �6H;�n����$��v?{�o��{���(���[�Fx��_���L��"rp�#7��+>[V=S����g��m��T�;U@_2Br�p�z��?v����Ge�@��ꚋ
���`�$S��S[�j�������k��5I(�NW��/�'�}���}h8C�9�n��8� ?��B���3�*�\��n�K�H^B�m���*���]�݄�K�ײ^�C�kDНu�$�����Qx!;��$u�0�)4��[��V�n0��Q�~ς�B�:�� �S���v��������<�ʘcB#���/QV_�<.�h�M&p�������v�_��q:e��h�'n�����WuQ�;G���)�/=�6���GN�?�ִ7?����l���>�� �j2D}b&��*��Wr�ۍ���P�*�
�{J�^ce��H�C�+�QܯP�=zw�~Y�o���X��Z($ڕ�՛����CĖ�H�����<~����[*�ݮ�������n��ũ�3�]��x���������h0m0�5�|�^u��q
�q���</��Լ�����J-�m�D����S4î�8��E$*�Hc!~�u�H�[�qQ(�������`��G����X���*N��G��	��p@��n�:�2��q���s^��Hρ�C�G�/�Z޸S&HF$�+���hf��Ӥ�8H���0�̅l����6hQ�h�#�`wZ�N*Q	����h ���:�e
ڱ�1[�6��"����%Q$|
O+7�)u~�	�Q�&�0r�%,�T��2��$�m�2�?�#��	�cs�����P~����ݫ��rGu�I��K*TH�I~e[n�CI���;CAa����X�ǫx�Y��j&wԲ���,�F�݀~$����.ڜ+7dh﮲.�XMl��� ���0�X^}V�wlr]�ن��i�y@j�+n�p�+ؠ��*���V�h℥��$s+�҇-��+��F(�7��Wb���kߐǑ����k�28���4�����d^�QT�0��J����T����������F%�Ɠ��3#�e��$��<�ü�mѧp��+�#F�Rw2�s\���H�F��z���|4ܷ_M��薵POdm�0��O~^T��9��uV���VA����Z�.�c�R��H<�St+�}|#�
0 �rP\���b�(��Ғ3]� ��ӕ1bu(�o�Ci��|�kٯ4���h��u|>y�!c��i�)Rȿ��z쭊�)l5�8��p4o�_�f ���6�=����MĐ��Q�
�a�!Д�P7��Ƌ��2f9���ȶ���z�{&��]�Ǘ1-����Ӹթo���:;U:�Pa�'dfNa0��Ȣ~�wۭ�R��G8�&c����������� ����{wPr
���-�pO�p�>C�^F�*����a�2}�X@t,���(k�Ŭ�Y�œ����Dr�i�G���S���s��b���]2O���� 2��t̓�zg[�C�W ]?Ɏ��=��K~���i�7�-7a Ȋ�������1�cm'��k�b���|�R�63Q�z�C�;��{����r�<̛�xql&�+≿=`�ʂ�o�O`>Q�	J�����m���P��{:�&�Y*�F����}7�U�{�}��t!tQȰu�%!�ϑ�햃L�A�Ԅ�u��W���_��m�����]*2n�A���ښ�>g�JMġ������U>�U������&�qZ1Vz�%|�c2����' �M<J�$���S�Ǧ[�g�D�04ҁ��>�h��iD�.�k1��0澋[�c����<��y6���a7�[�.�K�N��c�q����i����M.���ufq.���8F���#�P�j���� 2NgB� v+����i���]bmNF�	��R�HG�xa�v�V�DpNQ�$��M_2a�F7��9�����Tr���
X9kT���r���D�����C��[�W�-��dI���ˤ	~��E�-���`�W�uĪ-T]���f)V��[�R�)R߷fE��T�1����W�1��.�	e<E�00u|�3a�S�������]`ĥת6�\n�.}��V^��Ο��?BGD��zAd�2�$Z������ JH��]�9��T��$R<\�0����������3�e@��|�	��j:��:n2u����,�I�^��>֗W1��(xX8w�T��nBW^����ݭ�,�Q��Yr����>{qX-�8�`H���k|��Fl�C)��[5�)W�+r�s �KS����D��h� a�[��d6�r; #�Ң�C��e8ޕIhމ� ֊�*;<��&��py���/��w�p�ã��BB�tz��]@��lX�����RƮ	�E+����6�?�.7���p�:��gF�YV��VMx�p��f,0���7�%�'-=�E�/�ѡ`���MJ�a�.�L�e��Y�2j���O��B_:�-��D;C��3�/��/3 �%�29:�uݼm�[v����=��A�ֹ0�k �>��,�Wr]"6;�9��W���q��Lcw���C�~�E���БB��w6�%����
f��H�t�;:�:�~� �����F��?�,eh�*t+h�z�t�kߥ�h��渹�u9�>�p	%�:���f�Y)��������K�<M���ts��!�#x	�K��q2kR��θe��C0�.�P.�&���X̰��62(�@��I�f�m�B��;�!�x�ZO=v� �P�Gk�:���q8�f����u�
Q�e8��dd���(���B��7v$�[�`6� Ͽ�T�\ Y$��r!�$����4�!湕,�c��U@y���Չ����c�P겾���p^�쮁\��s/K��\�����Sᙟf$�v���o/��%��}�z$�5giZ��F�c�P)������U*�c5��K������z�AQM���8��16�b�+��V0&����0�<�gsl���w#v�N�%�, ������8/��h\��hq[�WԱy�y��ʃ��i��eS�Hd���ӽ̀`;���`�w��P܄���Xh$������0���Eؿ�si���C����+��;b�?�ű?�#Ӯ����o^���a�!����= Jb�XW(�!&�\��;�*c��0?QV�?HP���2���K;���bG�MoR�d�Je)�/x�Rs��6�С*K� R$bд�e�h��ΩY�!J�Z�b��T��q��MTJ��<S��J�f�'������7��Z���"xB	]0���S�@��C�
�I������1��k$��8>o	!�ޘ,�ёW,߻��"QV��E�K�SЕ����я�j�2C,��lP֔'q�\�*\}��`����7��ԾH+��2��␋���[|�:;&D�_��1U{�"�zl�0>.�iM��%"��t�T 'd��b�܍I���������U�'v�={�X�" 3̼k.�}ߙ�1}�N�B�۔���gƷ�AG̜�?�mŮ5Ee�P��KG��0�/�VgNt���pc���za1GT��E�.���K��+e���:�����0�����F[�uT�[_�?6��mKBL������T���8F�	\��x���6D�=���)��� �"����Vk������	�
Ȁ\d`Γ��#��G��n�E�>�K�,b�v>�f��b}g�Q"&�y�����V�W��o�̾qZ5*�����@q�;+���w"J������,Waq<Olφ�43��_y���9���.��Ԡ��� �\�ʋ-H��T��G]��*��E�χQ� ��t�z ��`�/� ����H�ܽ��)�'�h�%�g�N\�"G�6��v���M�����BE��f,K(M���ؾƳ$'g�xȵ:��#���AlCxTyzƹ_u7�(XVS#� �\Z��!�T�E̲��kZ> E��޴�+XT(��� �,��� �ٟ��f�L+���F�N��L�7�*�yxB�$\�Ge�-��N�����&�q,�?C-���`�,]���}�&ў�vH�R��f�f��A��)
�9+w��������r���ܪc�C��Q9r�Kޒ��В	j��J�22���Ҕ��AT΃I�m���e�K�Nb�� mWD&�s������J�Rd!^G˧���B&� ��B̹R����R�@II�$�cֲ��5���pl��R���u�N�yѲ�C��^~�3�fAs�M-^ԉ�n N�W�Ҹ�_r�T�Ҷm�y:p/ᆯ�(�:�gΙ[b܋���v�K��췴ч�]���;��֭y��DV��Ոy��8�P�|��G3��E�ϸ�O��2q.[2���Dq��Y�>%̩�*��a��Pw���H:�| F$(�V~5l�e���������F�g�mIإP\����kFO^v9⺄���k,:�f]�MEDn�|�����+�~�n6�ߵQ�b^&U�Qu<g\3\0�e�+�=��+��}n>S���.�B��Wl�oȸ��h�UZ࿓E��>8�fR10� ��=�\�i���幤��у�W�~�V�^+����k��bM�֭̤ܽ���%��A4�+ �h�>r��+�=�v��H��������+3�\)V�
��Chq�X��g=�1��e�p,������i��q��%f_%��l��d�����������9�*��v� ���~��?`>6��� �Q��@��ލ �[iH_���Mr���׸e�Ñ�ܾ��X��iz[�].��1�?ڢ�T��%�.Vq)@T�Ai�U�W�*'�=�F�f�G�[
��"ڤ��[����a?���K���!��Ч�t��h R؏<$�����k���~����CF߯�QCϷ�e�f�����n;y�ɚ����9~�"Ú'ށA�Q7.~���N��k�~`S_<>�ѡxD^�X*�n[�M�L��m�wY\�5�rM�^HQ�nDm8�����S(j�E0遟=�mZ�=���r�(��X2���	�A?���H&�	����G=�#<��hQ,Uo��ss<�i��&	����p?<^T�X/-�-�b|���&H@dt$����l2���bH�F�2�/R���;h�]7	�^���gnɴJ�v����vL9L�(��7ݟ;�����;&�kC��a�C��	J%�0I�QS�y�Ȣ�<~E|��ī�����;�F�EtL\���$�MK�a(���>>�T׸q�4 |r���dR1@�\���~����a?� �ߎ9�O[R�7\�/���$7��>��`��=7y]�Vn\�~�S����q�����L�ĞN	H:vG&��������ID��1n�A���6܆(�eI��U���z(M�V����c��0�s8�W
�������r4�
em{���yR����n'��o�VO�1wqk��MZ,5'���s���O���*W]	O����!�&�ѓ�e��O�E�w	Łf���ph��b�Cyia��b�C�1�?���0e�i�c)�~M<��1ǉ�1'[���?�L��3|�je��P�xB��N��wUV�}�m�c�����V6�ˌ�R&n�~���찄�Z�\K�S��>z4��O�OE�s�Ba�0X�O�B�{4�]u��k �*\�Fu,�.{���k��{�xu#}D#�U(������G��=r��\�v�uw�-DܩCB.[��\*�<�"�0�k���������9C<x�@�!��fN��Pq����Zlwk�ڽA�J0�1�� R�n�+=�s� vpy^`ҷ�:}�}�*ϰ���	�+I�v׺s#�+Dq����J���[�L.����];`�e�����6.m�����B�:V�[���	D t���~$ߩ�4{_g_7E�g�>����0o�"�9����M!������1�_���r��s��c60yrA.rk�~�&��j\���M�ň�:�L�{P�x*�L�;5�NeZ�d��P�(������A�_k��l�|�v3I5	G+��D��N�S�k��<����
_�(���H���䷵�7���L�O�'
�h)��_vqiF�wK�
���7{�<%8lP� \�;�}���"�n��"3�\�9h;=�9��ҋM8h%��A0H����&�e01�etN�sXY�0QBx������F����*�>+Kj��>,��ʹ�ᕆ��m�ء��{vm�����>�Xf��m@�CMo]�d�JT7o�0�w�q������O��R�]���K�%����>����@���iZZ�z��%)��;�-f醧���^ ��S&��o�<V3�</�s�U>�f�䌛Z=��/���<���[\���t�aLb�uZ�|Jͫ��J��J������>�l����>�X�w�lO���牰����ĥԦ�-�kOR��ߢ��R����S�W`;wXە�`�u9�;c�����A�pI�
7Uu��3 5wb�j�|i�~l�'2&	g��EU�E�������C$���b��&5���e�8W��qĎ�B�"ӷW�U�W�r
�`�Ҷ��d����ϫ�I�7�W��sH6��P�_Ϥ
@�z�&`j!ܠҲ:ot��r���A�7��j���֤ �i+[1�6,��U\F
��#���B�^3f���^z����u�ă� �Xދ� }�m��
^ (���Z�ަ�!M��5DΦ4T���-@��5���{����͋c�����*��I{�r";���(v~�`\
�}���-.��'������\���ߣ1�@$GW.��eYA%XmU0,�S6�/d�?.N��C~ٯ~SV�1���`s���~z�t�4P<<�0�UJ����) 6���U}�[�PkK��F���'*����i�&���X[���b�*�фN���&��e��5=喁V�u�/��Bs����O�zR�+�����A�T@�e�b�ڌ%8��L�Ⱦ�~:�J~�1Aq���4I���V}]G�V a�p�
MV�ţq8X5Z~ǶT.��a�"���!�c���x��ċ�VԜFHݒ�f����\y���͑�@����;m�D��O u�2P�^��X/���.�7�%���ES�1���g�lr��{K�u���
����h�̲{}��o�a}�J�0�A�=��ч)g8�L�廊K��"�e� �����J�\��N�����ϵ��޽W�P@�T�o���Z��tu6r�nM��,�Lr
<����j� �|`Q�z��t��k�Ұ9�\(#��:�}�t sj�іmAxz����`�k�m)<b�N{ �֝_�t)��Ք,�a���6���?�y��|���L1�ΈU}���yƄ����/-N��'��-��d ���\���_��{�	�;��Mr�>����aؖ��)��dJ�ehm�+�ĥ�PW`�k;E�T�/;$�KŠ�[o 0
yw�Sz�fb,� ^�4��{���W�^X�,�Dx�!�מ7����ھĂ(�p�Ԯ��d�6{31O��T�Z2՛/�vE��h�=��,�<9g.�����k#��3�Z��K
C��;2����������3��f���/���\y��v�L���>1:�4M@)#�������7���`�d\�U�`�{x��/��4�^�&�Z��7H_�؀H;��u�� ����c��De��vH_�dvdڠQB��@�lEm�y����L!2���Mj�3�A�������B��}�~i^�����,�9�p/2�Z�.��Ф�
 ��q�:��(.��̏���R��lF-*�t��^�Y#2A���q��,�(��ٽz�5��ExWs������> �;��%�_��������rb�p錂�c�><��Z��a�7�+�p<��ф�q/=*�t
Mǭa��������zV��f����7K��C�=C�m�\f��/m嬬�_�.����������_���}�Ϡõ ���
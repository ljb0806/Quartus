��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y']��=�%��]i�5��	-{3=��y�ר!�<��(�!�(AR��W-�$ff�P�7��I�8��z�4�iox�[�Xh9%R��KI����Dy��uz�0�m��d���e�|:Q�i�T���%@��:���J�=~t|u����G�J�jp�Y&�S�4�C�p�}��Y�%��K�pe��*e}V�\����<�^ǄW��r5cL0:�Ki-��g�*|p�B4g��3K�l��P��]��V~|�h�:�9\�RV��PH*��[��-��$��2�@�H��r�/|&6.�$p�����cR"��������d�+�ҺK�*��hT�����xΎ�O��u涠�8�f�$��S]k>�8���$Q����P&����y`"n���BhY"{�A�/	� >�f}bl6�ڂ�Ш���3�FH�U&;z9>�i��r� 7��߷�y�FM۾PAPj��&�X8D���x��*�� ��Gy2��0h0;��M�wjA[$;�`�z��yJ��R����/_��p�;�v�G�j�W34D��1&	�S?�l����tը�tUZ[|{{p�G����(�snSC��ܔF���w"�saO���dF��딣�r�cV�3�]�j�~�n���i]�N1Ae�M��@%���0U�Q���/[���2p3ڙBnM*��>j9b��h}�zM�Q澻t�tc�����?�f�`�z�N�����y�5cB�O8�P��F'���ز8��zz�ʍW�Q-VwdQ�q��Y|�!�dǗ(M3���$��r+�V�Ҳ�F�K��p��	�=3c�")w^+]����*_�Hv����3M3� �B�����_ن�Ņ;!/Ͼ ��Y�������i��T��i��Ⱥ7T�ف}�G�g�U�ꥬ}]�6�����n��o� / �+���jQ�!�����>)�2�y��^r�-s�9v��9������Ix��7��ܥu&�F��F����:]}�&��}@�zŕ��м����'U9��߰��N��F}Ճ�F�ө�7b��(j�j���;4p� ��tb:v.$�/������N��"y�(Y9���@=�����CAh���u�;����ؑ��-�i!ٖ��� y*���fY�9{vm�2�O�G3��3hH��q�t��d�l�or�ۖ)��%��Bu�Z J�y���3�������\�Jp5؅�����>���濈q�/#�����t]ly�5�|���:��`��% ȹ��2P��OG�?�;�(��d���[��%&�Ī���i�n'��²zKfm���S�|V�4g�Zf�(0�0��*�eEE5�E��ƁD#2Q����'��=J-��x��2� ���R�	4��'�1�4e@T�:���I��ꪝ�[��#�����o~F�ȳ�" fv�Po!ut%p��-�WL��tɯ:�oc1�����*�>-x.�@H��£X����׈#.jT����e0�z+ �%�+8��[Yp��	Ȕ^+�wÌ�4��苐��@󼔂8Ǿ�3�=��^�m0G^p�C�d����Wxٛ���t�U���<&2��"bzK`џ$ʫGٞK���%2�y�#�Mh��`��Kw��с!A�M�_gj7���L� ��ĵs�c����1s��p8��ύq�;ec؞�]q�^X�@C�6�(G�/B7�o@�mE"J��Bׁa�[�#P@굁U��>���r9}Y���pb]��\r�[<�4���yl-u�<���hn���0���%���pUǉ^4>3O]��{�;P����l��=&z����\�U�VJ��B��q���;���-$f2ؔg2�u����֛ܴJ���t�� D%���7���H�$�'N��?Js��*&�Gz�]A\��O]�@˺��94��O䠝�3�7dԂ�����_�>�/X:����Yx�8˓>����PP�T��)|n�q��y;m:���
C�?��y*'��\#�)�$���.̲�\�Գ�\"4�%�k�+ܚ2b�=�<�low�VB拣:r[d�#��� W���cY�{�F#�n�xd�=���.�8!�����<��a�P�rh��M���� G��!L��61f(5�k�6(�;�#�~�V8�ҡV��ʳC�pʙ�$Y��о��,����I�:k���i��Z2z�������w��Lʦgl�����L,V,��q}��8L�њQ�2mm���]���z#m�> �nB�G$Z>{�e�'~h�">���i�cAE T��ꗼ�4vNh
f�ز(YП��Д�ML%$k��Z�#�����C�1!
/	~�tI;(9r/lOfZ�Ďy��_��΂�rA+��b�a��յ.���X)Ҡ�G�p�Ƈ�S����1�i������Fu����΃��m���VZľmk��%����`Y�e�MG��-I�$�*fF����9��Uٛ�LG>K��4O�A���P��<U2���Ȕ�$�5���:(Kƫ�a�i�EQ{��z�׉�]&
+�*S5IL���)���mV��2��P�',d��)0�I�H� &�Wn&���G�a�KmE�*�r��D���������W ��(��;��	��z\�I��|��t|!�$�����
�.� �\��3�Jd�8�=0L���J�"�PT+��ɐ�LD� 4Dx���k���I�;5G�k��;�/�EVQ�.v{��ih����?<����}�d�$Ё�ա�V�l�F�z�y������P��s ~v1*h�cM��Xd[43�>�Y[�4��ؾ�7m�>����&#.�W�a7��J$��'�?k�������s)[Q�>��>p4�G��2'o�s��N�牀�Y�p�n��>�P0W'��w�����Mx��Fi�'el�ࡻ��E�I~_ߡ7�n\�Q#^�;�p[@�F��n�$�s�@�G����y�d��qYy��t�圗~q����+bd�4��K�-7������\���no�hX���w+~nؚ��9gx�!DieQ��$W�/`�(a���?�n�f���MJ��	���"��� �A��?�=/F΢��ص�ZM�S�;e��#� �Q׋�y�A�F"G8�g�T)x�����ks7�;�ސԎM�o#�Zg��h��w��tCr��c����Osа=��<�N���1m��拿����ZY}�	ʲ�R��/��h%� t�#��ca��b#��ft�A\��Q�
ڮnK�q'1$��Q&�r��{kD�#GP����*�*�VHE)�!�ִ8Ie��Ҋ�=^~�`ƅ�G���~���gRh?�T���ǀLM1��z�B��S�vf�0.�7�z3���ι��|��>B��G�z�d��2��+	�q�"XF�,㦦����y���q�ؙ�VRJy�X�����Ѝ$�y�+2J����� �x���5,���<08�����k���5�.�>_sE6����� CVߡ�H�^�]׋���՜b4L��
r�w��&ֹ~�]��Ipip���-p�9�*pW����=h�x�U�U
�|Q�@!�s��t/� ���t�&��R�y�P�Q��șS��	�A��V���2�&�#���m9R��.]�R�D��_6l�~& ���*��1��W(y����n]��qq2qҞ ��h�0U�}�&;��.�,�ʹ�R-s(Z# 3�P����@3a�q]p���Z k��"�I3�.�C7��7P¡� eX��4�W;�IhL��7�m����:�P���.����Ks����.w�X�F���C"�|c�} s�t=�A!�$�v��Jҕ��^�tx�K�HT㶷7�[h���O��8}�\�X���N�os,�+���M��]�E���1��1���@ب�Q��udK����ɢ�Nͤ7�H3 ���i�<Fￅ��-Y�3I��=o�x�^�Y^l�5�7|��A�v�+/zVp�I�o|H�J�u��wؗ˂�-?�>6��<[܎����E$���#��e��g���qa+�e֬��%}�T��`Э(=;>�:^0�0�\���qT�b��*T�(�1�%�W��������R��g��G[L���8���V� �������ܙ�3&�:;�&60�2�g���������o
�[�L7��VpT�.�3��V�t)��d�RD����꿵�,0��+	H�}����!���x���!a��1�M�t`��0d"5�H7����l��a���/z�����<��`�s.<ة���:&G���Fe1�n������!�j8�=��md�ȧh�'����짫�<%�y1G�K&R�]���.Wm�i��$�"6���E���.VQ��-t�kk@QX>B�ַ�(���*\����,:��qL��_���L\��K�UǞ�0<A2a��p�FB��9�9������oG���� �p:ߜ�f��Uϼ� S���8�,�.��dQ�W	7��TDc��%�(=�q-��G�����֬��uv'����2S5kiǁ1n�^I%�vO�XWa�cU���2
�~�o��-2-e�J�	e)�Z��Ց��`CQ���6�^V���e�D����P�F��h�$!l�}��h�X ��LCȴ��B$6F[�U�P`�
�!��A��.I��n�w�{ܧ�%�g�\5�a�-{���X*p��^)Nѵ�R�J�������֩t�~�$�Ġ�N�*�{Z��Aą�P�C��$�#�
�7:��t�(ҫ�!�7�l�"�~�N�-���FI)L�l�lq�
vJrA��>�)�Z��:���b���v�N�B-�$��(Jׁ����jH<"v���`�:�T�#a3�F��,��z������j��S���3�r��b�8`D��
U.�+��cp�ev������ �aT?���vߙ%!8Z�
�E�t�@���N�oMc5��k�B���Թ�|�e}�9l��I��������F�F!CHbt<��l���,�J�4��8�񗉙�w��$���l��O��x����̏Bvuj֩�ډ�'<՜��Z���!�s�މ�����9V?r�ΰ����Yw
7�u�z�T�)���L�`�d�JCL��y��N>�'6�椇�G��@�/�DC11PA�'&�EL�ϗ�{l��M�\ ��"<���9�p���b�f�ꮻ�X@k�������*w���?
�Z/�ϴ0Ǣ==jq�������z&��uFv��{�\ e$����/o��i��	4T{DWo��=�Ec����M0::��ت�fYp�Qk�	��5v��~�M5V�5��9=a�����F�Ј������ٷ��:�O`���ҍ�+�g8��dI�Wɤ��e�����N��R��m�����KoVp0�S�[y�.�S�f@*١���\�jf��͑qDՊ��9k"�F������G�_�u0C9�A|HO(|����B*Ƕ:�!um����b�����x�����u49CpKn(�2EX���
D�q�=���Gr,0Նg��K���r$�Sv1�U�خ�C�A�x�|8���9E��)֙�t}M	��U��	I�R���������팒]���Dp9��D_��C��큣�'���-5�ɼ�^�� D�>�6D>I�
ZPA{�Յ��K `+14~��'�7�<�6�M��z�U@��eϲcN�]���+R�S���l�� �ܬ�����j��=hEIl�v,�r�qWA�E��g%_�1���ja��fs��[��([`�D��v� ʕq'������uA��Y�C�u�&��@�.���EUՅ)ȚIf�O��,�7Wo/�g��s��m��tu�8-�=�V��:�Q��}��?~�%��s6�Xi�C+�@֊�}�������m�K��Bepڶ|o�8�+/��fx��hh>mD�T+xŝMB!y�i���:�=��l����ՠ�4����t0!n��"��^0�k[���`�VG��#��WFHGe�M?}'L�`�w�RQY�_�3K��ˮ醞W�){8d˃N��־%�K�Ghy�/lJ'�a�{Qd2i�'�<�����������f�Kf�V ���8��q8�g��颖g;�\���}�|:b����z�{�'_���US��f�j�$�K�BSvP����6D쫕��c�1��/����N��|�*E�����-��EhS#�3��?�N+��:J��3�q����	�m�(��p6�>���7��;*�XҤ	�h�,o��_r9i�O�j��B|��1�:��g����Y���5kp���x:%`Q�����mc�c��{�\Sj(E�X�HV�%߬h�t{�]��n}	i��Dx���^PU@���=/�vw��7�o��7��k4]R��R����9ѫ͌�6�Uf#>���=?/�;��$�j��V'Y��ҟ�
���B̒Pܸt`�xFuN�1�X��Y��������*���o<�ap��D�)�����@bl��v�B���_�/�f�*��R�v��!+z���B�e񕝚N"Gf� �Rʔ����'<���Y�e?��"�VSޤ���T���s�5i������#�6�_�"�-ڍFF7H6W�4�0�=�FFf\�2 y�����d-��8*U/��#x�'ҫ�egY���OѝP[�ؾ��Pw������"�Bl~^�p���a-�П 둟�5�/e���
Դ �����!Iq��C���!2�H�2���;%�b�C��|5�����:!p�4��+��y��Ʌ/��vLJ�������^�IG�:}�f�O�b���P��d�[oh74�9�M@���F������SōР�զp�u�覙C�ҭJ}�_
�R�0�Q0�����N<��ye�]#&����8�gsn͡l�+����o�>e���q�n? #\'Q��B��&`���1��r��&�?��KY�`M�Я��1g�v+li�$D���������9���a/�~`R�I�z� 5������3����v�n�:e�X�V-�XI���';�(>ڵA�r��gJ�G-ㆵ�=�>��K{S����Z�a���1d�ؖV>�����$F�#B�)-���M
���GG)u���Bc��_�9$x�ؑ�����h�7�ߞ�?1 Ȓ�$�F-S,_��1�� �A!�4ژ�v1x�!�.��!ZM9K�q�}�p&�צ�=��VAC߲cU��	F�v$YyN\5-<P!ݸ���j��O5�3�&�c��1!�%
G`�.iK)$܈\�2`#�.���V�8�.GEC1L�T�<�RSֈFY��hk}���w����V�(�:����_�,M9����9]6��R�L���_� �2_q�u0�&@F�PN��)�$�o�i�sZlb�iݗ�]�V������[,����p&u�'D,�>��L�˝�A%��_�Ǭ��	-[q���#W����">һ�����1�Ł-c�'�|亹����FduY#��4���wY�b)�Y�J�ȴ�C�l�h̼ؗ��N�]?ҭoqtv0\��2�B�ad�CĻw�8ykR�ۈ���7�ĈP�|&�J���W�|(��J���M�1X�=��2��&��
�� WHڝM�+�����'��y픯.��1D��\�db�G�� o ?�'-l�y{�b��R�t�N5����\���S59^H��	��P{��}�N f$*�\jw!���:�Փ⳪vk)/h���}{EW�:��� ��j	<��^P;[Đ(���Y����� �� pAu��@�(>@����=�؃4N�P1�D6�]��Z/���+��.�z�����r`�u�����]��s�0����r�BOi�+!���>t�H�u�R�d*����O�����X���Umj=tΑ�lU���Y��!�[Ee6�����Zǈ2���w�8Jn��Յ�� 荅xբ%
��|S�Ѷ=�pSĖh��U�9�=?�������/�������d�O�(��$�~��d�tZ�ٱ�y�q�~qiW�E4:9�FB�2Z��,rz���a��m>2Ү@���w"H��3-�:o]1�Qa�>6(2���뇁���%�x�@+�z�������=��v�ğ�@��
e&�5E�j���ciZ��u�!��b>�qEC�m�
"��{���]�:i(�L�gvq��������u�mm��1�?�c��HH�7QHw  )4	yl�lvg �.�jIƇՊ�O��e��gY��v���� f̧���i�'s8o��⾗u��2�9B����^-�޺�=���D�۵�'�emr|��}�t�jfOK>u�@b�a}�Fmq��ہ�������-�D��윗������x��>y�,�O=Z��):;]�9�UQ����,�41Y 8n����,���v8��[]|��-����g�����~����,��o`��I}�c=��W�:7礼ԆɐҾ�Y�!�m�l�r��V���x��TLn���FI���c�0)��u����+�lh�����<]�xp��0<m7���{IT�\�8��E�Z���k��Q�w����墍�zhN����R���/vn��9�,�W��'�W���W�6�\B&�Q���(Y �Ѯtf��|Ɯ`��9}NI ݮ[M=R�Wڀ��3
�|���l������׉�@)[{�W.47�}F��[s��~b�k�Nᅮ0!|31�S���}�Vs�,�q! .�������O�[���<��sy2acj����EEȘ�Oꨀ�2��>[2�c�MO}�sE��mL"��H��/��H��uU�)���
���;��7�SŝDQK���7�uYB�s��VL����fxH��Q�J�F^@���	B�����%ϥK��l�[��eOI
�|�d�q�����Cg��F���Uuxު)]MQX��E�0V�� �쟲#h�)����&�v������3�{�wݦI�g���}�n����R�G�EZUT�IF�-�<U��ܻ�J\.�-�m���}5:�d��^����|�ف�
��/<�px�5���G��/��̱<� ���t�U%^�Do@��j�d}�7��@HYH�ܵ�64VQ�4��bK�K*-�w��ﱻ��E��\�R�{.�q����;H[�ġ��d�G��˕�E�R�7��:�$55%7�.�5�Nɲ����9a�kxP��r�p� ��-�P_�D���o@�����V��T��o6�И���s�7[��#r��Ty���4�YW��AN�U�{,�^�I&kT��1���*���������>�̋��L����3L��g�_h��RD��Q�M�w����t@YV;�ae�޳��*�玘�|b����E���0>���ӱc����9 H���1& ��j�Js'���������״Mj��#�(}��~xBL�Jካ_$�
IVɼ"T�8�vّXP!�f�(�8	p%��a���1C+�řW��SE����#�K�=��p4e�]����S�~�i@%��|��^.��bg���)f>�}�1���r�*�U&O,GvF��,�Q���]'a��;حި�[����*�d�d60n�+(���������T��G=�2��~<N���(R��ڮj�7��m�c{>��}H�9�ZF���\1b��k��F�#P�Ӷ�JwI(�)����_���X��䉏��5(�������O3UG6i�f-��,�꯴,���*�;�}rD����HL\ Ϧ`!���b�� F�R�҈P��H����`@@�\����c�7�t(��˼��n�_�=Ql4�*r��$���@�q�����Ŕ
S0?M\}�|�\������#�o_�h���Q"����_,t�����Ah�ٶ��7��H!g������ݟa� ����X���m"�eI@�kØ
fl�f=��B鋽�������c���B���y|�S�r�p�\�P��]������<p�Nr�����)lt���$}Vxf�ϸ6�-�\Ň��$�m��[����tFS�ݨ���?�R�%k�k�Fe����/Ǧl��5��O�m(����͍��Ŗ���j���>��EQ�p�w'�ؑ�ڣ۫|y���7�1�=IwY-��`��7R�S0Λ�ʖ�j��K�a�s����?��l!%f�t*��h1������OK����`����v�n9�mVm�=������г���7>)S_��5�4`[�x�F����uG��Ǒ��{��(�E�TB�k������B��[�3�B�����0��Dd5W�8dv!)_�Q�!���,���;�S��n1�/}A�K�������qZ)M�-4�v�Ѵ�Gb&8���B��d�D��Y~dnP������ו�Ǌ�wo�;�R$Ʃ`0��W@s����%KڛC�0��B*|4=+�а��?i���3�MO����_�/,�v�t��N"NL��E���	
t�m/���`XN6�~�1^�����I��4����~(�-D��+tJ~+�m�CD}��eQ�E�Q�V,��:JWx��C.S����M�)V?�v&��!�ɱ�0٥*���g�_R�#�<�����J�����T*�� ��q3+~{Rn����4)����W�c�!�ı� 1ݿ��Y�j��p��+&w]�L���ۊ(:E*��DM�b;Y�!b�	�C)o�Z<�d��i��`�:��?j~:�TbCc�Q�3^Sr����(p���gf�	+ "G�i�E�=͢-��0��t�	,��iۃs�
W�IU�僋ً�xVC�0팚�1k�`A�@�N� ���k7�Lߙ-��vG:n����e���C��byd�bI@�tD}��|?�,^c���D���E#��?�w׮Ov�Bhp^<x�(w|8a��b��*�n����M�h������s4���a�0�IZ�,-����'��us��߄���6��`�9�q	T�T4c�^���X��lK`m<�������u[7.m�H�h����8vk�
�\ݓ�����>�e�ҹ%q�Vt*,��u}=BG7��ƃ_D�T*'�y�T{Ί[̅�7�y:�?�,ut�	�iŽh��3Ӊ��J�tZLH�rh�_\�8�6�%XX��s�~��k��a�Iыf�{��(@�?{���fm�ݬ�m�\�͚�q3����F+@�y���;�����y�3�XΥ<FL-"#��bh���7�+�Ӥ����AbJzi@Z�+I1�M����Y'�)7�1�&��&ܯ{���.p�l��#e&�:�Lcp��-��0Yp�y6p5����0Ѿ9!#��[���y$*�pʍ���è�W߸@�<V�H��8��o��,q]�J��H�����e����H�/]0K��-m72�t�hIAD"�^�8fI"׃U�������u�p����@�f�ZO&�fe>���k%���EDK&��@�w59*�<�6㿰�rPF�)oτm��c99��BN��`$���q�"NYC1C'�>�^�@���m���Z��]HS�V�-�y�wٿ!êja`'eĀ�z�BBy��O:�ͻ.�;n� �A-ӎ�H��������e����>*�AL���b�o�'��}��Tx�뎻<k{Ve6�=q���N���7��&w`���[�v!�a�}�yC�����e�Jwa������}�V�:���A��w�W]j�7/<X�Ov҇{:)h+Q�K�ˑ�ߝl����`!RP����M��U3��p߀�\ᒮ^L��7,�
5u�G�WҀz���dis�*�������'�8�UNFU�����1����Z@ɭ�^�Tݚ�ra3�����Ѽ��ou	��t�8,�Q��L��γ�3R5���[���%z��z�G�#;P&�hWu�5>��0�;�Eqth0/����Hf��Ƨg��
��BWM"���bk��0�W��m�t3J{��ZG����G'`p���T����
�:��������b��U�������t5ݝ�R���ytKa˿S|r��V>╳Z���>�H����=����e������enX����]5��3r}]�f60{�!3�fszp�b~��纵�������y�kb��{�Pb5~q~v[�}��qM��0�`F\q`���6���z��*�C��d9�F#$�x<NߠP�7��pq�Sx��Nw���tg(ja�a,��U�M<��Q��R���@x}.]a��~ݕ��z��w�0��@���~�R|���&ģ����ر����,O�T���]I�3��fnKY��:�Uɗ��t�+[�Zd�6�7?�0���M�r����t$;�01�I�L���|t���Y��lU�8eAG�~�v�g_�����1�;��5B(�rE��/�0	���������z��.B��-��?�VR��`����NE���J^وh��;&4�CC
7n�L���%v3^�[�"�ׇ]�r�\��U	o���������
�TL�N���+u�1M�b?P'ٶ˅܌���r�ۉ,W��<h�={��a��e֛��[�hA}��d�,����cg?����UjAN~8;x�Yn�2K�_��ce�
W�D���y������ov?��r�Zwp�#�Q��$1g~_����1K�[��a���|��ax���ckvrQp��{]_/��᷹�/�\�.խ�aA7����,�+��W����B�b�� G.��^p����mB�L�T�4��ڿ�gU�	�MxD���ç�淎3Mh��.����N�>~�z)Q�V�D��~zme�~��2����ዉp7�����lZD���ܬ���}h�X�؇� jp� y�NǞ��7Q�5G!�D�FgH��W��ܻ:=���`텥C�:"�- ���Dt!��I2Ӯ�%�s��<ei�a�=�	��ٮ��n�Í�J�����a�q
�+
gYX���s�K�pc"�5˕�O��C��C������#:H��˕B^����Ɯ�q���a�����4k��݈�#�y�ΕjR(7)�T��b�"o�������O����W�}�
 /T��})��(\�Q!B�޻�/8�*ُ<��.kE-����G*�F���\en�ѮY�m��~�̝���~�sy^��Ɇວ+ b/Y��n�=�A����Qf H�4�2�:c���ת)��BQ��.VJ�8;����.�~�^�EF�@����P~0�(�e,�(�Ǵ�!8�(v��B�,�p��a��ְ�z��b�"xQ��(�8:�6�D��#s���YML'��9$��rvo�o�V	B��m�i�5E���y��"r���`wS���H�Z��r �}�����q ��� ^/h`G�]�NN�#��'�FaB����i�䇿�2��a�q����=Ŋ��	�,yW;����G��������)1o�n_��4�f֡Y�8��f{����!f�*0�s�&o�z v�5�Bڃ8|/�K�X��"�(=�@_v#��wq*k�N�����!�QV���)V��N���8X�Ҹ���?+g������� @T�	����1;pq�m�h��
9���%ǆ�C�i4�y��|�Q?i5#�P���_�_�s���:(r�<O���T��� ���HK�K4������%u��UGO���}LTّ2�k��&�H�$9��Ǿ�JĐ޼s>��#�ko&w�#�,'������Yg�!%�и~�5�'�J�$�Ӈ��sM�r���`ap3-��Zt?sF,���b#%*�f§���n��DC��j	��$���$Ά��akB�۔����
��|7glJ0��m1�nQ�:���|��+$�v�����v�CC�\�.6�M=�}�x�>�?ZGv�,<�'p ��o�_�����UI����x���rVCb��G�
���(lK|���F1���B
���d��Μ�J�K���4c�������9_>�~	SQo��)�C��52.����W�ˢ�
��@��^��S�ܮ�=i����|a�CϮ����']L "��4^^S����$X�z?��n���͊G��FJq��oVq�v1 �� ��*�&^T���$� `5@�����bɇ�<���2��z��Yk��ߩ�`0�W$J�ιnI� O&3d�¾I�vg��\0��[V�*1��\[Rl�\�04�u���(����)���s�����鼊��%��b��&M�bvċ̒�$�¤UBr���Y��׎؜���ѓ��EU�:�ne' !����iP�����1�0��C��h��@������$.�#{
\FqG�);�Nn55�������Mc�k�#�2*b���6o���+�v�?�e6l���\�sl=�4e��AueRMպ�'_�89�����L���&/Z��%�M�����y6�����>���(�"�&���Tdt��3����}A@Cx}� �X4O�uY�zOwl����,��O��2O�7m"��"�x�ǐ�g��w�����~�Su���F�?o�G�E��Lb���l�_-�t�"���SX�Z0��N����5�#��7��j�L���TO`KF�7����ˈ�Rt���ZU��6)!�
ήc�t�7�*�i����Q)���޲��Z3#k�HF[B{@B�w8����/��p�誉��^���r��h1������%*�8��k3�!����^&�
ML�યk������,?��9�u�7Y9�nT��s�e�0��^DIk�2k�7l���=ou�Ɔ�*,.M�d�1�A+ѐ�K�!�.O����n"�%c��������\�qK��jV("c�;��k��A��θ�胠���:�V��,�ج,KG�u�kj�MG�3U ��DL2�q��|t%w}H�}	@���.�!�������H(�,Q�WV����z�߬/f�]�=���#2P9�UݸAr��n�\�?�!qN,z�8�b����4$��X쏭����CX�^L�.d�NB{'&;,,ڮ{Dȑ����wK>Қ����F��{c2Bq�ă�Į�5Ћ�N��D}�qX!�̋��X��f�������k��H���u�e���N���1���+:�q=Ιi��Ԡ�}K|ՖrX{��)p�	����Ҹҽ���tYm��򻭀�H/�0 ���Ro� $0��o�Uw	��t��`�r�l�ݍ���r�qb�����4\xY�e�wْ��� d%�Xb�K�9�Qe��67Ny��ڇ`��ʂ#G95��2�G:'U�rЂ(B6�Db��S�!��8�!��F����	��o�51F->%�x�W%~ױ����:�cix�?>�:
`��@�a
btv�>�����`�Qz��3�n"QQ ��d�=jCe��b����|\�NP�k7�MUʭ�(q�H�<a.���~&��e�e�B�=R�)�R���/L �ʞ�O\Qpdд"]�\�K������׫���`2�@�dI�����?��b�מ���a�_�&G��
%Κojv��I�����TP/Lgqxf�k4!�]�8V7!�hSPn��J��d\լ��4�5ѡ��Gł��	�-3^~�����ƀ�\�i��v�j��;���;�zBA�}��	Nc�U��O��Y�MT"S�{c�{�����&Lc]Ue��Ԇȉ��w8���J]�c�����E���?"%�������A:���������/Y0p-W`�[O��`��U����D��� �9ԑ�b`X�X�cR��lj�!����C�->؛e9g�9�	���\~�0m�]�ͤ�a��ۑ����Zf`�z�>�p�rh� �|ڸ2�х���"�6
��FԵMwAH=z�Y��y "��V[Z̻��ʄ	�Q�p�4|�"6Kv(-(q\��G5�FCg���9�)o�߼j*Y�4`�����qj�=봂��S�Zd�tIi����^�O��<���ى���oy8�ڲ��=�8l��+8D,0T��2�s����雱��L�W�S�-�V�M)���mH�L[��y�Q�O e��IsK��{5C�'Ĳ���7��Y�>	��E��в"~ع���g��SԶ�Y,D>�:1\����3F>���|�s�.�����![X�X���WA%��S��H����;^t��1���C ʗj��2�ﻁ�;�n��|�p��:�a�)@$�+)0h�ϕ^���A��iJ�eB�{a��Q%�]ǼM����F�S�y���;�`ko�U�&0D>�<ӂx��R����E��\�]���ܚ�
�����`��K&j��h��?���7 ���o�N]�T�l�ql�"� ���e�v!�NH�P?Gq����C��+�=��x��'�r2��R�*���%�=���"6��x؟�<��lX���*F���`ׇ�
��&�Z��f��F�?�֯��+��>�$��Eq����Z9J=��Ԗ��LW���Z�]��?V�9>>v�٭�[͏���N�~��O"�θ/���ħ�.�C�:���A:j�!C	Yt��P���ɀ��W��ě2T��r7IZ�{@wvL`ћ����n�{*�'ڈ\ʵB`�*��?������J��ê��Up�!�Fr��!;P��~(z��qֺ��vRsG��Y��ζf���B�L� �Pw5p�Bߴ�(��x�?���Gϒ�R�����{UH�0]���{��{�wݛ��i�S�!o��N�b_�"B;�udX����[53kTd�3ePFg~���I�-˲p�
Y�_��d��!3��>�Xh� ��p�yM����b[<�� <AN��iQՕ��29vJq��R��L�toJ�m��Jy�N�~��>s�).Dj>I^��h{��M����;�m���s�`���e�R�Í�;�v���7�}�Z�u\Nf�,r&l�/+���,~�̎��G�%�{��0�j�r\"�b��}��u[ᎂ�x��P@��7Vc��s��i޸��Q���U���Z����^D>d���-��W�/��ȡ��#n}��{�N)�=INj☁S^]s�Z�� Mb����7@D*TT�
m�NL�O�g��1�6�|,q?���2
Ԋ#^��3��=�i��Wư��9����xqc;�c�l�*G`���s�/��N�/�]˺TJ;d#��5v��ݠQ-~�����*�s���$��!R����f�I�Iϑ"\���}�o�E\�
��T���{�u���U�0ϕV,�y�F۹R��+b�Ɋ'��F��<xh�!P{hÖ5ԉ��T�#�f�r8Q����9~XM��3�A;���(m~Hk���j�� �ܢ�Î^�
�>�{��W�{v��Z�pº���p��H������h;�;�{�r��� �hC���b[�
���cr�^�e������سy�`;��^��b�|�]��Y��ц�5�m�ЦŎ>����NǨG e^SBȷ�F�ca�`v�K�o�Ml��䅊F���8��i?��9��5�[��KD��(G�!iJ:$J�	3D�2il+mc��0.�Q���?����v��③�7�����=_��` #�d����Q��%аL�$��0�xJ���l�-�E����:?�V�������)�+�>`[��}�.�ϟ�M���0Si�)��M]6��w'� �+�k���$`+2BǮ����N�s{�����_�&փ�0Gx8�U���`�c.�o�p�
�;`[�<Y>�2��(	���fs`񽙘~xnHm
������Ek���X��5�D���6q�CX��O��+-��b�!<x����D��yV��A¼�6�p�m�K�_=ԝN�)ހ�!�C�Q���Rg�$�T0p�Ys@�|y�N�a}j�_���4���K�E�h�E$����ҴpULn�P����t��#�Ut;��տ	���<��
���ķ����pz_��S�q�3�:=ަ�w���+��&$��Ğ��L$.,�l�F0na�K�w0J*9r5��}ij�������'\�a���ŊY�-����q�=��Y�&&H�6ܶ��(��z�K)����-��+�2C%��,�������Pt�Nft�v�/Ǖ�)��3�U��wy�G�B	>�y3K�dH�XR��7�3��@.�)�eC��7H���x���j�B�-^n�'���$����N�����\^�V�.$o�!B���9z��R!�;[>��w��.'Yv��v���4&0j�n���)�Ƕ7+��]/�>��{.�v ���c��8�ɫ#gmh�:�0��l���V��� �8KyD6�W�	���П�!'�E�ǵ�<���|�+�Sn�1����:�h�S����t��n.���i�_�����D)q��e�u��1�-i`�����,M�m�^i��M=nM�ay��'��#���3�7@B�2m�2%��G���{8�W!����)�f�E�E0&��^`�?%1!g[Νiq�^�FXB>��0Q͘�����4�w��Fc����C~�)f�p� ��I���x,�B+�s�@��A�IYOn�P���&�0��� mV����i�b? �U~����2ϐP~Y� \���OŨe(���*���b�ێrÕk@,�a��_}�>v���k��6X���?:�S ��E8�E�u�<0*�Ϫ[2!,/���^�	+�J�7ʃ^�|awgi���/�
�ϼ�1��B!u2�(Dj=�k���݆�>�n��%��Cc]���#װRk<���J�}L��M��^�^q�����j�)� w�o"�#�&�ь�yB�C��vZ�t��&%/b�,N�N��3�e�5�����߆bL���G��F}~I1�'X�����_�)�� z�ֳֻ�lG���r�0�s(�o$�m|�=�f�ƽP>��)I�I=W~Q��Æ0�Y��d^��,����a�{�K�`��D ��iT�-���&/��³��%1�&����e����OB�=�2*IP?���M��ؒ\.��'U��B���fe2j�.�.�H�閆.-����I�Mf�����ة2%���E�qózHxD��җ�+�>{?��Xx�EK8n��kɤ���t���'9�P�飠ž���x�\��t0+� �F�+\�{���S���$C -��s[���M�`�h�*T��~���;�닚 igJV��ъ��j���� ��.ɉL��8()x� $L����C�|c����ℓ�~=6���E3^�h^�f<Ƹk��ϡ2ǰ?��ZK#$6!�m�����%q��O�W����L�5tu� Z�����m�s����W)^I�
8N�p�d>��F	����,v\���F�F��Eܵ�zm4�)~�a�~�;�#�sp�?Z&S�\L�c*G����`�S/���7M�əW6�pS��j!޺����q�~r�}�e���ﵿ=Q�[ā:B̩0B�b���nRߥ��Yы�(h�����6�k �|X����j���^�a�ؤ+��u�6`A��d�O�4����V=��1���<�cD�����$��Mn�x9�?[��?���XNK4�oTh?��UB^�;Z����T6�\�j��� ����h����)��w�]�:WT��r�"�}����)NO^�� y)�^�m�^t|��mW�H[�fi�b�^9� ~n�5j��]"����	��&K�Ở�ö
�^���:9�{�����)�(���� �-���&@�B*���s�Mtx����s�ل�u�eO7�h���Jl$R����e7��JR��Gڿ2�G%q��;`�^�B�>K��H�e
�3���gP��16`��hJ��6���%0x��x��Ȋ�J�'�W��n�P�K�^�X=��G�QO��r��dW���H��1�Fs]�Cq❀h���il&��Օ���`�0��e�%��=r�ɑo�;�ˮ�"0�{��:���J�ⅆ��n�ΰ/��>���_�>�EˍOl	i�ay+��t��8�6~���չJ��+�R^VL�^*���]���d���ɀ����5�'���l�1Њ����b��Z�Hv;f�D.�(Uv��˻�Ovz�bE:���v�� X4�b�sI������ţ�^�z����p�ǋf�6�xE��"�1�XG
��c�)�	��h:���֢�-���ݬ.���T݆�m�(���9C�
8`t��!'������;-h�����Z6���w��R���bl}��}�#KB'��O\u@�-�o�XY_��)�UŇ'�&
i#�����Ї�1僵fP�(��A���验.]n�{�,�uj���L6E�-�?����w%c���nb�vbx���D�,%�����AZH���0Bn�4��
R ����Ϝʆ1���b ��A��X��Ms��^^�+����K�8M����YT�E���'�=Ǩ�-"]��ձ���gM�x�	��s&@r�MAs$t�T���n�t��o�r�ż��|���T[�0}�X0-�0��Ꜯ�\u��j9Fx��j��}o�J|ij�4F���%/�i�yI�hc(�D��'qs��E�O�{�jkM��g�+o�Ҝ�΍ ���mw�V��S�x�o��6`7�cь�����+a�2�������Ih��M Ѽ$T���s��Č��X�y�h����
�u����?K 1� �cl},4�.�*��$Zs�3�y���PP�G�c?88v��X�o���^Pۥ �d,�Xj��	a"1#)�{VN����\���E���1��֤"\yXD��A�>���M�#��[W����A��e��V�X�7�M�Y��z�?떊��`O����1	F���q f��1�L%(�/�ӈJ�q�o���`dib�ˇ<apU����	�Ǌ:B�5Hv`�ikE�ʔp��Ǥ��H8��
=% �8EyP�pB�&V��F)��p/ӄ�rm*�|^��t��3�$M�=������Z��\N���7�L�j�_��NiF �?zC>H�C�A����x��?W����q���/L�_�w'�~�1F������ߪ�'�2ĕ{��I�l�:,|����S"ۓ�_��2{�3�	4�-�A���b�̰*R>�A��O����[ǤP��VC�m���@[�x�\t��P2�|	`��7�Z��T�I��@�I��g���>�m�޲OD%�u��K^�2}.���{c/i>si�9�C�,��9/�&EXq�&��j%ILu�����P�B�;r��/
EX���w�� �l���2���+Ev�Y4*�@zX�W�m���%ɵ:�c~�֜Ӹ�}�6�Ia��~����u������/�S����NT���1���z��ZG|��s�N#�<�����(Р�v��	��Z�E�"m���2r>��'�:U��Dꋅ�����z|�z�6�چq=�-���މt	c��@hD6vk�P~Q�L�3�;�;#�<�=�)�or*�RzoEе�6��v.��H���o�Z�?��NC:�NOC<Xȏx�Ό��7;g�lg��͢mB��n�x� #?v����n�^G>�
��,C4bQ:bM[��M2gH.���]�X�B�T��Q]d�<��C�>��; �Le��xY�����/"�w�ٷ���{��Ж�ģ2����ޚC���pg�P�a�W���z�����ܐ&yl{�����t	A�dlb��t�T3Y�J[�AL�m�����I��<�|�2t	�,��x�=g�� RM�,�O"x��:�t)��$���U(���s���э���#f��|�݋��P�P�sq�nPm�Bs�:^��8�x���λ*2���_-�2�fw���JD��^U�(!c�;@,� �V��6������\/:���S��oo�.ݲWұ)چb�� q�h�wk�G�W�M�
�����I��+�w���S�"=J2	�~����Kd)ܕ�)X��%~��b��Ĉ���ә(�yd;s����j�+�1R�<r�s9Od�G��a��v3a�83���m/��c�K�O��o�P�*z^�+�|�\;-I~��5�8�"�j�?D�!�8?�%ؾߑM�£xëD��+mǊ����-c��7�*�ey�{������XG�1�Qz������^ ��ŏ��������JQny��͂�g�?��/ư~�t��e��z�G�4�މ'H+�	'�����S<��SEH����{,D��8�ܽ���qk֬�p����=9ׇq�����;ʙ;�#�聲jۙ�%����L����:�Y���"�*�',�؁��⤈�ƅ��'x+C#�}2�w���Tq�0w0ў�}*��Z���U�}�H���)ʳH����a/Ş'jk��Mb��Ԃ���q!���	����~0�)�jn>)O�YM�1Ǒ3��%.��~�5me�&9K�]:P_�7����M����>P#��ge`���W^�zGV-�B�ż/+��������'ǳ��z���, �9�M�[ш�������E{35|1��s�-��]<e��Du�ϖc�0��_ =�`�Ci��x�� н�}����2_)+������/�Z<'�><�Dz�Gt!F���%�[6�?
�d@K@\x�se^ �V��cz7���U��-���:��L1�I���%0����j���&D�1d������{��<�g���fd�ٯ��^o!yT��sl��(,ɼ��E�7��S<�c����_����Om�a����p'��l@�~*(597|����8�$���k�&*$W���A۲�&?lЌNFҒ�K"��n����ڈhd2Md|h���Ir�,[׫i��i~�7�{/ ���:��R1�2��}�g��2�����׋�ZI�ц���3*q�f��Us�>(����X�'7,U��n����!��	�y&3d�6[AK ���
�]��\�?�w��J�61�{�:��������}ϊ��
m�<$Ǜ�Kl/V�����ݘ"��k1������<�E��%��[S<���Sa��DLv��f���)�c���.AӠ����G���uo�r�!�Y�ƖK���nC�d&4
�j����A,�ٗ)�K�g9�2�9����fP)9��~�a�?:��t�
T��D���5��' 7ѝca���Fu-�ͫA�����c���^>�%����� � lʏ�m��(�0��ll��mq:لz^���*�<�g�Nv5;�R���=����\�-s�u�_?G$���[l�S����� ��o� ��k�ƖES���k��9�%3�o�'&���E$�鼁�C��t���ǟу�(������z?�)P�>k�PS�O'r
���ڕ���ޘ����I41{X�T��=�&��u+ZK�IY�|���/?��$-����4g��5�"}LB�T;e?�Xs��*�&U��&0��sy�B2�t��1�*ǒ�s�+O~s�3Qĭ�N��'Hԁ�%�d�搛Imh��Й"�	���� ]r�$������Snڊ�S�
-���NjKVB�4��g;&;�*���nuM�k�#TI�#�j��H$�`&K!G�����M�����>8�'�W���vt�;+&'u�{���uՕ%�ƈFw=-3�f2t�@�+�}�G�"�G�lX��'/�P_���d�w��U�"��ed��l|��S!�꿔�Ɣ��6��Sv�찑y��s'-[��
*���Xe����\���q�B|�{*2�6����ߘ���Sv�v�-�s�M��[�_�Euq6_��e9U'EK��~���*���F���q9���hC��;���>:_ }��<Z����#\D߅kW0�٧�-Z�FT
����;"�t/�^rc��H9����dc �L�N�ě���#���(P�Buk�a�a7e�k�W�V��p�b���j���]�Mn���ьϒ���n�,ş+㘛��:�$o5�غ�V���e��M����`�a�)����,��n�lB���q �m����_�}g��[v��?O3���b#'���=�7��>���@�����o��0:�c���}<��J���]	�y��m<juR%'G���F��j�6IeڙaL��H(+��G�Z0�Yۧ��I��ƺ�A��B�/�e�]a�"����$�dZ���ا#������@�G3�t�%��[ڇl>1Y��;�J
�%<9+�$�C�e�e�,���pj�t �t��q8�,n��Y����w�ڻ��:�n�Y*����ZA���)6����V�ӨحXo�@�fpx�J�6,�l�z���7L���&!�,	"φ��%� �=o��Ct��2-I��b������؍�,"KW>s9p�� ?Ƈ��(���I��͋&�P����S�^��R�#c�9�CA-Ӻ�{B����~��|���|�ڄ
U7�1v�K�;n��&�KL��^+-]!��K&�?��[�}w�-u�cHf�P-�P-ާ�AkW�[sP2�v�����¸Xb�$V&�W�/�ko��YZ������ ��='8'¾V�ȫP\�aeJ�+cO&}��U�ZǏ���n5��K��r�*�dTHe���->�Y�Go)�rDX�؇�*��UI%�������V/�w���'��آ'�NM��H�A+/� ͞�����p�z+���ʯ��)��ee�U��<�%-�*ul�Y�@S��m&��B�'��X����$���0s싳�Mՙ�aV��[�ܳ�Q�xu�n��d�k4�PR�v@c�!��6Q�+���&)���mfWA܈�G��p7f��?6�JG-��""A�ue��Ʃ?�"�4M��^��T �Ӕ|A�P�� �R�I]��5��rJR���	��2��'�#�#�Iy$�f�{m�gtfw��0�b"�,�Aa����@hsM'K/���U`�00�#S#B�sfm �����(��yl��r��e�N�ݙ�b��ժ��S��T��ub�f���;a�7%���׊���MC~1 ���2�dZg���޻>�GHv�7#RP@ݸo7! KF��f�'�d�~�2P��i��k�$~�=�=��8폞O�ɘ�΀i�̙����Z	B'r/��m���d�?��L��䂕���Z���������=	Ѥ��0�x�ы�R����r<�D%��īF���O�$n��M�u�\K�0��Pj�c|��\8p�`��]�4`2jYL̺6�U�����Z��cI����<�-��5��7CҤ�_�;���ׯ��ف�8�}��!`�tp�����n9`�A�)`��?��}�]w-^�'�h/���E?s/Dq?��c�����Ce��kn4��(�!Ǿ=-�ϑ�wb7�_o��UR��|�^�౔M�`�������z��3����=�O��6{���	D�L�� ��nXĈRi:B���F�d
: ����z���?����Ձ�����:�'���q�ױ��YVUH#�=W���gG\K�,G�z?���^�9�U�SDr��z�vě��e��h�����C㵒������i�X��{~VG��c�5�:b�ُ�u�>k�a7�F�1�����4{�XKjں3���A�!�R�-�n��8&$�纤>p7I���s�B�Kg����:�d%R��R|:~��t�������$��|�]x}߬�~6����ֶGt�P1��ɈJg�,+L��%ݶ-;�˧�0�̧�%�E�/f��B�B��_0P,h^a�q��J�ŝ�G�~_��k?�GU��"A��M�x���F�
��������N��jU�[7u�(ְ�T%[�&���A0��)����>�ۈ�������ؽݷ�ܺ��	*�k�{>�ysذI�x��'0��[�5�&f�|d}�oju���s�b����r�0O���[��?� �Ц��`F��K|��|�)kܿ�eQ(w;S���-N�(��;��A��X��%�5P�sу,���b�SjD�����οHģ�jx�W��o
~��ڬ�8��]3e<@��f3+z�YY�%��<@�*������N�X��B��F_4N��-Ս�`-m��h)�6OL���Hٺo��)�b��©�v����GXB�7	;�DJP���0���j���7»��d)N��C���D�c]����%k�:�����ܢ\+���ohaɽr���h^����NE	^��!׻#��F��]�N$�Dt<���l����y]\�,�ER!��e����o`�i�$���޴������ӭ���DۗЮ��R9\�m�+�C$j�/�S?+bN������[��3��v�D�EjBX��L��	�ܕ�0I� ���%+NyF�=ᷫ_G�\�� `�P�>Oi�����+Wk�␡	$ӟu�-9<�*>\���)��ʚs	&�-q�?��D��`Tj���'n"���|Aۦ����2�YTo�"�hR�ݽ�e)�ʄ���T����P0��G[SE�XP�i��`������y+S�:^H��y#[yI���[1�}�6���̾@tɚ҉�Ҭ�TВ'O?q��K1�6A���`�~Tz	q��Ǭ�P��Lߨl�&���95���|���CH�X�}���h4�_�'��V�R�����BC����υ�u<'E��5p���~E�܄J�Ʃ�mk�@�G鋂��BH��$͜
~�?�!B�&�e=��w���k�oT������uvS�-�ʹ< `jWr���dG��`��K���RC9�x&t��]�%X�=�`FpS��ь�Fk' ��Y@��ɟT�a��؋��!��	�N�4���V"������j�g���@`02s�3$ 9WrX3FN�ԇ�1��N�S�~��O4K���Ғ�c��D��&aP������������%�JHޕ�~>�H���_n]�>���jמ�}U�p��[f`����q�l�:C��d5}��AF�\�Y��e�sCDpV�&@��������Yg7�P�k"ˑ��
�=s�5���A?��� ^�K|Xб�O
U��
�Y�Q0��)��Jj�'��;;��f\����]ӊwPZ�-�i�k���V��~���;�"nV+�Ml�������B��
�^�,ǮT<D��2Cj<9�EQ-����A�p�N�L\nB �+'h�)Q�T���>��d�*]��6�0A��ny������A���������l�2�M�Ж�b�x�:�b�����&�<G���v��� ��	�	�u��$�]N�Y�}e�;����W�w<�ՏMJ�kdȫ�QD9��p��I4'����Ƨ�[z������b������G(�V��U��uQh/����]|�V�2�c�i�)@*� ��m:+9�Ȉe���%���~F�]�gS���x�;�0��c���tZ����0����MTϯ�[o9c�ZP��	��@:����c/tNw�ᚈ��i����#^�{xn�E��hO��Y�/(2��e��tG]s�������[o�z��t��LF��X�/�C����K���y?现�A���CN�Үͯ���w�P������q���e�~�d��ҪT�!(y�e�4w�@h��0��Gs+�Bf�Dmps���d���˨�k�����e�KK������6R�c�4�����Q�����^��:�����u�[�,�(��Ӷ&��}�b�"�c�#4�\���EP���ѻ����R�ـ�)(�Q� � �����a֐yė��kR@O�\י�Ϋ_�HiZ�q��¹����.Ɓ0�pyj2"|�w�B�ʿ;�:�Rܛ�j�DS( ��-��N-#Gc^�m���q38(�m�%�7U�:�b׮Ku�����֖�EI�q���W+��k
��� W��"��K
n!�ϥ�9nhE�s�E(?ܑ��o��X� W�%�i,#ܽ��Kf�_�ѱ��tg�SHF����34 ��g��P�
� ->Q��ƹ$G�m��%1Bt�!��\(h�py B��J6���Mk
��h����I�p7a�!���(�)Iˑ[.F�m�00_H������W��Y3볃��)��a�% �0Y���,M�^���Q��#'�B����:N���Wca�g���JzC����8��"�i\��a;b O�

�y��?�`%�l��r��(��W�����0�]t�pc珿�Jx-�
��-1�zdj[9&����2+���ޒ+a�Vgy���
	wy7Zj?�����l+yF�ʎo.�B��S�D�$����sH�}w�|�o� >3�A���מ[)����*�[t��m��Um}�
t���߅C6�Ƽ���SPƼw��SRz���Z��l�$ԁ�zI�m��~٤���*���A�]t��)��m�J��x�L���3�S����YO�{?�x�g�>��
��,�?�T���$6��\�	���I�� 7��^�RA�����kKު�h�h����s�jm��n��/�l �|���M�z@t����c��=�]�g�N�鰼k��Q4+0^.�fzӹ�谱,�����\�(�U3�Œ�O7\�O��Pu�WB6��n_�
����>0(h>�f
��鹶�<���hl�1�O�glS�=�S[���ii$����[+�8iaޖq�U���A���R��5��po���!���LgUe��HX���.��җ���L� �/nHʪ4m`>H9B��2��`��A���%n���EJ�%�Ҩ�"���$��q���k<��l��$3������dڿ5���멭����9(\R��5Q;Z��܍@��9��Rx�Y�,��|�G�N�,A�����7ӷ� w�L��I=NŲby(�z`
��HY���������x��#�`��N�5�/�iR���i�9E������@��uF��I��^lؙ�����kb�1M����zX��۸U�3�8)c�d4?����?�L��OY�w��p���u�?��p&�5�*'��.����ި3-���;�
�P���j���>	��.X���F+2�k�;��u�c=��φ+�'*�i���^|�Cs��7o���^ИU�pPp��.��,�54���
�ho��,��v�6�y���3���3<"�@6Y�Q��������0�q����j� �Z�����AN������*�jg$��Hh��}=_�u��tDd���`�Q�<.����&}異�o�c:�����q�dR}�ԅ�±:��$K>*����Q�+�ŋ?m6�I�|�� ��?[���=T����VAk.��*'���e'���T������>8d�L"w��,�6�d��Ή,~M9�M���'��u�34�2��ht��~��v�Y�O�FJs�:�5��Z�~�Va��_�]�q�qwg����t���4�*�'���P)�R�y+�hPõ�b��u�~2z�X�b#D�_S���t	rqF��&�U1����Pτ�i�e�m�b:h�ՖD!�W�/��x�� �r�����l8��G����"Δ�p���.6G�w�f2��T������kҵƉR{����F6�o_����Q|��(om�21k��%�4^���{ I��y��1�H�P��:�
�K���AN�O��:�k�P���~'�.u�GF&�<��`�>M1�����V�#�Dӥ����Z�8u��O4L��{�b:���a7�v�#P���Q��'zB�-Y��O�o�X����z-�'!�ś4x���@bIb�RT9��b��?S�[y���/��5,�]����t-�i��/u�g�4E�DPdqi�s�����g���E��d�ek��e��=�M>|�8Ր�1H��<��@k�g�"F�5����R�v�k�2Qy�κ]�����E�)>Y��c���P��)�z��C�B���(k��Lb�=S������_h����I҅��0�8[��o�Ov'*��lUy�z��f�6�tf�3�8������ϑ[֤&2S�2n��e��Ϊ'6���t㝾�'�P}�J�f�`F�� t�]�G-���fZ k�c^��4p~~�ޱC��p�W��z���6H8Q�M_�I���<��CO�|S9��{ר�T���s��E|]W�/b�H�8��;��Cl�FN�^�g��i`l��gܒִ|�%�����8�����r����ڙ#��l��g�8�S��
nئ;�M���l�֞;*٬s�	��pr/"dL��}Vz���H� ��|i���J\N4�N����.Sפ8?8gc$�Ėޡ�$�U�s&C�4�_�{8���ZK�a9`{3x�20e��lO�_����\}�5hr|t=G ���_�6;�6��b��b.�����j�Pǀx,���پ�/���-��F��!�F���4l�&oF|3�\9T��}�W�
�-��X�p��vL�i��i.l�6nP�nw�*���$h`z��=��\]�l&�"{
�;��H�ZB
��OW��ⶼ>���5a��v7����Da�qן��^6�E/��E���7t�<�\A%����[3l�UB)a���,p��U���(���s���JD_mu�d���-�]��*�,)����F�I/d�p�F�mI���Wv��y��G<�j�$��XRI8�Ѵ��NN�(o�M��x�%U~�TL������A�,���uM�E�n�.�]w���p�1�a��5x�;C�eR� �If-�郍GC�I�i8�߆��֬l�=��{(  �qh;k�w����w^Sò�-���m9B��%��͓�2�o�|?�G�����p�N-�7�-3�����'|y�b�~1uCG-pP����H��~_��%��L�EΗp���9�(�+X�4?�L��6��bQL1��>Ս>6��%^h�^���'�>n�N�V���n�o�P����}�Q�A^�)�RUJ�@w�hr�:#�hfi��O����V�H�{���۳M�ׅ����eW�8x��D�i�:���R�-�h<���a���	�`��Q��r��5�\f#/���0^I�� Rt�۹�3y % �~Q��K^�V�RJn�����i����+?G�AK9��G{ݥ���h�|fKl��{����22ϭ�𓤑���7n;��%�a���-#C�m�����m���b?�!ۖ�^�|��C�4v{�i�&�;ʠ,S�1��G�?x6]I�^-��*���RmӪ��x�#�upw�2���ޘ�<۟�PDY������8�YnS�r��j���g���gx�N��Ԑ�Fi�^=�^mB^IF�1��ؖ�<F��	+������FM8�@�wW�,�o�W;�f�(h�t���cW�8��Vw�,Sk�6��\��|���Ǻ�/�|�q�%�C�jӘ\� �>�{A4��"��7k@֡e����/Q�	�>u����%��2�k��#0���05�����L�][�iE��9s���U�Y7`T��q��*�XH�5^��j�
|ݣE�cn��W�/k$ͻU[X)�KiN-e�x��dbs2v��u�]�/�u���pbv�Q�h��� Ö.>Y�O�|ƾc$����e�F��:��=���kQH��̻��0�y�uD+�r{��~�֧"�3#������ۦ��SIڻF
`���_V��jF���5^j�Y�\�b����L�w~G��7
�����n��Z�����2Dv���2�X��w�����k�7G'^&�y4߮�.F(�7��$
V����ٳ����]j���1H�ʍ��vua��U8�#�ŰO.�UI������?���e��ວߜ\n�U@�����HB��D�0���='U�D.E)q/��/�B������sL�-��,�'�
@ٜ�;���M�6"�܈�6d��תv��`R�_��/��+OIay�,����c~W���X*<&ɧr6������
V����: y��ۏ�a,m:��n�^�A��$M�=���	Mt=R��M����U$6� �Gu�kF�rB���T�Z�	o��B��c��*X$���;J	R��K�#���mр2��Ѫ�¾�ʻ��jhu�����籓������	0��r
�~RB���e2??�C�p�ۮ���O���Z\m@�[�ӏ��ϻ�8Jo�gD�G��^��<
�Oc�5ǻ> 6G.{�Ô�t^�uSz�|���O~H�5.��`a[
�Es�x�Ѝ;�NQA'�o��4��ߑz�B\W�����
n'�@2���L(�Eh-DqQ���p:~������~�kP�ػ���o������5��Q�w�;T`���P'��j����{@�d
�8��Q￸y��2Zj����+�3���
�#e��ց��l��!���at8���K *�j�}�d?X���D���Ug��}.���/pӌ����h�5]�Uv�����/6�	�.�����4lA�{>M�bW��x�6g��]��OQEZ�\@r0J�a��h,�*�s�%e(
�wE�T �VM���K��;�t�}������j0/v,Mm:�9�Y�U�?$�RXh?"\/\�5�	&L,Vi��[�x̛0ԑqD�����O4�D�(�_),����y>��bU�QL/}��<����zHV=X�>������<WJg�;4�_����mvA�Ʌ�__�a7�J��[ci���ƐO��i񛂹��x�P~�V]ܕ0�Y��=�Ѵ���3���j'�����P�� ٰc]Z�Bj���Ab�[z\k��G�9��c]��*��p|�2��(���(�C���EE!u<�p;�xэC�>������hJ�t:�V1t�u���1����al�Ej'�ԧ�	�ɳˠG��/�!�U<m�]��GH�nGu�	6Pۣ[�cx\-$�)ی��Cb �p���@��F��o��Չe�?���;�^��hqT��
E��N,��=dR6>���J�w�b,1kqc�9�`SU����	��5�Zٓ���0N�_�1���*'�"���b ���RqR?�����%�9+�"�]�V(t��(U��푴�g:M�5�}&ΏZ��{�"��T�^���N_�PE�ű!̆Z�d�����ie�*���Gc���n^�he_%�a�������������C�[�ZX����V5V�j�І�S�.�������c�F�"B�իf@���J^�XxN3ƹ+%��������ľ��Ao.݉XJh,
�����#�yIJ �Nǿ��7�
t̠I���v�@����Zif�P�^Z��ͣ��):6�A�E�"Ԏ�ҝ��7��ǵ.*��+םߜ)��;s�]��%��M�.����Z�M��Ɓ_�i% ?<��=<�����;qy��U�k�N��n�%V�D�8i2!���~߹V�Ɩ ���Ƣ�
�[�N�&�nKi8\"P�_f����ZP��lM��ʀ�]�����0 �y|2�!�(�x���qP�&�r	��kƲ�"�YZ�?U9�.��i��z����Kٟn`�"�e�L��P���g���6��_�qMxZJ����h��15B����?[�=P/��i|T�a�>3���P���Z�F�z�>HP����\�|����LD�*��H������O,v���+7�'�#��/U�Bq<��-��1�AQ�|�200����e�;�}3ݦ�9Դ�gSP��4��
�]9t:���~�SF˦�#��6-�i6z��$D�)�ȱ?�tkHl��p�%���Ӯ3k�ۦJ͂��L��N�%�];dþ8/+������g���.�[��?{sR��K��=M+;�:.,�� l���p���I	:7�ߢ�4�~�Ho���r R��0l���Af��Ⱦ%��y�LH���Ͷ�ۢ��`�:�3��f9v̧l���xk�bT���U���}�I��� %��=����cv���u�V9I>�X�Np���4�hh�����NѬ�J&�f�Z0|W�d��d�TS��g�Ɍ�s�'&�ӱ�>9n�$�͏;�6��˼�b�B\ʔ�Ϗ,%���a�F>7[`�B�`�Q��TG7�|��9>XG�k4��mG5�����K��G"�h��6��؟(Zx��m!F(4
L~΀�R����˳��x��q�a?��.Î*
��9����e B/�5E9��]�K�aYO<��ʫ08�::ae�ˠ���4�o�=a�0����a�m_=7�ؖ��2��%$ʳ����8���lCH]�	L��b��Ţ�MNǑF�,{�Rk׺��/������E���[��<爑�b��_5��R*~nU�U_OrKK4{`��W2�Sb�������/f7��`�/+k�3zvR�*�wt9]�"ɲ�ˆ�#��źr��/{"!��dwT��=t4#r�y��h�p�!������U��2:°c�& P���Q������?Bu
���U�IXn/N�,�˪�k�P��/��V�R�|Ê1]-S���[�/d�e~�ٮ��uJg�U
����R�9�0��c�央'k)���7�k'|�^p׋w��t$�zd��W�Ъ?@w����9$G�Y.�� �䗪7�)��8�OYe���mXr�����'щK�euP��j�H�w��W�z�/��xs�� �w�L~d�~�0�O*+>U����q��O���t%+v$*'P1�^�T/�"�Q��s�S�$��Բ�Nm�J�}���E�Ō)+�o%��3X�;�HPfa>�#9�g�=�oֻJ3�f�!p\i�$��6؇�\ 4��X��糹����z@w��-��A9?��g�������3���`�IfD}�z���f���Se<&,|�=/a��꼯�3'�ҀDӵ�a�8�-2`q��1��n.�v	7�FO1��a��~姨���}IS2�fS<��_�bd��ݓn��W�B�?�������E�X�FL
�0sh��6���*��;Z�j?���Kq��`�\��v"��v�2�r����3ET�q;��m�A{T���  j[�=��È*s��Ph�f�S�f�g����+g_<홈0��ļI49 ���E�2�a���SQ��LJ�4��n��Gy�#�I�E!uK�F}�7��X;,��,���� �a'ͩ���=��Xx�Pˏ��@fBӳcu�K��#x&�]�k��s����Àe�A���\��q����e�q��Dob��' F���e��U��"��`
÷�{��/�L�E���Ō�2�o&���Z�����8�>�}�p���	�v>�S����5�C�m���3��7��ܿ��-]HI�
���ڟ
�j�Iܐ!@��G����r<�w��`<Z,�0�w���KHm`I�Y���9r(�|�����;��m�pfO�b2Oi݁�\�k��z���~㳺�!���A���+�*aAz�	e�\s��Qeޢb���JBX��#'�w�Wa�	�y�dޮ����k����a�{<���ܕ�\�W��9pT,���PrV�+/�D�TVM=��k�gUc�)fG�Z��)��[�����A&l��oa�ۏ$��b4�Cm%ra�hB���'V�8��V��KMp�AM܋z�x�19k�����_�e����bA��[���XTKHM�r�;���P�cr�{k�����#ł�z�����q�'d RG�2�U��qWu�;��z�ZxWs�:����d��s��C5�ލ��Y�$��b٠`e�R�C�
�0�rO���KԞ�]�͸�Q�<j.e�k��(��mP�P��G�����!�~[w6�B�%T����<7ج�YV<�N��ѓl��
��i[�ֿ;��j/PT�u
@���y��Nڜ���k�TV%�W��T�"���.�:�gXՋ����^~����iQ������L����MM<Xx@]��{��='ZE��3�RC�����*�Rŋ������?V�x�|�������>�0a�,j��g��Yõ��?��XԱ]��O$��rp���4�S����̠�Rpgwj�A�2ҽ.eh��Z`���nN��x9�s5/�8�6�Dؿ��Cv�|�l����� !��"�E�
���y�*�8��5�V���Q+5qm�tUhOo�7IHHZ��Ij�|��kS���.�h��5���_�yS��ȕ�T�� :R�����X�W���EwT�������D�.��r����wҪ�yV�	>��mH�SU���Q���|�؂��$�c�<o��@ݻ���+���;"	"�1��*��O��D#�B�QX���=(�v]w��_�Q�K((�缿9��K�J���}NU�hvfk��'����q}'��|�`	�\�n��8�]�Y��
&��^�'�К�h=R�4��"U�v��{�0��2Bj�����?����Ĩ<+NK[��Ƕ�3��n��.S�Ҽ��'#��N
O��-G	�0� ���co��N
D8�bɅtK���ki���s��d>h�|����Xw �^��u�Uw���~7Y@�tcC����K �_U���%J*��O�R20b��bx�L��<�&��#]�2�Y�d,�YؔJ�2׋Z����-�_˫2^����N����-��UYg}L��H�8��8�w	��&���t�F��[��vh�*�}��ܓ���1��Z�g�t�]\�kM9�|��?��3oS��|^�[>��%�.Ꮅ+C������X�)О2��<x����
�>ڥ�˕�(�#"��\~&<�<6���>�2�'����ɎQ�~j��}�J��;��0k�Kx�@�=��"]F�x;i# 
v��QZU��p�ju2��N�;
Op�Ö`O	���x�ӓ'�Nϡ�K'��W�Z|�בK��&�	����v�U5�����S.�/l�����uQ�}q�Mw��P�dUZ/!�	Q]��i� ���r
�+j�WQ�~�'\=����j��%�`�#*_��Aߏ+`ҹ#��� ��9�_Y��Ղ��&k�2E7�����51��E��/Q&oA��`��G�����RzG�u[ �����mI
�X�x��~�p����6����*��3N���]��F1�%��@��c$�� J��#�쀛�^��DH�ݿ�`b9��^��ݽ��P�GSO��<�����3,�#���'�(Ϳb����]fJ�RQ�XE'=��3'Ů=Ng��+K$µtc!H#���,n��q8pE���q������[.5e�,7:p!ޜ��j;�6�U����O%Z�m/�8�+����Ϥ�\��4D����{�H��Y;=���U�ׁ�g�t���S��ֳ��ڵ���ڵlD�����m����b�4�b��'eӁ�/�㜋�a�$Qэ�"��k����tD81�Q>�|n�bE���� c� ?�i�r�ё�%CO�:Γ�3���AsL
����16T��gݛ���q��_(�Ļo6k�&F�2�G�HɤH]g~'V /���sؗ�s?��}�})͈�d+~�,p���j����:J��Y�`~�q"x!Ŭ}�עӫ��2$tڷzW6l�|"�Y�%п�bfj����~����s�c�<��<N������P���Ԭ�ѳ����8UX�GyTS��ڜAn[J��v�r���YSj�ȇh�bsm�5�~��ީ@��;E�*	[-{����b�7R�D���8J��*�!���N����3ޯ`�crѕ�9�i����? Ӧ�V�z[jkb�#����a=�	9�����_xZ�JL�O��!�o�\��\��� �/��*��U�J�'a�%�_qC�T��^]0�u��O,%QFʈjBy���^�h�j��bd����+��YJ�＆��>Zg��>��$����?�(���C��ݓo�1� f��-.�R�q-_�DbV����`*ݎ)���,`��"}Q�=b�n Uk=�"�(�*����Ԭ\7V���5�D���7�&�I���5c|�gc&�T`�tE�.���uC*Ec�2��3Ӗ�]372qؾl
k�Y��xYT2ڠ�'�뾯�w�(ǕQ����ނ��.�w�핍)m��:��
1��{�>AUҡ/ՃJ�)��%��=N��M�'~K����*c�lV
�=e���S�OV%#�"it�F���O�U�*�� ft�����R�8�\��x?��}���ۋa�Ј��������[���f]�r	���훘
�]ο��5�Pt�J��:[�Me&��;���6�^�TA-��~q�\��CI��_��QoE��z�"-Lu� �)e�U[ 3l�AT�����j�C�V�KG�Fv��R ����0��V���ns]��Cq�hQ����V�I�
��ʾ�V��>[S��[�� x�	������i�fny562�<����/��VM
�K����Ҁ/3Z3��{
~�h��B�F$w�}��G��Í�!��2G���6��l|���3��i>��\ҳR�?=�ԅ���Q�7�����09�k�.��Y\��.9|	�H%�����%	����Rlb��{�U �����6X�� ӛAi��;�]�Z-�#��D+T�ɼHN0��:wL��30��o?s2�\����,�wl�<�),��gЙ�>�7<O��9�'-@&����˦
�����vmq���J?|�yw��B������sQza!���*�}cC�l�Lٰ�����8�'&v�#DgL�WV�a��.+��G6[��Sɚ�Ac@e2�ap�zӟ���$�Zϐ+�����	���=Lseh*��(ȃ���r3#L���X�g�����h�ICo(�2#Y!O�mf�Fw�Q��;1�Tj����õ��<� 
�n���1`��'=�&{O)�;�6��qh��:�!�K�=1���S#�q
@�O/�A�P�6�"[q]�`\�R�E��� �z�8LSb��'_:e�#"%e��x�o��hc{����Qg'�H�f���D6�+?H��iن�f�.����:�,�ͩZB�� ���ԘC�Tm=|=��tX�ҧXa��t#�8|�J���f��f��L��P$��A-���(;�6�?#�2*���A*(�V@ˑ7�_W�)�x��q��K�Zz�.gˋag��#u�^��8�d.���X�D}�:���FƟ>
�hD�'9�K���2��ϐ�¼U�8ƙ�X0�By&����'݉��v�0�'Tv�kiP)���V�\KL�;c�;h�h�̚�vM]�Xy�4�Ҝ���](AEە�IZe�T/b��Ǡh�u����+h{��^º2�;��X����Oh�EN
I���`��VX|y���c>@���܊u�Z?�~,p��U��F"��u��<�;�A��A�oH�o��e�կ�f�ۈf1p�tvx �KG_@�{ed����y�����n:~�����~K�f�
�_�g��zD���l5��c7ˤ��:�l�1g�ӫX�Iu��y/+����hJ��c�g��	�X�h�]ࠇ!��`$
C.r�$����)���GA�����TM��αI����-+{h�;�{I�����飐D�E��Ϲ�G�A���o�t-�g� �hjVtn)tz�'�(f��f7���*.��QX�]Į(۞k����m&i��<��faO:�Ln�V/�]H�/�Q�ic��Ө4��Y���83
H-Ɗ�L��I����j�p�L�3ݱ��)c��8�vo7[f�?y�I��Y�;�C���ڪ�
�bM���՗�9�f��+���5Z]?&=��9��e�*ߢ�پ�� �#�p�"W��8�IP�@wm��$3�0 ���\�X�m�c�).ƬUU������n\����BN�f9�g�������6�o}h��G�N�"�(�~:rW+A���ϡn)�W�H�gH8+w�ئ�~��|�/�}i���� ��J��9x��������e0�zuE?e�a�/+���f�l�ۿ}�jZ�\��t��^ݳ!�S�2���b�����O{����l[!;���`����2#�a':���0PF�v,�;��� ���4�ӿOi��`�iZ=�O���3k̰�`m�(�2�`
R	�q&����qX��]���hp}���y-���6��4}2g�T�� 6�S����c���4t���-Q�����.V��F��9��w�\R�>�;�M��KU��kۣR�a��*��?��3���kc=�D����+N�&��ν��ۮ��?��*{O_��Y�q�ٟ����"�~#W�7�A�h���-��ee_��e��B�����<���i�E���zڜ�
�Eì�^��9C�m5�K�C����������M�B�c�ka`�v/��V�.l����*���<����YhI�*L9����d��H���&r�D$f�ҳzɲJ�Jb�$�r��ٯ���g���QIG6��9;ayr;��k��wM�g>�|���β�&�-�/��h?���ԑ�ѷ�F"nE|�%8��p,����1�®�j$�V	��(s��1?����+��i�]�!��`�y��I:�5k��|e��M���ey��G���j�{ξ:�'�����?�|��M ��rD�+���'�����S+�J�����A�$�f�N���s���e�0��Ѷ]��ZmRB�o��,v���P/V{�k�q�=Hc��'p2*D-�KI�Xͣ�Q2�_�Z�Dd�Y$�Gl���ଉN�b����Į�v�!N�s��v�bh�giYӚ�[b�u�����b�������L;Gf�dU�v��4^�pZгĸK�ʚ��Ů�f�a��N���RXG��?���[����.2��3�u3��|���蝉�T�r���{G�(�Sں2�'����N]����9�5�r���!ʄtFt��tF��`M��$ݴ'�R�����d�K��x��10�]VY�I�Ȕ6����h@�Ti���1\��RsǼ���F������GT	w�u�&^� i�Izg���l�S�p�`H���
v9�͕�M���U��Jn-13��&��M@ �����}2wSkuj�1W8��K9:,��ƚ�K���_epI��{��6J�CY����`�\]dED�E�M��*~�j��P�+�2��X8hң���`I|Ƴa��[P�ON,~���-���J���xN�V{TJ��P��Ԗ׶���ĩbw�"�:��8yR)�����nJ�Fo,�V�5Y|:D�n{E�n�Q,d:;@'��I�O\�8{$�ιn�������D�_�Z �KD}�%2��B����'�jF�Z;��TFx-ѥ{�8JvV��4�'V�.�N�w��*,�=t�zO�3�F�5�9�3�6����_�1��Ƭæ�9�#|�����qW��ٰ�K�$�
�+!aS��%�A��U�+��-��TY��w���^��I��w��{+}��:�>��9??�����9�&�3����z%+���H�V}d� �S9�H��o�`�CI*�sD�h8�zx5�ￕҷ�?��xu�0�
e��'l
�zυ^C�Y���6�F�[x�-�]f���m����._�i Zfw`M���=�G���c(���q�~�!���'e}4�ԉ��Z��)3�!�Yo����2����e�uxֺ�����C�~����>E��u��Ow�5t�Ƶ��m��ݺӵ�0�;v4�Ʋ�8K[`��L��]���\�rr�U���L��<o�u»g(�p%���`9���<%�A=M�"�W�y-[��9l��uui��)?�L�$�}��mv�;R�̞��3��d`F�%��3�fm�����P:�gхQ��ܟ>I�%��-�\z#��8]��»���/^��?s�^6��&[_�	m�D�Kt�I�4��^^�ɝʢ���=�PZҏ�U�����~�0�������s1TQ�/Gcj 2/6�K�'Hw.;HE�D1�p�B�!�n@���h-y���#?C'#D�P�`5�9C� ��U����6O����Ӣ%���_� ��5�p�:�0��<��c7ˁ1C j��Y(���Zv��K*�}����Aِ}}�l�Ji��å
���S���i�M���$��_��pa�h��(e�M}uۦS!���UB� V��)�	�T�΂���=#��)fF�s��˼W��}&*�0a��|�l�|�y3Z��>U�q��Ev�G
�<��vE��F�����i��1��]�gQ�����n�H����v�c�-54yt��u��@�Q��!jS��������9��>r	M~_H��]����N�o��K��yX���U�떃
C�\�[%J�"H �r7t��R`(8��1�[���"a��T��Ҳ�0�;�`���K����rg�UC�uaݗ������wO`J��2�����r~�� ��#ȃ�dSjk��D��`�P���:x�(�����N��f�ܥX6Gx�f�#��e��15�R�C��,��[�������%��(�$���0f�W
*yA��E���䫁�Rfy�1���W�&'��H�4' R��᷻�e}D�p�4��F���&o����_�%��}su�'�S+��ݕݰ:U	쾬6�����������lB9鎈���o�� ���oe|���a�P@Ԗ���ۇ�G����?�-AN�Nܥ�QGb�z|�s�6�םFfU#��r�π�u���.Y�bf���e�8� ʆ����l� +ȯ���ﾐͩ��m�/�J�����߮aW#K���X���R߱>����i��3��ޞ	E��Lg[vQ֔w���ވ;adCQ�0i��{�_�={�&s�x���<�|a2�f1$M�5>�,h�O����Ǹ��"�Ґ��]����k�]����|���t5�M@�7�>�8�C�O��Oڨ$1Ҙ+�dy�k"bF(�V�5�rU uV�����c*������kA�a���8����o�������|w�?�&Fo�����7�R,k������>��_7&n���g&�o Hc��gwU�)�B��6g�~nѡb �3�@�� ���G`��C,���͙o�U!f���^�����7�������uj��׿:�2~����>��~���v6�M�c�ˡ�L��kx�p����j[�P��X��G{yY�:�1��U�� Tn������8`x���f�V7��{���{r�ėw1�4��^�&�3�z�
�ҽq2��q�]������)�o�Z�ra���*(�k^���̙�6�b*�1�ݖ�&S����>���&Ԝ{@d��o�uɕ����@�1l~|_�T��$���u��lA�>OH-Y��䬥�BV�Ϋ�0K��d�P7��VntG�����W2�e�#E�*h{����^٩S�\5��c���H�iδ��G���ڛ����l��2�Ք]��,)յנ�>���c�����;m�C+���<z�̚y�x�"V���j�����8�1USn���1R~	M����O�D�[�:0�[���b��H�UD�����β.��ry���(F�DC��9۷��Ԉ_��ol�z�.�jT���D�na��C�I��������+@�l�����<k�ӳ�o�WL)6�2A��
�OYO�-{�0��~S'�G���[�@<B���O!j3��=�ܐdF����CʷtJz�`@@��m5 r�d��]�J%�V��I�\�Q��8�ޙ���U-<@;�Na�OBo|9Dou>=��]�12f�9k�`Ij
'���P,��z��a\�Y���&K%���A�d�y9���|i�4��_�qC��{��P�#'���n�����B��
*+r.��*�9'���g3�|�ɐߍo,[��T��5ue��{E��\�hzȃ���Ğ�.M1]��z��ּP<�t��L�����7�����`M�@Ҍ���1V#��"�a B�xߍ�������̽�	m?��ͷ�m6�]k��D�����u��	��+��F��Q���In�x�}k6N5�����H�f᩹&�ҧ��)kԪ����JE{"��&xLE��sjഈ\�`���W�zz+`'1(����Uw�	�b���QT��Əb�{��b��>uw�2{��G�8����T��**�۲�1������d4��8~��|�����`v�M�ے�X��P���ðe���\F������u��,`ټ���]8X��kJ�$�t���>F�1��9�^$\=��n�ś-i֝Sl�0��k�����o���o4�x�0Nރ���#�"�Y�؇���y��o�]��e��:�#��M�*�F���E�kb>���I�eY��@�4)a��P
o��������}UC��]��(}����z�A��i9���RJ=������6�?��b4=֟�;*�2}��#��D*��\o	&w�h`Tmps餩�w/�f��<���'��N<�Q^-����6����Y�����`�K��6��������8]�kh��ϡ�	֕�UB/�ѩ]��$M��>�'VN�i�P��SL�%5)f�#m�!4aB�ݮ^oy��|�z��7�+,�FT�P9z��o�����s�x�o ;�)��Z3J��{2��#2,r�w�50������[���aP�%(��8���|�ʮ�x�#5߬9�y�_+���Bӈ�H����(:t[��ߡJ�l���ĀFaq
v��}M5y�m�:E�в@��M��㠶�㽬�c �#SLwզ,�R�#.��[AaB��,�$��RD�PJ��T�qE#h�Л��u�7� �?D>uc%aT|���@�B�vH������)�fyV~��a���$�c"vc>�	X_F�1��u�O�O�+�}U�VgC{�	�2<� �`�j�����ܩ�0����u���;�tڹv�������e=:n�N%yN������?m�GH��9�kR�P{���?�[W��آ9�`ij5�������L0 3ϓ�;6	�A0�ݎ�����d&�Q6����yH>2�q�@|X�
�����o�Β�Ed"1�F�α�2?j�(�k�i~��!��=!xv�j�Ϛ4
����]�	�:���Oლ����^^��&o��6���\)��j����"�9V�^�S�H/'e���	�yo�BtBf�K!��p��b���<xٱ�p��F�ixۃ���w�f���u�G��`���}`�6��*zY�ǚ�jbyKSC����� h�]�X/A�}E,�4�,̤�������{O\�y�k8����adďR��a��-͙�:�5����0BN 5�$z���v"ܐ�1+��bf�O�$��qa�}�(���dQ�+��=c�¢B��x~5ᜟ���Kr�;u���.В��&Q�}�đ�b0����cq�qB�6P�s�^�bA����a�w���;J��Pt�h�.࠶�$*�E5�3r,o����(��+��g���s{�q���13l�驓�"������+P���Vp��|���wb�X�N�xΖv�\3��0�.�)�n��D�/4#�(���m~$y`�����9#º��[[��GԸ�������^�7���ݗn�Y?���;�޷��S���!x�6�����Y,f�.㒇#�C`z�T��!�� ��c�����dh�}�9��[�f\I.�k[##�P�����ֻ��1e��7�z�~�}a���",!��c�阩K�vCzV�	B�F��I�q�uɃS�~Ob,��S)�� [E`T����.���S�����)��ŔO�B��1m�zE�-���}]�6�Y�j�+�y1�9��̂"R?\o �a�����C=-I����ەx9�fs�%pfc�>�D�!-"��|��m_�2�(�4�x��Le����"7j�� hv��81oz^|9W_qC��t��c�g{�TF���SZ�/9htyC���ɯ�6�0|V�,���y�>:\�{�X��5�i���ՈR$˩rF���5UW^`�Y+�<;~��{,��������ˤG���('�
%o�\�V:���D+`�a~�����Q�C��z%�\���tG ���L/o����
�+�-&{!1}�����W��["*=���ݜM��輷�R����ѳ0�;k���X&[���<n=��f���3�L��fp�e��~?{�8,������]>��qn=��%��m�?�Pi�z9!Cr���	V��{�bj��O%�og]��tc�5����H�O1(soR[�CXYb��+�1ʴB���b> �!��=����tEp�̹	�I����5�1o�PeM��)�o"�nm{AY;S�;��0��)9Կ}��P���2N�({�xb���=\*�C-��jS,]����ScW:!
�}�<	�(t�;c���<�[�s�]P����;H:{ (������Mn��"+4�މ�x$4��c�':�v䮠7sJ^��� l����\+�SwK8)��=Y#��#�3�K��\���jw$u����*-|7�H��3"��?�rn�X̨���8&��~Q,��f���o�,6IbC)3$��?Ŕ��U�RlK�ěc��uSם�6���{��$�(��I�=��Tv��2;U�p�F�i���͔��E�K䤾
� �we�J�K*� ����؀(m݋o}nab�\M�U��R����Z+X��vO�0�]��p8�i�h/]�i�Qo�;��Ǆ�cА�X9���`ʱ����%`�V(N=�e���T�
P�8X���-��:�Ft���2	O�i�	H˚�h-���Ƕ���$��㺗�f�%J��J!z�P(4���S�X�e>����3z>�m��,#)�t褒����i�ν��1��{�G;�#䡜��|���?`�qv��Y��|w��o���:��	���+��x	_.!M3�M(�?�<�Rw�a2$�d�;�;Tvې�va�t���\�M�K�\��dt0ꑿ~�|���r!�R`bQ-3��ѐ�Ĭ�4SB����l��X)�頠�y�۵Xt�P-\�RVO�ޅ'��i�[��c|(l:ݹ�>�/t��t�ƛU��\�����9�ǻ�i���C8��">\���f�
}�Q#�g��]�7�f�3�:b��DH��� c�r]rlVؒ.-x��Ia�4b y��ʢ�����P��{�i.�j[ c/���5G9�^)�p�t4�N�b�*�Ó��֡2r��� $����&�Sm�`�0!���������E�.�؎�81]�D9���]W�;\G�Kٴ�k'���\J��k�h�_9�W8C�=�?k&�ǊAJner:����XUPD3���!i��:�724/#�(���{a�ƍ���ͻw�-��*$�^��Qc��"���{-e\��/o�TI���y�!�x�ez��{h6��h�]��d9�����U����O��b�i�ֱg��^s�X.�� ��v5JEg.��XA�ω5�7ZdD�W�Z�D�J�=m�&ŵ�i�r�Opٲs%O���r��LbgP��+��õ����ȟ��i�Y������].�Cr ���e:�����l��d�/����<ж=u��o=�ɱV�p�	�>�]n����9PST��]7�P���T��`�90Y836���dx�,'-�<�}I���͡����^�ƒ�V!��H%��?����޹ޯ�V��)\�h1ߗ~G.�j�dOo�ۀ��#8��İ��.A���o��I�ff[Z�Lu�8��$I)O�V%��C�f
���PӄctC?�D�e�&P��Se���5
���Nw$F�i�2��'��4���(��*�{�u.XQ�H*Lݎ??J�*��A���z���V"Z���v�<g�Jc�r^��`����e������;��~	!^b�lB��2�ڹ{���T1�QD��-2i.����H�o�b��g[��ղ'�C�W0��}�S$Q�@�G?�t0ڀ��C+�e�5M�=HZs��}�Y����Lf�ۈe�j~N�t�X���2C@��I������ŬtY/�Ғ..ٳ��0�6��VN!��I���t!�0��XI���XԎGq�{Ig�Ί%�S�a�,����}b��L+[���Z?�i;yAԙŻ8���+��\�
����u�7�[]s�f^�3ꉇ������6O6�PC1�HLW3����\�쵳2�N��^�Œ��_Ԟ��U\��qt����.jR���/+��m�Re�܎��?��T5nJA0��佚=wow���Q"+�_��P�T���#��V��Í���	%wU��qK0?��p/��p.�3<����-X���Lm-��]�I�[8��ַZU�w�Q�.�h���+p�#V,-�w��b��?������5�U����^�Y��Z��K�ӽ �y�( d)ј��k���
(@M% �Xh���@lȖyU�y{�	ݳ��id^������B���[�s�.H���F^>=�G�t8%w8��'����>9`=����4Y҄X��I�`64��<q #��WhҬ� �},�BH% +׼��uO�\-��?��K��y��-�<��nj9D��Qߍ[Zo(�c�����NI�R2x	1Ǡ՚U\^��G�9�V�o\�e�[��R[��sқ;|�-�6{����ڍ��L�k�g�<�]�%���jT��&Is�f�B$$?��,�+`$wع�ZL%A)c"jY!��~V:�H���^эtA����T�2��[3r����QU���k��Ec(o�c�8D�џ=��.Wm�ߐ�h)۪s��'Z]Q�f
�})%��7@�E1�zL_#���.4)?�Շ�Bs"�+3Cm�����ze��hIУ�D}Y��H���/A[�/��v�t�Q5��:A9�Ñ~^{����RA���!Jj �\�1��'E4��� �]�� �C"���B��0����U�ub�e�
杌B��6{W�OU��e��ge�َ-+n����d�
���&C%����L7����Cڍ�'ōh�]b�~�/�8��w:-�n�X���8��{��x`d�>�c�Ŕ{���("~�ECZ&�T	4i�+����|���`,�	c��ւߛ����%�z(��K��{��x,k�u����LjW[�2��cg�}��r�W��,r�D��բcn�q������)��k7�&��;0���
�0�i[��Ud�b��!!�r�:;rd3 �����d��:?bE��<.)O7�ۓ���s���I1{7�35��]��i3�559��Ӑ��"���v�� ߒ0a����"�hh��0/v��Gܬi��/|!"�Ne�س�2v]��ܛ�CbdҞy��rhy�vfkn;���� Kk�j"���}�|����&V��M0��[b\<"rN�g�9��g��r���A5sRc��ǣ�s�F���C�hÂ:�#���l0��[��N�7ݙE����%v���M�[�	�,Z�;���vU�k&�ւCͳtjM��Z�����<��2)��=C��dn����e@X���]p}�O�ຈV�w��ۻٜQ_�H-̻ZU��k����s�9�#���CR ��	#���C?S7�
si�s>����(=�H��-�H�tN�q�s�
9)5��o8"C�hG�t@���ȥ��=b$-J	L�0@AC��R���E�"�P7bڤم��X���7���5<^D�Ͱ-��Ԁ��d[�iS��2����!Y��vZzf#2X^���F���,��DE~��:1�i�>]�:IM6����� d>�������}����I�P� @�l:;��|W��ࠤ�~�R:�!֐ywX��]�Ӎ�3��X��l�;���SSڮ��-��i|闌/��jo��ܕ{�eڸ�C3��T���mfc�DS d�(�L:���D�`HEnsh�)!���K?5$(���*�J�Z���I�3!�Q>}�	����ٹ�g"�x[o���L����9sr����`�R�e�����2�i?�6��~�A�!|��N2�ʪP/���I��+��Jh ��	�aH�z��qF($]���kX�Cw�i��|g@&�/��&����orE�����#���pu�rr����T�j-�<M|��!��UA%�,+�� ��`_D�w5u�;�?�c&=	<��q"�0&����>D�q����g��L����������Zq
5�%�uȗ��-�R�|�5����3�r�nb���kDHl#\g0����@Y����.��.F�i2��	z���!����y]��$^J�ؚ��\f��,�]�S��#�C ?��U�]��nX��]� k�XLS̠e���0�J��ɐpi���S�������\TG�!cr20ZSm�k��A_Gnx�RZ��C�?(�{^Yc��j�xzb�\�Qr��x���Y	�\[��'���l��u��5̺?���	b6�G���9���+���Y�R�ύ7[�l494�!ab\����+P��QOL�j ����M��a��OUh���=���e����&?�;��T�#�	�G+�������rw�U��7�J�p����㬙*0S�@ >Ȍ���-_��f�w�`�h� �$aޱ���z:#�~���ذC��*9S���+G58�ud�o�|o�!:�
;S�u>��z/�Bn����M_A�b/}�WP�?�+pI��0�:}`�KX�O��d��I��{�ɳ�M��3�b
� �F�Wש��
A�Л'ǳs6��=ū���'(�a�7�p�L�:�@qL<�}�$r��Ͻ�4i���\|��Ƅlx������A#���"5:,����k������C�Aiy�B�p�j�I��u�ɿ�ў�/��Z>��\��d`P������2�3-K ��|��W"z�܍�y�!i�" J0m|2���E&�Ji޺g��-��v �7T�Ez}{Э�ܱQ:/��0+��ǂ*��p�bu���=[��[W���q��_] T���F돭�ByN�3?xt�?[�hBi]���;�!�J}��ͬ	<{T���8iG{�;�(��<����\�>-���c� WQ��F�	�� ��S�hP����!vI>3�h���O)M0Nl�H�D|���P;^"o�'?aR�$�レbSRO'�^M�|��7{��d;��P�l׸}2�Q�V5�7
��U����'\�W�cq]W��v��*W��f������씆G�U�GwN=#�Qd^/�X��0ۦ����bu��-�ك�1����[繉�B�.�c���ͷ�g�Sn�pm��2Ϡ��I.��͓��t�������dr��,�����o!�FVhJ���/1�� ����Z-�&OR���k���Q�\?X���Rz0�0�:���f���6��*y�F��|�>��U�k�dl0t&E>����

t�!��Gŵ�٤Ԏo��&��f�թ N�n���yy΀�n�� �v�K6{���ZI��X8KZOH�Q����� �UM-��q�R�x��s#�����T�~ ���{<1�Io�%���<?\�ZV*��bf����fBZ�9��n�7U�e�<&e|(�2�%�v�/�j��w�^�04��].w+D�who�=���ҷ&�ͽ{�W��z��E!�lB�M��`�&׍B��P��N�kt)~@V�Vg@#����m>�]3�dץ6� !�"h�E8��Q2��}�-�Y;�iK����뿬��ZP��
��r��+/+:�:zdU����V�W3��3�N��4��K�ғ��[L��L�|o�@��&B!��C�<�yo$��������z?� �t���v%�:�ľCf7s�H`,� ���E�1O���WTLL(�6aL�,ZKm~å��ӹ��T��Ke��M��eؔ5�x�݄3��S�ilC�a���h|�yV�fԌ^_OȃqFv)r)<���6|y4�T�� t��xX��Lv����&�P4�'�n��B��T����2�#�����}i�W�hϒ�q�o���g?{	A[.���/qqϤ��N6�D�}��X��,4�N��r^�MXz�E:��	l<�����][ö.�D'�e$�M�!�w������=]�VoH�ҩ�Uw���k'���܌FU�"gT���)�Lwn}���(��V�8����L,u��T��o`B]�5ڣ�L-�O,7��k1�]j�1˨��A5/n�GqȄ��ez����Y*M�TI����UXj[�bA��p<~��|�O��Ф[��x���§�vщE�/ "�ݖ��H����1�U
>���\�~����E�����^�0��Q���9:V�Q>2�E̤J0�����\DtΤ0Q8�T5���7�`���TK����I�rp�}}��f�n����1%u�������]H0 V�!71����~��\=U��W���aYW�����\fEU�l��Iz@��0� �a�rm�sGQ�����\�J,"�����I����r=��$�}�����(l�)��*���v�}����|aw���R�1j%�&F�>=�KIh�W�蘁��<�"1i[qp+NF���@���i��'��Ѓ�xS�:ܺ����=A$P�u�vJ�%������g�oq)m��,,C�ы�^[���ի�:���C���@�|�%�b(o�4P~��ƿgb�oj3*���g��]{9�N�{'�|(�� $�P.�N$t�P}��ש��3����<��
���1���d>��ǅ��I�^ɻW��� �ǭEK�����X���b
��+㞒���OJ�_>ơ�J�B�{T�r�Id!b	}�7���V�I��s��	� �lx/��-������N�[P�s/)-atE��=K�K��x��V��vA#�ȯ���ǩH+h�{I$���G���2b"}Kł�xO��ʕ�:^3��6:oFm߭!�Q��>����'rob��_	�n�n��K���wm��:�r��N��NW��"��8�G�G_&�������<4@矨v�D���BÓ��I��8��j�44���ļN���
���X�f����xZڥ�\t��^b*�R��h��4U�b�'� �-6��t�0�"
�	���c- �%�|ε\��1Só!��c��}
��$91N�'���\�x�C�}�iҗE�����!� �E.�+"���h{F�t.d2��n��������4���L:���D��[�:��˦i'�&�˵M��4xC�}�Y� cỷ,��=Sr}vbgEw\�цD��N����.r9��-xK�lfE�1�x����`7��<�1��o^BbQ���,i'� 2�ٞ�qq�C��S×2s)��^s�x0iL�0���>���5X�~���ڥi2G�4��v�.c2��)�z��Yr.�mN�%Uq�D���E/�g=��tݕ@���Q繿���m݊����c]��@�I�����Ye��F�C�%�.�l���}�u	���f��w�2г��E/�v�UΖ��$��ѥ��q����l���+�d�R�����~XQ���T7N4��T�^/
s�D�;N�>�#���s�9�̞K�#��/�s>�|R'*K�z��2���=A���K��c�� R��[7�9��k�.H��}?bzӞ}D@��Js����7@�Ѫ�C���a>T[l\c�dqZS6��N���a>�U���;�c?�#��:������ra�?|r���K�|KN�x�)�\[=O7�In� G�t�xx�)���ym�cK��y���S����wd��2d�Ã��/��Ի���6{oh��,m�D�).���N���q��A����i�Ix¹Y\k64�j�Xl��r�rG�DR�G��p�c�&���AV�5{�=���	�i�D 7���0�Dpz�c#vRoG�������m�h�05�Ѫ�ֆ� �|��P�*?�|�n�iն#r���oi�M��b�'l#+R�%z�0�srث��/z�T1����'�Z�>Z+'.~^B��￭�@�f�w�v�wbj�,�Vc�)tB��է��A�s8�|�S��pՀ�m��4u�T���v���=p_g֟P�l&k�5v��h2��c��dz���Obv�e���,�Q�93�s쏅��9:-�r�2�᜔�<�a�}�ב���G��Qj�z�I�%�U
h�i,И�������ӂC�oe��P�bDba� {JRR����4	ݾ��� �����W㏾���h�܋��<��Iro�&!�ݚ�P�7$��(����]P�*+�2���3�<�D��ɯw�6�Ģ|sfڕ�r���s�ֈY�2 +t��C�1<�9����J|��y�!ᖤ7���%%�ZD�>����ż�T�����l����>���I�3�������'`�e��h��U%��P<���g��d+�2�j�^�q�K=��[�B/�X�6�L6,d��l�F�	ϵRf�����2+u�"2뫎K~�K��1(j��tT��[�W*��F�"�ZE�nm���ʉ�rTkwQ6Y���5G�c!yR�S"�!�^�C�u�M
�<婛k�t���OZ�p��y��D��3�PD��CI��B�����B����a/w �ZC�X+$K���Y۟������;���DC�|�ݝ�A����w�c�4f\�LK�u0)�q�J��DxkcՂ:n���w�+:R]�=�Hb���n
��a^8���K�-闕�2	��:??D5Ƨ�=Wp}{�E
��_}��8���X#�V�R��T���[��-�I�:Z^��_��w�S���PHR�D"-7K (�ـ��8����������,]@"@��-��OeΛ�u�����J;��R��U�QR��ʜ!nb#PܛRdԜ<��N�O����H�T�>�Ws��a���@�{q���x!I���t)���W�S��e�qR󙾒m�{�|�h������4'�h�wD��q��Ba[x5Ȝ�c�7��O]���[
5f�u��|�Y�d�;l�hWj��M�ˉ\��K� ":���uf��d�F�f�Gi6����уǹhזi�
��v\f	V�w��@JS�K��z��6�Z�-I:#v󸥒��2���y��9���daa�����$��[� G��F^Z�+��K	����U�u��l���h��E(v%̷�3oc���9>�aV�t�,`�Fd<1-AA�����T`	Gü�F(Ə�}��DqM���-a,Þk�u��K��:����rW`2�0��K��s����<~����+�`vr��)j��Z�6�)�X�Ӂ95�p�S89>�813�DB{-�W
�C+Nu�b��'�e���C]��g�Ph%�S��չ��z�/�3��KX�����s�o�2-P�-���~�Z8m��O��X�Y�xT�2����8[ď�����rlA����j��Q��3�p��+AV�)�e��\��-*�̭[��WF�7*�2i��f��%ڏ�4 �y"�혍�r)�K��	~��vkd�~�:4�/��#o�K��P�	|=����,�h�9 �H��7� =m(�Xv-��Z�/Z�3#��O������!��3�.F�W��M�&�!)sH�]-%�:}���`>W�,�܎�_�JD�=�)Vz_�9�=�`�a�P��
�d�\7^ܤ�Zݩ�;�r�l1S1������P�lT�~��\Ě��\�M�w����?&����g��gL�q��c-\y���̃��7+��b��a5�eM8Y߻���,.������I|<�S����	#��L?tc���5 ����n,�Qi�̴{��ّ�6�ư&����"TJEX�OH�� ιA�w(_9���]E�,�S��f]sم�l��
�ϟ��t[2.��^��e����}���O�dڵ�"�{v^\�*@=��
���4p�arTs���[�h˩g�3�kBk[��kZ�/i�.��@�����
U�7���[���%l�p��<#�/��N��>�����.6�A����K:�����vO���$"
t�kr�'�&�ѹ�ܘtW��Qwm^^����T��������_ED�@����<��A6W{&�\�W!F�Khٹ�$���Ҁ��C2$^>��Y[�Kc�l��;������MMXR)!f�$Ik�z7��ہl"W=!~��,A����,���a:Jvn'O� �+���-u�u�����W�d
nX=���'��r�4�t�m�|�q��g��y�}N�Hz�lnY7H��=�b�Q��sm1{�0H �\�,�	E�>�k�%��lx��;����c�)R�":L�'�j��W�
G��D[m��~���C���N�nѨt_��Ҥg�*K\�]ϊg@���q��cمh�D���e�+���):@FvĖ� ��q �`}��)�{�-�tQF�	zF),6#��64OE�KD��Q�{�g@�0h�bG�y��Cj�d~yS����4�ރlH��(�1Oy 0aVs��F�G54�B���1���4�����\�� �l���=���#'L�ڽ�P��u#�ax�����
O N$��Q@9#$�����#��K�����$�(�ʑ�өc>�0�B�����i<�d�|��G6�h����V n���� vZrl��&F2w��1�>o�s4�I�&�������3߁:���"�P����3���s���|\W�bMJ_�]P��L�.�]�~�	|��{k%��((���~W�[9=��؍l��*�B�N�>_�A�Z�>��9�W���}���8����0Ѻ���s����A���zȲ�k���줓-U�x��}���8#$LW[��B,��J^s)H�!d0ٰʟ6�q��߁0����s��T
��C%�VFi�8�7>�88afQ`�,�8�A�4��ӻms���[<�p��J��	V��w�>�׼�		؞d	ԯ\��
u&T^PY5�A��H���9��xcn��T{�7�Z�B{O�|Ї�}'l��Ҟ���p�i�R+�t�����g-؂���S:b��1���yZI��~Eә��GDF^Ky8�����=��ݔ��2����՗�2>�J�~�'��^[�$��MU!%���/�	R�gtX��rSP\O��W'����� ��Pa_�g'p\z�)���^N|�vW	�q<�`2e8<]������'�	��w5˦aT����΍����\(�q$�I�7k�BHA���M�����0�O.a�����~����6��K�͗����x�t��+�*9p+-�<5���;��v�]����|�E��$�j��ߛoh�d�:�q���*���_��۽>}��-���ؿ����Ѡ.|�$T���6aw޸6��Φ�9��J P\=)��`���UFw'�Ȳì�
/�l�J@w�D�wY������� ����=��tk�M����D�n�i�����X ��A|�d��"t#ʉ�����^d,@~���F:׏x���cR��Ҝ�?����� X��6r�ʘ"ĳ��c���u4g� �؆��A�0�ŢA
�J�r��:ѡ���~�VMH�ş����9`��a�7�$MVJ�
�Χ��W�&1Q������p��\nQ.z���#8�͟>�\�G���mi������8z2=a��0��jQ��S��p�0���ux!f�G ���ډ�ب{|$���B|S�7 �� w�& Cc���0*����<����-w��7Q��iaS�*�n�fucW��r��#0 �|�x�ݰ�H�0#:~t�z?��.�ᛯ'����"򁁽+�ٺj^8��w��&�p� �qY#͇��ٛ��gv{L'�_�X�w�{�8C��n��Zmt-���;䍂.�d'Ru�k�I��Z&旲n���VDF�u�!o�[A�֎���μ#|jf�T{�Ð�+ѹ���1�a��f���Y��;}4%U�1�=�a��E�vQ�cR�x�:�r������tݭ�q/�O�@,<�Rw���׿z.~�ˊ�R��H/���ٹ�f���GXh�f���7�<2�|R"r�b���H�VO}�]�~(H���dtZ��)Ih���[�^�W4:�H��~?fd��� ��b]xa�B�&7���#F��M�A0����{Z)��}4�ނA
�؟�I!�ξsW�����m4�X,"�P�R�.���#�[�2�$�3�	4o	e�qh2N!}�����Ў��H*��z�޹�v�`�d�r�|��˃�?[g":X�{o�G��(cJE2@']1t���@/� Y=�:��sK1��d����(��ѫ�TA;�Y���d�����Trb�%$�O�3�\; $��<������T.&�UUϳ{?�Z�N��'}
g ���f(�eh�6VFf\{.�g$�5c�$����-�I)�L�\������"2'�*�)��Y?�hOHLy���a�$�� �'�uL\�i���<h����эG,� 	ƀ	ݫV�(���5�?_�><~�6�~ �2^��xN���КVT߰X��zF�Џ�P�T b,�>�G�1ׁ-lm	j� �ŲCW�r
����%#�P�k��5l\�t��CL>0w#�$GkW�j6����5:�N�s��\�%]��EL���tHnD�Q������*מ�NOH�&7|<8�&~S"��=��-{�c�h�DS��XJ1�`ZT&�EOs�?cU6l���
�e5���eL`�~�s7x�{���f��{�_j�����K��eʬ�qzS�p�9��vA�j��o����ռwy1�8�1��4��r;��O��T�Y��Gx#c�W�&Β72�H�"f���^\3�.5���l��)�����~���#�Rw�%�U[�{��~��s�:��2�޼�=Y}����Y�з�=�IHb������LՒ�0+Z$jlJi��F3q��`pm.S��m��=N�s���F�3�>��_�n�_,i��(���~XjK Z��:��@�va;.#����X"@�O�k�wU���C�P :P���qǆ6�s��S��y�T�م�T�#�0��1 ��Ǵ/��}�k�Џ�`3�~ˑ^��_1�"���G?�eW~�d�b3Ek,?�Г���W!�e@p��������cSS5W��8��<�9c`� >դ#CM�����GX�]��s7]��W"^9'��O�� ��D���^��
��Ъ�yE��w�>�	\H��_�5Ы<�����CO�A�J~�i]��=6Ȳ�T�3�%����#]��4_���+Q�@ ��`;u��l��]Cg��w�D�ț�X�:�z�l�����c�cOx�ǜoF�Jf��S�9�Ђ�u�S�����U�"���蕴���s�ݓ������������iF��͋���c�H�f�__��#xW/�ޱ�x*3�9Rt���K�j�i��(5�#;��q�W+X����`��k�}Q�U�4&E��9e����w�C;�h;�Z`�'/&8��r�"	�|�����"V�}������ЍL�)��K]�}'QS�ɨfot����)r�*CK�0;�Ga�pE�%T\�Ǘ±�*�e�Ū}r|j�"�g)	�ޗ7���6bå�_�v��^(�����0z���1󭻱��m�@W��cV���6�7JA��|(��_2�*Ɵ4���)c�ӯ� ��L�Y�K����8�k�\~.D��a%�2���c��2zH/�O�a$�Ѯ�,I��
?�'p��M�'S�I7��<��?␑���p��+"ʟY�I*������|�}�E�'.H��~o��I���I��Ǉ��uc��G��f��*y�C5�#*�71�O>,Y�G"S����G�s����c`���a�:�G�:3J�јPg��gg�PC��q�y�U�B������Rr�N��A&��fW�#�=ye��!��M8��<M�E.��N�Hj���KB/یZ��d��X����ހ7;w��-�ó���H�/�uSt(x�|����"ВQ �?&��H��|�� �(�rO?����	�<[E�(����l�;�o̕��V��_楲_N���r��M(RY1-��<0�4����to�$��F3h�=P;��Zj8��gyԻ�]<�x�$�2R�l��m�S^`�Y\-:c	/��a�3�M�u���+�7��9��:�XZ�f��!��}#����h�(qQx�&ߕ�z3`��晸x�~��S�������z3oW�;�?�.oLA�'y���U4[�"[Ү3H&�\;��.�M�z�dC(�q�U�Vd�|$Q����'G��ş��L�RC���mo�&
Ak�����7Dngd{f���	+��CWZ�[�OjZK�����<q��A:���?(�-�mn�i�u ���0��,Gi��[ry-3r�<��������w�d�Q{���	�!�Aׯ4�G�:b���DT#U���9�+���f���w���e;{�qa�vYj�+�ܵ�\B ����}?J-��׋��x�{�9w{	Ȱ\yD�對N��'��; ô^"��d�$352���� KB��4	���8��Y>�5(}c]I�!��S��~����̭#�)���_P�������~�v�sq�R&�+�C�X<�?{�r�rrç���Ic�>��<�:q����-��'�D��8�8k"�!���b�O��z��Y�Qs^I֥3j�D#΀5)����P�R��Q��$��f��1���m���R����4���rg9���!�z73Q;���i.)�-5�4��*G>>�??97�9�Pz?~����^�g��3���� Q���gq81D�c����u�}i����U�s ��M҆�aZ�P�S+�$�a�_��CQ������t`��@��l�.hמj�&���y�)qG�ǜ�<v�B}����{��5����D ܹsY�i��u���׶�40ܺ6$sd��� H����]e.����T�QxŹS��7��^�<�*X���2o5`!V�2N��)' ʼaJ�V�6�ϟ�Z��~=��i0���-!�u��LP7�b!Dl�;2�m2��d+��U�y���N��=�g�B��Zq��4�˙�Zd�z�XDS��cU���
<�[G���1Fm4~`.)j�Ƒ.#�@Y.�/&��j�}М%�礟�#������h�gF����
�(�I�!�&�HxMD��⢕��Ip?q��:��'�R�cu��;Ҝ����l�! t�����m��!�D��k�I�ʚ?�߿�s> ;ܡ�9VcY�پ�'�c�
U���ȝ�*G]�!
�-S����U�|�Hy�2)׀7p����vȡq�sݹͷĄK��n��D-�E�-�.�p:��1⿣�<D�
Mx��T-��\)߀�Ŋ�݀���A�J�����Yh��&I���`tNu��B[ǔa�mꢓ�()�+"�띊)��EK6���O:<�vg��$����Tr<�ֳ�(���+��B ���� U��鵿�A ɹ�T�	��xL�#0�6o7&�^d�Sʣ��i��S�M?���|	McN?��L�UG����v�ׁK���*��(�'���I�����Q�8���x����L���\i3�6Rw�`����FӖ��["�C-<v5F$=�9л ̧�� �׊*<�x�N�Dz��ii��2M��F+I��p�Fc����=Y82=��G��q3=C��]�0o��1.�Z�.k�&E�"gC�t/�IQ���E�k��i>ݫ���_�_"�C��hx�����&�j��"�t跙�.K�7��G0.�@81�4h��C�B:���$:�!��U�\�4s!���I�ol��i3"2�0�DKe��,;Ʋv����f�/�`��M��|��S�׽m�'��}��;w]�Z� ��w����'�D!Ͱ����(F��(KG������L�$G3w|5�=�W]�{���M"GM��.]`�'4~���$3�Q{��)�gI L0�7��P'�@�!ʻ9��_��zbGGToP���y����>��(� 8�"=�(�����!�]��jAk��,tݩ~�.xȚ5B���Z���8i��-� Z��*P��AQr�V�R�1�r=��wؼ����7n�s��6ߢz!��,M�_���#�;uj���R�����C�2�<OC(/�� �~3Z�ep�`n9:ا���:� �� ��i���`�T>W����H����l~�eQ���*q������~�8��[��V�� ��T��,�W1��$�Q��`��l�;�&Ϊ?W:�y��_|�I��k�W�����"R.{���Щ�:��E5��+�2id��Y��f����9J��Z?M�H�,w�T�Ps%Ua�=����w�O:? @
�����96���0�<MZ/�$���'�Gx4F���w������x��ҁG�U{K��R���.V���yH��Y��s����J!kbφ^v�����3�����y�t~�aS����f��$\��`)�ܺlռ��@���b���%�cC�S��t���U��鍗�r_�3?��=Q�+�G�D��⾆�E��p���`b�T���4�]��G�l�W"���K/���]���B.�E��o�����Y�s��X�����(be�:>U�#`�@��U8�=���{S��F�瘊����CʸLI6���U�GYǢ��D�P��ظ4(���<e](u� '&~r%h8-�����B�^;�{^f ��tfA�24���^�I_��N4����y�R��,��=��)`�?��<�Y>Bw'�Yi�]]?�y^���1�
�.� �Ţ�Ti*Ԍ!�a3���MD���YɎ�	t;,f�n���h�6%u�`#0>փy#Y�%[��8z��-���i�S�)�$:���6��YAHXA^|�J#�·�( 2��W4���N�ou��V[�ƎhE����틦Ff���|��Җ���e���_�W:��^�+n����Vi�C�m*a{��|�擜���E�;�-�5�����;�$t�eUe/���ݪr���y%XcTjef�̅O�����w��������M9՘^�/�����|��e�9�\���jL��X��MD�w%�3N��o��Z����nԩ�X
h�͍��:pޔc7��O{JE7fߊ�&f&5y����d���W��x��z ��9)������2_��eW.�yG�a�-���Z��,R��0:{>rb�V��lh>��J*1Y�_�o�^eᡐ	M��"���ϸI�c��^#nLo�E�]7�m�̗��Av7�W!�Ѐ:�\�% ��8� �0�`Xҁųvej�m�����&��GL�
x��,�f
���v%��b�"dd�m�JI����P
� S�nH�D^�	Y���¬T48xH���Zr���+sS;���3����E��p�#�\j�6�9�[�������L���pF�U��P�:Nh�o�'�~���>�TO����w%AaG��Uz���<�N�c�]K�i��9b�h���?�EYYR,قEψ{��F�x�w^{KkW��ǄA���[?�uI�XO+���!����p`Ϻ*���>��[���\d�$|p����U����r��~�ᡦ��Gˎ��\�z����s����t��+F���Ȼ́�S$%��T�S9�?"�cI:gT�3�ɒ�0�����d�N,ֵsξ�E@�[�Q�U��S�g[����JI�(
��7߳C�Z⪩���~���/�$����*����i�RQ���;� ݩ�e��i��d��U�V�gjng$c����Y��x.�~�
�eW8��8�_��G��K�|J�E�tF5� ^k�6��.�������b���� ��)�K���7���OʿE�4�| l�����ɓ�"���k�?u_2�x~\���B�%{'�l_PF�����C2*%���EmU��{bWG��& � �������L��NYn�)p��d��������� �AX@���3M��>󕝖F.E��m6�ă��>�Y�����_O�!ᤜy5����g���S�:���3/���~��@Yι%���n	N�.��O�X�!3�G�1f��M����S�D��|g'����=@��É�P���*�a�B�SXy�E����tS��&9�����?��,�?�^d❆=2��  �}�R�<�Ю���r�2�+��q���1"�����J����ɛ��nm���ν��Md��ݣ���!U�_�;i��E��<93��&�!���X��B���s�GQ�)�oBW\�����x�\�ٶkv�M�8��^�
�ꄑ�n|
��'X9�~��d�V�cgU�MF��B/`u%���� #K��HG���w��""�:������yE����������.̛����Q=?�ʋE��f�.]��؂��u�-W�i��K>H��E�[_�3d���K��z欷p��˺����#\ӎ���^-ޠq��[���肕�K�+�ǘ�Jo�4���-��>n[�º6}vs腂yaK�H_������2���Y�?^I�����x�-�`/�-��y���Zq,l-���h+��XM�lO��ߪA\j����FN�5�n촾�_����y)Vד&����6�S�|�1�9��U�l�'Td��bA?.���?��E���z�iz���jK6����N>B����4.֞�}vvJ�g�yU�2l� ē��2~��Sn����%���o���뫽�+�h J2E{�bX��Il�p��A	�qqR�p�i��!�����.�ɲ�u���U����w���H��|�
}b�n����+b8&�c����6+��Ǌ�8�༺k�^���_�=����C�u��+��L��9�˫W������1��lߪ�ժcq�X�C�HI���������8C��n�c�e�F���ۋ�����2F6`�K�u�`��i�ȚԺb7�����'
qj�/��q�bHO䤪oM'�k�$U�A�0e<��B���F�<���IS%��bb�y������_*��e兛��)����E���e�U��'����К�X���+�Hq�w��?���߽7���ϕdP�Ut ���`���G鬖V�Y���L]�A�.�4�c6}�]̗>8�K��M#�N�O�BSH�ЯLĝ���!�^�6��=2��*I�'=�;ؙ��A{�t�y��J�o�@�?cf[��.V�������e:c����n��\��L�M���g�qpy[�3�s��>���t��Dh��s�D��Y;��+�ɂ�����w �V��n�'](��z��Zd�n������|������izf���+Nz?LfZ@n�S�(s(�,~�l�
�z�v:�>�À�MY���(#L����/0����lc�U��K`�I�6UG�iƷ�໸�%�Ge�
%�T�(x⃜�H������Ղ���,0)��}a��u�"�[[��".k�G]dB�QY��h���2
{�m�Uz��軘��c�tP�H�"�EEb���7(� �榰3X�K���?�$���_a�n`���2s��ɠź�s?$��u|�lьS�%e� �_m;����u��!�
L��l�#� |������r�l���8�.�{�1Mͽi�B�)�4\��ĳ����׿�>hGDk"T�V�}{� ���ƗFjr�.�f�%��O�c(��Jn�B@M�t~n��N뾫�m���ʟ}���k�4��*S�>����3 V�����@�_��]4�I|�K�u���%���C�G�\$�/#�t�M�sUQM
�V8t��@�������_x����h�8l����2������������]깫�iQ	�;��3.j�_�֟;8����L]����7�%��+���R�ǚ���UQ�VHq���:o,�j��/%�p�Ҙ����l(������f�BSo�ۓud�@|�#j��(Ѫ����]��
�_�8��r�N���0#?�W�Z^� r�v�^Y8z�4,�eLEQ���;=\��-�ӷ�
����Q�s�&��]ܯ��k����~�?�k6re��Q:�d�s1s])܈�dYTҨ�皴����ǲ���id�N��G!���J�����h^Fx�n�D�HSݴ�O�ٸ0�]���d��u��㎖�.`�`��<4�'���56Buv����� ��B�H�oq'3��o�vq�s���m
|���E�Qg7�ћ�R��;�؄���N�y�0k�$���/Z���?�c�H��x��p4�?ZU��Z_0y��n����Ʈ��x~���Ӑ�1����DFv������C�����M��f~.���9�b~�>������&U�94�@u`p:�S]��c�\�����w9�)j^@KPA�Ը-����,걓2���-���(k���q����o�"��!b~�[���P®�+��X��_�����	�MZ�P3�����i=>p9������
u���ȭ�xx�|/�a��t�{�<�	�hR
���l��M�7&i_���B��̼���r�)�.�n�*��[^�_R5�3cdu��,k�'*v�C��@���>���^<}�"�}T[���%���Ύ�N��\�`?s� ⸝N�&p�L�0?�&�}[��/�_�d��S%��(���(y��r�4�2�6�����G�1��[�ج%ήqY�(�sl .�� ��VL���=,:9>�2�ڧ����W{�X���Ԃ���V�����{3 �0�-� u,��U���9�ħO���K�ԩZ�ؔ:���S��Ã����f.ڔ�[�Y5���H���YX�󂆕��`��I^��&��&�y�����F�8U��s��ȩ4��ܮ̏��R�꣤Ǘ�h�a3�E�ƶ�k]�6A�S�n�Z��:�<S��C��pU�ƶ�W�GE�#�� �%
�yQ�ZWrfB�9���bAc���0�iz��ie�ھͶ/��K�Y	����a{6�^�����a���iԈŎ@�G?�6��҄J�։^���gZW�F�F���C�`�&�M�(���x
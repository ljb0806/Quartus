��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB���G ��[��ʩFF�8Q��*	W�C�V�MEEr�u�)u\4c_��_0��WW�"&�s�J�(9#�Q-�LZ�3�v� ���T������$�j5��QS�m/%٬Q���`M����Ř�'6�Ɖ����=��, C $
a�Pwi"�}߲�&(� �+m7�O�X^J�9d�}����U��.��"b��V��s+�b���v�It��8�EQ�F�9�`pU�?;����F���\���Z��4�1$�k�l/9;���*%��`��5D��j&m�b7Qu�k�����a8H���!9��)�!��f�/�M��%�*U���E�"�S�� V�3wJ:a!��պȃ�si%)p����7*:�5ӻv9�e
y�3��O$��4��>�i�m����]�m\�l 7폼P�o�7�Ȭ�3}���%����sCBn^0�s�.�L�S4ϔ�����X���y>8ў�4�� R�D�+����8�o�@kl�������	�����t�y��-��c��Rg�S^���	2���O��6�,�Bg+�7��i�����H.�]O2ʗ�x�4�u��f�e��A��H����Imգ�Ł��>��v[8������w�I�-�Vժ:FI��7�ƄT����{����G_�[�ѓT=�E�x��Q�_�H����Γ��A�Ʃ��OC?�,�&"ӑK��G� ��P��Ls�
��9ZXD�WI:U�[u��6H0Y���Q��zA�򄞓ȣ������G_2,���i�%b��Bm��ۄqUt�XbhI �LZ�"��cQM+����x	YZ�	+�7
{R��[�7�w��|�'�iLK�۬��κL�i��؃�=�7��SUM 8�j��T�=<:������1=���qy��oS�2��<�ř��7�h�]Sk�x�#m_˛h>��~���=]�8#�jW�ZB�ï�������N��(1#��Z�U�Z5O�2�����q�:���"����'��������aUwտ�* �mA̉e�]�Ƃ-u�#to���*L���V3eI�s���p@U׈���<�ʨGz5?�F�I���N���[jS�.p�w��9H�I!���	�Q��a��YFm�p���7�`9h.ErxcN����3���b��`z���,�Ҋ+�0ؼ��{�a�/_:�X��߳Pp�q��KA�#@�X��6�E�IQ�f֕4�������g��Z�:�~&^Y0�� �n���w>���&�l�f��vj�?��O���Xy`/p�ʗ��U�� 8_/X�n�1Bw����_�"�G���<�=�\ �Jk����FVċ�z�6���v��2�c����oB�o��h1�qj J�<�Լ�"�v��=��zi�˸��V���9��U�Sr�e��w\)��s���F�[��8��|�jx�)�c�I��>�ڏ{��0y;}�i���[�1���T��(���ZlvN��y�[9ȸ����F�^�V���i:������,��֟��B��3��~n~]�L4M���mk��p���Lo��v�*Sso �c>���v��%��HRO���(�\)�	�����AY�M�t�4:�V)��%��~���x�[�z%`���(6���ّ�i��t�"�I���S3iޫػuJՁk�/Qo���"P�'[���lp��ah�?￷�
�$z�%� ��p�[.R��c{���v�tx��x}	W�F��9��CG�N�/ft��`RK,�F����ٕ~�[��5Ev£�@;OM+��>(*ɶ�YRl.{�g�.��w��z�_ڥc��)���$�X��e��:�?��0s��X����s�e�
��^����u��ڬ�;�����#�u��@��gf����I�Ne*���(�>C�;�4���h�b�Y�U��l�⮮]R���@�H�;l*�3���jb�Q�_�Hra��hB�%�U�����_X�����b6+.���W�e���˴#�(�!�![�v��z����qz�3�Qa�z��o��7�ə�+.H�����G��οj�_ cu�dj��;��p�	c%�|w���x�W);�Hho4�}S&��'e�{�T�Ճy�;~z:�(�#qMp�ȪD�FHۙs�vn8�ٜ����}K��(]��$K�Ej%O�0��_�M��~�UC�h*�L��;�ېC+h����8�h�x�r�T��:Р�48��C��UU��Z}zj�|��B?}��T�%�����c�j�ק���� u�� ��^��ܪ&���B�<wZ,l�j�OWs��;oP��%�����2Bt�H����1�����߂�j����f�6a3a�"���,��m-�g\"�Գ;o_3AW�����?6�[ ��B4�rl�R~!3�S���{ ���X��x�`&[�`c�:�0N:t$}��9��+g՞[3�x^�J�J�V3���n4���l����7f�����ѥ�����
���k��8|�_�N��n��yz�-�����<�R���a*�p�ce��x��F�:|Va�o�"���$�4鄴/́a ��	�kl�̔gƠ{��xċ�T�s|_���"�O5��n<}��[�RW��V.M=QsoIŤ�E4q\:M������ٻ�� ~3��_�� �q��FӾ��9��k�5֏-QB>L�?��q_y��45n ̏���CUs��~���067$V��[�<P��xi�ЕO��{۹�<��K� ��AʭlƄ��%�{Y����Z�P9�4pE9z�.�Ľ@{�\�@����W��U�֦+��Z�Q���R���_������$�U��q��z3"A��J����P֬'����=xѡ����b=1s��XK���>8���	,��,c��Axy�M����hip����U8_������f�L�nJ��S�VhD���@5;�f/�a.2�d�{�����������0��!��c�M]9m⽤�&x����G~�[S��F������\A�����W���!�q��v5��|MGO�HDjqpܰ��5��Iw�ʰ��~�:�[ظ��t#�ߦ\�u�� Js��yX��
"�����Dx��Y��g��ǙÊU\o`v<�ݑ�˄�i8��G��g��j�f�F�Ӎ@� %Q� <�٬y����H��Y|��3�e\:��z� X�Y̆�Ѡ��ʿWN�H*���	�Qc�J���˜����ᝨ��Zj���d��ala��Ks��"�	����Љ��nhf��
���V���߃���,ɭn�E��!8�{��!�6RT�,��g���Ȉ��(D�$TII��B��N� 3G �E1q���<���������lW�fxƳjp�jk@��,���q�������5N�3?�g���+' ��]}�6�B���6�?���La�m)�v���rMQ�;�W���D�%�=cInǤ��bj4���[��̸�8
"C��>�,ζH����k�����_2�>���<* G6d������
�J��8"��U��HV*MFn�C�L v�z����*�x��#S]]k0H*�]�3+���3����k����u�F��kt�+}�+k��
��7���w��.&�:a^[�^����n��R.Ŕ�L��?�JS����2<���p=�{�I�ae���n�o0���4>�By1�;��{�w����f���Z���Wn=�3]>�}�7}\"/���f��x�+>����<1pu�Q�/d{��V�xCQry�,P1�}��I��-U�Y&G`8j��A(�< ����7~�<Wdq�p���x :I��YJ̔���G!�]�q���vX/���ߣ���5L�  �(G���g4O��ٷ)����X�������4�݃]\�M�r��~ɵ���C��<�GG$����;�s�ou�,DCF�Wc�٭=�݁�V���.��?�]a��1�� ��� �����6��^b���<29��@�fbhO%�1´_T��~����O�������=k16������rO�����{]��<�3
��cM��U�-�'e�8=�yzEW��rB�[y���"7�[,��;�Z�r)\�@]�~:5+���%���W>����^��%ඊ�`�IZO-vV��x�e<�� Ė�̻*�l��5P}��̳g=���Ȅ�	7>-�k�˘��cXM�t�k�W�����ِhO~wl�Kr6֗v�٣
8$˅p|��`C�L�ü�K?�6�#MR~����6)a_����4�8����T�%#�R�Qpd��Bf�]���J���J�g��(s`;uS��T
�P!��\�!��+᱙�y���DG\5�Ĭ��T��n_z��ֈd%�[A�LFw@�	K*3��N�[-�)���c����U+�1���R��s�������{�\2���>Ò�ӂs��N�u�(���}�]Ӵ���U��	C� >�xQ���F��-R���J#�=>����$����um�S=�pDٮ�TLOY�-<C�T�F=�����\ܐ�ѫ�ݑ����R�ʘ�5b?����
%$�`T�9A��V��/�e3�t�;T��@����GV!"�%��gZ����2q�����Y�9$�%��ߟ��K�={/Qj+���S��b�)/�4�f���xwV)�sk�5�M��..��R�f���oۛj�>0����'�Oܳ���gn��F6�:'��Z�g�AKEQ�DV���˴._��v_'C��n�L/K��*�*�^��^c�4i��)7���|N'��a��m���HIItc�V@�2-x3R�¼�XL4T�B*q��Lѝ ��x�p�X�n#(W��9f63���˾���hO'�7
@T'�P΃�$��k�%�o�I�g�,b����;|Х`�O��.�5��>����dp�ny��Ѓ!�D�SǷ��!P|��;Ʈk��uw���T�{@��r]p�3���;�@��)۠{D/��Ѐr�X�Sl����U[��
6��a������%-R�4��Z��=�EڛC>��?A�]����{N�MoĤ�I��s�#����Bfz'�l�X����,E$OgYǩܼnh��ݼ�O>�>z,��v���o���f�D�M�X``��d������@X�O�� }�2:*C�I51�v,4�G��<c�A�}
y�ESe��L-ڄ�/����-�d:*��e[F>d�����n���Q! ��]MN)�J�M�����N^|0�0�\��nQDc0�ُ�J��9�2Y[:�HZ��}�3�T+.�&&#��h{��-�{�%_��U���:̻�i˴��Մ��*PE�/%ΐ��a�y���G�����/؛���A5 �e��=��"2t�i2y���|`�wh*�M�+([|#��[��l�[T�)~Ɓ��]���1:�"A��i}|b���������Ot��H�\>/��KϦGw���UM�h%/F�CX3�5�O,p��x]~$5�u�/Ig�L���`�7ʻ�Yc)}��d�.�[�i�D�8�:��c�k�4
�d`��>��p���f4~�]^��0��_�o�huc7�Xv+���Zv���3�`3GF����y�r �GXϤ͂�T}�s4��/��T c&:5�[���N����]��g��ް:O4W2@��;�N]@;C����ɽ ,��`&����̼����.}��φ 3.W�K9kOz���ҒҺ��I�}~�J�Q����Rp�"O�7���x��U�H���(��z���F�[��ἂ����{�x7#�ěE�����E��.:������6jp�ӜI��Q��%K$��bM|5:(����:��&AY��ۧ��S�����rl:}䙊��d���S�4g'09{��o�[^�O���ZW�%�P���rFk冨M��G��pC�X��`Tau�X?N%H�MDI�O�Ls��%��py'�R�(W3�����̝���U$2	�$�ވԠ�t/�a��7?�U��I7EV����>T=ț�14bϟ�m�u���nD��>lx5o���xX�R}��I��3?u�BǇ��^j��K�{*�7�N�?��eg|;��dsS%�@bl"f&Mgv~n��~�_���_W86�p%^:�N��I1�c�C���H�
M�G;G|mʋ����'�1)��h1�&Y��3��l~x-��2���{ 1%*����|�f!����063Lg�hǠ�NW����&�f`*�λ��i�5������3����se�����O�[���S�.<������"���O��Y{��t����]f�k�#�'�Crr��A��a@���;O6 �d�'}���R�53�9,4�}��S)*���G+ ��V�.\ʛlFf�d��xl�P���/NQ�ĕ>Շ�z����*�ΙSoʀr�P�Έ�
�i�ƕL�Tލ�7��͚�Y`J��pئ�L��`s;�en �3���w��t�C��,�ٳ��l� ^��?���J7��G��3MP�o��V��M���iEG�ICZH6�T�r�U(�q���_(*]�x�+T��Y��L�68�,�T�3IHq	Ýg�-���w�/~��t�#��~�-^��Uɧ�����p�3�'�������׸����>:���m�1r8xuļ>��H˯�G�܆�h1Yi�U�4�B6[1t�������㷳g�D�/���S�*Ӱ !%nΚ��Hs�  �C,T�����TЭv�Bi3okr!Iݬ&�<!��f(<g� �z������[|J������h�8���G�]�آ�Cq��t_�� p�}�"'h��߂��ߦa_�-m��!t��+.�4ql}�#Bt���d�^����
���ˑ�˨�O�ݨ+��5&0��l�Z��S�d`ʌ9��c�C���sF�I������?�p2��s��Q�|6�֕&�i�V[.�u��0�$��=���"e�L���~Ԣ���MC���k��Ŧ�e�mWݷZ��!�.���,qx!v�h��l�r�ٞ�h�2/���e'1�}!
�c������
V���i>_��F�NE�h���=�B�$��������\�*&�W^Ӑu�skc��8��B��HGy8])�-��	���g�$�t=>M�;J}֏Z��"��ܦ̀���e֠�B�#e����k%��?���N�n3%�4=Ͱ�_���r��
�-�U��}s6Y�a����V�}��;��H\�+p`���t_Lf
 �D\U:�NĲ�sk��mة�@?sy_�4�d*3����ZA�n�/�Y�UdF�Q�Ϭ���� ��>�ܔ�3C6E}|F����	��S���sj6'�i���qq��7i��$Q�pCu��៚W�d��Q�E���	�[1�Z���S��0�����	9r����+�y���;����͊H}j� �}�b4u�S�{}KH��t��U��'��<�'�j s�q�ГX��GEF7Z���3;�R��A ��RD��A��O�)��&���m��`��GT��Z�����\^��8V��`�Lj'���It=�ֽQ�V���b�p�%�ȈD�j��hP'��
��� ����h�P�b���ˑ�P�M����v�f�*;ThYOS�9:��P���k�:��_�)��{�U��|��.�-�|+X�VE��̥t��|����H��,ce�i_kKy����M��l����
�"���|�!�gxU��$��3��%�+�����㨩#�6��Vr��ך��p��/���)�
utIHVv�ѧx�n,~�P�^c�!�����Oφ��z�����z��W�o���C��U���qZг�Ón�O5�(����!��\��ۏ��Ȃ�0�������{�R,�.���t��{"�����*�M����� �n߂�G&~^�­�+�ν�l �am:��7~e$�M�-@�}�Z]F
z�T����G�j�z(��quG��ͫ|�%X���olq������wIoO��)Xi�`����d�L�w�ܴ%��U+G�֐�Ʉ���u��uY��M4p�kP�Rkt�-;vG���<хh<ɸ�v�n�I�!7C�@��Óo؋�]u��w�XZ��.-�U�_��3}�?�]�����_ڨrbl����ZWļ�@��:[�O��`j���&�p��k�C��g<��dDCX�K+��Ye@��%J���2���-��g���3+��և!d�gy�FA��]f��8�
-��z�u.���]�[�,<�DK���
����$�Ε�82���a�b��d�� �7�S��!�`�*�t��*F�,�(?7Co�uF�r	��c��E'"0��0��u.DT��E�=���׼� d��?��7��d�K�ã���;�WËЋ08Q�� T)0eF��w��$�/���`%��P��xr3�!v8{�C�k`��45�򊿾�Ns	�<�����`|T��׾�Z����.�y�������q+TO}�Ĭ���{-��`����кa��;�Yg�U��ps.B��YV����Ҹm��;� �������c��-���c��H��¸����&u�H��W�����5��i�6��D�����w*�/V<?���5���`UZH{���;��NQ��_N�ޝ&�N?��h��/��:f��Ƽ��U���"�ڭ�w;���i%���|���nA�>�@�ܛ��;$�#/Y}+�aC���:Ƴ��5dL���7�����^������Hi���P*٤{a��<�c��Z���BK;J�T�oP�k@d����R�lKB�{3=iOq�.�.�U鵡�*��o�D
Ȭ<.Ӷ� ���Q��ʐ�;Y{�2o쓕LG�����]�6 ��6�*8%F��!~���
����V�����+���t�13�llx-6�a���ٽxI*�6�ӑ48� ��BR��%
)�:تi��%�?�����L)�ȿ"�90:�@0\i;�$�w�
����^�5�!��ߟ\}�0	��	]�
�ר�#��|���i��fʋ�@�L9�=L$����� �F;��o��'��q���(@6y��}�������J��;��k��%4�Ү�4jy�� �W돡�O�*jT�c.J�Kk��O��㫭��7�9��2�k��")�;rb��H
�7YP�+X��A�_��6ϫ���<��n�����j�͓��U���{�pE�.��g73��8%P��6���/Cge!����A���HL67�Zr��j�{Ka$+"*z󎙜��%��BD<X鈔�Z8��=A�7�i��P�gz�]T!qV\yӔ#���o�η��<�aY���9�����'�$T�T��sA��h�m���/h�e�Yϐ/Y��4A��%2��T��9���[�)C�����Aw@U��T�mty	@�	u��Z��~�
2<*�n~L�E�cj���e��~**�����e��'��%��G"��!b �	-���ůuA����mH�h�۹ �Y��m��*t]T��L�b�X����6�V�r����$�{��mEzGY�^��A��@g�͋�;	/_��(�����Rl���D�2�J�/U���1oY��c����ڥ�s8�����OTgJBvB����b��ja���m'��iq� ��Vj�-��o��0������%��4�mS����A��Ϟ���Μ��DwX��3��#�D*p$9�?F"��xi{���I�6�
`+���r}V�P6C�tE_�k�k0��&mg��X�;n�?Օf�� )+���]�b�P��i�?X��b|��D���zf���A�qf^X�<���|�a�^�uZ�P���E�S���ԥw������>�G�C�Qy�����3���z�S!��N݆AMoʼ�P�H�.��r��"�6-�K�p�=�a+V�RL@�X��4�d��e��t�@�p�W��u3!M�[J���o�����1b.�A�ҥ*b�=��-7�D*/IA�sz�ep&�4�#���hT���Z������$�zxu�D@Ww�+��雷C�G�&�T:#�y���s�bL��u�f�4ј� \� 3���W���e+�i
�r�?o|�-6����w��C`A�6� a�+(��_pYمX��-��&	(V�Rf7��1t���9���7p��!h9V;:��,-��B��/G�/~�.��y8�����{��������y�?�8�����Z�>��.&왗�ވ}���r�3^r)����������,�Q!my�]�a��ٟ��Ru�PD�c��-���d�:��)�t�K�����%`}�w|��m�%���0���$4�����5HD�2ϧc�p\Q_�����?������c��z��O��f�����:0�͵>WM3x�Da-�LHMẐhaM�2�Ő ���p4J��/����V��H	+�p��p�3z���x�0WŲ�'#��,�Gv$$.�%�_Z��8�s��r�?�?�zcE�8 ���j��O����_���s�W-�̷-yh�P/�i�:̂�r�\�L �6=�� s�s"�r��b���C
Kwڒ��!9u73W�l�рTdx/?��`�e�W�Wz�F�h䡱��ٖ�
`�	��c����E �mk���Ф�,2�s��kn�G����j.�lti
�&�LK�W���cI�;�x����WD����Jet���>c"Ex!�!��:�Bh:R09S��VĐE^��V_
�d�!h�cx^����0��$9�4G�����9��l��l���5(�&�f���J�^�|ڮ�#�8�U��d�s;뱼��+<��zx����D{g�`](x�j�<�`CVA���W4�a��=5eY?c�����b��QX�����\R�3�[����.>�-�)���c:�z�������*�Z��#�>/5�u�Tc���u���H�� �9�nL�ّ�(aGK!&�E}���r�G�}�
]�m���1T�[�Y&����Jj��熂�7�cu��C�@�}�S��ZMc&��e$f�1��g�{pu�]�5���g�"��E*����mt�1y8|[pxt/���Q8_	fRwm�Hk V��4�A�%���o,_��j,�������Gd3��:��C_�e���0Sm�l�{��,�ڐ��L�R�!����gg7��*��3a�
��r�:L��o����:�p�z`3�3+��#H����R&8~�t�e�Ps����Y�j��N����fm�5�)�M�{�ҙY\��
^j��)�wn7W�1�k8�̛P�S�]0�����"��"����f8�AI:�����f�K|�&�GTDe9+�>�E	=׉$�?i�$	0<F֋PC����ȸN�U�@Si	zO_�^t���R�J���u�1�}Ɛbf���
rؒ^h�+DoˮҬ,�G��K��q����:ۙȆjN?��Ak���vO˞s{MIm5l���n���2�Kg���w�M��=2-'n�_fV���\d���X�نO��r�i�Щ����ϩ�jv�H�]J��{�_{P
U��"ƭM���"ش�c�tf�vgk�Y5W���$�
���>_YJR)�� ]����zq�c�SEv�#��U@.?qJ܏��|��"�{���C��$�i��u���f�oAo_G�$��rI���]��yI8Õ�����$�86�v�cL�U��EAX.��Ӆ�
��� �ľh���ZdE֡���M�eq��H�&'���@o�(���n�CLCE5�x{�n�
o��T����γ���Q����iXl؋'w����Pr�C! ͎C�$�w��:�MM���Uc֣���2�[��UH{>�J�ʅ����_�>n��x}i�NB1�i��)u;�m��G�e����g%�!~��L/��-yOAV�ϋ斃R����s��d�; �f��껶�Q�*�S�	��2�r�%E��qk��P��cX����L`YpxǷ �/�� 6��K!L�ơ��Ё��C���EQ9(�!;*�Q�����J"w���ב�X����t����O}oz���b�Y�xO)e�t��C܀X!�B�v4/�p}_�]��R��j�u4��+���//�sxU����6&]�b�V]�=o��b�zm����[3	E�Сs���Hb��}��@"����^��*�ۜ:*��@��W�>E�ل
n��Wo�8�+�]G����!Ě�R��Q�e�%�RM]Q`�J\��4Nz���6��� <W�Q6�4Zb|=��'VqIKB�� �k�LD(Z�ٻMl�e���f��6[�J�>c���huńBd�����{��cc_�H<qǧ�Z)��H���`U����/ "s��ڽ踝ɡZ��#|W��s{\a�l����-��
pՉTB)u��9��<%g���ftL�4?�H�� �o���W:��ӷ��l����(S�)=����Ђ�+��˖�V҈O��!gA�d$	�pƀ�jB�S7��3>����I�֐����B�k��v����K
�P[���$�Dl�(R@E�SU羆/ȃSjf�����V1q�x�3�F,�;�ȭp�������mq�Ќ�o���Y�O�B�S�o�	N�9���&cS��!�ݪj�'�sCM�����@�O	Ҟ�(��.c9*����\��Z�~q~ �=7l\Co^��r%t�u��Fh���Ռē�p젝�!ʽ0��_��-3P�Km{si}r+B�0�0��4���c@Yn_,�1��?�j�]@G����Ol�������ӌ��"��P�[zk~�H��Ｈqpx�z<�1��{1|���vƛ|��T ��K+��e���Q�У�O:�t�*k���n�/݉��ݛ0��{�&�v�=>�s�o�ܞ�j{�D�5�P�.�VϏ��T��Y�;�%;!�^40d�91�+��EA�{��h���x��FT~��Z'�\+*'r�1������2�9,�� 'K�M���Ş��.2P�׈+z�[�!�U�{�����l/jQ�J��8��ls�xu0�`�'w���5ݡ@���4��u&��e�D�ۦ"�G��n��P��7��]���Eq:��ƌ{�K���|O����y~��?��]��j�&�n�ϯr�_��������a	w�B5"���Q�$���.��DQ#I6�)�=��}sq�j~�4r��� �;甛��}#�M
 �����9��i�����h����wAs9@�_���3��C�����]Jsv�^ɲ��2`Z�%w�`H���.�-�Y����o��]�y�v���X+Y9`aw�� � '0�	()�1�2�N��w3���`��浼�d%�7�X��
�2%XrMmٸ����=g͞����__���1�1��]C��=��ȉ>�*��q��k�0�K��]�iY�$�&�9msrjôy%{��xP�8��w+՚��:u ��e�
�!�fX���V���}�b<[��K��x�B�'	!�����h�L���3�f\'(x�Lh�!�5$��П�N��9�k�q��1J\�~{�9s$����C���?~5�mH�9���y2�}��V�V��i�d�*�D�2�841��P�a�����T*�e��nN<`���fe��@����{�5!=K����4�ܑ�*��e
"5}6}�j{ǦۏJ����������a��w'��?��L���
�([�=���p�����q[���+���k�o�O�]����dC��|��2)�
��<U�$p�n|th!��8�$P��"����G:�Agj[|/BU=��OM):�-��(������<���o�1(�U^�pXmD)��u����%MRk����Κ�Ǆ��޳@o�<�5��|�I%�@������+
�/���/�H�e`MK�;�b�_��Mq�͕�:�����Y?;1����薪b;�	�goB����Ot�?���)Q%8ݦ��XlEm?��w��k��O2.7��E�|�g���$H�_��Pw's7��=�}<HY�j��m;����[R�q��,��r���ee(�~��w���xu�~���җP�	X�2^�9&R��|��t��~aV�8k�x����	;��2�R�QP!��_Ń�ш|�I��7���O�����e�d������Q6?G��j������]ұ�^e��G*W6|�S�z\Z5Y�]���bZg`�Bl8�I�ͣ��"��'%�6�r7B�יY��E
�SEr�� !�;"u�|*I��L~D��[ [nF3v��D2��K�v��O�>Ej�.��Ky��ҙy�����S��^?��VQp������lH�B�n�N$����]Brx8����/�.<�� �dyY�҇����YHW��!�"��fF�nT�Z���rf{F�1г�j���*�1��Ī�҇]u�<v��<��ƹ������[ђ����>�Z~:�IdYc��?�(7�k�aB����:A7�L2!'��Vq��#��ծDY��3�&B5x����?��=&�G��� ��@�a��N�S`��BV��t����\8|:�f��[�!I�AT$�`��b��~�e��*�cϢ7���]�9fWi �_%���Q��͓�N �;��5�Տ��?��s7���x�Oq
^�1ꄳoQ���:�J��a���ς��w`B`B8�*�s� ��շdf|	e�ynWu�����Ěo~U�YAs�<����S�J*!�5�_3������t�鍬V���R����)Z��P�oTJ�sh+��1R��
����8��|A����q���݆$Z�J�ie�� ���8��O����mL(>�=�Q�Z 	N�{����
K�8ߎ�jD�9�d�_B�w�μH[e��M�I��~c���rI,�S*�
�|釞��b~�\��չ(�[0�Sc�>Y�j�D1��YR��[���C����������CI��k�����~w�>�6�<sX��`Q��{U|͕��ÝI5��TM�@��i���_�ֺ:�W)���?k<���[�5�d����b2��Z;	�5��jlRK�r�v����XO��������X�+P7���i���,�����FU�b}����t�.%���܄����&+8��|�������j�2��[jpi�.�IhƠ"�
{=zp��$��+�=Ȱ���t�|�]w>밉�1Թ��� �Q�����:4C�����2���� [: e��}�n���yĸ.�j+�w�?�+��(� �B�}��a�k�@�BZ���R�Íبé�Y�q�J���*'�^Q�8�X�\y�6uK/�6�8����Tut_y|������4��}  ��O�ٓV[ X��h�1�{��6-�j�/�VK�G���;A�LV�u����!�^�=bl
��n"�:h�����/;�!� ���
U����j<�Ȟ�r�����{����p�W��.<�8�h�Jww������9j؍?T�{�]������$�\��`?�6r�F|�/�o)�@|z=�.N��GM���-�&�Y�?��u���{��*��Ϡ������dl��"V/��U�ʲdF.Iڈ�� =KZe�+�3������r��t)���Wd-�7�ig��LE����Qp���`C�>⓹ׁi�qF�-#F���ВM��K,UX����x��Pj�@[(���	��i�M���ȩ�e6��x��<�:n������&'�q�>��`52�+�YD\8��qdNF=6Z��q$����ݪ(��c��zK$�U7�v�t��X�}����.�$�����*�5���2��@��ꭷ��ڢ�6=N��3H��I	���H(|�Y���a�f�i|�zK�!(�h��>Ly��߲ W�`0+�َ���neG�h=,��-�@	�� s�����ʊ���ZT�7- 7�f���T����%���G,��(;�Oc^D茚���OG��_c�0���)�G�XG�����d/,)e�m�-P��NH���Gޣ��@JH���	A�����b]}�	K��+A�(&��V�Y���ג�B(�6L�(�<�"9�0��_m��W$LJ̃�H ��فӁ��^��,	�Py$W�VL�\ܪ�]Iw��� |�]�����r�x�|�D��"�u�A��q2��Ɇ�Q��2 �Ā<rq7["�F�fs�� ����գ���s���p�bg���Rյ�����X'���J���e�-�
1�߅Q��+ǘmPG�Xz9�tޓആd��:��'ѯB.�j�����c�͊����4�y���.>�!�ͨM4��#���uO[� z�+0�6ԾX����Ob�����6�Yw��b+��!�_�Õ��*��"�1Ԇd1������Ͻ�H2$}Zٗ�m�����X���Wh9���ĭ�&��Q:-��e3����ht\��]	�L,M邂JA`��L�q�����u[<���i��Ѩ#L�D��( ����_���]��x�x��{r���܂�p
��z�B�8�w��e��M)4/��G�I��E�>x�v�T�F$�pH�W��K���F;��]p(�a���*"P���ޏ�(��
��PJ�Dj  ¨*«�XdG5�@�./V�JjH��P�L�ۉGFͰ{D��|(a���Y����F�sR��]��3��S$E�B���L����x�`�&�6�,�$:~�B�`0"�����5>�ّ&g.7��с0j��.���Bʌ<�^�N!G͘H1d7�>�O��5����U���\4NzPiG�d�[��Gv|
�j����\�öj���U�l�ٕ �"+lEԪ=@͍'<`�!�2��uZ���7�mbg�z��"�K	N�,ǧ�� $�2uw+K(=�G���Z��+�唭�=V%%�0�/	[%�![u'*��j?�L�Ł`Oz��r�K��]�$F��17I��\�;�>��P*=1 ����2��+w�\��KیF�@��&�����&�Tb�
�n+�҃:�ź�'��0�CaB�F�
R�s�c��»s~-,�_�I�|�����C��]c�<9����H`��F�F�wQ,�Lb�\g�x�/�2��]�i�ֽ�p(�4�P��fpW6L�4薧�z�4|���4�=��w9�q�Ar��QAV3W�Fi�5�HL]�ޚR�I8��X�[��6���݈���/�!���!�À����_L翫S�f$�g�#�ϯ쥷��?��D0��K'HJQ�,N���,x�DBX�'�i+G?8�(7?C-�H�d���J��l�d7JҚ�^��t�?YQ[�'��#l;�E����v�]4q��5[�X��0�@e�'-Е�,)G.L➶�W�x�ݬT�Ԡ3M���ٴ ��CB!c{����u�aym�D��Ϩmi��-e� {Dύ!�[��%pzj)XI��o���r���s+liJ�z�'(��F5��h(�!�u��Q���O�������$:�G�:�@�CX.	�9���Jq)�@�>���7Z��w����$	�vv��~�R�@�
�*v�[&w�,B5�0X����?1���tG��B��K0�/�3�n�������>�?�^��J*���T2a޺���ܣQ��+�i���"�,�Ey�T�7�ohBt�) TQc2�� �I�]�"�r����m��߯�m�����^BQ�-�ێ�Vw��t�K���Yc�m��s�M�*�z�ByR���0;�D���#Bׂ���;e�*@u!!V��Q����Z�>�d����1�c^���(����j�(�c V��)فg� ���#��x���_�+N�9���s#��^����f�U����9P.߽�����%p~Wg\�E���j�/�B0}�_: ����b� �j�Q���#	 � }^�X�i[P�01_9��<w����T�!� K�z�1��W��"`��p�ۅ�hqs���ݫX�FZ��Si��-�\���|��� ATa���Ι��͙�ћ�4�^�^�c�$2)��#���e�iX{�9����j��C���Ӓ��S��E��i�s�mz�miz���x����"�T ��؆�Q�I�ӍZ�8��H�r?}���C6拝t4<H���	��*���T�ui�����Uě
��;9!�����7/h-U�/�"�7��ъu��������m��mR� �"�!1sF�)?��x=�D����ˢ($E�@�k���O���~7��^'eLK
W	k}A/ƚ�?rpG��Pm���T�:�w\����㋥�*!P�ۮ��W�@�=޼������(p�4�����q1��ٔ<a���� �Uw#ļ;��!!�l��f�`�6�UR��J�������d:�,M�.C�N�IZ�ˁ
FA ǵ�I�~�z���T��֍F/��r�M�`������b�lF5Ι�TJ Ǥ�'b���A�RM�|f�m�������'��g�Qci�2 H��.K�9�zH ��P ��;!�.�,e��z�P�熪N�<U�O�v }p+�9��a�v(8�T���ow�.(�Ѱ�x$N���h�b1u5R��2�)���x��֔����4=�X��+�~�v?	���S�DA�k]^Jވ�����ƺ�#n�v�6�JΤ�B�m`0>���'F*�:����B�ď�
 ?�,svD�h��k��3⡱����?%Vc���-MzFȟ�y�:U����p�0E��s�C�e���D�m �D���yL<��[�Y+y�*����Xp8mN��jb�ĎF
���{����x��I����!&�(|�}g�)��g�S�Z�a��䕓�%n�JlPA�ۧ���I��wino�WO�5�|����h�7i�4f&0�^��b����w��L'��9ѡR�-�=���dv��^g�4�#�)��GS̔�!�V�Zm�;qϸ=��&I���N��S<Zw.��C�t[�S[i�xY0z����rrZ�f���}I	敚~�:�GX����&��j)8v@���%� ia^��	xT)�LN�\����E{�ΪP�(��S���8T*��$��`��!��H�������w��͈Aeπ:�;�+�W5j'�:R���>�n���	t��m�:�q��\0��]5:M�zy�5b���k�Z�{���7�ɶ��%��$)��<%P�k�z�-o��ʣ��'o%��9 {p�f;����ύ�7M\=>htT4<��	ɏ
��wC�ޘn?�.����ɏ������Ú>����ܠ����\����%�����K=�c��J<���?���rZY��'�L���9)4�mߙ��<���|>�l�O6������/rd s
j ��x���	/��bz[Ab��h������Q?�E��q��kEi��ǵ�3���Q�;o��H��4�qJ�`;JމF' �8&O0˧}�~.�)��`6_w�ނ��QX�����l?��J�w��������7M|(�����a�;��q�<_�4���hK����.\�p�[�7��\��t�N-|A=���2S�V��漐�}<��ԏ�*f��{e��UF�����x�%��͙��oS%��� (���gټ��i	�� hm���e4���]�p��9i9Ϋ���!�,���\��wE���$Tꔲ$=�[O�8eo1)_B�J�q��
5��z�9���=lh�*`3�Cb"�ٕ[����C�A�7H"����8�m��!��β���>a���mɸ��M��2UMe�LVoN�,X�Y�CE4
l��^V�a��[O9�l-*�V<�����_`�vC�Mk�%�y͆�к.�
�w�>�~�ì����Þ��y�R�ɗ�	q��pӦ�I?ۗ�A�
�����L�Kpo���$��
t�����g9	�f�x�Ť�
Ci�@*b{_3����=ߒf�so���X�S���"L]����q��Ϊ�f�ޫ1�bc�%IÎ�~�W��ڭ����������]WW��Vv~*��$T�nb��pV�;ݪk"o�H��E�)�4���ĬT����e^y��0pJ�j̙���iٵdu���?�{��Y���oA"Ý��I	+(�@��yi�MYtp�ٻ�RE�Z�N��J�S5�3jԕ��q�\#�>�xQy�JL����k�@b�*�K��#�����~&��,Y�C���e���t�:Q9�V����j�vچ��o%��JO$���[�@^��K85�mV�Z6���j�FR4,W���DA�X��!τ��Q	<Fg���E�q�	a�0�-�j�2���8l��U��ɘ�.{Ib�	���?�l�ZKL��~�
��y��?F��mz�!���෰p�O���l�)��������շ�&�͢]�ټ���v�\��dvOXB�vQ�~�N��ߌ�
��2�bQ5������z-��f#��;i���ܵ�:��'�(�ˬ�[��!��L��cJx=ȫ�����ܣH�bK.��Hj�R,w�]�n6-di���j �)��gدݥ͇��C�YN�S�����!-#J���&�6�Z{�i@�� ��b��L�R:/�/�6���(26@��A�����b)τ��$O/�a��E��{VѾ�Iُ�[���{DP�H������8@�e�H�~Es��M��C��z]�����?R�W;S�)�[�j��7�%�'�Y�o�Қ�yj����F3@�������E�������D�dV�l�f�ҹ�κ��W!�F�tT$�ӆ-�'��
Q��mV_��I ��Q�"�E�� �;��a\.M`����i~��6�a�li�޻��|���D�S��� �j���9zmlٜ}藽	(
i4xod�\�{�f+�Ϳ�܈�E�n�$�,�� �趷S�uD�N6���7�K�>ky�do���8]�7',r�{{*6K�ЗF=$��3�H[��u_�����u	���5%�kB�f𼵵����Y��n=��+��iy�U�\p�$�}��0��3^�j�x*��^�tC0�o�F��k�k-DTϕ-�d�?�
	�����11��C�{$��	��{����6�@��. �U�lJ�O[�W���?Rwkos�Bf�ݷ��K�R�J	��b�yvh:	'�����W��h�/��>��̦>�9D�C�JP{�a�x$df�P ����#�Kf�D�ZP�0��A@�ր(�����'G�7��Y����ʰ��6�|}��>�]���)jX޾���2髿~�~�(�"5$�$u�G�)%�q5)�3�i`a�m5�`�doN�:����I� �����^�b�Bב@��p����qL�6�L��E✔(�i[�)'�5~�0c���Z��'��:��1�w��d�ɬ�8C��|1a�t'J��4����������e0N���k��}�u�\/�zA�����
�u("~79��r^��`B㛫������ǔ_���"Q�*��2�w�-L�U^�lf-��T��\鸹�ι�-8�bݛ����K8Ki{}�%���U��9���sr���|���?j��Lz���E��K��GD
����.�OU�2λ��}k]Cf.��J��������pTi�%����[	���YM4eD����aR���r��f���n�a߄�>����E���[Yx���,����WF���V� wO��΂�Z�b�KN"�����2Ӧ�^w0��$�e�4�x�~2�&:��!&�܁�g��H2����j^�	�F�z1����[2v O`~�\�y�O���Ö��#I	b����c���A�b:]�����kD�g�(>~L�H]ě�(��z�7O!�bB��[t�\��_�s�Z�6�>�g��;;�/Z��)�&��`�G5����3䃴������B����9�o�(!́3ص�a|���;�p
�kb���S�2]�^��M�ڧ?Ȼ���	�88��p-�=:`����V��s����B�"V�6o �.n�%S���x��f�m�B��!SB�.��+,k�Է@>��M����*:Hw����)��ͅ�.x�&E�����\�s  ����i�	=q��P����*��T���"�����v����2R�Qv,Ӥ���5@�+#HIJ�+�YR]��y�*V�9N�>*�sX��T�,�A
ԫ�r<��u}Dse�1�e()� ���Pg�+�[��<!F��bv��96��@7�
�CO=�)F�rP��}6�����%3����m"n��2���-�Oվ7�`�����	yC�|��h�ަ�aFo�s�f[��s�uY��V=<��z
z�s&E�bH�b��HA�e�M�U���*����7��9��C��CԦ�4C���2�p���㦟��n��a�Js��B��b�2Xr< ͦ�r�Cz�0��Qu�7���1W�0�l�"�9m�9�6M57�G�\�����F��|x��ZY����fH ��E�9�
;���gF��+�S�%W~�m	ob���k�;he�[(����n���j�_��+˂V�A�᛹
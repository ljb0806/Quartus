��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB����]U~�_u}��
3��7q{k�m��s�Q0�Q�3�iԮh��!.Bk�|�N�j瑥��9E#\�T�Jxt��dm��w�+w�_��<�Ǝ|��ֱۘi{�A��9��>��U��w��E������cB}x�o�+�6�n�G��"�ӕ�R������ĭFK���[�ږ�Mǔ$'�����yd���{��W�-�a��D�{�"���ٛ��P��]����O�Ӝ�>�� �SO�P�$X�@�H�)p���`��+�i;U��O'����o��dԢ�m%̃5���G���V�����D|U�6AMir�橦�0Yh�"�Y
pFj��<����U���W��ܕZ�.��B�;<n�E��4|�_�Q�,����cms*z�K�%`>�G*%D*=�W�����ɐ,ܓ����;�@�/7���Z�TqS�Fm�Ɲ���^�E��Q�����)��^;�Nn�@�3�׋�[���a^�C��ωZ�����ۥ��&V+�lKq�
YR�`G��;+�4d����S<c���7�i�1og�YW�VEwgZ�%��2�)�\��w`���`�]�g�?�:�>kD��F�l��\?r^�t��(8�����+燲��tj:-�9�,��~*��B8���+ׯ�4����7l� k�UjF(�@�;��
���D{r$��kL���Q M���M":}2�>z����XI0_1������2��Z�Wص����ˢpb|�kq�����P:����[ȣoN@���-�
�>P�X�w�)����}��Opީ6&�RC,V7'ڹ����%�9�^B�$�
�h���;D�Ufw[U�^L�����2fթ��J�hy+����1�*����#��Z��wwm|ϊ�ڱ���]�����|�E\��t�Z�--4d��?gb	������so�'&���쿅l�����x���M?<��������R2�vKiW~�J��4Ft �%�l��}��P�F�C
I�%���d�H���V2/� _|1���'�'��{q�@�tE�84b%%����Y\��L��*�|$��,Ħm%j��]�sK[2y����W$�t�L��M׫A����c�C��'/��	�x�\�-'B���({5���j���܋-��[(�9�!v���+hOA�X�x?\&aą9-��S��YP]�b����-��~Bb�_��a`8=��N�����ކ�%wę��ٳ�.�� %'��8�2;���q�U���>
�Y�@���6<��G}-�4A�{ys.����X6a$�`-\�Ҍ㒃��զ���f���h�h"��J�p��N���SF=Ƥ����3�oA��P����ZS���P>L߆K����F���c1T4�)565�Nc�e�HJ��@������"��ͼ�R7C��v��㧜IQ��MD_4�Ei��H��w��rdx��� .���Yb��!D���6Vq�B�ǫ߭ϯ�,^�5(�E|��;E��I�����@�4��Qq��XY�<6=�g��I��zb�O���m��,/���}����@�lR�$�gx��0dH7�	���?������`m�Z���hY�(��j[���p��_/cL�ྰ�\�9B��:(�2�}@V�i��4-wu�@�oV���Tf�:"s���y'�tU���$i��Y�0��c^hg�U`�&� �o��⋖/�@�J4�՞����ň$�"���$�n��}����@��ہ6y�^}b�X��F�a؈�����+���ߟz!~0��U�6�e2�.�v"��%]bC�V��{�M�W�~8�[��e��)l4�@��_N�]T���)3Y�fzy��8l�`Q�s<�����@PE����x:�&LB(N�tA:�SB��NP���0`����SUaz�y�%��w��˄��ڌ����s��ki+U��i�a���d���!Q�5�2�I�q]�4�*/|>���R�e�T�+įc�1�g������%�5�d?bfHbax��9�x\�u�m=q��H�2�|���z�ͅ��<ٿ���"UC��t`E��2υ�'g�2��F��C�����{7w&Ξ�[�]���Ԟ�}L�A�Ba��c��%��z�H�;�����>���~�'�s{�R�c9���ME$y���?���̗���ٔ�3�.P��5�4�*�&N~P�5�w�q+�P�ђ\'��]4ƶLz�2�F�9hHa�>�u���9� Q�eJ.�ď/�)Tƛ�����+n �ڑ-�$i�̤p�"��?S��pBh�#��J_���-�3FM�4����s�Ԩ��Y��Z���M�]�Lλ�H�|7�����uk������ Sye�5��;Q_B�61�j���JM��<vO?A�Z�eZt=�S��P�;��R �)s�I�`�cEB�~�[ӽ�Ea�jwt���r�*���o-�J�8��~�Ʌ[3씑lf-��F>Z�G>�:M�w��c��I&bf���i(w��P@������d��h��ɓ���'��޳�����i]�n����^���w�C�a��ә�ϱ�L(�v�.�F�7���--k������;!�Y� ��:�5�J����͢)$��^�K��5�0<A����2f�ѥ,�N����t✶���-��s<������g�f����>ܲ�&U/wD�/��S�n�X�T�v��%� �)�P�픧������M��;{8z/oRx���èٛa�O�h����坮iز,z�]�uշ\:97����):���/����7�Ǫ����.養K:8��P0���IxJO2l�B����r�K3.�x �A�.��j��a�ԗ����J}�{�$\r�0{�N���^}�� Q<ZDP��o�[��8�N�!�3�@�-��Հ����\k���}���ఢ�a���i�	ڮ��tR���hx���ŉ�K��H�����}HO�`�s�v�*p ����B�nЭ�ƎÙ��c�݂�7��u�$@+��u�ؘ��2�k9Cﯾ�,�OxUH��N��� &F�{M�uM⚝B���h�N�Y���>q{�.e�8\��N�3��>��ń�~�`��f����H�u�w#���l4,���aS�mjyO��U��oUܾX�"�UE,�U�ݲ���SN�,����W�~Xj�Z'ޣ�1p��3�u҇��Tle�}4�'���?*d��q��h�{�cՄw��z���3������A�����w19�g:U�q�?�B���w�T�E"k�:��/�����x��Z����|�d��Dr�<�O����r������7������̘_�W�_@� �?{�g0i�ԁiC~� ,��p)6����Z�έ�({����ʕ�0(tB�t���ν����t��//��=a��ًA!��u�"��91�Q
��+Ԣ5���q�E����%��г�F�D�3G�&˄��)YYp���M�y#���Y�Z�']�Ă��R>	�X����˲2~��vt)�S���`{N�O~�q�ͤh��@g@�j8֓n�j���2y�t��B�'D�t��:֍��f�vIe��CU�G#Ҝ�x+��f@-�U����s?�t��ʲ�e �4y-�W����+
��?6]{
��#����bA�����`��*����7I��D�:���B�"
�Y  ��~���j��@=�Z	�zq�-=�њ���'���g�H`���d�&�꫑���Cz8jX�\���,1�w�I���_I���7�K��Ȟ�0"6��D9���{f��l��A��(��+K���P0>��uG�a�oEt���`[��¢��G@v׾�'�������>���f4��`zѤv�ץ�3��b�{�b�E����N��Ie�[���?�[d]{�!w��ۿ��|Mj�羧6��6H�S�ER9�2�*�_�z��A�^������_0���R��{^���J��_r�)W�'>y��b�/Y������e��=c�0�wCF*ڐ3�g feD��+�����M��4��9�4�!�?ķC�6t_�<ޘ��	W���d
F�P���;Ԑ�n����?�:4�t:K������{�g�����Hk�e0'T��q���t�6���N,3���� }tV皤ܗێ���1.�޸f��ܬO�R����a^%!�����/�J<�
Xa�+?�\�>:�V��P�d��\��r�m�={Ǫ���M<����B\��yy{��5Տ?�s��+�"!�H�&OS2�X;e~NT@�Sy��I���m�0j���h�]^����Pf�����DKll�*�1�x��,\��*����������V9ШWk�g2V�9oR<�]V��sF�v��O2���m���m�[�Q&�%4�!��:������vy��'�HT�~}�����C��eA��!�g����0�A@���N�{U�N��X��KZ��)��5�@�+SǾ/Y�#���r�)I�S�H�s�����}�/��RcAH��Y�ɄK�\&r[}�Z�QJS��h�j�@�=|=ҭ9[U���MT(g���`�xo��G7H�I�v��9*gَ]�G|��ϟʦ��}�_8�3gf ����Yekl��%.�a]\�|���cm�H�s惉�����\��4��'���b��L5*����F7�'�gP�ʽ4�%֒�b�����o<$��5a�$�EG�圲3��l�fAvZ�Q�E�:�:B'ŋ�j֋�֒к�5o�'�*{��� ����O�5W�N8��V�����ƙr,t��آ�]��0��{�
�,���Y�[���*�0!ɳ���kC?sV��J���V卼!)�g��	23��Y����?��� ���W纎Y�u�9�Gc�O
8��7-�c5��c5�T�� ?����b�"+h�0+�A��Â ����.��!��rw�;Ǽ�"QL�v*N�m�� �'L6M$��Txk��Ȥ9U%�n��K���ŌɝG*ឭ�)-;e�I���~���v�^������BL4K �@��Qp�@�4Z�'���]Qw讀Q��!����Fi�wi��~�bX� �q�9kr�A ��L�dc�Y�ȁ�-��7��`�ʄ�^3��|q�١���|�#�E$S�?��!���S~�_�Np�)4��ݘ���Z�r��+M���n�ȫ�[m�z�v�+!D��>/a�֝'�m�7���cAz����R�.�7/]�&�J�@�Y���@2=1o��)�R���D�Mn/%I#��8�@��#�;	�-�[G!��G=u�`|�_z�j#�0",�}ok����/��P��L"�o١A�=�+y��[�K�μ��v�L�t�������&&��ܼ+�f���?	Т5��Oj�B&Q�PL�W}B#5uS�|a�:`��sf� y-��9Α��D��]���$��a�j�q���&T�#�K�~������aO�j�zx�M��
��_�F����5t�n4�p6��lo����vbr͆(�����ja:Y}�������%\O�ِ p��cM��	�q��EMY�T�.���n�C�K<���u�KR�TM���
�
��b�~����jzy� ��w0���د`#����6�a��!�c�3�ƅSgQ���{)�y�R?cw)ٖɾ9��޼�~�]=|,C�'Z�����n3G)�����"R�O8m���\j�U⵲`���o�f�:~�deT�TR,�qy��Ve%�Sl�cѺ8�Z>��&Wc~� �n.�������o\� 4.�l������#��g{'�4+�\+`!��3�^�vUWw��E�%����	TP.�c(�����'2�H����B�����UP�Ǖjq��w+WP���O��\;���U��l䗯�i!�܍�,.%�P���p��!b���K��~~��-B�oJ�hQ8�9?Ӓ�Z �3YZ]'KO㹠��P���[�v�I����1����1�u
S��Q3M2��b8sMALlS��ҏ�@���JS�It%�n|�W+5�!s�9�D��p5l������^��"�K�5o�}]p7�^�E���Ƌ��6��x5�)��׋�-�����SznJ���T���bj�*� V��h#�x�9�ʒ�2��@�LԘ�;i��g6vC��&���%���-���Q��{c��$fU�jV�P$�k-HjfA��F��N@]�<��1j�7i��6�8���D��;q#�ym�B\n6R�r�3�-Ӹ� Rd�*��o��QL�hWV]w*��H鬧��oڿK�O�23��"ΰ̡��Y)_��"�/��}t�H�+P�A�{�=��{�K��{u6��~0;��T�䀐� �Yv
r�X��HI�A�]Ε3rߥ�D�~�stF-~�U�/�չ�,��(�@��bs�����*MZr2im�	�\u��ι��Ј/�HHjG���j*,č��gV�5Z`w��2�9K��¬,}뾚��q*���Nm�\�:ib�g��g�ÿ/h�]��������(Y�{�0j�^�b��8l��K��f)�x����c�mM���A�����X�X�K��|�`��x��5��	Ta�z�'! �T��6jb*~�ݵ���?2�\�:��	��k���U�0�*
4Q8�rW�2m�#E�3�� w�Xsk�����~z�
`�7���uщ��kw��ox�n�ɚ�@�f+�Q�r��l��������W��:M�mC�x����h��3��幺��C�,�͙�`�	����J&~Yyh	�#d������
.��l��%�G�σ�Q���}4X皂���6��$�0�Z�o�w��"p�\���'�]�(�a�e�cu���@����
r*͏3� ;0�����&�>�驞����|�(5�(tóH�^�+l��Ę�ǂAj0�"�n)9��@�2�X(��������zV�k�5��Z�t�I�Kb_��ZoC}��Gx_G�A�֥�X��Z6�l{ ���b�)�T����F�j��+:~%����/���4���4���D�#��!�=�$�c�s`E����pa����ec��ocV0@}(�%��.Ad�ts��Zy0�$c���S�����@�����:ƒ�ճY��ua�W_I���V��f�j��1�;j�	Q܄ԅ[I�S�d)M��g�tt��0��v^Y��6g%=��"�
r~��},�C�(ʯ����F����TѼ��M2e����X~�o46������y�������X["2H<�q�U�gysB��N�y$})\Yu���+�ceo?�ѫ�q	��$����#���wW�LJ�,A�׹�=й[���e�g^����7vn�y���s�$�T�\Rk��/�<��FK���if��_DP� 5�B�&|�}|	�~��ܪ�EE�/�hR�r����T�nI�������C;v���=8XuUR���O��)�gV`��%�y���E�3�j�jDv��/1⹈ɷ�1H��h9�P<@բ��Nh֭��_�д��1�!ml�ŧ�.A�K�	-�Cc�;b��\<�&8i*dL�;+�!�|_��t_�ѥ�jFa�8`��N�jfţ��F4>���$QZ�#`��m ��
X �g姟�cb�ut���%���}��*4z��S�N(ҷR��/p��� ��]��"��Z�U�C�M�AJ�糀�2g-X+/���Ξ�{�ߺ��7��S��F�5���p| (��(+j},'ݏc+V:�J<�X!t�'9,ӿNn�;�ء����FD{�b�i�Wo(J![${ Pl������L���4�Y0�,�p�Z���I��5~*v�p�`��Z�P�����M�FG�����NoH.`Ge�i/۫9HAi�4A(�"��C�?�3�*ܸ�S�J?`�357�o'�Q��Mo�b�T�^�
�c����Z���8.�F�&����KlDR
8A ����q����	�gM�Jח��z�H��j���K���Fќ��!�;�-�{�H�ZH�ymb, �l�i-AP�����l�w�%g+|�V��E��#�>����^�XX�2��&�ٱ>gP|O�����e�F�R��b8�.��/���ci��"q@��(�ˊ�@F�w�'3s��BiX3.��Ǹ�%(R��
Ptm����։��ɽ�ip"�~\��6��+¡t�c!h��\�V�GSQdP�k��	ٲL�ثǖ
n�y
<�D�h�N����%��p��ZY+� -���X�׋OB�G�٧�Ce�W�R�X��1A��7vU�f���Aa�i^oTN��&�H�α������r�]��G2tn�Z(���r3�2L&�K�&���>M�ò��~��_P���tf��0�O�D�c��Nz��Xf�0��3���mu�#}n� �� ��wFI��gΟe�ժz��O��)T�-�&P��HX$۫��e��ՒRi&�˩}����������I���[,���\���#D}:�f�ej2����aw�"���ݓ�TK�{�$��� �-�{���bbo��U���<x8�� �6������k?��LR����d��K��dl�����;=���? <2���t\������T�Y��k4��V��O)����*��ol�U0u2R(<7&�l�/��\��?Q�~�>��8>�̡�J*vpp���n &�nb.�Mj�H�:�-�I�(l��8��۸/h�:,{�#�]q3��|��wo��h5��!��!G�����=�7��������խ\�JI?���ߘ��7�oD(�읥��7�}N���k
��xh��Q���12�}u����}�u��̜�Fu���i��wGKh�=��*cS��.m�Z����(?�Ťiv݆eϘ�> {�0C7Z���.��I�l�y�`V��С��k�-1�U;	i��7��vs��r�\Zk�zȊH+/��Rgh\�iV�/��y�A��\�DED}Ƹ��h\���R�|���Y�H���D�s���3�D����O���D@jc����>��"_߾b����K��
_R�E~*�dD�[��>ve���Qa�򎇋'N�Gg��<�2���nǂj�jC�n���#z���_5j&�,Hzs�Vm[jMq`���$��82ڸ~��>�Xpn琙sn�""0q�G~���:���ǿ�A�p.AAWA9�̅Qr)ؚݼLy��/�h���	V�ݯܧ`����t�82c�V�Lw�!�~j����kH�f�ތuEzu��֣t�j<ĝư����95W�r3�w�zМ95��=)�-�����2�o���Q�8_�9�2�b�e��<�#�_ǌ�ƊΟ$C_�$�P�z��(|��������du#~- =�.�&�3���yB�k9&H�5���
��
��38v�[�G�vu;�����=ZL�c����t2�?)K��:��"�M�v%��1p�D6�-'F�R~%�qVC�ga����A3y��ʙ������-�b��	�Bdْ��_�Q�R �|	M�;�%W�{,a;�M�z�_2 ��]LP�Do&ɏ.Hy��,.p��0&'b�4��(E�����Ď���`mE�h�#=G� ��z�[@u�6�9�����`8c��K�v�N�#X�@N�~�K8�=���վ!	��_زiD�63�K��ҡ�7�'��
�M�8}�R��;6#/ ���[���Q����Rz<�b�b�-�J�,|q<EU6 ��mj�[e��ہ͵W2�w8��r��1���$��H8��!�p�	�b��$b	���(Av���b��q7�;�-�ܚ��r�]�pjJ��,���&U�嗀;�y���9j�aÎ� �	B�O l��F�	���[�͍���7�#P�%B���."�#���a} �;���Ӻ%Q�ye�q�v�Ja��y4E 5�E���g�����CU��{��Ϡ�>)�X�y)�����c���懤Z���N�ړ	�Rb�'�q�L�y7B��<SJdS�x��`��>� .�=�L_�|��~�j0ql%�a����M�k�7ij'�Nob�)�Y����얫�ߛu��yN���Z����yDyPM��r���qs���!���E�C�q�g�89�.d���@�{�P��L�۾���&sع�Vk�C_�ߜ�.j���2(�G�=@$�Uʅ��*v��9Pg�X����c{��6�"}u	1��o�2q"�70�F����V`�3���ۓ�D���*0�*���׳��*&�#�B���$�V.���PG���CP���j
h��q��ag���eY\\?�B���vRe��hp<�E�;��e��xP��w<aHL��Ԇa��>�\'�kRv�4ŬZ�i��0MK������Y���'6͞y����C����kA�s��??�rK>XUa�j�a�����:RS���&lDl�A��gԳAKޑZ2b�ap�p~*���%�� �]k���anaX��z+���k���^W�W =��
)�p�Ճ>FY�y�c?V�8=4Ѻ���T�fh_�������o`=�2�J�<Ew�@�iɃ���S�V�BVj�������_���Sy=��ީӑ!��m(l�UΉu��[i(�r�>u�c@db̽`�.ЌI��\�\�V^n��HW�i������x]O��G�o�2��N�D��n��{\��|L/�7wߞm�'�A;��/x3�k�$o�è����-ހ���*X�F�2�/p�X}{D1�'jv3�����q<�ow��#�ff������'�6ԋ����G���*Q�־WX����)���q�ã��)*IjdI���i��}  o�����*�����������_�]N�����՟�	�]�x�p�������I��~��w�+9���B8>7��|&��7��x�lLE1��:�I���������%�J���~�<n&U��Ӆ!�}�g���C$}X�`92����<�m��[�k!�iN@�ޖKM��iSq��iw� ��HӬ ��)���	h���	  T�J��������J�԰����Ϣ�e}�mӶU@�G@bb��jôo�Q���	x\��AW�i�M󅈧� jr�����mR�%C��9�_Lȧ��c�h�6�⊯� ���x'��f��ݣ�cGHZp1D T8�-��.�\��W���7t��7�y8�|��g�uc�E�%,�?Hַ@�p��}@ۑL�=��ɮ�.���i��3��%��{b���>x�G�,�l�_T]���g}t"6�0��$N����I��*��K��?1�=5�ĩ77Ѧ�(N�pό�+ƪT�P���bz�� ���5��<�tJ�@_����r���HB�O�;�ҋ�qfB�8#d��P�/�����>�5�C��6��a������2�H4}����G��D#/���a����AӾe�);�ݻ?[li�����kr+�hf�>���ڻ�S���F��T�i�c�R���]����0J䅏s!z�<�oF)�e�5�p/Ҷ��lz�/��{e�������k�;c=���n9h��.��=��,�a$(����v��gi�;4����%/�|�Z�Ѩ�PY��u��/v?���fQ˧F�Zn�`V~<p�������=\#16�w��l6���O5��X��h��|ŀ�ֈ�|�[`U)=�i�S��n�(�'O��]�	x�w�3��g
�H�F��P�-L<�Eo��cH��<+52ь�Gf���g�|4���(ox�m���S`�F���JA/�Ӯ+YW�tk�+�?����N�v�r}� �7�8[?mj�R4��Q�2^��/Z�����M�ޙ[�1��g��hZ5�V>�|��lV4��\L��5�oɡ"��Sb���&LM�"6V�w�^��,?��|f!-R�B�e�&u�=N�͌Η������j��_��>(~_�x�+�k�:G����􆪛x /�B ��9�K�����Y�s�o�Sƙ�G����c���	���u��K1P۷�����I�g^�Mέ'�dbVAH�
29(=���6�.I�<P���ih�R�`֌�+3����{T�Z<2�w�f��k��ό�K)]-D�`}���yԃǂ"��S�ȳ�����s9/)|v:����s|���3 e�׼ka��$��i�ђM�E��+u�Õ$��칔��:R!u��i�*��P[��JJQ��	q�*l;��MR�I����?��mf����H�G�f�TbRڏQc��f�/<�G���3OY�ѝ%M��=�F����. n����Z_i"����)��������gSR�sBġ
	yKxu���.?����Ǵ7��5�??2��S�޻<KtE��p*���&u�n^��AJ2Ԇ'v����M��LSg�u���s�@dZ�iY�q��o҉k�xb�Ԋ'�j�i��	3p��7��n'�*���n/��T�Ɉ"��	[��2���:��#­��$�r�*'��ߐ {�k���ݐ�"$�[�k���v�fmQ�Q�?+�(E�$�X�l�d�W@���qj��ɕ>��0˯�3{VyJ<@�� �J�c�hC��,���RT��cA��0:��l��~�ʓ���b�>�[�ײ�(��}Xْ
��D#����Sya}�&PsB�TI���E��(<�^>�:EN4���95'mI��V�i�RȘ�������?o����j:����	�Ft9��m��R�E��&���~mm,J�a{`����x'���V��f5��Nزf��
k�hP��a*���b�@oS㯐�l=~9�ژ�4�D`�&�L�W�?uȒ�Y$�Qe�����efhٗ:�g�'���M}�ꇲ��'�ͩmh��ȷ̱�D�Br�4���d��H��s��9����&f�s���qO� uh�tN�-�x92��~��q5�a�Za>{� �rz�jk;J��~�YM�.�x�b&�W[�3�f�e�?Z�������I^��a��:�P�g�G.�ʋ@s~ٹ)) Ӿ6�"�-�oX�۟��o2�C{��sT$�"���"�vҕ�iNY~h\��_k��L�eyg��(��l{���a��)�kT!N�SW㠗���b�mWYDn��*�t9y�4�B�²�=~7!�Z�S/�aj���`�#�AVǥ�J��o���X�Dǋ\��e�����ԣ��1��.~N
��R�I��?�+¼{�u��g�*�|�7�2��ƨ�t��]m��'w�
-�ݮ;2!xK9����YU#��3pQ���cz�C�U%��8<!�-�6-G�f�3���'5�Z�D�^3�Ğ8*-����><U���@	���������+->E��jΠ���x�!��Q����d~���+���#*$l��ǱYAn�7MX�ׂ����,�������>����J�"�ͫ�����$��� `�rw��p �8>h+�f���(-\g��}���f�?!9�Xm���"�*�$�����������ր#�$��Z��g t��L�Zk1����M������CᆥR��yݡxt�W��HYP�z!���#ы`7spm��@ܣ���N0�"�����/2~4��$�O~�ڎ�16H�r0U���[���Sm���
���%2�o+p;;� �;C��6��R�9��CJ�iJ��\�(l�Ƙ`rRgS���ki���(&l�>l/�>{���I:7[%!,���+_�[E�P��ܣt�E@a���)e!	��5椇ը�J�a�ֿ����ja0X���0w��I����΢���q��d�G�N�<q���0��,X���s$+�����w/�)������4e!\�DA6�4���|.js�-�f�?�����:��E]܁���2H�q���:��7��}���m0��gi���n@�pt�;���8��gR����2�dm��=/�݉F�U�ػO�Z��:m㪤����0\��F��v�-Fl���ҳ6��C$cpG�jz�.���5l�J�o�!/Zut83����~��?���"������<3�u��H5��k!X<�#=�z�^nk+HKc{�f՜�2(09�<�����_'�QHix ��� �(�Fr���;p)!(F|�J�a뎐����Ͼ�9���H���JV��ؕ��ߥD��H5��Q�X�nT�0�{#��~ҿ�Nh �E(fE��c7&�ږ�Y�}�?R��s~P`�.ѿT���46x�$��H1P.%g���Y�sJ-�g=�i��03곰U�7�1f�E/~�D�h6rQB.�bGay/��/�{|���>{�]m��@,��L����r^��Dj����ݠ�O�?NI�q��0����>uz��<��+r<��G��v�e��*���Z��+\�^�z���q��$��]`)�	��%h=r%%�Q��oO�l� ��۶*��޶e`�%�t��	 #M�^�-��ok�~�H�$��
�<�F�%�k�6�}�卣y����+C��6�����%+���۳g�o���r�H���_�I�=��˪�B�w�&�vVfܣ>/β�<: �4�18��u��d�]9ůa<��h�'Ц[����yA�T"�f��7^����-��U4���C1<~��Y�7���.L�����!��������|�r��v �`���8w�H��?��y�DC�`�y-�ߔ������?��|r�!?u�Eĝ�#(M����ԥw�<�D����4���èK�>�xM}T��kP��r01��X���Go5�r��v(��*�>�؉L��n��l=_�s�Woʗ:�R=R��Y�	b� �,���Q1V�;8Ԯ�ܚ�@�� d~��7����hYXlЬ�ޛ�+���	,st=�b]A+fv+|#�K� ����})�ƙO.�����e2d��Vv �{_I�<�Ȥ�̈$�(pe$d���m��v��ܝ�IF��i��xG�.��)����d5�ty��m�_��F��u�oΟ�gÖ
H� Yy� u���&~��uv���W�0���VG�5?41?�)�����1&��׭x��vY+��"�&*�v��!$��:I��$���+�?j8�[��Y@K�ш ګ���}�hf�MQ�������JoW�ʿ��ǖ��n�m+#�i��A�����#�{���f��qM�i/l����-�D�+	�&�����w�q� G
e��&4������H���(������ƉQp�YS�p�b�@`����@Aá�<�}
��u�,�rz���{��#�0 [���+i�Lsn���;�)��Ͳ�'�Q�J.����U�a�}z���J=f��k�7���b��=)�7��W>ʰ��	��^P�c�A���PX�}�	D2z�E�`�1�dpj�j\lC�%/54VY���b&r0Z:��@b�A��l�L
��h�
�o3AGK}ȵ� �
�����.[QMJА5ǻ"P>�����w��象�@�c�y|F`e\JF\���6����vDӐ������em^\��i��Wc.%�Ŀ*���Zo���:�yDh����$=j���hw�8�.[\�j^��h��rn7~�r�-u��Ft����<v��6t�}Q㡣r{�"���	�x� �H�j�U:ȔH�y�D6Nó���
�����Z�����Xq�҂���� iw/��m�Ǫ���NQkM�o�IuU��}Ƿ8�C|�_�g����)R�m�Ҷ�0�@Uq��R��o��-�E�wwS���s��eĳ���(k�!Z�C��������ۢ����/յ��W�ZT�Y$�p�qm��o|N�����h�O4|5�P|{WD�64B�z^q(2�#��Cw�~���ax�K��e<ef^Ł�@��DWh����?�	��"/����KhP�zkd#�jr-Ć��m$�o���ȯ����c� X��ez�
�q��XL�>b޶�$W<*�7U�_@���L�-+ʍG�Y*}R[�*��I߳١��iw�(��4!�����ԓ1�)��W6�/#AA�w����m�2[<ڶ덳��������u�/h<Ҏ�V�#\�>%PE��q~�@�of�K~z��K����w.����������xkb�/X+�T�!!g_Ӊ ���ŀ�:���8B��/����e6�
O����q+�5C80�*�x��v�wA�?4��q�N��k(�� n� d��rr(1��]��}�Q�Q�����-)�E �P�*��B�ZǸ����B�`+ ��B�N��l��*3S��ynF[�g�9Yh��1a�S+T�m��d�@���9�2���J_�̞q�>i��ǖ�9��\D��o��o�j4v	�c�����D1�anc��Q'j��,�J1����SO�Ddي�~���!d�6� %���k�)lߡx$�u���ye���G����t��S��jPc���v1X/VD����G\�x�r�5�:X�;��Y᩟us*�<�1��)h{�Gbc�ؚU=�S��ӥ<����3�<K#���T�8qR:Ie�Åyr�*�~�)�T���NZ鰞ef�v�1L{��q��Y�<�=����U�D�z�3	A��O�vUӰk6�>�Go8�hK�j���vTj��,��j��`ܑ��+u��AE�l=9D���*L=u�h�P�-85�Ȓ���K�m�V[�Ț�rs��\�)�>� ꜹ�a�>v^���<��,D��'W%$��:�.е��P�B�Ԙ.�>�����F!��{��*��bk[ĕg@�Me����%�p-৅��d���PG�1��� ���{ӻ������&qI����F��'�u��7o*�\��K>���]�`��A	�G�&�I�2�@�3�x��a���s$�Op⣻����H�2�\0mR:�Y�E�8G/�=M$k���rZu3�n��M�I%�5y��<B�Fi�u���6N�P/a�TR����b.�MJ�U�O��E�μ��d2��E;����<�H����L6��O��xᦑW�1�1TDPy���.���7�l`r ���	�H�xK���q`kz��QU _�s聄4U��*/1�=�?���x�l��"J_Y ���=��a���ǹ�����'�-���=�ъ���#{���Oo�,W�pFj5��)4��/���NM�|)�'����F*��$`���"��Ӵ)}�H��_*��WI�|š��	���5`��g���@����LX��w�Ռ�D�h%fɃ=�r�\��j��l� 2�lK�*��-��`@�c�	��(�-�>��~��Q|O� h6���������w�p;]�� w�<�'��C�r���;}UBZ�?�ri����ȹ7�k��+���[EdD�&�$lBt=�u��L2q��,:V[�sp��w��+Ɵ{Tc���b|�_�Fa����\p��? Cƌ�uL��hf��F�/��^ݤ�1T�x|�Ӷ���z�c	��x��v�Nj�l_����T�f
}G lu!d�p�F��^��H0�#�z�^8Lr\m��'w��*;}4�Z��-�j �tb��DJ���̖�M�'?[����R���]��	W���i`k�@ش��!���C��uﲶ}�V��)�j-�Ђ�H�I��}Gב�>���+�C����,<�iL!SJ�k;ح:��\%��8*���2�N�B���y���3��^l_��R'6cv�t���ˆ3,�X�S�x�su>Z��j}[��P�|���f�OȆ}�̙eɥt�nn��qV���.� x��4x�!>H��U��q:�X��:aq�ې��]��Q��X*�b
���"ᵬF�Ә	�{Ѭ�Q��E\��5a���l|	�q�(�ј��Ǧ�X鱖���*�v��]&�%��"	�35�E��#�K�.���	��J��[���X���Ƿ4S��ѕ�O����I�OvyX�"��׍(A5��� ����O'!�e(9@�����5�+����p$�T7UW�2�N�]�|���ܺ��n�/�޺[ .p� �*�VL������m�^�Ik4�t�&���@-?����F��0���R�����l�'�9�h���>��#Ñ�R!ձ�0h��o���xoD��H-3���p
��
�2�����k���zel���H���b�b��Z�~���܊˿� q�/p����is� �G� �%���Ia�����v����M�7�M��&D꺪	ą6*^~8ў��c�I{�C�oG������Ӫ�i#ļ���B}2���r�uO��� n��,�,uQ��@�������4��;Fɥ0P)�|)�SJ	a1R��;`(H�M	 v�ݖ�{���_&�m� ��lkӟ�����+%&�^�	/��^�Ĵ������]J��M� ������x�~b��}����3�2����d�E��2�g=3����t����oΐSd���>�CVy�f���ʆ�@D��N7��#[�"��BΪ�@��[Ft�;��G�u����E�ϹP�]�!�����-�R0N����*��W��s�G��H�~;u��Z���D4_��Y����;� )(��5�>���l}��H��եb�ߕ ]�e���2M	h�S�Qe���pX�J�@�H��ڜ��{�X� ���_ �g�F����bFM�P@��V�Xxoπ�1#K}�8{9���)hz<[��om�����WY�ҞpXor��@B�ku8�7K�H0~P&�
���U+M��/<�.�a�*��#R�(#R���]���&j�S�߳6�M=�\���=�,b�փD}!��#H(3��y�n�<��=�8��/����@���I�g�1d"�9�lFO�N�tV(R�3�� &.����֫V����D+��1���?���ޚA�|�̠P�!SA^�_��T��wL1����_R.���D�W�T��ZUhxo=��Q��2yCO�א�uK^�Ri��2 ����,��B$h3����VtuEz� �������*�d}"�&�Zt
#,۱�f����1�%ԓ`�4�'h퀏RP^K)f��|N�zm��|*G�r?$�;������wK�����2`x��Y9�i*���J�gJE�o���d�����t{��k̭�7�Fr8��<Mf4�#��c��C�":�SU���2)���!�/�:K�s5�:5��l�Pt�em�=�fm��W`=���o�N{Wb}ɕ���Ҽđ�a��i�פ�<K6&�R������:��-�:�eBnfw�#�Ă��Lsh���)щ�/���yO�1E��}5�v��Ʒϱ)�=w&�������Β���&F	CWS�_�N�,+�u�l���8���V����G�o��aIf���8��V�_�u^�n�yBD<�X��	��D8MB-�9�hRZs��e���047͝���Bc�z�S��>]��
]���̇�a�@�C�Jtz�PF����M*�_ʵ�m���$�+B�>� ˾�}�F��Ԧ�`�0�o���䷜K?��d��i���6��Ӓ3�P�8�W���	ĜN�i\ݒ��ƞ�����R,���[�r�t�bMC��8;�'�=��ULW
O_��k(l���8�^�AɱY�s��3n��Ѿ�pU$�~9��i\�ޑ�p� !C�h}�˭��
=�����ɩ������n�]�f���b�o|_i���!_ڰ8�Q	z�
co��0��}�����j�I%�0N�y[#��H�)�뗛���!�a��fK�[NcQS�rv�|s�A��}Y�p~�Hb�6�T��Q��&��4v)������K��W�AkC���Ӗd����-#%PD�g�?�УxW�L�؎	x	�� SNcd�� _��f0F��]\�o|��4V8���&���`RN�U5��V��خ�U[�:�ɼ8+`={�8tU��&k�I���)$��/K��J�B��ݤ�$���<l�5�M�� ��Ѡ���h�(�.�I�r�fkQ��-�R6�U��R�������p"9��H��8>��W��T֕C[�ajW�ĸj��h��l��G>��4w0�Q����}F�>�G��x���Y&��c��{�Ue���+DM���~U{��b�_"����k=C_zu�v�Û�+x(cj>�?�z�9(FR�tk�n16��Sh��B%��_�#d��߯�h+���;=6m��eL6�qE#~M���X(w�����i�&�e��w�p�Ԏ� �#~�"+�T0������ˣ���TZ� iP3.�t]�\'��.e�FC�;�Xt#Z�漨�U�Q��Ha�V�8���T��
������^Ԥ�j^�G���\���(s{E�7����{��qu�S:������v:EE6��5ȖFG�IĔ�[������A��� CH�W�|��,����Z�7e�F2�����([/�l��z�Yņ;(��f�\t���Ϋ	�򎼋�� �4�+�3���rS��������7s'd���3AB^�דby�� �b��7�_�a��5):ڛKBOmҿ����\�Ij[����ѯ�*�)=k��҂�:3�@��jar�;=�d�K�կ?Y�/��;��z-r[�*������V������T�a��,PU(:��|k������ �š	�;�N�J�׉Y��lsL\����f�w5Ί��mJM�����;�6X9�t���/��n�2���Cڔ���/�͂��2��h��I������f1Y=�����`~G���#��^����>�Z��/eW�IhA3�~ѭ�O�?{,W�%���P�v.��Έ���"3�N���	� Ɲ6n�c��s��²�	���O�kn�t�C�:�#�W�OP��b���P�-�Q�V<�l~%m��̝N�ݨU/'�/<b�|w6�kP�%�-r�i{��[����Li��tY��f�즟���%x��n�iocmiaB��j�N�d=*4�����#[���`��P��2�t�xm�)�8��/M�?�W������&�ov�n��ه��/0����`k�I�����w��������YC�`\�	IL��Q���]��B�}�Ί!�enq�K`���<�>_�t�ZoI�}S�J 9�* �S�.Sv�B��o�r�,��.p?���Xlul=-h�m��k��hqUq�`��t���Բ��9��]~xz>{ޮ��շX@�{(�w���Hs��K3�V�/7m��_��s�l����B�,�:�g,E��� �H�I4�^�:��?#�O_7�1���P$�������zO)R��+\Rk��3�$�A����ͮ��Zx�^�*��f�[�!� �ȵ�I\��	x����$e�����#��@��I�=.PJ�2�T�݌��뙵�̜�͛ ���m�ݰ�0��]c*�8�vx�
Ͼ�ۯbܚ+4e��ү��!�y�;�NhME�X��X+8�����~%� ��`�=�4D*h#�>B{�5⩸��\jEydش���<�Jtө�2�J�l�g�&���8��3Jj��r=���2S3�m��􂷃34%טR�b��ܣ�7�Jc+Y9gȜ:�����������~=~5(��_ۚ"��f�%�������<W۵�Ձ~�U��K��2����yl\���Yn��<� H����U�Mq�c�MP���A���&��4���-l��!�{������gH+�-�1��[Fb�\bϊ���+�ְ�N�fi��vw��<����K(IP2n�p������]��ٹ�JA�y\&�B,��7.6x�1�R�o���S��x�/R�☈��XV*�BLx���$C���`������P�N�c��/�j���W��4�#��zu����[<��*�x_M_C�`x���ӧ��<w�|X̫a�O~�D���c��9ѐj�R�^�J�&�Y�k	-q��.�Pe�,�Q�Z�噜'����`�͐�����4�]�7�d��"_{n��fޫ�\C��� �)�(����_ru����oޥf.�D��2�w���j���s�U��r�H�P��4��D�v�y��	��IAY�qw��ߣ���h��=��Zrhl��d�gѻ�F�f�	;e��%�(ٽ<n���O�!��]x�A�$�w�!�hI���J�{CHP��7ʏ����f|��u�8~�À��p`_y�e���O��z����_W�׺n���!�XP�$8���LD<s5�6���B�)��� ���~BSJ�̸��]|5$�VLa&&��#�-�de~�*�\f&�[]Uf�A�4	�.�d�������C���H�* �2Fy���2�9���']��>d���
��i|�O��a�dK��-^�wQ�����Qn���A�����A}��ek�ZZR�U�jz8\����7w�P�^A�|��u�Ư W�������F�Fby�Z��"��a��ڀV��;�u�g�������pulg���'�Z{Qc�P�dAԨ���?�r�K��G�n�O�شDA��P>�}B��:�����g"�k<�� �zF-�>��y��dq�α��(K��^�)f������~���ߣ�M�]\�� 5z}D��^�1�2�{�f��y�n�p��rX��ʞ���� ��c��{����Jȉ��Z��e�c�����ubw|�.�7L+S�H=#fU� ���辪��1f��S*��q6����k���֖�PO�XV�����o��A"R���Gs���Z��N,�L[�*9�C^h�ĩ�/��([��Q���8�����j���R׺��M)W0��3��h1|B4H�kWJ�����=��4"�I�6�y<g#�p~)_���l3Eu$���O{��JY��dr��a��
Ne���6vXC� ls�_�P�-)�(Wb���릖�3CA�WA�#�/QNY�D�"KA.�{��u���B�!A��	�y����;BQ��fk�z���hmmP»Dy���r#:N"��5�vۧ^�$2�K\���JoTmi����uy9�"���X�K���~�:*��9!�������bS��j�NFə�x����6�gEsH<!{�I飋��.��6e���i#�:�7+A��V���>�x�
�!�:�10Yλ׳:�}��|���{[��8�����gg��J� �6H�ԑvsd���D_�������+3�I�$�����&�0�����X��q"#���"ҩz$c�?\a)��w�	����~�qpn�Z�/�t}Xi*�#�.�ä`�X���� x1>�<lt:�r�|؈�dʠ�0t?�>��j��L�U��7���#�L&8W�4-��H����jG*�N���퍑"6m���}�.����T[�(��ƕB�骭G��O��R-)��{�ZU��ǏM	Uu��n��m�p<<���m��3~E�Q`�5���Sj�4ǚ�9w+��-��`��$3e,RI@�,X�Դ�w/7����������
6�xq�f�Sr��~Ia��Yj=���3|�#y>�Q4*��voE�za�CQ+L���l�b��p�l����ЙKؒ�r�bI��{�zb��?c���|6�����Y�#X%n� �h":����m)���|�����g�0-k?��A�=��;	���P���B�1x�4l�u.�L�a������a��5;������b�6���.�[����Jv �C�e ᅀ��5�)�!��Ә\5)��k``��(Q=_r��ӛ��@:��Yllf��xC��=C�������,�ax���&�VF�g]V2%U&�PЎ_�HӇ=e�0�p�w�C�&ކ��i� �Ѿ��B�3�6�{��1���|Px�y�J��h�Fn
 �����[�3K^�I�HwR��wD��#��0e���+LJ�l�yY���
��V�m�%8���4+V1%��&/l� Ms&j�NK]�=���)f6���  ����Q�}�HOj�d�7���C�r�{Z�a��+D�kd��N^�T/cV8Q�W���!¾����EM�d���^���
 y	U7��ϵ�r�}m�aJ�¤�9g����L�OU<d�M�ԄUb�?x�Tp��~���Ӓ	:xh�pFWYP2.e����I�b�f3���|h�(t�I�r�ѢQ9� �=D��'8L�Dh*Hš�o���	ΛOW�;�d�H�����nXH!!|�������cā�p�=5�c�pJ+}�V���j;j3��|��Y/�5:��@�5#�����~#���4dtN�
�LN�Rѝ�ΐ�5<��u����߅�0���K1��� �G�	���W�����]���}����� Z�N�c׀��&C%O�QNL���-�\@0�WiAr�;�	�)KW�u��>�Lh�K�E�	"7��b��貂B=���$S�2�˳��T�l��إ�g��n�A2c � ��\qN��5�~��ŝ�?�djZ��~���T1���ߤ����[Dƥ�!�K���k�'�$�Z*&�K_x^�c5t�y�����S�b��v��ɰ�j�
�Q&!�<��y�njȑ��ٱ�K��=Kab��)�j2b(ZX�ҵ���;vNZ�ƍ"2K����bk`W2���P��v+A�CA�F��Adx,�0���bn��ׯ�w��(���_ϔ�.�"�����[T�.�V��d�y>;K#׎	Fr�+'!�޼ӳ+� �0
 T0�~�~�S<\S�.,�Z�� �O��ۣ���%w�h��b�2,O�Uy���Z��o����n�,1F���)��O հ�������2���ak�έ�Gs&�6��+�̾E�r0C�x�U�l,�����XR��7��w�kȇ��,���UUI�c��]� �ψ���Խ*�Hљ����Tr��H�����9��u|	}~�e����	�f�U<�]�+[�c�٬���٢']gw�$�v֟�����dW��P��2u4qh�Z_Uk`(I��N�Dnc�f#=ɶ�@S���#k� �]���6e�$�y.$�}m�҃$Aw�EܧY7��x�N��w��ǌc��[
�4|���D�Si�h� n��0��Ѯ�����v��.�פu�y{׋0���|ܸGz�x��� чR�:����Y���:SR��B_�kT��2w�\1x�?��QH�@��T�,ܺo�1k������C�n�6f��h����s��w�����&C�i�P8�w>L�綹ؤ�V1V;Fw3��Y!�j���[�P�}�����;?W�b%q���jR�䩲(c��3�4�m�x��H"I����Y0Q2��F��5b�[E�]�O�3���	���K�4B�Ǖ��$f��*�kh��s�3���s9�4������X�0�;�mN+y]�Tm����l�?�-�����#�"7��W/'N<`<^��-�r��9+4"A�Ì��k�0����K�*";C�Y��Sظ�}��F�X��8/��T�z]ޯ�@��V���i�g�#ط��ǝz�H\����k�^�k�(�e�ܴ�=�M$�����#�Ό}�7�l]}p��-�ߪ '�-T������%4����տ0���ݒ��o=ny�{�b����$��:��-�@ֈT��B�_ϭ4CHv�	"�r:Y_T�Q����s���F���vP��L���Y��ɟ����k���u�v9r26W�9ߑ��K{�Ź����xe@�I����`f�I��I��wD�����^����X)��\R�.�/w[)��K���Aqd5�|�ug0m�(%���O����ES=��_MVsKaPzRiu��CF��Vm|b$T�%��c�h�)��R�������_�T黗�4 ��\�CU�xB6�l�.c���'B7^_��GA�}c�6��8w@� 9)���j��L��_K����^伛�^k��0��d��Z[��M_���s(VI_I�w�`�$��zJ=�30��Mڗ	�X�DGLC4=C�5��,D�7N�N�J"Y<���$Q�O&�M$(�fY���ήo����
�vR6gP�`�˵D(߭_bג�ʥV��@�9��������,�3!���gfX�ڥ|���(<�k�Z4<1T}�����4C��^І݋�q��(R�P�_�9����3�]�V��tL<
bGpHx����kI���浡�gL�´���5�� ���u_���l`�Y����-���ƃ�!��{��<$���h�-5�y�l�B�<G2�z5�ݟ&��8{P���
4���W>���7Gb����cgL�)���w����\V�,l���Ukg��VX8Y4�v������W��a������8��m%2�O�L1̌�y�\��	T>z�bA3
G ԍ�����ھlf��c4ج��"B��7�x �ؓ+V/Pנ�Ò~̽e�mE%f� ����6 ���C�*&k��PV�6G����ݵ�����{�S`�^׈�������,,c���R��Rh�a�m�m^|C(�R�C��x!1�b�����!t���Q�`%;�/+W���	k��ژ����ޞH�O�����/Ua�Oz�>�H��и ��}�:�n�\��
K��놿��l} �)�c�讛��ⴘxF&��fҬ]b����D�6%VS��5���� �)�Uv�"M���I�Z�E*��KI)�j+v�O��!�c�YlL�&�=�W�jBo�ñ���}�y*5L�W��]�f�AlJ�
�[F=��J�'�;��O+1�emS��ι�r�@�r^�&�p�5�o*al�����6Z%��9)�}��	�k���F��ʈ�����M�W��?��Z�v���S.툮�bl�!���du�o��s*\B��|���l�Z*$؛�OD�1�d�l[}�o� w���95������_���b�*C������,K\�U�Ş���#Kp�,P<�v�D��tRvI��1B�����P��ᗑ��i�>�b3�dxET�h�>�
��D�3˝�������#�@�\�GU(o	��t�~S�����5Bs�Ik�P����:�G�*T�H��Z�@���Ffi��+إH�D�*��=�b�a��DŐ���ۍso����x�����ʠ�4l>��_���o7#�I�3�������9E#�SE�.�|�W�B�6g�H4�[$��B@ �EnҰ)w"�q	tq��\���I��~�<SmU|�z�_l�#�Go�w��T��d���X|�@v��4P	"_U��!�&��Ƙ<�>�jhy� �4�UM���w����
�
�
n�G x?�#�O=U���才�=�4~�� b��W�G�+�+�O���-��	V�b����7�Y�o܏?���H�ݡ����I�wf������I��u�}ÈR�\C��=o��!�8� ��>��\��Ѣ�e y��;�����UT���\ }�2II��p�=#/\�i�>f9�`_�H��2�x>�F]KI��M՗{�j��l���L��Z9�R/F���ҳ���׼�j>�>��W�޶�t�1���1d�Wz,�����f�=�>ZuW�Xs�qii_�M�h)�3f�$����ĉK�ȩ��NK=U3x�w��Ox�6>?<��>�M2f*혓ce��x��ސ^db'+W�B��U�y!$�����=o-xWPlr)��E̤!S�աJ�Z�z��I*���:u�6�#���1�s��K��Ka�"��	0��qDl��9P`K2��wB���eyX��(�|�Em-"��0C2Kt��=v�����&q�F�%]�+H{ޗ=ٴ�$���-ç�dd	���$���:������̭�!�h�pg� \�
�`ջ��\"i� XrZ�x!�)�LL#˝��p�PIl��%}�FJ�ԡ��͸h\2SW�~B�`�I�iX��E��v(�u�E�;_:;��q<��3��:Z���r��5�l�%�^J�%n��㪧 �Eж�H�E�N���\q��}U׈���H���ju7��}�@2g�������w	d��M��p�pXA�ng����Һf\��i���!	�I>+������4�j�s]��]���u�0'��7-�*�r�:�J�P-cu�;�+_gjj��_�#ב�(�C�'��](ũi6rn2�m���X"�������'ЉL�ݾ����M��LD���0�2{9�bÉ�CR�n?�0G�"_~P4ޝ�����[�S�%��� Z*��	 ����!K���%-K<���o4���#��9�d� �Z$d���eg�v��}!�+p�uS��t�Q[�L���5?����]�	�A������L�K{���=�m�K��R�F�06����5*9y���BA�4稃"��Qj�S��c��.M�9j�������E����MT����D���7��Ǝ��K��)U�_p��ƍ/���:c�*��(��F��V%�(6���ܘ����$g�0d��@D�s�Z����'_�]���'75
t"�;�9_�S�]"���+�i��J>��I\�A�����\Ҝ���HHY�X�=o7 ��#�˖I�ߡ89b�%�8&B�Zt��Y�!y�2.��6J\�S2l�m����ĉk�͟7&�V��OY�bK��J5�6��KǊ�lR@�W���k�r^�T\-J�H�l[���⥏wxLd$� %��!F9����G���/*-�0�rM�]ޘl�?��^L��9taH�����Β  �E-w^] Y�)2�ݑ0Le:8��ؑ�$����+�N7#q������ԣ�95hV@k�>4%T�h�a�'#�|�!��[�@�������d����@e%��&!ƎqAK1!l�g�x�����_���J׫l�����k˞����f�j�v�O��'pG/���f5�%2v�Z��>�V��P]g?�����,ʺ�G�$I��*o%d;�w�J"Tw��=�Q_���)����L2�X�w������[|��Z9@Ǝ�Ě���O{��R�j�#����D;�� ���XU�ٿ����0#5ll�_/�U��l�1a�H��e=U�j�zZ��P�-L*gM2;2��� Tt��gw*��B���_�U"��Z�t�O8���Q���t>�$5L�5��$�@��|����_b�*���mq�I�֤L�LQ�� ��q#U!?axk�4�@\��F(��w]s����ӲSg!,��H��b�E�<P� ��Vd*�� p)������������I �
���ˈ�}��BgY����-�sW�`�:�沮��A�\ENI�IL����� ������؉(-����	NlrB�Xd��'}�J[UF^��hf�ɝq�*�F�9�F����k�h �뗵��qK��r��Ikdc���&�M|�N������w����ɑ���r<�N�ߥ�-��ёG��<������A!6�_��#©�Dچ���O���2R������S�s[�m�EEݺ+�hi�ș@���1J�l��f�ut�
��ܦ�l� <�Av0�~��p�+��O�ͨi<Z�.�#�4�o��g�����>P6��n�߸:/�Z8�_<@o0��<ؘ_�ַS:�[0��G�Qfk���W�I�:%Zzݼ���lI��H�Ke��8a#�<��l�3����"Fz�ņ&c���<_�!�5����h��<ҽi�6D��� Xy�$:Q���"�aj����O݇-���M�st��&��.W��?���4,�v���9�CdK����$���N�&��tbU��s�b������Rc��Yk�&�{mrd�1�K��s8.�xQ՚1\��t��2�K�3z0L:�q3.�����ó���ꁏ֬� 	��k�g0�$aǊ���>g�o;������A����������rS��B��jm�� snj�64���#+�u�����M��������B���wPO�n�67H�J�/8��2�y�h��X>�I���j1���k�T&"�YI��v��ʴ78���X`,ѯ�� �s%���x�͗����*}�=~�#}���S{�
�C�U�hpM�	/캕��l����l��J�:�c�
�i��vOE�H�;��O5�[�AL��)�H�q+�*tMť���`�'i`��z;�~̫��8��λ�
y��z�(y��Gw[\��+��k���M���ξ���tta�Y�cF����W =���] A�ү�$��P��h��?
6,a���p�+��Q��}�+%�7y��$+F��6{��'��xۈ�a��_����k�!��t
4��X���#5�V��̩6��J��(E)�*U�ah��!%����S}pm�3�n���zM�:�v�U����&6� -�}����`F��zׂ=F!��u�rh~��kX寋�p���e�P�B!
m ��w=�cHm��,�լHdBf�M�+S}��[:W����qh�_h����|~ o�3���I���v����?���I��ӷ6lK��ڮ𩷳E��5�:��i��I�SC@Yy�a/���YcWOΛaLZ/D����`����u[�ZZ��>+3�%i��څz�'sw� �W����]~�.�(j��V�Bi��~��r�߃/-W��%$y]O�5ȥ;|��u`�m��G��?m2�\���I�����2T�P_�q�D\X:jp_^0Hx��.�>z��qx�)��HVOĩ�S�#h)b��d�^%�w��#�C��yY�V��DV��{����u�ڋ����H��Qn9M�s�M�,�s��i&؍
��FV�s��kM�H�waNE%�z�| 9�(Q�%����E���Z�EA����Sc�  ]bi�QNn�����zzBϛ�>�V����r���E���R��.N~O~A�	����ZE{��ۉ��=Y&����r~>�j�up�e�YawNS���C�"&��OK�= �n� L��W�&�ql��\!B�mmf(%9�����e��ٛ=�������;%�<�{�F�mMyhA�0��^��Q�V��p�̲�+�8���L/~�审�0�]��LC��Wf��N��d�ޠ�e��S͜R�D���}]�p���OI� ����al�BG;~۟����)��{u� �Ň���-�m�������fv������!ܭ�C�)ݐ��!��=.�w_��d����C��>��Ɵ3�*껐[�����y�`�tD���r�'��z�Ss	3�?����!Į)��K3�*��P={-�b�1�9�G�%����� ��񾮋����qDp6���k���;�)4Nq2_�X�) n��$e�v2�t�3|-��h�7�dP������y�gÜ�������h�H���.+��m�#U�c���%�� ����^nmU��D"��U��l�Q�0�v�7e��i!6ߨI:�Kz_���m
��v����{�f�W���|8R��s�g�����MA@�i5��P)�;f��y*��{�D���+/9��FC�zv�tpb-�w[�?����'�{?Qg�g��HX}̯e�Ƽ?��q�r�~I�PқgB6�<������dJ��]t�ӎw&� pr)#�<�?U�W2zͿ��Q��u;������V�I!� ���/e�U��%O� 	=K`�ɖ&���L�����"��M|R�2��
�������O�m��bz���T�5�[�i +S^�����A"�l1�Ā%�ŘԴ?G6.#���}+�\R7U2j�Z�H@�-U��w���Xo��&��hQ�
�@�`��?ɰ��B)���M^����8]O�2�SwJm/q���Z�o�^�e֌d&u�D�y�
�?{8�\2�^��ă�<�s��f��Ҟ���]pO?�{�b�����v����y�J��}J�]푳T�"l��K$�6:)�Z��]���a�k�s�W���ܪ��7��5�w����S��{kGy���4Ǽ��l�7�8ur�����,C&L]�}ʐd�:EЦm�e��ԗ�]?�V�R��O�0.�,
��Ӻ�B#b�5�$�D��R8�VTJ=$Ú��8�\�e�>G�$|]M9�6+%犯�WX#���/w�k��[E����.��S���ӽ�Vw��Ѓ� ��D�Qos���(y6�n�����Һ�v<�tZ>��C2��HC,��ܝkHU�a3ƳT�䷭�F�8)���Km^A���"o�-����A��,�h	J�u���Ȣ����;����>��?'uO���#�WːR���.�4L�1�ﾙ���KCL�o揦7\�[��� �7�U!�*:�p=�@q�&������m��Coƻ�D���qA���� �D��x��.���B�D-�dx 8O[{��[�Ѹ)��ē&���pd8�s)��`PEݍ�f�-N�0+&?�jZ�!��FI<�jW�����<���4|��7g)����1��I*�����}�촳���ۗ��ہ��S�[�[*�9��:n2��4<�& K��	X'<L�`N�����îp#4$��%�'�zW���<B��x����jI����Ǔ�)v��A���-{�j����NF
<E�@[mWp@�`�:G��K�)VB��T��UZd�ۙq7�-s2�Q�Kqh7�7��P�}�Pu��l`���7�`��XL���%\VI���7�v�Fѱ���(�ޱ���H���A�}]�zbJ�;����,s��;���:����A���d�?<U_8q'c�5�X����N�W����-;�ư�g�J��Y�4j���.FnX� ���EH�⡉��1����_j��/�m<�����6���g�NB'�
\���?m��%�X�c��Sn���e�e���yjw�z����d<?�����<����_R�DNYP�RW�(�r:�p"K����	��P���rP����v� G����ɶ炵��3�&�ރ��5����!T��"�Y	V$��#��fH_�j'�h��nt�$��n�Ek���F����)b�#9�bU�w��AbSF��Ň(��ZE���M$y�⛋��j��kjPq}�dt�EݎZc]ĥV�k?��N�wi�m���	�퀬!@�<�u���Q�&�����h��y���
��R���QU�{�Oqѿ:SJ�K��wV��x~v�9D݉:�bp�#�a~�P�]�p�#&u�����r����q�#<t,g�~D\ʇ,"'���"�	I���b����k���f$7����,Z'T�����lF������Y��}�{]eu�:�]|?��G�͈!��.�jA��0�]�Q 50PM�lve��ŧ�{?ה�o��{�]w��p�F̵��R�� !/4��^&���W���<F�y ֑(�ad�Rx�� Ii#��Ƕ�M,���k"X"�h�R�Z�E�j���!5��sr�-f��(O4��j�ͭ��MNᇭ[D����w|6<�	�4ޏK�I�����X�7 Z�bnT�c������q���D7ojj�\fnN�����"�c-P5���X��L#X���a� �U��lQ��Bw?���n�'ʛ�q�V6_�n^�k�.����G�^�3Bv氐������`�XT����<�"�\`��Nsd�f����cﯞ wT�u�ĥII �cϘKƇ/c�����=�XT�ά���ns�y�:��fj*W$�,��]�D�|n-!5��pBF��	��K9K���q�}��o���D�C�ޤ��}�'��Vqk{M_����Y�V� ��׸++6�1�:���DR� ��_��@ٵ�����ܮ�KϤ��k�g�Rg�<�`l+L��W. ���!� �l��O�E�o� �U�!dW�>j|u����WuD:��"k�T﫹oz���:���\k��%�	Pa���5�����{�������H�k�[u-k@�ꇢR��d8Ҳ�L�qWkist�1@D.tD�¬ky�6汒�i'���FP��z9\��~ẵ:��:�y��/1d$g��^+�*��b�����ǆ�xLn��0��kiL�3�4��fKs�L����JM�{�EI���çJq��Ԯ��1�}�:����)�v�����8�͏������J�v� �E!K�#<�>.���?�3����|sP+ŵ�_��{���z�cI'�!�Sχe#�n@cņaz��m"�	����<��`0O�O�-̻Z]�q)���M]��j�N�/�#��T��*�X�TU}�t"�a� ��z�yu���4}3/�����Gѯ��+S�1�p�&pb��f���X@�S%5����E)��`Ra`�]��n+>�`X2�L�=$��J�S]��o�G��Ê�,�Ғ�e�Y�=I�O�y�]��H�
�䳛��`-@!��Y�<���!�Q\��Bju�o�QpT������j
(�dҺD��7KEFT�SQ� ����o��� ���Lě�
����+���#Q|8FFYE�X�W��w��|�Ē�ۅZ���q!� ���a<��
.ױE��I/f�8��K��N�QG�Qm����3i|/Y(@����&�����r`#��g�i���H�)�:��4�<�Q����1�SY��
����(z��|��h!�*InE�2ݎ�!�6�9��Om����Y��]�?켄�Ѣ&�������.�X��<_6���e�ez�%ҁr���4S�fs��=��i��5kM황�O�+��N})t�ى�Zi�� ���6����4����\��{S���/ �lf&7X���C��\#�2�y�#7��:���I��bƌ�c�h�_\�BT>�ТQ\��e�o^Z9�cZ����K�;��t�����+�m�O�1]�0*��؅�2�:�0�ފ[]ژ�V3���|�M��pue讅ݧu��V;�(c�}�0	ж:�,&�EkR+��9�b�]+����`h�(����L!����Ǧ,� D�$��̒>��UO��E�-9����Oކ�}�R���w2IH��Pv��p��Cy��p���]��6%���o���0���4�J�Şi���9	-�l�I.*Z,�'����=V���X=t%��)�<��Iu�<��VRS��F1����蠥h�J����S�����[/ca��8���$v�q��-��ɩ����}/7�Zu���g���[v�eQ�W�-;��	��A��E��e;����,��
���L7�:�*��#"�[�[��N'����d�jR�³C~�N���f�*�G���@���ߺں�'��h3�[bJ���2�]d�]%ƀf���[&tRGGB���W{�WZݼyp���s�������UAY��j�^��?:}Y���\��z�� �G���O0�5����,&~�f�T��Q��oT��[o���:�����s���@S��k\`x@)!�5�wo�ѝ�mS�-r6����dų���%�vВZ�~І�J
�R�>ɨ��Q5�L�h~M1\L��X 	���z��Z&�jں�
ch��|T����b�J�}���=���1e����⷏�X�c������_��n��U��	gr���kȨ]@���r��	� Xaf��
���)��32�`�{�	���c�e�9+ha�R��Ca����h���j��N7�E�$X�1��m�Ә�X��nx|��8�Y��.���S�4�#��)�eiW��y�
������-U��P7���C)����s�D{���2k$?�j�+i��o],�Aˌ�`�+sS�|,F�+^e�?�ܹP(c-�I�w�΃O���H��&��P��cה�݃�I&�y /�2�W���f�^Z	��Ց�0�k�4Z�� 9)��r0wǴؽǅ
@Nu;\�]��ϻ �+�;�o�Y��,��K��Eݹ�pe���)X"v�����\�:���.ۮ��¿z��Y[<�
U3E����9�
N����$6����W� $rt���:$���Rh#_h�T�/����YHy�'z�);mo�z�q���#t����Gx�[��������p��mc_�6���Ǌ�%km��ҢHm�v�3��d�v�� ��q��٣���3o8a�1 ��c��o��{��U��QH0��M$'��Y�Re�?o��q%"�L��nY��d e���A��<g�!p=��&h�sa�E0Пx�<��q�6j.N��c���E�y��P���h�V�j1T��'�012�Ŝ���	t��<W�#ʍQJ�=\�ʐ��6�i����OD���T��Fƣ��m�1
�d%-ϝ���u��}*<'�t
)t�K1TJ"ad	��	��\�Ye��[�g��yHˡ���B�b���;Io��n$���ǔ�, �ww�ᨉ�L��8Ƭ�b�y�;�T��+����s�SЎ ]JXt�UڹU댏��`|UV�hQ��T)g����lZb��Tޣa@��
Ł<F��Aן�9��ĊF-�Ek���=�Z_-���֕$�1���p��Sa�
	2�H[B�}Si��7��dCǙan��� E�}��M�a��/{D���Dg���b�3������|�	£D=���l�
@@c[���68R�%D���~�G��BW�6��eyױ8mHPL; ��}�SmQJ�\���� ��k.��O�n�(�+���}~65E���>*3#����pK�3���7Ȉ}D��FxE���}��R-���6U��WY�9$�F!9$�`����F�[����Ev*K��&c_��n}�d������<j
�:���J1̑�Y�4n,���X�m��)��fOA>�@���fD~2����E�=���!�Ļ>��t.��we1�G��]��!��}���p����<�#�+c{e�$�z|.U'�`����lb�������~$\t�6xF��}��_7�}���zF��*ƿ������'�_.�y��8)��~�5�6�3�<�1q�.�g;���nYh(��wv_
qVwI�o��-�C� �������0���޶l<P�tW��d��R�	Ŗߘ��XAB~�PjzK�v~-
���)��)mGR��vuX_����)�ߒ��BZ� W�Ӌ6�}Q&���,�WH�D�M�����y8�?�E��uǛ+K��ڽ�G_�5��-%<g[�AK�
��sQ.B�k����t�02kv�զ�����Y�4g�h�چ2�m�`g��p{-9�l�3�_��J±�ۣ�HS_���F��Z.�ڈ�׀A���uB�r!^�y���g��.���޻g��S��Κ�# ���^l�ɗ���M����tb۳��� ��s��GW�=�#�� �����o��:�w���ЕK�@�:{V)�FD�f��_B�l{t�܈��g���]q�M`�����c{_���Qt��� ��)j�
��G�s���y����pQu,��GE��gY��S���S��F�8��y�,�M�fQ������Y��):���Bg}x��z�u�T9�Z�(-K @V���m�6q�e�	V:��"I����Ρ������;�+\c��$�C.��N`�!& 
��c�85˰<i��ڄPk���UJ�5	PWoԿ%��Z	24�n��Ov� ����r��OYJ�iu8���2��Q,���BFh0�iYP�F��>-�)���ʥ!����r���>�U�;�N�lQh�H��x��.���p�g��#���^��+2���@2�l�ı��q��G=J=Oy��j蠿�}�N��,�{ѩ�2�0�z���ڡ��@-/c�m9;��,�S���˝�D�ĊK4����	c�e_v��^�OgS#�j����TY�꼔�u|{���RE�*[L�����.�C]f�����(�*5)�)����'A?�`Rv��E;�A��+�=�o�Ju0��S?�or�7��#z��9�󁤤�@�c;R�����8�v��c.wlU8A������ǭ�iA��dr{��8�儰N����1���$s&�g���3Gm�𰈏�8����VM����\��<�4X��̔b8���g��ov��b�E���p�y��)z[�`��Ⱦ:���άl�DJ{�9$�������L�]�&�F{p(��>�X��@��®�������d�-'i���tmܭ�3C��G����<%!~ߨHf��,[rh�{2M���gX�� ����)���_��Rz�Uc���|�)��i`dA7S�P�>�������t`�ԃ��w�@-n����I�<�r}p�p�I[�N�3,�i.N'�Sz�4?���;��%�W�p9!"e���?q��K�1H�&�:�ݜ&�#ԋ���ӹ���Ǌp�0>�b�M��s���C#9/�����Y��~��P|�Ed���e�v]���F�O��K�
d�fB{v�= 6���k�7���H7j{�*@X3a����W1|�-�şK�C"�a��Y��������Ov�Ɯ{7Ηu���--��*��~�h�ۛ��V�o���E�6Th�����54f����DN�/����b��p��c�
��ܢ.$�fh� !J�&�'3�]���g���\�/-4�Ee����߬��-��Ф �b�]��X椝*ߤ0c�����x`��9��6Yn���fw�w�|�po��;	�6�>T�[�캸T�9M�W���G^tT+�X�j�lA�����$Y��o� ��j�n;��20!�'��S��3E�`��M1�`�˿���<�̖���Qq��L�dw`�SB�C�URM/���Ϯ��
xf'�t+��H�n��g�O�ϸ%����MK�}r*7�6Օ8«�Fx�}u��/Z�Z��ެ�U��]�Č%I�� �;h��7��t8{����,4I�����&+�>T9��y1n�sk;��J�;��M�|�Y%�_ź��'wN5z�����}x��U��,.���~�uЂo�,��n�����>���*��ӮIG��e�S�kq����6�h+��ĊC�i3P��aݡ�'��[@�<啼J(%���g�\��\<l�(�V�_]��8���0���Z48�
?d�v�;\�������r�\-R�VO<��gW)�]��Pa��;��1\?mF����N��E+@����2� DRӑn\�n(��N
�E:�x�>'4W��d�D��q�I�v6�dFݐ@�5��+=\$���=)�������>��G��q��<����i���P so����Z%<��a��~`���^t<4C=y7L���)��HK��	G�h�2�Y��6�B��?�w���Z2�q�&�� @���fA��[>y�y&�0%���jG�S@+��F/$�z�Pn��7��#�|�۵�1#H��m��H�">��D>t��6dH+��qu{� {8��N�7���9kUv���2���ˑE-��^�9�(7��[�<��G˪0������S©�s"��Uu���F!���{%Z��Aq��0J/� /�_�
o�=�`rI�#iW�����+I�V3�R������۟�7C�9�m�|f�࿈�;�^t��p�<��'���7�Yh�L���I�[7nW��n����p�������k�)5$��7���wuzM�z�@
�s<x�f�N#���W�@JB�+H��h�,F�hxZK:`
:M�2XN,*��[d^&j���2���{��yx��2P��/JU @[{��-{����Ԁ�@��6[����į�-΁=�\~a���l6G<�#Cs�"�>��h���E.]j���P1T��f@M����#p�W��y�X/U��U���%��H�P2^��|��'�)���lWd��}�}���h�LOF���G#�K�ZqT�*�p�]Kt!�����E��!�����b�qm�<ч�Ƕ�R=��8$��!��e��,���5��7��?���t���(�I	�}��j��x�4g����L���Ę�#<T:��\U���f����g�3A�FF��}ThxR��}����M)N�L�'b��&�6U�7�7�|J:ev)b���j?�;��(�/M�����*�Q���oAkhU���rH���>~���������;-+p�W�&�ޛ̯Z�⚂8���aC�0ljf�V<Gy�����H��%j����%��ۯAn*�Xh��\�Wu��� ��@�ň�!G���U'5MwE���_@��X�Q�P~D��b��58��Y5��{�X�w���9!AR.���T���v ���l��V�m!���}Ǭr�cY��5z�p♝�e#����i����4p�����X� Y�э/_��Z��:X޽��篙�y�Z��Z���)�eq<�k��~�m��f�5��uJT��h���ў�J��7�u�bϘDU���L���r�B6n]�%�UP��M&�Ŭ�t�ŷ%�XB|<�����~Ye�p�K.�����e@���oRA� �lٟ!P΋�FK�K��� T�,�H�y`;=�s��^P��F�����=��/����˧*l�%t_�%$*g�_�[R��A!�.�c��fK
lw����@�\TՌ�����j�*7V��GM^2�΀��2�����2a��E���O;�:*��wY*�6�k�6��	��p-�1�|.�t䠵��EJS�qʯ���.�Lj�p�<\:ad:��I�C���(G3GG}j$H�v�<2PHxEm�o ���`��4�"�I32���;�M��by�"��_���K+z�|��|�L�������@�&@��B���p�M,;�X��S{ֵ��l
�'�u�!Ѳ�'�����קt)�'�W�_�2S�i�n�-E�)���(�Vh}�`N)�\����	��]9���p6���ʔ'���?'�0aWܢ�P<fJ��E !|�T��?Fˬ��k-��-�P�y�aPm�������߻���Ķ~tK>�,��9�/�W����h�\zR/�� i(� ���3u����n>]�QZ��}鴻r�]xgeɫ��W*f�Ц���1t��ɮ���c�``E�����ԩ`84]d�����XG^7��	f�I�m�:�a8j�P�.�D!��Ϗ�1��>��J;a�u%8`\���D��pS8(��s¬T�r4��e��Wwt�V>�@M��02��J6/`}����	XhZ`z�YrD��x��F�5,Ԧ\H�l��:�P�V�V��V'6������h=�����:)�h�v�^m:jd���	C/Bñ[G_�=^cm�S��h"��Eu�Wa��`>e�a ��V\&�Cs�e���n�%��ݺS�s��+�$��kn�k��>�楡��[*��_K	�8$X�VC=��Z��/$q�/�j�BhV<�������ԅE�l©�)�w�B��9��L�����@���tPFU��'̀�sK�;OB���=	�|��*8�t�+�2�3�EK��,�@&آ&����t���ⓥQ���d"ܘ�����{x�CW36t~�v�}4'����n����&�fk�ۜ�t���E6#��`���E3�Nc]�s�0<l]ye����R�nw��J���������N4��P�� ���5+��(Ŗ?��w�`�o$�7�� ��T��V��#���k�Bz$��}���� ;��rj��z���{̞C�LPye_�(��6��E�A����JX�m��b���:�{t?���xB�UgQaa0Y<v����*���f[���Q���a����U�UbU��]�� ��^S��K)�&�2x����[������E�>���ĝ�%f�S�<Z$:��(��k%�΢�}�2�P��d2l�e�/���*ʺ���K��a?��ou$6^JA@ɦD�Gk��|
�AFh���(��]��MH��C����7����h������U
���/p� =8$^�&,���ѭ?�o ;ܝ��֢�����E[yt��z=�O��j����t�S?H�ʟn�IFx���yK��rB,���H���ު?,UFA��9�]Q[�{
&2G�dI�D�����2�im���>�����BO^h�+
�V����*�DI@��?����ԃ�,N~���5шp˾����r��!�϶RL��[���4��q2�.��NI�[��h�Lc��Qr	��otDm�˂�k��?WBi�.����������]0䇛��M�m����7n0#��a��d���phyl+��go���B�>��NMG?��l���JB8�X� g��\T�
��%Jw�r�՞�����A��0�\���kI�`i���3��Z�(=�G��QP��Bh�c�m���cq��8�}߉\�Lh�
Y�!���9o��
9��W�����-�e!�A�Ȑ-���0�F���`p�\���Fzt� q�r�>�����;��"Z�E�)�K�7�s�`G��gAn
�Dy�����9!�6����{��{���7C�1'�@a��A��!�-�+!f*�60�SN�J��g�s-
^�S��ayD{$b�G/q�=Ex"���=��&��c|�e�o��b!�n�	����"#Y���Ê�F>{��;�u��K�g�z߻hys5��UGz0b��2
n�1���`�����7%�X8U��Gv��u�t��;tX��,�;0��]��jXb7��_iLPy ��E�iiĄ�y��ȹ�p<+������;�"z�{PK�CI��A�l�H�-R�R)��
�E�ݜE�↵�dԹ�F'E����6d	i�K�E�I
0���ӇgG��$������!��f�zFIT�^Qf����L�W�y���t��EM�u��^�H�0RC�D��ł�>WP�>��b��t�,�x���x��a�������媉�#�Rx�3�j}k�L�>lHI��л�4�Z���-�}V܌�=l>��I�e�~�����v�3�+�"n��X��u�a� 9ńy�PeB�D��s��ֆS�H������sK�#�|�I�+����۸�����|_ڭ9�$�p���PGM��ڥa�qհ�fj���V�l���gǦCT�C v��h���ހ͇X��p���:�����vp�N_ ����t_��e���r�C�)�eg;�8����M4Ӌ�shYi'Ѡ�O�
f�����A��mc��T/j�#� �O�$i�'a4nݓ��]���,^��M���G'.Q����A�4˻G�nM��0P�<Y����H·�%��_�x���1��_y��%+�V�����w�̳�Ϩ��y��X(�<�䍄�5`Z��ӫ������a�ni��a������vڀ��.��C��>��R�9�7�e[��BN���Dk#}K���'����֚{�<k4^Ҧ#��d�I`�E���H	t�͛�I��{M��<yy��'�I��"3��ځ��Vza�1Ǜ���9H~�W�hS�v��+'n�/�������V�	~�l������*h3��U�4ܪ�n�ؠ;��!~@�0����w�xx=��2RC���P�bi���j���W�Ex��@��?iS_�b��J@��e�3��s��}�$� �D�v(t���$r�_�B/;���8�̢խ�Y���X����I��wuۣLA#��e���4�ǝ�s�S�)q#�o�";�(O�#��!H�:�d�!�m+M�*]�OÙ����&��)�C��I��S|̠٘�ص�nM֙�Z��d:�Ή#�g��4�y�lP��2/;˩&o]�䚃�|�Au*j�)��ȅ3��㻲�x���s�G�Y��!6y�D�-9�Bsx��@c��L���aZ�=�`��U�"�Ct�� ���xV�����t�5�q��������v(�r)w�m�h'�[rJR_�W谻>�h�����Ʃ^A�YS�:])���?9�ց}��F�Y��s�ܠ�n����cj��܊��*kǞ\�XV�]�5�t���$�����\_}z V5Q����}a�C��? (ؿCw��`�p�Ms�	�M݁��z�4�__��F�+��������5N�F�r���6ʵ�63{�����|���}��\Oݲ]��+�#1�� _����uP$�zph� X��+ijC�'�L&���x�(;��Njznd}+9;r&�%r�]�;�0RԠ��ﭒ���O�G�L���det>��ˤ�!qy�H�����$���ʸf50���O�`�(ً����3��]�_�y5F�>��!q�5=ǹ7�n�Rc�%�d�{��lj��_۸�M��OCV.'"7����G� y�(�d#q� �|4v&
�h�{�]UI�j#C_�"�����q��V�:�����?�^�`��k����6��S�ڱ���������r���sW��O,a�>�P��z2Tp�9B�3�?�i�C7`Me?˛�zc�s ����xꎈ� Q�G[��x���`��H��5w�p����H	/�������!�1�I�'�z�����N�9:
�4A�GU&x����4�&��TTpZ�Ď>�h�m�w��:c��l��_-�m?u~�� t�����_�k>L��\� �Ϭ\xm&tnL����F�*�S���p�}gە�8��	�}ȻwU7��$f:�O^7G��}�ۅ� ˽���� �q!�8�И=m/��A�?��?G�u��O�U��(пg�lUx+x��QV#�e�O����5���8'�'q��.Ku��].E�,6���������[�n]0x��P"�ʦz�v3u��G}Du����h�6~LTD�/\��37��'��ϥ;X
���c-㔕LB*��)I��4��a;l.��!t�#�$y���_���)��R�uW�n@������R�$�ٵF���t���8[U��(9;T�0���I&T��/� 営cZ�W�]r����ctW�Z(+��#�&ڙ���	]H'�ݥ r����M,j��RB��%�P���h�Rd`���=&����W�I�_�7���0�g:R����1�ǉ��}����d4P��]uEȹ�'Ŀ�9�?}���2ߑ�cO��a,��k���L�`kTT�'�H��}}T؏=p���!�Y'��T+)01�+ D�y;���v�����<�0��P�2�W���w�;�W��z/++��Yk�d�ݢ%����S������+ӒNw�oQz�ʁ����Z���PX~Y���_X��
��L��<mu%��}䲞M�2Dr��N�OiE	���0�B������--��Odb�}�6�����T���b�]���mO>T�_�F��38��gE+ߋ��7�	�!�������E��e��U�l�F��qa������l6��.�$Cm#
C�{���;VV�z�%-eN��x��cӰ,d��c���V+�#�jУ�Ozv�=�fb9]I<����
��q�NM��9��xI��_�q�ˏwz��D��Fh�/����R=�30?��bK�#�)�3W��3���v�X]��2>z���E�`�%��5����v]YLK��V�F�9������V,��#���P	^�	@3�I�����;s��4R��$Q�X~a��'c>��z0c+A'U�C.D�3�����40\C��-*{s|y�L�F�~~"ᫍ�Ǌ�y*H���猬WCޗe5�:�����}�ki��~��[/���������f��S�#�Z�
�~MysO�1=Xg�Ɵ�v:Ó �G�}Q��,�m���bx�m]Z]��XÒ���Ϛ	���<�.7��ҹ�\N��f E�&��+lg���8Oz_�w	�ݮ�^��o�
��x?�۴D?��[�֞��.HS���n2M�oOL��A�ysG�O_B�����<d���i}{#0�}��L���X��Į�FʩI�#�2B�1���*�ׇ�j��+�7�t*q5��{��C4:5�yg��)>g��X�G]�T��<����P��G-\ �"���Ήͣ� �z�J��ʣ��A'#9%�埝��J��TRV|ǈ�Mx�O���4��?��^%����8}�ITp�(�g���dɕ�C�.�4�<O��]'�����|f�31ޥ�8�<�� �<��,�&{7�Y%o�g;�-�7���w���Q�;09Q'~���x9wSt������0r������9T�Z����(%>��\�7rP"9A�Q����Q=�ʈd��ϧ*:P&H�癑$zD5ۛ������A٨��_�2�V0����#��TɐD5ϯ<�i� �v�5���{�)E)�^��!]�P��}&�H6M<�cA?�"���S!��%�Q�Zc�I��H�46����Ʀ\%�~(�o#%��
B��8�rSB��/D*O9�$�Mi���ގR!���0vI*�OcDF�@^��&	�ҧ^G�B� (�}DB�k'����ے�eq*�*&ڻY��L�lZ���-N�{p*����\����ћl\
�O�e������$��HuŊ����=��L��<}'�}p��Ђ�`�bo����8�^��L��^�f�.)�_��hU׼�T�/�:�E���j*�XgDb�]���m�˄sRk�f�C�>+�\��-��k��ѯ�L���E�� �,���S���?,�"�Lm%�_���c�g~ ��[:.x &�I��OQ�*�+�J��m&S�d)�R�J�'�/StQC@n)ߥ�������a�Y��Sd}I<�3�?�9��Q��-kǡ.N{z���L}�O6��
�	��M������y��Ɉm�t~\�J��yš�.Q۽O�����]�=H��4o;^Z;}ǿd�6�~��k ������':��0Dhج-�(�ǋ���ъ�p������O��-[����]ay��nFz,T<������a�8�w�t{�JH�UA�e�f}Z���z�S���0�a`�s���s��L���;풨N�Al�O��_�T%}����"247�\�e��Cc�LS
Mz��� �?R�3/:��Eڇ��d>J^W����D�����CI������U#�ɛ!,�Isp��!�G��<~�;����i�����D�6�/8��):��f���� ��y�gb�#����O��Ѧ���wA��N� �������	�5��c��-�"�iZ�=\f����*#���mz<q�ƹ�%d�a�HXK�������$�`��2K��й���������C&to�:٥[��#���}�B!����� ��ף4��u����]�5��܈��Bg`^�������wrN�E�����.�50�q1����W����a/�Xf.ꛠ�7çi5��#>צJS��Iit��`.մ�-F/��r�i+�:�	)��6�s;�ƓOG���-Y&�*��4ʦwQG�3@�V���x�0nU��Q���d��n��K^�U�/�n��������d(�vS*#�c��^㇃~�)cήe}\�A:�E�h�ur�j�2�js{�	o���"�k�v���l���������g6�+) ��q��"�<߇H�?=�i�����~��^��M�^-�!�<��=�:4�'��[�X��9Y?ьX��sQ)�{�68JE��~*p�1ٿ �Fx��i�,K�B��,�KI���5\��v"R\�e-�����a+p�ȩ��S���%�\#�<�|%��Z�,>X7�
WN�S�l��j(�Z="���BW�&���IR����2�"��a%; �a.���D_�ޛ.Y(��l�ޮ"��BY�JaZ&�)4Zxߠ���h�@(�]��N�Y�>����dDbW=�Rx [K�-� 
�u���^�@����5ԶX��@�?��~��{��x.����~X�a�s�F��y�t��<`\v�t����TM|<�A�j�B�U�W/đ�*��Fz��@wq���Z�P����dL��+2Ѹ		;�v{0�w�����V�a�Xȩ��u
��=m�_���v�'��o����s�O",��9�� �7'�#��
��G0;Ģ[1�lJk�r����t�󇊱����7��1�+�Ȣ��g.� ����yxQ����h|�Q�;��Z��l�{^8a�D+�5��㇋�m�gL~q��+zb�-�80���宸�,��+�V�Ҍ��٤��{�r�	���}�c���CoVA�~Ъi�wz����m��L�7gT����Ř� �}��q��z$��v��e@�$!�1TN>�������o��"���SU ˚�L>��h~8���ure�Z��O�=�nI���E��y3�yO~�)��;�\�p�����D��?�f~�9'�������^#͎�:�m���MT6���3-p�ʩ���(�A�C��_4)�8�u��)�:��k���l0�j`B��	r�Φ��?�v����M�*��^�J�t��`��<�K�#��od�t�G���u*/n���
��9��>�rf��?��o��]�l6@"��nP��p�xɲDK
���u�p��c��!x�k��������þC�e�X��v��^|��_Hb��%r�.�����%2̮^]�}B��P;�8��|������]����C5)m6��e��p-Dl6#iO]�r8;-\�@�o1O%�jA���PP���sv�Yl@���bm�(0���V{D�6[^<��s�g�a�(muf���p���w_�RW-���˪�_(I:wQ�d�q
 �$RO/.�N��f�B!B>�	�_-H[*�*	\"x��B�v=�m(�sxK����	����E�n��-��țAD8��J�ǒ���!C���f�U����B_}N�@}��� �O���F�ߖ�P��.{�Ԃ<����t;�I{�;��PG�T�aE���wR.���,��V������^"�0[�[�.��5�fE���\iЊY����͔-��80���_%A�3�؝�MaMH��@do?2�-��;��ߦd���i7<w���.��������C��Stޫ��@�W>���W������g��ԙ�'�$��� DS޳7Le�M��aѾ4 S�q�����I<����7���v-1������V�˅V/�mߩ[�]]Ld��E-��Ooœ�N���1�8���̢�
�q�Hc�������,I�� `l$����T��d�C�wI��@�H�V{��q��YM?����rݶh�mՇ��r�m9dK_BGž]��9�X��H.�Wl��i����Ьz1,� ƻ�Ua^���,$������%8y����B��6���1����'�(=X���r{z/V�Gel������Rn=�F[�t+�����Ԛ����L�k�/��G�<YP]�dF!"��;(�*גlX�3�f��d�r�<06���T��Ղ>
�oH=�E�b��b�$�(,%�3d�~��\�����g�Cv����V�K&X�~&���؊f�?���[]�ޖ}�0�>A��4\)P�CBpfOEf0���v�M2@M���������ա{{��~�#��[&g�ʫxyb��nI�s��|�K�C�Jl)ʵ�iA�d�P�FSS��rM�U��cC�9���-wN�nl\�=Fp�0�����8�<�~V���H�^�6�߶�� ?~g�qx�8tK�L���[+ُ�5����Q�gH��	d��q�#��GV�12�!�/z!�z98[����E
����-���������M#���ȑZl�x��|'������R����hn��J�Zj��e�[AC��&�a�+,�Z8��%F%T��� 0�� ��n���vI�ϵ�OH"�/���PiA(��G�u�;���8����-��ά��Hϧ��{�.�j�,�D�K�Bm{��X���a�9v�	F�I�	9WE�2Ռ��l�cj =�V�<�jD�$n�qL������*��}'���ܾm�x�G����	�='F��Z��B;�^%�͞�S��l�C6f���ԋc�[�(Гѐu�7nj���Ћ�0(��c���)؋�;�27�����yK�>��6��*�6����:>�_�=uii4��ϣ���ա]|pA��8I���OL�G�κW��fH z�-��/<g�"�Y���;���_Pvc���uiIm��N�Cv�=��z��տy��7��rf�<[J�х�|�۵���%x�p�]���$Ϭ1�Zh_XE	��ڇ�ח�w�'s�e�H @�ՙU�k&I7[��U�bӴ�6�h(++�@[\���Q���|H&��F���a~F/�q3��Ta��򁌠�U�
�y]�� �'���� !_L�v�U�	}9��Cu�"*�����1�mc�!��I� ?�H�<Qrq0�A=9<6��9Z�Z1Ȅ��2y�HC� ƸG�A_����.,�@�R��ɐwv[k���c;�b=�� �}Y�b°M�хq΋���Ăp4��>�r}�0����(�l��g󝩧�؜�V����7pz �:�ݚ-ɠ�%��H��T5�����D�<�� qq��߮M�w�[��n�F�\1Pg�V���
?�'�h�$���E9y����Q��b+������ /?Θ��\���iB p���,�~�V�H0L�S�h���  �����:������]�;{�B��5��|A��_j0f�2���w��LA�u9�O]g��)A�>��y��	e��E������#<c�0'?�$��Yj"�uF�\}��%�As���n-Ķ�z��Ms��C[_K��Qk�g"�����a{��l�ء�H������>�n8�DB	�h�kS��fj���W#tb��ӥ�L��Q���$9>�r�s(���c��
��ڱ�F��c�/����M%�B/ԇ�K�h����}s'6��B}�D�MWx:�Uk�æ�F��݉>�n����!MNs�����CGcGBx#V"�/m���sh6�8�G"7���5:'i�u.��P?��:�T���W5���42�:2�1m�~]���H�Ǐ���u���l������ Z��j殩|�G.�x��,U'���5��gkL��4yJG������ȿT9�������������F�j/y����K�^�0�3�l�ψ�Mؐ���x}��4e$�D��L(�_
%�$r�
�����R�=�q���(�U�4�z�;���&7�ϑ�2����7Y�`����kH�o�{!-/�oǚzU�,3����my����Α$��7b�7Ίjc~B�и� JÑt�[�i�L������&cM�yY���K\,"U9��uG��I.ɶ��.��/�
�l�Fj��6��Φ/R�������S�[˨�6��2��L\�H�Kk%$���5����})Z+�;���c�xqxm����~zP�r�egk�ޟU�p
ZS�!%;�zZ �c�SV%�O;��,Y7��9߫�p��	]�nz�t(׿���S�����<}V�������ֽs�P6-�X?B�Y�������y�:[Șr�Ew�9��FǱH:GOd�;��Y�,\`x�g:�d��$Pq���(9Ŷ�e ��M����Q�Y�9�}�W��H�@����I��#	��/=-�91�����Ą�Y�Q�n޾h�@s��Xgbs����
���_�VK{�~2��A~�+��SD����I�d;�^��h�J"�1���)� ���*�; �M>s�{n��@�lU��r�o.I����Dd`=���H�z��׷1z�g͍��6:%�	i�^)�mA:+�J�p���2b��|�`����������$��y�V���Hf���LM9U�QoM�m�z�[�V�ݺN���;����q���m�>��\_�3!?{�ӻ��@���>W��L{�HE7H���퐵�`��Wce�)@{�
n~���y���|�ٴ4|��*�T* �`슰��':�{��/����m, 6�b<R�8��b�%o�k�F0v��J�-�z���$9����q�{��JgY9���C��|�$V�ȭGo�~Hx>&�-�8��޾FS"K��/[�Z���Q��A���<I&�·oV�Ҋ�; y(�?�%��L��=�p�l��c�����Gj�Zl9�x;�_�C�3R0��R�N��Z̠�(�H��m�Sw�}�8<���E�N$�m��H̪A�V��DԥQX��s��a,�u�?�% ƈ���U�`��h�:E���1B/��H�ڧ�w:��hM�Q�dc�p�'��m� ]��{L-w�}o�&�ˑ��WZ.��(�E�vϕ��4�o^@x�}ٔ��5�3��	z���/Pi9M=<z۝��� �w�A"雾�T�V�5/��݇M�<3Y߁����kU�U�ʲ��U�%xSp#��	���Ɂ��{\7��c}�X��%���l�_��b�
��.�>�������oN��mCL[�F����/�����D�ZM����Ϋ�}��Ӌ� ���e~�E=]�|--`;-~-�5#	�J��,�g�{?��nTY�i�ϵa{�t8L��	vV��\��g,�?e9@���v�l������cg�1]���#�J�7N�f�K� ?!'c AN�\a�#A
_M��o�+��D�K�Ѥ��%��9�s��]���8��:�A�h1lW��ra��V�:��b�0C*�\l��t~��Q�Z6�$��9vW�L�ŝ��q�q�s���Gө3m}lv�Z��o�D�A�S�5���탕�o	�������[�߱p�z{~�\��<ĩ��~��-�ŕ���)*J��������ס֩��iB�BCS]D~�7V���	@���S���5̠��Hץt�B� ts��1O�ֵ�]	�um��
,Ã�Ѳ�eW��]�a�f���5B�9|�.���;�����݅�M��3��W�
�k��/��$�\���W�
�ng�.�aa�m��d�,�SI��t�"��41K�`0�Z�d���T�{�=,��[C5�'f������%��O���F�;
ݩM"2ʟ�JC�s�����-c�|�d)�H���:m�C�J��t!޳�&{�!q^�Jlt��񾦠 +��	��1�k����oFG/���?�/`C-���	ϫ��dp��"})s�Irm�㉑�v�ܺ���{��4��n�v�
�rJ(���QM�NP�.'<r]6�	j����y?�x�V-y�j2���s̞��֣u�s7>��49�Ӹ�X��l�D�a2c�k���w�:�y��ۮ3W�q��G�e����e�ئ�r����19�t3z`U����$����x���D7iH�u�S������.x�ܱ��
p����uJ�̢�2u���L&_��9-�a���P����
k��xn�h�i2n+�%��G�Ja��J���0Xҥج`1���9����󼲰�;��xdL�C��|R2�"�|G�Ӧh�&�ijy�BF�f�(��έ��`4k�$dJ�<C�� �41�}�-���+���17���������[�atq��z���7!	>ǫg Mq� �ޜG�0��S=$v�z5G����	Y�]\�Y�u[P��4��5+�Wr�x��)�M�"��Mb)M9�
%�u�Ȟ6V�m7���~�6q�f�
�>�m���6�~��HH�iŒ�����b��ɍC�g��Q���|���{��~�ٜ��2Ku�w�R �׬���{�n��2���0=�dc]�nn|ծJ�����/�s�8�Y�a���B���.Ch��m�l��1}7��oO�iA>�w�j/��0Θ�|��y|�g�#i.O��e��*b6����!�-���B��҃V^��� �J	88���%��	̌F�cIYB�__��i��ҡOVx(A>1�q
;�&9�ҫ��({���R��p�w��?\"-��R���T2�S�WkͰ���/�����VI���pA:]�UN@\��[��5�Rj%B�MI��%��}�P%�V>Q����u�lX�Y<�"~�Ĵ��*G	@7DSԽzZ�L0�nl�����[�`���'��H�؀�6�Zu0㇅d����}�G
��Pn����E�gi��X��~K�|�RN�ٸ���Β$���)�7jM�~=Jcr��d��bUJXE�[�*r����C�$&����v�Z��Hѹu3��\�t�'���L�����q��1G*N�R	]����rC�]� �> +<�d�b��-���GOK�Edx`���6bM�M"����vu����o��\TOI����{�U��bc���&�u�J�&Ct@1,d?{B7���������aJ�"��Fw��������|��/o�>Nx{�2p���������i"��|6�d���"R�8<�ȕ$����c���"$2�y�}w��6v��y��(I�M���dh��+<�'��^���oJm�2<���"��
�)��3yD�-!a���~ʉnMJ}�A���le/ i���7Mi�9I^#]��!�UE�Go�dpB���M�I����V	X3Qh���6!�f������DRe�,��\�/���:W�eE����%�|���Y����V.`��"*�䕫0"9L��fW�|��Q,Kh�[��GV��� `G_?νE
a��G1=n��14��zqGgAA��-���5��l2�a���_�% \�ߐ��6�����${��u���yl͔Tw!xG�&N�\.�k��!'�=�x3��v��X�_��V����4.˚�3�CHIg��RQ[�f`q��,u���o)�\ܮe��KGf �
�B��[9b��o�w��o�4wi���BM��ü�Њ�ۦ���&Û[t�-.�QW�����Hw��`)����w�M�h�x]Ԏ��i�ҶF��o]��)�˵Z&[��#Nu�s6�G�Qt0�E{`|\E�,/��.Pq@+orS�t2�(��k_A]�55A�I�����k� k��'�T��_=0�ɂ�V{��Q{Fp�7��;��= 	2.��a�^Oe<�[}#{�sE�74:�mtl�dS=glz�I�It�+�ų�8 ��x��&P�h-�C��"p�<ܯg3b��1�b�e)B�85]��cK�}����Ь]�� �@�n�l�-3�^��V����:�k��o���}i�SXE.�RIE��k�$��ASbp�J��rO`Bg3�*�[۰�q8��?�YN*��7�[d�I�B~y���Z��y��iohh�sGL|dq��t���Fj����lb�Z�$�XhOW�EWzg,��V h�ȵ�K��/A�TI =@ݍ�Ρ��Fbw8��҈[����lh�/�5��̵���H� ���z���8/q�c�x)��7q���Y�+4��{s�a�lf�aƾ����3���4���E�ۍߛ���g���ɯ�rk�f@��/�L8͔"��Rp �ޛ+'.�6��7��XAJ�7SŤ���M�P�ނ�:�k	9����*�t�����Z\D�@�v�氎�1C��Ƞ�F�C�#�+�mBo�&)�y6rDwT@βx��,|�\yՆݿ	B������wfϡ,x��!1��UA�י>Ч�PՑ7O?�~r�x[�y�+lͬ�b�l��R��t+����\��F�,���ܼ�9{��25�:q��d�F�2�PT
�8����P0�mf��x��8���bt�0�$�5D(������`~�)��WFS4�HE��a��kJ�������΍UG
^c��L��|��O�o�)6~�&�ޕ�mD�y�X�sk��3�ٸK�ށn=":1�x��C��FF�4L]"���8}��f����z�-Ʀ!.s{KZ�sx�l� b���j�7L9=f�gqvѰ�M<������<���(4�B��K4B�aq�]V},y4��X����c��� ʩN�7�����>MJYI ��L:bph��hAI��^�0�uC>#���n) ��K��\����r>��?PV���y���D!�8p��֐�C��;N����1d���^�����X�#�$���{ݻ�:����;�tR֩�� �ܓU������T�U��\����My"^�/a�Z��M�X\������\��WA�#M����z�꫶*9Ű���y��t��/��;�k���(��[Qw�)�O�Pٴ]}� 9K$$I���B��bLo�\�WVc����:36�2qEF	���i=��'�މ�"_v1t}�ir��s���=�C��y�㮜��[��R5�+�xZ��Ð ��+{�����H��sJ{�Xpp�!�R������R��	q�ߋ]���p!��D������"'6����m��k_W_�� U��YLbM����#�/%��vN�@�c�v�Ҷ�����r��PeeXz�ܲF'��dj8��˼�/�ty�~�L��"���y$�o�ov�3,@�3�3q/��[�ig�:�i'�b�{�p�q3�f9�p�j��·�^�����V	<�l@��p�E���'�������X����_W�(��3V�k�;�4�>�!!���Ǆia��Do~����u�#��$k�ӽE���^!)�BL�F	���EIM����@��e���������nN���Π���)w���'�n"�����X�6��NM�	 8]/�yٸw�٠A&�}��h!�5�&��n�k&Fb�%���l�8kD�����sO9)U��'�}��1�{l��f|��;�r|`^u[,�Ծ����-5TL)�3C�����Ư�p>}⏄D�3p(���ʏ���[�Q�.\8�˒��C>�i��i��w�C�$��R���I/����N9��@K]�&����t�jz�>���!�#� �h�l0��M�J��Ec�2SB�Զ,�B4"[/I��_�Ht���]��y�;�S'+j褗
�37��L����=⦣ҙXmZ�1t��[����(���1Ң�����(2I��
��{R�<�F�&t�D���l�r�D�l��O�[�l��b��ԱXoXB9#h3���|���OR;
X��wG�z$=w�<%p�؁�����>>�W/C�ʏ#�,��$9t���L�g�b�f���K�E�!Д�1���L8;c +�����{\���Y�����VXI�bn��= K�.�q}�9x��RH���j�'��D�g	GU,}�9	Ҕc5��M�pqC�ӂ�ОwP�\ّ᪥���e�o}Y�/Hj����9�a|8N˂Bu�=�1���`z�I�j��uP��al�6��+�۾�$w'���+�U�g�}�J�\��	N�}K�	6�i15��8
�LU���e�Q ��>
�Ï���or.dn:}��TI�OLu�6�P�~?����׼e�D}XU[��������xE�=H��3�B�.� YjV����ܑY_���r��἞:�ID{ƚ`��+R�A�ʜ����%Lc*ޘ��A?��U��܇z)��&�'��{�Y�R��Z�!C�����7�q{���p��oSi��q�����O��;�9<�z�k{l ��Wl8,E����+;�)^�.K�G[Y�Rr�V/i
7�]�F+v��
�/hVf�����406՜P�t�*>�a��~4��������릊�vP2O���B�A���8���+��yIg ����f��� ���S^�)I�8X>^���������~r�-M?oe��ն;du�f�Jn�@{Ƣb��zA�"Z�]�²ц�[�f��z�ꫧ�|H���4��U�4*I�A���bA^+~F�};xT~�n� �^�H7�C�N��c��C���fË4
��$��^ �Ά�K�bM�N�>n��X/������T]��� ������ؐ��7��8h��%���i\M�1�W�Y~h�f�<��M�'HꝮ&�����ޫ׫V��Y@���9Χo$�utK�t��v��
��J4-?˳��-�H�B�>�?~�9D?l��;�s�̑3pU(��N�O0r��L�z%^�/�Mn ���ތ�=s� S����|��F.�&(@��b2$��|���1�ʹ[g|���'a��$��4y{p	"��I�f��곸�J��{�4���H�~Nj{�����@n��n�?A����Ֆ ��R�;iDmR�1k8��0�`�i D�M��P��@�]9RRh}d��ʴh��M��N�qcM�uX��Wvq��0N��	yU�nH�Bn�X�O�n�����3��~CR9�5hU�n�ؿ��X��R���.>{Ɲ/^�I�P�\֓=�)<a��;7�`��պ�B���-��_M���IY����%7fU5KL��/�����E�������#	�ѱ��s�3Tb�Awc{wq����y�d�Y�l��Ǎ��}i-鰌j��=_I�^���4��%[5�����}_x�?�y����"�c�n��i ?���(Í�IO36�jK��0x�(54u����X�Z)�6]�[z|�n���;c��]=5�+rK�D������Dzh����9 kV������h�=�P9�27Ɯ��{��Z׫>t�O�ƨO.�K��s>/��{����ڜ���6�B�O/I5ƴ[�7�x���w�'�xC�z�&>ꩴ���v�u�#�(���8�J6'ՙ���Z³+v� �*��NI�]�@�̙�O��\Ii�;��Q��|�0�H���X9��&��h)���2��5�D"_�T���%�~$�< ��8�j@Hu�$�@���]�l/a��~R0��Z:��q	�A9	��0cy�}���;b���"n�]6��)��,Vڎjy�|&�hx�@�p����[>�N�D�h��� `���M
<=�GĢ��}&���k�2xΎ�[�����d�Wĥ�����QeL�|� �3*,�s(�=n��N�Z�!B����찰j֥�B��pC�g�fo��G {f�;RN��L���bۼ��b���
{{����|���#�+������l�xG�"TJ�/�"�&�U�%�z�0k��)؉5qn\Ս�����,4�{n��8t�>�5��m�����[CѺ�����Ǆ���#Afu��:��;@���)��
�.Y�--m�{��/�]Y3��nU��<=$J�;"Դ)CJ���C!��N����M)���6���mI�<n=���#����m�F�]õ?L,���5v�K7/f�(��l��b��V�����//�qޝ�+��m�gǃ�_���EHo�x�7fr����y������C7�_K������u;+2O/x��Gn���.�h?Ol_UkyA�x�5�9Lݣ�&%M�V|��VH(>e�V��"~MѲ�b��c���Ż��g��t&�H�~er*ߝ�7)�K�ґ@�
��<p���'�n�{ArQt��])�9ެ�Ė�1C}[��Uz�9v<�H�6��q����^����UO�I�>E�U�іތ���/T��+�X� 3��n�+����SA�.��c����-[�zʭ`]D:���1�u�<�?!k���kN�K2id� cM"s��pRV���WGOڠ#�fc��X�]���3�M��54��~] ��gv6��JbQE��'�~Cf-O�D�\��]��	ܫ�]��E䠅�w�a��S�ɐ�ҍ�cĘ�݋�x�D��ٖ����	=7����v�}UUv��@'�8�;��WȮ9���#ف;x���������ђ!��^����챷�����aI�$��KW�!3r�r�Ⳓ��X�+h'���S��B�^�Pܧm��<q��������c��ȿ��W�/�ӷ\o���:
s�`�d#S1�oz�#<�|E�W}߂�	�Ҁ�J �[�Ĕ-���h]����=��I�Ė����[�ο �x���@�,)�;�y �D]�cF��k\`�����5%ט�U��Mq�f�G�3G�af����+�����g
�бbB"�M�W/�.up�Uˇa8
�2}&Li�?��Hk�-$��ڿ�	n���o_ŦR�S�m�ﳸOx.]�_ϒx��� �@DcM~�Ps�j2�2��Yu�x����P~r1lO����.���xPqi�%�_X��B�G��5Y���u)0 �k������j�z��	H�p�$6�R�j����J�f"�}�o��}�2��M5�w��Q���t�[Mf�5C����0�^>x9�	���mo�U�;Blj�ȳȲkd�6O�y������p(�f�q��VP'�e:�%Ǭ&�)|�ID�1}��/c��"�:�<ͽY3�?����׶��)��8,{)=J�~,�[����A>aAoU>��CH������p�t�0��UTܗ����Ұ�WD+|<�
�d3�8�:[��C����!#B��D{���wI��s�G 3H�������%�ӧW۵����ᰊ�j-���SR��Ҥ�V�J�����w���������qc�s�%�Ƴs@D���*�p
��a�����vx���Qr�m�'�'��)b��k�ZE��x�%�r1b�}#b��.�{�mBԊ�$�����jA���M;fRPzڋ��.�t
�Ej�2u��E��˩�	��a�R,B�J;��F��:2��ϼ�̙E#lͬd��#T��4�{���m&ʟi4U5�:q���@߈�$?�1���^F���]�/�$���C��+��{�4S�����Q����y=�m�D�,ARx�z8�N�f���G��2XB�L�'Hv�0Ī'(��t�~X%��r�ө=�p���>���4��~!9v�K�0\-ns���J�z�n	�sY�]W����$5ޔ�ZY�i��Q�YN�5k�a���cw����DV�6U�FmCn���)�����z�"�0h=��}zu|C^���qR�qLQ�*L��#��'M0B�I-ѿ�*��(F:�n0��D���%�^En�oe)� -m]Cц�!�d�/��
�t�9�D���7D�(�d{�Q�~�d���7���0�-�m,N�
A��F(}�;��²���Sk��Uc�1=�V`�:�˟x�\�6�v[���k@��̧��JE������J�����3߮�Y<&�93���?n�z�G����ۨN���`�<���G7�r��q�Jꨐzy����d�o?����%�o��\(��oor�P��	K����E�b ��YZ���.�]}��5S1�y�!��1,������Ż8� T!�y�b��5�F���f��P�r���j�(?�v��4���ي<��fp*�9C/r*�s��t�i`2�S��H�t3R��t�k��y�x��	*#g9�Lr�'�塒Ox]x��kdT�����\X�~�&�G�k��%��	�MI��$L���`�����7���w�ߧ����a���6O�C���_}h,I��Ν� ��S��}��\5^��*�$MB��W�k%X����ևvbl���+���/?�X�'������.WCܴP��2�<�:��ѳ��:��^�9���ֽ7^�X۹i�6@u�녔��oLC����@���sȺ���R��m�&�[��-+��l8[e���U�
xnG�el<��)���~��#�H:�fx­��F���*�"t�'�G+:4N�hyBS�N;��=��ʈ3�k����+ޜ���*�aj��HH�LE�;��GY�|��G�����d��'���HPb)�E�z�$u�VB!���$宷XU�r<"�3N���A�Y��ߜ淮��Ղ���zf�h��(��*��,�ّ�!jL�шz�j��m];�,��4���[��H����$�F-奞��x �F��T;�ܻ���L"G���(j�-
O	��@�Z��]�D���)�����zʩl�q��C�(��>�M�a�^q9،��LYk~t<���;��9u~�'7RW�W��� _iN�a7�|y8��8z �ϋ�p���*t���o�78�oOuDdՍ���54U�-\��2�EnJ6�[��v���n��`?z!r�;M⃬oC��ky
�'���m�������h��5��c#�pS�X�Lˁ!����VϚ\�L�jb���ubj�$�@g0CR^��H5���3��1T�>�B�����2�d0$�d]�F"����L��DZ��ě�u��*sE�l�D9�e�#^u�tܻ���d��%���&�6��A�(<�������״�<����k�F�Ʃ1��Fd��w��ܴ ��D��k;F���	Q{I$� �͓�:�w;t[�ޑ�hEr��	����ug���I��ez	==݆7A���O����Ѹ��?\�6_��9����T~S'j�vcw���Hj0tr��S{X���cy,
;�t���Ƨ���u�OZ�d���W!��C�+)
%����Vn%�DV{so'�ӧ�N"����6S�*��|[���3�<D���|��I��&;�T�����;k�+���p�;m)� L	ʇ,�!��8R�5��,���>;�h�I�[$��h��n<t1o�!)�I.e|�E
���>:Tp�X�)�N�`�t�ļ��	DKۖ a��.G���ߍMO�h�=��l�+A��b��P�v�9�3�J#�Đ�/��$�),�>r�1<�{Dc;jO�1F����<����Iw�PD�&)�W�ƌ�v~�A�
(��ۯ��?��țƜ]	%8Az�dnT����+��3�	���:,���l2�?G���w��7����ڑRD�;��W5������r-3 @f���bIh���ǖ�@����O�̆$މfY�s
����d�GLP_(e����SE/�ȟ�X��L� I��gk�$�O��Aޱ�����z����@U)N���g��wq"� yךu�|M��E���yc[O��
5�;_�����5�����%��&1ʱ��n*.�Gw4�T�Κ#��zu*�5�]=@��A���v�������j��f��?Q]�-4�o3����-X�4h�b�H�M�bK���[�n|�tbrK�2 OFҠ�嬳�����C� T3u^I�:=	E�O�b��y�����	��������� ��o�:�f�v�y�&�����{�sk���{;�t�zw��I�||��~k�\�]�]&(&�ċ ,����%�f���"4���<S;"�_��&E���o�eج�J�ix��`���ezs7�R*[����9 �-����4+�,�m�����x&*�'�J��}�p�w�p��Q�$���;�f㧉��IL��H�7��dQ�+�js]��zG��E̺{�,�6fF�+�ٝZj0�[xfM��6�E�_}~5;I@�v��,	��N��r�]t�0�4���_�C��A���bS3$<�"���t���~[t>��mB*����K��<rU�+��A�7��
&�x~�]*T�ELH�����XY����7� @E�s�7{dCX��	F88���X9�y�E�Fi��BS��St�R�S;�H�/�lk�>� w@�Pxԭw�+���C��O����g�,�~����	>��EQ�o�f[<�[�ts�����R��0�a�g%�>��f'�	o��Z�
ׂ(�ec�������s�+�_�Zfd^Ud��`qfb�	t�Z��P�����Q�-]���C�o��rN��w�=D�N���cLk,�i���4GϵZ�m̫�ډ�Zo��͜�ޣ� ����!"�T.KN�`1��D� N���;ßE$1��j�ܯ\������P���QX�/>�,l[�*l�:��$��N�{�� t�h_u+y����j@�W��'vVc�����`܎�p�6|f��^��m��r� �!��I��6#����+w�q�e��(���fF��>���m�Ƥ��8�C37�wVWa��l��R�9Д4���E�u�Ô��i�WJ� ;�ry�6Q��)�K�?�@rf��e:V|
̂ ����v�Z�+�j��k�E*����'���֟�e��)�ZJ���c!ʷ��y�4���`��B�p*V�.�5�S��p�hQ��D��bJ�\R��^�F�{���]�_�� �f�� ���b�
�$�"� p��m�4��(#x��b�쒦z߹Ei�8���%o#����&�&E3�������,ve�H���%͊)�~�=Wk��aGp�(<��N��f�{�`�����tE����2�ޔ��PW ]gy�7 #��t�HWW)r{�;�3�;WߙPTB�=�d�~z�r������w�Q�nfQ����crS����<yz}޷S��6��J\��~#���e|zj!��",x���?���=�e�1�����F�c����s'�$lXb��#2 d7�?���
�d�D��r7Q����ZSl�Q����4�o��"���׾J'�i	PS�	�i���ۏ;�9�_1���������,��\��C��*�V�~jJ����A��+ןդ���Z	o�O�����:�D6�42D*ʤ�\�Z�����P �>�?����#��e� B(����.R���	pU��l?�Z ���R���Ũ��e�3D���1	l&�x(��ь�X�"�%g�ǩ�4,��O�7}0N�G@Y.E�rr9"�ldkk�yq���6`���(�s�,h+%J��_��c�O{�w͈��ռs�_�>�|�l~iU�i�F/���pJ{ g�0��f��#3\g�t ~���bM39(y�:�|���t'焇����%�m-�$�0��w�/�s%���m�o}���u��\a�q�$�ק�ҬD����'$6��.���$P-W���P��"�8ד�]`r���^���SF0�0�{�l�^`엀B���s�Ҿ,��3Tޱ�j���9&���B����A� �l�J!����j�~G�P��zcf��:%ǰaȁM��T�}����N�"u�8NAR��A�G'y���՗5�˧�<dC3A�}9	��. K!+#C�=���o����{����T�d��@�~��&yT�'��ޗ��\��$iD��ҹ 3�ȁ���ú`8�&����-{� X.}��R��x a<��&�t��?k�t������Qm����1c�O�0x٪�R�U����qZ+2�_��O8vScSË��a��
;�7&�a���3Ŋ��+��7�"�0n~�(�4z���r�z"p
� ���v5�a��3��A��u.��8��"�ѷ4�Bvfӵ �D��%��:����G��l���e{�ܤ�5���ݗ̥�e�|4�����A.� ��L��G�VFҝ��Π�J�%6y��yK�"���d�!�$���E`�H!��6�))���>u�����-ċ�\Zt�Ж)B㛄)%�n�{+Ů2�o-BLP�`�̾-��^��׋p�\��E��q�S�0
m���6� ���6���̝�E����$��Дz%�� (��Y	�|�3���UȤ�n�4༅���L�|n!�z���4AН�>��\�]�ǳ���y��9���6�OD��@�K�"�zӂw>FU��� |(V� ���:^��m�A%l1��B���Y�:z=��/i�߂ǉ^��?H�C{҅ϑ��Ɩ���*�d5�^Y�qKa�@^����X�	`i~�@��b���P%"�L�Dg�2���Em��by�����D1�ߦ�[ݧc�&/�4�eb������1-&���j�A��o��(����/Y}��P�� ��SimfU�"��ք�G�HD�_�d4B@��n�"�HV�On�RK\f]��|�@���J�ye;A�+�?��E�O�P6�Gb}��c!+92�$ h�g>�u�=>�?�L^ ��	LC���m�l�ȱ0G���lڶ�8�I;����Kw݉\��x�G�)��?i\fQf初�)��7n�LBͣ���a����C�x�x��F2�����]
2���P��X1�V3�������s��m�����ZCrI�
yq_P��~��'�EZ�� �lĽ�-7��f t#y׋.��K���B�{�&������8���9ԯ����Y�!b_�6]R�)�VG�l^�����P�����!�� ��B�� �tuv&�y��cdZq����DSqI�l�6�p�����$�[=�y���忝/�;.j�"J,���"ƣ���;��9�i�����3�h=����Jư�����v'X^����� �3���a�Վ�|�12����T27Dt��7vh���Z�ˑ��Xi�(�psBK���H�$��.�g���g��w�{��ٓ�=��š�_��'M<� E�t���E�ϑ�~����~Z�%�?N[;�|�]x�]��[L?�f�Y��c�]I�������1��B�8�P��p���"��XZ�vչX��(�(6mZ���Ixu����$�/�4�ufU�������x�hA�3E�b-K9g_���N�U4Z�����S���濖�Y
�'�=����oW�!���B^���cAH�m��(;���@-�+�A
Z��ܖ��֮����@H:B@Q˛jG�QX��ӛ[���$�[�4�g�g����#�P�a	:��Ao�Ǯ����}y5 �3�t��٭X|��/S�[�~�S��g>��V�i�T� ��.g�$�I�;ِ�c�X��θ5�M����)���X�����ԭ��1{�f��Y�[��p5.��۪���n��R�������`Crb��$��1l-2��5L�j3�;�{�����Ԉ}�AX��Fy�(,#�@ R*$p�+��3�4� ��9��I@��0�d��dΫ�o��l��I^ЀRn�L#5�ǂv['�ґ?����R%����D����B2���������̄l���W�{n!���N�%.��H�nsu���I����h��7�=Rq{����toN�\���	�*�;����Ń��j�S��nI�ﱝ�h�K^��c0H����%y�ee��kU��es����'�\����u1y4��s"O(g��xD�oO����$�u�Ud���V�W���?%��;���̧�\	#y-$��P���JoI NP�ʑ2ޚ�f���i+��}D�i�6D�O���^KeU�k�?�g�ϫ�8$��%s�l.�Ai��e؄�X�ߎ�} �9Q�d�+?G�*�"�6Ć�P�
:&�n
.��2�/)q�{P�6�-��k�<�!7hn�e�/���:U���?�/��8ơ��Q)�Iȿӯ�i���1�D�W���~��=���pL�����6���[��V�E絉���y,o[�g�uF�O{Us�p�ء��`�,p��R�)���(�T>5�d 
���V����Jaׇ��l�d����^�΁�*b�K��P�"�Н#Gx{��'ΖU£f��c���H~|�cS�uK�������@�QL��gx�.8P��Ew�[L�*&�e>G���/�Qx�=�ُ���d��d������x���<�����?��9��}Z��_jE��!�	�x	.�\J'�Q�d��P�I�	9rfikJ���"�#��e/m�D�X���Õ˂���I�]*���)~b�g/Mz"TA���������Q�!!���?�+X�JR����g�y&�e����ҧ�� tN�'����4J�� ���uሊ�Fc�J��jHCr����ڲD���]y�� Ә�q+iP?�qM�Z��bq��THԦ]���k��� ���}LRQ ��u�c��U5�d�x#7��%(��Qse1�<�nd���tj��2t����i��i��	��1�h�u�j�w��a54CxHH�_���B2����]�~���o6W����j�=U~\f�:�����5}�er���GY�P�� ��>�8��n�"��,mO�p_���d�:�+w-�[���H���r�j���^��+"�v;��i@���B�ɩ�F��W#]�D~U��1��	�Zײnُyr�T-��2���g3߯�fWO��ǷgR�j=��o B fmd�J������*�c���,������#or��q E��Z����e�����d�m��3�԰��1I���-,�C�?[����������]�l�e�96ʏ���$9?��༴��:V�	I@�]ց����D\c�߬f����E%�f��r�����U�5�Ố������S:k�~���HӐ$�e��[aQ�݄�I��A������H��/望p�8]-X�@;����g,�W
�ޥ|]O^#_c�45e�F��yP�f�[�)h��`�y�I��aU���>]j���x2
}��k㱌^��4�xv�d���ĆW�=Pú&mEu�&_H�G���(�r˵�MSuwF+]l-�$z6��~*�(E��'i)O'gQW>q��뉃fD�ֻq)H|�1�,h�ㄛ�t:��s�&�4� �z@w�j�խ���J�Z�������Y��<��Ԁ�u���l�+����v̌7.�������U]י
=�[��t��kKƓ�����gh@Lf���d��v��4��i�WW�!a�����w�����.w4�0��]�@�Ź�,��:��WN)�+T�	����}R��V��<�t὿�\��bvwp Y�6����@�����k���A"�ypO׍g]��۝�z�[,�r0�ƸKN�V��6M8�<8����bX8�!6�H\�W5�Ș ��U&����{g\�_���a��գ=�+��r2$���4� ��FVy@��n��G�F�Q�k���v��j�Ҟގ7�j����7:��ʫ�N ߱��;kˁ�4"8m�y=�0�=g{�&�7�X�]�:���>�?��\��%��uZ���k��O2U�y��L��@2&i�i?�6 ��61�u�����B���~2BS�	��m<,	��C;3�֐�s~�/?N�u��oCn���c��Q��@1	�[�߂�B�P=jȷ2�uĞ�ʤzvAd
]�q6�	�+�%\~#���T�K��]�*���#�,`����NR�!
��2�E�p�E�fiei	.��.wN!�����W]��D;�6�Wyʖ�
�{�V���\"M&Km�A�v�����H��6���l:J#;�'�	2����W5I�[�-���>����?��T������mv�	q�4A�<��P�h�Kv=���ǃVO�C�]yN����I<U"��=���$dF��� fIđ�����U���=�Ȃ���e&�b���/��37��O�~s"|s�"�|�4�D�m�sz��~��Iiș�_Ș�4?��o���Cg�f{�u �f�Kh�`�5َ�P�Ҵv���em"�y��c��)���7��d��W����r�)2�5���<{��R�����R�1:�vL �����7���7�ǂO�Z�v�(�u�G�
j.�����QR's?r,�u�,]@V���_F��
�%E%���pҤ��#����O���)����*9V҅�v��{-�������?�#���*��D`�D�^q��-�l
���Q�L��x{.Ʊ���>��52������g������<�xp�|4-�i����59�[��~y��B�����2�Su�DsM&�K�r��$��wF�CW�����m2��\H�c5����鞒�Y	%��������LW�X�u;/�$�>���Y���A�1	,�(hD*sW��'b�C}�t�/mof��I��o�ã��,%��8o���	����*����a�K���m��â�b~��K�yc��}��2aࠂS㊀�K�5�&{���G,9��D�)�pIM�̛�4Ș!D9szU�zZ�7q؊@��� �'>
��[��Ty+s�ʞ�q6�s��ण��ps؊.k��D�7@���1K?��:�w�󴸅��uN�5� D�(��.��Ҡ�%U�B��,�rz�̠�����> ���=D}��jI*��c�ԫǟJ����!m���冗�f=ƺ�?�	C�{�q�m f��?�⩗�fܼ�j�H�}M��۽�m�CK�8L��H��[,�%�y\��e,�t���3��$g�+,��}��
��⪘�����`z+!<&B�t+��o�AζY?o"+�>֑�o�`Z�c��Y�����v�b�x"��@��K�P_ol"_�f^�0� nE�Pwx�n%U�:G^��Wmr��&\���O��!Ɵ
]��''DS�p�z��Y��a�Ŗ# �+�P��hPxw�1���`�vİc��靽	���䮝�	�� /�޼`w�bP"KR�NSy"On~֕��L��L���7���[�^���C5ĵ-��lV�X�����7����o��~����g-t��b̪�D�6_U���U"]/������*�&h���J�W̑�X3�b�B�-�ع_�y��� �o9�$�QPcm�}T!����3�e�<Q�����7[�,M�׋y�����=p���]�V�nyɋ�f	����Ʊ�Zܾ[���[����h�H�.k���I\x|�2����Lf�&�������?+�Vv�v�ʠP�Q�^S�o^vr��K�л��y��s��}��������d}�۔R�w��P�$�����k��Q��/���tS�	y�~`� 7VJ�GGa����s�Re.�m��I�����k���b��%�|1+ؿa�n��ڒ�#rV����ϽiU|ɬ�+q�1p��1C<`S���ݯ�+�u��&!9=���7�?K��^Ќ��	4*�a0*�*�o���;��U�r������]��� *cl���������H�k�t�f�����(�o�S=�r�m�]ȑ��	����]o��Z#G#���X^C�SeB��p�:?��R|�u�=~%8�Y�fb)�����6�cF^J��Â`��agh�ܵ&��^���8�K���B)�M����-Ͼ:`6u�Ӆ����X���h���b�ZA�W�xL�8_�����V���S�|�/��&�a�Ů��(�R�.��)`\Ԡl�RM�C�JϝP*ZSʰD�Ɗ^�jm�I8�X�O�)����Ѧr�[���Q��&z�\�E
�{X���A�����ه3�^��/�	��%��FM���3�fn�2���9���l/A"����x�3��&B����C���|!Vwr}qnTb�����&Y�" ��zmӿ�9Se!G��Xs,~o���E
����Z�yx��3�S������#��T9 $.�#�l
l�c�vF,\ϭ4Xk��-��?���{�*" *����Uq�49v��wR=�ك�2"��i���
���!��$ېw�횉�>SəgV^фDe�q�"%��ך�a�~��6QQ?�����Hgfb/�	���d�6���@Fe��*N��@�"��a��y���X��DD���lg��"\��Ɂ&���w?��D�o1ڻ�b��i�BG���x+E����Go�;��2�������?ɦ�Z�>����xʻ�"�^L�Y>Q�6�vI�Qd����j���L�)��{���*�!��J}�Z1�ў3M9ѻ>@(�4�����Ɖ�L�V�ڈ������g-�
w�����L\�@R�CW��;��L �!R \
t�u��BCDMh���WT�n/�j"�Ր�7޲K�rBCU$
���`~��G�וyzt���ha�}�R~����p�~4�xv��}FO:۲��F����Eo�4�sԪ�ܽ�{)5�$w��{i�t�Sr��$��w�Zǡ�ȣ�����3<�In����м�� p�@	6��G��u#�2�4E�ܻP%�b�c�ixC/��Y��Bdr��v< �{Yl'!��r�M�7�.�,�Ʊ������2�J�BB<���K���=�Q`���]z�&oGG�h�6��Ƹфƛ��ě	�O�Nd�Ӫ<��=�F;��9�$��S�7� ck�h�o;p�׻����;Y�C%��4 ����/M�x#=RV�֙o-�9�̏?)w<IzH�h��0���1H��}�/d� 3���`m�L�xU��6<�����W1�s��^�C��*�l�HgSo�r��P\�F�l���6�T�]+?ˣW�;Q�a�� g}׭c5J`�m�������U�d(8`���OH����w�Z�`䘹�!��F����4��X>�o�g�aI4(�����Ϋ����9[�����Z�^6MK���/݊&5q�s��
� ������Ձ����u&�9M�;��AU=Ҹa4�Tߕl2mc�9��W�_�*��VXv +,�3F��T:XZ �R���Ϣ�p~ν���d�'Lŷ<!/�!�d��hx�y��S�x�����#��v���SM���(�\l�����	bI=�:��R���v�#�w�-�M�����le��9�~��l� N)���Q��͚:��1��-�uk�U:��L聲�?���B4�L��Q ^���kRX�:�!u��c#��Op?х�$����X�SMC�h�UK��Gn���D�ݟ~J&�1l�2|xڪg��j�����������Ƈn�x�~4 E��,���N�,�؛D:�"������.<Ĩ�M�����5r�G��2b��!QF0�`�\�F"�f&J�`�o�����;~�r�BŘF����k����rE�V�5�P�;�<�A(�b�a�y��-��u��_r��sz�Go.�(UY�,��?�%#�������k��瓴�fr������ȅ��VD�#	2j$ĉg�3�i�u%e'�%B��o���H�񫄁���_V�~���[*RvohG<���ٸ^H�݇8t!���2J5Ք���G�=��O����ëkq�-�-��,!Ng�S�;�S�b�*6b��"�_��ޫ]��C�LP�Oa<i(����j
±g�f�{u#*Bc�ݡ���씢�g�ܐ"�=4��#�$#��9F�� �&;�\�0�!E��it������/�4���Gwߗ�t��S���|:���Oki�O�S����T�(D��;�H��XF��N�m�8�&�������N����}�8ĳe��X�b[+g޼5��ÎMu@������;���0�����ż��%B�_B��e��iW���xϹ~�Ƌ����
����'ZuL6)�P�Ow#]:���.�x�@���M ���'�I�������u�Ɯ�X�(	�w�F�?�}��Z�H�}��y��@8T����>1����# �Q%�x�T��Dx��v̐�B@�꼹��z���9�PP�&��G��Ηr��s[�<��(�hP�s���޿�=w�}.<���������d
8�y2��2Ń���j�kӘ�ƶ:Oye��CL`���1tSW-� �X�A/]���Y=w�EC��Ӕ��aL�@/P�t�m�<BKEv�)�1hf5?�u����R����W�~֔��+�
�Â�n''���V��܉zR9X���r��N���f��M�PK����ۘGQ��W��@MnC��-<�
"rz��]z5�φV���,B��k>�zm��R��e\���%��N�C�@��*DUo\����;��.�G?s����1��>=W��85y�0u1u������ݙF{[�uv�I���v.��W��������_Ij+���p?��9��Tu�˅ǭ>��ş��U�{#�\��mf<Q�OyՀ��A�8���^
48��6d�!ߌ�'��&JQ�;�Rw�?�O'��2p� �>-�9�.�y�#+>�QL����f3�܇K�a]Ꞓ�j�Ay%Jeܻ���Ɇ�q���"�"H�n0���@�/\����܋A��\:�M����!�)��30_,^HB�����)^��v����1A�rk���T���-S�S=���;5��cF�#k��"�CY
:2�,�/5j�Kb�հAg�aa@��S��}�	�{l�<ge�U��˝���C�@���1�dG?��/6���{�������f&�4y,��`�96�r0<�DV�g��q
ORb��]�=`� �*o��̷�-eٓz���^+�����s<0���k�#�A��.PpT�eLe�W����ի�\p��[��yi yU8&�ّ�?9'þ��~�/�k��8��� I�;�U����b��%d.�r,+u�Tݍ�$WT=i�n��	� ���c�w�x�a���©�~�ca�Ck�X/^�^��_�G��_F��I�<�P����ʽb��1"y�b���7�;W�Ԅ�J�:u���(�m�Tn��4�F� U�M	�,����+���+�:��f�	��D{h�
�M:�	�c���e>�b�X�R�Qr�Yj��K�����h���m�A+��&�5��YlcD��ed���~�: �Vf*!]]i�K>[�gF��q����]�3��NJP1o�Ƶ��F�)��IZ��Mj�v���,=$&0{�rů�B+��}���P
Y#�)�̒dEjmI{ٌ��I����â�U���\g1-�$�?�.z*�w ��x w�9�� �C��#5gG
�Md0����>��U���:r�C=�*!Vk�\��q�k�.���wku���:<*����1�v&���Ѯ¹��44uT�.3ہ�>��?��1�$������.�#�0cfҸk��P��9_]��"SSe�v#��k�%!ڛ�nK+�z ��I
�D �gg$��g ��F��5�'92��Y�&G�8X;U�ӤQJ^{kt�����\�n�8�
Tc�ɿ�kVh���GD�o�`�x%	|a�
�̡��0X���Y`�'�-	�T}�五�F���N����,)=ŭ.��C���^���1�q��m����Q��8~{�RjI�ʓ�����F����R�@�tZ�\H���q3��.|Ga�昶��^ȝ�_yIB�����ozr&�<B�:�H�xu5�t��AB����p2K����\Pj��-^f>�Dq�`n�D�;5U|``T��-��D�Lє�1�J*��^��*Oy�%|X^+��X�
�[����66�ȳ|(ą(�`	��j���-E�&g��J9Ƀ���z	���87.�NP���|�
i�;ӌ�a 9:�|.IP��Esd�uԌ�3����5&���wC���d�[��B8w��r��ά^
�N�}nBq�����)����(�)�W]0杌� �	W�g���Wj/�b48'�V6}Q#K���n���!?*֠�ݽ8�h��x>�E�!u���w�UXZ��#;���%f��	~�Iw�&�g�g��{�~lu��D�ymY���x�p�G���S&�.��pWq[�ptӕ�Y�5��Pg�V&e甘b��Ʀ%0x@,f�%�%�ZP۰ia��eamc�:|?�"�K��O:Z�#8���%�^'R s)YI0�@-kJ[F�R�%1�#���t��������oRKIQ�4s0rk)����;\�)J��fi����Bm����W���W�i$B��%��~��F$�V�TL ^L�t�wy�]��ysR�����'=���-��Ț���y��[�u�l%��e�䇖��4�~A�;t�.|[;<)������{e��+ �,!�Y��{k�72���ݨ撮��a(���Ow��O�:��C��<u���7�L#%b�i�O.�&v����9��微GIt4��<����"/E������rR��W$��Ű�R�h�nT|�o�ˡP�\v�*�Mϥ�N2�.4(;H��m؉
����;�/W�����v�gK���$��"��(�,���P8K�0!}�}f��eu'Lf �n'�r��9�y���Ѧ�m��v���X�״�,��M	Ƕy�_魃��$#͠�R�`{�Ҳp.C�a�sp�0<��d~��;s����xr����)P7��a8&�YK����I�n�+n
)�!��9H �b��_=��6�#Q�5"��spM!���V�*<�P7�o�V� "�}l��O���*ߡ��3|�S��6:C~��f���}����n�3��;3sYZ��	C�ek����l9��v�ȟ|�C��[�z�lkz4�C��P��i���[&.�b�-���2.
�R[<ݛ����
�}�L]¨Zɕ�����>����j���o���������ᮐ?vk���nƆo�t�aZ���]�s]�|�X��*����tK�^���f��lO�૘gu�q��������ZF|�*�l$��ɟ5u�&۟Ǩ�iߩ#�D0#}��G@?Hp�V)i�^L3G�[����Q��_f�Ǔ�R��V[F�S��k��Ϳ#�~N�W|�4��y�LҨB�e��<6���rM}�����~7��e��i̽7�0p:6ձa�R�^ �@-q��)�M��E����m�tr����K�����WQ���&��a����a�A�*���by��"YL�M��lg�NV�mEn9�sqE��}����z�����`��s��]0�C	S�V(��B�NC~I��v��S�H��t`KG��:�)����24-���Yg|�[;U�;j/5H��f5�X*u��Il�����ȻL��m��yw"�9h�2�1ΚN��,\�� &�2��,�7��R'-%�W+i�Uu�5Wړ�3�ڪ��t���C��o�I2�_v�1)i6%�y�A������Kf��w�j �`��m]���ճ�~7e�Xv��;X�P�^�H�>6w�:�dg8�^�M��7��a��+���H������R�aBj'��͂�j��M?&&�V`s��jӃ�sb^�Xu�u��ʔ���6>OC�%�K�A,�вR��5z���G����s�c��:1;W�h�^���&�v6X�]���C��:YjE6"�E�17��l�??��O�M�"�e�Y�)���Ο�,EG2/��bI'�Y�?Q�ܺϱ����Ѡ���&�H�D:�ӭ�0/�Σ]ʱh������+�Â>�қ<ܮ���9[�+�W������3���ղ_�����%�ʆ�t��יhٵ��QE13��F�4��4Rw���<k{F�]�ʄ�I�z��{x��	���(?]���'�!�j�lju���[�5�|�F�Ö��)NܫŊo�E�	���hS�7�\�}j笯���D�~h�`��@ �,
z��΂��pS�(�}�TABu��>�9���^����=�C!�.�~�9<�t��͘�:tȢ�e�9����S����!+�/�A�F\O���6���M�ڟ�&�0^�؝l1$}y J��HQ��8�F��*�m{�¯�I�c�C�&�
ˎ����[�c�XmL}`9�;E�
���� �"��;������9!&���	��4�:���$r2�T��ގJ=�C���H��.S&�qP..9��'��������v�}��TN�/H�3��x2!U$�BC����F��v�:���#�+S@�]��ų&���p����L�I�����2n�Z�	��D�:^nU��c���3�_���V~�Y�o[z#4��&�;��R�؃���D�"{�`�����Z�=t�֔����p�{������ݾӄ�/�hPN��xC����}x�5RG��d/��:yֺ�=4L�� 5%���u��7�%��XY�9�_�c���w�X>�YO�����~�y��}�հ���h�p�'nz��BL���
t���{�q���5��߄��7��yd��U�ej���k%���̈́W�Ș��̌���4�<8��R�����JNy�n{��E�r����1�
��q%�ٟ=jmz�E���e�a��%p�ρ�Cd��g][�����7,)?V(".+�x�C��%?�B���_O#����نU?����'	��h���@F;L�\��S��q��4
���pv�IyO#��"+\i����6�5�i��2�aO�+���Y�4�U�u��UR�;�7��aJ� ^�*��5���?��>6� UwCjh#M�\eaB*�1�|ݗu_�E/��6ӻy�Њ3��[CN�u��8L�z����U���t{���F��v4u�X���.n���<��=�?4���u���e�O� ����'s�߳��_t�]���#a��߃b��@"�n�b�7�.��kP]���jE�� ���r���V^gۂ�,�Up-�PD����˥�;�bXf�.4���}��/[�Q҉*��:0����a�xN��$~J6=�V{�9.%�!��\l�"�0ABL�k3Q��Z�TA<��<�`�����h�a1�1��Mq�ų]��@���:��fH=A��hM$�K�ecu��\�q�E\�r)�{�vC)r��w�6�/\7�/ ��5`@�֝B3E>�iv1�J��k��kt���/� ڢe��@>'�&&�q4s;e�	�#:ٰ��;�U���Lkˊ@��ڮ�#Y^1����f� ����M�G�V�\y��Rs�,F��L��)0�B��E��Y���5�����,GH&<]>A����S�x�e�O���i�0��
��a"(���F(�S�8|�"j�ʔQ�/�;*aa@��*e��I^���L(�W���ZP�L��~% OF���9r;�{��[7Z�ʣ����ʟ�t�ˆ�pL��w������Lr�f���1�E��+����w����-t� NPH��X;d@ye�E&��s���b�ǋ\�R����q��),}	R8ـ>;<�$緊��ڎȫO2�"���oWM��)������z�2N�U���Iܞ��|�	��_݀Y��]֮3��e�co��-ңxK�H$�L�Nm��X�r����!49���Z�?�tA��d
�{���:���$�WG���b8i�����@��@rFG:���w%$��Mk\}�^���������
7�� 옘����IUL0�*�`F���/����.�S���ҳ�QW�Z�]�����'���Bq�Q���J*Z�^���&����H�/|,i�I|tC�p�ۯb�F�:*.�gw��࿵�c`{�㗸,�����8����E��'�_��>[�t��-�wv����+�h��?�J����J�I
l�M!3"�@��]L*����F�$�8B�b#� �����H�#�.o�-Igr��ĕ�0�謶�]�"�xK������B NI���Q,�c��_��=�+�M�9�V�T� ݳ����ш��)�r 㭥Dl/_��lͭ<��w5n~��ɖI�2i[+��߿��7d���U��рMy��M�bU�w�p��د�P��`�覇�lhxe9��_W����ܦ���L�ݡp���:p}�1���B��>p�D�ʍ�W ^� ���H7Ǧ+:���'���H;�x��7�W"��l�U�NC 'лL�:�Y��!��L��h�(��Bi���?���2�j�uh�,��:ve5b��ǉ�6���'���K)R�l��EȸR�+�2j�P�bJ]D ���1R�˘�8a�o��LD70?�s��IA�D3e1�k�<:��I����{�5X��ć3�p��� "����4^�*��?�"��X���Nݧ���>F��>�x�5��ӚƸ��� #ޛ��S�ϟ��]��W"��
�7"�j�ݻ�>�	��ϣЬ��ˏ�M���)ۼ��nz\|���nY��	�%g/`"DQ�:��J;7��c�LR��< �.>�W�
��4�2i��ux�R.�� 	�>��"��n��;��jt\F������Y��K��c�!��p�����`��^zCQ@�jCzR�≮����΄�npT��ϡ�jj������ę�"��m��i����7���_'�ۮ���mU�aT�_D9߁4�l��	�~�:�*%mګ���@l��m�Y��^UP�&�A�Y$K���g�~���υc���Κ��ɀ����0o�6ZU�.ܸ��[���������ꇴ:�M4�^��p����~:�q�?�ě+�Zb�*��2/��i����A+7р��[$J6>,�6/@${s`�Y�,�ݣK��p��+�g�҉9yH�C�̫\��:S����V�o������}'�]������x����u�$+~罅��@+��q|C� ���md�B����%�c�f�g���s�ϲ�
�GV[|�PN:�+�\VsJW�����*9uDg�$���ڡ�� L�_�+7vf���ʻ��>گ~��<Ɩ���D=��8��՘B���Jm.�M/H�����	j�@��`�r�wr��h���~�X�&���pt�H��?�,���a,�X
��(��݈�A�q���/�l��֪�a� 1�
��b����ke���lF18�h1�0�#�05�N�b��84xf�h��z���F�嵄?�/"�2k~r�O���3����--�z������պ��\zJt��[�d�Z���T/	�H��f\�C�����x���-��Yi
*�4>��[�, �g�FQLu�uL{�C!O�ɂD;����@w� t�!N7�!`m�Ҋo#}	u�	_�q���{=������w8��+vM]I��o&���ZA7+�C��c?�@o�����gV� Ƿ�$)Z%%e3�=:�ܸCd~����aqPB�/L���PY<�w��ky��}���n�����F|6��p���G�;����L���<���2��{�R���j4���rS35R�A�y�=�r�## �w}�ǀ�g-ƃ2*�a��mǥ��J4���pfv������b^p`�5�V�3�]_�}��jR���4W�0dY�;��=	M��π��b�㷿��� 84_�K��b�@��9����MMЏ5!!���e��D�#�%4��^e$t㍷Jcԇp�b`�ED�3���I����7v� 0F"�D'�G�Jɞ;�=B��<1w��E��(�U�ޤ�f��
#�<2f����ȍ���3��@�Kɉ���<��ť@,)(���.��%]y��j���[.��ʘE_̏����Rk�A�h���M�	}k�V�L!X�Ņ�"��}:Z��j=��9���I�a3���y�����o$������^��_lU��O�_�݀@\�b��q@a�x�e�H��k��O��\xAd��t�=�%b5ĕ5>
�ZF=d���Ӛk�H�x�����뚓F�����+�c��rE��	�<l��oT,�rN�j�T +��pF��#�v�U
��u�������j�;���H�]Hc��A�J�� �$�M+���M�[�����'�;���/T�$��5�2Gu��m$��ߒ�	 ʣN����R8���k	�F
���M��c~��ӥ�+:x�+�3ʹGt���z�=H��r{�'��5�8���Qe�uUY[Ea��;-,�Q7��߁*�S՗!�6ԡ4&��砀D;E`�����j�K��Ce��S��D�Pf�:�Q��J��K�\{ml#����J[>��1��'�O��󁇔X`�b$���Xq�#��A��M9B��o�b����2��L�_�c��M:$�7�5l׻t�1�y�Oo�4:�o�$�~=��)QE(��$�r�阄��������GrEeP�����o�j0����`�V�q���B��Z��j6��>[��o��U�����]EY0�G���Gɒ;�9w�>+NZ��{.I��	�<�j�p�T��2���m��`d��:+�6�r;-4z��9���h�������/>�s(9�=��_�����"�4,*��� dR+r�4��jEؖ�7m��ͳa~@�}�)s�`�:޷�8B���u+�@��ߵd¹h2r�E�|�v�j^\�Z��8a0�]��e��9R��M�'ǜ�hk��h9�y�}u��P�W�-��{v����A�Ct�52ꃫCznؑ�����Ohʨ�䰇���h�0�n�����3�P;50�53T��&��ww�ET[�����S�O��c^ʂ.��!���|52�T:&Uc�y]SnH� �jK����Ծ2 ޘW}�������a�'�:����=��͗�6`ap�s�9�!a_��z�B��G{�"y1:n_on����n�Z�s��OS}]"O����_1 I�(��C�tM���k����2�IF��|}�8T��kl�{�������>~��'��SW�^RSH�&�$������e.{Y��S����|����ȭ`�XB�Z�����k�������9z&�{��\0D����0P�
�q�Qf��V������y��Y|mdY$oL�ͫ@A"�Dԣ���' �sL�Լ���oRH�����2��~��8���T�3��x�.���䣯NN\�bP�B���#�AU�Gb��<����gi�냊�\@Z(s�FW��(�$}?~��/'��e�׽;����l�$��!����������p4X�qw��ul��_EA���MK���ᑬk��[�6��
nA>��d������R��>;آ,���i��f7N�U6��s0��7ӥ|�to�����}6�zm ���*�6.WuF�tM��lK>��(߯����vْ�jX��ڮ}�� t�r�`h�X�-&|�W$~/��y����e�M�;;�������^e ��_~}������ ^�Q`�K����*%�yJ ]8u��ڒR��U��6x݊�Q�ff�7Dz�M��v�&������ߑ��B0�a�NY1SM`Z��6Cp��E#�����f[��c W��S�:Ҡ=��"F�@�8����n*�g���|�����\�o���[��`z�H������P�����0te'���Ɂ*f�i;�'Q8?���f�'��6����(�+�Y���okZ�`�n�zS)A�$�<����n���Te\�Є-�ʃ������=^r2m��v9Ha}���U��E�~c�Ax�Pe�u6P��������y���l]�5YM:6Cb�A~vJ��p�J�k��Wh�����W�f���W�Sw�v�7�;[Z>IvKe��Jw�M��	{����m���_�'aR���O������}���n���G(0F����|�G�+Ze��l�;��
L�	-f�gh��'C�gё	��up!�h7���ហ�V��'}�b�����C�>�I ��6*��Z��LrA������F0��C+��cJ{���C�FU��>��R��_�O���cM5�ա�I�D���?{��g(����G��M������0�� ބ�%?����^\a�i���N_��Yu�j�K��mIV4�k4vǓN����}Af�>�t9�������.�qz�F�ݨ�4�iLR��K�Ҳ�^��SoWPR+����a��S�unRp�08$�6����D~xhy�c19��E�8��)�C~��+l�kۻr��?ڟ&.~T����yM*m�5�Ô��i���^H~�a��gwћV@�c��ۛ��X�l�u(a���vC�0y<Li�3{فW�
z,�	��ԐU���Ә&H:��IW�Y\�9�1`s�Ƿ��ޢ,�8�W�uxN�}�I�p����S�2f�4�P�
*�Qv��$��~�v�U��W�b�/̠�8���NY�a�`d�"x����o�,1�����B.t��jm�+78b�X�"]�P��P�Oh�f� [\f0�*��t���-R�06��g��@��]�1n�y1zg]@�,k�w�'���P�MW~�wp����A�!,��&3����m�d�q)��d���h�ҭl�ԉaԟ��$!cLfZN7�F{��8Ҋ�������f��]�-S��N�+R&2T4�R�8ǌr�=]�W7��@ưni��xџ��&o*�B�'�c�'*?L���N�H�$���t�ꐏ��b�=�@[s�e���SE�o�� �M��ԃ�����	φm2~lw*x��c�����'w�V�?Ho����g�Cy(@,Q���s�rx\��`�U�A(����jw�N�'�r;巄�Nj��e.Tl�F�&�(��G<�����~�"Sa�'�]b��j����}q86��q�D����e}l�a������lt������(1�wt���Ȫ����_�
/�o%O� BR �f�1C����"jS����e&��e�֭8�Ȣ����f�FSoP�XI#db��>{�V�A�j�qϮz�ID��z.��ĖW&�́a��V��D�d�09�8\��y©̂4��y�v�Q<@dm�����W����93����a�;�j���|�y&��߇�ʁ!��]}�F$Ye�uH�w{$�O����}��z�n�F��Y�u<�Rz�%���p�f�ajA�#y���0V���Hfw����DPTrꟍ��	���_��ܯW[�ƥ�H9$�N��n	gy�9�Cj�m-8|���[;j4�_�8��iX��o ���Ko���4�1�4 ���]M��j.�fd	�<�-'kTƔ	�9�Lu��M����7���r�<�:�*F<c���	P%���{�5Z?I����?1�7Q)��GC�/�;�[���i��O�N������]��������P������{h����b��`��2��3��ѯ���^E��ӔgE�h2���	V�����	�A���k��8}G\�hQ�00��&�_\p/����hs:D0^�o`0$*ӥ�q�z��!�V���_�]ø�z��ضk�o�QbI[�1r.&Ҵ�����hQB��e��٭�b	Vdtj?��F���<��6�֟���Zǎ���.�֞v�5��0b�4�@���Arڠq�����/��82̏p�'ޅ"��8s�,�"���B̉%E�Nd}���z�@�b�xT�r�U�E�iA�b!7�$Ug��O����1��0K,2em5�,�1xsN�ۯ�|��X�`���W*��={�(�D�i(���2ۼ�#Y�Ŭ�Tw�_������3v�+5ی�_U&�\������]"@)�I��-<)5$rf�C���ɕ���D� �eOCC2l��j�
M/�M�:  w��<�U�H;�\?��ͣ|;~����Z���%ks��J�7�zj�H�����1s�������x�D�����g0m-{m;+���D��s{�6�@��`�ȡ��c�\5L��<�#A��&���Ϋ�;qkj��]�~'֯8�����O�S7F��9��5��p�q)f�C9#�Tŉ����Ќ2�H�"i�92����R�LQn/�uS5I�:h���ԠC4�؊�hC#(����崙�����$�I2u��1y���ǧ7�[���R�	n!<,�hi��:o�k7�`8M�ҿ;�,��>��~��!���4�Ǥ4D_��jL庲j���]+V�t�QY���#���n,�Ⲹ
�5�P��a�qG� `l��&�rS�-� �u�D4����z��Kǜ��%��8�������.*��6��#��@���`h��=G�����'>��m~��H��7%1�H �d�/���=KAV��̷�'��NܯL�M9�W`f�f�uC��[d���^��NpL80>�%忖C�'.�����<!g�_���mM��åw}*�p+�M������x kz��k�ؚ�Z��Ⱦ���4�q�\�7>�:���U�-G}C�@A�p�(�:���Ks"�%ƻ%�����ҭ�p$�[�~�~\E��0L�>'�s����8�����]�x�9��������JU�0Ob��hGA�J=�i���Vh��H�ƏD9u%�/tr���9�\7�s�284�_����nn�:�z��S\oJ���x��@���B'�E#�k��e#~T�R��t��?�9�%�F�(��Pܔ�J6g+,��Y=��
W1����(;���菽�v�A��r&$�׌f|�d?.7Y�|��@��K��Rv�Z+�����G�1n�B}�.��{����5x"�N|/��?o ��Ӹd�\��ٳ����g<PE��Pm��!4�`WL[�R�E\�L<jVQE�fںs���i�X�ށ>��,��A�]{����������dR��G�����8��Z<�"��~���/�,�d�c.�n��W�)?��D��4���c��}&&A��1�L[[�urZs�P���B�d�gx�c�w�%ư��qM8�l����2-��5�]1���9V��H���D^̚ԕ��.y������������=3����qf� 9z`��[��`��xE�6M�[y{�S��f�*&����9�Te�w�yǃ��_�	��9�ѩN���{%ǕX0�l�,�wN���G�,�3�!6~��U~*{7A\fs����K!Ņ�=��-�IS��LPo.�R?���C`
Ȁ!;Vh�gw��"��E[f�5���n�l6�C���e2Y���JIJds���F�4��uڄ����$�i8Hc��c8z��0�y{�_g��mA�?T+ �d�5�i}d <$Gi�v�tj\;�T~$xܦ�甓?��@������a1p�~��6��IGv�ݔ��7��EZ9�{��:o]o=�e�o&
��:x���,��"�{�])�������b	�ẛ[F�`H�v9X��=>ɓ�=^�10�w��U<~��X�?�sC��	.odRd��������f}:/A'1L���P�����DxO�����%���SӤ����SJtC�ֶV�MSp���b�v`�X��D�Ӗ^�S���DȞ������q��_����^�� Rk|�G�r�#(��6��v�~c��;�b�d������(�^p��� HLB�A��(>_�H ����
��g@�vZ=6�d/{�����]��8�F�V=܎�%��
�J#��c�ɂ�}�?�C:_E�
g��y�uBM��m53:i�:��27��+Zz�?;3œ��N����=h�oHë�ل�x$u+c>f�#"4�P���iFz9���N����9M�:y��)�����]PSe���,�D�@羙�.9���t��,*ŵ&H��G�pjjof���ʀ���vgM����A��A*<��S���r���
iǭ�>�,���)�.
� ��9��P&�Bgk�.�!iZ:똇-S�f��8��dѶ���@k�7�"0Mm�~��~*=D���M����l�R���bR ���k�/7��+��JZi)�<�r֑K�͕^�jK��:�~��7�����5�&��Hk*�K(O|��١&�b������˧,Qٟ���i2�K+$h��,�de�X�n3z-���p�j�x��/����6Ʒ��(2��� �=��!I�m�@òу\;5,A�ކ�)��[$t�S����&B<XG�( Ϋ��4��va��/K���8<!�N���æ��0��$|$�p�e!�Ň�u{�4��#��)�%囲�p��v�ˀ�g^�V���G��E��ٲq�ς����W<�ϛ5�R���7�v�6��h�X3(Aw|cV���ks9���H�c(�Ey�\u��Hg����7\�Va��N��K@��8����i�~�n|�c-��D��������$~�dީ�A^%���j�8z�kJ��x�Ц"
�HF*���G���5܊�=��['�X��9f*��@��I����鴯<�z<ߌ~���x탨Ր�:�ƙ�����r�pIat����	@����p����4t������� j��9�E=�\���CU���Fc�sȮ��Ǣ����&B]@֝�iTZ�;b��f��s�Ŧ�ۃ0;����<��s�_\��@�V�{?��k }1�5Pd���"�|x�v\XG�����)ב	/����L���:R"�9��V�/�4����;7�,Vn��ë�����/,�K���;�&��iWs�Mq������$��`�X��$r)��J�?~��>��2�9�e�Eh<A����O��Z\�N-��'1��������<��3�������~�/��q�'9��}00W'�����ݔ�-��1mϥO��n׼��R��$;��s�V�1�]�]D�Xv	�������1�Ƽx?8)#HIQ#������*sH��~@�'�E��~�u���\1���i�9M�\�|����V�wpѷ<��t�7��2i�I�?�,��zg��aKQ\=��!�t^�Gꊊ+�'{��� wWR��q�x[ς�--��^��J�'Y��_���0s�5`�$K����S9
'�G��˓����	w��w}�2�8ڿ�{��i�<ۣ�L��dّDOS��aw_������! ��IO͔��^%�8ا������~��ʔ��|��6�'+�M?Ʌf|�?�A��Q�j�� ˤ�v�P��e �vqԉr�`�)��0R�"{d�3��4�+��Ի9�
k�+�F�]��@��a������o)�&G�cK"���J��מ6����WQ���ֻ_GTO̯������mO8[]6I\�r���(��� ���=�y�K2�v $�������,�GP3�����v��]��)����t�|޽�]���j�;���{��%"0�~��8�!:�B>"�[�Y�s�R���v�/� ���0�^�h�C�������(8b�*c��^�n�Y����C���*E֚���cX�@*Z�NډK@yz���V2x�
�Z�g%W�$��%��������%Ϫ����r��Ӽ<�
�@P������z�52�}����Q�!��1.U5ލKp�[׌�.j�@k���՚�CC��"�@�0I�e�����I!$^\>y��r�����#�]��D#0V>�ؔE����3H�ly.b�^RHmm�⓵���bA�I"�.�-�$��7��$0t2Z����	�M?�3��F��F�Vݗ:-�Ĩݰ9��Q���������ĬڼM8'��78,��jF��o��Rj�w�E��Lyq�3�1�FHU��RF�̴�$�^m�_x��q�͝���X7#ƕ�hL�_|�>�8v�z����|���� �b�/���gPa�D�PB�'������ω�(���P�O�����qA.CTNj%�Pi����)�'x��O�L��-z!��
<ޚ:��y`�@f�J)v�i�&-Ӗe.�*�/���WH��:���O�_(��eK̴��n��\I�:��
߇�rܴ&�mҐ�M��g��X���Up7����Q6��U?��p3��Lw��*���󄘈ck7�Q�Y��%� �F��B�?��u�t���t�t�F�&�>�0���;|x����e/sЏ���!Y��e�kIKZ�m�|E��"
�JS:��ZO�D���V�db�ҬQ]ց��f�Tfr'��yC7�$��qp;t�Q�"�}X$5�b�6��<����#2�]�es�1�j������zC��N�)PQ
kP�h`�cJ+vP�dBO�ռH�P��'�V��޹��c=�~I��!**{�s��T��O��a��PV�1[��W	W��d�o�@��+���'v��Cr��V ���Ҭ9$�˜sϋ�
��U�l9���D���m�.Ժnɫk˅��80%��Sw$j*�'B;]�lײ�z4�V�'���ī�;����3��
��f-Ҡ�� �դJ����H�d�F���X�Ѹ���W5.��l���MP�L�=.$X��T;0��mgb#�\�U�(`�#x��T�����4g\&V��ZvtJ����v��Lڌ�t��C�R
��ю�0�@E�g��YD��̐h�B��=��4U4֎������@�j�9b=�W�E�%O~� ��k��L��*�5O�퟽��07��7�{���Ο�#�]�2�6�~˚+aؗm"&�	曷rM� ��]�j���^��i��)k�O�D��}+�ԗrbry�fQ�V�
�o��0�L�ɐXF�=8&)����sH��ވg��=;���>-};������@	A~�iX�Wg���>`p�*�������U����M��;��u��Q�d/Z�,��K�Ir�n;8C��0�A������k}��鴛��;�la�=�A�
$�WW���~�k��g!a`Z�P�i��b#Ѣ?$�X�=��k><������>ċE�	�.���4�.x%�t�<�<r�'�m:%��!��C��qy�R��zΞ�:�-nok�Y�TI�2�6%�����h�Z'��HW6�����~��L�Y����4��B瑐M_����,'����38��'amo����B�Y7�c�p�
}��B���v�����267���f
V�h�p4�YZ�Pgݻ�٫D�~r��1�%%�#J���ݨ�u+P��4k����<՟��Y�c�M�˅`�+q��ו%C�4���O�F��w��?&
	��S�QX�}�?��J�xr��0%�q+6C��Q^�#�~"[�[�Rb��ސQ��P}k��zp���+�B��r�0wB&��9�O�� �RVk�J�əv���4��)R[s�O��Ɗ,mP8�Cds�-��엮����OC��oU��wB����:�)�%�a�� @�z.�-�@8�HX�bj�O�K�a��kձ��nu�|�o=1/y�7���Y��bŴ�G4�X�����ّ87�K;w���O��$d� ��lUBmY}��8�nLAC]����Hx��&�I�}}����j��j�3_Cx��]ǌ0\��j���gbH�1f	�Y,���(u�[��p���D>8=4}���j��;2�y�4:� e���1C!N�@xD���-�k!�X�8ƛ#�h��ϥ� �8cC5ƨ�p�s����$��f�Q�",0~}�{�2�k(cAJU-�f�u�u�:sU��� ���w���G��/C4ޥ��^��u4�v������o=aW�5�����9s�R��p�����,m)���>�}7��ݎ�@n�L�^���){ga9��S"϶8��%�Y�r���h]����Bf��l�O���b��f�3�+�}��Y�����f'>5�����NP�B�~G�MB�Խ��95[���1�N�1����hi�J�`�FS0k�0�;%ʇ�>���
�O(�lK��B�T%&Qu���[x�Q1j@9�F�w����?[���1A6�{�u�����U-ͬ�a#����E�)������ߩ1��+6^]f���7%� =��u3�QC���4��uDG�Z�YÌ��çu}�L8��}���	*�@�,h4ťx����}�b�����'��Hن��ix�<-!K����-Eś>�ֿ�wT����q݂)<�����$}@�,�x�5`j1�����2#>2D�7Qsw��_��P�T�CJ�]���~=q������1��Dfg8��X��F@���+��qB��n ���E�&06����,g2����[7Y���D�������*�HVP:�/�r�v[�*E�Mm��۾$�/<�Σ��1�b�34���&���x�� ��j���돍��w;�uR\s���X޻;TK_`�0��n����㎵aT�c���1!Ē=Q}���Ԣ�|�����B�.�����f��W��Y�T�DD;����CZ�L�U�;G�wI��s��ʐs[7,
���U���\^s�N �%�hF��_w&`pp�&q|�����]r�] v�ނ�RJ��:Y�d
�.G�ܮ���Ӏ��D,�l��l��}�:,�w:ZHSEa�g�y�������hO�ڇoƲ�F)�xY�"n|����7Z���n����X��0z�#`U�}7Zn\ֹ��'�WC%޼ ��t&yHn�0R�m=�˵�O��Ή�#|��M�9S��@��� )Γς1y3�zv҉)SkEeé��2>�y �����vIj����$	�V��3�EԒ�1�"�z����w��H����/�����U0��Nyx������(҆�8G6�_�FuA_�q ��=<���{��*��L��|���`
q �%ce�)\��x�׽V�RW�0��hOf��t=����UTmY*9�t0�C��
��<�?�F9�e0m��[��{j|�/��tB��q����Gd$��
X���好(�n�X#_�~���ܛb�qT�.~VNL��A ��Pea����e!q7/n�������p`���($Q/w�MC*�W<��@����s�sg}��/)���&*�iqb�԰�:�A�cG�p,���V�W��q����p��t	*�l�yL�ptC�:(j�0�2~ �{GH^���}wŀ
�U�?�_�"}ޕވ�[`�����RK3����Q�غ<����<H�$�ْ�Ŏ4�Z�m#Ō�U7Q�E݆1���7(���AV��P� K���İ-?�8�}�*�T�����Td�bĶL=2����z�w�a?I-z+�v��0֧;�c=�zҏր]BXy�WgS�r�7��G�h&��!���t�Rpށ��p �����c�^���cf3����1e|cN�1�P�g*
'/�,��T�:��0��ϝ��jh���o(�~�oϢ0@N��UL���C��E# ��a�&�b�,�n}�e;�>�9d�
 �)�"�jfa j�m�2�$�R�G�2Nx �	x���+zod���-ML��*�'{=����-$�����Ұ�#*XiO�O{7�CS��nG=8�V˯�U��;��a�P�R�����t��M��=��-��2�tV:P�3�g)�����0�$`o�L �t*>`x�0+���,���F��ٝ����)���~<���C��������B�҉�5o���w]��n0�UWSYM�O��EL�d�/E���Js����+���4�b:T�MUȋEK�m8W!>>��q"g����O��
�|V����>�*'j�Y�R2�)Ԗ�=M���ms�c��Nz��_Q������1�D������p�����wC7KA�Y�u�4�2���.k�M&f�5X���ƅ�:3��
�w>��5�ĴK���\�j��Ȅ�2 p�:����kTQ�Ŵ%� E|Xt���[b@�D0ٯ���$yM ���BtpO��[� �g*$s�-��K=y�Z�ߒ�X�
�6����
"���۷v�ѕ�7��.
Qa�a�K�< �G���/��dC�
�־���h���]0�Ƴ�#��M�
(�	�܏I\K��U���e��Y�L��l�����j�毱��/Xf�CK�:4���h*���Y�b�Ѷ
'�U�3���}��	����VM�����y�1u(	d�7�'y������H�|�4t_�
Y	4����u"�	&��C2p�Cr������o*;��_�n�<����[~|�i��1&�:3V��H{C��P]�����{�mtA-�sܖ��i�Rr˸Q�WxI;w�'��ߐ,�eg����x��	q��	x��k���Jtq-��2�>؎ ����\\{�}>-p�n��le�)�=����g�uʝ��}w�UH9�m-by���b"QAx��P�!8z/eO�vW��0��-&������aq!�.����Xq��apjx�YX�*�a����$���w�j���o�I\�@��g����۱�_^msk��D�!v��P��;V�5�fM����4Fc��^]��햅�;��w���=��n�`��8�p%g�+��5&s�J�z\[\k��f�:��*f�K+�Z G�[�\����8"hT;��F�#�\em���ޤ@:Sg~�Ɣ�#hKG�;o{N�|��|f�x?�b�[����yq�s@�o>�a�HO����]����<��� %M�>���p�n@(�2}�p_pb��ַ�=��gG�C|@�I%�]QA��ael�H=�?H�U��xM��+�2+`\YWoԨ��1�#�VWӦ6��^5Y�.T$�����x,Jkƴ��},����"�LGZΊ_~�
"��q]Dv�5�eN�Σ�G���^=FM��)	C�a_���gw���r؂�-�τ���#	����X�(�SN9ŴC�Pų�p�"/��=�eO*P�0⿄:��P�Qֶ@����y�4܆���t@��('����[�,9�q�P�c ���J�G������mum&2�5R��Ag,��&ӍE�F�&��1kQ��F�:V�r,�'�8�$�G�L��G؝<�bwATb�P��N֮9�M	�wN�<�����dA;��g��8�.
��#�jT%'rv����&}�w6�^gy�n�h�o��=�,�"��P�(.��	��]�9N	ƔRr#W&
��	�ɍ�
�5��#_�J�h-��/���B�~*U �W��B�+��Jcz]�l��^?`ξ��ϓ����˺1PŔ]j�ٹ$�,�|�Oٹ��0��Uz�oz ��˂;�� ۪��Yk�	pz H��ý���L�~�N���:��D!_�Ӆ�@+H��!P�Te�M�I2�4��q`@�8���P=>��	Ȗt�j̕����RrHG@_ռ�9	-_'��x/w}�td��@�����(d���|ͽ�HJ/�n{������Һݰ�B%�J	����X�.���feI�b?�s�13HWqT�{C��iA�����7%3l(�`l}EF4<,��iC�qbCH3{�9G�WW�/��ӕǈ|@Rn�4ϋ�=*5�TD��!�t��o�G�nϔǛ)�����$����y�-��FCe�Òd;B8^T��Ipv��F��9��&�Z&[y�K��>X4�TIY�򠐒K@!`���K�a��U��.�l3ܜ�Y����prD��K��~�Y�#�k=������K˷Ņ�|H������t���t��p��t~�9���{��%��rl=�m4N�-�w��G�:���L�y�Ѧ����������oP,����=���^J�&�<c�VW��Q,A�vߕ���זBIr��?�N������Y�7,�� _`ܳ����2��Y�0M�9�46N�<�Բyx羂����AE��Eg~\�!KF�>�r�"RE�ه����~�z����t3]��Z�tF��pM�Z$o�Ż�����1�$��F��4D $��f���>�Z����D��+�>=_E�D���砤P�����ٞ�<�)ɸ���M�_q�0��-}��T�(������[�\aH8����]�:��GH���T�?�n*�U�� D�t�M��j4#�u'$�~��r���'Y�<��q�J�h1JK�)+��)ո�b�/��׼�@���.�
���7��	Q.s�Y�P�1k<������֞m�m�Kn����ء/���|�Tl�
)^�O�o6@+��]i�O)x��m"\L���8�>�8~�)�H0~���5�"��*>t@nq#T��\�u��Z�V�]����I��f~�u��E���3��(��ˑ���t��c2]w�x�|v���; ��댨�$	moy�m��X݂u��\��^M�K!%}r��P�L�ݙ�A�Q��r����*�5x��8$֨Dg��y�T�1�UqK��n��V[<���q���lx���x�u�i�1�o��h�\���E��E����ħ>����imҧO��n�Rĕ�	��^��>T���@���$*3��a��5td�`;��n��M�5l�\I��ͮ�R�%rSA���16�	���|�<dǕm�z�F�V.�F
�	>T��(Thp�d.��G�B����Bb�3tQE�}Mp�j��7�ؾ���]��h�:�R)�φ�63�Rr��bK)XaE�6D�.k��D�G�KT���*��Ӏ�5�$�C/�*���O"7(�[l����+�5S^��;����+����5x�#�~O���>j�qO���|Q� �>�y�'w���������ǹJշ�/_�E@�vu�s�6�]̵��l &�7�æ��*����e�;x�?�3�qԭn:p$(?��K"�5X?������DVg�����Qф)��u�`�!�؉��>���hL
�4��S�#X8f���4i���lw�q�����'�&�$��X�6_-��;]KM*��0�M�����������T�"sL[_��Y��,*�8��(ʫ&�Vn�|��*�an=/��`�VS9�ee���u/��fU6�:\f"\���g����4���J����e�3{	J&̆7h�A���gsY|N,�����O_!#���$'ٰ:�˟��DO�^�����n '���{W5m�ܯvv7�$`�a�(9�g	g!u����V%F	ˉ&n�ٟ���	��,ɽ�G�[�l��Қ��A��/]����E�I��˄�Aa%�3��$�lȬa�y5_���-�|����Nz��@��[���������$�*����-,M�����e�Q:��5����{-��S1�a`5L�bW��{�	s]���[�A�8z��\D��"J��r��M�G=�8��(]hwF}��1�� �P��z�yz<
�a68t���垤,��9~�v��e[5w����'g�{���(5yɤ�9��~���k}�n�aw7!S��(�C[��ް�%Βx>��R�"bb�b� X$��� �h(�ˮ�HD��+K�Ԏ��A��2�S��%A#�+��lFs(	���Xb�*IQI�!.Җ1eUdh�;
4]����
|D�@�����Ok��4��b��,��.�$ ޯ��}����@���Ą4J���ا4�6�5���t ����c$����>k���ua��ޘ�D��	Qw�n�'p��X-b��H���2I�=��y��x ���j�ȅ��/!�l^�<;�������2F��f+^���*0tq��M,� /��:�:Dj���E�"��-^o �kGz���:v+ �Ɣ7�X5��n߾��.��vU���FkK dey<�r<��$%��:��0�m����G:ό�^@]iw� �4i-@�c}fB����ł���=�טu�_�ɽ� ��#�uc
Ɠh&�%���6�/��U4*P�e��P��>��s�g���Y�E��*nf"��
�=��UQT^���hQ6�f�G	��F@�������"b�Q� ��P�CI�������&%����N��Q`-��J8� �/�Rz�>O�Jr�n����I)g��`���z��k2�F�P�hA,'
�?��+�S� ��>�%��`\�C�0�-7�%8�B����g�|U�S>m�AZ�if�ɫ�,U��P>���ʶml2�!m���h�_������'�
��x��h�jl���y��n�ap�~BH����F�����/������_@u"Wd������z�b�6=���x�$ߙP
�����Rd}ȣ�8�J\�Lg����W��F�%�H0m0��6�b�L�-���Z_�A��J�Mj�y�r�z���~���9(�d+%�]7���2�ܫ���+66|i��w}�清��f-�[��{e~TiK���t4Pn`����s�9y���f���
��r�v�\�d�΅����dZl��]��o���0 es~ R�� hQ��_����v~9��DT!�r��!�"�,�Jy�\I�iT�r�=Y�jdzw��v A.�\���?J�Z�F`�s�/˂��j�/ր?��ѡ�9����F~��z5GZ�bQ�T. /�w~G�	�1F�z��_J�Aq���Ddb΄z]J����#�'��ԡ��j������������ �9�YT；Wd�
|ix��MK(�)Ԣ��I,�R~�!���/�X eZ�.-{�]�q�_��� �J�bp:�/��Y��ic*�B��R�ۀ�}���;R��O�����ˤ��k-u�Q�ۨ<G?�?�w@C2���}�s�Lh����F0��95,<�gn����'f���#��m�6K������tơ$X�XS>�}n7�Ys��IR��	WΗ�f����L�G� '�+Qc���ivQ��������}>)@���b�L�o��L@�����Y��.��%�cȴwg�f����A��u�O�����J�s�
=L:	��<���\Q�|��")=�E���8�-����I''��t��;��S%D����ݏq���l,D��՗Ot�UOy��f�3�L���ӐuyP�.�ZT�}�M�b���8�~�MبQ��d��	��-C~��T3�^w����\��g��G��U�9�g:�xm�Hm@�c]��uq>�//�J�{�qE�[t	60�ĩ���n�EN�����;�*4��zi��+d}����R���Կz#|�$1��/k6���^5��._r,{��O�W�訑��IL͠T��S�H�Nn[�y�e��d(��N��/���y��I1�h�'���o���Yzo}iʳ#���Re�g_e�1��ʉ"N|�X�'l#���,�Ȍ�Y��_/e��$J�a��xCVz�m�$��#����={-�3 ow�q�ϯ�$�����6/�`#�1��1��a�Iv7M��0�4�.f�O����{a��c��.�^� �k5���%�I#2��b�uPÉD�2�G �7�Ǜ�'!�Wf�Fl�R�!~V���|��X5ѷ�)��=m�$j(��)�qqI��D#t���������֢X�?ܘx���S�LN֚�����01��b�Y�Fwn�� bMSꜦ���b�k�� ��P*�iX��*�c�d���
�3���I�5�P���פ/��exT[�1}�FwF,���u��\A�zI��;���]#��>wə{�_��!�7��X�<�e���FӺ��]J&�.ǃ�#ǿ�k�)�Z/���}���5��Y6��v�T�'�JӅ� �X�X�z�/��M��d��~�8&�E{ЧK�w�y5$���� 6���4!�$[;|$��J,z+qHs�=��W���p��1K��<t�_�4-F+��-hCo�GA���LQꔕ��=g�v�FȔ��s��A؍�wf0���O,b��n(��ָVF��9�k)�ҷu9��%f�:�����m�x�^��}�&�@��c8diS�d����.	ج�fe� ��3u��tw�N,�A�..�^�:ͭ�� )�1$L>�Ũ��i���Jf%u5w�a�d����ѤXl��lV�wz��<D�S�vb��9J��,��C,/�d����e�)�Z�\=*���ͤ�̿W��Mؿ���-ak��,6�֊�d��тD���JsI�RW�7������5@
�&�,�)��BR��~��0{�;AqX�x�S^6�F百�KǸSZ|h��~�g��
�~�<PZ�؀F�� WR@�rF�IiL�[�W? P*d�t�n�z[�r|�~�RR������-w��Y���k������k�Ȧ`H��A"w�����d�H�De��O�8qk@�	-Nf�7!�bd7<�Gu!;�{W;p�El�=���w���`�_C��[#p�΢@��Nu�Ww*1��8�U͎޳��]|�������-ÜҒ���c G�vb} !��H�@������A�0�x(�6�;��ݺ���X�y ���r��%ϩ�؋�\Z�Pj6R���7����(^0\c�4��{Q����öl,	FD�=L}�[�	���:�ԧ�o�̷���:��ޟL�&nu��~Fu���������M�&d���Y}�;�r}�0sȀ��|f��11��N@1�G1��ƶG�7޼s��Á��/Y�Ur�2��y_s:����O�a�[����`����3� [���vŵ��6���
�ad�h
�^�Q��O�1�r�R�bX���_�R��t?��W$����kqt�Q-r�<��j`N��j��F5�v�w2�rD���5�H�I�y�$�<��`ے�Q�B,`XI �z�&���
3h����z�>GPw3\é�̸��F�b�R»*'��*�̲���`$Z\�QG��cpa�tLb<*���2�zɉ�s�!��Z��+x2W[�\���Ϯ�w��y��U�AD�lғg����8[�"�N}�|����Wa�Uq'��dۓ�S*��{�!RGhn-�(� ����jt�lȏn�t���fm���/�U>W;f�������{zw�H�Xo�-��,��,�p�x$�,��ܛ�M^>-4��bF���Q!@,��� ��H���M>Zx-�pg`X藇���	;D_��5n��ƨ�>�5@�
J��:�p@��w�+e ß���S���Bh�Y��H���%)�mk�5�5�'�'�E�8��G�{�婩�/$e̗8�P����9�`~o2U�7��#���k��ܧ��)X$c]�������
�~�qpjpǑ��}�	�e��3v�a��r�FԣGC�]�5^����L6W~��S�Cxi�Cn����"Ј5{�I��iZ?1�� ?-a��ɤǓ8�B7���_�ևp�|fSt�ɽ���б��]BQ��:;YF�+&�k�f b��GB�8ݵ��Χ4g�/�jE^��t��bg�4^L#ܥJ!�ܹ���Zړ1���T×y_�9'qϟ�e�?'��|�yM��*@D��R�m��B��pf�"���_w��Z;� 2�(�Gc	/��1�5����z�,�	�1�vg�4jm�1�\�O�/�:q^$Y�^����S�K".�Srө��%SW��s��5Mf#{4Dn�o��P"D�j6f�F����+�L Z��sC�֮=�>u!��V1q]x���CoR��|�����?�p9ux��-��8���9�υ߼'t^�Rd�A�H�շEy%���",���8A��ޒ���K���6C�zH���}g��>�AdX|1�����i��B�������O>�����y7J��&� �Z����s:NӘ��J/�3�ܒ�J��
o�j�jPZ�DT���`�aD�HnuL���:vn|E�Y_c�Ԋ�K?-Pk16�hjǨd�G2;���:D��b�x	OXFuF.�Z�eY
|p�̗�9Q.�Uik烾%�����uW�K��CT��Q�A�^�d�M�`��? �:ƒzlh
���Q1N,=W��c�� h��ʴ:�$����aS|�,�jˣ{�tK����"�i��	���ag�&��\��t9Bܕ�=88�;*qBj�ժ��:p՛T[c��T�0B����[����v���L�zP�����~�M*��<QJt��}# cꇕ���aCR����q�/�߉�}UƸ!����m)2�xl.33	]&�ϡn�{�R@s~�WF���f��7�V,�`��p<���6gGc"�����@kI;k��#A��6>A��Q���4�o~��S�]D9r��Y nQ�,P�w���IH�V�����*_2d!{�pĕۓ�V�Ôw�b��I�8
cY1����B+��nS��t�;��"e5P�to^!�lXT�{ԞਓD�p�a�U����v��t�d�W$$�; d�<jqwmS����cֈ�i�� ���#��`�<A�2U�*j��7�?��)�zXV���کc?i���ْ
w���g��q��T{�;O��]�5~��1���㿒��x�@�l��l�o"�Wm5i�@��Z�<J�e��^�gʴ[�$V�e��g�'0��r�2��k/PftD2P�w3�! f��5��\x��5��4�,}�G&�yj��m�s�E\K}�D�M鞝�u=����s���{h�U0��gfE�
诘P�R�Fg��˰�|������8 �$_ɠЌcݙ�<|-ξ� s�?�5�֓�=� 4d��F�V?�G���
A�<	�<�v��G���1	=g��z|����O�Ҹ��߲�������'Ӧ.c���,�zق�.�y��5��/�B*�~��,T�/y�H4�?����/R�Z~�%��=����tEA�nH�ṇė�V���nB���q ��Y�6K�>}���>p�� ������C���X�SȽ)���NC$�k?�"͔n���p�%�sv뮺��_Z�_�W�nq���#~ijj�A��u��v$�ݫ�{�OJRRE��6LZ��jqWz��m�vc\w��v�ޞ�Ѿ�;M�T�R(���nq��d��op<A|9@�����!�*/T�/)��|&���v%�־'����x���P�6����5ljrJ"��^fI�g����Vpƭ�:X犟��-��z��fm�0�t,����D�`����w�r���+�	R�B2��l�Q��s�� �x:�ݠ [�oYF0�s��w���"1M������|�ȓ�仴�T)7��14��
%j�:�m��"��֖���B&�#��s�[��"�'��r"�Þ*]�;ӗ����y3%(��I��6�\8��Q�a���7�'���j�K'}��=�s�)�S�κ�Y�u<�K�%c��&�#I|�pf�rfUt�>�X`�u��A���5Q/��꣬��bQ-d+ja��T�V	#����	�y��v��/�y����<xI��]Þ�d���c�C�1�+�w{��F���Q ^0*���|���B�t��
5P<gSV{-Rg��F��mj�,堟w9A��b%��I�+�R�guޣ��nl���n��M��yrܣw��*?t��yi3��{��>D/P��/��D܋Ҁ�@7'��;���ф9���bss�8?�B�ѳk�(7nm{wl-I�$#��������*�Y��f(����}�����oGk�e��1��d������b@�t
P��O$�mWV��SΣG9H��ޏz��z��g��n?ϛ)�14���a��|Ƣ���#��DX���&����P�4!t��|�h�R-.�mL[JG���[�SH�L��W�3�  N����5h����8<VZ�4�c���}X��kx���ߊ�SkUM�-i������D|w7P���E�R�� �a�U�����{c�	�A�[��#a"\�O>,Nw36�ܯۨ��޾�Fb@��}����6�l62UE��i�T���J�����;S���QFY�+F���A"g��@롅`������z9,�.Uۏ� r�%X��#x.B�-��	��4�Ryx/����k.�m+�%:n�T�)�I/S'�9�U�x���Hv��S��yS����Êp�� ^�[Hr�
�A'-uO���x���%T�/�߲73^6��"�(��VrNlI�L���S��$.Õ��59�ubÜ�����w%c�Vȑ��Iz�0�6_����{����*�*^N�lb ���>,Mt��ު��6���	��]O�i�#�(Db��Vu�8U��,Q�	��ͅ�h���������E�~#i�ޢ#�3/w�%�G8G{Y���'bo$�Z������l�pߵE���3C�`q�"���3��YطL�N��;���nn�EY�C��AK�l�D�[�S����.���6n��Q��*g9���^��X��2�Z���hpv�
gS�CB�13ܸC���(B�D�LU@-b7��όi�V"c�N�Ny�G��<M���A����7�5��6�\s
�nl#J̼�.����[QTļ�+��q� Q����$�Z����@H��X��
�q���N%��#��c���|�y.�%��F
{S��p�#%q�&��5F٭AfC����{@W'DX����3���Qo��:��:�z��מwh`�(� ���
:�z�%;���/6�Zvz���Q��0-��r�Lh���$���JM�,Pu�ڙ4b��OYV`���wܐ��t�߸���Ĺ����a�(E�#4b'	�/�C�5�L6�C�;��U���b�*Z�0�ro̜V�4�U�U�T=ě��*3ص�h��|g(GC��e�*�XHi�1%BjU�Ƭ��t#2��X������/rn�+��A�&U�����h�͓-�e;��{	S3���#���`��=��[O�8�ra��r�:&џW��<]��4�{��"�~3����@��=-~�Uw4�u��u�yS��[Ȥ����XHf8���d���㚖}R�9��*堎M���7��
ϝ�o�1��>�,�7�����̛3L �`G��xY� 	5+���a�8�Tx�fDs���E���zo�sm�*MY�T#�Ί�6:�&Ma��9/t�n|�h{���e{����n��Q��Nx��ar��\:/�ɬ@��CG��#na�iD�
s���-]�!�6��H1%f�hnp����LCu��_�َ=�WB�7��	�ǲ�qS�S�p���Cc}���l��b,|��@��"Nd9��m,=?�F��>����$��ɮ��=|(�QQJm����V��G�i�TiB���� /�5j�9��� be��0eߥϴ����c��g��tW����Ϛ��Q�[*�5�J��1�in��Q5D�=�e&�ԫә��ds�<�;�����;���c��L�����Z-N�3��8���04Q��GX"R��<��Qۘ�2�)j���M�Q�E�����N���'��N��!�����M��etH�LE�j��Rg�W���i)�Z��ߏ?�P+2)�[��Z���=�3%\�\W �)>#@�g �*�3pb}n����^�l6h���JdȪ-��Ǖ��RL@ɯ(F� �=D��P~�)��=�6Q�������3g�F+V��_�u��&L��G8����W�`^�d��=-�d�[r	sq1]4�"��gɗHe�Ӭ��n�(�R)�N�{kx?4��q֒N�u1��|3G��'C� n����4nMsi��1[��,	�T���L�)̓9u��Ak�O� �>�sN�;���N�C�`j!J) Q/8���9��)8���n"�&}�HC����)DPOT"��#�V.�߁��3�o��y�W^V�=�JPfE2���U�(���\��'�(��M/p�>��$*�e����";���t}�o�8�r;/�=��Za�G���j�g�`��9���0A��M�	�����Q���ѽ=�M�T��O'�T�G���ƻ{2aj	;Gs�E���S��rk�|����>W�Y��⼡>��I���8j��D��©�:���7�e�ٖ��ѝo�	Q`%���6R3(ܖ��4��*����ߐТ�mu�?W��8�c��w��GH���v���(�B�t�|2���+h��M
�Z���G���?����ˋ����s_/��!V뀤 u�I�>W�`9�k7L�xd��G���R@]�)�^�J̩���9@.�V�wG����!�{��n69u�X����D�_%��KO�%��)�J��J�d�`��,�kx���|^��-MYs]��YC�1�7"�IM����S��1nu��3u^k2'���c�G� �_.p������w��$�ȶEm�£�l�e�ơ��U��yzB8��{�;Jr�K{�X�?;kY��ދ���0* S�S���ھ��|4��[qM�+��	Q��oTEr����rA�i���v)��iD[��Fp>R�*�j�2�q���Y-��&�QO�CD8�03>��U�X��
����<�@� �匋�p[���֐Z�]�˽ݎnh��+_��0��8��ՄÄ&9��9�x(
@�����z5K+uC0W���3������,,�	���;ކ���)	%a���l�  ���dJr[�z����%�_������$S=�V_O��������)�8��&�N����	�B'}�� WbcCL�Ãt�nb�V���@6�@�k*`�E#���뎆�T��.�:�2��3U{^��Am�{�9�k�寖 �V�t�6q�M�y􋹲�$����Р�GN"1�-ARp�}-��,%���D��iC�M�2OH$�ac�}�HyE� z��n?d�26(���=�|��d�]f�Z����785����Pǖ]��4��{�)��q�����Ǟ�L�P{���ji��W)��7�P��4[f�:��b�W�a����J�a{A���z�8���@�#�P�1Np��.�[蠀�T^�~� ?�y��M�G�|XS�ZF�j7��Zg��d�|�Y$��OlHD��1��ù9X`�A���.�)y�(�:�s�#4ztj6& �.����<W�����7x�ߔ�V7�c4s����W�tr\��:�q���/1/w�w�w8~N
]M�~��:���M���_�#�[5�56.^�w3�tR<���a�9�����#'�d��B��xJ�)���:d�H�î|���B�,,I�Фz�j"�N^�E��v��S�(@���iBЍ��4"cYf���i����y��cIV�9n��� �8Zm��^��`��Z������q=@��Rj�f��f���-���c6]}�A�,̯c�ѰM$�`�-�K�6Xb���G\;h���F7�q\3bY�[I��g"o��v�^ۏ-!pk&������cҙ�\�ِ`�J�y��H�bc�(n/ד�I�k���4{u�4*��?��kE1��x�RVZ@D5�M#����Ҡ��e���f
����c�rH�`l��J�� t�P��Cl�3!Li!��.�^���Ǧ�n�[���"�N���6J�y�W�v2I�A�d�#��Ej9Q��Ճf�72&��R���j�k!E�sZ�;��K��ZU)8���cZ	�`��[\m�w��c�|�a��?�'��Q��I�)�y���8�h֟UI�1u�T�j
M�do��PAvHF��RX`Y��3�3o��]S�Σ���H^�TD�i�M`������OC��U�"�c僴7>��P+���Ą�X�jm�U�� J�ud�ίM{HI�ԅ���('xђM�C��g��Ds��~x��rqyVp�^uЎ/B�Y����lk��Ŋ�?�p��nSOn��a~[M$ld�J�����Y�U��a!�D#Z�3a�v`��\+��&,�/��w��Xlà�"'�`D�3�l���k�G�
lo#�߈#����I��@��H����P�n��?�G���C��XY��	-�8�ҫ��YiD�Z�pr�0�n6�/;Π��ꈉ+�tT�s=36��Y���
��~7,���ܶ�	����VU��B���/*�WLN���X�jЈ��G�s�O�1 ��:�u>�M�T�H�g0$���7���ُ�ߜ&��wT2���K����,��)�6����*��_��Z`�+}߸$�g��sQS�W_j�A�r���¸��`rl�	�/TN�5�'��\�\cq�PuK���f6%!ʐ@�U�_��e}�ֺ�m�>?_�h�y�'^'�lLd��F�����1�)Z1��u�3}��V�VC�L($v�"�w��m�]a�ϗ�> RĢU��j�YHg�uœ�,@i�B�2�U8D���H	�s&w� �T�Q��B0��%����r�o4�ml�1���~�]��_$�CրO���F�QE�"�.��S�D��8r5�ґ7�u*7>�o��%M��5�OvE$�5/��)�x(Rٜ�&Z��-V�Ӯܬm��b�c�h�qW�o`��T���d_��n#�呆RȾ �K�b��}P6�E^�<ʅm��z�̯�c�x�p14�2O���F���؅�,��0����l'c�No�3�E T%��&��� �u���}	ҤNVV��"�<Z�9��N���hl�#r\�~:��N1�m{Y��9���l�6Ca�G}�f�M�es��;"�� ��I��#�N-}�V]���}G���i��F��'��ϓ4��
ކ��k]6�:�����z48��o���$ݢ��զ�)�'�e8�ɓ��"4v���"ʚ��������l��\˶^Й=�B��Yz-jb~�TW/�h���8bQ��ET3�W�'�*�cTa���h�l�,�%]2��k& Y3��#��p��st%�[����Nz"��s(3� ��0����雒|v��ݜ�Ɍ̚q�P�_'5v��;��;��%*=��!q�[*6wV�#�t�|p�E���
��(��ϛ&3��PA�[F��8����c��p}\����e׮Q�C�ʡH����T��k�\ۥ1����J�k�{�ٴ�=s.@{ ֨dRή�˯(�~G{��U?p�6��W��ꘝ����o�y ��84���[k��&-����}�_WU>c���Q�]r��y�}B{� [��d�T��A���Y ����^����Вk�3Ȩ�v���==��ĝ�܏N͎UT�Ͼ�x�Lq0+'gN���f�lb�b��� �H���Lç�u?L�bF���-[��9e��}��Q���ȊN�� ��Gۑݞ�a�>(���n�>	�7�N�:�����ze�]�(��t�d�㯨=i�<9��/�U�]��2���s�(�$�y�\��r�U�>����_�Ze�"��<_�餎�ZP��D��/� 8���zS�ğ{�n��rw��jB�l=�H��F���ۚ��o�Z1ގ��}]V��Pc�X��%�������ɓk�r�1Y�ц*]��+6܋^ř dżYJ��l���Rt��^��+]�h/��@*�j�B$�!�M_�mI�]m�9��g�\n� ��
o�1�W%#|&�U
�*��d97�}.�gz	�t�d4�F��yV�ML�5��\~�dE��s��Q�P����Ye˸8��jq���ѫ�����tBV@�q�d�;����PM3�;,V����ЎR��*�D#o+p�Ab��p.��So�U")�ʋ�)lD��}��;�r۬�q�`=�88�~Z�� �C旬t̷z|�з��"$�U^�Wd���C�
1�d��R��Wc{%�j��J�.+��м@ �8����b.��X6GB'�L6�ls���6E욘~�)m���)I�ӑ��3��c�˔e]��7��ޅ+��2T�UZs�~/3ճ�	�,
Ui��:�EF	
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y���U� ��խI0���10uF�vG;4��������=3$�����n�C	��qD|�ƺ��pW>���?&����|dڅڰ���,?}rrL��I��ئ�n��L���5�/�����g{��Dk վ��r��Qd�H����u@����-����(6tw�������)�ִ���҈`�O)$�M�s��e?��������W��qG.��mo�yI.N��_�hY&�8��V��p�t����jY�=�VЊr�BK��[��� ��#��kSlA�G���:*wgj���������R΁�����OQ���d3�c/��p���qξ��v `\�v<f�|�
_͚c� �>తX�4��+�ñ|E>�}�H�N�� ��->�Т�n\eTfC<��˒'�&�����R��h f8�ѐ��A�5�������&�Z&3�m$�Z���E�<}����9zM�3�gt�l����i�^���:X�fg�uW���i��0���eɪ8������q���/�|2s����}66zK��}W��a���_��#yQ$!c}��L/�O�3�Bz��M�'��-��������56��@@��L2�8Z92?�_��ַ����z�2˿�D���
"̿:A~�{�z��W#V�d���P�t��p��w.��O�_+o��r�?Z�ժ^�x��8��hf�x<��R�tg�S�R<1��Z�8;�ѓ������]0W�>�~&H��]Q�.Q���[ٰ��I@�N
u~�Y���M��SPAM�[��I�R�K�����O�z��.&Z�7(D5y>���o��������LL�ӡ���;q��|=�w���z��~��>�{Ԃ�Y{���77+X';�-��9;���$w��.f2��<Z_��FB�t
ܤ ��s�Z/z�W����>�!d��S��G9%}��ߤ����w�fA�Q���%X���.s�7LX��N�W�X���0AK�2lp��ʛ��f� �ǉ8m����P=u1V_�MH��O���8�HT$k�z~fW]12Y�>S��V��%���-�^$�2EZ����b���Q��s���#����;$[*��K��_9�Ǥ�t�6�Ho��h�P���Қ�g8�G]y$6��`��@��=h1+Vi3��U�j�=F�W�K���2u�Bb�4n&�K�}����!P{=�.ҝ��<�ŵ���,�� ��'c_�q>z����z��!�y�*�A�y�P��ŏR���|	#4�;��X�l`�*���/^�'d_AW� `�m�����).��3z��V�py��t̆�H2[2+�+� ��a�(�F������Q��+A�-�ʊ,Ϲ���� NU�����fSr8$�=�]�a{�p���$�����$!K����i��w�?�?��r
�u�������!��	�����Y?ͯ��(���;���
uêO(���9{soc]�#�PO�Y?�MM	�������l@��֖�d���s�}�~���]3�{��V�nağ��w�vm��_�����F4�
�S ri����(�J��:���t�m#�s4)s��(z�� �ҋ@�=�
��ǃSzzQ��h%T��FT����N�3�ό��u���&�|X����H�%���+
˶������ O%� �n����	�8��Ot�h���K����}�5�NI��g]�������z�yR�@��*�\�T"�����1�,��!���F(��rP���� +7r��!H�'�]��QD��RB���q:;�y܂\2������6.�޶U��V�tk�/��7p�t���+8�e�g��?HM�x�ӱ��y�*ۥ����F4��G���1U0�{,�F�9�|4��^i_u��L�aЂ�����`��04���Rv8�����VeU�8Lg� o��쳃Y�a�N��p;Ό�:���mE�"�8ȑ�a��Q���w�c��o=JXQ��T-�Om�v��i�+�X�Rĵ��A��P_uP�:���T��0B�Xfa6�@��c&x�,s�0"�z�|�'^�NO�C!���	Y��p얠T5��>��rEuM��@�Y���"G�F��l�A�t�7-�/��%V2`�h������'��cw�;"c\ �_�^���e�����0K̟���Nx�>��A�v���#�^獩T��~@@Q3�L�ȏ +��l���Z����-�;��e�����A ��^r�f�Z6-���	,{�a�M��82^:)�j�^ c����F�>�敓J�U�: ��{��.v>,�\�<����$z5.-���r�k(���/�T�/���y�ޝoAc�*��g���x�����j�T������R���њ���Z��H�]�Vu�����נ)�(�ꩻ�XbE-�3݅��l�V�q�H��^{�=Ŀ����:g��y2���r��B�&y����X��M���2��+������dEÀ�zٚW,S5�}M�b�2�����ݷ�P���d��e���^�N��V�zտ���C����|�f��򜹘=	��aV�xk��BD���Q%�sP����������4���h����f�k�������%iTNR-��/6�^��+ ��K�ɀ$�T:'R ���'lR7x�09ӝSu�M{�7x�@�����E@hc�ڔf�kF��&���7ʋ��7Z�L.W�|K$�g#�,��^�v����-t�Yw����X�Ҷ��cX���j�`�� �_/Pi?e`$��ʼ�k�[�ow�p�ѫ017iC䫛5�b�!ݳ�5�}i����LPZJ�Y$9���TW�o�Wn*�?���8ߒ�#k=H4͟��S�����c�램����.߉&.N�l�{M����dB�Jz-�EH.�]Y�,(F�ٺ������!���M�q�����&�}/�mA��oʌ4	u���Fn��]��W�B����X,!�.�!�}䱓f�_�1Ƃ�w���1��P_$�-q&�R)K�Ij�Z6vA�<��f�����c�_�:P�X��EW&���)uuJc�1�Cizs7x�(��b�������=��U�����/&�C#�o�����5��R�H��[��,.v�u�E�ҺwO'��������Q{r���oL��/��
]�y��؋Z���D�S���z~��^9E��S�� X�P��r%n=^3�����nΦ.�ݵY��П�z�=H�hQ�s���7#/�G��ߏ�J�M� BK���N�~uv� _��J��
\͌=��6쨱���F�bDȏ滶�1��c6Hҗ���W��sH�L%�G��i��8&ǯ=�Do��rT�.@CY�Ve�_5/�.up�*�ڮ"%��c6X��+ s��Q:n7�=�ww� �*�T�7��5/�Ut��Q�r�(b�,SЦ�+�	�Y�ߢ�X5 ���0��8쇨 a��&��7�?-6�ƎO��߯g��I���ޓ���J|���	a��q�Dzab����8�?�jGH_{5��S���u�'��u���y����C�0����b�@ڼ�\`��:��S�ι�G���/����1J<@���ޒ���'��ֲ|�ͯZo�yN��?e�	�f0�N�!+�mxEoCj�h�����7���G��'�k=As}��h��ë�˅&لe�R妙���翚ǋ��Pq6}%��;/���*t?�o�����'6� z�^\��ą�Pj��R��>�!M 5��De��^Q�
��6Ka�TphwŮ2������"ZlQ-��s�ɅRE �t�@��'c��@Z�lF-�@Ӄ��x��煔��<~BJs�����Q�说VlD^��^�D�/��u%����8ytM�뚶t�aE��L�������fh�%��L���$�St���s���9��(���jJ@�0�:r��zq�k-t�V4k�ȩAU}z.(���-ƛ�l ��ߍMM����bZe��?!4�RZ�V/h��:S}}�Z��F��~���	@��X�O���J(�XO,��@���%���7�Wo!�hQ`�3�	��l5��0p�$NLO��k�_k&�L������_�ks۰O{dc�Y�_1�d��В��c�X�(�,gtM'%f\��u��1�J�։Κ/6�a?.U�������n����sU�=SGlR�oբ��wLEF*�@j�Q�[�U�Zd�a[: ��!.)D�ש#ț8�v�N���Fx|�򣷿��H(�`G�|.R]m�9W�����t�\��o�.��eQ�ix^"ԥ�E�w�a�4A	�n���V-�(2�=�z���,�Q�o�
,"���%ſ���ַ�[�n��tpi�Q�n��<t�+�`�?����.0\O�~� ��D��t	vgq ���2;�	*�1�Z�����lҷ�~�Th��A�F�?�-��_���uzq��_�	H9�	{$�lϻg�1<p�@��4�8;ggTݩg��h���6d�u����Jm�\e% ���$�/��3	�� �1h!��$�o���Ԑ�ζ&���_,o���P'�X�7��_F$.uNK�A, d���1)��Wu���|E�(����,S�O�7��ŁI�̩�X�뮗��mX�bF(}T�4���xHT�5��CJF>D�W=�e\���A%��X���ZQ��ZD�T,�VK�y�+nB�D]������),�����Ǯ���.y��D�8h|� t1|Eh��C�_So:�>I�/�;��lH��'2�w���+N1��'U�B��W�3�c�{���}�B�="�����{xIi��X@��='<��G+�&�P&䃨ם�΀��w��&�y��<1��}�t��2'����2����Z�.
0��|�� pTRl(�	����)ϕ�)���o~���^ؤ�\�p�k�#opȳbz>
Bn7fU���K'�x2���d��lk�[~�
�Tl�6�S�JC�����3�Y����6�=�$W��)��m²s�,&��0�;w�|q.�Y���q��Ԉ
��'^�PZ��9���5����ư���b��n؃XBc���Et�P�%w<߷T�?�7��TtL��-��.���q���{�O�bso��`@C�W�v��)톨�T�*v>�I��w�.9�U
Ux}���5�yS=o��)�Nk~p�A� S�^aQ�\�ӻ�2>h@E-K��$"Q�f�qq�[�d�g�p-ɲ#2�/to�o-vCÀ1�V�(��H�岩�i����<p����,#�r��Pe=|H��a��P����9kfh�h���[�LS�wq�;	NW�vh�y��C�)U_2j�O����-��fq�׼�Fb�WE*^��ȹ�?�[ʳm1��=�浫��|���o$�!���4j��rLh���S�x��	*��,;4-:��*�� v�rЯ/;�>)�)��l#0�%ye���['�[lp�k���7NE7O)����!���y�6����#����gLh��B4���ס���4i[+�}���\�: �'��ŵ�k�H~����Ϲ$���$p���"1�\���*�COӽF�Mh4��sMYR�'��?T!��U���ą�g'&3sݔЈ�'� t1F|�R�g���3J~��o���[:B��T���Ѧ�
�zt�K��|~���>[�u|_�c��z�1𦅲���M�8�G�=H��H�A�#�2%)�ű����t�TX�����n��z�(B��f.�e��e��~�-*m7_G[�\���&�^�>�� �k�3��C]<g>��ȏ2�N�G�V�=�K0,�liR�	{[�"�_i1#<�n�\�Hb$���G6��dz����P1��!�\��d�yG������>�XD�#ۋ������)V�(�l�E(��Ӄth> m��6�Pۺ�_<⫕�:�2�5�Ph<�Ύ��z=u
������J��&p��g���q��x�!�G���,�z�D ]s#R��Ѽ��*�g��>l���ëZ#�g+g��)q�M�L-���`=}K�Y�!q/���_�5/P�"֪��jV�i��X؛-��j�^���-�6o����W!��q��=F�n�c�.g'����X_�0k0&f�%��xE��Hnhژ�ï!�	A���� �<����G���T��[�3dQ�oRa�h�6���{����Q���'�Z3��߭!����=����:N�dvM���|pJ��"�Wo,�4��f�����2 $���"�[��^�ga�h��ll���]C�_*�Կ]�i{���n	K �w�N���Q*��b�� 5h>D�[���P����y9(�	��Â�ǑH�i#��p�}z6O����i:���9�� ��V�1��� �zip#�j�0�ɣ�^3���*�(R�z�u̺KY�`kȆ�fa����VeY;�ᩂn�����Mn�{=�O
�2|n�rf��_m����H&`���!�����8�w!�`��{N�E��33'�!¥=�10��"wcҚ���2��7��g'E��K��倆S��|��l=u���MC�WGÈ��]�։ʿ�9�Sm�M��M�i��u�@}u�PȂ`)�bY�G�)�4Z8\P}H�Y�2C��}��/��_�e�`�1ye�x]b!'*ׇ��o_�����<i�����qUGTsRS,頙uDaP��<���rY%�E��n���\5�AR��4�a����6�z�|L�b͖h�����N���Z1'�M�؟7�'M	�����a��y��{�$��O��mD�S�	�Q�������9�$!�N��'p����t#���4���\/<&> ʽ�\I�ĜCM-���[�Hh�1*ME�5�t!a�u�<�s�ȱy�<tU�^�2V���a�?����g¬ǀ��^�s}��$ "uߖ���*N u}2�9NXH�����d��A�yY)(�[c����$8��K�z��2B�����Y�c�;.��Nx�E"��x���G��?����'�`	�kL���ۼ2�z��N��j��\:����%�rE���y��<%��>9'U@�mX�3���߈�F~~�bY�S���n�wߦGnkIW�c��xL�%�JR�r����#�<�
�6<��$F�`�14�Ama~�V�"Ãb+Tl�bx��}AZX�GÅ�(suPn��ݜ>����Ce���]���ǂ��L mΞ)�]y�`X�#q�q�T�:	�fcc���n�LmGWap)s��Pי��G��M<EC���B�`��GO-g�=����dt����y�~����1qb�w�x��
5�Z�̫>�@���!R�R߼7f.��8ڀ��a��Ė`����>Oy����$�E(�X��A:xi���	�گ�5����r�����8!?__�:~r��k�HS�N]�������&g���ȓi�G���Ώ�Q'0���S�E�nA�uz�)3d]tq�(֒��W������3�JK��>��.{1�Mk�=��Pʘ:ͫ�寒l��D�������F��$�#4�q�+Z��R;�~p�@�~	J G��_�B6(�ibZ�?ŏ�����ڼ��z���6����ɜ�͎�Ջ-�ax#N�`C^���39:-��~�JIP��� 0zRR=gߍ7�� ��਱��b�C1b�vB�N�L�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�M��T-dV�Ze٘t�6ړ�MfTA��ȼ��p��y�Ofdd8Lz0q�!M���),��1���-o�d��=��
י!!�k��ˤ��c2e�1��}[���N�L�n��ǚ��������HAr���36ji���¾Ũ�	����3������ŎU�AW��	�ȡ���&�4#�N�������2��K3U	qt&R��N��	��&��./������D}P䁺��2�Afp6�Nu�z�Mm� -K����lU�z���K"�@�,��z�uC��9I��@��>ﵹ�vՙ�`�t3�݀MW1&�!H���LatM�U�C8�4�E	�O`NBz������0�+���y�����U{x <ժ�E_ҚpØ��O�S���W3qcmu��HЌh�P���,�������ח���K��p�a@�Ү���o����w�i��q�Rh���)��t�XVZ�9�k�a�C��ipsҢ =�B�������d�3�D�������Q��ߜe`��e�	*�D6���Vo+
r�"u
�EU*��f�c��UE�?��;qU}�%lԎ��}*vk�y,|Q>�l��x���� ���v�&p�i�c&,@�͞e惯��M�4����r��o'���U0࠹<�TLZ4�M$��FR�<�dk�U�b���>��y���g=8�����V��s�p �oc�{�(]�L\�_$:`��W��9�ϝ��j������A�,�;��q�6)��Su����� p�s��Vo�Y4�����牸��~u""_��P���/d>S��[2yu����Q�+�0sd�ȥ2�����0R�;F��	��M�-��`)���R���H�����k�ʇjKђ4R�ųr��- ���'��u��F���������CƲ>/G�b�����N��D��27����y}��#�C�
'�,ڣ�LU�jسq�ִh�\�(��}�FQ)��%!OO�'���M�>�����i���א7��s��hb�dn[@o�3Nz���P��=^N�7w� ���c�]b�o�)�ķ�.��[�ֽ�	k�I�?�����Qf�7��+���2�x���^6��x�r�e�G�Jͤ]L�G1`yg����\�lKu�zU���D��+EO'4f'A���k!�`{._/�[�oh��X�ݟ���i�(�Io-�o?���3R�2K���Эk�S]���F���{�c�:�ܲ�7��<�z�����Ff���L�m|?
4C���
��e�G!���h���iu�Β.8w�<�O����'_��'�%B�;櫤�.�tI�CV)7s��K��l�La��zÚ�;B�YI�Qd�����C�7�592 g��Q<�!�V���N�f_k�"�2��=���#,��(U�PT�h���F����-�(�\�8�s���~�Mr��/�b+S>��H�<�f��ٚ�AM[�<�Y,
��V�����;�ZNQ|n���0)���J��z���tL�~ YO
�`n�c��A���������g腊����q���90N��D�p�}�� 0+0pqn˞�����m�$C��/i�j�"#��8�교,F��~O"ek~9�o=�Y"j���Uu�y����o�ˍ"��J��L��=���-U\M���� ^�p=�^C��qh5 ���h6�FA�]	��=(�`7+Pt&���Y�C*wҫ43S�p��.3_ٶ��{H��Ts�N'�F�H��������S��È$:f����GF�tno�� .,�����F&4���}"��`�.���������dm�`Ȅ��������%?T�|�Q���b� �^��a���ٔ�u���Z��K��X�!�j�B`a����I���I�j��OT���]F�7W����E�@ά�����;�H�	�78�s�;4|��$��b6*'*�����N�s �6�h��?"�}\�k�
(=�����@�Y_�R`}8q�B�9=k��Xd䍻:�N��ڧ�ʃ�I�U�8N��B0�$أ�w_�w�gW��W�J!t�d%�m�5=!)ѭc�r3z�R��2�$�=�E>2���T��8Hņ���9�n����'X�M���_R���;�% S�g6V*�4W��E���4�(�G�%-��p�=b*�{`����c.��@i��įL̐�|2c���ꤚ��}����w�{s���{�!3-��x�p���1Ky�W嘞l��y/�ݸ��r�]��G2��� Q!)C���@uL����	]�S�g�	l���cW�׺��'��htO^nW����pڼr�Ot�L�_����0���q���m�E�@^�
z�θc��f�[��\�ј&�Bl�ň�snPm (�ބ��J
��h>����^)7:l���Eh,e������a��M���٢�;pg�L����o�����y�:{y:n�%Yu�#�k�����	l��Ȝ�����v��<dG�L25�Y=����էs�dh��D�;gv���Hj���M��-G�#1U:��s>o^�I�!�[js���Ca�ieg~�K1�"�����M�^�x�ܣ�f{��Q'e���f����|��X`�CJ��T�s?�N�u�!	�_�%1���_��|P�A�������#�������~*��V�{H���=���a�z����붕���U�����=���Kz��O9��t@�lH����ڟ�������c~Fs8�|�Q�~P���W4'8kx-�
�x�\Y�_p>I�\�3]p�4�`��+"l�L���)��Y9���1x��Y�ɒ-G��)�?9NY8jI.9wq��B������G�)p%�?f���|zπ�.y���_,Pb� ���e1,�?�RqU:����=��4Q���ȍ�:dlamJSr:�Z!)Tp�W/�"&~5��I������ �O�Щ�t1��Ԋ��6��w�r9ڪ�X�_"�78�q�t�<I<D��A����0b�gr�D���]n�� �Y�)�U�W���������uŀbJy�a��AFSRu��[4��̽ͤ�b�>�
�<.����a�1S���Zʎυ}��H٠�Z�J�4�h��j;y�<류���᷵B�&���aU��͂�0z�+����2@���� �h�&��c$�$'�ԃo�Ej���?AZ&,�#�}�;7�0�ā�sM�>��q?K]�R��^K�Q�e�;��G e�;�̽B���m-__���2��A��MW�VD��X������U����7O��/�"aIyn�͒v����7˃yZA���vT]�����/����|W��ju�_ST�\ox���<�N}0�ܦ��<'Q��o��@#A,f� r��8gU�o�ՀKT�sJI�Jַٰ����O�҇b�qj�7�ԡ��55f�7>�kv���
O^�-�1t5er+���Y��_�7k������D�� ��?��@@�Kx��_��Uۦ��=N`sx��PRs0���+N>)��=����)��^�4� �Kn1W��@���A�8B׈5IlW�I��[�R����%7c���ֈ�ޢ�^��}��:��`~SK�-�U���+���
3h��\Hې	f��e��� �I��D��7m�'��R�U�EhQ����Z���u�X���	�����u �-�Oϧ�e �f�h�;��r����xi��F����;��왺��ݳJ������f�݇>�&	4�d6b}Pŭ�ᑂf����i��r?2B�{6yͣ����ua�9��d��r��s~W[|���#K���U�k�37'�>����ؘ�6Ν��?����D�L1%���,(�B�a���Dh��~w�Vk�]%���k˹{�P��\�~5�_z��ӊr)y���
�]���gm4�����wn ���0���{���$�	��5���l}4j�.{u5�mT�
�fS7�K_�΀�@v�듇�J�����ց}��%�`=w�ꓨ�IC������{��_X�z�ptK� 5�WTgb���SP��a��C�_Xx�����S®[F�"v�O�3�z�x'���2cv�
Nj�]2�w����ڜC���Z�\CS��f��z����ή��	/��M�Jk�f�:�^g��l���]#�e��Ů,�kmw�1��R.U�{l����αͻ����~��̟��=����y4�$*5�ۣ3�bp��w�*�t�4JR|����]���O�)T�����0@:QmcC�e㢂�C��}4c��=��z C9}�F�-lH��i�����M�"���^"���6?��]k�S����1��Z�V,�;���)�<x�p�K�m�����]T�Ef!cޢ�����?��`�2��9��޷F��=���\�u�}x�ӐY�S���@����E&u�yZ𦍘R�.ި���5�Q|�)�	�Q��=��k!$�Y�4Gm6���K8O�x��y�e������u�ykO���B�s@�?���s�޳�L	���3�f�U��Ho�4��[f+���D�qWB��U�j]�hy#[��3��?d=�r��)-�U�F�=��*	F�㣙Zu2���?Z��
���u�\�`L������fٕ;+(.J��+@�Jx?y�/hh�w�'��5��?�R�ԑ��#c_�R��!�F�C	�,���B�!�j"fI�[Rx#O4.E����%��r�J���?���
���n�p.uD/ /n ��
��l$�"�)�
	��P"�_�0�`���P���F��:�!�?��(	�ǈ����ym2��&��%�|��rq��!{U��)J���U���a�_��ġ��*��,�/�'����"��<x1օ�J
GkoC�u��:;>Mm2|wP��&��<HF��C#��ؠguuQ�sO�r෰�3k���toS���$+�-uֆ�L�r��'���6=�0�U�D���=P�RIbm�n,�i��=�`�68����4������X�	��H&)����-u��[e�a��X%��8:`>f{�G��F��8pa��uv ����r0��8��8�� i�lX���r3B<p���Xd^�>��{<*)]-W%rB�i�g��V��b�C'Ώ}�b`ig�NR1.��-$��|oIYK�ޅyf���b�G�*8X�}*׽K�4�yA�V{������(bz���n����t��K�0&>�j�̎_yc,�`4��hM��#�2�� �-�`���AU�[�q�]`x zT%����.��9_�#C�ә�?s ���Pm�j�����oM$� r��!��q��i��[H���rr�t�1p�yTx���o@�sׅ'�}D��И~�^������l{R+|�\y�?Q��"%�l��: �S��x���X�PΩr:E��R����i�'�WD�^����0#�h{r1� W�h���h�!b��
Ĳ7f�$� �ltV�P��������Ȝ�kI)aX�89���n!+�-UqX�1a�>�l"&֑eX���д�2ރ���� 1�U�E���}���4+/~QhDw��b�����Pq��kt���@���N^�<':���<ުA?��
ze`JhF��9Wt p�+�F��7��wԣ��C�J�)���J�{��G=Z��(���(��/V�ޫ����ݽ��R���lʺn]X��P�M�е�%x�{���a�"�K"9 ���Hsmm�VU̖ʠ������>��&�^6��I���M&�{�h�o�)��x)���?M6%�!F��"��f4�b�����6��26b��(�\ėQ��K��5)*a����D��]��m?���1v�S����jR4L�b{�R�Uq\���-0�nyʤx�w
�hJ<���j��a�Qm��r1��&����R�������R����)�8��s�����GUׁ�4Ұ��p�%�8�-}&����;єG7C�!��"�?O���jsI?S�͹f ``�'�x�&p�145k�Q�&-��ôU蚒p�%�Z��L�X"�O^b��<)L%ds��ɯ��Ư��
h�89̯�7H��[����?�T��ӱj�<��s`�ҷ�gV�Q���A�k+ݍk^V0��@�]�~��[�l���x*p�V�Ll@}��ϟ�֌������������8����H��,��8�7�<�	)S&��J�d��f��/��ݽ�-A��Jf�"y!�.�1�bo�u�h:4%�M#\�v�ۺ\�z¤5�W��������:)��4AXcژ�� �n|mS aw��(���N�O\s�!5�Z��`נ�E^����tvA�Xq/��3�J���?n+��ډ%YB�{k��Yt>78F��)b�`Q�!'�pO)�����xE�f;��<x����������f��$k���"�i/t��;�T�Sz�����P)�Lcpp�����`.�e����x�������4E>~(k��T/6����3�Pg�w��<��5�gS�Y����BtHvЙ6��/�PGx࿱V����+:�^��SF�������:��� la56l�C�7�7F�9f��Ǉ.�2[�^������uh]ؒ�U�jʴM�G�6����&tc��;�P�:�[W��+�?��F��zR���@�|�b��\!'hw���%�	������!���	�_��� -<�����c<.�@���2k�n��T8�p�.4C��x�Jh�)�9 �`��C��*e܆�W$�@B$J�6���X�`.)#8s�7�642v��c����se��j�cP��&�Z���<���`6��<�y*��r�O�᭡p�̿�Y���(
�J���}�]2�y��:\[�N�f�E3Nas�������<�)��׺��!����>Pi�m}x�3y����&,>�5�,ڀo�,�M�)�� ���U�� U'����QF�+d�렼�jޭ!��t��Ҥ��w).#���OAZE���&^S���U�rPW���{���H�i�+>m����$����W�Gw���H�Dǈ�#c�P�9]�H�N�Z�0�Ym�c�G�!^�yY*H=Gg��
n���M�%9ٖ��ye�\�RD�_�^��S������d��%kO��3�u9r�Z�`�Jd�x�L�Ȳ��9C����w����I�\�ƅL���ˬ�d�2?8�y�+ޔ.��goE��t	��g"����j�����%v'd�V���]��!$Y��UQ��]yV��!?�B@�b�d��*zI��w�ևE�yT:�&�^�h���+}�o��o u,) 3+�I���o��:�6CI��~�K�G[��/�^�LH�K�Ai�N�������pp�do���.��.��;���nD������@a���C���5�JvUOBi˃�"�h!p(+�U�� ?�DG��כ�1�S�/5v�4[)��@*L	�9�����=w0$)Q۞k	x}�9*��n�c��O=\��CCb~�ً���)��4g�	D��P,̻9���c3�^q=OY���Q�T3(*��g�Y������&ͻ�q�j_!��K�MR��4�/�����R>�D�9�9���i7�Ͼ�WȜ�\��ZgCL������N����5�bR���1�>��dՐ�Dl5Ȯ`�n^%���1A*��z>Z��~��u����V�� L}R��ӓ�\+Bv� ���<��C}5���յgW�<�|�"˫������ ��3��0��N��ȹ-���
"�3�NN�D8��NE�ϫ��yr�3���A��/����v��MA`���̉�� ���6��cW���%��H$XAG���3�,�%�H�h)��1g΋M�N��N�_@�W[|�����%��N�;�X�s�ic�'�3`!�J�ϮX��@�(H�n�G�U#fT-��[���q�iS:9�z��P����֢�"�uR|l#ia�O���:�yJ(3��iO7Ɵ[;)�0��w�1tF^�'M�^O2���\��s�Y8]�h`,�+��/JM@0_��?/o��ԗ�vB�G�f3֐l��P�(@%aO竝i���G´jK�_7�`�\t(ľ���=\�놎݊|G�;i��BM1�7��N3N��ٹdgNq*ET|"�����Mٵ)�}z�pgV_./�� ��t-7&�s�%�z�\��(8<������{k����"���TH��y�����P�g`����5�1��9 �%W��	���|b�K�qeo�#Df�Z�7����cH3K��s����O
:O�)���xgހB�����{���a�2��D싞�=&E���RL�$����������uM�N�$�r�����D/�	�o����W��z{x�[�v���q���5$���Yɑz�nj4�ׇp�K���|舆SL���dJ�	=�k�Չ' �SVR/�\�i�ǟZ�C�r����4<���<Ϗ T�F��ǲ����_ K���y���4u���л��]�`�wv�lr�nC2�3���!J�d�=��E�
�R\��h[�r�$	H�SQR¿��A� Ir��FDz$�)�a��Tߡ2&}���dw�-���9��7�i� �F�Zh�<E��9���je�x�"����N�i1��!Vp�p��{,Z��(Zy���EN;d��D��ܥf̄f����	 c|��eh��O���b�(g񵛩Q��2�����<��J����!>��׊���ŉ�A�6{��^>���T�&vf��ĢX��@�&<ĤSnJWK@Y�f!d2@2�N���L��ͯΞU}Ql$��tX�*YX�`YSX#.�c�.��4��}�q����23d��D��R���FY�T�!ź(c�sAH�l�����]gڊ����Mw:�N�J&��&��e�WX\���D�_K=�	�2�k6ܮX���Һ�p�?PA�Y��Y�ϵ1ᒊ�7m��5k��mr%Ƭ�B��7�A2��-7/{,%���f�]ͤ�)ށ���3TA�4�H,+f�@��@Ն�L�凰M.3"�i����䩣/�a+D���S�*��Y�S��R���h"�B>'gU2�v���W������YY�ԻĲ����������1v���Cb�Rr4�֧��L����_�3����y�=��Vm]�n'�����QD���qD�ߣ6.�'`�:�_H�hH��DN��+����Fa3{����Zg4)��U���t�<r8���IutxB��Ƭ?�<L<	��8)���R�9�ƪ�{��$BO��>��_&89��_�aŭ"��z��Qe)�y�0����:��}bh̬��'6�Y��xH���̋H�G.:�T��'���ǿb
���,~�e�Z�J��亣�$�?b�c�^@��LMT����i��l�_��5Dγ�U�A�˹�IN�T�Z�7J�^�&��֦�:p�^?V��:������9~�d.�N�w.�65�\q��5査c�
W���K��N^N�-K���rP��&�響�J �� )�Y�T�����0]�>�V6�18f$JU�C��Lg�'�����[M�%�;jI:�����Z�_"y/�f�������zqF��z'7��q�Fb�L[���`W f7+p�n����b�M��y�zz}�VT
�3U������y�^�QC�+1���{�uh�Xql�s����ٿ=H��?�w�웑��Q,�S2�� 3��Ok�ֆo\K\��#K9�ђ\�W)-z����>��욕N�[w�/O4���ح����ok�m�'�R��� ��9jPQΰC�Z��;�ͩ信��)f�H�]�/���h�a���L����o @Ux��$��pSt�˞�ak�,�
R���x���9�T�a�w,٢��.(��J[U�4r��C���@�E}���
��P\A���������bm��z� �Bͭ�����K���hI.��%����z*���1�{��b�����Z�U��w����r���	���T�����i��շ0��d��F������56��e�� �D�+�� ~-">7\�j�R��
��ɵ�Z�l���'n�<Gj[�Tr~�!���o�)"wE�\��p��JO\�_;GD���'�#1��E�5���,�է�s�J��X<
@�?i�(́
�M��C�l���R�򑎞�F���9Wa�qQ�ߗ�$�b_���&|R����2�ii��CarY�)~o�H�di�4h��?�<�&p|a���V)�MP��^i̝	�,�%<� _�h��΀z|���R�G�;�"�ů�4{�O�re� [v��x�rg��h���	��4�k��%�����uv�T�'J n�G�`�;#�P����N����oE0+���46��u^�����:K����po��H�2}k!MTG�[u�+1���p9.Y�ܳ�F�� gM���z����h7���8�w!�������$*�V����)ǍS�f�Y����9��$ذ��v�悠�@b�pd�N����z����P�.��@�@#o���Rj����߼��|x�]	������<8�����K�܁v��Vc��q�i�)�P��8?ɟ�@">oZ�҈�5<*�qm��
��# ?>�vB��
�@'T/Z��:^�rl�0��}�r|�Q�6�vk�
���%,��]U&"������c#d\zV�YB#�7@N����S�ޘ��h����q�,kY���J<�"�(Ҡ��L,]�y�nu��� K��J*�h����$��W�̔�{�1%JeO�`�L����wܽ��B	���8��w��ku�,�L��@^�0� K�MP��Vg�H��Ζ�d.|1��ZD�tDNk�>�*�M�??.h[��K`@�?S}�"��J�k��S��Ұ�)tR
A>�7l	���\i�Ot�˧ʈ�D�L�g3;�b��l`��bKR��6t3��g����v�!���a�s��H���K��vv��;�0�|t]�gS�Sp?�k�?."@�Q��]���y{3�B�JXux�]�9&#,�����g�z�t���f�ny��d@�ؗb�����n=�y⛋ৎ���tF��"���<���x�C�~9�ܽԈ�"�Ӎ5���؇'D;\�O�и��L[���a�3�Q�n��	�@�����h��z��.�~GF*�5�F���gQ�e�9���a���/a�}��gTu*6��<[�W��2V=��,8B{���Z�P����QT�����G@	}��$ $����m$E�S!9N��4�ߗg�r3Q�'WS�k��t*��hf}䓈ߎ�f6+���_�h�"Ӹ����Lj���� ��LF���b7P�RyD*��i0*+�:���0��n���IC�$�% ���7�QqM�Y�A����W��#}r�P�8=
C��]�&�N�J ާ�߳�Jם�X�pS8�>���7��z�5|$�N��u�C��Z4P��_��mh�|����W0�$�Ni�����K�7ef!6�.畓���y|��fCc���{V�~8� !��1P4�_'������
��;բw5Y��p��^dt8��ւ��ɵ�q�5sWa| �].�mᖷ+�wl�X�'L� �j ��Jr�B�u�C���?
�=� �٦0F�2}�+���(~s{k&m�^pOC����nwȿ�j�pR�Er�l8�Q�uqë����r���X��{�c`�����x������h�F�`ESP�~V�8�5L;7d���#Z��M_3���|y�n�dTC!,���
B��Y�,t��ug1��|?^f��f�p��
��H�MƳ:!t~��V�E�	B��8�V�����w��2$���K��B3��S��5���٭����"��<��1!�p��&̷�Pz9�(̛��w�ϳZ*���R���
&��l�ݪ'�Q�	r�w���]�tO��f�.	�sZ,�_$tK�(刧��$�֑X�2�d��tnh���&^��!a�b�Q�P��p� �k��e�T���^]A$��Q�tڏ�J��JS�$�wu�XXiW��1��ucH=9a;m��F��>k ��f�e�iOB�ͷ"}Sg��MgA����9`�	Ɲ�A�&ԅ���������N�C�Tr	D�Sa��[%~ퟖ�-������o�N[pY �7[Ai��ʀH�Q��Nѫ������>j�3#�w �up[V������to�h��m?�����͈����$�2��uA�\~:�(�͊�VM<��{�M<���ϲ�9��^���Qn��K�~N������i>�|0
���:�؋�R������ܛC[���G�s�f
��ШX�%���������0�ڀ!t&y�
�i���Խ�R!�u��ȪR�F+\����9�,�I�
Cĸ-���\{mg-?PT��9�C�*p�j�s����i	�PRY� ����}�HF 댑:S�4P8g�땇f�Z#��H�����w4Ku%�!�YI���3ߕd)F�[-���tm�Ϫl�Rϼ���d,}�ߍ2]�N��<R@p
��͚P2:�vG7�=�!Du�g�Pt�"���9�'¢����@����E�:��D ��h���W��N@��O�ЍSE���FX=_��c6�PA��gM?�Te|���;�o ]D�=����"��1�v>��R����b�]��!�܋�j�2��͈8&X�lN��h�G�
W��Ơ)�q<�E�zLY���TS��4�ZbF/mǢ].��0�}���I()~!���y$��7~���kU�*S���[J!`�T`U��_��~���������M��[�&^���cv�΀	�-��`6���_!��)�s�=;�@���r�e*��vl<~�ܖ+��]̶�eYq��j�\���ɤ�������N��TnF�oi�]�����������[d��xh�8��!����>�>�/s��7f��R�g���Ȼ�F�a�<��%R�V��	6�MDF�×����eEr,�_y��e��B��o]��Pa�5S>u��3G�QO�{����O���&1��/�CkS5E7�\;BGu�yA��#Q�2��%�<�� �pwU�0�a�ц�F�ܗ|�CC],Ȧ�X�����!Z[�������[%i���l�˒���B��$m��R�!�f�/�mix~� c
���Wp��Q%�	V{0uH[����f</>*�7���0��%�(���갣������0տK
�_�kZ,wI2�y����H����)8qyԱd�KN��UY���B��W��>$��c3vXAC����.I�|�"��� r�,���ꨕ`�۬z娐:8Ѫ��#��"QH�aS#��w������' £,�E�cL<��:]Wb��K=��k&���_w2\��pߤ�/-����;�O�c'�	Ģ��$Z�T,���@!�j�bZ�����Fй�������Gt���[� �Y����VX�?�Ѹ�+���e���d�	��\+ұQ49Kѯ8#5���р�,B�&�|�(��a��Z_T����-(@R[z"��4$~c�� ������YpGm��p���z�� V��Z�y��EFeN$�
�#E��
�MlŤ(Q�5��,r�$S���C2sS������?��]ݲ����'9&b�L�}���f7�`�_u��� mSi�U����it�2�Wu�P�W�N��I�B}���>�rG�ӻS��9έ�9c	�w֘��ߐLej����JY��I�۔�2�.Kp��Sq:-sK�V�Z�ZMȶqw������t������g�)r��!�5���0S-!I�Q˩X����c��6^���C�!�m�M�2� �P�-m�%��-:�k�|u����
�\���Z�޾7<�'x��jD{�ğ�08?^/�=�]��t[����U�.֘����g� h���{2��[�q׸]Se���̛��8m,Rqߌ��3
��d�W�1~/�\�}��?>0�bY�^Vɺ�n5��*��^�u�ՓE�����>��tw#���<���jӍm���]���0�2��3���a-��_��Ɂk������ɷ��<X�lXn�r�/�p%!bA�
��dÐr�Iӥt�e�V��
�������9�$ae��NPy!q�yDQ��2��
)=�m�9,#$��0p����.~��}"5�B�>)S�� �*����7�m�JGYrr�8���K���f&ڭ����У��?	~��+���B�̂�����|N!��hPD����3_��]C-t�����*�%�|�2�LZ���i/�y܍�uu�a~]�D��T2�b�ӃH�lH��
y�%���b=�r>&���6���*���o��
N��gzJ5�����CπR4gEc��܈�&j�?ʩ�����ĉD�`vd�!����c�X�L��3��ƴ�������~�*���p�b?δ\�l���*�Ɇ�v��Ѯ!q��X��n�<@R�����l^P�K�./���H�͕��!t%�_T���<�!�������
����Rǥ��'�����wF�����6lF�k�ۆ�v2���/�+��gBQy{E�P��gkO8��$�P\����/o�;Ģ��)��a\BL#JT ��&�JL�ש1�L��AiF����>9m)�ml�Z�#��2xU����t!l�y}�h��G��=�D�B�f�V���Z�)"�q�U�G�'n�e��gI�Tn����gF6ڥ�_�,�5���u�i��9�6{a��c8�R�s�h�1m<�{8)9Ӛo��r�#o�md�������NUi�l3���wS[A�Б]y�zNX3	�[�4�R�+�{�#�e�E����#��o�gJ�3�R��p�ȫ��c,��Kk�P��W�����p��+��bX�U�L������8�R�e��G\!.=��Cء�e��3vM���:�V[*"��v�����j-�r�V��^`�Q���Nm*��O����9|և/�С��G:���V#T��Ԃ"��Ln"���Swf7>��0�����s^�'�ٛ�ϒ*c�"��Î�)A���el�Guy��Jw��c�5 ��=F������<���TXr���	q8���((O��B�C{Qb[�8�h��K�ׁgK���t�+V�$)�֔,��a=d{mR��݉ϳ�Q)"�H��rH��֋Z��9��%�4CDn�`����.b��a
뼒����B`���p��2
�Ά�PY�m�0]F��!��QK���Z6���F�O��՟ف�L���Q���G����ib�R����}
�vH��Ld4��;=Dp6/;�� ˡ�rSq���s_좗�-�J�Y�S����7d��&W�\��֘�/��Ŵh�6���W�y��}` ��x
 ���s��[{��]�?Ikvn�`�i7�떅Ԋ������๽(tn0.�/��w�}j��e��չ�1��V�4�
�䂪f,����o�nle'2)���.�ڞB,�ךi�K�yK�=��ss&�⏖S��J/6�Ztk`q��a��-�L�C�_���>j|w,&�tM�=�21�� A��-�^J��� T�d�Q'���0�N|�Y�T�l��~���rI[�7�R�U�e_�J�.���Q2�k2��r����2��5�ت�7XE��;H�n'�'�A��]0G�>M��B|�O,��P@�JM���j�;�f����D��e�Yz��[������8� �D����
{��W�2*L�*�����z�)���ْ��B�\�nY���!���8��Q�������\��.'����C�B?	�����HIW�:�'%�qCES�������$��yd�5�F��H˚C�q�փ��P,y���4J�us�7�R5'f%Γ3����)��[�La�){Ǜ�ƒ�N(�~�?����cXo��8'��M�U���N<E%�p�q�e<K���<��nHbF$2��g�R#k鐋ĕ�M�qcE�F��^
�q�=Y���nlh1FF�)sA���	�e�$�V�y�ߒ���8�Q� �׷���ɝ�Եzbգ�x���u���C�6��n ��	X&��r+8 ���OG��>��,����P�����vH3����#��Vo�Co)�)��F���Z���iF0���ے*���s��Cv��E�s:�;hG��hý�Iњ[��d�--�4�F�H�L�l��o�����*oc��}��� A���s�V�;:�	����Eih�FraS�4��e��[.<��k��jɮ��/<4�{�e2k�ޘ?~��6W��mz��Dv]�0���>�� W٘˧=��xS]}�H��_�gܼ��䉄�^�#2��62n�O�Z
�L2�|\8�8t�ԃz6�n��:dV��<��&U����V����oZ�ԬV���s�B���d�����r�����w��T�v ��	�O�	�+�_��ˡ�.Ć�6�2����?O����"Q@��=�,�Tc�T�-$pA�lDs~��g��q\����G�qƻ���[�p�����</�>@]��N�ޙM�QV����4ɬ(Y9���0�q�~���R5� ����k���tH����	k�m�ܝ�y0���˨�p�w�z8����e�o)b=��tdI,v�V���|��b�R���?k��� 4Sm#������?�R�a#~�2&=7�k
Sxj(��R���9���(2����o؂{�E��)��<GJ9Cg	N��e�Զ'C�,{e7ߑ�g/t��R�c+BVx'������*L���j�8�وO�c��� �ee���_��髦ڸ�ƨ:C(y�	����ё���sH B�Q��j+��j�+��j��6C��/\7��6��p����$����@B��S~�
`QZ���ҏꡉh�P��h� �XU���3��)v�Si��N�(h�T��i�C��VT��Db��G|)��.��r{�� ��7���w#ہL�]����_�K��B�"�r��F�������%"���G�����_��L�M��JQ�gÁ��+��uÊh}��NSkQΗ�sC!�fʘ��aY����n3�spV�To�P�a�?�)a��~R��Zb��JH#@��b��+k\�f��˭z�� <�c�>�/Qsҍ��D+��o�dN;B�[9`�w��P�j���6ӝ�>�H@��_���a��Ù��c�?
��|!D�\3@�XBΆ��5$`njޗ�WF _�
q&˚�kib8����g;a�.OkV��0��
"�k�۽�T�nd7!��8���O����D{p�`{4���k��x����^��]	g�r[��Vq��NDi����ޔ��jB#���/��qg k�䡖��51QN��Sw���̡&��n׊ȶ�3}d�I����;�ٽa��oS���p#�+t,q�c��L/�,�U��w�q��p�k0D��D^�"��c�'o�}��� �1�ٱ�{�ua�{�@���<�>�U��mX�D��t�+ɬ������f��\�S}IoqO0������Y����n�7�8<�e0,����r��[�9�x�\��2�rrq'噼֥�h�"��% }�G��z77��X~v�b��U:mn՞�D�R�u�}��g1�:��	�<�^�6�7d�O�ϸ���������<�%�9v�2�3��~\�-ϙ{=����$Z� �NN+�wp�xT��k��?2���~m�ă�v�̐3���9�U����	�ƹ4I?Ԣ��gq��9�;�rT�UBկۗl^���K}w�J��7 ޚ���4C�`�H�����ĉ�i2 �� Cu#bp���FK�ÕA__��ӛa[��t�tS �U�OJ2�l m��m/��1� 1sc�Z���;����e���X��m�����@h�r�	�iV�'�]摄(L'�a�U�J�Py�������ݺ�}X��i���1wZ/2��h��B
��m:/��ʝ��xq���r��\k({�}��ǭ�������6���=�U9[J���3��d�n@���}�f4���d�4,-�f扎�=�{��D���F#�W:�Zӱ+~+�V��F��5�����^��G�#��څ�5�v��Z�S���q�qJ���������ǕV���1)3��7��߷�:K������=B�kd����؎N�3ܶ(����if�������M�"^��ܠ��m���r��&�oW���O]D�%�\|�g�Hڷo�)|��bd���� ������uE�f�J�x���QwW�)p�Զ8���A�����)26s�~�~�3�L|�tC��0��{��b�L�!�U��0A��ն�"9��P���	��7���x��D��;�������eS�"�X�}�|�i������F��{5�a��]u�x^3"�s���X;��}��9O��	�#�P��ޚ�U�j<MA��Ȥ�D���\Ɲ�8����!j��(�%[\u�A��E��$��L֖<�^p��'TʅTT�,M����v���vyZo~qs��LV��I�]��D��s�`at�^�ݼX�S�R��6Es&�ے:2򌄍aݯ+�W��|��P �(��c�_��d4�=/���[6�$
����kR�Z@�fy.?���D�p��O�ԬA��Տ�u%��b�N����
��{aM؀��N;��-�?q�?��r6p2���P�}.����ОJ�1�Hh�Q2�s��K#ϽX�w7�Sx�j�ƞN/U�: y�/���k�}����Gh���mwwSk ��h:c���P~p�DFyX��L]����F��%uE�,��E56��?--�M~�]�q���8��*�E���[����dֿ���5�#?�G�ņ�c��)��p�c�1�
���[p��D�T�Cu��:7��ʪP~�t l�:,[�:��DJG��!G_FKr=2.jr�*8�PRZQ��U���%�wk��xwm�� ��n��OHy� ٚ�����OM.�}�F�)��uw��ؓ�г�J��_�Z�tf���W���d(�!h@�K��@��aa^W�l����S�9wg��4�Q���P3[g^�%V�5�
�{����R�k�㈒l��U�3����=����� �܇�A�O�a&����J�<ڔ0��ǳ ���!2l[d!�����F+Ry�-��p��"o�:�JP�\��������u1՛���� p�M�vN�>�P�:�2>�n�M9���3��`�Ǐ���ɭ6�r��B�Wsj�x)��#���v5m�D�	��Ep�<C���������ȡ�u4#nyF3��[�J��o�3MH��@���ۺ+,0�$���[�h�MW#o��_u�x֘:��B�(�(/%�A�P���}�*	<���`�Qz��Κ
.��5�����|V����"��9Y��N���C�����˱E!K���	h����u2�b���g�b}����^br	T�@�m8�����G�!� ����՚=�xO�VI��-���������aT�����Z��^_*��-���X.zab^��w*F0��C��Ǚ�S`=`L}����o��������wY^Ұs �����U>tdf���L�XQ,��A뀉Ӧ<�?r�����V�)���eŸbך�_���JU����Z\�|gR�雱
0���t�@J���#6�'O#�E!��7)���-C��4�r�5 ��A٧��<)��;%G1����y]9�X�1��La���i��I����P3M�@+�V@�X�1�Ae���uV���7~���j����C�K�V��J�+O�����v��P�ڻ<j��!/�ܩ�>��d����6G�E=T0z�=�(����}P�sm�z����MYV��T������"�Ք��Q�Qׯ|�������)6X9)���0&Z��"����3Q�{A /.-�jz:`�}�찲)CK2��Ѹ�aW*v{�L}�;�N.��'|�EU�3��g��.pC'_z.+��n�X[6?\�;Z���|,���y�̸�b�M�5�+�:�KT��'�&$/�0�?�\�?�-<�uL]I�t����-���C�K����B����/���:z�x�Ok�AX'll�5�j.I����@��q�b����yg3�N�ځ��S�G�NG�.޼���, z����e?�sKw״�Y����C^]�����t�1�r�>vZW��q>��j�����ԏ��3	p�ضH�ʯi�����s��Yk��X>ɲf�tDe��6�G�n����2u�O���v3|=��o�K��٠T�ōue��x�M��}f���2�e槹�G��#|����-���Ű����DN 
o��o� ��8�2S,���
�w������P���:Ώ�����)g�n�D�g E�%��b�J����˛fJ���nU}�1��Q�'��;�����a2N�#)܌�(a�ǖYd�n���YTd!�j|�dg"_����yE����ӌ�a�b��k`:�J�'<]&�$�_�,[�%���<���a��B���S���{"	گ�K܉eN�7�y@p9f�)�zxi�ڸz�����`gR�;������>���k���:@�0)s�����V~,�&�7�F�s�^�����Ŵ�3^~�~���)f�DcL�
/v�?�Xo�7��^���PSO�>e�&c�������/B<��.`XhL�bF/���AߝfL6"�M��FBc���gzJyS��e^+U�&mȗ�v��W0A�㲻-͎���Ls��\�|ګz���{y~�*���kݻ��Q�H(,˦K$��g�/������փG�j'\zE̐z�8��^�����<���	������jC�2ة&�;����@۴�4��a\�]Ҫ �~f�)�0�]�Ժ` l�!W��|� ���kzLHv}��rV�\��H���6�a8��V�k�Au��@#�s�l�F��dm��X�/�~O�V�F���e��wP��=4f���*�	Y�R ���	��D��t�o��K���'�;�c�X/,Vi�Y���Q1e�ՎHz=�a (mnVWQ���V0��B��i(�H��4\�m�>˝�N����'������k	���<����ӝ�/ec����F�+��V�_�&�X���?�_��UQ������ܤ��X>���U��H����S
o~�h �Pl��U�6�1�W�?��� �U3���)3�1��6��������%�R�^���3�KAF�"-5�I�
��?���ʠ/l^�w��Ud�H�T����B�q�SF�Q�8���D�)Q\9���p���-g1���dQԥ������L9�&u�*纖0lÓ'�e��s�6� �t��1�$�^&�gB|ơړ]��Q)CD�O�R)�	��M��d�6z�����9�`�*z7o5��~f��p1f8'��d������ٶ��2�{�~d��4I�� JWj��PX`��f��Ӱ���0B�o�Y]'�w\`�RK|w��>G���<^C]
"�7Y��� :��<w�ghHe�����^��>Ӷ����8�U�[J�S���5��Ҧ��	���I��0�@<Pޱ������o���Uò���h�^����D����ڨ�O����	,�e�[#�Wp�]�Y�K�/T69�}�q��7�5�_Qx���u}e:��h�0jtyJ���
%��I���o��oC��9j4�5��+�؂�ċ?�3ݚ٨�;ٌ��:�dQc^j�7��]ϴk���ׅ	�6�%T1�Erx$�~eТ8�ؑ�G	�	�.eZ9��琍D=��g/�E��l������_0���Je��u�:��RC�{��a�I,��lU�6ʍ�����/�gD$xM�n\�:���״���A�&ć���@�es��k�`��{'Dm�j��8���撇�d��)�L�v^����,�Y���O�g�������2�<�ԥV�IN�]|�̷�w܆���#~2]fp�헾�Z�WB��i�oj=5�N��Y���gʹ;�*�=��Ar��Y�A�-���Ӭ��uU�MB`���-:v�0�2AIջ�d�A0���(�J��pں5��� KK�~�>�"c�E�q��jA����9�Y�N-'RW�����
���x�B���p�;0���C����U#�lkBu�n]�'9y�~�˃pW��F"7�VE���w�1�9�A���zdZ����ՇpI��`_Ȏ 9F"4`O�|�*��0�#�h��Ɂ�*�����b^܁�w��cb(�,r3ׯzrn�|��PxP�'E�� ���\}�,EZCo�e�p�Kq�������xGTO����g!��̎��|�cmp<l�]���H�Q�`��lNH�IL�t�Q�yY���7��Mq��U�+%�B2�X���� �R� ��~Q5I9chͳ0�i���Z����ȝ��/�Ԟ�k�t�A�FP�>��7�U��V�p�Z�����)M�%�}�/�r�h[��l��!�f7�z3k���R�ְ��<��>� Hab�ދ�C*�'�tK��r}���Y!��K�c6�(6�hj�`&�K��H%k���'�7�2^�r�j4�'�����k�O\�Ί��L�����9"���|��Ī˟O�b��#�Ue�R��g#�մ��6��k��ѝ��2�K�;a�N�D��4���� �\Fyi�!��d ����Σ�p���&D�jYxZj"�vW?lm娊6���]��b�^偉�jګ�,I����-*!������ ���%�B���1�'
�5Yٽ�k){[BS�� �q�b��j2?{B�4����r1�������s����Oq�PH�;JRW+�v�ȇ+t�\�	��̥hb1�*DABn�,� %\|&��Cd��b����ݣ(aq��"*]����J$^�$weR�9B�#�Ƚ~A�=PxHd_D���|)t@���� ~��l�7��7��."����E�
|S>�5��&M���"&[�Pٓ�>�}������x�n~��Ǵ��-\�n��ҡ~���^>�����o�/VCHѹj����0>@�ɗe�/�T��I�����yBf�d��ޤo��Tc�=6��b�)p���(��x�d��+\�+���/�Nnް�17�#A�DVJ��6��v4���h��z�ctM��ܒ���@��S�p�8�޺�r@o�_�E���ڌ�l��FmT�ȎgM�]��!�ݛз�`^|���~�����f��3�߇�c�}ثm�{1�[U��`��H�b~�$�C�r��IqG1l��	CU¨�x����ɡ������652�:'�|R{�V�^���Z�Mz�ݦ����[����5����N��#�l<=@���u���̆�_�5�x��Wuȳ/�-�(㸕���)�A>�N"�O�����'�T� �͝`FpZx����n븱,o�m{��t��B¢Q"����<+�z t�]�9Iqq���^��O�g��J�2�|�D�O���ۚB�3}�b#�
<��z�6��!�|��l�IaJ�T=R� ���*��X��Hɒ�p��r� 6z��]��=�\Zi�"�r;����V��ҙӣ���Z�:��O�L�7:xv�	)>O:�O;� N�F��F��d7�/MI��hOw�>�QH�M�ʬѺQ��_����8؜5W�{���E����<�P�(U1짯U����L�a!�z�\If4��V
||��\�UnM��k;m�{�h�f#h0e��a��
X\����]Cm�n;S5z���P G)E�������h+lh0��g�!;��.� �(c��<]X�Q���2�a��(̺-M. �li��"� ���Rt���		ٷ{)�B7c�0G��=)�My]{7B];T{����&�Tk��Mu�b�S(s�������]��3pʫ5�B0X���w����~)=G8���r��C�T�{�۱�*^�zln|#�4�%��.|?F2�\W�Lj]���5��9�V��W��Z�v�P��Ύ�:�A�5��bs\QF"J����"�c���m��Ը��i����淅L)�)�윋=@N�(�������60�X��oG����q-�R,{�d `}C�ٶy���"�J-����H��$�9V��k�Dw@���na�F�Pr��V{hW<���(%��B�`�:]{����UP\^��8(D��4W!	�?��^�f���Pd�m����<�$v�qC�hr���>��V��k �ƣ����z��n���~|�ŏ�x�"���p� 	�f���P'�b.�f15 ����a�l�?<���u�gz�n����Z���E!��l� ��$K��lf�0s�B���r���?	����
< ��[o�N�0�����~㓞G� �0���e��ب9a��Z��~w�5�~��`9T�7�i"mv�!�#�UsF�l��$08�^��dy��H�a��K��F]�� f�8�#Y���Y���r()�AhY2�E�$hX�6�|e\�x��zC#���%�;23W�6�8�x^w�k�$V�oJV5|R�C�+D���;8�m�o���0/��XƮV\�B�`͠���m�*�\���{��޺�+��:��~�Τ��|�-�=IY�"߅��k��/E̦V,w�}�M8좜蕏rbv�3wiw���dcn�G�	b��	�!}?�&�F<�����nX�7�P���d4���
����)�]�%�te�m������_䑽8���tW�梧,u]�����!V{w/�R�BRk�s���4��NY;��q�4#�<G�k�pE��me�p�K���eCg�s���"Ҕ�_�Xc|��]\��z����bL�geϛ����G�������'&��r�l��XH�h?p	=�E�����⸉͘�1lb�0�5�Ț���\��`&� �d�4�E$%�+��] &����:T�qq�j��b�F5��5�cH�9DXJ�o\�C9����88b�_3W5j���0����'��Z,����t��e�r���w��&�ct"����r����
C7f����k%�-�A��^*�{�y��D�2Af��ә��`c��#� ƙU\��������g�T;.gJ���A��MjZ�Dm�U2���(�%.>0@��P� ���^��e�Wk7T�k��sTL��~Ai
�Z���y"�Tb>�7E�D���V�`�c(�&�\����F8t�V���f]u!�@�8A�s��dһ[��L�4�H>f��!Ӷ	�@��R�	�(T��4!2�wc8;� "`���I�C����5��3��G`Gb������>�	~�����
tV�i_}�\'�8��Q�z�'�"��/	Z�cް�X��!*)mou8i����@��R�M�G�tna«W�n���t��~`�%��4��h�&k��[�SG3��wѩ]N�3�1r�F�5G������o��R����g���'�q��?�)�����rg�sJ�[��(<�J�؟U� �Tv�G���r�/V���T��os�������}:����h��G\&C!?��;J�[#�f�:��X9	�F��YU�i�f0�H�(��aa���|��4��Sլ��l��/�u%$;�y�Jl��+6���p�,x�#~Uע�g	�\􋵈�5x��xYX眼L-27i)���� ����������t��؍|��0�j6�r?��F�d��W
�`��,:�%��y`�f&��94.Lڣr��6�[�bK�}�)�(mG���0��&��h�0'��:�+�r!��Wcثԕ��*����5��q�[�G��V���8go��P'+�ݕ�G�>ݰ��W���I���	���o�~2}���|�J"ƃE����v�
�eiܧ��"�9�ж�QIW5>iWe�݄a����=E���>�"�Ȇ[vl�ᤛ��P�����Հ���&�	�ptt!p���`Ն��p%����t5K��X��HYW ��{)���ҵ�Y�e�Li/r��CW��$��r
F�)	��v��(b5r*����7�����?R�K�M��4Ls����JK��]�孡"R`6
X'II�F��	���w=;����1*Ϥn�\&�m�A���1�*�Ʊͨ6ƒlt�>/�G��i�Ri\�.P��"��;O��<ȩ8
�%����ȁ@���D�'��/̺�s�o���6[��M>���S��B�(Q�uL!�'[������3?��&7�.�_��}ɔ�;WB���v�t��Unut���pg�T$d���y�������"^�l���g���	��z��P����-�<o9�v�f�syQ��{�}~��뇋�U?	[�"�"d�S ڡ�FB����|�I��K��rȿQM��ę���!n�j�\�Po�m!"��wLb�����L ��p#kB�:xd�Yl۶
�]�?)�2]4m��y��\�u����Q���^�,��k�I�@Py�C���Q�	+!9�WĄ*�*6�l���f
Y�� l�Q��}�^�ᮩx���!7k>��9�/o�C8���9	ӃXBVR慂�4R��Y������(�f��'�+<���x0���*���}������vz�UtTN��᣼rwZ'RQ�E*�z~�z��`�ğ���V��-u|��,��}H��@l#�7d�&SvN�G�����~h��p~7�8F0���E&��9@:�Z��K��aLO k��,n�/D��.��G)to�,�;C��2�_���k��.��%s�DIg�p�ɛY��:�!�����G�݄m%aʂP�7��;B*���M�PR@�߽DK��,ϼ�J�\Z�#-��cnH����oG4�А:��/������	��F�m��qpAʯ���<��O+��v`!s�n�NF6����b�I�ia�>�D��aO�o!�4iY���C��O�$l;��	���D����4�҅U'���� �\M�k�d\k��`;!.r����N�&��c��D���iA�)�A�I]���Ep����Qj2Ye���M�9%i"Xfb�
; �o������n!݈��@w�m�ɧL~_��,�WE�,� j���C��K�	�_��i��Tw�!�Nso�c/ti>�qCϮ��+G4=���(�����?�M�ʚ�I��DZE�qC"�:��$�Z9�t{Tr��U8�ϛ+���`?l��աE)V�G�9VI��ms���oפ�{;��E��P��� P�C
z��.����8]��ǹTj����U����5_z���_@�,�Űs�a7��h���E��l2��2�L�o~8���T����c���Z\�uع����ʯHz.��|���H�Gq����'�a��큝KHEt��`�'?ڡ�����T�Q@�s$ ��%b��5#�ߏ��0ϯ��P}���.����Y �.*$�(]ܤ2=.�K����&�A�y��i6�w��Sbf7�w(17����)P��\Y���!��pY|����۶!�z��1��s���jlx�J��_�1�A��ے�$p�����r��)BZ��Khb�X��E��Z�=��Jx�l���5v��0@H��g�1/8h����Kb�3����J�`\O˒�P
�;���bOOx��9	����.��$��
�J-�9�w��b�6kO���A��b<�G�P�ZFe��|�yˀd� �^|�T4��Q�����B�;I��Ĕ��.ƈ$MsX0OGvl=���*g-c�g�Q�Do�o�e�d�ʓ�*n��5D�y<���������jV޶���ԏg��0N���8�����rX��GD��CÃDo=�']�P�]	%<�Xq{  �q��	����БM�s��PE�@(���s��p��R��M�~���	��p��L��fq�\�bPO�����7N�1� jV�*�����˧�Pr�Q����H�ԕ�i��G�EL�B��U�t<�ӥ)u*�z�yt��Ff�2h��'qGA4�9W3Js$��I�$�n�થ�!��p�a��̕+�HȌR�o�ÑH��8Ya�.���&���u&m�^ +O̗̅�!��ײ����*�S"l�m,�����id���J~�4L�iy�aF|K��ڸ���HaѥIM~T�w�%4�2�$��+>(��-[K��w���YG��	d:EҢC��ƌ��\��; *���
^�WUKfA$�|l\	�r�O#�!�=͵��xx*ͨk]�
Ѐ�jV��� thB��أ$�Ǜ�oH,2_�m�a6���1/��7+#�6�/wyˋ��{w���X���	%��**8O��S�K%g���f�ɏ{��߫�Y����:ɼ9��
����+�fZbF'��&��@��%�f_�Wf���2�%�=��u*�8FᏟ��T��aW9Kl\H����.=}2!���ӟ޶a�cp�TG�a[���'-*�[jjn�P��W9X	�����β���VyI�͠+�.����'�
!K(.�;�-�p��*ea�����m�2���`�qY�ڔhR�B�o��@��K���LVw�;M77NP_P}�^��٫����0�L�w���[z$�~p7 铗gxOU�0��E�w#;ʻ��>�Sk$����
��D)|�~yV�m4����4��	j�0l
c��V�I��'RМ�F �^��aY���||>��WY�Q��1W�і�u��a��O�W�M������(����#$
���;�w+%2)��ޢ�M�7O@�5�VQiR�J���23�;ベ����s�D��݋����Қ�2�==�� �G�l��9\䓀{���Vd�%�/�"��&�� �'Ӕ(nW��!ҋ[Ʉ����g�Ϳ:��L�Հ�r-�ŁL�0T���x21��	�D=�	�x�Pc�B*Q��{8*�����>�z���[Á������'��eT�u��#�|Ro��,�6�"P@�!FYl�s�c̕"Q�b���Ď�DS㸣�y^ߌ�����T�=�k��\;nMt�@ewl�Y׋|�2hP6��q�?�^�3� �2"*�t(���/\�켵\��r_.�=�6�G�$�;��c9��v0�䂁�C̻7�����^�B���5kOJꒈ���aZpH<��AS8z� ��\,H/�f��@�+1b�t����q���������؝4J�k�I�CjlK��D�d��ʅ�?��� H��a\��.���^�I�@{�gn�u���a2II��c����9G^<�@O��\\�P-��`[����Z	���8� ���ʮ������A��蚛�C��'��SU�dGU� E��b��Ы��hbHUL��9�txVV���}t}wqljyg6���z�"�.�z��g�\n��*����4���e/o�������K��^�,�	춼�l�c�M�峟��E���)�5A��>���(p~V���r�`o�u#���*ei49�TjPA���z�6('UEc'���.� �._d�M��͹񄋁�ɆW��M�uf�u5�S�{��1���?	�j{�͓[-����/o�5�O�<˃�[�oE���@���Z�7OSi��YI]�;J�̎W'�(�Y���6���=��#Q5EQ�J�wj�
�m]V����/�=#���c�0%��A鲍8¿l�$5 �\� ������Ҍ*�=e�� n�M�"��\ޔ5D2������b:x*�T�l��@6>2|���}հ+Ng�0��	�:yBJ�No��q��nK���B�R7/��hheH����G�կi��L��SE���5I�����Գ�W�礷0�L.a/� [� �Ǧ~9Fo�$���C{�ԛ�|J.r72 ��tp[�?
2���հXd���*�fQt�Wf�"r�=x�+K�S.Q� ;yږ3���>2.!�Ȣ�cJ��{�_��U%9��k ��$����8�Q��OFό쮟c'�S2����R���@NH��!۝\���g}\����/�M�G+����~ѻ��!AI)	��?&3U�#�;��f��^���=�n��S���TF9���\=�&U�!F�)󾒞���Q� �3�j(<��M�����Hm�Ec���b�<��g_�M�@�]�]�"*\���P��}��Q�7�;T�%��q��R{a�ؠ����Z˫0��~��SPX�4�něKWϩ��O����)��X�I>4�Ub��hˋ6E��R���P�p����u�13e�|B?$���LsF.*7s�{���\:��I-��N���ē��4���6��p��N�Q�²�����(=��Z�L*�o�s��J|���[��lX<��ؤz�d�e@2T�A��Azv[4���y����p_Oڶ��ƒ����4b�s�|�(7�\g�]M�a�x(T��V�S������T#����U4-�C�����各�&�v:3��=�T+��Y�t��A�!8�L�t%��(�s�7�`OUc�^�L��R5A)iRL[��I�8��'�m2V��!�]�e���m����}7&~�(�V�G9jb~gP�7�Dr
�,�mS�3щ���7o��&T-������hgYk�OӞ���e3�r���t�&�B^�|����0�bj��587zN.|�*������X��;��9$���C�ꨰ�)p;��WU(4�#5e�3*�~�:�Y�5����\{Vi�n�̻�honSK�W8�ofjn`g�6c�\���#�0M�(�*>�('�<��aL�L��Mʨ8k��"�wK�?R�:.�e�pao�x�Sk�u�6�-\0	�q����Љ V�)�|�(S&Q}�)������H��d����(�(����s�H�?��@���.�n٢�&O+�G{}���6��������V�b�5\��
����JY�h��������|I]z4�����Gw�8�a0Z��W�������ۊ�T;��"\)ۄ��DM{�*�����<�v<��(�Z�T��6:�E�he 0,r�?�B�r��j���p/P�Ni���������QV<n�[�h?U.�.�D2���<��e����/##Е4�yV2b8m��/;	@�x��?)��^ɃG�aI�L�$�	d�z�rx�#�{1�<=�⩡팊$���"�pr=@�7ۛ �њұۜOA>Zj}��eY�M)u^6b�>�FAY�w$0���VE%Y�kB�OQ���X�yD5'�|��]RRCh=��[i�q�DEZ*FO��]�,�������j�鏯.�:#)�v����"���᪎-2~q_��V����ZހL��Aij��䶅��T��S_��#�%� z�w>I����o�`[x�=�e\�?oj������+�m����4�VO��u��G'�X���r�!�K��;��I�ɝ��^*ްM]����L�L-�Dw�(�4��q&ε��3�^���GAP�6��y��c�}Bu��ݘ�;3;�[v�QD�)J����
�Nל�iЃ7]���i(`����9�J��uht�5`��5
���n��tR� UY���Y�|h �Y�PW� 6��f��l�uY��{��{��b�=�$d����~�0E�|)��]|�tuMۼ���U��-�e1�ת3oAI!E�R����X	��0R}�6ߋ����W��ņ���xI��z�ƛ�L)���S�f�`��9�G����	���p�ö��F����7��ѻr�P1O��(�s�&����(r�"�O�\��5�4����thZY�&%�l���nF�Wf]�����Y�l*wW�������5�W[�0y��$�u�.����:>Г�n�������)t�D��W�1E#��?��� ���Uȸ��[��H
>J��RhW��iX�4����Ԩ�aƄ{K��.s/�ο�r������h`���pd('�\��؈�n	&]rI?�Xdj��s���a�����H~�s%; S(&��6�_'���?f�.��X_[�����=/}�e�����j�D���ˋ�1VY&�u�`��T���==��C�7��?������$#D��W��WNI����q=p�ħP@�/C������ :/q���&��Í-�����_ʻ���2i5��>ZҪ��VK
�P3��	Ƞr�8�j�F��l�ɍ}����i@4�('��Xre>!�u�ؔV~Px ٳ����(�������B)��h���=��������r;���,9��آ#Ɣ4&�:kԏ����!��Q�n���j��K���74p�%~e�R!��0ZO<Y\����E�%Q��/�� �1:�����@��i�-�u,[���g[��9kA#�����%
��r�eJ�����2��?�uJ�+m����������MԬ�A��vQ��^���g��	��)v����=[L��>`�\?yam�zo�>b*#����f1���D��q�R'� U�������L��cI��a_� �v��&f�Н@��4=?��&Y�� 1�L�Ϊ���ѵ���Ŵw�N��}iE��n����÷��9y�rW�O�oK�Re��幎eh��K�� %yxA�'I��H�Kr��\g݀�ud�Y����$�l��g�6��$�j�j�����Q���kq���s_OD]:���?h���gY������@?�}���� Nx��A���s���D�)i����m�F�3�b���~�!*Th���̞K�6)��Ȃ@P_��'V ��3�H�ѷ�	+L�oS6�Y̗t�x�~7k�ǟLM�6�A�0�Z��Ζ�0�j>��Pd�Fa8P+�g�!������X�n�`F�+�hw]�������d�/G�U�6L!*�.��#/�[�0��(Y��T5'�,�N��˴ϠѬ�<����٥���o��TR�r�󸛹��A�e�o�ᕈ�BF M���N#�D��Dh��h,��՘�NQ�X(eT�{7d�́о(s��w�J�-���L�¹�&��q�lu�)���WG6�t�uCA��^�B0���I�#�����-+:X'��`�}�A�}�z/)Q�V}������S?�X�:nYV�)���J�Ӛ��H����'Xm����ǵ&����O�$J�DU"�]��k�;�4��H�V�7xdH�E~��h��N�3�+G�Z����j�re(��'$��<Ӥ͙��ƺ��85S̸~Ь:��z��w1��t����B���G��U	�F����W �RwYM^4n+��jY`���j���&��Hݿ��-��'PmS��+�?��)�Wm�MJ6�Ԭ���
%7.(����*u��TO�2��x*�9(p�c����`j��$��'�&�����1#����kdh�*�j=
C� �M�jC��!9�ˋ4n��ѽ{�c�r����7:-d��l�p��=f1,h�wȩp��͐l�+���GL�D(ῖG~�j�������ˮQݩ��_�SO9M�ãE�Q�qK�����5.�%������`\/����U�:�c�:�r܋	&'K�B.̂��,uN'�Ѐ]����3���Q���k0ꪀk1ߔӈ,��7��ԺbI� ܙV�0�h��V��1��~
����<�׉����A*u�$6G���/q%raʭ% >��9���j�%c94�b�;�"���YR�U��}���mD"@�g���!�{e{v�P�o�H����b��
�]��>4�p�cUuA�FMhY��g�IU�ZOE��=K�'�z�%KC��i_K��q�L���ww��{A�'Qz��DU�&�Eb�$9^+��2��PfE��a����C�1�4W*��.�d�_����pZ3whk5��bN�����H���b��iZ	�U!��"p�9/=f��T�`
6^PA�,=TYJ}�A�E�z�N�A �eU�y�T�L��K�\u�KEk�aH���(�(�  �,��@_\9���^�"�Xw���� ^�|�j�3#�t�Q
��Eۻp��Ä6���pc$u�� |��w5^�5���>��LLv��BQ{��^C���)�\�w_����H{������h K��/�*��a��*4T�$���ؠa�wݢ&�ӻ#�O����@b����g#2�
����Jӣ�Q��n=��f�\���v�㞓=SW9p�� ��ذ����$�1�$Y��ր�k�1�C���ݥ'�S帧bR"MO:��ί�/1��F�A��̵g�_���.�����`��k��x|K	�m�L�n�d�䐒���m���V\��4�L�~�DM"})Ӹ-c���8�u��.�ہ�H�E�2/`�w�h�O
�THY&>Q��� #�rf�U)Ӓ�[����B��twe��FF�ڌ��3(���2m4>mAC��$�kr�V�:�}��|	{���R`w�O�ʔ��`YDD-&%Q�̘0��( �HQ�I<B�k�q��F�p%
���KL�Ğsղ��z5e�} �a������\�g��x�oq~xQ�1�>5��'��\16�V@,7O4ex�8$�sǙ��Q�h�EFQs�P
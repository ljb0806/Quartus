-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zN5yP7XGFJTDFXD6HqNlCY9yCuQwBItFV/ibLzSZx5V0eEG717kHUO+gWoqXnVxvz8Vuuwl1B0ti
r0zt+9mKiNKexI+RusaLrrjCwXNnKorLyuz4p/W7Qob+1JU7n4TjFue9ubVOr8cH/D4sj0QK5z4x
bwpNCh3jYMDIaSSI0Y0v57et2J60eKjVV6HkYAisqxBigFu4eiQeMzCd+GyMtcAlln80dLWUobHd
BSqTGtBxGc50lq4x9f2GieZZHEZQwsnwk+pYX58n7dGEpC/hkUDXzcjhsluvCsYwwPjYTQFesVuy
AtmMYf2dojjw+sxILxKO7kvctqyhLfFOywUBUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114400)
`protect data_block
0wPTxFmc7gSzileIueTdfxFm8AXieR6OsbEM6vuTupRYz21g8Hp9Xa5aNUFYoIFxeCKsb1GB1ZE1
xiGkTm9B9TcwrCCKDJ9ZRpHhZ2lr2ruzPKrIQeVE9uzySitac02UZxYNUw0bKcWa1MvUM/dQnF/U
UmMJsr+ZL4DQHOIHHqfnsDVVr5F+ef3rdzlT7Jc7+3KDZaunlCObDRJ1uV6+lsRLPTILHCeDT2K0
K+rIId6QXD4LOt4hqun/RiAfglyyS8WjTVbL7JRRfvPWcIlxOAsm/b/Nn1csOkeLkxtbGOCWfO+H
NDb72NyuvDE5m/rDYjp4b23t8F5HzjWJrGeG4xwfevgU38psjmwgANn95pCiAM762fk6cAhyC8wB
OT61lC176tbq959IZ7KNqpT7fPz8vnaTIRYp1jAsR8pkr/iBTbPeiaO8oPl7Up8EjiP0ISAsCai8
5tz5MgUOXf5+JAH4kqe+7B1QM1siBwDvzET1n7LbEkqnRTxKLu1rmbba/CxPZBGamcNbpqSzWVkM
KMmyoFTtnD6G14LrhqhWW+U+lno18DOsLYoR/4L96ADXtlmcyh4p/2undzB6XYSuZ1wqB+wgN/VG
OlCiAyE8pCzunJXVxdsUwANL9La8P5OAF3DMbn628m5KxbmhxP+iF429+imklcUVmcekNK9QVrqi
7amd3YqHu+7IkbQVV5TBVovIqphfm6qc9v5/qPSuQkcY/dEataA/YhXuwzaZ1K/a61qfJCVcI3MZ
Kn1o89FcDVPZm0hz5mGlQ/6rNIPxr1kbOddGsiUEnhQBjJQStch00CZQCCjHcYi/88piKryTDGko
JzqgoTDal4m7oa8zTfIQRyfcCHTy/5EhFq8y/4ajBwhOipuE6N8FS30emqfbDmig6xt1Z8+MOTBa
yLY/A5SALnwBkWWXCeWjqe21qhi/9VVi1jIfca17/qSkPIToC3LQ0SRSmNZtONy/8tHatFFhCJrM
pt8gMvN9DatMDIv/H+VE6Age988IFAoHMmgyHnZvEeqbpJt49gn1dCJLncQcEC+yJbFimOjjHylN
cf+mDSe5lkzMs9t9hr0ldIyTcyebJJY9pUuD93HNA+y5+uN7zY30nNWrLma2vA4GkU9cn9k7hILo
zIFevle5SFg6L6K4HzbjPZYhjECaChQ1DBzkXDe0a+0wms8RJxc+gKjMhb6VNUf9XWuKlfxV3x6k
68Kp7b0jXXCVwg8dIJzu3vBoxw1gqKAjkDvJFFLLltG77XeUNoONB2iaSIg/zmVXVHFymKi2gwe5
Fj6Gvkr0z8oHz5fuWX7tq0Q05s1l0ZEtKQSrT8HDRhpqfacQchmirXjkMX8CfYKhIJUHpesUvtq/
amZD19rwtiz8/aCWrLydCeZZA8uQJnfgBciRHN9vJDgxc4wsHzUxruI6/WUBoKiJgxzqbdDuzF3R
XUrXv21/TaP8U+cuTcPixYi1OhKa9nAGXx3ZK+Emdry5aka+B5baJHvB6hqZVyVZo/Q9VzwCmlgw
LJYYV3T8nYGY+4Y31tDFukR1Xg7a/Ug3GXfz+zDCr1Ee0Rdt4HPMROGBcBpo0m8wd8ovbdeWrGNi
XQsxZXXkuQ2Hruq7KJLeiB/zLJpA9941PU/T1lXlYl+0XIUaN7elO1NojLOCR8/WFVIVRQG2As2g
59pfiuJTlzEEkxLw56JdJuiu9i4wpi9rHEetSebzj8Kowp/05E0gUWXN1zxX7W7iLn9/ViHbDk1C
hP9Wqw6IuUMIr5LdiD3e3NXpc1qebkvl1Z6wK3z2+WeYqOA3feJ54SDtAWLm7dis9cJK+YDyrqGd
tu6sm1KJS+b0U6aZvTMoZeTdUSrdNfzSNK35JFeZZ1FzPL61aGJR6cN4j7iuWJo194Di2EI/KpeY
V9R3hv766POi35Lx5+8deX9Jmin5S9gxH7GB5DSN3lcv+TgQZ9AFrfzWB8sdCgd8C7DWlvwWmyet
+jO+3dYqD+oVF0ay1DXJ/4EXZDc26MPIUys6uTXEaGsRYRdHrvsxgEzhDxfrRXzjIZ20iNqyi0c4
PZorSeByc2kpPSmejsh0UeA+tzf0F5rWqnbOw0mslOw2ZP6HhT5fNXtqH1KbTs8jVUzS8hmc912H
7n9Kq5qqz6rx9T9dW2F1ginWKH5Mxn8XrTIBXyfjpfJZX9cyKmk3rN2ZTqe3SZN6S2aI2ZBQ+8IL
LN7oDFO/UvjDu62qS/vILbEcBoOW+SWDKNXgN/XfcdQ84nicvg4vSww4YEosYt2zTqru4OVaxAEg
1rtwsrIY5L4Dp7cSDAxRhJCqUXzKV4ZBDLe6r13EXkdzZA0lK0Pw/MuU+DZo8wovyl2jzNOa4AH2
R/gzGb5zBKQnGaxskoCPl4iRHnpuM564SLq32bc7sAEgNXePr520k5vWTkqpoj2njOER2BSCJ/5V
EKEh5tTXS3eo6ZZ51vERS9xQMOK+6rNFUaCLLLNcFEdR/+FxiDW/QgaG196jPzfOBYN6k7joQFL1
OmYL9KIIF+trZZLtgHMHczdiCXtgpwjDTc9LNFyn4GPqV/lPVsyTRrg+zElFPsIShzwrpcrXrJH6
sjHDcdY8KmmtjB+cY89B+eqEIBooQgbX4JCkuBduMpJhohopXgZeDIR5AsgtTSPCjZgb7L3gpT+x
wvxhH3ezFC2kquY5K4MPMrfGftHNnrttx9Uj9CAyB1p+Ln0V8Q47ooEBUUqWvWNO2wjfX27J7BDp
ozwnuTr0mDcKUwYnBbvwLUhYh2zjbStbHH1iXygAHyYtGnu9lpelHq4ExSeaHcsWnh7HrWPAEjU5
GvQzy2tFwglJD+y9RRi8I1V3MMt4lr2UI4+IDkeal9c/1XhYmv/jzn7l0xMRTvV9MS0hUh2uwEZZ
zUZ4+U+l25RvHVAufdjj1BWWoJaZoicpUspysRF9/FVos1GCL1z8Tcf++0VvK6bVKCsocGbgjD+8
r8guOVCqufdmaQdzPClhzEQIkq47xVCpSIzPI8X2hN0aoghiXAp5V/nNTW/LzR/urhNi4Oo/WDSp
rzKFWhe5cWVGtEGk8Mn+RivJR0pp+HAHvoTxHMVJZfBIKLZD02IyMYS1LYdccWd5qLzG5Ay6lWYD
U3MvdaMAiQqqUv7uxTkOHOkUruMk1xx6RHN9uCmf11hWRWGf8wksWRCkkaaeiXhQzjq3bbeHvxnq
0aFKydg9oiXll3zdNiCYfvmj8qy9SaVTUqR9xu45Gn9U6CYutowNRKfMDOauZrIz9dJomz1dDyX2
NscFH5vMtSNnEF4soqI2tkcdG1xr7hbyK4WsafARJT8lZ4AXKIUkFoGATffKnTz+jel4c1z5yhjU
vvKbZfjnGr8c5hSerRMSgCQEs0M621qgS75/kjEHGMQbCsQLvQBXChUn+OiEVAIfqaIVRlAImb7E
0Cjlh29egfddOH2yD/78BD2+NUFdvJsNbBZdLdU9D5Z/nF0h4mjwvtqQ19Qpd6ZVeo+6rMZDv5tj
bNZdRzU8uIKc/J4BnkH7SeKn4twuSpe662LNrwp1lPRAXRazUr7JV/qdEU1ALdN7zPtGEuMOY5K2
2Slez39jda/MvPodTlFU3PQ02vSVpDIMJcGbYx1uUeGmq8591eK+TpAWQ3vC0Pokjxtp+GsrcPLw
+gemWI9uL+IQ5YORmOGL5PQ4lbmdG3nZGofKUtH44qbuvYy5m1RvTsN3gplyW+/yNgg28fLTeFMR
9QkZ3Tn0DLrdafrCcnJewvil4kx+4EtbMgX1EEtMTiLqIYaPnhh2fYQT1aMgwylfGBCtlbMoQG8G
mEi5CQqbaqfRzc32QvYE1LE+o//IqYfzQjDGe9lLOPp0PnicKOx9Ob6PSF1AiEIivilUB/VCKlMq
//AxSFkhJBcAAAwZaN5oHH0urjsmSl+NQaITDmwMgriGUUfp9xiTClKUasr0L+aWpTuFG012TuVB
V0MYDx4Xwhy8OxGQ2tZyXRpJx4eyA1SoNxQsY7Fay+F5DoxmDr9lnBMhfE6jz/8wxu/HkIxug92O
grrtYscIqc+QNibp2NyE6nd07XQ0WxDv9pJcI7ZZkb2t0YmCD9wQbhhSI51ADuYEE9AOJvejQG+M
/FrKCxoLeuulwpSP1aFWC+DJwnKggLwr3XEW+O6rswIkaK0TeSUiLlYxqHB0bGtvI+qpoLqDjouR
kaeFON7tMmARq6BKIq7iYfLn2AlGVCQs0PyyRjLZvoEe1fCK5KGimOrYe5yXrNtcvIj3cM6gjfx3
DqXxrckCJT3wNR9uAjxL0xQQL60+Dt15nzxz5jIdPY6Pk4rvXTQLWmlWUY2HgM9YkvQwX9eRZ9Y9
1Za8lpdr4BMYhTXPUeT9/TWo0vHWFVq2VVPyhL69Lves3adHjevqRPspljYbjyUK5o+y/jc2OEWz
/X6kgGTG6c37bSABsnYABaRI25vEB1wikRIbyzPFmQ9BAQypz1zcVomhfTnbOF2xpceTou7L4Bp9
Z1+sh6h1AdEXvj8fOR9Ao5JGB0izUHVefWbqDnGnfasydz1RrMILALO6FtS8AhN1Ol3XxEYpsXDQ
whbO3D0TLl/IspoDXr4cj2MOWEgtH5xs4q5apa0zRlht3ScJNgzM46+UMQXGlANlASxFV+neazho
EFV7mrcNn6DxrDX8gbgkMo+Djkv14Cl5syVs2ghjDxZEdqf8Bi4a1pycd5aALX84N2WIBVM4wxEJ
nogt/j8ooDswe9AUv/IsP3wmKFWFoHrbYr2OEJQARz/qss5KZn2NU9gC3UXT5eTYXtNs2QMg8oNv
94bfrvEWu7DY4EX6niBzWFODZY1ImSMkWEAcbY8Y4kKwBI1ID6v30DP3sS+Oe6y0+hXsazeao+kF
GzQDO6DYZMZS22eNNOExLyRqdIl4RDi10zvJ1bAU5Zfg9nRIhSxm60GvPwgJHmEZWt5vlGD3RnRo
4eJTcxgmEF9KS8am/4bv8tV77rwV5icGqbwMMmVZroNVHSryBTsfn5rx5hSN4GaqUku5h/3lG2aI
jN/khgirSbbVCTY7PHX8Po7okWo9N07Jcs+he5BTA3vnl2PrurFMQRqih7c9pL8NS4EEZISBM0ew
KkOdrMMjJFMgndhqm0IZ/hBRPHqwA51ArQN2R2PiJ0m5UwKg4kRoNC/IIJpJEnR8xuTCAyQHBV7E
L9SsKtBQioFV+64i33+kJA8yyeZUdvAdjNcpeiNzFIbia5FZZ8PR5bB17g1SSwbzidtdkmJAY1v7
aOwFtSVYNg9qbY5xIX4mRhyde9xrn4m0aMwom35S+s5Zr9vwnkO4O2DjKj066xRpN/h6VF1lgWAC
Ka82LeaPSOo4GZSDzwYJaSR+P5rPy+VdJ651QK79lTUAwwXOWXqZKOFQ1WKJaDZZ/glu8tG0ymB7
5XJJIXKzJ1/CyGHskIe/SerL4Lzvc8TmEmhKCp3N8y16fTvpo8EKMSFJ+pP72y8Pgj3ifoBDY3+N
vUbQNhUUnN7fBJPTMSiHz0qkUPij97zSDRZC9OidTAxXPE+PFTeeF/Josp/ke8/j5LsAWkLrciPq
Ds8AQPJUgBWdtsLI0RlVqB4H6NLpi/iOu1XAF1hQukTIjpfXu+PCvK7y4bm2X095SmpdIzJ2m3ZD
QsOnw1W4fPr59Q7XJfiOS8+lCKozfUFQ1Xacy3DSLgC07wsM3FwjSFt5cilTjno2/xVssdMhDjiu
tYlN67Jcl6ual8H+z6EvVTxyHmVs1BC1ftar2sH4ZoBRy6dF6O+lXUN54EOCYK/raON/z+KW33Jw
ROyAKH63Ow3swuJUlt7GBQeKP7uauP3yMXo/pfQUXiRO0hpzc2rPfqMy9VxCdyjehvNhAOIiKjtw
xY78bmhuUeC4RDY7D8QgWhBhvpWjAEhsVsVFWHspUJxD6zEwjsfiun9OCrtEFVwo2CZx4x1849Sc
X7/EXricbzT6LjlormaKMJDy4KRkQF3dFBom98jBHEPV+2017QPKdLElL9SIaGkF6R5q3cUqn7dl
nELoMANlQOzD7nCFDuXk3uJD767f2/TeUhuuz4+V8t8hPXJAfExTMR0WEEkWHAHFH0QwG/zGgGPT
Vv54pEnNrZsCU6fVEl6XK44oHo0y9zR9x6UJASwPs4dE1VY+rxIYNk9Bpoi1nSs3ZLieTmNtLa6n
XF3Tve3FD+UxPva3mlkUsyM9OzA6aefG/SjPOhFOj6j7dVW9yV1aavgRjO6CuLEK69cXZE+mtIPz
TNqigpSbNHoK+ml1ulJOgrgtTFKYDM9iIHSsW8Yz3DZCz/Wctg9oJ3UXhnPxHIwe5pzPhNl6nUSA
zDU67qvGT90VYQJY79zY0m85Audbx4sMUxV80pwD+rgSzEmCa4+HSGqxkd37BIO073hIbNZG70Wp
KQ6pzN6k+EbMiIsu0OAAyRNL7vpUwLKMJx8N2rLv3dLw7yYnub+y6TW6Hv7N5mmX8lD8glfv5bhU
w0VVcoOgEeFY0gWiLeilklafiiZ9wOJAaNp+MvfqUxxiWXaGhGBrN2OBzeimvW57M4XvJxYir8hY
VVZheDlG1gG6/O5juGBn8sv5xekdNCXUEYsJNBM4LAunGvrHOH1buKD+QLJvTfgSdAC8wozhWTL3
Qj9WaAsgZ+MHFQuUOgyXtVY6+Nwi2pX6vp2CpUN4jTQ+i+UtfZkB8Xqox3gyc68GUIH2d5+Fbl6D
ii7bptGxwkFz1DQDFDwFx89ppSaA+2kL4DjE4svZT6mmD5aPe3NJO25jjXQ566hKQwflRcnl+JCw
QxaP6XPYu0uzGPnfHdgGWAKQ67ieAtxKTq6VLnnBepOnHPyF/ATS4X79uFw4bPqt6w9Yo9mHNiiM
5U3N6oEfjQQblVVULyrNVzNn4xNDsqR+Qlbpui7RcLqUdMDtUP3R90B40HNBEDhjpUWQXlJMoBo0
akJEAMtxk1OmijM5n8+D3xLJlq5k1N0juIfRCyB1pDqkW2uLCHenAupsSehnfcZLkX27vzjWfcGY
AuA0URwiEtx8rsPngASwwUKJ1OmCRCP1jueLBpc8NECmMalRJk6Z/GjvHYfpGM9J/No93KzNTB+y
wnfmVDCPRB72q5Xsf3XvbUWEZghg4rQwDkAe2TrPug9oKAkpktti5SuWxXxjkhv/WsP3E3LcoCMg
dbYO8EbRnihPoZ/EXxR8QLZ7xxAttMnGsJJGIppQIrQtHkknqkGUNL4xJ/fxpovq0Mhbdc+ndQFc
VCuq0Ur3O08GndPW6qhdGwe5ttXJoe6h4mllrhZJN1WiG/kg0/BU+fTH83Pj4csMPHCP4lUyq+H5
NBR0a9ZtWm9qasQ657WsyrLSH5hTMAmahsG9PKInYDoFU3ODdcNlaSuEQvfoHWo2fmHIaV/24p/N
lyZg9UtMzu7Pb+5xbyv4RBWxw5iYJkGE6IJghO31tvu0J4JoAum9TPnu0raOA4zpA4NnBYNTplyw
XmucUTGsdtEpLMyIxgVRwaA+RAnan1Tek0/oRJcYz6B0ALO8z7ao9sJmcp/0shrCv2JZZDsG++9I
IUiQCAh00M9Bf01Z5zVlg0Z/f27V5XvgFS/zex/UhC1jAwVgijPOvm25iSOSgb49APlFihOMM5So
RQz2V25+RZQNqWxCSDd4PclTfNjeDZC0ZMcLwVdkiRRU6RFi3t8I+V/+ot3WMdiBIfqiYwZs+TFj
9T3uE++IEf4/nvrehpTkTNEE+/qr6dcQRS6qqauSEFrLuHpSs0pvMiQ0+Bytyew2xnPcE2BpDnul
uOAJV/0zYAbmpsIuO+2bNY1DtCj0l8QH2uNpKUiefqfzraYGgcvUEwSVnXv2NPQTqsxRaGHNfkqk
+N7LGZKbFfvJ6iYJZDVf0fERy78krAJCr/5xhO2eAoh3bAjD7dx9fwjx3vHiaIW9c+Zx+klVRqNV
OC7bB+CL9qFkCvIOts5MHfSloKGVbDzCYundQJrewcDkGeTUs3TbC4iXtnvmAfEWlIK35Go4PoCk
JBtdGNnR25I2cdqk/t0kWyKhaOICSl1oGAlgZx+DpZRbFKb0XTWhicBlI3o7x9F4VwZjQvzRd8WG
5Kz91u6Cd17SDePUNPAUbnnDJkhYSin/qbJnIzQifVh8NQ5t9ce2X8DOaAyhwZaFc0CEU+husaAs
PvFdWGpNA0lKMbracwJPI1+lbJdNXeRKyzpHYab8OmDXLbO/GoEoOX+NNZDnru6aqIAckeA54SUR
vM+fUqjJ7iRBDNLgtrM/Lk+bwaB2moZ/oZ44dmbaxeYZh1EiAxqgVCiLCAqMQSkNMSyOWNazBBqU
Na5L/L0/aTjNuWNzk5TxJ54UhDEJgidgva9gW1Pl3tWyZUcmXwUi8wxaMr5lk5CjDQDgJTLysKbg
Px3KF42SGqXb5aV+1LiGkARPfWHRyPzeQY3d6eCud34Sbd582S9ia/OP5qO04CkjBFxJebNKUUw5
s7ZcF/Z4K850UdonzfgTbdhrH5Onf7OVr1yDWdJYHV4UD29/3U/RpRcjGFZpUqW00ORxu2AQkKiO
bFeMBDl0espmVi8p77+yo0HmjWN56gKkskvqWalIvklJpOLuVAhe/wXAqQ84wCw7Qlxygc8S937x
0v97gu6rzqBOTgeTijydJ2kxgGuQHwxktCIL/ISjvnFJ766jSzSJK3TP0Ylm+h1aruJdBYvscHpd
f82cTeKb9f19YgX8Yj09Pdfs73zAmdAUmp9AHaD6y7Nz0aArc9wADJbY9da84r+uD+XWngJJyTP+
8hrG4Vx5ZRmEf9tHyI3XJ4VW25O6c+Yqdo+nvZgDFj5XBbhBNB5kXY+VQi48H9yldvdTc7IdkquJ
uk0bUMPto7gVwY/WKtzbwN4a5yRhh9PeWfiAzegTx/tof51OhEPmcg6RfAty6xUMJZF5vcYSHYg0
WHuuiFQis+akQWOtefgsj9hma2Jxm7uKaivW1WmmbTaWpj04aphq8y5poh+jg4aiR701gERV5Gf6
EFeckHo4jQmPVm/K3tWiIybXS4UUzMBIoxpkBxiz/+6PT2PMHOIEgvPoIkrq+WfIGmRJ9K7huL4x
iPn8VWBI/j0jKFbZ1/a6sP4LqysitEMM2iXdv09ie8QqyO1OlrsUFKR1HyaNO4rBpVHH9QIfDXAG
Ad8wq4P0aSeVdo1tF4pH1Wsu94S+v5krbVmWnMcPI2P+Afp3X3Q5riw03Yotr8+X0GJEwie8Wxci
U7Za8QmvCXzUR+i/WXUdARyoMyf/AsFOszVkb48yRjC5ijAjlccM4unV+AoONkWBPQ+G3bsflCen
5H7ASGHXR9TkraG48AMLUyljxCUw9kxKbQ1X37JUFp1yom9aEc0wDfMEo0WwDnUVf0ron5sLoHBx
k5/2WKFL7eVR2bp5PCofk7BVG2OiLKdbzD/QsLLcXBba1C9+3CvydArO6tYW7FOEHHOMTL5oxtS1
jR9w23yXcJgNv6VuNpGnD5b00QLSdo+jY4afHs3NZ9R/70TxLKABf8SmEyxHtJRxAuIZPF1PJVfZ
a+KmXkCaqpJEUdnqRrmErv8HpHoIoUiefAKQ1pwQzYEDIy7bj12Yi5wn6B6+OGzJnIsMTDnlTqKD
PAKzeCz+lLp0PtVZGIEeX1PbUFJE5F2rJJlrJTDNVXgvIoicqwOuRGfUiywy8EkNAt9/1PVWGeiu
+fwNAesCYB/sx33j/DFdoUcPciFFJ2Pcl2RvTmADAKo+grLsTCOoQRUE8boomfvb0lHu0wRDSIZ1
FEvExElWR4OLmf84788OLaZruCN/G0w++Ix6BeKeaBBFaE9vRuiPcoq4GWwWhBQl4eIY3ncK+K6a
KN/gPQOzv3ITxdA4zxAnw/WjkMbHDIO4Q6fxJE0KWASPzY7l0bbg6G3Cl88rb1+Zy3vkzA+JwvP/
XQkWYP9YKhIkps5f4GHKAAJyZ0zD6FFSM4itFgdPYDUocCvJeACV05Aa1YYfbkuM7fFGH6iTuTPL
2uhrCzpppXfZgceg03vmlZRlXfDgxT5Zc7Txlh+mbIzK91IRMSXkT6ePTQpGvwyuqPa7lftdH+jw
fa4NzeLXX5t2bFtlvb3hUK9RPxXlTq/JsRA+XR9sDNjqgPfPw0I+aViyJWtMEfcV7fH86SM1mjsQ
7IwyyEqOiFFvoEm5xPERqqM7gfJGBqTtgihWi8Z7YvZeyySkTFfy6dUOiicjvplmeK+DZtR0FaGj
bp62o6+ba5iVc9jeIpvMiTka0EyAacnxsXFFdqwHG/N/7we4VwTi6hfeDFJ5GJtNF0Nct+8TpFHW
NIAPiQ5XMC5h7v2vyqbOzqmWQLvbJI707yvxUzKxziPFEHVnBfkDT2D3741cACxb2FQ60wvkDoAk
rfqQ+ByxDXPLw9HqW4tr3xJuNXc5EX50VaIVAD1I4L7Hv6nBySHRuu1dQRv7bsrC4xov3wgHfXKU
epolLVG7zI9xJxdEFPlyWlct3iAfWEg0AwMsEoBUYCojf/Gqu/vLYjEVPSdcTOInubXWPgI4oBIc
GJ70R/dcB/FFAMEXc49dHv/Ant/I2MlRgfm+CAhqKgs/JtfqJN4cSdMJ7jeuu4yV05HtVIpaqHAL
5lgmocFoFc33IdxlyuIeEBZMr8fObHoaXJ6uDeaCjGMuygfAoZpxfJtOKrvuK5HONm2G/4TcJ5EU
wjMYq+hldjzwIIlOyVrd3RIyt8+qxA74e//wKZvGK9OHbFYlNKyZ6efCQkdPNJtKWkyOk9oF+64J
pb9sj6avysbKIqCwpzyBuC6WoxIyVITZCKkmxT4kXs4QBjY/kjkLRC30X18IpCX0F+zsTmzFWOCX
P1Ed0ObKK1CJFcOKb4G0m1kCVI1GA8nehZ8xYvqz8P8WDuYSwwBB833jYibaGa/vABHdDHcakFZK
kpL8jUzW+c8WXBnwA7Vju+mrYZ1PXRSxR4sEeD3X9Tps5kmYc9V31Yw3Gmm2x2TINocbI4gc5QyV
MK6eeyxCLyZPmmVlvruRHCO9GXF1+0xWjwxgqzbE+i7YJwVnIqmSGvbeTKfEJE6ggUDy4tjUy2Jz
cZqW5r90F6ABOSPJIucxOWHL1ZxvK0CR/GxlMrGu1IfOQcOnPcmdZs2KLBqHc46S/DwZiY5V0PQy
TaA+WSlhmdYYHvDoYYw7fhEXtUEXUlkZ36JmEQETkQ3xEjVyc/ZtNYXCUpySru7011AHMhATlt/m
cvh1FcfXiDEk7KPyQe3WsmGqoZN35wQ8BPLaxKauURgLYmye/LORAbyXUkZo2z8cHZDlYnMdNHYN
F2l/lKxRLNEaIPpFU5bl5hSVQwTzV51E1Mkt4t9XC8NXxzuojIkobGcjKeMmt8RL1TQSSqQoBxxc
fPDg0xclzPMCnwDBsd9pCMgXl3nlsRn8pbLXY0O/OO34EZ2WSVHAQ438jlgCzrdSZY2MBPOaPNAS
SvaB+8IpprDsaBueYJvcf5Th+g2lbd6uJhKaQUv6S6XkqDXwPlN8Ia8ryN2I9yRYXKXJm+2ivhRq
6+WXXvv0a3F7oTYEXpn4MlvgdX4P0tsY7GSq8RrlQcaSxlMIbdSjRgyFDRAcvqu2HMLB75ViSYKN
LDPNKjd26G62H6KE2yvoqM7Ou1SyNiXIHPBo9Km1wxAIrGlK4+DhibpUZpPEyj5TrVWxTBCy1OZV
fE16fy/9XYlRY7PcntGwoa8n8TOPHf8r9lbn4EdsQszHoxRC94l/vsn0iLxF7G1tyRi2yF46+Saj
sHs/iZ6DK1GMs8y+t9C7tZ516JXwtz4T6OHRxd1rJeY2wyfp1XyZL3RPfYadCO49066iIEyX/i15
JXrxtorGJhXzP03SBydbzECkG+g9M5tJKiez8F3Vpfq5Kv8vS3dvlM3NdRKZe0brg6gxQ7LW89N8
pieUfVe28xjmp6bihZpCRnO9GoNWOwmPYQWRDlYXP34s6yM5+0rV0T7gK0CAvK6PVUfR7L/oCDpm
sDTGmd1nehonxzjGRqwBuut0XnRkDKe3hy/+qXvVw51obMC01nKc5tiv4sNQwcsd9JXOdOHQ1YVr
525mt9Yg+66qkDFKrWghYJg+W7NcbYvrjtki8F1SGRN3PNE1MPAjIxGTF1lNPvjvaRqWf6ZhUcF5
IHXkoPLke8hHnFFqZ3eA9T7CrSbX3coNM0X8Bk0g4TRw0oJ9b+tvJIQOMt6uzpHYAdaswJ033SNc
9843DEQ1LnSHzoY8JfhcIu1vdqmfC5JGvZgcKZH5LMi+3ESPrBct65uhHx/r5cAAjs3hLJ2snzdO
DQSUXLQwDK3O1oADazlJWOIpJOVd4TB1MfC+3fyAt+rDoVg9F5N8uscn4nfbHPX3X5RWNXC1hjVy
lVFRuU/LQCYal8CIYse82IUAPwYx7oXlQzhmioJDADtjoSXB70S75lKJv9/sfgNubJbCJJ3hU425
klEkD7ReNxFyIL0RE2l3aVcNXpvpIZabjeiwyd6ux+FMHPU6ayoJtBu2lvlmZHMUehjXGzyFhMql
1qaV0WEbPlMBeuotmVPS/mxlWHgqgspobD6EOP8T2+PQBAYayjXSBBDMR71z3y+9HEkpAuRz90RX
b4RdEDymcZqbNLdcRPvctCoYer+Sg6d+8Oh17j5h4ydrThV0rGyhzCy8nJ4F/bqL5SOD3Mcg5oNd
ORcQytA9zaxgjAH5lRuYBL9Wsn3Y4WybmmKKtR3Q1T1DyXRlDLcL6NihJw8kS9WJzIQLQlvkZTKW
vR3xZmG//q4+JxhB8VYktjFwxNK5uEmmNi8m2HGxz7RseJrEcA4L6jRrl1e8NLctUCzMFVaZcHYn
fayY5kd4mSq2DkL5yolq2dw7dZaiUjB7qzdqREPT90EYdF+mQ91SxN0RFJMBIoYh2hRAuPFFiWLH
fm81TL++3fowA4J9lwyLDsO8ZblFP0C1Q4xxpXCt9cJqUTdEj1NSSZTvZ0KP8Yr3HwqgMqgm6KUT
EgQl4yYECXENewLkEBbXdT046SVVCPxGuVDbmMtoNIc+0YaPHeR60YRIrsI9Iak2XJx0eHZvEY4C
X6uYuzIPHASqpg8OvSplEArxL4whbfwcSJ9BhfaihxYEwQG2dvBRGDcGOcBLLjU3woFoYg2CUVrP
WwkXph9Fp/H7soHzFcVVXVhz57wbq+n38fDu/v/O3C3pSe3VwV5ghlwcIgr8gACOtcYWCJSa+t0A
o0i/3tMNZRNwQn41BGfbv5q6Vtrv3wiLbIWw2ELHOnv6pYQmbThBeemBuPCoDbrUloiwV6L2g4tA
PM5zh2ZOTTHFia+/jj43pQv9mJqDIWhOIkrnJHL3Yp1kwevOZhztEGCavo4PTSq88u+CoqIXBdXh
oROGyk5s8iU9RvvmTN1EAn1KcN8/wb4a302mBllYCYG77i4w87lV7tUcDKvdaHLnz0vht+P0+Imh
AYBTmaRQ68rJL8TiKRQGmkcy7oF1IBI4avR9T4vG9BdnwKIhngik6j6zG0lnY/FN1noS7qMVtI8Q
5hdZxTXI38we9vZXVmbvbf68/BA+PFWh5tbfnKy/0dEwYGXIZxJdpw7Z985IrwvLix52n7BkXeTY
bM+vtXfqEempwRICXYrCp/XCKjcEmU3QrLvwJMQ1mI+Jw2o5C6pmIkp1uernijEvXI03TgD7kvjT
vMxcGYK0C0VWSbpSce0kudd8VQ/KW01h6eS94GiX60SNr2VuRuDTsh/elctoqFwa9bX6UwRq6eGS
1Ar3zR0EdFeKH1dxjipt1B+tMA7q7rqtQxx4rpOH4kQfwIJe+r0wjX6cHbarTnyUHXMybarzhmdx
dC1iL6CqknNLEgSCn5dw7rJ2/SF0jP+ZHBJUECIp+xbIRiWrZHq819knMwb6c2kCyj2UV5BRF86O
USMbAHBFurKHyiq/HaVGMQ8K+iiKfWK52HYCjlxYjc8PTTKRjXkWmAqxr2wXTEmX9dHIpaSv6opJ
1fBARK6WEhVF/GySTwLP2Yyb/ziP9z4+7IVj9u6ezbw1B3mdELhU4gPURliOiZIv5RlaYrbfYrNS
AwrbhtvnKao40ssJ6KSCib9m8J5ptnNu4uoHSMdKCrXepQ224GuKihnnTdZDXMNbjoCyGYxuIiTi
I4NKbIL8GY7iSL8Vi43FxlYAWMZYiEIvGWDVowWxYGbV1jJrZ1rP6+xTl1K69TkW/PvVyz35EAPB
Ll8kXhg6ud6G2CEK2ufSHyiRGbZfmaLWLy/u+PS0LGmp6PvsBIf4J+pG10VdjTaqgWrs1tTKNWgu
21+jYH63izuXwnv4NJy5Poz8VbXHZiCermg5JuegvWERy1+Xh7Bz8fefJHFOxIYZBjh8LAZMxh6f
iyoUegHoCRpunEo2zsi8rYUGGJEcywMFsHjFpD0ershitklbQV0fsAoUpgYMCLSUuUvFof6PKy33
EXuCcnCV7j9VwbKFAWOQn0aYFa2bokzL/6bL7WYN7mzg6ETwPeD64Tth+i8MYlo5+RLlYIMlMfx4
4z+fb0dN2510Vdr8nZ4WYDTJfbNZn7LY1iQ+nyl3zqqGejN1jzzsemZ9bJQo4l+XRzhADcfKotJJ
xQV7FQKxwlFD7KBfjnNkSE6IBsq/qC9Hkws7LK8hgY5Qy/9lU0r/OxBD/BSL28mYIPV9ZsJmBqnc
DbZlpEboKda2xb0mkj0KLwo1FVaJ3K668g9bhHlKOhUmpDcS/IvH4kxOERpausKoE1QXWSuFA4hl
FOrBC3KMp8rzMOH1S5TrtQhyCRSSpz6UwB/KQR1DBc0QzAiS77+Lw1+Nkdroo+putIrHFJ0xVRvl
DZfw/G2lTJ87TBS8I22/n/bfd2WtliQsV2/rHDz6gnqZNA3mwHN9BdqxvpnSoTJ/Ieis3/2/hnjE
QtQhW1U+1vOH99GGmq3dvC/T+kNKMLj9MztKN7y+OhxPw80q/JS32wdYfnx1dGN4eXOR0EC6IqWP
YgwG5wJpiVPcVgO3r1+HvYyaXvHIyeW3PG0wpM+JTznUUGMHAQVbdr1EMAmttntwUIACKDSFZSXe
ZjSz7vCA2xwwsxBbduDFmFfL2aCPDlHRcOjowfcNEmZax7b2lTcIokN9+ptRdvtmGJoqlgymmS5Y
3h1VK51V+MKqK1t6rzBDh59W5ox769fB8sU2duxFS4mg+scVaGaPYyJ5Cm4d9pJHF6Xa8gJORKcv
mO05kqCbZM7Jri9L5vZ3mxjB0H78GD6hT7W9S1jaJm8UthBzdU2wrS4/3IqnHnwmWK21Hf52UyEr
TIt5FPPHhkVRE15hm9nF4UMjmX9c5Q7vKSe68r1isP+JL+c/2KIDtdSS9ZQJM76YjSYB+qepw07p
+SKSnSNLyY2+khz9OX3STpwEvgXIgJVpeOrG0KuDrIzhvFlA/epQvFH1Xsvb98nsa4VMjCbRtjMZ
HEhN1FaKh8QD0UfLuMwF/pJH4PKcrpP2+T9x/nRgLApnH/LvKC38s5js1BQgHVJgdyzsOB2s32jQ
WV2rtFbcV1qzVYvhy9wJY7LSHYeH/xlqW79mRug6GOg7maKc84zofUffq+kN7GTlgWMLm9SXHF8b
Oz9Ho/4IlreSKCSPt6WeisM7+m7OGgjw/N2BWPFyYu66d/sVxqXJIR12T4TAhjjY2EH3Mt0SbTj4
mRiZmBy7nhxoIu84s9DjwRAwEY+FmhuWO3lpA0AoRn5vsWgDvL/iWKJI6CUj8L4HvGrjTOTcHg7V
sbQ/8Uqdqk1aMTJK1kffwJqmgs/rkdV9pxhb8G57hFUAEh7q5A20s4AEXfxVlrlHu62cHH5Gkcab
mnIB2gmKKJZEL1DkqZQi/Te35drznGYrnQjRuIL19u+Q2buWPM03Irqs5LAUdpzqIeEPx2VJ+CGf
y2zyrQW33XYZP5kc1/Pu857V06e7LF+DF1RthOAJLrFRXv8Ln/y5WnHkxa3eynH2bAKYXwaAk6+z
hX/8Cv0AkEUhqW9Vzlz9dXddUFIErxtm2S2lQve133QsX4tdLHRGnIURb1Q6sK6axnZkKlYh6LKU
UO+kEtKXJdneYX2FKJ1r39uaKTdL4YwvCdD+cp5bgxyUsIQaGmtZXmsnjD+skZBM7fgvvlGNTmV2
BZcQLAU1yG9ZAENqAKYEw0000brFmL1Y/eDa7ZpiTXpW6ZdJG609eLa5kLWVuy68TVmcT18FicpC
2KM9mW8EdtAYQgwDXdu6m71G1AHyRNPhdw9x1trxlg+bY8BwszCzfKU0xvjSU3Uowp0pw0xFSCJT
lcR9MrKuhvNqtSWUw0ux8Kzb/VfAcE82zMyeueOJpOrlv6WOB6xJqiDdp/8VtgzitZqdvEfIVcuf
t9aae6dHkKRSW9h2MfoTdYhfvkfN880yslNZXRv4Q3mWZuTsfLbjfEP/k/b9b9eNpArU2oWfAjzU
ZCx69vsrZBFsY59incU+nBIoi73rBxyOFLDOWwyPuPjl6SpYpXUwMV4WqGEUg77CbDnibiYS/yCr
F3udRC3RKRKBnT1OmrutboVF+A/KQ+L9nYDZF2FIDGPuhDCcvdD5ub3vJp1sK35EwODkzXD5IC3b
kEXXWY1dDzQXnZQMRuxPRsJtfEJOnGgF4QnLki6ErChhIEWi2D1DIIC/yNKscoC4iePrTabCVkOC
vh59yWqM9DB3tWGllK1aSOPQSTlVCP4bQcCKtjMzcRWB2P6axxR3BQf7odIYkv8HnpcJYcNWOKrJ
i8KECkDF9BlnfOS5vLNqZX5LcGWC2I2Brle4h3B+upNtW3xsLwOpTggZ4bJwsxb9OkusQYifvCis
JCZatsM346R3ZAPNK7cBHiDGCWoIl+cL8pLRrOW0g2XIRxqhCaBTpq3rWX/X7Aye0EE75ycwe45U
2sepv5iWR+ALsthftk4LFzcfVonA87WOswmYNiuA7EDZJ10fXAhlMv35CNChGWM+IcTRU+6c7SnP
CgbtBdxPZyEnBSyiDF3obs9bzGxouY9SWUvOZ1yLjiW8t48e0I6PAz9ppeMq+wjcE/hsclfhqVRz
JPz6Lmfj9rA+KmFyw+kjF4AjKLvJV035IiCucJn9XFcSWhMcaZha5sHIut8GSJw31tmJyO33saWU
6216YZuurq4wI+wPV8zKyf477KAHcCimwcFCr9adXFAfQs0WP7/fKw8VEQGnGLIVH0XasEAyoLZl
15cK95rj6cKFPp/NkRDoRO/rQ36EixGlPJcc64rb38S7rFq72beEAHLkuC3QRnpB6sSZB7/PYLhg
ySgPz2WaDIMYGMbtaH2Gb1wTWKQWH9B6rClVPkKVcS846ZLA+kiDrmjrAyIQCKoHeISiJpc2kCuo
HFCPmxBzfaFWu8IKFomvfyWaaIByMqI80yRFn+hCPWS0QmVLF0jLgsQB2K/IRQuMEr6GSkW7mz6o
VHd+fQsFJ9a6ts5E/jklYPB5RLVZUBXBr1j212Je0K1ZEkKBBoBywJC9YlPZJjRjwXn9RjBz+IBy
m6EPWhcW20xDTDZxeQFhV6GVgtmmA1KBrHMh/T4nWZw5YDGSf+s7DpT+1wmFklO4CiFLSCp/mQNG
m1n+y9WhTQlv0MVIw4v3BYOyP/OcFya0bHXH6JIyGKwCvRx8JKBFwgvXUlVBeXOC+ESCDfPwXH5h
g9O170YS4/ZHiiaNJaLJPYeA8Ln1biYp60eibSM9oeoY4NMGHwcOjKbHWXu+mGs0k99IdQhKV7d+
2VqR3RiTXn4BxHKKsFZtb7ffs9HfloAQFVVebWQrTvBy7WS3z12eLZ42WahxfIQsYfKN5UyQ8KJH
ev6mHUKVyQTFp9pFd8oaGEZCdbOQjHlyCKgv9VSk3iLqDClNWYyNbD1JAbR7RobqIJs84Uet1Ohu
0LY9jLuU1KLl8VewlDZUk4sot9kqaDPIdKVf9teN3mtYk5kOHL604X2ERbS0aLXsa6zKt06/FsXA
Bb3KSNqVyubMRaHPg7N0GpjNjTfrQ6GsYSDGCzyeLBqSI34kwoiduRHRGGoWQ7Zqs9U8X6y/LoqJ
trJBt6/0Tc8e210R+vvNZlFutkmElnwiQs8Mw7h6KUEfeXzxA/E6L5qGyRKZ6lFwRjkrc6GV47/n
MXSo+KZZKsdwc9NfRnUdBrovli4SWqYkTITxdl80hBMtRkxKsRaMB3RLmdVCND91quDEV9atfzY4
RPe4MyPYjJUGrIUbZG2M2aZufQBXlaWwZIN+gtV3E4g52LLkoo7PTKTCemAW+fChT6j2l7Hjz+0O
u5SKucMBiRe8twmepD6356s7OMWMOH42Mr2qoyhsxA5gVIYqmD5amxhl5q8VLfKmk0aGNGStOuNL
pVR7C2P13705Z5NHPpDUNGDWrBCqaGBLO1WSu/2PwX7vqlCtYgRiQNw4Z4Q2PJb0lGNr+QwoFdMe
8KCqsuMznvgLfZluTDHtblHs5qtMNEaz7JBuxtoovO6FEWtJ4Nielp+XHmcTtDPDQ+kz7VUpcJzj
F+PYBDc0pQvapXBZto9IzNuWE6MTjsogFz1LKatCQ1zExn9cVQitv21XmWy00EsKGWwD/hDQFel1
pR1geMdZAB6DM5bDpEDI40TNhdw5U303l0J4aEz1k6bwdOCZjQtbuMTlQP1OpSzr7Bs/Ma+7sm7l
JUJbANNTfbkSkxeh1/L4wn+idWXoDtj5S+4yiTn48E+9b6YSf0I7UhW5NFThCf1LEGrtWZwMJloC
eLs/MRYny17yVtmigM0XoGew0NShVMJViE4V1Hot1wgZ7gmMBmRIWMJEa6kYzuFeY37qJt/b492T
k9roq0jsQ6G8N4c8z+r+drws7IFfyS3EVWhTWTvrLzrcoJFpv0Ny/IFuqu1XxcEbrIv+HLILBjW4
9J6Z37kNpQ2YnWyt7QtlyhJj4xGZ0Yz/Eho2etB+Dafi7I+aF8Kq8n7SMlrq12DAtx4nJSQPqtuH
6k3qUJXIBACyS8L4rM/j0vXOXMyP0GAVpoaiKUp5ydpo6Uel1RuU10P8uqAy+yqx0JEKWvy0jtB2
MgGfbsziYkDBpc9XNZS2AaOiq9b9wg1LQq/T107Qsu0cheZWgsapdgdgV/dJ7u0BwWS++vIzo4+D
fl/uXcyPa/Qw3CfWGk9rReKtF6CWs3EjuazAwkXhFYkYvyv+ReJ3oosVvtL4nGDVAeoLVjWokQmC
iw7pR+cht5RQQiM9jL05OnrfqBOv86QS3QolPJo9ZCynsTlXWTq2RltWKd8CdPV4BqIj90aIW72f
Z7lBqjPJojuand5yZTAMciOPH05lzAvI1HiT8J5czLBJBS+42LTO2ml0uUkN+OCYY/7fhC6CDsoF
AVUrCqEYR7VLN7s8lSC1zUh09Ts43SQXqVktUhAAtms9s719wwtxiBfwkYCxdA1CbjS6YJ7nkeSv
ZGo8/zt8gwWeGY5xWGFIMF+HV8cmkP03KZRR6kM0dLdMcFCUP2w2/npHYB71vXXxZOeVx2FU6vFV
JNfyzve8+aj2rQMuucejqGi6Jfhgin+gn0myygCY+pQVmWihJCvFusBSYnqzjDI//mC9KUSfpx+J
+yaJl5ZCgutYjgl1PJ5TyLZlixjMvt1sUq8SbnGrU0546bEb01/mDjqURI0Rx606Brrhq7HQa+PE
nP47BUDVyRpdzWv7IAs/jn1wZiPXC5DeTDeXnA5EUfQrjdWxx9Eg9EMeXjbdPOhNXhF8gH+qX3Ad
Of3ed41fkEs1Ie/4/FEeSF0UiBlQAQb6ruj1KDXoEIeJtxaOzctSgGiwwL/zLkMPt6tHccv4nOkr
ENJbnLS/HzIeYQ2bbEoqntA0JewzUnVjrujJuTj4uRvXELiSfNS0XCZByBHx6q5u7QpvSu5poxID
eoBdd5ZN6n0Vssg7IujZFgYE7tFxzdTbP32748j7iAP+AxM2ofkYsiOywV5C0Iv9eHGPEd3dRjpH
VG1nW2Db2OzpKaF6xVQthnR4ucuIbRGrJ/UWNP1C9c7QkC7iJxgGNGdaYUED7qfeujKumIqLeZ0D
QCwnfebfH6A3sGM2A9XJ/13ZPdJq3pc2rKV41JrmSCdfIcynmf3eMJ4l+eHwd2wzghk9oc2wgA6v
LiPAJp5N1GWbhH77jM5CcngvNrQzXI3wW1nv1rEnQkvDY79HUahebRMBxYLnYAbDPavlzAqu9B8J
JkKh6EqGVlp+muRgBgcNTNwvmYNVt9vH8LL1nUEcKVoE8MYOTLU8iKEzgsjN2DK1nXKu5SWo1h0g
d7/EHyeiROs37tM68H9273sRf/oA9jdpbj87KXGR7WE9VLMT7axYIFtLNhb8pzlzG5acGMOIVAuQ
Rzi3sLimNW/r2mMPCNkMNDMHlNUq47cffwKagJMMZcfJisyWHKiaJgqCAUs7sOyWLqiFQgYYYkVn
0bs+GNVOZpYQpHQOS794nSt8fOlaiJ6xZpD9OvhdwI83BQqBKnUaVyEeeAN+yY6hjWHfuHAbw1GF
O5CZN9B8lFPWWp298sDiHSCbrLwt+NKgmHCMgnOfczea8dmlVX/JIlBcfF5ovSQ7rsZ9dDpRQsq9
pYdgLrBDN88RTPHrO1VFPulpB/MkHCG+hSZJICrUB3ObZKq8sQ22Wrxk8EVPmUjHkZ/iYAVBdH+t
S4o39SkRbyu7TGrm7xX7v4p7Yfte8Yc8PbXY3YrZjcVF/FgCCokQoOno8lBCqSludPeSZ2Uqv6un
TE6ZSN77dSCRYD1cYRUBTpvzGYsgvRfkd0mveWN16yMMsvT8EBzckZEaRYyMnMCqdnRVWinYhvYl
qi5KDuzMaO4d6BOCmgQn1suV0G+vmdt7dgbIwwuHYlJbzxc0hCR6eiLSqnJBI+SDgiy/9LJdwOsM
vzGmfS/0iWG024JynyXLOHr+qivvmtCImWVkbUn+sQp9Mx+qdT1EDMMAdd+v+xc/Tk4lmmxqWSR1
eDyKxkG9d63CZZm46RMCaG7OoNIHy3mC2wZvZUS9WG4+QccamxOZHjtj0uJN4Ykd5YuNkLeFAoCS
7LTfQ8HPGEyxIBS+S/HMa6J6c+iyALyfqln0UcQljk20ml4LxSGhsLrWaPR9JmIhWmLRPK1HuYgv
7GWm8p7/f9M7iDa7RbB3ckRPFpA9xjtJy4V0KhMh2eZZYV3C+MTvrZUzD2Qb247V8vUL+/I7aZkG
t7mrXQmTaqkoz926AO/6C6lwQbPRodsRV9P36ui0hnIyuac11FygdJopXHCcCyZ2pe6vKg+6rtvB
mRWH1LwC0YwebDyAJClQhFaUCL+kH8HaF573N/zFGQSFHia+rAcE2xDLNh2ZCEEAH8m+2zeLd+0M
j4qLU7x7geOSXhXkDjVy+Fp+wiHL2lYeKPkmNmYrF8hECKqURM147PvMdajGQ3N7vhPUulbLb5A7
XX8I6O1nQWalqsKeQd0r7jqpkdGw4V2SS6MzOpaf4vAI3avLu/QgBAbp6au6wZiEagOrHGyiVMKo
LLjy0c3DuxrBIRD9PflzCxdtR5NvHKjdv09kRkhCaTdfOiRTlv4uOSkVOk96tJjs4FtU8Zta95Ci
djDKso+P9jK82zTR5UAqYvQ3y3MFvMFQ/Tusxf2AUlXtC0JzooULsR+RY4rPNqyDdOmrGG+szJpj
2nx/EaRr62PEJzhqso6xEC5+iMG5wt3ip+iYfhn8HWs1X9ZS74YDxCjoFmyJrXs1prkmJZiCCjDS
9NG8XCeO7oT1so7mGfPsRb+udUSIJdDtDlNYvsNVwcIdzBRVh9eyKvteVY+jvr/WQ84SC+M6Cs7h
qGDZzDsIWbDrjM4QhelAvl5RlTAW/O/8xwE8x3liF7PNGMdhWPyun3bq1nKgAwhJ0kjUnD0G5rYv
e0JnTRy9uXohwfo2Hyum/nTEMQKagFi+QvO4m9e6VTpWcbLFxNflRj8Sas8M7/eCmVaCv1xLfsBp
sxlxGCJcMQVyM2r1NhSDFpLW4NmROZwm0WIG9JyfeCZ6zkbvJXOBrpyVGXcMpxppMxuUPsF5OPDg
bVr22t5L++sQ+A9yLtTitus4euDl2fWIG1tNYSBNo970kG/nAXQR/DNYWLt3L0ObZPaYQsZ+vl9L
9q+ETdSXtGrpWAzOIfmWrBGj5LzX4tNZp0YpCnozBhpUjikN8n9y4IucY/k4GFMkDKoptjQMR8kN
UvbAeQKA4+bBwaUfM0D4knDn5ok1WBNvnZ/0kaFPZ4SCmUMit5wqUdIv+B86dHz1McKdpHZpTahC
jdPQGDJE1BOGqio7+WmAndUcG4aJ6ZLJsQfB0sMkarDHVE4u4vjWIlYTKuBQ1jie4UGpPNqmmKLX
IPWBkun36PsrQ/d4M1UUFChtoVUS2RLTZdg+NeJWKXd+OeiAx5VHC3giRBY+cmocZWuEANYy7OPN
9p9h2xEt5l+mOVvts/PrDD5cqRkwbKQNowfkKSjBdbMEN4hP8SnJsgTz0NsE0iwYsn6z0Fr8qm/Q
K0MbuLIXmXUBFnDtStY5iUzPudfhhgIiZwUaHCvO/rRnb9t/jo6h3cr9jTw84iAtRfgwNIei9gv8
uWaSW7Y+OetzlCAQHvVWYsqS+k8vd/dxEq271BVN7CETnKtQpp/OcsCZBjPywoTlTGJwIyfELXT7
10VlCkSC2epdNhdrxVY/Cl5QL2MKb2rXlP7KNuAasExgYdCSvPiK1/0dVY4rsFvD/nC4J6jVQUXO
yvXQjw0n5AjTCF90KeuRgO02GpO++WLt9XS0dqjlDanhTtpfUeczYZ7lz1BTDqzagteFsejYtSsk
Em6K/zG3zbmVqPOm+SP0k2Ywjn9qXOPPQuCTl23/arQp8fg5J1DXQsNcOPeMFuqIHWLzwnDoeF8A
2ZHISQ+WBqMoAh+TYD/n3bV29eeQCOyrlBHY7RN0A+50XGhU9OjiaIbkkGxH+bGh75Fj8RRaVshV
S4yDmj77ie+vt5cJAlWuOhwV0OfVmnylQywI8C6kRVOMDqMeA4naG7ZaFnCD086tuVdU+UBEmxet
rrMFRB/Ak/X8ZUjltuEP0u9PVtHsTCGxNTNE0a1nMfrGNfL3k8SGDJ9DmZ4xzYJF7ZRwzDyd655E
T7jTu9WOBW2HMS33xxJHSQYtMDDMgwsIb8S5bcbv/fPFMd7qBavp37gF/xpR70xtTMkcWeyD8GrQ
a42i6PuODUhBs/pmC+mqQj5v1Ybgua5N0i8oVoV6av2L51TABMnxQ4tGfYzuwp1yWq2xN3rCtWLw
iYsu6DHu2aPWGdn4EmpSj7V3i4l+FaX5oBmm4XFxF7xp1NBGHqJT6nGUAXAHMpfRid8A6udwzZwh
cwe73Z+FLkBDT0k550OyYXd/ZQrajPjZ4UmVZp3sYNc2z4n47ylfqyhA7k2RJkt51juCN2LFFR6C
ecwB9lxSpI5UII7qSBhL4LnMSGc/oigoLpXOtOiKYvvH/PfpBjUgWO67CkTRvCwDHz3n+VY/OIPU
ZVL1BoA3bMKjcavkD0B9FUX8k6gRsfMzhWPyyDlR4RzRZYOB3TOaxM7JF8K4V6J4Isj3mBXPVIFZ
pSpyLXDEcPJfGGUgUGd+PqxP14qikTDAwMLD+W/gTkN896T0JslNOfILV+FrFECobfPH/F3WkHfQ
9CLIs/StLXsTOke9TqYPjQPwcqu+gz+vV/oCwuxYVHmSsKro8F8jNxmkVbQuUUOGsZ/jD1+LU3fr
d0bX0NCnLg/J7QHLaJkZ3Z6UdCdE8uFh/05f2IydQZJXyOCTw9zSbwhGtNX+NWzCtbcO3Wwi4T+3
/qQRQOEsC4MyDWX+hafLdasCT315UHilbK1CnDegLKZHwqVX8OLXeDeR/JahD4H1bIHc3qHvcNSx
gIRFg9oadeYW1vq+4dFQnYDw+2iGmrhiF1ziasrW7pK8l9eGilvhR9OQcdECTnGtes47tmY7agbj
ScS+KECc70pYKVQHNWlnU9mxatogNqagSKLK/ufZqnkX2I0srY4JCgVJu3Z40LGD5JkHIzwYlc55
AxZo89h9aczg53FwSPZthrpWOqtOJUXWs8VmVInAewfFSetAQOPUfIxPgBXM+qt6vkGpT9YO5bpO
8+tSLABX3tCi39V8mDUbkDQLGuURj6XsHPQupMwSkbYVgTYR81Oz8gFKgdHr/Fay07cbQEtGxE/Z
AxCg4qfjqBNUyI5D1bSVJaa98aoS7eIT4Ru3tdCtrGQA6M23sU+6n98DUBn61XLf3g2FlGu+F2xC
d2cSdtzyStn/Uck1e0hqtnZcHos11Dhhbz8KKpg5kAYfg3fNBarBLdE3xCFfzjyFo/5Cr0cdi6fh
1aJ63YYLdr5OJ4fIPTFf1C2Am+ih3Qn6kNNL+HmKzuNCcrZj1W1eo9kF+w/n3U+G4sjFBfZlZQSM
w8ZHkR/RYx3VgEVxpfJ8qPQwKJMkG9UnP3D+kDcYlUNuMX3/Te0iizbq3paE+fo1BZUlZCkLS3rA
gWz1wuu8ro3OGXWWsJOemuzfcg0faFHYQSV8G0HI5/IDQAzNnWKGY4i/8BmrND+OgvULrRYc9WLl
fthw33ahQdCP/IjQrQ5BnJ+mHXywXLqrNciXL+YwkzcpYo3D3KtKaC6ORCRXBVspBXF1VjUvP89y
doPUeyYqkQkeq2YRQD2+r+23OutpLynFuDadNTwXj2Yf3W5shKeygYwZmx7cIV+99Fm8bQpxcdAi
T/n78kzj9eZwvzSS4JgS40+wQjuQVea+CzxGr5QhbPvfuXKzkXU151ikfOOISP2EFGHwCf3i7jwl
Jw+XFfxqAOsTAjQs5Z2KDndn3JBKNdx9umWXlZCzYA5AFYC6/QKHBtkHw/yN/0h7oHTKJvHOJ7n7
pik+Tyfl5bfH2tCZr10DTsc0+pq8zr00HgpdC5CcPHcrD1OeG+uod5OKeNqFry62ZaYG9fvWzoBY
3/FTygcM8PilVTBzwxpTLjosjzZ+C2TBxf1rEXIbMUeWjjBx0NXSHHh1mg6XYcR6AUS4CJxdH2lP
anz64XUL8nvH6qfO44u39a26nImQ9MUgTA2YXoTLwl3czcwK5jjc/qgOQFTvZ0O3rpT1breKD4Ig
Ke2WkO1MU9SvSHDYx1So/vlVdSs51O4wucLVpQsKfVFaJMQa0Lm615VAK4eOfaBiFT/j+TdVgVK7
KmMuKm9zW7t1o4VHZmpM9dc6KYHuopu6h7BvvKd96XOuQuM5CxQi41V3Ynbo2dmqFEqxGruz5DS1
6JhImLmuJIubj0AIuWeycd4hXPV9kTay8S1NIZi5gK7FhAvTBb+mFkJr7pDJzUkitmu1MPLWaQvr
sqhKaUUabccVRK0rl3F/kjDFe65rB+GZqGZg0DZFLsx9ASOQDRTqZXVIRZJN8AnlUZzVaufmz9fB
yrs42MiywWuXSAQCF1ViseogJto5jI1P5Q2X6EYrf9aokSbESIxFcB3Pmw1N/QUyStxCIPdTcrYx
pTeXiXvdJB1shUsGNLVFeO3C9flzocLCiUJqCniWfq8V9aVEEA97pGviHAiXsZyXoN4jQUXT+ATs
dVfkW9aLLy2zAWoq6/RKsHXdg/V/ups/TopmGST62UnBLgEj1V/HDFj5v1gJa9DXcMPsSwMXk7JG
9o+Yf5oCilzpde4nwdlvSpO5qPCyxvvcdQvzLuqkiaUNB1BtBLoxPwpsUkcIL+fiKbkhiu5TopHd
6+ZqvHodVZZ6bG7iaqZMJFUruUpwL4DyeqHO7wuNyx/NV3vO4dhU37L+pGK99nrf9GLCG7dNoECq
14j4F97ujEh0ldoWZ15sI/5G7ggCBXRqj3nUsvGHHk9Qjo2XNMmnbQWHgaEAJnqqOeDRF3ld/RLJ
jh7zYPiog1GYyFF/jHxBSAbZAeu/gMNJvFg5wTn1zbPWxG4tVoGH6btRELsEqQtiPGWYvhUJz7qq
l78yBHerOoWVnH16XZr/MzLaO1ICXKIDJl2oNTemcTLWJLAkNxtL7GFQJnzNgSLOAgV7rFTPGe7+
7dxoGNflRRHt5VfHz/sb2b+6kJOjNdAKvW5RudyjN4B6PUkNwsA0xRwMK5RMiH+IuCLCs1AbALAe
9ilO4uZGw+C2C/a1xo7cwgXXHFRsduvMJkde6EVnvMy0QCapD3PQccacdOmdAsjyTeuwH+YjWY7F
Mf5g1FVIywPx0l4flLS+jZM2+3DHRGmQjXneVJpw9JbBS9qmbSURTiDIhBENz7NgAR7wJvkLRwkg
TVdLWHu824Y3avP6I/2TK4w3dpZ5AY0R1lVY/VrXbFjMKYsUkiqAM3oSYH37htQa2isejWC3nCrF
/KiQ3e3g2L4gejsZKGiwfpSDgsGzNhGg4RGk3+CycXrVgvSsJAipJvAfbuvRKE9j+sRsBC+kaTXa
qOmQvfn+le4sx7/sjT51MhVmTLlxWDf4fVswfTD2cBtX/yXNKadIlak+liGPjoHc575vawpNt7mS
+8UjLLTwqgFPw/FRyC4ElMJ/NSSwzwzuXfbZ2c94HMa121PF6X11hvhYIjPkz/SVnvrTyVnFWJDB
dtvi4IEos4P79K579rU3KhImhNsJc0VPAqRh3Dn7FX1ylJvr/l5j+6yDSb78002/y+ms5rW+XZGE
J4sILtWDA+233hvWTvQR27R2Vch4UoZFXlCJYtuGPvrZqusVVZXSec1kdXYJR49MBTzjvoGWpqMr
WlwBhlsZNwgvaJrqQSgc1j8kxH31sy14qlS6eJp5OiSQLkFTvOsEx2tDQZLjtG+NohHfaFpbqx5h
QqcDartZb9UMV30wa/W5gkyql1Uk6FcxVDupeJDjnT4BhZU6LIphmiqbXjiw06Bakmndl0/OmUhI
EHVvgGnpWoqclF8u3GiwZ0E085WnUjjZnCYF10Y+dbdl2wtNeyh5usnhcfda/G03nIQcsK7go6Kw
is6zdfWeRrH+9Weew9AyZJuIGHEgn6ZLEpj9xeJDZJYN2XXfIOrOgsdlBhkeg+JNVB6USulwPEpz
2LfBToYsBIXZEoyiYkSIosxGFWyDPcqnYaHLp0A5hE0bm8rrZ6MwsdQkbwPx2eqXKwCcrJeQcdaa
XAvXDKcqCkX6CF8qBbrvga1lVi2IaaHa+0v/uHT/Ac6YWO9izor9oKssoPtt3eLWYeoJvlueKTkc
3ik9p0TKbHXTqudmnCMewiTKO9p3EV8pc/Tf354uY6NfhBqcw+bQ7r/wrg7RDNxAYg9+FC96tBkw
zzcZ3D29OBG74NdgT3OQGmVyjZnFqz9LsLyiihLJF2wnkyoqEbj79MpCvno2dtIVGQmIjNx/xUIN
2nx/MEvjQHoE1kzNQ0KcEqyg/wSGQvBZ5VOXAtXpoq6byDahIK+qJUujl6QWYXmoNoJkDByG02Zg
NMziFoH3G6V7wa5NC6aydiLsO9ZVYQqXWr7MmijiMZ7BHBIJmgWJ/wYUvW65i0Z1jCipWI3zS9O8
of6ZEnpIyRYJEk/reIUKv5OYvD3RBeFDk/wrOWx9QDZoUe0tsRl1CSt3hQN7o+PExeGmI4IvbxGC
ZZiCiVFUu0aQUrcGsjPg8AN/6ZJDKY8CmfhPqOe3e8AAUQNfzXFnPDdTR4F+q510zmD+q5PMzWX0
BNaVCX+/9SrM+X1efJyQM+GOkQLElCnBLXKTbcxI5p1YmsjJlxXyfMyomxqy7fRk+4sR5tXLxhT/
Hbv9zH2fjFC9CvRtMmfNXizMBrkOQSxtNDT7UUPNyO8yjVgE/XEy7NG34avB6vGtFZXtLyOBM+io
Qk8uSjiUrXtqj5XMME+bsOIg1MpfUc4Jp/0fB8JHuLtxQmce9yrp03N53L88NiRQB1VUoCvQHUoZ
jVV4s8jmu9SUcmu5xD9rTm8n7C/GdlJOfMQZaAc7PpGP7nkmWygCK38zaHKwmqnhvNCV5AdywNXy
r5vxojh/GKDrerHqtOmalzE29cHBy+iRi2Y1Vos+FSml2X3ppY8RjJ4OhgAVAqzzz5GHpEmZnnAj
sadtU4NhC4AZBJ00KzydT5gG7QqnPYuTXMSna2GCaZC/FKGDMjcY0IXyXzvHOWrwjYaKlfcDmWWF
QL21g+9nj1Gj7MhKw1Mas5rhYtHFwS/xj+ZJ56v7DIsy8yLYJU+e4t6KJ9XKWlePaHj3p5IIYmEJ
Ze4KqZHzq9h6yh5jYQTE78mMTyQwuwaN1sn35gd/CO8V4RgRGBBKgxTEzsTg6uVqWbhynr3fc2wX
Vwd5Nl9Y505I6fOmc37CEVJrPvCH2cdqS+U6eikZmtoFNPBd7P2aYrrxjR9hlj94rIRfdoSkN6Be
qXP+5/GexIxsXzDpWk9yJtnCdRwFYU9XIFHnaZ+KfuZZJ8wDfg2aLer6Gfaj0Q9uiVsud1pIPov4
Hml+8WSx7/AUQeuV2BQnGfCP1G9Rlv10Hhf9gKHUb3IgNsv5FZAi893CfTi8kAtpRQZEx8k/v1S7
BNnjFTYztAv6UmuzBB6ZQTagwdrQjYRyKvocMttH+1oqZ8urlY6m6bcbI/QkUlbfZgee8d0yaEjW
9daTDonXEBbvHUHaQ+mIdX0MpfPRTaMbA9GvmwEYUxPDtIFd1T+6vN/VcGkcLjlyrzwzRM76U7Eo
yJbn7/GcckI2WW19M7LHwjuNxKeU7MMPQhLk8RKc/H3DnBsOpeKUUzrYDxesKP+8363mXKI/XKKq
Z3UbpThT/O00X7Chfymgd/eyBxKx/e7XCaeb7GY8256PnDJ2YJmbg1f43l57G8b6VqJ0UqyxHnsK
ltRw6KcNrKEWNpqPCeWCYkYJE6tsZcn+FTPBbilRszMc9+Wz3bMW6MRNnAY1k4qJtl30kNIU0Wqc
HrN5cTdvyT4Mz3hAYWH4N7v5MyCaA7AmnmQhO5xlxXyjUYz9r+exs7YBCcvJxG2t2A5KNuvOqlZW
F5rXsfQ7VBRcBZ7ao1EWAURlcNxKhErI+fntcVkCrI10zAyYVy456skn1pxwN19F/HEjbOg8/Y8n
u6lqyGfQbTQU7rEVe5ay8JMqo54NT3DfA2VfqFPdxEd90CvT77wkbZc/qabtVNdXEu3BUPFlHjbC
0tMSP/qIRLgNpzacSJFyUeRvVNgUwNUyMwWKV2BuaC7cfpesrw4DYPiDPAaNPh6uYsxTrpEOvkUv
uqCRHol4teOHTbHG99g1W5XjfC+t1xBgbmA6fZAZwHCLvMwUrI73b9DZdScmld3bMbszR5WLEMkh
AUqDJdtCWVl3rXM1EJXunOLjs5Hd/T2gub5pj8OnRgNq2c385ebvt9Ehk6BsLE1kywM2a9vY2oyZ
+u89KBXUvzn6fo63CxcRvyRHVifGPB4pzpQ4SDMwgaiPAjRpMQoN4jH3QnenL2wBeslgRNZPqL1q
XjmWKPsyG0Zs9YaA7oB8Or7mi5KwRvtjUWSjMfBVQI3Si1j4/62fglErHRKPP+283iwTq0CDmDAW
dfMw3/eHETxHRdW5UwNk1Ns9S02oqtoVv/YMxO+7+1eELK7vcOInT2tc+DwwqlT4PgwtPHMUKSra
5fVi4cB1L4aIeqxbkJ6JHGHf7SfD9Q1V9SbGpHRAb4TiE1C3zoJQYrTo5fEiR66g1bpTATjSLwbC
M0MVdxQh9IAMzdcw1OvPnzlwhiMPxyngyJYeYHIJiybHnmutL13qs+JFREdKfNLxf0QSfnB5cJAx
7BfGD1BOIHdIPyxLnL/xjxtNVhuLA3yafVtY7gm5zV4/W6IAfG3gopfuK1rc4WVs4U13d+4bjx58
e5Q5kk85ybmN5MzyoYol8bmzqRljK8VcIIGIHKDagfANH1/qRQTRaHBdeWnoTKZTzCdS/Z71vPJp
EsL9d5R0oQwdLJc2YpAvSiDCyDVSwk+Tnd5HxKj0wkFjdZ18Vn02kLri0PzzwaDRxo9G/uEdNEqD
cK4PWnG5xeOfr5vgnnXGcYb0ngXBYxv4POL1HkYAKHPimJqVr1FYrn0k+oY8AiScEVM55uFYOuKb
rsRhehFCkweMDCw9I15XiNvUJMz7mUFlAVL0LOqkW2gfArx3s/ZZYb3KJkuVtGoeF9KxyJb7cPZ6
sVYDaMGFYuZe/tr1dHwRl8HjHUSDjxYYqg2eIil55wMIu9t03Got/ArhkKgX9R+ZTCyEEA4OwC3V
dKJB8BlXI2MTLyPYFxwDnz171+4i2/x1OQAtBChaDHxYFf69vGSeo4gPnqgn8T4vspy+aqR/RSYk
j94sFvgmrikTHPHHU8gMOni2uvaNyWAvT7YfKNXdxQ5879qyFT7y64R3l8XtOnkoOXihD7j0Jm9w
LWCabVK/Q97270GlaNS1t8iXe+THy0nlQdBaBZoWVBt3SzTFWjyMZC9uL28dJoFhxXGbQWEOSiY0
rIbBi0m4FPiLk2IAoIw45Bfi2EW0HZKPhG7geabn91PcgBmCqxfX/7c4aGN5LQ27TxwoQXhLOPeD
pD+eCmKMg204RrJMVsl6J4oeU+cIJSYB/KKQ3eekwS5J3HpTq7rlBqaxbVvGSHIZTwYv93jGxvZO
kPaxPZVdMEEJqUEY5i5LW1Rsg27VNuc/jy57htXRJi23/+Us+L4gv30/2VDcLoraviMKlQTg1T3c
3aMR9QdeF8H83MJNI9Oe8KpgsK9UPNJqOErL+IJ1n2N629dQYuSsO4kZwozPCeC271vsqA57I2D2
j9OMYc9gmKgH/17KJIIlZAwG2+EnCk2V0eKfnpP3ziYCtq//Q3ZW50dzkGUUXiSFhJUmkwjfvizo
JSfXe9hiD8RFmLRpr0HT9WyYvs8BV350bk2wf6RgaIpFxxRvbxWlNRPYCvKAO90OrQZIaT26cWV7
PfcXhrbjK0mJRpiGuRPYWMc1Ja5FLOQa3Kswun4cSO81CXE6J2VoieoXXJ1zvuM+u2S9A4/g7m0M
8XyB18iObHxDb/6pxP/7Wwf4bjfEWe3eUNz3byrfPSvxYO5cm6dLpAavyrb3OrSaF+tZLslQK90g
uru+MDHdo7LCPfBjq5Cz2eNOWQSQm37ceoXZEc5ZJPqV7nV29kHMY/D37FRiay1b3P8owxXFFLMO
BNTD6JHmd2WPrVavejDndw+jZVOnjibpKhguXnNG4NEPbNAuJZTDj0plDxyNgo60l8MhB9zjVUz7
iZbvEx4IEiPFjo5y7Z5fT1d1Pb4CeE6UaQYAcOiwgFW09CczpW/PFiEGTdeDS2xK35F2gHcOt5jv
ZgGYef7Gwk2hE6L1AOf+pp7ClQdf1vKlRY06rerFM6VMJHYdwt+j+sKyRS7hvy/8ZsCzLM2nh72f
IEbEgV/t5OOoyAHWp7DFKB37k0YpSXaojalsUmRkjScVxYpnZt/wbMHC6k6WelOcU323HpGp2I0a
NcJ9im0LdZNS++BBcHiDYZa+dCShpI8a/N5jvfymo8OfHpdELFFZhRbPlIv87asqK+PSleuxwCen
s3liQutW3U32xiMFdVmYCBnNOvgvXrjqkUx0nxSCTbPUN04AetOY3g3zMi+6qL1PXB3Wb0bzblTN
ok/lAtSSVg9D8aVbBxh3XwKT7tMPY3pEie5zdYhZqybN3VzbK3lwy6jfc9Ds7X0v7HIkkdiuWLDs
uqzBLwToaETOsKYD4i4GXbIwK14SPcHChpwHowDZSMNyr2rad3cCElgDfjSYvewcgvr7gqU/oWIQ
VQ87sYmeqz2XdYF2NwlCC3tT8+ZiIY/T4im9/clNDnVkocbSIPtjekzrVOQ97paVhjLnjXUWJEQS
nUYkmzuSTJ9fhSOriRr0vCIqTUnENJN8x6aYI5UoppuHTFC5qpCWUQduW8yNmu8QNiFDyluAwhM5
KK2piXupdpYFl3lgrztH4bkZ8kRkDoFBPEZBol1+nS2fk27HAD92xo43vOAMKd6ERYadQOTyL/ks
OrGag0wXp788FUzSKQlAr+fsltjSJkbYXykzohVXiYaFp6+pF2LHdeY8DuIZ6GnbfJiiswxDegzA
s0i3hGc+J8mkOnnmCUDh8YOIkg/v+9Xrw4aIPGSi3ChaFrk4Js1wiWx1XbBDq7Ov/1WrcznJd2Aj
h/GI1XaH+Ci+hGq5cApj7bWj/3kqYNY1bM1n8ynOHMvWyCXbP+fHdBdrscTe/nsorDkwHDjCWLNg
ZZrLfGRI66wWa/WNokjGAZpixUL+iGjtkqMlqAuHjJH18nq3CCVMwsgXwg2D0cnqxg5hT8HmdrNk
U9ZFl49Uo2OEkZIw1Ju0Z2ag+EsbK+PGA8TKggm8YzoaB2Mh5jZspVgASggD4H/OSXH01CaBGv7P
9BJ0Zlbg8AxBDKpujldxcJz4V/5/x9+xfOZQVKJfLs6m06LmVQowdTzBbKwkFKppEW8RVBf8b3Y7
aQt0WnCBtDRSoNtm9FB9q5sjsh7la7YYCGdl4OR85oM7DrVwAqmwFyM0YoLLztlzTszB9WeIWXCL
ASiRMB5qSxZBTlYUdGx6ymsfnQv7OOIOzXMeSbqIXQsfZ10WN1/yacW5au0YTQMv6f0qGSLY4hCd
uinqyrUi1NG83E0jH/F1elwZcTS6hWE+hcLiH/u558+q5R2GilmbeP0zBtNkQxJz3a2yOJO4qcss
Iqo6Bk2nZGEgaagt2VkeaSYj9LI6xpH0SEekZ5LA680cc/QvPkxFwtbapwq2QCWSNDmC8sfCjCcN
Fp7uDryq1r7BTLoQggu7UiW07XxAT4GMsq/+4cZ2mhcmlOcBfCoMdWArsjzcM9U+rHTOyH7yh6jV
RUrxVM7/ZB3QJi4jvaPZ0tQpoFYm3iQ2dq1DGDhzfPOMl4EBD+S0ch505TgIX180wpV0ZjcVzm+Z
4XrEgwe4kvjThSjXwJqFaNVPUWjXVHGk97RBrK6ytXZ9z1Q8pB2uFudX7Yzk6LODjoq7MDVHiVdu
1qsi4X9xNmryevXYTcrgZRpxTC0LntjyzlJeuzzaUGKF+8ZBy8RgjRDNSdSFiiCqIu/6seWRE8v5
bK3TrdcVWdJxLLpBFH+bUC5f+Y6uB8hGyNDiebXgIRE7QL0FMf9ibbH69RPYBmm/0bo9lLmPf/G5
qIRHrlQcbr1nE+n/piD5YlJUHT7gNwYJ6C2p2kbVU1oromZP/BT6N7p+DdIK69Glw6xSf31l5MPK
PgnWjH48VNcb3ShGUXBSF8+acCRadl3lAbSgSwi+t8ood1HCA4prZMCbYj+UfeEPb92Ke68J+KQ6
ODqlf0FLsD1hciuBGMR9t2zChQdAjYTmZ0gZv3kxHViS83swyz/Coxo1ylC4ygruQTB/taI5YXLZ
fomKMY3HvWLADg5fHoKvmLugx220x9bsodABiG/FTauASr+2lSUvHIthfDlhll/DlWWrPditolNE
Oc12gZBFTLfKQKLqzztbVpimhxWQ3ZZeeZjq+VRriOxF3jMRjPSibO+Djn2PMmXZ8ChVQRpl2iba
+iC+0pp7BPiKGu3+ctOIqlV/iB2G1hPN07ptKZToqGrTWAq01m8Ds3/ImVON6s+MQPqD4coVS0KZ
EZrBK0h7Kso1YffK/CpNVTW7voidQyaeocKoGxUsNo+ewDmRfNDXAki2OVURbApyh+CnAyKzU/mk
YUxMxoVzSLyqcY/x+Op61wdM0nlpnxOk3h6Vkqw5ClxssmvYK29Wkj8RnIWuzs+ZyegZ+0RCc5oB
V/U9v/SPQgwkSV96xJvtpi4IW2w9UOhcRnAx5RIHEiU2hBO7mjDRMqyXkt4BDU2++PfhVHRcXxeT
9jUYq1IOGZgHcgDm0D/uO9n6ebdzl3LkZMEioj+vYcjbT7jLwhOELOlhok2IaTcYtWM/W3FAIXml
6+C+urA/7cl+yAQdEwrSuuf7lkiWrFpNV/juo21XK3FUMSPJsTgAn2WwC/1tGoDFcb8OajUGcduj
hLWVhJtFwAvMiKgT6MDfncWPBsg44wC2pREDoS1K//3/9rwKg91lejtsIzGd4aS34ayzABA6vGxY
1uAgziKocXRUJySS9NGrsdQ0t5/JoJgP3niDqoDlynhdv4Fhp8jh/iDsRLByW8lrv0cG9NE+QGGR
/s34MP9vmSL7m2sEupAyXDAe9xdOr2tw2FJNZuVmU0e+Q6DXL7YKU41cfWo8DpwwfXp0zs18G5Bv
WbuCBnMsfTgKSsosi49yu7+Mf7LdmOnhMV0EZ6aj7/V6BYyvUhRa8t2AaZdRi/CVlKy54T7OYM5h
spiXgDfLkOvfkFmtg0T92Ebji28r0RsZahfSiu2jR0wKJZH/vk5u7Fd9k1zwmQ67YMGMBPJfaaud
1kTkpq1IUikB6LqfD3nBwOP0U1uQ9dEhrwz1N4NfibafTq3qGOkxhpS/PCdjy0pkFvM8oiDLA075
xCir+BS61Js6jd4o6xgsLdl5dEeMCeVpD3UpCPBqCiUIdUC1FXZarCKqPuvVGNKYj2fyOn0pHMwy
e1TQA9dYFJCxUZb1ZOabVwgZisZMEV/S3kX/uQtv6QVKIcSwLE6VqqRbtkdlvRR8pz+wAKrPnIDD
Wj31CgwHS0C6sQQHKQk0ft3+Ec9HH6h7CI4aQ/vjZ+IeAEknHOgn6XCnUlgb7XO3ADHG81wY76Qa
rXNKdsEmIGGXmmlu970RaQ503Sx6vtKFKrfG03MwS71+1ShoZMZV5fBWQF1Du/QpbVikSLhI5UkX
rqR+sVCWqqKgmpbT5us1g3gsp4Zl6T/I4l5rvIWILLk7SGiVqyDTCN3MVsXJgZckGCyowoUXVm+s
sgXWyi+k982X/c2j8dHaGSIAchZ9fgh372XZ3bVS0mAv9fMvRYy+EdxgR+xdpx3CecVz8Ij/xgjv
hb7D2hSoIniUOxjMxXKgGcNZGX55MBqO5M5iTFFSJbksTPddpGbS/HH1PnL4tkvSCzUcu1RHvGOd
kfhmO3hEUYXsdnVUR2Vo+v05srItfY8Khd/m34INv9z/Fdm0qNH2xPjCzDNc8H2f8nL/rsqML1H4
iyZlWIadestD3uEHfznCZ37QBN+Wa88f5iPcJI0SWKZpigfTM7BI8KedaO5z6sQO4nI9AIQz7rTi
pSR92dtuVfkhHXEjqQXYM/dFKfrCsiOlKBCt3aPzusa2qb1rhWA+c8ZUKd8qh1fP9LiQUimmZT15
ljl7nAcqNh8nW2zV0p2IfPQfQWmhaTxaP6/jzsEkAz+I+LIFpT4lv2XbxjDNascmjWgrEFylb4lu
Ebd+WW4DvN6RGVKbdZsXVRIMR8V10mt+jRgWCV+g7qsq0kQwumO4/cky2pxThklKNFOXAgzKKyHK
IcYqN7t9oTrmqrsqiQEdXmH+xoIq287BdM8wKdQUKmYdEI6IppYssMltsK2egy9geRNhHiMQzI7e
MvWuyXwEKQSl1xG4tcml42mTJ+m5W3xSAZ3VBmDmGjYXF3iHz/efHctkCwzthJaVRtyb1tIbRTjC
Mi8FWPU5kwTD/2NfwxP7Fv7yomWaYN/QNHbw0kKOysC5OGVXH6vkomwcqMBOZ9NZahYUA6reUUU7
h6aZDrYmxtY8jUnTlC8WmEUDPEtz0vYMnqn7bS/ReU78W3OhH45dfmDaUs4dRqxLslm26PTv8zf6
5CFuvx9O8q+SM+sifyI+OD78iefzJ0qjEvgq6Oq4ZaGDkPaT0RR+bGZ8XvpFphkTtN8YdDiAqCoP
rKm7Mmm5f228LJm4+IbeckU+OTJVmy4Cmajh1n14JLe0PGljL2i5iIRbZHUWwZ5dLFsMO8tQi+8t
82GfoUmb1S/0Yk+YirnEAkmQUVa39LbkqCxRYA65Z14rcXZOrUgbsBYUaodod5r4PLS5yygkU0Gu
czgG4WNlI3Xfx5yVseFLRptBHRUhYbTuVPUauKTu43YkLjPLGoSqMXAcHM38q+3kVbuyb44MShiU
s1v4HI/gO1BYbkw8QsEeoHDDKE/Jkz1kjWnP245uT85uY2jhMd3cTtlJ69Ty7NJy3KhFNHJ+yf6W
s2Zxfnph/6vnSjGMX9YotTdwhhZjFJeYCU8eFPf5cF749mOjagMdWU2PlbGZP8+FJNnIokwmGfEP
l08MTDBpBB8i9D1NAfto4LFNv8ZLSvTyMVx0utTqCCqRWB67b8qeqwDky3mgDgUBIVhKK0eXelEJ
CDonsexWmnxJUPO8WEBS4EGAHGfv9fti/ChWVwOdGFu6USIPEfM/Po4cD2Gq+GbUCV2hAFecbffA
FulzbrO+wcDteZnJE7Vq98exabhDK3iwXicfVNjEHij47rvNoQw4uhBgGuRiD60FDPvOFoGmhJB8
cqHYOZeGtIktmY7FmpzvF7AY5c4KFDRtH2u1RMcTMsx/FcZVgCLD12HTgwlTtsNY+Sgjks1bCzjU
mRAt+zZ2HMX3atoPxz/stxtkbIH6zGJdI5GVkX+3QQed8Pi0RmigGb96Za196WMe2d3si+wyRrWw
6gJ8s8V46ODLXNksZ4G9rL7zXszUf+j3bC/cHpwB1j0Ey0n0BMAClv/FS/aTFLpvdd/jM+JZ8UDM
x/5a4PXR/qrHP1mHB+4Opnm0gG1K5HpH60Q7ANKwPsRDnsMeB6p5mTJmaPX5dABDGmH030Zto885
vENqslRwSHGh466IRvBxTFnaiT65JPaTH2wklw7UMpyIOqrUpExoP8NiZUA+QD/rwGa60XNMBBLA
6Qc+ma151JBcbdEY9UVas03hcM2roKeH1SM2UJqaJPSu3oyO/YX4Qv2F7OjjA9k+Zb2nA2pVRpxW
y03UT8mo+qmKcZfx937nZSU9tefe51wb5x+zAn8H5WEDbJPTC2XdZqZhIi7QvYO7Dyajo9JT7Nku
ar8E6rweaZI2gbSKNZJJ253lJUwsLmxcUl0lV9SUL8XnOydZdiwQxq3rhsF/iZCxIOTwsAy1I7EV
cDvl9GWg0RRmnIb3ItyM6oc8HfqakRpw9SX/u7EMYKJn72c9gNpB/hbniW9zN90X8fqqhPe0sdJT
zhqpRb3ej1I4VvZBUcy3fVqnf7Uhmho//fUKLxX84gVC+bGDQ98tJU1EBVd3B4u3snZPpWNEIYJ0
mc2tgVwk+aH6aDex5lwZ2uZZ1tvjmYCX6Gg2tFY2gTm07eHN12ABa/2BzLlXlL6NeBulQVKKjB7Q
MutfOJfQ2AK7dyla3KC7oPjlPcdj1eUPGZjs/jEAmMygZGDB+ZWo9whUVdDSn0/Bl9JVZ14XaVgx
Q6NJ2Mv4vkLH/5gubm+X1y0u/eDcmTKeT+JA06RyLORTojt5USPPjWBmZjWzSiR2ZbG+EM2IR1LR
Kr8WXpLSV4/WKk5+UpwdmEDJINtqcWo28QpY+PGhK/bvhkx0jYQ609BFJyBs0iW66mHuGud64cIU
V+Sc8wRIkeX5WDgVUWkkGwawkvVEzb7wcmklkf5q2pDpdTCUdMmKLSCGNjD3PwddsxLsrIQxR5Sv
ZFGX2cp2IrJDz0mZ/5u2F0yBhZdD+KC/78m5wxVEcdcTh5TigYS7Y/a1racP98y+3M+iyUsRLgbd
l8KGMhrcEMjzc923Vi7LMru/7SKa6W0AZNafMPxSpyt3PTzNJH9MF4hS/PqZojR+epBK1m0Y8Si4
MCxlqFw15QSZCICj4N5htzmSl526lG3Shk5J3uebUN9MhbOUQQqDM+0KW+Nvrh7kcVed7sJhrzn+
bNgs3Y94Lri87I8s1GCk4aiHN2uFWEdI0JybpDaZ6/Ib0yn49g0dRciZmf0sBIawrV4WcXyApOGV
SlaB0My7uoABqOa/mHeVF2Q53S+qNQNWFDCyxsp49sXoqcex7fOJ/SsbHoRnptE9g5VteQPO8q8w
uWQP7IUki/Obu0NLhUOT0tTJISyzR1ypCPTHk17OzllMcAO6CAUdIcJRRqY/YMSpzeRxvF7/C0Kj
nsugIKYI+A/gayJJ8Pu1fnl9QHxsF/y2VSL52lqn6Hgcr6LLpJOTGBVYORq8uvTVT4RuO4ha176I
LLouKMglgitIVFJL6tEFPxusELMb8AzlSl4sFVqurzdEwtR6/ijJWxSJbO1qQQksAF/eVof+2aC9
uTyz/bXloTIiHfOzSZ/yxUr5p9imCdbOYwG61u4F7xc1CteaZvORfpN709l7jP/S+UqkfQBAAg2p
67Ls+APUgeC8I90Ji/u/HUkIFNtCVdcduuMEBLpUW/XkXCF/eQ0rHbSirp2Fg+yemteFKPW3bUBG
qey6qufwRTiIOn9/LoAl69RC5l4+UvU32bc1m3pCtVKyVT5Fv44xLSb/XgPeZzuXXUp19kPLYGUF
aX1/ziote7HPhIicBGs5sElP9sdQaxuCHiPeYg32bJUVrlWBflm3DiRqeFb5XXvpUkBuBl8OqUTt
yQB2XrSk9+zuZ1DsA6lXqxlbsll2Cg3C9LHEmf9YQoZER9sGkGQkKw7d8kJ3zuWJUhAKz7eGAdPW
hV0wbgwOhPBt4YTKXeNVqEGqCnFXjBSDqvuPeZVmvrpKNeDOT90izBq6ny9Ox+TAzhzVmNLeS6iS
n8A04ZKKuTDYZm0gCSuh5g1WtWyuDpz4Cn3M38k+YjnvMV2CEEuVvP1weefZigyik93iyjUCkslU
yRoh14d68AZp7+3oSFRJVJ3oOExyQDx9BkZzs57KkwgqLFCJGc2BK1nAAk6OYsFTFfrWRmPj+2wd
WQnG2NC0PWNighSNeeA33g0S37+GCD2IdleXgn6DMHtWCx/SYV2z9XOOLEXo8H9LqpgoNDjQ/nCG
E3O3c7WSC7JAkBhXiCFx2BQldT8NZfWvXV9L35Iu2s6lwi8F9q/raDkfOpvICe/46jJZ3h2xRULU
cgYKapjxWuqqH0OLcn7qx9fVHVtf6+D0tCQrrwriupKdA0udGb9f4Sgy84mZAtjSgzCMrtIsZS1P
afrxIg60mgEhfE/z21JH1Bidem94bQHEs+iTJ+lbWbQIe8PE89vYQCVu/+htFbBh1LyW4jrzuT9q
Mz8GQdY3woEYaAyTOTO6NPJOMvx3O4dBxxcMyBikkyof8GBUk5IofsM695HrA2GgSH8dhdmWWxH7
veZDfMEpB29E4qgNbZ4j/DMDsGLxaLI7Wt9/y5FZUbq5ymNPVDhFHW8H7RkSwPRlr63HyI1G4V8X
5bLeoT73Km9u/YAwtwdt/LmogyroTDfXEZ7guj4pK1TTzFIFB6UPao7Eqx/PIhUq/U5vWPWo8LzY
uTs3434oYR3nY3M8ywGXQbbHPo6cbCf+1Exs6oL5PKNMqSYPwEVtYQlwyZnamUFc8HIfSLyaDL8c
G+XXE8XCcCL4Zy9ly3dySMDj4Lq3rCr9nCBcUjsVwCWbmQNVkpPCGi6m4cRGLmFxC/P1u9uuEPQN
bKghmHYYuw4i2HhImLkI8inGLbLYVmjZ4Ryr3QGJ+de3qdOQA1SvLUF6kVfuRYbYjUrprzW5iPQL
ejDmFVZ05VHcUQw4irBwZm+3sQYu5XSZYPVNhmfuXGXM9FV01x7VDebilYXEq3Izv9jg5g4p2J3i
/DJSQjvOJ47rjsSTnlUS6Uccy5esqw+W/g/eKvQMRc0birRgbkkEp/IscZ2xL3wPAAPowQYZk9jE
B5L7sBMhEzARo2lcch6QdUqkN/s0hzRS6JZCx6jkR8Pr4q/JDlJz8XzsoKJP/dEYhX02PvN+8VNS
PqoVAn28AMG9Stab+J7Y0uXpeV9Dqkt3w+0zhY20KbeQUjtyalus+kOzR79JNqUQ7E3gwdWYoHFi
4p1LWFHO4VGwXJjc2G9DAvgUGq0XvHTYp6RVnnIShMjFXE4nxfROn41YQgT1FH4z+4IyMZx5iAsq
uIjFPp9WYx1jQGhCjnMSbvfmbdVYl2GHWVBDsu8LM2VpZTxUByodzp5gyb27Yk7wbyp84pVsD/Dd
qXEI/n9ko7qGbVBogcHBhJPwB7Ch8UyOfnDIF4Q4yF9272Vuh1+8hzyWn6OPJqKmY3ze1PlfO2EQ
Z9tJvCdCmYTXa+9tkfibXDh0HP6XtCqgPTtib2UADcT1SXDXVXwcZX6kFWxEOSah4KUL/3NifzHf
2mU5Nozqj1lMk1seu3cDLzSoaBx3h7KcOkvVGRjk/R7/l8bogGZ42SLDsneuKlxIHjuOpoV7qM2T
BHvoPO9kBV9JCjRWRTMIIWtkmE4WCJuDXztOAwx5yYBjrd1wdxoB3Gqbn/FWDBiEwuGyZS32u+bI
xpiCBsUwCKuvs3K5N/qLnFgetYCUq3V18J6Vs2fZqLKosDpSgDY22x7OjZTR/kIm3i2dWuxVQnYX
YXEq5MxIsLW/swx7I494R/mgDgKJBt4+ZWLpOjC3lbGkmLs1Ag33AKCVgawZxApReCzSwaoPZQYF
qYnw1RI0YtxQtOI82nd6awOAvbMxdtYLfKo2eVlwbrOpBO6K5RTKhNCF9C9ptMKG0mVZMsnlRzf6
rNUovQY7X5VVrgT+TW7AZxQg2eXO4VodxVzu6X5f9ElQpxEVKBALFab2fF1rJbSi4eU2aQZaIAuu
5IaQw5ehCso81PoXRaOjR5+ByPguR6ntaG2juN6fZosSdN92lOdw+ibpyjXqnunzl5hUzZsy19qe
kMlT6OCWfPp59P6IuS2+XBgzLDekq3UMZJHXm5N1pVb12JymAAufxRTCewvYhsJbSENR4ZBUJ/Fu
ffoVhiqvZ2PVfAllZWE4//WFGkKJXhjW0jtQhH6WS5kprvrLLK3rUyuxORaMinzxdICCQ6lQWdp7
LXYMII7hRHH7dP4XvCDcrUGGZylmrvNtbyvp3wyhLsAo1VXQtO/QCv5gVASBlBXGBSyjyXEOWEYc
uCrob2TRljiyczrAPWdSuHbDAi7Q/F5IgHTaveqyn2IrwDU4F9iHeMSOw0MfVUkvuyYJyoWqS8FT
PYjj87KXyQ3PxDY3EMLtI9lfSIij0JVvfeh9sPSR8r0v6ZNZ7gwAv3wLOGN9kWzmNInBUHfGNVSy
OHwx/+zo0H0cjGlStD+KssUpM8dVHDQ1Zsky1omQIKseTY08wHbHc9NwTYGoZdjEGr92oOXnuaQ3
+EmfuWGPAqFi9aVOMDuPSKm/aGD3b4W5fNTgBMRfZXPG3Vv1MNb9U26wwOoYQj50As0SyIyIUPWY
9VlvqFn/nBt1XUJl6BD5VaPJ3bMfx8/9I2sMQSrBF04JppfyShfQ/vKQR9KywCcsbrEEv1Pw+v7v
4tPCGPYutcQuYPWxYaX4LUy2dDPIX0fqByd5vs1JV+h698oYH+GqEsWJ/u0Hkjbm3tQSlk++mVEi
VF+F2kl/mLAlAOQVpzCvfHL2w1kWaBhm0zMFiiBbdGq5AGuiI9NbTggysReSAKsypz69S+5pMTK8
33kn/1eY/kP63qCuuSyI3H2B+XZ47JEm+l1MC7I5SpnFQh142UITtFG8pDA9XtkB5TkXSVvzuym4
DW/WQc7IZU0w8MrD4GzCid3LUouiLy2FjldPrpgjEQ1Yw1nEfavobZVNC6Z9Qf/+MQusMD7rWx98
GO5IwhrjrcvA34hXISdnC1Bb0K9DheKCMQaN8QYET+grpzVxVQKyEUuKloUhbY15Cym8Z2ZkfcY/
mQGHaReIFu2znYG5rNIzJUPJ6PUfp8xwrGd8BuhZ500lSWlN0Bk9fPE3yTUmfOqQZIC2EKx5vybv
oGV2t0pszNMKVMxWik8OkBilKE2LcMHVrQ8Tnuoo4ZPRsnkf8eme2mAtgk8Banb77LTTD6t1V10S
k6+oUxEJXlWnZawWw4eFtk4zomeYJPiZk3oXHabPbH/kDBqtm7Yn8FEom31C0YNEmwCvWkU+LOwc
LI86yrfis6iq4dA5y1/fuANU5Cxd2Bd3/nkumBGNW0ur9l/au37oXYMw+1r4oDc+0TeBbn9SbvnL
IqDLzDHFpRyu0cj9/NAOSCj/8LtDjM3tLzM7doXca/oS9zNrQY3YFJgcAc/H5sofZ5TImnJJOtKS
imNUJG17Y/kG9RgNXSQ5U1SjdF4EFbegkTznl4mYiT3/Zukjj12njJ3B4X4uVzAiIaAAqiJDrELj
4lDLdiMljMKAYcz36tWzN9nFczjqjGTCBSYnpxw+7wWcTTzL/XT/cMEjG3fgX9ZCFg6xEMnKq6Hl
Mj0CQ2sSqjJXZEENGKqGOLdhBxMtsGYouWo27dcaoGNFIPhOajtU0rn2PHfH91jGHfdQktyxlnKq
2UC8uJnKXnJYXsupWkKw0ZuGLRM4X/Kg2YRy9G1aS4QP+XCobGA5VzEX/O0fsLqRUtnDW9zs3ai6
yDUUWmUX5dApQITmWNTP8prRWWt93Xc8DOSSlZt5UAZPs4yksiJ3gfn7wvZsDxdJOMFl8TqOUm7n
KgQCjVTtPCwpeI2SSm7Xz5Q2FVD1OB/zl/8ryOYqc36LxldfdEtnPQfVK29upCgbkev32V/Cpz1w
xnSw47EIvgDittQX2pHPepg/Ig09zrj0bfQnlfF/WaNOYb/ObMgkyfK1j0TGdYoHXMLpzJeElpFz
VH3ZrixklcDT5CjLzZ/nqvMg9KZYNn+1TBDxvv6yvaK0qDbHmG5Ci7m4ulfODp1CD32NYne+0N2O
s8rPAAW4YMRcUpSwKczxPW0OD7CS0ZKXGfxUrCA7BbPSjIGEo9ZpLiwQdnjo8kEpda/AFks38Nnj
ihR679F0nrbl3SrzGnRioXq2WWp6een0RhijHhYKU3lSiSnrDdRxTI8GmDylNNX0F+hvfwKZE3kR
4ueql3aAxWFsvF/se0y8uKwknvJVq/YLnKJmzJGgXJ4Slgu127fs+6qBIPZAD4NooDC0tDmwquWM
IDTPWar+9OQlHfTTwmgIRj2yWAxR7JMoovLnxtWkQ7rPVuk3TvxwupbQicdpEDwn/hF95GyTQV7W
sWv68O6x1ftrJ9O9SeziG/7GPXbhy0XukuAIle7xZIMwIglidweK8tTDSbHidICD1DBmA0eoyfyN
5KAHFEBuyTiTESaHIqE5tLtS8sfMdl099lfLMcYCZd74Q6i+VD6BnpM7U4DVEjmBF608Dq4qTO9G
orljaBS+YKR3g1cCQRZD3I5bCv0wdstR+vsFEBYZl5QF54PMlPf6x+ccPZ4dETb1cRrpx/XJzn7s
9uUc2SJvx5GE7pfaHm0EpjG+ite8CXRpAuH2iPsE2ynGQBKYBoWKKFkwwcBbaexS9EGg4tka4JLl
ykMNWT7aOdSMTjGNxpW9DSghXJGINnrG01rDx8V222beyhNfDG57sj+trjalPJ/rK8o1I+H1jFO3
s++QIjoOCvMRPgvKMZihUADxUKiHdeMSIu0/LROPDEk7pqQk7HT5FpLcDMhV8TJEcz/0qE237UwH
amIajRxwJZbQ/Ws7sq2BFms5B8LrrYiq9gwTVfsuSsDhLnwfA3wSTv1rFjXe9Z8K6AhYt7HaxKZV
KffDzWW+RM6mCqMc5VA1YpT2en7Fs/4EuQCA6iXyC+IKB5RprKh/cEG7CJL4ltpNlg0vN6LYf/2N
3tzWZJs9zwjSTswE9IwtLYfpWBMNuG7wEFwxgjBfg1TAzznIEXSvA5fARMBzI9qcW9FF3NJVJ+FS
U96bZbJtOw8I+KPh3BIStGPNg4AxxpztuhCpp1Y9AKQZVusSTH8KdEKW7uRX2SIrahK+U9fTQO9J
csd+yn3NG8kkTWEnyEWDJlDOjW0DzE/rLKu+E+BO1S0BC49NiR3vWkqmBnNp2RkCZkFmNE11RXQR
sHIz1ukmGUyEj4WradYLdqu7cazdO9e6YLT+77/vlyq2PVcwj+MkT+vLEG8u29aKE6JKiuSDE+Iy
MO2n6AbvrImPl05OoMmw2Wo1R3lJSF69iKKBQ0q4NzxhyGTDU7OvrRfwRi/+bW/P2wdmGjib2vqY
HIJvCt2RltbKaCZNhydpwxUhzPO3jfw3NwdF0jxBVH1sZJSOjXNRfb0OFAIY/g3xa5oEth6mG18G
hQ80vJnH+YwM6/USC3o7XIrIPZyF2T/SnZL1sxdhx1ioRtsZdXtpYLyOT99/mmisMn09amwUMuJP
IaaQuD8VRSyTD4qHBt32qEENPQDJpBUqNc33BlUBddT9/nkYKYB8qPb454EUhjZ9HCd05stEG5Fb
sFDIv/1xfI8uxj2CTpndvSJZe246MibptxhIE+RnifdzpzTSVz4Er3E8Iofaz8UjCvIeRUB4u+yf
AwzWt4kxIxsAqTol+dIu7Z2INEhtGmXEGk9kKwGlm4VRdny9prP8JNgQfb8DT8VklwM7nhLO5MyF
ynQJhUg43A3/9o7zs1BTqxhxwV0KsAf6U/DqDSlPWZBNpkqyxTW7JZ6kTBqboA+YrNEbr1vT6I+T
VRMu/NYQO0RwTi7Rj4SzjCZ/XfsZSbYA4iqmlHwPB7h+nAaT3Fm/rXpFZs739HA6sYmcjB28m5vG
YegX10ReYRIUH8pbv/nL5DknthZy7tc2MSwRiAOdYlZrEZ9JY7ldyVdOw/OK+jC95rZIyi2y5N+q
ZImDaNFasUvj9IN38P6YikVARBxCPRdjQ2q7ZCAeplOELDOBI0jcxlx/j+BIIOaOAlPQ0I+xx3ef
8rGHzXkJ8lLEShniLIVJqmIvSnTvm0pSPPisFdtod/yKd3AVkSqmyQAWXCiTnMlRhDhAy/FOPLW3
TNk7bzSBjBS1TkYBaUgtTh9fTxo382/SPOJ87UdeTENRg0mnsPGpLl/jWXMQezsRGcNTNPmWh8Nz
rj253UC1GXRw4CmAM+oHZkowIAKo1qhwXCE7WRLeZtLWq6tJ1tjMDmjDVijDvn/dSZumJHmbiQYC
pRr9rD9mMGODW4yIAtovxCfsKfivuy5WVQmHSn43aexFcKSyfoIPi28pjupufNIDWnNAHMPiHkNO
EpFMJ3ZoTh6g0gwQM0nz6891HafeaxK06dKx3ROPWHTOx8r3NSyVx5mk2K1dEEMdI7sAuqFXw05O
Hg/q5LpFQCwweAP7cl3WGlT4JKJYksjqLuISMeIP08GibdKZFEMyU5s1T1i3fypJT1jOMlOZ6GgB
h1Ues+M41yYCxePFFdTwv1ebVEzqLem2sVoeIrd8oDxcPGLpqVhD4tC5ix5hdpfSjVSSZdNvPwFQ
X9WfkCV6CRgXtkvDlhU+lugVNVxxSkgmXDPLfWGW0nAl/nyaCJkEUQykK7SVtVpVQh/HG4Egc7xa
pMp5I1dsT3NqWSeQpWIqHBj9zusP6dIMBzpEMcngUZkUBychgi7W17XKC2MoM12bMAAzHXuN7xB5
i+v6XQLWxUoKZRTeJE0QAzZugI34BzMECVfAvpEsuPKvKGMRmG7i2DZDMmTCxZg1AjfDdPn3sRGg
v8KbD2IyNp5HyTuuiU++N0osMSL61kMieg5IaPYpihKEqYdSmEeAoVQroj1VMzCXkybq93zkbIOX
ORL749dT9ct1v+NZEnnisEl/adN57QzxgEvXuta1ssTrvBIk8pUpgMQ778qbLoxQOqrim6UnBU8k
TnVWdgjlZ+p1++PJexEKOyrRWAHYhVgAE/MxIdHz3sFIOgAyx9pdfp5pptop1PyEWdRYoZHkf9Rh
r2z8dYu7EP0W7SHaFGJ1tbaCrWgg8u9zLSLVeJpzv3A090JfYWtW/MoXAIzoou8Y/bnW5tC+DEY1
mALCnf0c9jMaL6RxJbYw2NPanyfCn26zt5SOHy8YnkOB8xyAyhPhygJ+fyAmdpKlB/g7/1Ck2QXw
wcnL7DuTNZRB0xjJASh1ylzbTUW9EbV1n4JTDd0MqsGpu0zuPDhD1AjVHZtiSyGt9eUpNlTV0MHh
tbMDfdx06KVbfJMPAe6pS7lKqXzukmmxjMS0d/SFcEG3wsuUnhHZm1s6obmHg5x8y+WcyxVlJBeA
pHnZ/uzOYYiyVFc4yEZXOpUBzGuOn7iocwa2muUuxP2KB2wQ+TU45c4paCBncV57V+vw+vulKmHs
H+5UGnipdXQLg5PU90zrqKvu3Qty6MaseU9h8sXwIwToLmwy9aiGtkDzoNZvbBj4Am0pslDPRvHn
EQfhyKZovGydkIjJ8OzxES9DN5x3LM4ME+zO4fFzdM3z/A3Z/BzJmi227UQccvzZAc4jLMwk8awu
0WFRygcCxtzB2DvDOGmi/0yff6MJSC9cy/jju7yUosz8NyW+JaOVBtg+7V0NAn2LJlqUzj8LKY6p
R005qIOrunFApu913yt48XOXF4dXW8OOv/fwmnT1DqsGWIjlea6T9NynN62Y2rxvt4hT3nNFFgSg
wZHJ/CUpQuc+wun+FVaiUljhL0rlCiwLbumtzDsfF9YEvGTF90AhQW3uQJoOkU91O1BRS1ivXN3w
V9+tbeZw8uUvRNWRXElqBtPRcA0HRx12zBWK81K49fz0mOA9sN0NByUtGKbUc9hrEAdV8EG3zI6U
41OHyYbTz3XxRJUrHng2WM+PbgGSdBnzPxoLVOERNZDfUFs6RVrvsaVKlCLmM0Aa+dPGtBlmjAiz
nuiu607upoKT4ldwbcha+782Gtc8/cnyFI4VFC94ElrRMIMti5k8t6/y3v0NPejnzP5k8/fO/lyv
WYN04laLV7JhpZ09C2ZWDjLYTZi9iVmZogXNiH9lV7p3+vLD+56J9lAsfR2RrP5AtJX5BvgKLL4J
SYy4st5XH1sPtryP/3AK95w2aBzZcaTbfmcoFEbpAQP0MxV1MRJw/ArCHC2pPAWGBVYelqO97hLa
tYN3lKt6H9Abkbhj0KWoDmo9xLTP2l6eIM64JEA9+c/SIaF1SAJmDiyZQuUHOEXekBFIUG7t72D8
tuiZCdE0KRZf5IisIMQm7t4VeuXTr6SGn7HtAbY6OOZI1heWE5SrHV8jfYDK6j+QDU0NxhIn3nGC
aykFlmahZOyHdHbhs8X0JxEKcgA9Zj9ZmmoK3VhOUAakFOvRMtOL6oY5tQsRcNRA4M8D9jQCgGnD
S/2d6DIS8OxT0GtZRt5Zu/0LrJoPX+5STKL6UMMF41ipqKge+rXvTCupWXVuXJL0MMsAgyaVwIFM
oz4Pf6aKd8nBVF6Cs6SWgTzrCG6mvkybTmGYhgMQfKWNLnnAHQrr1/z1BDtkndY/7OvaXlKh+MPT
IWhb37DzvvHsAxaxGmXsnyGiRH4rbjfUf07HNBVDlrs4BzHKnBgtvauTRtbndEHZ+2LVMtWGa+1D
HpSfXLvnn8hOM5S9PONHRl4Rg7IJWWmIyOHVm2KEVercUJahXJN+jjzEN8EwCF6TvuojB94564NB
d3xxtzCdkFCSIxP099PuZ6u3l/ys6mMIg+NuLg/epIUY5WpCEi2vs7NWNIHvybhY6txJSKeKgXzw
lBDFKpK8vj44hmbBfVL5VP3kOBr7GMcCLxwp/fpGesTPb9jiGlp31u+NZx4kC3o0quxjYoa/+4Ok
SeBZJ5Lfr3ms9E0GhxflxZpXRTQ1/ApkJFbecyWTLHyVhOBEDfJ1Jp8gXiFHPEpnDImuKfrgr3dK
nPUxi9vnvNNnB363P8QbTifyanLjTElDLrOEqmHLIhRfC9xa+rr2M10o8E6JtQqRVXmgBTRi5EOi
tEcTD5T+QDserX2Ms/dzdr3xOA5VySUUDueg1pobxEAj841MpaIt/QQolcW/jqyFMaR4tz1XaG47
Y9+XQAPRI/8ZV1d+uU13bXtZYKtQX97Ld/r4f5lOBRg7UgUpKDQO4pNAABmxSDSDSfmn9wAvq2se
5xHNeZgDzSaP+e7z5hKfbzYINixpmTY/cZeioJyJMSm65qL6zKGq0y9WXSl0v0YYqiGCtWzLPX+j
HvyaLAxF6TnESXSZu+CINAXSzUZhPHiQ5Vtri15X88k0lYAXIzIxNQ9F5SoYz59VAG78zeufuvnV
ju0hCtW3GyAtipdBKtToDyHdHgxLF4IoocZRowm4lqpgg4f024cxPFIBR5d6ViFRuZ0s4lgu9lyX
3iqKHE9l6vMHKVxojyjpjedbXfsMHBvU4Ug6Yb8HAkZIXwiI4jwv7otSWKezLLjEOmaQSXwanaHw
orKK3DrbKVffuF38C/5A2auK8Zahs122cMGWIUfkajW3niQEThp0v5IuU6bAFh8vVP8tZlXzT364
XRaDukOZXWmkjK/wwbX/CWt31bZ2A0/iQcT+1dhGnHctte/1ytuHFr0/4QXZMn/5GEcxjr6GDd8T
eu2GwA8fRC7XTxW/kIuel3ZYpK124o04GvrD7T2AQ+jbjDb7fXSFiio0GQaBwbcGDHt1ygfUYB1j
CbAj34JT4A69yKHx5zD1gSH6dUOL8yyirNvgi4ZlKwfnbbTglUocIlD8WK1cGt5lfpx8QBCVy9Wk
ADKNnFIgr2fzSWZmxquA4q/+UBZ4s8gE5CtdSYGP1m5wfbOXn18M/pDbtR/0i0vYMG7moM62gpUM
QuJ1pWzppAsAFbMn5ifjT0Nvv6zZfCjfiVaHDLtjTNizpAgNYuzs2Gonkv0WuOq8B/ED5VbgvRor
pucMiOE9lXdLlSX8JRjqmdqw/993snd8S4UPLSYH+MwLAt+6yIZcMA5hkHMghYHn0z3TeYsSRKZr
NmUNrE0hG6NNGHfWqlCl1bE0Fbxe8HJoWneZepwG6kdRFKJ0SU3QUk9bMEc643lWPPkURKBJCHOr
E9i3Ow75MdOiJnLmMgU7iNMwRwMhPSZK5T6IDs0ofvzQdjfVQMZi2nlAs3ZBREl+V0jrhWuuvbaO
3C6+iYZXunFopo19w3oHlDgyRrd1Fn0VdNKVbwGmn88AFwIPOXXAfbRdNNvJhBvKo0KbmU7DqsBL
IUO4pT/SvB53ujbiLFulZoYedQauVzHFT3anmbDK33BzgIzARoH0+nkvHXrzwMctZpIdAlIxunQR
OhDTGbgtxO4eqQ5swkGdGCrdndKlDVV9ibySpeOdd/n3ASEftqI+3wRn758S9MJyW9LloU8Tf4GU
tp/8r6xfJdu8eUZyYQZK8attsXGcDaR/FYQotNzbH6jXa7gvZICPtg8m/dUFHjma9Ji25wbCJTV/
HjYaZv6QyWjKXlbIxQ9ieXDC9ToX25xPm50UW6IwFkUQK5OMDTy9Py/G7J/RD7irAWL387sCOlR9
djFSNmdxppPC3yJ2LR+h5v+XQ6cfSFE3pEEQHCq+ZrSvpNdrii4+o9/J5/7/1zmWgKA3pwKAsCUa
M1TOE3T1pXv0tFMISSp7zyUDYbvFlUdlRqKeMGUjquWVZ3ATTU6mB9v7EOl5Il8GLWyJjKOZ5UvL
UBxW69L9GHVcrETdXPdMJm/txXi7l7VKFSguArP3ISAVflNDNYUGQzFFQOcf4PVOU2cbqnS1NbF8
5UbKptigG/hlq+/6JofwgasfYkuytd3L3zdOSNjWyNRxGLdjAPaygEByN9f6fImcT5s7nccem3Dn
N1iKwL7Jcjesan76qU42xpKoOR/n+FVTrYAtXm0RTDZ5pYSevZkrAxmhETA176hmp6V2tCa2+4Tf
C3zM3I3iyuL2Mfvu12xSzlBBnRPvSG6f1tmRST2OBWYyILb97BVkJS2NS2efZv4wG59ID+G0/vqq
uwTZ9iluXWBV3EG0vtDh+pTN5Dd/g9IK1PlxXlcso2AOdWU8v9JB4vgqqIWTwoepk7kk7hGw83hl
IWRfUIEf4DHTGxmiTvmccSbdQHrS2cYQ1/TexX51BRj2AUQFCi0vmmsaiVfZLxSn/S1iIZjwayKX
U+zO4v48LKbHp90fFG7wyT/iVdAfu1RfoNDsy3NACMKfCoTXhG4rv+K6SZhu5SmX0l74I2NM3qxR
CuJ1rfyCuFh+v6xEuzMjcdB7ZdVTn2yK8suOBgZJBfX9aGcZLHVBPKEe+F2t+LFi2UdnASi0aj8G
n3emnbAE0EDAykawxFfBwlY5wqXK3GHuSRC3vD9jELc1PpknP84+PtkavvKcawvso1CypB4FHcwF
dLeOssx/D5yHyNiCazeIDKauKHd/q3Y1RsuGz6VuxP/EnvoTPs9phIAXKe7z1ar24VBDssZ2Ml16
ARHeuywpK+Pakekm1oIzLO3E+nySX0fRhfSn9HWrX/x6dVfDbfM3hkgUkot/mvzg+ouPywPWlTo0
M/B3FM8QUBME0kRtZIwQuTsxxCLU4RmFxYlMYvaDAd2tMB2tSZE+1JXtszqqEtecFjDLNvr3FKO9
JCBPymiTWKHM86rxbXdNeMtAlJ3mlpa9idyA6FoDMzJjFh1dy0c/bLvUFaBueNBSjFVu2zSGCpu/
9XRVUyNQ7T8Jo94bgfgFrKVayl2oPw/anxjxdN27dJBLWlq7zVUbaOjel+OHKpHGhcxu1EzS9eU+
ubI7YxB+ZJFZ4VBTMMXHF8uMCIUMgy8Tku+0L/uEkeARFGMiG2qbMXBEdBsAXoXNF3935wcQLe8w
sPrLy3EV4crH3qwIiaNEkf8Q3Qh+rx5nki9kCknCtBlouOoOywdw7jQ8/QdIM2jA5FAdRrJQIuUF
xdktQ/vqUimYgjGe3Zu4MlDVOxalqQRWRZIXz9b0rROPiRZXEsRXnjqb+87LoiLa5ZOcMUB7zKvr
1lPKVZ4GoDFGKrWtKUMSTuxxqS/Y+GDcW3tAiW4IHDLqZZwgK27BedpS5Z6WAJhMbJHhIxJgYB5w
V71Wkmjl2u67u845AIsKEHZWhpceUJQ3CMz9bfDiEYSf2Qem9WvPUFdsCgMK47dYhmoTmhu3pJFa
Ehvmrt5pxjaiACKpeGm2bb1XbfxnfnnEQ0bIMjeYwvNfsH0FnwUugZaStoM52Vw702ajrVimEspx
1U4L8b+g4P/1/l+57fMyHmk+GLOhnz8z3I1hzBiJbSlgqFG7PUQ3jjdtHFKeEGfyDlFIhCQgSEEQ
EZbzlMYePD+tY42NseaFDSZtxGOSsGa3DcwKaiqlvxVMsmO22Sz0QfU1y79uPgL2J/j/K7M8rr1y
riXqq88KvxVWbJKgq/N3JASFkCjS5yrmv9/vunDJBXcUuGwLX3LcLFbNb0Lhbz7FO+Ai0lVkKD2I
qzKyUFAuEFxVg872RwKUr5Bf3XJqpnzeI6tKcZ5b6fwBMvGqI1XWsljqhrY94Je9l2BudRuEfv/y
zJVzG2rGGuYYWYXkyIFPROS/i1l8FFd3LGP2ODLyuBgxvraADP45VD9wYVtfLOCxP39/GDiB/JNc
/pr2UJYZky4AZO/OeBpZm18YaAfJ4PNcI4ZBDf/yEtwPfU1kk0csfXpQGygoqchg4qUs4A1nJzcy
fSjJ/OCaVgzvqIRB4oyWDoyzHT638ToUpMT+CqHmjGenYaunvqm95afAazrmNSbUoer+nPRGznpm
PVaZrOG8GvcApzrA00ecVwvkqUFgh4Tf8fhl3pYG1gtl+YOPj2NqpTuFnVWlEOIz37E4cG52iWFp
RM3XBjj88yA2/o+n6icZ6zS038ZvOxq9o3eCeDA1UbSfLRdfn8SjCsM4UpqB+tEInEZCxHduv4h5
VOVpGcwqt716YCSOuUkRy4d0bLan7udwPJtM80yua8BGugVMzttm6ZR40Hrvz7K9Q+Ql61p0JfAR
0kDlCYOfEnZG4SL0K1anbcRbc4R9TnQRgj923hE5bRNA7iRcGRlc1Sl9LK2dnk/dS6TSJjTdC++o
lJ+ntyRhgPqw4CXDRDBdK5P4rWyDE0moor90E35Y+F3HQhVMFvsVyTZJ51wt5HpXOkcfV6zEGXQj
+KDveQUz/Yz49+/LLRtFvqrWJMqw57j+JaWSXmSepCMkmdAvlXCv6fodLjEe8i+J2zyP9Gsee6vm
ykuF+dAdpjo2Q0HnLDli6ZFyceUlG9WL/hIdpP6BFqOpowhg/nYwFF0+sRg0njfWv1cZfEjgUQWG
WFjcj9KfgFPMUWaDVDXWoYalcivC14XIULPWYQ8CMV7EAxJ7nbW5ZheWhCRQULtcEzTKTQ573ryZ
nOvNVurD8/6Zv7jitnjrNbONFaYiFrHpCeTTmouZAnkEQ4wxDEM35o6r3tGFm00E7vkms5oPLZCH
PqqGUDAip0N7A6R+LQ0hNziZ8zGOBLgCw/W5EPTGB73lwkIuaaIC26d20acusgzbfw3qc3aCSM3G
HKBGLGwKWvFY4eI3GF8WjcRkN064+FTIfTCdYD27FRZ/3B8b/FsUldobYWNQ/AYhmFq+IJb62H/h
zTne+oR2aytQtuBT2SZxlYYHHyVznysrqJLRndYMSn7EJ1orJB0p8fDut9SsXOKnji9KVPnDFhEG
SNyFNJ+QfGT0TGFXYZ2AxLug3b1PkXYaHGjHbGqVU2AgoDauN4E58pP2XpItGnfyyJhXDWI7eloq
hCwFs0F4MzxLps0cy803EfWOC1Nq7UvVEq1eg9afAS6wXSbdw7urgcbnfx+WJ30Y613ypfBZHrGx
f2bz0LRB0GC0EMCtr0EM7UBYyQtKNtq3mfbCZzvtj07Pfjw8Ep7bhGt1DXX3KHls4qB+/IZ4pvzw
Nbi1M/yW3MQJCv+NbOsuo6cYf6Is4UWbVls39bK6BwGYlp3vV1TA8jDLY+68vS9l8epl2+5QBTXE
6+fA9AlFuVjMYAuMoZnjHZ3081Pc1QNXvtrd/jc267PimcZhHYVSNMo68q0qeZAVuSMiEzpD+BW9
gYADfUs2obrpQlnV9kQ+g2YvGDieNx1LTHdRY7NCTFsMQddK4uG6XcbLskBTCLpUPEPEuG5D0B0l
NZbiVbPGJEoE/LW8EpgSZaZ6SKytPy0SyQystnXvrb4dcajLt29RPWwJAC4N/6zQvmgw4aGtVRbe
btDzjuIXDVodnvUiiguBZCbiGcyfrm59Pf4aHPJSMbYU/Cw5BClJmQYjkqHYGZfFAofD4XbRfGia
Ir7bRG4nUGnGPrD9oLN4ObSz/Un8LZi91Eg3F7ZhCP0FOP3uRSi1e6qeHcwUmeaDSLWRy+Ch1Svn
W1dUis4J57E4EnotbuziCQHjLWphvo+y0KubqTrl04nTNoyqAtOVj/Wz3WFqZMJ34Dy0w9nnU92Z
ETPFe/IrHyP0XjcWEmi3zJy7aHBgH0pPK0g3r3MgJ5HLIAaw02HbBbatxbmvD/zdVYyN54M7/Nhd
ebUvsEXFq/nBsF7x3iGF8cojpt1hl9YdTD8dRYefzbv5tFcIJlLdbMftCSWB207/leLdGMQMQVGn
VQWB1H693M8U6yK/gg8jCmNT2bIsXKF07XL4Q6K/ow/kndU8VMk/vdJ7N+j8j6Kx0rbuaLdW4AP+
3FFAXMq5qPYKbdo36Ni8lxKMIlwnlkFVe2WCUc+7u/fvIUwNV5OnfSZysXmr7RjekJ2UiSqWgqqC
XlnoVYXdeykKU8VY4oPBEItHpPIa2Jun9QGIGTV+h8+P1bGEtjo/zMKDx6k8626J8v84y5VwnWVM
G9RffqM9pP6Qui0CJHuiOwtTdujvuzygFdfsPHlTHQ3zBO/aY40MxQe11c5uxeBD78fH3UUUnToj
U6AoolZU2aJ0kZMfb9lvr08foG4ww4Rqrt8cJM3s2T0jtE/Y658JpXhE9iWCwJVM+IEN1ba0/BiJ
eMQFIvhHcVbI20jkkMP4fl5sfLubMwiwOKmDW25BKqL1ten1PpQPads4X8/TNb4yvQGrd6ee2OCI
2Wp0RYXbp3kwHGahJTd7E2Y5OXvP8NnA+gFGJS6LQUYDnK0lus2Jr0l3JaIMUWbmVH9bM/PeQh21
lS+4Jd/Okjpyu5yQEHiRnwdT0kbAexawQHm0qdv1jQnZC0BCS3JBJidHz6LGPJ6BvGzDAdm5vCh7
tahASCVVy3WeaGCe9BUl/92V2nNyhr2TEQ5kGSCs833tRnVlWCJ1whT9b5lT4rTX39xp2pE5gjpl
GVUp7kHmXkg6KJACQQVTM76kGEh9s9vTMEP4IXH5nF7OPxjs5A1wjmW60oA2g0KE1+ez+QS3c4li
JDo1C6Gjp58kQM8kHwLO6peqhkdWfKHqpSDiNycUVALhYIGtOMvlgV1p8PRzTKcK1wA/lAQ1LTLV
zvaQ7qAlCGZvME/G4WYrXD40mjmHymylPD+iSL3hkLKA5Ex5BkUoY5GTxihVrdqgx3zZMQrs2j1C
WtSkkF/pd9JTZOxIT/MBraXougEnAVJ7XDznt4wu9AhmEoHDdYltnt3UONXKJGQdeYPEvDdEGhXE
2Y3WuDekUeHWvKDy9/Ica+Yoph5oP4VfUaQV6TrFKZJZA/hnUqj4vcoZl622Fmca96aRttcVBE33
deZ4+ChmrkyQ1Q5hDTG8XBzRKGLjqjW3WJndc1BDxuSa3vdJpE4Jg4o/jFra5xKeJ/EYwZT/vh1N
+miwX9jPt8lPJpKZhHBGlhJ0nKf6XAEdLO/cfjQA4EACePunIwA6G56+68gNC8YBda88DiE4lhDU
+pabJClvG16wTa74R6+sGuL4LWdVtzBCCYmcnMhJzt/j773ALFDFMRbc5oHwj4N9pwxiCkj1gqqL
eYJ4nkNGMEe6WwMowOjXuwkTiJuCzDHGlDOeZsF/p3FA6UK582j0PMa/NHHzbihb1ph15ki+JNIo
MDbEA1KBmPMkUrf/W8/xRU3ZkrxePA6YP7snOc9cdbVY1GnIUNGV+N7QvsUFDO4OK3hAv4jXI9ex
4+xQtZazVGewl/dCNnSMxQ+zEy/Cb29IvBcAXbGx299BVD6on+/5bdCQDfjs0Oi/OOtaWiTysO1c
cNydwH9RrdIbtbbSu86rWJO6OqBanZ11aC0ZoRoeMWXQAU9GuGj78uzsNTIMQKzR4Z3fTHKuYrz9
VWD5PM2V7Z81WZDDV2gHP8C3YYsAUWcgvImTcBO1UIZZZA8171Km8ZKcEFBvZrtglH3xDXieStXZ
jbvUGzrQmA2GlByqkvdcasW4xGY1OExWB3l36Y/7aE214+3V2kbsND1wQ+UhjfgFqAPJuj/yGytH
Fiv75VxzFmjd4jYNgybv6Vwex9yP0sKiXttqeZKg/tMMFI16VWSmjPULF+aF3my0tT5ekONW/d9K
fMng/AWGPeju6fzx61XPm4T3IHbTAW7FGO5bwZVyQAun1L0cqoPkHx275Pk9gkc/T2ZNO3xjXWWe
HXgY9Y54jR+b2mJGSZGSZevC+qXBbhMUlHlJqSR7ia1IOinR3Y7y0qISC43l9kkZoGkUCOih4/S3
NvS2Sx1XI2jC3aKAy2Kr2s8zh8wLUVs0M0uUAUaTuzVcosO7PsNFlYL0HSocyl0zcoINiXgOLxZd
CAdpluWdEgIDs3/mgANi0LvQQaxZWBcXd/g6KpZVX4wNLbg/BV0oQFpM0BpfB9G6nHhcSGo8Zn4e
fRfL38NvwecL/YQ2UbKuXC6FnAiuXSH7WX+A55ISaaXTozoB99FooMTGFH7VA8kz86RNi3+HmnHS
pR/U6cc3YP1H8zj522qNTxcT8slS9HuhGqAuSa4ek4PuhU0dPpmH4Z19+6hsTfIeEb7m9wHmjC0l
NA/lEUZirDSHV+nTjIpk0lMQ20V0XsoDRs+/vG0pEij6BZgqjCYGqfyMMnm/5Wf/+tLBLu/clroL
pzz43Gp9JheO6W2eeY17zLfUp+k9ZSZct/O/hJy6ECSMHUB4aw7WlsV0O9T+DnUO3PXrwxt5/i3U
k2M8NU4cnHxhjgyBx6lB4+5AUlQdTXjx9r+4GBgfzqkPy1XM8ZjkgFwyjG1F2TKnmVEZ+9C+jEZx
TaNukpnrbL+cILfhVhV9/pNtU/A8KMa1hvMxlmObTVqA25uDGyQL1KbnVN0aPRstaQt9LY/Fl2BO
D0GE3uPzzgBP5xPFpm039J2aTc0MP4x3wRxWeENf7UqNBNDj9rcQFbr0ty4mUaM8TUB3soe4jxax
dW72ZTqrbgxsslQ3YGjC+fuSuPyJrOeP08oV2r379CGizQHwBAo2uvzoSXJuDenjQ5LlBx524o9E
NEUEqDUrhltG+WKSZI4QBl+9zYOxU8/HqgZhP4U8QKukL8gDxYYOI5NmpLnu5oebX2w9ssoaHT+9
huUyoaaFI7c6OPbia/cxfvQpYaSK+uXoASbnssys2cBt5/i070LpjcbLzi4COdcoKtEey4stbr82
NUs3+8QRECLIx7uxwpzpszVJydFr7Ge0lG86KOK99wIMf2mShBS8o3jG8p3fbHceNEqlWQKVf36C
MQ0VXQlBhAS14ksc08MquM/ibunnFAYbp4xmgz0p+gVLInCrJKieSgkSmYZoXBeAGXJVxBqzdBNA
HnabdEtxWto5Jq7Q/O4gufaIcvPPEDLg0sVJA14boa3hqQR/JYkniqmNnOZ4H/7lAicJ+0vD5dmU
4DKEVZpHU3mcLNrVDuZyG1+sy79Q7u6h/xpBicsAIqWoxzuuAfqm1VExTggSgLxVBx0nlQhQo/b5
898g9oU87/PAErxp4qXhY+/EOqob391qTOxx3ti6cdiy+dBJeA+YihY/0j1Jhvupp4dzb1g86Fxl
L21zQtm3eH6SZxKjV2indzttHzkRhWul90HFYOEzt4IFY9VVKFY7JqGFZUslePxRN6aw/R1E0E/n
qFgEoBxvrOxDgayOOU8PF131IUnt/6Sdp+qt+QVRT9MtOUGIQ0byM/AEZb7dda1UB6Bc3OG+stGt
ATSCig/x+3CO0+pt+8JX7oSE5LVRek5Ne9Z8kSkPRVETT+SzyAgXV1dh5NRajoRl/Yv3b+37IYO8
woxtoZNAwcRcLx8Wcq7ArIqO3mRa5cUFhevbLSV+6Zlc6C+LxhmN6TOiGbT00HSTBkqYmMaO9e14
6fuO37Hyub6TJ837iHrnjYpRzv3ttw3zdgMbhhM79kTab6aqQ06U8lIUW5rW6K2XqxaUYRVLkegT
JCaIgJXCx8/XGW3upXQ12nc8DNhd1ZY+SifNFtLcLI4uFAW+4OJ0VM00dQm9ASqGci7FsfT23rym
EztftH3uBbPJ+tNYpdKdU3px+gETsvwpkUa205AUJwSh8TDuzK9QKOiIoSfca52notu2YrIRroS9
9ncj3LEz9VEm+RWQdQzrtn9KUPdh4lXSi6REIaGswepPOgxa7qblsu7lqVqe2JjnjRL9rO0tm6GG
8DEVtUVW8PImVshGD1ktDbdtScMsrpjBpXaxjWY2QZQOhVef9hvKHYDfFFuAe+WvLhjtPG/98U7v
Oxt3atvSmBVMzGgt/YryPIsOIpASUIXZQlYtl2ZSGlal05J535RqcTGF4w48MoQLkbXUS7S9/Bit
OmLHrWGN1YB6W2TKXgKVSN7IFSxUqhhSawbtkIA6b/ORZHkkgHqQuYuBnIv4SBycFijSbRk3Qv0c
cG8baueZBRMq9NNCfKU04eGmy4hwyKGWG2yMcvrJxlzeIpAK/CjA9VAqdLgs6gAyVVe9sh+w0Rzk
EU40VBErorWn1QVBgYvdI9/oKPqu43tsbg+IuS7ZaI4g6YK+W3CF/CkHyJoiso9VaENJj6ZB1LKZ
3Cxdbv9GDpsJ7H/a0+gszSqeYHkk3zYdWPEpI/35STPxkdbMcpmCg/l/8R/WWc4KVlSuspuIZ0UO
SoQlAMFZS43iVIM8K7rMVpCCne7UV5aumd/ahxrS0/bINY9vjw70FcwEP34JrGZ3INiCp719qoZG
w/FSPsRk8+4fWI0yhMgnNha5R2dxIKXkHmiwqt++MAgqFxMRl2WJyYdtwnMc5gE9KCwtm3R2HCg8
RQND5993GVXQTDAFXlngYQlscvLlNwvzSJuEpl+YqwsWH1gC9TroL19kFFQpUwIwkfFQcPExRbqM
RFsGEBO3S5vXl0jlR0UoPxuTn/OQtIXtXlahlFWQGdTQI4EVtCpe9Znun3qTj0ITGZ0r33UaFPdV
T+kfGO+azrGCk7v/a/Ki0ljP2RApG9NwG8A2AASiVZr/NrBT7Zdwj+AcHZOcWLUMJFMomAzfpy8q
bFsS3Gd8Gt3/4EjVsP3Xf/KXhxUmk2I7jXzA3d7shdZgryNw13ZJ9ovG+skGxIxh6oiYzCyiGFPI
apltb+cWwGolTRn94iRFlo6Vz+1c6NuEQdY+XXV9otVTju/YQtOqWtt+QTvOZwqCPn+yoGyJHA3y
xPlTVNhUQzGvUfEZ33hXK8R+le6S848GEuLe0yIBcjXtf7jf5ZJCdL9ddLXA/RTdA1Ad3NJkdXLr
Tr+0J4LfEwhwmPoOuMlTvPDoaIHc8bJKdFhzlkwGEBaGkjZmPZP7GSJgX/tGPX816Fyw/GH4d7gv
Z+M+WsXEMAaGUv93xHW/mSJFnR9U942I+DBvDl6P8ihlzPU4kJTd9vwkjNdnLkPiz4YjZrhCTzXg
l5ZweB2kQyCQsWJj/6WL184mWFhjDtDG2hOD7yNKfjQZtKiubsKivBuy3W0rfvFKaeZ1pDtiGSAp
Q+ejQycKeM/0NSf1o3IQBPjz6NrgV38JKNuYhxUP6a28IcanX/LWylnVNVlycq+LeB5JReUr78Sx
dsG4jj0XU1U0hA2AsABjXc7cFQ4qvGlSfFUBWLQY8CeGxSZbeKVz27RULc6XGCt7lZ00+rCrG8LJ
Dr1PkSFV/wuMS5zQg9jWPawKT1BySopAVLQFwjUNrQbLaU1PP+qMGohXv3wN/D9eSXav0UypB9jG
YrYvwlnm0sIKDNvurpUT2VuY5JTGQM4FrPm7uHeBF2A2pXDvhAlEmweBAa+ACW+4krcoX2G5WS6B
Jhn9V6hFAcMU+aAagy+YUvEHACns1gx2tD7yhcKWse5UMMkce71oXiliK/mza9VCebHcZEiZuQ4h
j7so894Wy/oXHydbNe4z2BYyxVLIUMMai7iLfIs+Yzk4MY+Xtt/5AzwENTmJ8BZp1kilFj1E7lAw
kiVErkCmm011c3m2xZ6/2x2XRRJcrXgY/oVIv+fq7lFcmMiR5DkVjsSmfjgvRsi/e1lzvd9QuUN4
ySe7R+voWfSg4E441X21r8gxuvlfbIJAA2OBLXGVOW1Cy+8ZZggEyOSR1rVeRxaYgqxBFgSRarVT
Gzk9Y5o5niMWNP4fhXheBsROETMAKpb7argqZ7j3z53ssteZacGt3mXdIIC3+roekZxspmY8vybs
cZXqqJUlY3ZuEnQJPT7ERhaF8695hYRlnaz8WpvFjnbowhqNBzq/bD4aH83IAN0F/VNV0Ul6JbME
Y7yupI8tqgxg4J94xelXVEBd0oqJWk01TKt1wb/vOph+XunDoo6K/Z7RNhJxYFbHzxI+2KYN+sFQ
mXn4Sx6ERTzi5ztubPDBJoT9gVx1tSB7NxRIeiE+seGzClD6iVleRJ5qZIT8yZdGzwJu3i3I2nBH
mumIXuc+s1pVfJp9QpqEurwsKzGhBKLOlm8FuVx0M117+1uynDGgwRAt/liFuZb3HwkBQ13WUY21
cigmz5eg6Y6lKJGpePfmY+ipjpSUqsXtz6Xdxy6iMnJk+Ly7jP4OyBbapHR8WDF7NWOGDfigFmek
VQG10RlaV+PZFKOtcruiLbKt+oZafLNNhSyQMhsrpHyF/PFn21U2CLI2BYUA48k2pHfCU5sD+8eU
MvTCk7k53xntHR5dGwrMMrWSk5vmVRSuQ09FGqXh2m/NMYvtaZeBpdCJmpLkuNshTpL+BOMFU2JZ
zSmPq2kPxPlggcagSN2QL0KzK47SSrgUoMOOcDYui/jhIv8i1sfI/51T43CViPre3pyGdxekYJ3I
3VASkWnNK/odmzCnS4GUzr6GzLUBtu3p6JzPKA7OMOCSHRc2+zdgS41eS/soWiCJzRGfkhHrkpwC
VXOgh0zNAuVnCQSNqGqF+LdAZMdkw9vq8dgsYAPAOymsTkkYVJdsL191xkgSndlAZ2I03guC49IQ
oPGDzvKUd0Q+vtuVlB6Yd53w/SnL1Wpb0alEYyW2Q8bUOH6mGHlCp0gDZUxMWyvq06VXu5pgWwUy
PbhX4kSlNV6RqCvznM3+aug/FWm1IVgVYKWlkouOhddH5ERtv2L4/U3Uuckk42CGKYFv9+49BSLz
dekUDe/gY6GIid43pBKJDvcpjhQOcByjoVEv9+KJ2LCcvX3YFLXis2cn4skPhuOe7Hi2pPeRi+ii
BqIPRBiHuUfXndvvH4X5wT+GtFXW264M59bQRP7YLa9OyW51M+5VWzhM+hqcYgeXdRpUAfE1zMFS
Yt0IpHsUNZ6s31qKR7dMAKPVoYhZ2F8amcul7W3Qo1yBnsmm1uN3S5rnxzneGr1L5bI69Qw6zkjc
ZNSbmyEdoLKxCG4pEYseUFDDKQVTVuUdkHsIpOebyFH8dRzx0TGTbTQKn0X/rfDAGthwRWQjInY/
4OsklM7IegWPFNOWkInHdfxk3aOyaDU0lPifz26uPHte/Dn1t2RZuCCR9EEbx1qdp5BYhD3xjNnt
czK0HgWu956uhd3IHApgjyobwHQbtJTiAg+QEqWXEAGU8zPr+2d0Sym4rTtDbipmCBymKRPjnsam
OxDMxq5bqO9HDjgBDglH4hQ7tiZ0br9hdSxpZ0zayCzDTGysuu/qkQKtxL96APCngDN3zsKoNCVx
qyrw8CHfjYhsa4tt+6o/vxF+LtYZxZktjZwr38HJrVIsGkGvsrtEiFj3rNouKsHPh0MMp2O33ZN+
dFo9qiKFBCUWhiMrhJnZgO/C0nz7G3FbKS8n0kcokZHNcR3jiuQreEOPFrYzeDqtsaoSMRxk/Fog
Zur5Vr26js1+XuMQH6BZ8ZHV4vuOWOICYj+FRv7RLIko1OVdCrJ20RSWHE+WLeJJR03cry6huxeM
RQZVxpfZUgOuj2BK057GLTQ8f8PnDNkZAWhOt3VrELcyqcEB7zbHs1ZLDFEecyHhlxgTF5/2DfdI
4WQGvevYR/aWRycsRip9GCgb/GFBIWZOiCRnLDs46yUwsTyy0aGfK1lcDUYhkhCvTKSo21A17piz
O03uV4E03d++b5L4ITXjCOdjk7rvFO38wpkVRwowkK/UZMDGOqPpPorpP1MbRHSGDZdBDLZl8BBX
qzggiqc4H817WbyiV/TRlfRCNiHKzDiZDFEipg/snLWKRhzCduu0308Du/lZDvhAVdUhNNybZIM5
EER+zgNqrmEcyKQYMX59QArMg/ZlScY+qTautswBBcI1ispVZY0TlnigzAsLULBEXu61DY6EJ5iR
mtS3VwORC7D3cmCHUzdNLRGo5t8xb7UyHWUYNdZZ1ziiPfbhmrekNWARbjaCFehOPcUfdknkI/J/
A8jv/yo6kcjrLBUx/BLIRMGqaH4F8S+x3zWfr3XEFGTQqqaX9Pi+qE1dmuUCTsYznZxtyZJlOTPO
csMnCbJwKUvohqyWODjIq9TU0kgs8ZSBJt5Dt6kCtMBwIkNMOVigBgdEIzmAKZgiSHhnRnZZE/Bo
ahM9N/Xu3F+Iuo2fP49vrTrh65TgLdeCdvHcJogQbyUBr55Tp8R8A1r+6niUjIdQZZ+zjKq05seu
XQhgrKS94PnqFhBWVyJ3PNajbjghEg+ofcy5ZCpNS2zhlSYlcUAWvXaLZ4tzX6nIIwCTl6BbAONC
ZSKXA+hVon14q9UFqNmeXCZK2aYBqnMrdsKt7K5bmO7fBVCKwv4rnNSldzvZXsmP2f/i+6eHtm+X
2F/cwVa/i5Nk80jehUPjPKiNinMvPl4jsNmeUznFHsI9tgCmkEeBucWG+DAVaodvq+aXFWlKaG6f
5KQU2b+muFtaI+y8O851+KuAGi0l+43XIsAr6KVmp18XtHFKWrG/T0jhe48moa991KCWSV7dfCYW
BBeGAWAy41OhAHApKKZkAiLrbmUOWjo7IxiRY/oZ/tILEH7Ef1gXEFFJc0ZfRIX37w6bIPxUDRrx
AHddgp+KKoLwr8OK07aPVKVq1U3pzPMP6lCRMUenYEJCNrKfyKDe51kjhlz/ZkgDsK3Wc4sECrHt
0N9TqP49t7IeIcvLl7WEnb9tNm5smbZl0zsO+tsOGmtQwFEtMOok/X2+U3FY1SPuG4GZf5A+tbVj
VhlLzRWkxESFMHV0RgtOlVki6C66zaozWuNKIR+f1yWnhY9QXUu/G6HqKP28h/A4W6Sy8jVwmjz3
donIGBoOwBpVFtB6VstSe4MJg/OsimFi82z4sxLjfhsEhLiH9l3inKppVgTV9d3CkeHYGlTz98bE
MAp9ta2HqPbyiDz1VmkCC7b4yV+9ATEtnehBl2+TGHMzEO0g+hKDnpOQg3yNv5wZU5TrEaPyFCZz
nBC7yuvr9AHdi/yB7IhSTpewOZXzZ7pbjPgOHBHE4NIjxdqp7LQTIMLMWVryU3iYoSkNvcgcAiY8
KxLXB2NAQm5IgwGgjfVbmfUJBKSQQXJhb1vJUk75AjWW0te+uomCGj7D0b+7rIA6ee9bvRyNqRF2
kb8lxZ83Aelj1K/rs1RcWWZ8j1ROYOsEmi92kGeZHvBbj6nya6T+dtfKhEC7iUShvdUtJgTOPRRR
6ZL9LZou/K3mK9cQeozc419FmVgUk8LaM1VvwgGm+fyVgeyGVqYAL4E2YZ8eCLX2wrhE2B8KdLUp
rziZ4iRbQNdKyB1+fdZWuZ8lu3oRa0xnquA7e9a2Q6xE9pAI8kv9XUmpVgnOK/Jim3uAZm2VvW+l
1Gfixt7Zb0dGZht+3cCd47NLHKeAh/ekJaYfOnZYGniXoJWxjn1c6Reg/omBF7IU47Tehruq3uuR
m0HMalzHFYhWm2/Pa7gqALRZYIVdOXe9e4vC7tNqT1vpKg0VBEjjCA4Y1Ud0PoZh8ainN0/t1crh
f0Dxjwy586pskoCCPn3YDyRk98qPIxkl74kFDKrZTk+W+yCSFuDLTPR/qoMRGahXR/InJPop6wx+
H9DTId4lJ7kWG7HZfI9Vi4mz2+X7BxDtO+s4me9IqQ09ZwR7Ic3UoX2F+GBjgFkx7M2ulFGyOp2v
V7DMVBdI1qi+eeDcPoyqQ/stUNUvxIcuw1JwSVw8cb/Q0avz+GQegvhKt8ZEloj+u+OssQw9ZoVY
hpyaIUVGd1ZN12jkoAgJqipyJkDb/O2vkhZKrRWdmxY5IZxnOwlmIuM3QcjPw9jh8frGvqV8xfh2
QcDPTaej7k6X7W72z/J+9m5qSnePkWp1uAMpxs84fF5K1k48o3UiZth0S1OiejcTsWxEw2iADf24
JnPveMV/eiYfPgQ1uS2RwV2JF05qOn/ZhJ/I/IPqmr3Qg9sXlBEXRLx6NdHBh6YZ1qbN3iyyuzbT
EhqXBeyFBY66Kkk+GmCOr0duXke/bvh0sBX+p0lCW34AgTsZgfBoP7wzkSxJtPqxytPnQy82qiGj
fVT6PCxz0W/vUpEwaQ7fzt8lv/kG3UbQw52sPDpDntzoaif0X6Y4C4ebPpFOCz8/Qpi9lGj6HO07
X8GXE1X65yhaAMRZVwBf9AMsH3rIYwKyZuIqZniMqviYE8sky1Zh/jPcPgS41F5eAknMVWG9zSyq
w8M4TCDBcnpuyuG6DCHPshGWxwmePlyv+gIwX2HPuUyrS943EJX7vkAjvhDcaoYMX+afb3G+3hD+
LiG4vep0/yd5IcnBL+TpWZZU7Qai8TumnCoQshL3h4Po/sAKZXauWF8bLx89O4d45xzMpJZuo8B7
r3K/Slml9oW9DDb27GWL+JF5prQAGjlp2YPvnZGiOg9Ibuw4k8y7+EFuOskvVhIqx+4/v1r9qDXN
kgJ465VIdQjUb3tLk6VP2hqj0vULaaJ583ImwfF7pN4xMTpdBwEWK41Z4QrGrXexkg+tSJ74L8uH
XGQA+F79QRrKiy+PDZy7ZVJ2/ol+3wLE8ag2V1SWhpzzh6gXmVcsuA1PKiw7Cfc2BBTZokQm7B4t
wIjP5whGwOU+ftm+CGEOxs6rH0c9UY83SWD+3DfDbXCpXdqXEQB34pBT9E0B7yaeJSyeNM+MYOBL
A5RdHn48X5XW6KOJPgh9UiYzME8nWkI8sr741Yi7Q0iVOhc5vSaAihoTYtjCdSFmuWucSErsCPRk
Li+GkaG7C3oiLDX7qH8FVaNKSHZ+JRMVXgRQ1Pyu1VQiUWuptjXwI9DlBdBV7pE3/VUpZ2eFhhf1
YDr9kNcTzmZ8eBy8eHylBLH0tW+q30/Lwa0ATZJjIcn6Jp7lECHl5RjfhMsTTz+6ziNsXAO11ok2
SLCmBU9oj23ozRbmFf2ANOMjy4PWVMyzmeeLwHPE+e9o7ZxvKw8VmbyUqgf9rsvJJoUqzTkI+NMv
TKzDBA19eTrk5HuGyeWlY/qKdn+tcK4eaweV440lfTRCVzqw4arVMnd+Y/HVHtAVJHbWclWsSoeE
AKV+XYz4GP69h1C+xojPiI8VCuGbIG/8VBYQQhuFSssL1lv+6Ym07S0f4s0Qds5Q6vAqNdbk069K
5+6/gcsm+UtA5u2RoZ7m6YYb3fRhWtdpieLS/dKuN3qp2p+zEUI1BRaeDsM+dYst0oLkm5o2BXzy
r8Z3i298TezvliqeVnoay/TsfDYarCdXSYaHZ98WMTKIzv+KGyLRybvrYUK9N1/mpbh4Py6JA19X
rJAgrTuaCp/Mz9TkGHL2mGc10WF/JMjwh5QEP+a2LB0K7C4Eu8k5ebA7s0N++fhjfZQ84hRIge+j
ghT0fOXSdCp8oszrSNVUSFJBRbJt7CJtijgE5V+FnZFfEqaAbKsaqcnuWbRQMAWGsODfNHyJlQr+
MjAptbdBSg3OiKvoL/KALYhCABD0ACJ87MNI8uIg++ZV1Qoc+rC9dVyxBZPOu/TN8Zz1f/7ym7HX
B98gKB59roAXC6Ge6W9ix/5FiR0+R9I5x+g9nISy6Jw42RVZGcOX3WNRGUwuOFJrO+i/WMpA1tUY
w1ug/azcllQr+GIzPxiIJlo4s/0FmqYhourlNzf6Xlsm8GxqAU61LOXpWqo8VnNkwzd0IgMjqRWw
Qwgj4Ip5k7MNRLbXTYqllgcPelgXdXUq/qWEWn56Dkiv5eH1pPy5WlcrRfBvMtKgUsCEYC0EnN3a
ddueYuebGttUAG76ma08lEwuhfJdZXZK4rQjia9Zev2xCekqk9ttVR1O6XNmxne/q9yznEdHWIUh
sqwSqA9yRrFuDCjuJEUgztKCx4WMVluzn/vy0T82876XyYgWFnlni+Fnk+DbBx4rcRXVkxaa8cFT
tjSASTLa3hccVB6OKB4rAQ+ApMgbSmyJU+87izXAJ93L54Yl6txfiGy23pSK2GlRc1Nh6Zf5D6fH
47kpKauagcKNKeWzVBFM8w/X3JN8ih9GPm+CIaW90U5FVCkwj9VbDdnGvfVTxRmmMLIDQ1GnBCcm
E/Tnq00gLXtCuRM6hEC6Q/Gj45R64cgNftsdpjqXJjUU5HIBrn6BoNT/vnO6pn37Epzdekep5s/w
7pNrjHyG2Gdlj24WmR7lxfBN5NH6HHgPV3iLkkG9vrDv7DV/ZVTC8Z+6xF3nlxvo9EM/7U+Af0+K
+eTy/QNzDhVsw77mI+WS82t1mE0alx043nDVUSqIe9ihDJvLgB/lC0aZfFhUYQlwG69j5UeWvoSg
NxZL8YSAV7r2GJlLBvUVwSUBaWZxFfHlt+NX7oPecx+9wboueIjHq2wdHvcSbI/4crR8thPngAlb
COjyk3C8WebdXHR+D6tcK7PVklFm1IFGkRZJq2Deya7NbgKAAlaUmJd7cXgEL1yHc2piyi04zPtt
f0bnBJSkVr8Kc8Ar8pj9FUcerXrIk3fSSQY8NfILvzPIofX+rsgsxFmg9+XUJURlmVvntVkEZ6qA
IAU2IlIzX7s8Gepf/Q7fs8spI+9gISp3MojVOHfTtOSFcBjFQR+4DH71D6G4HPXAeTmoC9pDIkGb
Tppcqe8eutcQkKqJmeahfGzY37sbqQhel3OR9nsPqEza31GWk2EGgn78KSdIwX43phI4GaxZm0LP
H2kUyYZfgftiJw2JudCXVRxqE89JRMXq+oAtFzfUqA2L2frAlyxXS1IKfvl4ahM5o5dsupxkkff+
8sWBOEcODayIYCZviic9MsHqlokAjc8RcOhnZQALHtRij9cztg8koktp38zQwL5MjsWZa1r4cqsA
K1YNm9qSbSIg/HVidh2KdOXXBg5GycL78stHRw6n0Ef64MFMc4M4PWk2/vPCxyB2kaRQnBlWEVzn
YBi4p8uJ/cvEYm06uBOwFJQKr1O1B79WDctA26bdz429sqfpsq8WF9DOoUV8UvZy5f+62Jx0uhTQ
tPmVHAQOSsr1hgY5AF91vPZvCOQ/CAQVl6yw/X6gpImjUPfN3or49S1rqOA6GKjV8K2O4OIxWyrH
kqaTNngUqqHOV9VgggIrNMags/KYQR0uSs40A4K4XBjTdCPQ3RVaAqj4d4DqYz02KR1QFfvAna2B
V6gu4Jq1pyOuiRj06gOyQJWtzNspi4ASHjiKk66DPLsbOyhYLb1PxtMtIWaJ8hiRe7EG6JXbEQN1
4NQWcrfdFAZtM5zOMdi9rd14mhakOjviiqYnzOPvJgXGUakR/a5yuz1uRwkv+mKEYdGkSaRWCFK5
Lbb5NTBiZ9HiWIhW70FTn+L6AuOcJ9ABhxMB2Y4TxMEvM3hWHIkY6FuG7MCpoJ7lOLW926eHEWsn
ZFwf+/MSwFJGgkKTNy8iB1hekClrqj3V7x8xsvb9uqlkMsxBd4QZFQbi5TWIzy075sp1NlRHXD2O
qU2Kk4CGMSdhrm/VCEzVJxQa/cAFtPr8YM+uI8MTqcvSofofZ6CWgDYL00RG12/87PP5QMHQx7BC
KZ6lZUvCEtD33dwCxHg5aDPStgcrpcP8UaoPm68wYsRUO/x+jo2vK3XP8VnBM3/UZhN0/eM/mSRx
TD6fa7/tE78EUy+zAdoF5dBoXGLDwgiD135a0ZwKSOFypTGqYcylKj23aTJ/Nm6x7Uko/ft+d3s1
zc2yqICRH4OSrVUkX80Ts57yh4l9CWBGh2eTa/LzC/t/RFQE7UYx0C7WSC+co9MwnQmCgAxjh717
bYQtf6F6dynQQ1gL5tqgqstV8a1dpfGGVCNezU8eJjoUuqebYBYQmp42h5lKx2Ce6DM1w4Y4VMrz
pDHnyc1bChYXoi1w6hLNx8F4900GimTXvboU7ssTtNSdWWfrXcDsK6wMmyqUG+6hnWFwbb8gd5uI
yz8LRXH3ZGb16UpoyYkYfPE8P10lYxSAjTbpmM42aDG0glgdUlnrNhPsjS8OXjnk86LbEdImTXex
I2EBGODhie/56ol6N8mQoBPFVX2FtQg84XrtdoIYLUVnAAEWxwSk+4B/fyweq8pNBmDnc5wxt0if
nemTwfrK2OUd5zY84wxK8wM+GKxtD+7/8rht0XqZaXrcGFDMOpqkdaqu2H69yUjUWHxzDgLej/fI
x4VxbaPL5RdrUUIy1D4MNiQfyAChEnyboHeWefdguQAYwIradukyMJG9u1Bmt4yG65B4Tl1dC3Z/
lse6QAbpI1TfyioXXyESuWUKy4MymHhLjklscYO6xaPsDAWSL5r4OffyKOyo0i1z+ONSKFJxtKz4
/CcHy9ptLy75NkldQ/JktMUm2gZEuFNjvPA45wl7pSmc+JHQ0TV2648P1uLH0A2leTCwpSivT4YR
K9GzEpttmAOAkyIjCkj8D2xAC4MyB9lyH+Bc2eemdUKVeAP1K3NcEysUg2J+cUXlvQ7okMKmMFeI
4zrR9PH/YdC778bWo3Q59IHzcHZbQfPVGmEoDhG6YyEZ56bSu38pO5YSEiMIISzFiUyUlob0OsgN
GPw8CcHcTdFON90brVhawIeqACbMN0wz40JIZRxC5x7fKY3PKUWOre7+PRjTuTMjYiFvsjoTKj2k
Wwcy6Lz7Vzyi+c7o0Vc4EkVfjHlW12yp1FulrN5LYltgx0Dulu3aYMpyWU684AAzO3fPz5G//AUd
n7HYwKtKrBoymPkbGWcGoLrixQHoGtCxWg6AbgkKBGYfovtk3UHx+tdXJox9q+QRqRWwCzkx87IO
9Fy0ybt4nDrji5cer6I4gIkaGBAs2avJ2mnvZgardV3xllXmsj6GRvTcIFW4eiC9Ue2CZQ0uUi+g
hRsfgL+dPK6My6u0xPLBjYsTS/6O43lGxHY3GTVdtba9cQd4vcZ1dqhLfmI/WS2KoPx2lEogE8DF
IXAXQrjcURrWS/cDKfpTz/jlG3IVUUxDtxWqMlZ1EMTEDHqCQI+Ha7qYm6Ba8696fv06dkXZlHup
LgA26y7xZUS7t847J0H2F52hrUzG37cwtcpnYBme6qfYsJdZLfiEibB/VfJzTxfLoilUEYJXl0X2
Dgcet3WMCSbzFv4qAWJyVm+OD7sTilPp3Y4XK84ErtRwXcMXH0JnPwX+AxyHI8v6lHyDPP4mIfJt
7Gl8KLXkeHexyllfLZeEDGtz4L9rkpP+KhcQjYMfvakKAABPnCqN4ZGM22TO0BYWQZmYQm71oCBW
RcjBf5C5lWmjjM4Yjxlyq51jGUjv6AwAdJRq0Pg12P5+MqTHBuuA8JCo1XapVVIpl20akvAl2UUy
pKgCQio/NHvzzJxxefPGDQ/iS+S3P5dpdXJVKD7ThIFpYOoUDqiSuaVlsydm94O105G472yLwLrL
Bi9yfX/5/HDR7T7wYP5evMf3FwkI+5lqPYE8Ss293M65JpMZpv/dCN4VhcHu1/WuJktJIekUZGRu
8laB6EPgaCAXFooE9J8gnr2Ln5z36WqpSlH1Kft3YjplPDlXnS1/jc5Hg6tqhlSw8g8i4AJ9dfhK
AKbWKTNHa/92DQkQgA8S7uO0S6218IynRSs3pyI5nTVIKmh0DZyznWSK+jKJxiAfLEjfZvuQeJtD
pOLkn0PfqqkL6DNvw6auPOPZavAmFeDbFIaiHvsAB+pNgNuEm75WPksDLy3SL84dEjYZSq7P2qty
NEI/AgfcMKHY7I66q7Tl5OwVn46rFukBYn03YSo04ltd05NOzUThbHG9RkU+uC6sbXmgWLysAJuP
3ASoKb8ZqxsXfpsw1/kL8mwYFsFG6qP1Ob8bt/I0ErRnoqg3DRkDcwyXOqvjlVueOxumHLwI6z7T
NLG4XLaAyaOMxE8re29f9zMjIoo5uaNV5InpyDvTSRNhPqoMnpE1f5ofr/aS36YNKu8xlxqHs1yD
2jyyce/laoDf3PV4N4XkDkOdaD9xwnUtK42lRLhQZyI3ZRTPIaCNOmjIC+Ret9Csd90j32ocL4zl
NTG+48Mv/qxX1ZgW2A3mPH0zzYNCPqzrbCDU0pDn+ffpfIoQSPHuejwM91nmraP0ux+bjhVBN+jM
0en8M+TX2xGVHh7z43c1mio7LW4w3atQyMDner874DDrj2ULx3cW76wgU8eZFdtVjUpv5mkw6vq1
yjd2O/aBhkstfryMj1ukaTjqRqOs6KLkwk9oDQyd71tALgckk4OQhRxdhfrjwTTd56bqKUD26cTx
+ELEfr7lR/e3A/j+NnEi4mRiyR2+t4zxtkJYy8bYKuAOpuiOiDCXwk/XnIvzwWZBlaYJDhgnjkPO
GHG9xs6gzu7Gm6CEZMY2uUJ/d1uKpy3/4Y9inDEBPrLbB93+He4LXxb1aOr9FjNjSaq7+lFKqArD
0S6V7jd6V0FPXuS9XGu3Js3+34dpLUV662s8fFd799CHtdDz56AYwM+pSvBNmFXCP1r8q8rhHI9U
rJusqXRYMOZEuy395xdDoQaTRgDYTtXwgdIf4QXotddoJDPvpyySVUTcA2EE3LnpJmsSuC0BA8tK
MddDaEYe4EC4PhdaG5bitkIjhLhlkc+Va/ehuQh8DqnC8n76SoQlVT7ii26nQb8wgCPYmrJ4/FQh
H/qssKDeKmkkUX28OeuUbTbqcl78F58PNeDashNSK5IqbGnCH57Ub3yMKmt8et14yAUqXGXdlkMx
scguk+2J0XBiXeZNsW/7EQLt3TgalLMpVeP2oro2a8IuxVHggRLOFramWpWKrqj0/N4SDstE0yyw
HnzZLGdOVo2v+PId63WYG4vp22bOOPelYz+5WvrKv4x7NiWE9iVfirxydyXg35/x5028rsLQaLfB
tCCk7AzTkfd8U7viPEgjZDHIAzJYKqQcte5jljjOvBOjXSKQ6PkIzHRPtcZtrGZdfI4Yp1Zi0jAf
0y2sOCwarA7dx8s4ZchAc78/X9qJJ70rquT9qe++eZKugMgC+Hktya0AE1XockLnxZ7nGZvD0wtL
1DfiUaqHvHqZbUNOzt2Hze6RfXR1xVQodapiRP3XURSjduO4l8d5JsCBT9jPf/6B8DO8kdpXyKbg
fLjavb3V/o0capLyN35dpvNPdG+s0F9zzqKiSkqgBAh8xpq5Y1fR7nJ9mrb6R5E/X6bwZDl+Ofyp
dl7KrVi3RecquI8bYoWBbJxwFeHSLQrWSYFH5B03sKxxxv6vbga/uYG7YiEWoYpN1Zc4pjXxyJKj
PFFwGKHAKNym9zrJ21UavCyb2hiJrPovzzrhTxPjHxjk+M99iAwpO1AZkYXoU1Mrex/V4AMtnSKz
yhjcfewavAFIXlsvlNQW9ucw2YfRKWIT4hnYACRULsoaPQIkIllZQXZtpINsMClX3fCwirITgp2o
2yYllQIt/Itu9Z+Ew78JRkKXwSysjvwS6NkHY6+k4a+Seoufmk+5JKRl9Fa3uIlS0ft0YltO/YLD
fZK82+yNOChSqAIQ7un2nE4yQfulIqLoRCNugZ7mjBaWJZ0ahHsBR3LTGUdTe2TVpVqKm9AMvtVB
skzYEMwSpHke+NSt5WACpDW+AgrO/2WidJeIW5M7cIIJNkIe/CjQwqIJYQbDysMSLBHaoYdOc4or
PhWlMPHPqvmr635ynZSz5Jfz3B9YCPSNiQNNprqq24Zrbd15JBiqqDyMPw/kQV+KpM6fq0LuIqNt
aTK/9savxK5nlZIfSV7a9CwuGXr3nbUcOOUElrHjlhhQeQwfuJdtzGAEA+Y8KmlEPzNMBoUSvZhZ
0b/019gJ1GLk2TH1XQ85i/8lF4XmT10cDijq3DeEcWql5teDVrX1cLhJ/df+DgshBJDm2YAGKHhR
qKM1DZhi1RCjLTGdZpyi9Sc1VyX8UCJFVEGj5XRN0w4gKnRenTmjfcROSaFcr5t9PmTGPGAATGY3
DZShMOVmUdVke8H+9eNWILqIFHecZ/OHOyqmWW2uKlrG2wU0OKaumHcyEErDUv1fBuJSdWvAAB64
k2iS15fcEprcB2nCU+H3GrBTbpJJuXcQDTitwNwJUk2dSfvNFLksi6IqTDgQ44P6TusbinhytuLg
0XT/l26m6DxlRyQvMz3IK/tvSbOrObthOABxT/yiqJssjx9NgXTp7uAhWRHdtNxDqvlrsELP54Hl
un6eCCmKXxGByKmT37f/2+8Ta6XcRh5RFMBLLcxKPlvqHLgcnSIaIRe3mXa5vVpqdUa1xcrNOdJN
qkI+1m8NTk0QxkRG/tPoubLpJ0j8XzpsT3wTtE5/TM2xAMICRCfVMz6q2+jtA08gDcKcovYrBUcg
p7VDmL2y1sSDa6/WLG8sFFwLj70lppIRes/IOaeKhtvzdxLihjOm8eqCkVYTNBKBJo4Fnifhw/pq
ZbOCOYZ6iFvtJ/z+L4mXIWsVhVsLVQnygyGvsAJWaaRnCjoKk+cmvCn2pjvDqVrb8BkigSqUhhYC
XkAtLtwkBnBA82eBDh313Y3PLR4w3S51kKGZlePDh0K867fc98yB1P0BbbA89KLGOrJGhrXw5953
UOG6pYPpw03pdmbXdNQA+PMgN5B8U8k7O5iVx+UJxcqD04E8mzhV37JUhiepnVQrI2epVRUqCWQw
qzz51NkU/bsiwqn12sEdSivlZ9llG4AiFEkdXIlOAM4tzEIUFl4aqfKhk45oxYh0+Hea0J3yUU4e
BkO35tcxykmd/rPzMZYiHW6+aDn6RtgXMGbYo7pc1XXP0+q2PVWUFARblP/0U8ed3JxTdlHuKy+Q
jCjQkk9GbJYoQ5oS8Se/e904YXsQ969ra+e8hFLqomfcynL5LfoALmsT78vxciT0ZkV5Q9kiZ8MZ
P1t84OpoLh6bpOi06ZuebARqHm+aR1mAergUs70e+n1I/s0bPw7BUZ5gh5K/TtD1R0MBeJ8c1PJY
mJTBX8R8/YpWcGUskYMzQrgETMCF+/46l4VTR+kEfQD+1Iml8RUCMZ58IeG50hG7ZMtHtvvSyb+1
TJx6z0SJ6QmoaLslBdMysdYGsKI3nP45eTPeKb7+32Yzq2mpALVTQyUpCUSY12ojr0lg8ui8t6qh
NxodID5NBeecCV68zu/X7adH1AGHGWAY7qLWeSSNbd56xlEwI5moFinAd21YBrV2vWpjlZLl400q
FiRyywrSKxJIUHSqHJ/sgF4EVH/Wf4erUM+jsOcwFGRFerF/ZTxYGeIQpQL/bjKi8FB7WNk18VCZ
4Zf7FRJDVdWHWgb7JBrOyMSm5GQH4tiEnjUmCCVtrlW11E0sbrt0N5LbJpdWWNDA6mILTOyhAHIo
6VNsk7OjPxUVI3n42XNAnp75Dpji6RkIXfA7MgZ9bT0NZruC5dxfRxI9MVwwyOh2L4aLNhvBMU8S
QKCwznAFrILEHGDo49DzMb58EjcLU6pT9nQb86jPQCiDKgpLi+zXVgdNwr5oSMu4btXgJvG5Fu5/
JrZ6Wqmmy+53Wsidx4Cr1cMYR6ouM/+LdoKhR9v47RXw+ffnvrsAbkoBG8AEIDSGE9G5X0y2ltaG
Nba4moJhit9DnKhZJlR8rJrdFXr4icCO+MNYBaa7mDO/LymJJNDhG1kZlDjX9rB+PBWh0rxTGiG9
PTlsPJycwzruIrlmrcWQ7QU3Gi/rIwqB99EldWaBdOlFgnCFtHBrfMXljNVyd/oypWfujIElqZE7
5vByHErixN4tXXOCn11tqIzJ6tWozlTSEtzjLbX9b1ijWBE+M4RUnraX7zGPxBsrvG2A7r/A0PPX
7wCVLmdvVLrvgoWMyuyct+KVhGSE8aBVhHZn/tiOPgwWM2iaoGizF12k29aYf0igkj2HH5qhcAHB
tWH+efaS/R5yCndL5HQIHNaz84mF5SO0dfnDqsDlpFyHd6gKdJFfpgiJ/BCmf0wo0mU58SBE7NRo
mRUuZ+CkS8nvNZHQnnofgJrpizluByusdZ3MU3mV2NG8N26Rr14Uz/gOEMqBALiIoBSKUQ8RKZnp
6/HdhU0L7hkFSbOk5DEvYcA3ILfRmTsH83jXxO6dGGgoS+xSQMP2MWhff/mBiPa8sN7Tt4ngtUx5
Zq4Y5q4nuWoBWKhUBUDdmNvWv4J7GJbH1K64RDRjVxxdXD8ELHSyUvfYFXU3YwkVhhnVAc7S1QMf
XErncGWUbwyqzXM3Wdv6bRNoTFSYsQ4AeUq1YN71g52aU9JDTuppqXc8rswk4AWzGNT8S3Cyfc1s
OfaN/Y0spuhIrgAp+OvX7uIozcCajS5m3f6wet2QiHPAOM1Tbzrfih2qeEcAQ/aQ0q3+Xcjb6xwa
hOT0se+vT2hR1i8QT77nzeregAK4kKRBOYio4Qxfu94eH/ZzT47fEzGb/zjOLiUs+OMcZhEW6hVd
CGWDXpi0VHwsLhJq2xl6EeC29dA8kakLIKgS01wefQE07hzj6ogjbU29pXq5atKgplgSzIsuS7mj
aScwlwiK/q7PRb/UiQToII6Pk4Rqd0HStWRpD1qaMD7TwgbyIP7m4jRq+7gxX58Y4mQdYFCn0NN8
0YFU5RLnU28ivd7yDGJy2zp8dYtIZsdkCoIa+kOsfH2umEmb1Wo7EdjMhXQEhxf55Q8gcZ+iOl4y
FpZOyKZZBwjj8ENVowpC9oAVp1gNbMWm6xiH7ERmAxOR2/9bWsdnfOnUM26sWuaHBLoiWCUNW7rU
l80MXexWwCFzrFKdWCDpnDNSdsGbvdmKrC2Bd9ZRjLDKQS5AUuxxflvWhXC9251MN+DXFQNcTYKZ
jmMjiY1lCo5BETi0SqUkd6lbQ+TrJ4tHA0sHm4gVdfPTzu5OPueckg3HszpaJn6b5d2/Oex+0cAJ
lagBpdyjfemDbHpXmTPFoBNaAB3QpTCCA+zuc3XwDQ1Xu+q8kp0RKh1euhAOf/8hJbAk8/kJNqP7
0UfbMoiRRMpeETcaRj0tW6KbTmO4MfRpE6b8BRtBk74tsP9vvrKPPHkjJx12LPyv0JsBYAs6ukm/
XsJyUloZMezdWAm6xe0Jx9jxxvz/e0Nbq7BMZVJM5REl0gYxKG1WbBNN0ZQIlwEs+UN642kvmvQX
L0QA+HipO6aIyMTrX2tduG9V6hinPfgvk1r3HevmQDl7aM2E9/XOfw5HO6GNgi4VHGfl3aqesOr9
jT6wO0lW2bmpzTYDqDu5GGUavO9O6c7pBU1/sdQ7H7DAYbWVNhs3+NQjjA3h8wm4ogpDpVx+V0kT
lpdrVjrn5ztOmVYFbHnVpn2p/0Mzc7ZBW6hCb+CKEQJMxd3Fvgljzj5UkuwkvOya/ar0VrDcwO5i
1EMZzJtNqvejSWDh/HzFcn7IJzh/lJeT8/R+ZFDF2QSt4nKJCMO3r67Z5xtIkV8wlS+LyutbNbOv
pIk/FlgpX/2XOgKWkUW2QTU485sw/GT/7U4pgTh8ffrgYZlLUz2Jb6j6pER52XiGgDC2YHL+QVX3
yzkEGQdmIhCzUKMGyXQYQJ4iyuV6SF76W2xUIXyvWFW1pA5uiOKNZH8K58mJidg1bqwLSHRPz3sH
mizZ1HJRq6+TTWDFYH0r+nGTAFvgw8W3XHOScLIftw1Vw5LOhDLg61mNIpI0mTphkoijcWz7ragP
Cu0IcHSiYJUSYuVoqljJMrvSX2lA2yM9vpk4F2ecVySKlMP/wK3S3J9jjUsUgUsw/K5yZ0OeszHh
Z+ydf4hKZ0CX0oeKY6ekxMh7oUQ+qyLQceMZjaVz6UrR0jpmh0Ti/IZSOg+XG9cfNjGsy/3NejIe
GQhIWh++qO5i4a9Kaknv8gMIXl+Lz8+9buurf9vTequxbyUTsNZwgWr7D/pDVT/WpUkxqpTgwNDK
GTLpz2NqFnSm3u8n/Gu23VVuZ1vOay18SlnNgpErPLa2w8Df5rphzpW2IEslFQuf6v2Ktqo3K87e
JTu+k+przguzfJ0HCDxLRWziqb8Q1/AwQJcNj3/5WWg5Zfm1eogS+YpFscs+H/1QIFW/or7uQCXc
8wEvp2U0UBcmEz2//zqah8jzb+pHqc7K80EVhFtnGoIiRVb91zPo3kaGee+6F1Bo2fAd0dY9wtAW
wxRDAvcEtxXqbF4o+0LF593XKuxiyRxup+dV6qmUeZCYPfpvCBZy6jOIyjMDOStQJWXpnUu9a/uJ
QnUqYKFIXgdE3wXTNDSTAAP3xvL70GVQ+dQQojUVj69hENgQ9wg4/2hzFj0BHbEv26jYW46O86Wy
GGzyD7X+f5qP0WxrOV+BfagPCokXun8jmvGFkvHPTJVepy7GtsMl8WYNHdvc5NWZ+qLBgfdgf9Nn
ZXsn7xPjtxN+ihkvH2AoPuzIjBeWu3bwRa7FuowkjWEuF5ckDKDsk2Zl7aaZnt/YwIvarN7E6NoT
4Tty0G9oq0+ls2XuHxpdTEvsWyWN+SFQYnZ7hprKDnC/ojy3cI/SFXJEzlxwca491u+fim0+pWxU
3fWQGlG9jGsJShEMoEIqsqAw8xMoS2ysm+fXM4B68w8E8GYTqHxsdy79/oUvV+shozJLzcrWdISY
brOnwPk7pmzsUMNbz6g487VzlQDrldP0WKoDk+Pg2YEdNE5KlN+oMRKhdWU1Xmivn7pXctp6gaoL
i3FKZb7D6+cSLrrUuQkZuN0TrciB1T51a3r8ZkKmw+PF9adcHqHTtnFdZriJW5k3mSiRljAZApUk
acQNWnNp9csqGJ4Ja41YtVCo5a6Kv8cJ60jmQS0g9KIVdjM9wJr+DfoPRAHDXVl4sKbiwmk87/F6
F+JjGjMd31N2JmTTb27IowOEM5PqRfmkflj9Ky0+h4rYQcXHbS5lnf2nbREzbUbYhJPBQEHeK6yh
CAqPCto8m1Chjvpbi46oPQBrxFyaM2mWHWVBvOqPZ4yo1BPmucbfLymV2hYGW/xEXNFUbE+BUt2T
O2vPFPGNr8NsBRY38BAXpOkkOz/RoMi/7G+nBDLAUu/0YK3VhojyaN46WrQWw7r3w5H22bd/xHn8
E3C7sVmFOcIhHv/Kht86pRZcfzNdEEyhW3x4Vr0NoX/ECmStig7xwkiSb1YUZ/DpZyCNcmjXBtge
whU+c0YP1jJeGbxxMNPn0/9A5qGiNgOawxRICu27AxXLrVU3gbJlr2cMbSZZc3xkAfuZ8zSZV4JP
zlGwBAl5TWtdZtYOGiIpptoJ7OvQSkmFVg9ffbm335XckpFmN4i691hmyF0rNUhajftjXExvHw3F
/7/hzIiQ1c74wqi3vePVY337m2zq09qsZ5RKqVae3UdJfpQIFXYYl9UFVonarMPADDiHXBA6uamB
cGyzZyRGQyfRreHj/+hTE7m1IvWQOGiOVbw8ZvudTpvw3vKwGGIMZUtFwWFTTz+jmEtLVZ6M2OcN
Zj01XLuS8TPlOt6rebUtftdbuA3G6j4KLOq0BRtQhFr5TOQ/z1rlSGprMduBT9tYtXhg/8fpvlij
MJak53i519EbW3qvIF6SBKQ0DgUpt0rDGyZH/o0f8Lza0MxY3oSGgNOvjQ/0EVGf+h6mhpUFUbtk
iwmNtW32qNxbybyK7pbZncD8iCGu9OcCRsOe0rutDfN7F5OQJnXi0vNkWLBxAhbjzDvjS/TLRxc/
GzZD+NBIeEDXT+C1H0IrYV2eEG8KKENgTTQ3CoJl4hm0KSocTDJfVjjD+QrXDlCuI/eeQKSiYEuq
qRnfeBFSdwd/qfTJpYlNZtcKTl/6xmAej8wwD5jh8CAKYkoP3qGwdwsK6dJejho7/bwQ6s4c+6PI
US8IcB2jiyXtjSgRhtlu5Qe2VsQwyI9MDrcl4jPa/8Hh2LOAQkteF9Ux2gI4VhyPUGBczYMhPKM4
iF7jqERONkFAlFU42Jl/IljSEcGi+eimlmp/ii5rFswRKgpJNpXUUWaZdW7Jm9y1jzfn4v8AYVfn
LdIlVjGNC43nzmh5uFtH6VzRdJur0vULsy56wl7VjC+Qt/bMsX4Np7jNpG8ah9NU4PLfedt248d/
veoEcYRm/XNk0C1qFHjOjgsQFXHCps8bIAldQlMM95JyOgt2UKki0KjSsovnRNxX0KynQBB/vDTE
u4Aj0PrHHsrNFgaT5VlrkqI/LVzxDzvHoZI/1bJAoGtbfqf5UtlWs0whBBuzezPke/d1G7abNYlI
H4mfy4nKdT/jVpTPqbRr8XtCmXTqUbq8CU6gU/peRzWMM5cWN0t9KhfEGpqVENM5KG5Cb5pcpm1i
q5QbYr42Al6R4wppqHmBtKxrtEJGcYyWFprJZ4kPNuE5X7ZSF/UTp4K4aH/uKc1Wvjn9dCeHnP0Z
hS0L9yjiZfJxxnu92oQIC8/JridNVpKQDdrc/AxKnt36EA31M1Jh53xUkTyu6QVg0ZRV6tOWX1aa
1T9d5r4HGDgsxKmu9JltAx/inGfH8U39DU7cfop/3x1vu5HZGS9dzCiv9eZ9YxPwQggOzxO6QuiI
TR44CTl0ceNeTauVW/VX8PrJw3XPM7xRQ/F5LC+dBammPlDEI3JWK4iGFoszSFStOFThLcIcxUFq
sKUvnGdVHht3cGwc35GPvsDA/vNA99dGgpkhJ6b8tCFtRG3sBM9kZsbxYtvirIoc1KmTFBtHqxGP
pqR7PTrGUdw1l6XYQpxmRKUsAh/1JRQw4iNTTm70hejRdiLKP++biMyXCQojX5OqhR/yH6x8h/+R
Jem9kR0WKSGA4rZ6pFuHYozvxETqSvY1A4fVnrelEf1G4UF5f1kFKgqZVjUTeDDfZBM2XgQUDh/I
6Nf3XN5TMrFeKvrswJ6dCY0dFF5jZrpA8gOC+sutTcBPO08+IarREO9c+z6J7YrxqGJXIwB1sRYI
fsSbEu0UGu838ywZIOYwlTUiFVfwJZu/gq2OuAOfrplLHlb+/ICiZBWSf5fDQhZvc8NU11Sd9Xrb
nUkw6bVZGMOTQmm3mLdZJlrd2kqF71LaiYUF8dQlJG0OaWvQNPzRtUmtuj0o2ir2ODhlk+2mFXDG
PDQJRHlsC8MshBXrANZcAync7tyDzLj9qwrVpfVPzUUxP0it8/2KTlR0bJznTBmAM5w219gTxAM/
gZ56dqSumszunzroPpqYth2Sb020etkcJ3qZSF2pbI/qTVczW+3poQIMnmKofYwWpzD8vAnAzfFJ
tywKDXRExxUtFj1VDHjG20tU2eak2qaEae5rwSasA0UVByLElhRampItSCBk9a4qgjoohVrG6O+G
PyCs1h4sKx8BM6joJ2RumWyq8sbsvEOymsz2Qh0vT9vuc1xyi57CtYMY0TBKp5SmvtBFGpLA49rf
V9YVUDlpXdfZJ7i/LYmRXL2dTrsrjrZCfQ2QqdSVc/jwEbnQaRM6Iidoy5GjI/jcfV/IdWmubL6r
XidFSYmPesyveETLDWsvvpc1pXXaZUWI0S3Uoaq7XmFEH2Uq0XpW0bOZKgPubesZhfS0ttA561nR
Wl5ToPUDtDaTYmUmGzMYVD+ORKxCsBpB9yPBkFPFBZvkd+ZlCl4Ya7pjNReGt6U5SL5MzVOiCgtR
wlVAGD07xrxlFDTf8xQXpUoIIH1YYzYaVw6IPUNlmSXdzIB2/sZ6K0z2t7MorointchoHLJWDvXY
iGIG4an+p6ay3eALqRVU8WK2HS9Bu5aXWI6bfbWJ4v5bNk8u/PFkSIiXq4zOh3jUkWyfB7LEN7tQ
WoGvJohm5UvK1R4B+QxeqmnVPRONWUEnmzcnap0BHvlSUea+bRJTA1T/FRyDQ0Zgb3/rHmuLWxpO
Z1FRd2F7QfbStUWRmc+fvtNIdxgKglHSSiYXXtqL6iNExt0wrBBwL0v7rv3FAlsaOqhDS7z5WMro
qgfD9j6l4tvQlOobM3e85CNsp5/Gygo/29y/iyuEs+ejwBACQR+hdEF2nPC7XJD8QlDxnGrRyape
6HGcTZ/Jc/MBmnIeomLyPJYIGbHSDV6WlNtYiWkhM2RVy8m2gjwaf6xkSd5U2R71bSTzOl9+1Wkr
Tep7k586b/c4hgKEASeRHKJ2Y/4tMfhR+4UTuNn1OCWoOB/HKrX4Icc0HS+BYEWmptGZavcQWvJz
l2On05ORmlINZ8wBwlhB5VzP6ILVAcUXOcz3z5UKcycidiS22aQb1W/RxC0nbSNtE3c2k3H1gu6O
0rIMZHeymIPiRPhagxD1+7RMReCzeq40Xi30Kxfy5aje9wK8xWmhv9uUFPVPzcw3CF7Sw/9KVxcb
XTiVEdyejiPs/eioduyhD0znniY5MKbm0pT9GU/klYOyD+4+OXowppn35yNs1khaoME9Cdc+5/vp
FDyY4mFoLLk7CC49TSYcQdzGA09KNmKdIlh0KrzEnatfvn02wZY+ogQPVv8GJvXuPz3M5YWqD5v3
qbU+4r07mBQiMoTa2W75+swCFF7QCN3SObzNmcdj6dfwxyDoCe+l9x1kJEN6yHnVwLO5XNte/1m+
rwHz5p0JChp8EiRYbfxxpGF/dQeFm1tts/iHtVNrKlOXQpsR5rLpEG+N0QBHXt0rH7Nh1S2Dk1u0
tyP7xihB9ER6hddP4+vBF1EOkzF1ZaIO1T7FpwDY0mnzFXbFv60epCzva8OuhSUeKG9mjK5YbShV
x4N3omsdfetDVxx/8NBuYLA3HFMyfEkcBqg63HTMAWXbgzCABZZ+bPfxFbJwMF4hfxjAYUnSqm3Q
AKfjiTqQBLBM2Y66ZajfQOk3DksmhZNTXLiOE60nWcn3Fdbh1uNIILnHZf/uAotx+q2M4lPCJQSr
SeDeBIiqH//4MLfHjbgMD9bWiOifMWpdHoOzewZuekpaKiDgC1YbK0v1fL2WEv6ZuhNZFRwUQRQm
Wn3tSBM69r1/sjc1m5hL7GK2wNX3ouDJ9GamWwVg57QhkVTQj5o5/tiGLGA0yt5tIkmXYH5DTvGk
mvbWt8cDsgXsLQkzuMhVTZUpEGh81qNeFQrkujHye5qEhY/1DFOkybaFFb1V1rezzCWstUupG7NU
gvEKSNx4hjPXspzo7jf3sjSUxTao8KYahNpCNHP+EWEwzqJGhNBePUmA2A43w9cVeXrSQydV3oAr
xjeVtJFXh1T3LyJ8tKZ2I0qzO1i3R95qpOrgbx8DX4ZJ3tPBJNGfws8pvuiWdLIMdzzbwu7sFLlK
Z6RpFuMN/LgL81uSkZTzi9ja1hLpk32eTc/fl6U+4A98TV3/IoAY6YeA5aAABOIvJR1uCW1BxMgr
pLPHwUkRDQihAEIW1M6mkwfXpl4LAAKgwA1q6lVRs8wlpijQSxBtxxopSF/U6AYchufa/0hrdWce
xu1b3sXE7g51Hta6w9h1g7W6MC88MVrjY9eJ7oUWxr3S608bZ0a+WK18MInwDsjW1aZvyl0J21TB
lrn87AQHIvBREmdgfox88Zw4qaMXrArK/tyWeTxrs4tEFmftRTcrzBOz1WoXZQU+Z5esYG2f5YEX
7Or50jpheJQxZDvcXim8QF7uuyDmh46mw+egjLIbQ2SibfzqBZb50MN+/896Ep4fJlm1JKP8Z2mM
+p6aLvswlbNgqc18+3mFOS7aTHqDdFyGcTj4D4U+u1cvGknNkInyD7SwxS9U1eqHChirLZERznMm
Uwfr2/3dOiPhdi9VaLtEa8HPJWCdkfnR64rQn9w9D8HCRsv/OaFjCy1/lJ+gBCRNjksvZLSaqpeW
eyuF6R6OB1+nPGwwyXc+zWm/10xZ+HeJ++NIgZ56eeEi7lMyBk3lAF+625H40ujik6wUEzA5vkVb
sq/XDjDDv3QHiufEoZnro7+ubP672YdQyerhQfd4nbRgWb56lrhxARD2YNXKp9bvWmLThNaHhGG8
P2QKkXiCGlwBaloIDWrkTY37Nty486zw02/vmq58dhs2i+WnAKOYBkCwJyArWlZD5EGYVh0mboPF
Cx4vZhYiwldRZApOMD3GAkFvT7otsPUx9Kmxxprc6WrxQLtWi3yVMvB97YqkqdD2Ah2+e7XjWauS
dRG+LywNVsNoATjkXmzUmtZfyApwz+IslgopkTP+xLkL8pr9BMPVMjg75Gl/SuekU+m00xm2Iw/l
Lh2xmEQKJXeA4JPkDQk0qeu3GTaFsJ6cYAwnqeutYcFb5GWygNoqqAqUuczJ3jdEPTEIoNEWATMb
Ho4ArXYusRyLE1jiqQOdxFVaA4a3JuycYZ/m7q+tqyJza2WG4QRXMP2URl2goDFFSRi4AYQYzvIP
oh5t7W50TII1rCvjxV8rzpXhWqEwCsdX836TmvnaQekaFFROhjMc7sOJDPNSsm/8rjonwhcJ92os
ivZMoOptYOS3n8Uv4SWGmugZ7Xg/4YtQtm8x0G8Ulc1chxbH8WoQkmTa7KQ66SNuJdG8fNA0Ysht
TP9rVsrkDH9UwXea378wGQoP6G2zATJ7ThGTjM7w7sRiBcrBkeYcOmAuPZNWel660xyyneqRUXx7
NJ10CC0TS4HbPjDFM9n/lOmA8iDijLbkGP64DNwgXaeglVM4/QZMUG7l3vjwgExAV0im5I+jxYF+
0J6zvNeAg0INufpiUXHolW1RsCSukwAgr5MEQ0mrN+EKcRQ7u31FOnTA/MKKktg+A/241RIwNV5H
rLKhuUKDvHyyrXsqJtWO10fgTQeWJvVNP2wLEzIWhOq3Wihj37lZ7KOauplp3e8EhJJs683jZOZ9
ak6YsSVpcij4m1kRPE3RFtZhaqmrFOtK5DfAMxMtsVggRM8LMAg/UDi168G+jC9kl6jx+Al0hbiA
bjP6s9/o4QE8IhQViUfZeLrp7XEFcsbixnpY9TRawQQm4264LrVCC4poJFHERTvamYh9BUN2o0D7
KnvKevC1s1/RcwpSa34pe8GCWWldzPD7rKj+9/C5jTnaAi7CEQyJl3e6rqEu1d4+ZhOkfYplz3k7
zvX/tTHoD6w4Op7cmWaLkmzyivfKf7wzSPTsWBJOBOe7iXRq9dF5JgDRHnSuk7CdAYVXhAUFdv0v
4EhXm8Hl5Dsv1vO7x+xhnZvvO935pKa3DKDr6JeW8hSm61xrcvKBPUqYMNrVuvJUM4b3JQ83ommw
xp79wt7H6P5zWdh9UdDCxshLI02xI8AR7hUGKiUkliTo6Mucj9zXdRl50lmlpobErYX9rJU+mDJt
6c3TwqLs0ekMdXLbTVuC02s6caEbpasius79IjZVuDR4Cflf9iRCetOouZpH9mfK8xu8IWm/cjsf
V4midrLRJ9aGZRN/1ylh7Vem/TRdidfAAXidsD4bndmiJKkyMaYNNEQKTj6t4JEEkWvurWTr9eNe
DIj/vNtNNIWqXCSo+9DlYm+BnoNU6UUfAolgWJFxG4chkAAKhooRfdnLXWgfVKhh1JZC8IT5gzIo
l2K+LVhNYU4Ah3Ii98PWlm2uKN4Tq9PO/TGbFRAmySf6m99EEdNX3ZfT/qt0WRDtB+28s3GyJDas
0F2y4seq5MrQijs5n/97ndSW7NO9sVXBJBUTSAJuGl4NX64vc6CNui8S4VTd/nZRFwdISa62q/1K
YWA/kqeClKck/fhp5pysr6OOhwF5UuCkK90n+QRzJTMUDNlnIZf9gpEsXybKLrUyE2YT6mbP6Rji
gD/doUotZeJnAuordJkaU4ErweF8qa82phmIBZ3um1Gs0nypRQUJHPJLgvZNjJA1yF92dJKVoj0k
lKejKCgyfxOdLM6iZJ6eIBKATR0RtHFl+HcKlEgs0gVPaKsa3ssVF3ICyuZZYlimejuRDoQ2uBFF
wDm+TYLN+zSJyqkVnGvyLqXmbplJhu6khP/yKwKFtqcFTY4elSMUBsBM2S39xjZNMGSXwVCZPji6
eFKYMdPo1+xCyVwQ2iiKveCXWXyuLAOfd2N5xtLf9YwF0gHnOb9aNmuiSn8hL0LKxW/dqj7XdEgy
7VkT4v7ghWL+oG/jKxDu+yxQUlNfB8EYFWFWfujN8i2e/LZlTNf/Lo7qPfQtZNgpTiiU5x51qNH6
9Wj6KDKKjxzexskGJvyuwv1oLEYFpujEFtqJHe8f+0r62W7/nEiPP2ZcXLBEF/FS4RZbSjg98XM2
o/xNeU9iVwWMfRpVrq64jsR6STD/RcDRY+12JOZd+HqhOZGpaXny16oyFmqba73MTL0NT1V13b+H
1GFg+foBwH3Ei23lM7ax6HU436AONvBBh22PVDNNk2BWqxXytr1APEroxDp+qbqaKbXrkVS8zVYu
7R+yd1GSDB+bSRtH6XoTyr3DB+zzaJnmHndE7eriYxU+a/KkMlyQlCY9qp1I7tql+yhS7RR0O4yD
8JKp6IaYmeLEfuvwDuLqNARM/Qvx+E1QEEqdPm0qG5BQydmmwh/HC938YjZo4n9eUGt4/RwgVb/+
5QWu8dqB+M6Ot03njQ85WckBGmyBS3QkxUo1eKO0+4K3XdUD1YEYR4Ko1+iS73s/w1ma/ImmYdm/
CsqxKQh2mVYj6Y7YvKpLWvgB95nbhkZCRZQ0OCLj4saHYlshY4ED8ecpZ+CWFBhuYntstMlqr+RN
POPNylRKGr+2jUc9xoj5505qB1wpUvapKRvmJQSFjvZIpBvQFUV+G/iOX7J8K1qyvq4JXUEMa9PA
WmgGAtSCtbTm8ejQWFzcSXvzQTedw2NABydEX2XStOckQPDhcWu6v9JST1qo/abWfhqjabtVZU6l
AmUMG2kvdz9uHnOIl3FA2x8jfoWav2xlPcuIMGHf0CKenojtoVR2Me/oXeLnExUZP451wlhkBAPz
lKgK7PG2wQSkMOw3uTmZVyDjuKyg2gBcyMrNj5t30xEi7uaMQf4CycONN5LcIPwxmHespX/s1ocn
7wirAR5zLdVurhoh5AzftUJibau7KomznnCJlJVluQpMEYO1F/XXyqJwnckBCmjma/779gJpljiF
Zwc9fkiJc+zI/8adP+7/daFls5CHjvDoHJkb4EUO4Wdh6XAM8ZETjjOTZWPRCGk5OyAuQBMsEhaX
BLiR4ZCRLO4MqjgnMD2VUr55jMBV7u6NdI4dVqtCe2nx3V8/KSLIU4m4drz9sM5e/ULg2rWh6Go9
2nIm9cf5uKS3RNi80CINSj+Oq39EY7G17kuYU8hl+LQpwJxJ3XF8tvMH0NoPO2bHbm1KnUkWoz2Z
ben0Qy10WGX+VxiDKJym8KZSYSrNcdVBKvcXVr9SkMSw+I0aF9pkMdvRVKrpsGw6PXQ7kFVnCmdJ
nZyAfgMYrN5zkO/ViTBfOS6H9wiXF+2RJjaaNvb44G1YSDsMIEluelRb44tqCIWmldBfOGRtwXEB
c26bgPr73bu6Uw6YdietZX5TSMYgDEsmH7RUsN+v06KOShCxID70n1Zy1sr4lMKsLFRnMmZgItG0
0CRFvIbgETsTLA4xFE7QC/C1EpJbAkK05lIwiiA+wTye/6Aqdt48HX2VpS8xlZwPMIUX7mj1A4oX
3dKVLZIzsTbZInCeTIal+tNU0wig0ZkUMjIvnh/as3lIotuCHxwMW3IYGBfbXTNdlJ7mbcoqfkn1
1oHsxfIGgaeBdiBA+nddOd+8i11yWdG9ARfpcBAWzEvqkBG5+yqw2XcWBVj4woVR/x5c5mVKMmof
BY81Gd7iVmDiGhXoQMLA273DCb2RUUEddKekAY0izh3PNg0o/kAbb5x1jwkR7yJ+12stUlL1VeyL
YEglWVOIs0876U5uKEVlhpNHmgL/HkZp7UaRdRC+QjIPE6FZ+celIiAS8KM2F5OI4qvQDqSKKaOW
EWqbqo4p0iCE2wV5/gX4VZBe6qxZN/pcinGVZKw0xu1VOSsQgFciaqCselOBP2LSVrH/F49owasT
AvQeOoapv6ODkZ8ngFl6Jz13Rzcr8TehTX7kzsxslfkzwnc1613PT5hsjHu2lgktn7KSzbgeK3tr
/rYjMwOYMIYS+5Afg2zfS8UGAd3dw5CJ1ZauVAnqgGPN97P1K1SjcNDMLZcI51QylEZ73YB2m9Iy
fBWBoZBrLABkCYjimP6jb5UINaqj5GpsGR9PX4d3idxM6chO1+e1JfdgYJa6Rw8N9+XForozPy9E
7E5QEn43Lk7Npc8dX2hsjXubvfVPz78Ugw6/cfB2s0ZJua6pTwhaRrEVQErYXPiw15Rf+VQOg8QM
X7+3c+lFEl/tApjSTeomB5joKprbn8L6kiVv8NhuSv7vl/iNdH3dgLiwrrFZ1iExY42DVg1VP+hz
UaYEyCQ16f/v9UA2Q9IkwpgW4CCj7wlbpn0ezBmu91WNEcq1fGTb8jMCSTrVTNOJgU/d5c4gfoeM
t+PsIPnqSrYh5PjHwXeqIEOSRp354LZkIazY2+WXP3z9gx8yp5amnPNDlNfhgEIx35irS2Qdd/4v
AZ3vIz3pF0H08eDcH63V5sS4IYWT/fj9aP//5Lr0dw328hxBslUgzrn64J4fCzx7O7yYR0DDIp+N
063xILqHp7nY9wtj3ln8hEzNBs/Tg5FdTAviVgccscVjSlDWhWyDWzU4kM7cGo12Ie/1O1Ie3LqZ
/dMurqmfwp9Xj57Pf+K4mRIpv1YzTRAL5unE4TJGbPrOb+ebFVbXiZodybvMFooPpOJ9rYCPUJSK
49CF/us0ApSF7Vc16sTuNiElbc4d7IJknpXPB3Hr1NwXgJl5TI8YKv945mMIMYCBpyUtcMUpdxm1
y2tiVwS6DLnYqbczjUvzsddlT6Ik9ceNiDXcpWlpQS8Jo2rsJDP0LiYqZI6GDdkuZuTi1EN2Q8cv
bnhtY2eCvk5+Kdii4VS5QU7xgSpX9OPA6NzacTiOLRldGv182VsnDJd/yFd9MEGE5/kJK9WQEj4e
YYlnmwC34VsRm4UjT59MO0p3N+KsPYO6CcmOr3LwzvvNt6tUxD7yfycDUqa38fVCfNLmjToS5n8n
TqhcDWe31X4/N+Vo2Q0mxsNqGWK7ZHVRKXuqBWYKMKbN3f/1advMku81OVvF8pHTQ5LuLl2ZTWDs
c9GgsaayPwYkbCVwqgtv1nJGB6/KNh8fXa/T2+S/vQS73ZoEtnHhKsWJ5R1nj2uSSNlVwnDKzrnB
608pIOrxl4o4el19D9rlEux2dwIHbjNlJKgP5+FQ1jFHh5J8r3I2XvdIOogJ3cWrRgLlzr5q2zcK
lSeJ1ncX/Se/SdzXL8l4Mtp66D1Y9bzuGDtcIaFlCHXzH6o3xE6XpR3TVXIZ/7A5RzQMgTB+Q3nm
FsqeF+rZ7gNjlc91W3RdRuyEnRbrQFBCAJQOjWp2skP2Bt1lcfq1UsBtdsSiYt7pnV4iVl+XcUTR
QCi76AwwLupM2zDcAHYzPF1YI3Ss1v+mDsgAY7aS1506iypNlKPSUsORZnQWPUsD+KQUrOKhdNUu
2rMmSB+4bRWt6h4Aea1e1ei8LXgWwToa3gWPI1vTBDHoNeIiNXCj72uh2dQrqAYj4Py0uWitRzGa
FnuvzRAzrpuQ0iPxogtGvaE1rjW8npqN7AkShVvs8COob4tNnQJLtueTJbGVPEjuaIQ3PnKTe+rw
fRe0l9Suxs7hfUx6q8NqZREOTkpcDeWCyi3cTENRnVjk4zh0iW054Q0OKBogp5xdmJctjEm5Sp0M
KW33kLnUkJXt6NoDDPN8EkPFP6o+Pk7v4uuLYARIDPfi3MJFLIvIL6R0lznpsYrkCoF12Ynpyd3L
h1B2F66QkSnpyvhMhKuQfOblKhYgDouXK60FJdia+eV+HUThbXiMMnY9/50uLNkuXJnMghKKJ7Px
dcvJNgM5Rc+OLcEcEUsdEt118iVG+j6EIYvxwpmifOqUYtc7ru+ZvoUIQ2CbYQ0SMVUQHrhUK4zx
0tEW9p3xQ693RJ+XiTELH2lGnvucLbDRhBIMii5BPR05bxU2qDQ8vvge1HofAzJWsMOSL91psjHy
ixCCO4gv/SKQDYmsrd9nwftXbodCzM/dKDQ7MDLW7kbk91prOe4ReigpKc+3IQ791Z6ATL6zeCPR
J79WdB7fZJBiVJIVBn2I9XbJUDhLj0AxtV1GmnzjxjvMZpFy2ZGcCly8Am5RV7FVx8/uf4I3wEe+
IzEKaA6XtFqrfJIRWbF/CJXTEJjiaeR9g+PTkiDCzUfxkH+3QGs69SoPjf2RiEbuc4DkQ8YCXEbb
BKYmQH1WzzCQ2RpY0wmV94yKRUT86oW8stqZUbHk4xUAKBRXQkeieP66mmMkYDtQa3bAb2v/OfV5
ZquST8L6lttSj3vtJBHgFTSEOrizkxe1PC0dY92ny5zgr86uXGymFQJSUcm4jNOetJqrsDOkOYoQ
9BBUMNEBrFxP3ZHxyWRwbgBeFboxSo7RsN4gJ6IySWt/hD4eVDb0yTAL5SXvN6Z4SsNhNiOEiqD1
u6gp8bJoj3VQVi37v9X+nDOWRRaS9njVNQoe6YIZH/XenrM9y2mzKpyb4kAS+sGP4flG2uXang3i
J91fYlx+CQM14f+k8UsuQAKZjx58fAEGZZTdAFLD9IARXYddVovfUvi86ROQKhZQ1MyAGzhMRFt4
urOaVzpkCiH/+WXSy9gVWsZQwVtkfgw79snyxVG01RjED6MhyK7cDdxWchgskwX6w26haOjC10WR
BD1TPq6P8BFLrce5G64WmG57O+f9dvU0Pz7QwcWf1qg3+wAP5NRJyA0gnm9HDL+CLQrH0NL3nyNi
hKzN4qr7rp6fqFnCG0e3PZqohXWwleVMc7uGr1WxQO12/M3KdhrLuxTwKCHF7gA11jgRfH4vObTK
ySJfWmkj6kumIVuuq0Ip5gQR8oh0TnqBJKlkJifdds3DU/FWR8iN2YcVyhEAnL4DoV/P+waqOIC8
7hzNpedjpyZGiFf26RsSuKgrBv3aptSX6Ni8ZOqwr6KellYRtnxYqoPGjMB4Ue1sgay/QhiELGkI
/1Le+VO7+v3aUBkqdP/oFz/teLTuP5NSXbfU13va3AWbg2p9cyd2QhZjHe5rl+rcSSf3Rbq/x7xL
84l/4OE+dUNnO2uxz5LTU5qGa86IyIl9hlz7PH9OFTB3ZXc3jx1JdqgPE2YQL4n66KomlwKDTRJg
p+WLKTsIUVLSK6NoAY8v2qOpL1Y0Ukq2DLz6MAkmPAqZLpAU9WECQ530VkQtefjH0weTtWivWeYi
2UezC0a/bPzv4znb3rV/hjSdkOUOOrXeUDGSU9WSXYjeRbHo/NWDmxZWk5/wMB5Z9pHzIYD0kqJm
fzUQ3qTOVfetGGnSDDahvODoMmhrjJKsUaFoxpCqC0ZM74FD9yp+dlJOkgo4SntQaSzurb+t0JO+
5ADWKiFDCnc0kInsBW816ezS+MM3LcORB+3sDjKTR51QRq1wrKHvuQlfb2IuRsCYsxwgAWmzxqr/
HDn4pfMK9CuEISE/oTeGQLqW7uaCWeZhDv+KNlIe0ZutbLJ46Ka9A0iTnRHc9+8M5WYftAeLyMyR
Kx51dEwZTu0Uqte9uqpr7z6nGSj5lnUM/PFQnPPgSVST8frNjTRn2CjVQBjC2S1/h69e5SBIZb4p
1ng4Hb/IdqwHLT9di3TG/DgCvpzIgwwRxuvioCPXFHEpMFhy5dYqGYMq2bNDesL825PE+a/6HbsD
wOwDsIeEPnK2b4EGMnhJ+QTG0wU8zoKldt0RsbyuEYsMVKNj3WenSyEiqTh+9gX9UjuHdpPA9o3B
vpkoCCs13RW3mWduoN+JOq8HUpf7R/D8QFtTve1Qw3gdQ8XLA6+Up0uf4m3f4+fVP2vjbkWg418v
nSqT1HFvA+NIMkOVjLX0qPkDwDH0m0Ha2TclM9DXWz/pNwOTGbHHDpXxKGKfTDSeXwLNnwJMLeHz
gQ1RynAfcr6MDw/oLGWeQpcZIYbt3VcGxOvDTZIdp8Ql4yz5s3cxed5K15k8/2AkrgjBSVvmORzB
ua9GiW2Qa1X8WYYlxoJUOJ3FNPpPSd/onkd3DwHHSj7gDFKt3/EW3hsvfiXkkEWotOQbDNTjDfYm
0MFq4ZlRzKbOva7FbFiAWGAFzzOoI2rDK85vWvti6m9+45LJ6fD161ztVuSQOtyMsX9PCp1p5l5O
zeimcsYDkT+g5rbZR4Ubo2uSinUY6EAnQ+VRskwj5WYNt4AgvxConyRIQAV82KZu07ebpm1+5B2c
IWIW7G1ByzmbXQFmoHI9oyc8eAomQsfoMf/VYDWuvVRO0cIujgRA/WnnDEtB5Oeuu20nzk4gvUxU
r/ismD8nli1nUf2YDG71KQQVA8azhNmC1VWhTzfI1C4U5C4ervZotptMxj5QlZ2G1rSvGAB0RWUW
HLVx6xXDRuJXWFZwYYs13d9usb0yghIK1k+PqJ+3tiyKApL+ibo1A4rCGp/MRX/cFXpx2Z2SrWL8
tBhg8ZKFct6C2Lt2c2lBNApO1qgiiw+jnK6Q14zO9n7YzC4Lx8FpNE42Ao8obKTOKWuIYTyO/om6
O42F3fWNMqIpNd2U3YGB4HMCM+jQSL5aL9RscAvqNQqDGdHjZhDqWAw3bUarmsZKnw13rytdCOgk
0zp3XfMZUQ1JJlIZKnvvPaXX7byDbNPlev+Gd56jnAs7UKOxwcKT53mFZuE+QBUGVY7T3/IPFqVx
ZRNxx4e+0Ion9+4bfbB9GXX43gfdQQzhwqLpnPh6oi3i0uvw/usZHicwB5Ds/zmMNKz4SzIaW8M4
iWJhYGENkbFMRgslqLu8EADTjYRMV17Lw3W6GJnppYn1EqaVkgQ3gMGD7oormX5YPHfzHPXi4sLg
xeeS8yZkVnJuIIWva6b4thU769EjNQqi1Ab6IZ4S02WEB9Zw/uEYdfCv36l2sko3v2z0Za9/nsgx
bQL9SWBRPJCOqIBRHc8xtf8Uw95MbvQ4BXzBmd3wf+QmAsYfptMvrM8Vq1TWN0gW+Cduzs6CNEru
FC2poj3D/vOso7nogJHPMuM7rJ6AMAZ9Newr43scVkW1uIbR3xcDSPWQn+ZuX/8g/2iaF3mV1kp4
fcwcq9j8J1Sn585DCfo3Q8p5Nv1pCzx90LNTROnZLbHz2P4h1nIeChzeu+nnwVu0zi9zp0Cp2lmE
Qqi5L8TTfkT3V3lwwgZGupQRHFq9Wt1bb0JXBPY2L6Pby7zZLNs3ic2vr09y9GqikuznpvNb6fAR
nqM5otMKx7e+mbfGxjVSPZPLCguO7yO/2pFqHtP+D9XcHvoet28NVHxZXCY4EUHDWJ6WZ6SDTS+d
VMMckB4PRTkqjEHdkKkgod69u9qmZSMWC1TsI38GJt0vtwOe4RyYErT50ZvYDyACeQykN/J+R3xt
TXRseoiLovyYHeYMSSJ/mOQsonx7Ad3qQIrA6Kt0UlI1lk6kEnxvlFzy3FdU4hhKkcXEqdWBs/fk
Fufgdc7d+U/9OCVBdyz4j08NshkjgQWhPCzwWAqPmRkFiwm30qBRUFCwqns9O2Wrpbr54r1nM1uE
PuXB+ev9UFnQFoDGXrbuHyv1yo3ICRd9fGTc7jqxGfeC7YFYU/MvdishjITjL9vq+hxsstdtSifF
1ThG5WSDnH0uv58YqGfXPeqsB7/4KL8rPqZf5DpV5AA8eHjLw2LPGYEwAHwjp1CHrhXlOwlJT6js
szKQZgdaVE+Ny6s0IzDOqVIEuwpL7DCkQOpB1GT+mao+dhk3+E4I9OCMAGSTS9oNkjJT/TAkP3Mo
kwUMPVuD52X3QNtOzl4S/bJI70tLZIyEoA4rRSWkZBVBGPguCaXsxMegbBj8vZeGXvuVUVgusXy5
dEPsKbKZRaDy8RDkD5sc04Z2h19dlQGk4rdVHuYJhRsUYWAXGZcOrEfoeuNGz9bqWmVLuviD0Bor
VY+iP2ObmqQFw761T+GV8AAdDdyyH83DQN0m3Wr9+ixOIrbjvkro/hmRU4C7t1F+AA+oP51g5DQx
GXSY7jr6mRp7Lv/7fApOCJOsQ7QRUHVMmSoP7+OM9lUVQlDkqaFPiKoUYUePO4u6qjzoEghjn6hB
lvhC7JfV104S56qQYie7NsLsam3gpRyA/JAVr39mzm1unsX1Ox5Im/01tgIQmMx5xbwtJ3bPUhCY
ltdCNLyT/GaE538yv900bm38Rd/hXpc+0lH8Swhbfwxom66kqf6TlN3NAFs8c8GczJ4VUTN5iOeS
5NkTe/ULGixKwFkpZT8EnoGELOUdsy8WTngvxLzynqng2efWBn6QoquURSgaEKEbB4jZDTrzN1b+
P26LpXdrucABW+9fqK3LplEMIcIhknRJf7QlpDjVikDKb/dr15xYxmBqFvXmiBCPJmt98kR44gCM
Lzh2twUF0SRhbDmt/ixasWqE2NCdbd2rSciQ4yJJ1xCmbZIKG+zqCQ66FZI/epghhz93Ek82SRh5
nhleoXAsrzkFJYX4ASjW8vgjizfJqHlPKsvlJX13gfZOGN+DsVOg4ANIg1YDuZUXcAx800hP5VaK
jurzJZqobgrD/IpgWuIoTRmLcjKdABHINe7xWBY1ylkPGdHpBnMCsWO/uEe6zELI5IRkstXQebJK
QUByKzx78rahA2cj7L7vVZPLpz+Xe3yeb+bJCzuHHMLDG3q+zoFLsPoGQQJBnaiKei23z8jJ4C4U
xQbo9mrxhtMz1Xv7ZEdXQR+JRnNNny3x2Kabk+Fh2u5mTFx0xzx+mes9C1QFi+ljb1iPlHyupDad
v0HlkqX0sT2Nm7j+U4cQXMED1THoXBw3hEhHonjF56K35thw7+wFnfcct0QUSA0LmDz3AybdEBvL
uKMsnF8TIHJ7IEBRqDJH9Vm/l84cB5rA2tMBE9cqU9B+HdDcenQ8XKNi6Z3SQQH7wD0mtcfRah+3
1zD3Vhki1OC4+cNI1Zbc65k9GUiaA7daFYSX9YC2l8e5VyD5UCUT0b15Z4+L3ueMOrQzrERFMVUk
VbXVy8oyEXjB7RGTU3Z7t4UBls2oUmhbvm66J0/FbtahzvDTDYXMUOdLrE6AXtF8aixUBPaALLA7
S+ajnuMR52IBhYiIl0RMqS/gS1peM065bW3O/pfQWR70zd0n25s+mfPBZetpbrBHY8UJNY4aP+2B
+f6PEWiTqsBxcNZ7YAKf61Tz7DKvQ1hoYwHcAqe6ZRxEVB4W1xWa9VJIutBTD6Zo2ILlY6NQJzBz
lidJZJ9ZP7XkUXfChKyEmiLgAlHT0WjqWv/t5x896fasjafVUFVbMEDxNo/GdiGsD4EO36TXecY5
Z+rZKkhy6iWBYLlN+Uthj6vQ7aDoH1UBNz/b5kudFhH06mytfoYo2cHwqYcGWUnyQq93aHtA/Rbg
m829kbHCioI/Z/bzmVJRXoJiLDuebnP60rFLUNpwVNeFGK+TbO3ESoRTR89dFs4U7conBNM7RRzP
reJki8WXd3Smo807+JqzZN09+M8DxHnFimjRTZ+KW7ihFVKIyuc8h7CktSO9EW+XU6jliAB2TY6E
yIaZDERXCkV6O8Ox9XpVFa8suw2mSyhJV8HeUgBvuLLCkjVbRQVGSL+ic0R8A/i6GA6xY9XrUcyo
02CyWI1QvkoLzGRFs3JNUUNnsG4wDv7u07csTBR3aXGPnhMLqOna+VUixsGhcyTkUei54n2DVgbf
UDY1EDLL/QR14E9/8OUbUGVT6kVaaSyEd6Cvd7oZp7pMRVDUCAaQgV5iknYuBlvAJ3ZRIYuEwghL
esYuEEkzf/q4T9vKRdTUzWUgXOYGibiPJSpIvNnFKBV/lH1B97zkm2BQTrhSV+PFezJ6rkEl3H0m
03+WnmGxSTkyr+ZXewuzX/FYPRBw3kvMNaEB1/inolcYWn2TE1h2hMUgty2wi77e4lYpGxi78z8q
DUM+5TPGjkYMMJ5iODaWAmkuWYAvwKBLJRQByfYSYe2nxnhxWbpxTPGjRLaoTU7d9A9MpqfasPZP
pEwNneJ6gp7tjmXzzvKuOWCLBs0z2dEjqGrKQjfjLrtmOOCowlDRgynQdhWlcKS80npIKX7JyHdv
1yfbr4iS5aqpX7jSTx50LhdRe6J4MdN8jfJCMYXkHxQbEAKW6QKBgdb4mCK4v4gLRdLQbubNt3zH
U5Pqc/SU1oeQ8Lfl/jwVCyXxyDUu+DtLFqk0c75sRybpON6l1nYzgZXy8pnhbZ2c9mACyllOrZs9
lOMFBwA4zu/+sq0C3YVyaFHR5SMEi+e9/LfjZJj1haWwCEaV45E7dgimE/igW6ToYcKBk4XE6kZd
IIL0m6d3PQipa16mWaYvZNGRiYSMvGpKiYztMjpqIseMeYhD4R8Jem31Q66tTJ/gNKlhyj4wtWqx
0+9L87Asa+FgDu/vmvia7TwWDphh0w9O8IBS8HAXshWQvbkK2y86td6IV+ifJvc/51NFHvL+XL0t
VV3kAv3sXtDs/gKw/8gHpD9OnBpdOIr57Px3WJk3SH72kudGMcmccoGlZtdmj+afaOimva1rGhm9
DUsVUBQ4GBXrcH0fnOSlNv4HTlG7sym3NXpm3TY1PvNnY8bxa+5IX21Q3/+8Z6dz0R+AI3tdd5lm
iHh3rBznG3v3PoTYm+OF7sG6Oo1HHh8IXdVmiN1jqk9yY28lj3B0ukoy3zy7xJZnSB5rm0wpw9fx
0GjFJQS35iiCrHaV/8kCGpNuQ+j/Uvq97q4BTVEjmc3jGklELGwdpGChhSzmBzx2BEJpDNSnZXMR
VcaYqdHZZpRrEXdzlKUd8NNf15ga4ID38HTTNF9XfsbDo9KMhgG/CSwMUqfGcCModqVcBNXM8A0x
/63GAq4kiBPfVk0BqYX76xnYIurWNE+6UIKM2kTpWFKsrlHymFBQ/b7KJdibUnlhl/AH72OE0aFl
u3DdUzBhdRN2f9XYkbAMW1enAHSU57UJWpOiAzXJ0QXspye++htkSIp9l/benFoq3aDyi6UaiixI
IfYgf4YQNM+w0Xn2mNKVgeyA6W6ULuhwYqCICAS0AidGyuJKMzcvhkoGy3kEekYpFJ3heSQRM7N7
/Ph1PHFHdfFxM/ltbHq5bL1tPVp00Cpwhn+n+sDKBz6ULAoshF9ZRavW42nMlpCPszLxZH8b98bM
XB4Rcw2goXwYFSKWIR71T/hf40dawAP5LfmA0n8+QgWkYT6jaARxhte6zg1mtjKkEgbY55Zat1bP
f8Cfdgow64WkhawDvkBLOQ8aAqDOSGgfJjCEeS1PeXm6kdtP6dvKtc58tHwgdl0axOtaxbDoWIj9
JOrrVsPfRnKNLcQph6XmZMOhL3WtTWStmchBQkma7EqY0XIiiIXGKoDmfjGn5EaYM6rMlNuqo/z1
abJ/fP59KJBYLdNl09jRjEl6Uq0iEvyXXqWdfn7jfJsS9bQ/k5hG4baLJwJGfYcKZCUV6QAxPZiY
EUWf+czKdRqqJ9XjMVnr8tHOy/JokFHk/QY0IgJe/0AEClNb6x1TgW49VAvVoxik9nCnexllxNlX
kYK8gSNZ7qGmM/otTxdBbC/NuTRuLRdvD//GZL4yGS93+nJn0LK5z6apaCQ9/YDizdjVlPfcgFOu
VHDqj3AmeIBIZQ58l8yow9Mph3FQ9/wBIpgojFro4G6K5cf5IvSagCA6s7hq1iiC0FodHI5OW5k4
/8nbJwOmZrILtuQ1A1OjGV2RUGWL8tpsxRn9LWlftolwOBEOllJou24ELW80n7XUY1j3CEzC5r3F
T+ithIRMMtvjMZOyvZ3QgTHzZal0cgPUiPHWB816r5hoBXa/9xZHkQxmXcV6Czb0w7K5vjifbbhl
pa6I7wi/ZuwCN19O1GA4ShRAiKmiqiyOOHwESxs9NvrRDi2abfdbL8c73BKNpvE0DGzH8aFkznEF
inXtxcUA/3nNJN9/lzPiN4ao80sy8iu4jhSN7uJa9oq/S8W9im4pE+U/KaoazSjcjVsVYnr8DZwI
qFSgxfJFqMimRlSnzk630L8xdUfVTIWop/ezByv4jME931+2ojWOy1aVflN4UXiQNX7xsUKFPNuc
dR2NSs+STkiAfsshIED3x88J8MJTDcdhwUY9SpgorQmDk81j7B+a26AGxhN3ETFRP275FGiwA1A6
XOjePYZax1XYhYhV701f+JriCoQ8HVDzr/+Z6E2Cg/2ZSx3jJns4exLHAI30+3YnOXGlfzj+S5YZ
ZIDH/KT54jjo2LQNMLShHlTNJytlQWOeIzYdtUsHlVEtXa3KT57J7nLD52433WtvQkEp71lbc4n5
5KY3Dd+Bv1j7n6S5dVlqWrSryIqAi0edGmcjqIGnFHho0JN/Of4t60IcWcYnGgtZ+w9YTDwNCmuf
CGwtuEJuCUUVDuYccTx2APlj/7DJde/ROADBKANtuYHuETpFFFTTdAkvyQSfXt732HdrR9Tqh90Z
DklQd7TkBfhZDPrShZcp4DDXoMz7YbebmOGB0yJxcSBXsLlwPFh17lWzMgpoWjcZT45///Mo6x6/
oaBF9lcmuHZNC5lbBl38Ze9NZHUk+cqiLKBKtsJGS2TlQ6B2/9S1l5C6gyyEeC8ZE7/3A34pRxJ3
hRunHz2CPyaEqfgTvaJWTg2XYgi2eprFaiauhB5/wi1NNbD+nzVAW8FQ0pxQgEhlQlRYW3tLoSdR
Qqm8cDGN6KeP0GffJuLax0Z198aQJGmdCaw19W2soP9HB8sa5aMF9HdCwht1ZNbRk5uakXDhUkci
fddj4hrKMrrXwiSUyDrAQypm7LWsu4L7TykUAXj5axhnBauFImNyakmG65kqmlTB+NA2dST7+I99
GlKpbE/99Y/YulXxcrTSxgifpBKuxVI6JhAF18gquVmn+4kl23lCpS9WvRnSWKk2ex75LRVATx+y
jrPpYvcWEc+wS9hVmiKj78kyk9MrFnLp6zvChXy23Kjg7cMCzhtAq5T6hJ0QX0kPMeeyNcBJYcoc
DSSPhDLs+fXKYUHpSktCo/4DvbDDayyAaeWrK/nHXLS7cA0FEkOTb/Ht57POGCweTbH9PQ3adPwf
1p8xbEKxYB6ReIJg/9PQaXxRhuIdq1gcPba66xLLQaghpz16Ic5JAtCaRYq3tI2IXE4Jq2Pt4KJ4
KTkLm3rfDDGVNzIVqhdhYvE9DQzgLqkRJoAQv3xyxuUpi0QvNVoF8csPHppjINMqyubL3xaKi+SA
tW9caVZDqKtcM30ry1VwmwnhnqmwpJ05NSfV4t2bzQYZwBQN1f6vU5pp3Rje8WSfeJ+c6ZZANwIh
ZCHDryH3SAlZivKfmSqS84bSUJj4Aeb0cXZC0QhKENJTMLdrUIRi8G49dk/SK2TtAE+S2Nn/lTDV
CwjDL60/G15ZHwc9xCE3uFhECaecJUBAPkUHYc1gfQ2i/rlVW6v/tCuWP6XIDNlF+IeU41M45zLA
2uJDTGxL0yplW3OG2t1EdwoqkFzwUIbexpO9Ejj0vqyKO2Gr2TR6PlzM/QeP5J3lvaxYPq/4ul/d
jHThrY9/UFry5fzLzdu+Xx7O6tk6GcsT+uGMnCzlhX1yq6NJUBSbiM3Rs9xnZlwQ+HCo/RoSmhai
HublqaW5C/oMtos/4saKMVKMiO9f+dmG/Dz/94nCG7KNZkHipXRx3XHvZadKhVetVXWeA+UbBHck
d6KtOK4hRoq0Z6sviG2dlkv3Sm4OQVN6+q6OWHCFlC1nMXLsnEb5v9SFkZ8dSMX/U1AQf6WoYcbf
AFrhbrwA+KCSg0cYfEozqlvRA4VGXZARjD+YN8BAXlLAi5BxXpOVxcvTd6eETo4aFREbCZ1h/M1V
h9zBDj2hSuUtWVOsbhPGepmZBztWprweB3DwpZo5EgRC1eVLZUSd8kEhUqszQMZGdt9Gzhg5DAKZ
ASJ0BK8GoJFx6XPwRMtQhqFkJfUukgo2pGM/JzUlpS6+1HN/WR39ge/Awo/pWf4Hsi8BSP85puex
Q/Wd/wGLBAe3oWBKyMixWo1SMFl53ZXo96p29PVx/loe+Tt2ifjBKADCz/YFVzyCKoPLvipftu8U
E+5QJsesHWc4nkHcwOErPne57rbG7YgV9aqaHC3my3gNH25vuHPr1oIyR2JMr8QXzZWwzAdpIPv9
cnwLy4NvwfcUYgf5IT3yKPzg6Y1+S7hvnC1tL7bRksZqXIsuvh50fcMg8PA0wcF0e2/1fjvuLio/
Z4yVa7KUj8dgGpnK9ZgY3VGaKbLFGUeWgql1Dp1e40bz/to+Mtpwo667WmQnY0VtOJkAVx1YzEMe
YYqH9BwIBEIXEut/n0l1HU7R3yeO/fyCmzoS8rfWZL/t4q63fgopxlCNz7kemUIVyiu9AnCUvbCY
gCPo7kYCVHRgdA7RLjIyjTFsQN0IppgR7FHMVEZ/oXQoQwxmdjIfBRVqcKNtqkKovU1LEeDznmuO
g1uB18rQkauzhK+gOG8VV2Tqbe+3crVYFoKREjSs9sKWrXsqY4/sR5UtTV0ih5J8lXDkKvsX1QTS
S4CC30UoquqHM6QhRnvoED9I9V77fo82l8XUEYLVbseQY2FUudTqm6C0rCUP6GuXTHoiRv+90Xy6
8Pe6Ls55GRvyJfOqhi5UwbGjLtRZxWifvbdeHOrMNyj1wKBk/D78/5crJj83GAZkfGObyM2TemW0
wFFFZ5v4f0RFbHigxwlKXDhZPSJnf8NTvuI6Yyul7twYKQRSjnBrk5kmNKRx3sHqYsWWze4Ox/nx
eyJ1xCWAflxZtgBrqRzHJpzdrst+q59t45Xpb9wGR8VaZG6Fm6jnLxEHebm+gdUZ1FU9Hs7MfjXO
8bOQ6vfcgeNEweC3Y7n+q/gkOLUDy4e8WZHfJ//nyfp6qaF/Zq/VrkSbBtx0DUNhZI997c0/S57M
dHQ9d32LrFm7EqMQBgCkSrSAu6+93//zQC8VW0vOgPVVj8yhxazdRSnzcenzPE6RpF4Ny4ZR2Rzm
ErJbnaLbQm0m5ZPIZ5Ca4EPlYzQsVpK6nNPjaCQ4LWzXU6Q2OkbWIru2hhNz36y5nf1wif4YW1Gc
FVPq96tFRKUdoE/vtw/xZ3odNZrxqtPhtx6+22rRozeP69nebTtgFtL2fQMOBslgDrV5goXzRZCm
B4TlElw+utI0/WED5hEJCSp0rgh20TU2hThTcaj77F1bsdWZVRB0Gh32fl/JSHYCc9eV0NmTjTLe
RbiGhvdbwQGSTE9XcfbFs6gLk92/FDl/DH1mRQAxXJbeuQaN+1MZTkQyZApf7OkAmBRHTT+SnIBD
h5Y1Ulr87VBbl2+0RRJPXdftfPO5TeZc8c4r1tW2O1LIwVnFqGraWHppA0duQQYovNQaPF/GbcJa
mL4A8sIwBLQj4YPewmgbFpun3ZXoIhWWkRzIw9jfe5oe2PtwdLFgShOrx5hNexZMQFLcIHjFViIx
p+1+QRr1Z/8f5qJzEAbIsdQXgv3mO79qn9Yb6q21eR22i8NUiQiJoVXU4WTvLe0UCU28s2gmkaI3
cDfZvm1h0evC0ZlYTyoKjlomDjWRHHPoksjUX3atGgzIFvmxKpWGp/R/jMkGj3AtrE5q33ndnMWC
FWHet3shkCCNUmS12dE8DfZAHp1sRtHKS9MTp8hNZl4EXw4VmzRZv/Tkey1Uxj7C7dfvd6bw1gm/
7q66C+Gy28YoVTNcqRZON6LXb2gLJvNTiLlVt/fCrgklC6PUew2MYILLyAXnRVMH6wc1oO+Y99mx
PmgVruVLJa8FeF3+68CAmweMukHhPEMtTamZNj1y/PHodCMsvNd1/dPiCzqIsHDziKoZFfNHxBlJ
D8v14vvFvu1ori5vVB0KteXb9WL8r0m0NzNjYt2CzlqJ6R+A7eRmoJN7jymPeFrJ8VPIlVDRxuqG
V4az6rnnu3GQjbJz3dZUExu4TABBGFQQuIBeR0jml06zZ8J0ORO12w4uyIv+V6e0HMb7yTw+BXwL
T7g5iev/wdXSOVzvq204i58hwr4hby/pj84A/wFTVTlVCwfmmE/Muaiz1s3xJ4LdxusdOAJvoEWS
/7z2pxFU289eIPc9HWaEaQbR0Ga+/HHV6tTxLdrN/LXD0XzfVR63xbMZLTayu38lPQc044EBqq9e
VCWgPfkzS36bR92h3lqqqrS2lryC+OM+WiNA1TLaivd/3mFEwdA/CVttVqjbCmfsjm2FVaroHez9
+1RKr2/Aboh85k+P7C82MbDxHiK8ihxVLOSBw4xW6OtbZTCli4/NRkaF+Eic+WZx59FI2QYQbzjj
AhaXa6Oxx3p3R/lp03CMr+uo3hWua9nPC08F0WnKeEUt37somkr8zus/+WBrudhmDo+M9+8uPUvP
OI0D7Y91i8KVnEb9bSuvo2GA/XWIRK/QOqbHfNEAuPYaPKarWS84V0g5FeI/TtMBH7e6f5X31oXy
Vaccvq1JAGi1MV/bno2yN6QHimYOTVoBXFFN6c9wqw5cJE3wptzhLoOhpBaGks7ZeqBAVnz/uoJt
gRGzP26KQhVMPok0RMdxNIrrVisK6+cmKvXGm2Vsd9usuBNucgmzkZgKwTllcIqgtAe2RoLqw47M
y4G5zjXrwY0k3V9BFl//Y3sirKqye+qfU+S6yivPBrKNRLM/VWSEJ68YicUxd4dz0PmmEeIzv9tl
2DVo95eVuMxr283/h7SuNVtWHkTMg2PiJ8y+kZABSSurhF8n7+zE0fyXOIETXtehDUnC90MG6Xdq
BAC3BPcjNy9r3bYLmPyyhOPWPqqbfS+HNczNsRQDwQbgXxUT8dELw0BBg4OG2eJUfXa6/iNLbc8C
MO6t8MRE2cQar4Ce2m+WZA4t+T0CCKYMhvhXEdGQFob8zVE6vqSu0kJ/rDzhwZKkVu62ygSJ7YKR
URJ99FS0AxRgWywMG+Cpvd1H0bJreax08jYtyBBbWW0rMyV/HM0ms5rhRLSZSN333hUjhfdVCyIC
Fo+HhwtCtlmwThSw8RaJqbJzdowYEUQJ+ob4eGHWBnMLVE2Byp8pY9+X2dFB0kos5qbtlPxbBV+b
vkw0PJem9Qambi+GAVOBt/a2koBu4daioend8h3zKh0SaVsgsPH7aaLNNR8uK41RDDruNaHXjXnW
vQmU524b0a0nmZBaCkHP41YhY5xLK8KTLv2kCBQndr4rg5Q5rOlf18+2/jiUHIo8tLQhj/RhPX9Z
64VZwe83hF89roVNl+xbgJG8YbZ2Q2qi9Anxr8a2D4N+kOzx8l/5oCEfrbcDHcBzY8DBQSg/Gf2O
5b1Q1usjlGH1NMMTLyuwC+Q1QWKmnHnSBJQ19OiCrhjzy8RdoRIAGhwBHbDqnGdo8VBzqX5o2wXF
Wb2TbsFzlLP2uSX2KH0OQn7+NTYO+QkJ0UalEQCdmPm+U017flyBwVQR+LgjpSpkNguq+2PS9OK9
GUtnbEr+/CPDMXKaHEIOF0taB1Q7/Cn2mrEclmZY9FB5RRigTyAELisYTNtjW8Ocfd0fUSkim/Ol
j4e3C2FrhBVO+Tydwh9v5dbRbvi0bW4XO9Vt3L2tdihJ1njAvt1gba4iGakpCl+PMfwyR/6l4Voe
WOH0E8WS3Ht64wPAAmlIudR9eylaDkyY618Du7vBAc2mr4f1RSddRUjCl8HkvxCix6tE0VsBnv2O
4DKdEIb+o6I9zh56d/I3aXvH68a4qtFSeaglOoN0DnzTiCaDi2F42VhxkHJE4CCJavgzCKxkMmVa
vj4ZLNqJI8pzGoGDgVxnhS9xF984LcIPycJMtDoI7qWl8ZOWMxcUeus9oQM8eLCqN2aFPzq+IQLz
40Wm7BqmwOojB59HXL2SoVoPXEmn7VSBwOAUUBEhxZiEdghye+rfmuNSCeowfctvCMaru0tcQELw
9jveQp7r1Xq9Yp/gzyR2fMG13SrANkibZmUwJt+j/bBKByQrZt9owXjL1YfxiE/tlwVIOUy8XIqE
4lIzCE3x6bIbXat56smqCe9eY6X0mhEbJ41J1J5HPZtCHJpU+0HQwHQgEoLGzBN3KyxRzzgEhQj8
wCkEon1yNL9MqR9s7PH+J70vs30Drw8ktRBgcb5SfxCDacXwSASO1+caNZUithlnXUzkYwo40oPr
EQWviSNXx6brct4gBLjNJt6HTS17WSU1ueBmfkBhaT6tr8ATSa55SeUAYGHU3MUmLuKGe+mQl4oA
mZ+3vqbcQUL4b2+GNo0jHYUDDLfAHBSOTS4KmJiMtJGPxMt9uCEsSWoIxMANOU+3U67MreYUpqBv
XEZVOUy3bNtbDg3NtlPILY3BA0IH8IrG39YfdLmahINuKWkYJBf9TEtLfZHfMCgXmS8Ni2HxmEEX
+1aEIapmZG/kSkMdMs4PBCzycsB7UmJy6KzrzCR0pcazl6lJ3P97OqGcgOFYxLk2Ubp7KDiTfPLi
PPFEoC8USiyhZJdMeNCYY7sSm6uyrgxAlqVkdhyZaKaRVe4XyLT5lgTDCpM/xlJgHmGeEe9S8PvZ
eHt8bQmPo/dgzjucKPKcJIFknsf+qB4CyM4nyItKey54fVEsjhtGedS8WQfXIMv8KwTsvqoKc5+w
U48A0AyeaINC2SqlY/PEWaOqsVoV4l9AYvpTvMNP9yvYLSMwl+AI718bH8GiQF0NHImA18rQkJn4
LoEcOw3oKr8BnPLQnQeNCXCpfa8D59NvsPty1w2RFEQk8mXSv1X0PFluiaNXDHYtwqkWCuN8nZ3e
FpfSXXYtUjiFEE4inzXEES6lNLBsdj+2tp5ZVPAFtQQqxHaNm8lddl8YWL4361/H0KawJxSkI6gL
JHZDzFqrNnxzaKmigm4ObAd5xsoj0ISaXCDQs0qwmX6LEybJiiPsQn5s7kbpIDMv/W+2wtdURzSV
c+y2khnlQVbmNLCiuOYNDfdsEPwvhTQ4f6Hs5V+EvXMADFWZMhTOXOTYRrxeGOtTPY5GRHYMSprd
OAhJ/HttXYHQ30s0FWahtrNwN5ZkYmvxDtdx6W+GSGt4CxH6+54cQreKzTRSepFcR3NC6pIhhdS5
zkBzYI2fup0o5TO6q0HnfLobnJ6jKAaxuUtp7/Tvodbc6dZr9+D6d8hzmJjHeQCW+wka55JjE9JZ
oW7UvPw0RZiOuWomZWl/QluAlgDsY8oKTAru0d7biXB+xLgEMumJoeJ0o5Hze5DgibfAtvJEaedR
dRmDO44RyFoi3vVwPjU8PwCHAU7SDH6PMmedoI2fL6YFfH2V31RTWkMGSPe4rORxgBqrA/J2ZBKL
67Qw151xBdtce8pgZaCZOB6CdS9FxATRzO8kBIU2auJCP5pDT078nKCCTGLIv2g8EX6fNbkowoew
DtikY6qtqxTm3xH+1iu6XHkM3rWgnHRLY62IGNuB0osjAUaYu+X3w96bEfQtpAIIlqZiu8VCIAyP
1tTOYm98ArGr5gS6oo8wUhgMkX4nZdhSgz1lpp8X9rQq8LSIXg65S/zXxL6g3hG/IeVQFBXbp1S2
CPrx22F3szRnYxdY9jc9IaEQDEdOV7vaARZiAiM3X3RVNjnckB9IDJLZuW2a+2G/a7dD9QaHt07R
FFtjU4F5hO+uMPs4p8O58jdVs3ma1wpoPubZH2faggftldcdcr16S4qKfCyN3auAXhHjgaaIzAhp
pBeLUroWLqMKeY3GEBVhuFYjtDbc7QY5dy3DBWJlANmRNc4rsgXJvwPeSV/AbWjqVOymzAtJe2oE
I6rsp+uNMAHoWDFbe1Y32ykOzB6GQK8mqEH7KDT9xvip3T1S3XanT39jDjRtIihaJf4xuqempc6d
TKs24km9QoJi+B/mZyraf1UymC8D7itA8dORr/i7LOtrvSOBPQlmLk7N6SPHvgYGQ59zY883VyUz
tIBgRuAFf4EjvG0Ckakfcj3eWWTiht5fTvvOOWe8mF+h27zv+RO1EMOFjSl0SYq1aymi7POTdpF3
A4/8WuMKNGeRKKgxos+iJdqoCv931E1uFmwutVFQFru2Hj4OZo41WhewBd8tNUtGZbCs57ZgCzWc
Q+Uhic+JIjItdTR5wG/OoBSqAU2IyB8u21SHXG7BaHwkML2DRbXIyJbM+DKiryplY1jhR2jTLdyO
dg4uCq9JBfcahbDC5plMFZ+yJju39hCMMJjfj8LP5/SAc0MDCXj5C/ZqyaCJb63jjGY1+2lRBHgP
kzx4SLtdgZanjcx524DQRZEy6oyzV+rXIsAdRzLXFHj0emWWsXDSO7fqxOHoqMzHDruzhHTaMLbp
GARKXQRcf7MpwXI/xBNAsRVTVoBI2ZFk15R7X43JWfaQTkbfj/Oa2vrqHtiqYdNwLQV6FeejFuZk
GOydAEMbUnslpBEwbvIEeOs/lR9j7jmYR9ofspUXEfc6saTTB6evL5w8OL8U8AdfmtNcnqjyiB5g
VrxODt9WxZjot0+hy7peRglPIZ8U9GZsV/nDEvv+m7w77g0ZzgwixkMMcHb7VhtproEGhVfCKwuG
n+Z5UXO/KXp8F/lyEeHUD2+1NOU6AOnjIcPq+CdzWRHm7ebuGWwr/39UFQlcj52OxhJTOyWf0SC6
lhqW2y7Sd/0q3lzRYt4I+fQ7Xt0wbz1NTInE3tLStCajXAmgnivDpIokvCW07sXl2FpfYji7RJBL
ITIpa56b48gOw3s1h36rVszknv7aPH3qgmcHejuuEW5rxru2SIeOzc3P4ZudfR0h0GYhH5b2ZhhK
UzcHN47HcXQ92nPYs5oa+tY6+jTZ0ZPgy1V5tKLvW7fgcI0imwbEo+JfQSg2joOY6CtHYZqo3g0I
HF0y8tunf++OJitBjggVgMOwg68p3QYYjj9LStlkCo4W9r/RQmtRSsssvUc2zXoihpAOgBRFYxEH
tnnXlWSxS4wGK9KentLQFO88wp+IzEOOqblYdmvAJmJMqNQlgKZFTHb5XdON+7a0D47kJRpNlBWn
PDD8uPJy673zgQjmOO13KXFjJrEcSIt3MMOecCUsRppcEGcWJp6MvYXCnjSQLhKS6XCws3WzaPmP
8hRYDDYPPtTKkzxA8KjyZFzo9uAUTTvul/N3VRtajtfKKWZIRliKWl7OyrEaI0mmtuyxZ52QOIrR
CL7sCeufHLWh8rx3N/LfBKK33BH2hzi5cRraWxn2WytQR1SsABYWizgyPyzpFk+fGb79+Shp1XdH
E7s2ayaiWVt7m/fQggpprrWiATYq/vVU/Y/UI2AOfTN0gQ3w8QcygJeie3q3oVYZdQD/6M9IMbLJ
+DG7tni1BnTco9EqAQb05ZA+5BeISV0xvdvnbkVFGPUwOngANxdJqcay8L7/xf/J+lkC2s++7pnF
Q7CKTrLLtVEmj17nJHaqg0abMK0cQ3OJpf6iEW4De+y8hqV+Jr3cdcOH6aSGrzC/rcLa+38Rowka
3sJk8i1c/h9nQlQzGKUudxfIX1bdpPlBw200y/fc57Q4WyTpjngky/mqrESHNthwrgoqH1NTH0eK
a7FpRNtx6nm51U/UbPRXHTuMm6MdM4e3FuUQAYoqygvGaM2e+5HdlIfG2jeve89k8Fzu8ReigN8Y
9VGgFvqhgT57W5jRiBty28SSB3cOdPW2iV/K6vm03iPk2QTBJfze91M6NWTIM2kVHlFH6OJHDKat
5Tr9GkAvHzDF23Q2sg0silpNGIOkn9ji9mQdIuf2xS/SD5qHzO8CPT8IC8RtrCwMyC++t2Yhs4sl
Y6cMyVTUgZjbnO6Gy1GlDSLaVxuz2NS5jMDLhn5Fuo2lMHSIgs0hT7QSv7k/EaiqKwVkdZskzvt2
wEgeoNDWcJJaSivVyfu9I92o1XBmlp5Sm1F0/k0qOfdqI9lbKLljmBtMay1wtDS+Z+KqMR5YWWeS
wUCaiu/gIREp9Mr8a0U6aKdAK7psXrEB2afSWprv5Jjp3NC+Rq3jOvpCV1yGqN3wLI6Dq+PCfguK
4KlHcIxbiRy9ZKfTCPC+v8nDqGP4bUFlrtvKRaxqoDG6SmJdkV/Oe4qLJzbHw0vbuJl8NBSys1IV
UmJ99ooLZBvzSXC/GoYWAdjIm9XEOHHY/jIe4uOJ+O9GdNKm0ZYxSr4H5y7qH1TFWF1oLs0LJA5h
Njw0PhiUFByqgmOvh8yj+nKMFHFdVOQfLoHX6RRHPEc40gUxWkqgl1juAYfzVpUycgmP+FQ3HuIR
q6gVXt1BZATXVQ1kDhdlmj50B2+2FhjopkH4WIcpfJc+YHQemYgh7HeR6v6MQc8LsKEQW2K5Et4h
7/VbtsUxLVgUHzlPYihVRToeP7n+4Yoh/rXggzgEFCFAvygYHu3cF6eFO1S54rOtEbPG6G9pq9k1
H0ywMtwOzOUNo+FDLTeFJpQifLNRU3yJWqWvCiZ6uGxv48ra/Wg4lbJs8YBHBhNVJGFTMUGaCoyx
FzP8Zb0qXZo76xEN6Ao9utBiOzPVNPD/G6YG1VmHes+69OkOTzmJmJJ4tBgyiBJuFR6QA5SvQHGh
jrGH3DLaVYgoAY3vhuXbentlam9orkD6GAUlZMr8Wz9wzjVR0CvuF8+IKaN+spiQvZm5Eq0cLNVl
wpFqTIGw8Wz9NflaSOewJqucuH3EcML62o7lfQjAwHwpgoOX51iB6wCI1VRohkZQt3JR0+IRDjze
PlRFnmrqZXc0m+qJLD1gSUNgLY4wJV+RSR3nZ7PaXtEI7nqYQbmqczKJ8zszBepqarszU9iN3qpb
EEBMonu21pMM2v5Twnh0X+EVwxC/x3V8PuybVVioP25Sna2wL6deCYdgqNgRchOYNReMC7Wh5W0X
SUYGU0kngwbfOiROGP0rblwjndHf/m9yNhRmca7Bx06+6LpNlv0yAY3KXc8BXDuhjCnZd/lhoMOB
sOvTWkZS7V+Oah3PTdHJsTCZ6VpxPDz+1SKVobfMOAUS4Ck/dB0j2dYFIgPfroSjukPx1FGGb8O/
5UJUoF5zbFq+eTO1yGWD96+M9A4DhuaYUSi5ozzGmpMpKfF5sRKT7xZ1wZyfIrtqvh3wykcJo6yk
jrtGhTcdyDMToBx/kJODUgUbCoQ4XkWG8xo1KqIgHWZ+p2YujPoJpHD8zNQiJ1/TjyM0spCUjVs8
nov9ximYSFiPmm6rs1U92lNF0CSq/Kug8+Gqi4ZunPGU0rmsI8Nqcr1dJbifeeASm7loNn3ftBG1
hVUDqUtB1aYO/1d/BQHABTs9FOA4yssEfT4D40Rm8elkWWYzUR/kLj4v9gFI5Rtix9j8sy3vNGL+
qydkPswGfd7mbtUz5P3NrqRnlwF6qQw79y4DcQ048AXF71LAyoOzv7odMbxwDVJiQ+XjebuBdXTx
JBTQh/ApTeBQYKc8JsDYErBAcWpXGUmqaYlApqBKNX9/zIg3qG6r99k6mvjuy30DOcgHLiX/T48W
DyIVyaGrM5qhluyMv9M+GNzja1ATuJKJIvLDqMEdUA+AkVGxNp+OBzDJUYIqjI3pOg0KHZZhSWoW
5XwIuLHMhfQDFQm1y+hJHVCPxXuL/vV+NAfVjVhVZX7Bv2nS48gX2SVxTMLyKQbfn9mvbdqkLzQY
s59v9YBweHAOKHsMifQsDJ1onkUZib/Qr9vM9iCw6h37nAJMxzw/ehTV3H3X7300Ur/q2Hdp09vN
oSYcWWVxv1yJ+SwsuVkkx/aDNRIaBLbsYEVAVXQSEGrKdVCn06eGAqOMx+krEViY4CPjGrYh4VL4
lehdFn0mZKT/TNKiLCuT+bdIxVpj1SsLeRnwvpFtg/cYWYuc/5pMQPG+QWIeXw2UdEZZbS2ETiQe
VBGWrZsObLyEgZBfKri4OmiZv5/PqkZkJ36QOo24W6xTIEHGUzYANGpl5qSi2VVZEObkbKwfH/Hr
nObk2rvcxufdHoFQHWrD61+kqn9uHT8RVzpI3UqFnBVM7WPzd9//FLlBXxoNH5qP6wUNlG11DcIh
i6lKLLDtK0tmmBORH7HJXTjfjno5dBNGQXBuCb00WVlVq8z92P6xk1yfPOroK0x2V7ee8S/EalVX
vdbefk6W8Rze6eIQCsS4JyuGIpKXAIRnrPr+vpdO93rn814GOCJU0N7l+S3WZsp0GO5wGwvYoBGC
3d2d5FCca4fZ8KgLUOfnvnfbQBWlwJjjilWuqMKpF5XNEKCNni8qfBBZ6v9NDM4JZLK8PKgw4L4f
UryW+eIvQZy/9GM8bY3ZisdysZZ8S+mPKL+NyyTXBlLF4MH3VeZkEGhlsrdQMGuRLNu7+gEaxuRd
JDk7avapE2u7pZMu0p2Ns152TRNVIpfVnf9rAG72iNgPtWdBKFeSM0SVPreQ0psjMGmoqX81KD3S
8OX/B3ZkBK6z/MLlQBZN8YeSkvHoN3j80eFrc5MKTYwR6I8AD01zrSzAU4wOY6OI++aCOMSKyAx+
HCtG77U2Iefei0/Um9cqWfL3EBU5x7zjvScK6O2MOYL4Hj9kNRVTisJcO+EcbUCXK+vBWixhzofm
/i6mcdD/txedkHtHGMZy2ITSeCS5xCkdXrOFC+XIQyllrzT9U5QIYt7qM4Etdlz6OqyXobGfEszK
ajnTcKo0wRr0ObA5Fpp1l5PwYw5MFrnK44bCqtLf9aTE1Am2ODEcruMGBsi5z9qrqjwmwRHUkH0H
92bEBEz431Ygv48L2FIzIsGYU2+dZP6nqqQH2lVp7XV1s//Hy1lAaBOMgq1eXVR8FeXKy3TsnTIz
vUJNfxQPdlPVfnroKyvRXdkqpk3Cqxh54SyHCtwWdJ/LLW3MAVhaBEvEJn8rdO0co0CeXu49o8Xl
Iw0OhDB+kUuDsQ6QG+dNpCnRewR2/u6ZFeYwVO1ajV+rbOIDsnRJSRLehlC3EjcEfMd3+pVtekGz
vKTl/VOeaG5SG4NMg4vKG5E6OmnBSoBXhTPaDdNTyj77HPOMhb/gyGlZv+Er836ie3rl7GWWW5hI
tcYs6VFprqhUPPwGwk/tblXCfuar6/RzldrmGit7IT0aAw9Z8nwhWNFB1qbnvadEiqCji9ln0Z4L
cCy70GNc7LrDgbwXSZXwCfKs5F7Sa2FEYOP7StjhV9VT+mSciVshq3MYSAUhEc7lr9/iu7He5Njb
aa/X/c+Fi4/y5mUEtMZOuIVw09I4+0V4DHMo2E554mBRVikupT7Ctw8dYXg1L2Ol25EXydCkJAhR
HbNh51nIqLqkrIrkBtPaQHt0144EjcbIUBuPxVRpgqiJB1QQRAWlfilG60eKlSjFe8ghwydZHjm1
732wQxpMnSl8dO9bcacWoTWuRT24sNauKa9YIqXZ2iTgrr/EoFMzKI2tW2fI2YRTKRpwfvC5h8dw
w2NP4/35/elesl9N1LNe5RqZjuiphdsDPMq61Q3H8X1L+8Q6fXFBtinJHlJoBoXh4CMLTU6Sjb3+
sI/ryEtWlM6P+bLFRsqItDpxRAuVS3uYO/FdsLyLx5hpVS3v5e9HpwAFrnavad6GU69SKESNawi4
393iBsisORxdnD5gOxidiQoUr1GfW8ippG0rbx5nLl8+I1KExqtDa/mEPp3P2JTaGC0S2QbWv9h+
qAU3zkpDiPixtaDuf98qQ+Aqra9g80YVeNLjjDTG2xaqzfvTqudzELVhJkKthBEe6NDEKJdQ7nIj
U6awVDAYLYDRr8rTOhXSjIXDwTSnwdgAeXeq/exHHJksksMJRj985fPb5aWmhRvDR8yGSFirXszI
tkC1qn0hbxzjXSSB2b8JJvZXTGH1PgiKrj7utd3UnhZRIQxM7pb3XMfjZYwFr3NN2mp4mqRnZvLO
R8wqzdjlLaSyoRQUe//l+3c+kg03sJBP7bVEr7dVfY05TXWotyoQn/0YQyXxEXhwFq3ne+dyh/vC
xUc3IdQOWcOjpyuLONshtK85eRE8QymjP7vojSYk0OAlE9wvBp04twAHwSPQiKKyosuo/aCkY5Wr
TMKAREkyXI0rRpcDEUay2U7hv0uJyFyd+rDHKSEMpxpC5KvDwKYzAwlXI0XUXuBUcHzDsr9c6O4M
P4ZbAqRqjnrXmxA2fJv9TyAY7rcC8F8Xq1pV/oItTT9qsq4IncFAGjxlr2ZuHbIUEsX8Go9bT6gY
9bqo44argSbkKoBS18ZnxvlRVhDd+1wTxtJL7hyo25exsFPf6BxXolxtQeQ3vbvMqpAlnXh5Zw9Z
1c7bBDdwgCLkrhZdhmZr0oj/dhhUURRTJmxDnhdO2G/mmfF//VAodTFjCcDPiHI1oG2LbWx5n5y/
WjnyxxVD1Rlkki53PIobJdZv71bo7nyJgdqc/vgvYb26grTMx2rwZSKzw+DVsKg4ygf1io/KUWoZ
V2uyvWN8qa2BKa4H7JR+0Y8EAfZtY00Nzn+isZ/8XBFVJf7xzSSlbL13c95zjuQt5OwJXgfJF+3b
J7RsfFOCP4Hfg1XjfLJZ5m16KLclDzb3CngkK573Gwhrj2OSwN4ss+yqX1F5wvk3aQjSemvoqu8Q
CX6lzA95yUOZEQe1oFRaY+oqweT7O/enOGpt1t+EbMQyI/4cMm+2v/nLdDRIN4OkFc1FdfoDRTzv
O9piR6Rutjjy8IUAz89RdooC0jmvT3Ov/ei1HECPnkBj5U5ZU4Y59cFOWI3+uCl9KVz/HHfDsyl8
gyLq9tNYq4PHj4yrfdj/n9G8hLB2id0UkKfDbckZbhKsoayLBE57uIfXfJI8G1m7aq4VnBdIeWXQ
Y26WudM7ORs5D4D5jHlVnCFuxQk7yJWykOO+6XzKUbGU/i9hF6aF6Tgt8MUStkqDHL+tEw7TVftc
toQV6uTXum3SMlZvrz4xnnsnqPQHMKqrI1QvDiOakOVLaFL4WzyOV5+CZ/G0noscE2D+zXTv4Ib1
dS0D+x0qM7OK5ArQ16N7j0WV+UegimA18CJdRXl9M88fo7izZGgYlFsXuK9xgLgtnDHPfQ47peoz
quSdpykAbZDhfulSujDVMuLMzGhUcai03xRmJt+Uelxgu9Y63D3KG6+FwkGQ7+ZPoi+S0m40MVaw
IJBhVUAW32w1n2o3xDqP1tY4sx/jYWjH6OK/VswaEZNRlZws5DeU5zr6RIKfzxgJ4iMRghOjT1qr
9NixrI4e8tucoPvfJQNsWXJgivuD5F7NdQBdXZIZExhVTbdOFd2B9xKDATA63J31+gCPQpsuItuY
hD+Cw4bC3nOvNYDOdd3x/2l3mMkmiM9FkocRIVeim5mqGFvQvrJL7ZzXvktc1bzPjufwPCX4orx/
PLAmt1YQWKcFAYqtJu4dozrVGQ0tR1NtEUIDRFDPpmdmbp3w9hhY5SccfS1lZrHS12Cgp6D+skRE
2KkMAmGb2y6/OzO7tltB6g6FpBota6BMHrvlV6SEJoHow+LCV4oNXsy4BIasHhGaMlijTj0BFeEt
qfhl37oYlcnojCjg6RQoUXSu1R3gJ/7S9DN1ek8iJ+7fuy32fqa3V16xNDV7Ja7xa6DPwhAnrKAb
vPBfb6YyZnirV2ScrN2Gj+W3hCC5sRoNYkKKa8Q7Xi5p3rwRbeB+SMT+vVlBjiIFlrJy4HJ1BR/F
PSdG0qFmc+8wq/okmM74Uing2G/F24zjuVbTEIhgqG/l8rTpRGWamvzWZqV05yyZD37wuSOxt3ba
KmC2nNoe8PUtK43KcEU2R1FtOzkCgCDfR3Z9f2MvfK8R5pIjIO254BxNom53vJLkfBXknbT6NFjm
IxwC1CvTF2vGPnn2LB3D/DSaOwXGE1JmwYwpH5McznjRdN27mDfxIaTuQsSdcF4wHUBlRUjLQ2TD
noBh/m9Mu7gzGPjGhr3hb2DhF1l0Z82CoRbzQSguniGnSD+g1go1ikmeE4+/VaW7i9WDAJDQCQnr
Z8hnXBuenXPdIywAItKv6HaqJDLXrDXcLYMpY8VVmCGVoFO/EvDERqfah2Rkyr5xKzptlsraNnDV
GTd5obXhbwzb4Q4H/lKeG9TTNbw/tOzQZ+9x7vmhRAoTuKWfNiU/8xfCHLAHDeh0upbTHQ5yU6yd
5sEA+fjT+bWu42HunFKYKoSJ5gS5fO31f5WJi+GQdSHoAqFVozf8u87sYnyBslHsENx10UEmmQUJ
mfWRs9+NCC1+o2zTvg5ZdD7aDqoc9WKQY9GRbidQofDIieYx4BzpBcINGkdobIFESjEr7AFDV8W/
EtVwfXfCiujfBnKLFzeJ0owmn8E23nZGGm5h+ldwwk2fnuLOswY1HM3kIhzLjwGgtSb9+VSrHIMF
zLKVel+6xxY7qKSbnrWxGQCBUpBCP0gQkNyb6ybu3a4N5vvFvbjgUr8bMNiqQ/ZHP/TxRXAdo9Pt
rpaq5JLezxi2PvAEE6NlxfioSALqO0cFBuoAaXzwIfG3OjMOBEpGmdXjBur/k3jNXyIJAXHUkwhw
zPAwWmI6QBfXMZYRS+x+yTCi1DKQDvKqXeEpmPiGz7Jx5iOx/fiLWvLkeHnuTIvqlXFUV3OoixjV
c1KsHiiIu0MbwB0CpOMd9nI98Icl5yzny+BWrMYaf3llmMY0FlIU6obwo7VTaRd6+rGjxFb+kJRr
tmN2vNThEUz+1m+TGuYKmLi7+dwcvUqbpbo9QApG6qGsOSrnbtjFwDrJliKwVkTIwHT8p8qN8Z2y
lg5KxxNE8fgxEL50SR00HIIA3kBqFaP/SOWcq+r7Mpme0Lt2LG/5Vb1JFKo5mbi58MJSpDgGtZZN
+rcrQiLGavrtHWw7TUNfkeJw8tmkKMRXYWrCaVZz9K41giyYjENsYl4h3BTsPm1Z+qrDntKOvPrP
eUfe1TzykI9K2y7hL+n59tve4zPnpPIWQMJqtdVOKBTysv5XFZVW6q2v/LO54K7cepysrweLfS9w
ZP0JvJgPYP6LjDHTKxL8t6pCZ1sL13rYpgUOkRy9ZHh084XsM5RPa99QfIEOgCW3ZTJSktSa4zfg
xPO0t0YL9v7Xxnb/EimbSXU2qb6w+rNuGNTEU7KYdNFIqgXZ7jpsip/4FeZ5Jq2IYEE6LNr6GI1C
gjenkSiqI5vWFqO1SHjfwhFTpLZM0OefTNzXtZQDgbGQQeavcMt36gdSUnlMNNeB+wmKDUqR2a2t
VKqHb1rRY04vEESVFsSZxT8mKANO2g2s69hN1RVzk1WkMSi90V2U/tbpGPC7u6DGQDT0wl0483wB
DuoyUU94mAnfil4sUEK0++FukpUTAR5v5PvGf3Ei13Mormi6KmjWTxjpy93oHauexG2FaH5v2XQI
R0LmATP+m5sPnIyxxBPEneMv9QcktOoxr8bV7aQvpOIrJxH6C8qOgbjAuWy7WM+41uCTszuPQyhI
EXpXjRtBMFUkASJasT1tiwyX5jcUhVzmUpx6vbUpFgQSqKWbcT44VHaWGBfwT5Rg+T4OLuExrtrx
KYLrR7A8FmhHKiCKwnZ1zzSfXLpUfbHcyd3b0zAthLMtZ08bP3Oawp9K0cXCLJ+q7FTBdGMnGChG
s4RVXtgkFd9LAy9+MT7geKuFWTq5v9Mt4kn8WIQcaakAJoDjsx+GDG0E2V/VwhUlvsKrSmOGB0M1
7H0y8bizdv6I/CXtpPSNxAYdZ3zJeyahoC2hgZkhVEDSczG+UoMn1qVOz2VTpr6ngHvwVv+VdK4L
eJruiHR99JreFjjR+dxLFoIqFRZjGwrbaJgjGDGUdICGjjZSGDQAsD2YilTivxOFY7jm02snHWk/
Ez6PZ5l8/6+2F88Rs4AJ7+N3167ybwATrzqjkoEEvwE8RLR6OTAO93wROEnzd8VEJZUIdROBvhP4
3gCXMaeoklnQXBu7r03pbBBJNon7jc14V8uzMH14ZDOU33I2O8dV/ky4KcIyOsCT+IQkol2ZkyzB
BLY0cjAElTUMA9fYyjTQ208e3VwmkKt+Z5tj8iwa2HuEscz8ynzpfaUZMwLsEHkPeGjPA7hOXwwf
D+KxJ/wfw9SJ3pTuQXShclp0zQ7uMc+gC5w/jvhIyhFQH7xhMcfpLep+cEFiKaCZYZN/dni+0Nrw
Z616mMBJJ/dy/QsRMt2WxZPPPSwrQvlKO8jIONUb5zfxTv5blA0PdguT58jwG0egR7iHamPdrxDI
0JvJ2Yt7bhUQrBB8k0PTMwbL6DZHvEKkYhB5Wjo9/27U2XmQ5C8V/cHupIyQKCSa/cr0ftcUReaQ
c7XFHxiicDTJG8/j2JiQj9u79BexqseuTEZniIN+W79iG/RAElv7jXob04gaPtFtfKuA8sVFOPSc
Od+TWZwxVOH3oRj2RMg9qzxGOlie0rllZ07kxLtU9GiDDb3T7JDcGs1hsSknxv3z0FLhEBPAIKNe
5Y78agn/lJQxnAV31RimYbQEh/IA7+EELmhVaGBi9uRbpMBNQOOkTNzVzcBRAfX8bMdL5R4Nfym2
PmE3tLJb4ks6dFsXCGbouGQuBmNSDHr4r/WTM1Fpt3ylK6IQKROjgyyz8E5LKgqVEdMVbSArm94w
Y2mvJH3ElLYg3ykZWbzjxNqcv9S7eTVk/1001jRGjdYVpP4OrqDmg9V4ds4YQYGUzaFBsbSBaeqY
ScfeydWmJBjk3WAwRFokWWfSWOjr+6FVgOTfXtlyy2+J+BmNTG9qjmCDV/L87OXoGagZoanuJhMG
FeDtOF1rqY2gpP1YeqysDvqVNZ1GGH/IaV7uNKI6LFsU1ti/ASWXxCwEkY+FSKC/vxWBjcXz9LIw
WS4E66kbiW40WDw6+yNuSpv2+v759B0GDwjVgVLHkk2uvgMbwoPI7Cp9juuR+eUI7An/Kge/f7lW
hkA1kkH3+vfzNNv/uiDtc8scmCKeVIGTIX4+DMKmysZXrcpWobSD3Ip2SBuxGOFWszIzI1woLmOm
1lK0W2cbWGGYvu0P5AjGIiKDn7jyKK1+KOUDOO29j9e6IVFhv2yP+/pivvcL9aRzKdGxl5Nxts1h
BZsAuyyle47ybd7/9kmAlfnByJq5HI6pQvxNEk8Rspo0BJ7qJ1Jn4/x3yy8Lwib0i0ZvzR2A4Agq
BYX9/0iHJq2C2LqdI1DRn6fgw2I2BBNw2Sjf8NijPkQ7/hEemffevyyAmvSUKZLLIuznRGKBuMxZ
UE7VUpwyeoyJA6rz96+iNU4ivtvBYpjQKmsslji/6H8iJA++qo8GZbcay5OamRyepM5wdJs69jrc
G5UDXYa4oJguI/+jHt3LfBCVet3q4iEK89Xcob8OhpELuLh/E0BzMvM+uESfFao9eDdRlPuF9chn
JxOF5ZPpGxd/j6tGlIu9MbdU0hK7oN+TD3J/awlGav4KuIqR9ubhr3nQYIosbcRpO8uXC4IDGk/4
97CY17815+3s8GG72JftLs6KfvsEdVNXAVkyTEcfSdREElhTE3HaN3EOWcP2N54ryJmmvGypiQ0K
yXX/joFZ9f7TucMqoGdmXx9n2qkYpQ6HFmk643i5SLAcp/dvj4YBQ+0yXQNdYKWBq3mKrCy/rJ0+
K+k4ssC7Di/+mcLLWBky6Mgzwer4ziN3uPFyWtBXc9HepcQrIEzEHyU2P/mb/5VpoNWlDln57yAQ
1dqfvNhJfOeK0D4dGMJ6pbNO9uZNZL+RxRuWU1luqGFr+D10daFPZ0Cqk5E2UpVhEXLUHDX6+5gI
p9whr/Hjab/YEgByNR7vsBJYzyiI2l9p2jhVYX4YkQQAU/WIS2gJBtFFxjqMZCylghK7kSCeKodf
mhrCxe1XBmKeZ1osIQlxgwbtdbplS2jC00BpqETPCTmMnp+mfIIiz3HZJzyYB4z+4iU6EuJboz9U
YeVZkDIUC1GC6qLavi5bTCTi4873hLzljItRAwaisjPW/XBMuMXxjvcoh6GVoP1OA0VJM8FPEuOK
FFAoFcQxii7Ujayklw/MXz7fBao88BaJdBz2nLuPk5zn3ajyNmrS4H8lYLX+iKhvnxrnM0zsTQAg
hLSoq+PQ9Ldm2yVvYzZgVgFcgP/3DD6ssTFrcFuommE6girQW2VwtepJsu021EB4iak4dADgi6+M
ZMMJ/caqq5otV9mTRhZVrqpU3O8KNOaGYqsC36D7dXWzluQAGJGwnKFA4EAOfMs3DA8ML1CXC/aD
nWaV0GEPQWrCIuaRLk5oHhi2+5/u280LIV2+YOa5wU6srT+2JUPGGUz5ArxZIpGHDJtYYFxvJcX1
+zPSmyUWS3IXguMkRB2BXZEAPlxEI5tUXAdgAgH8B+6UQVumLW7EqDVvlaZ3J/0hbv5SWbqTX5LK
dB66dyQ2yPQ8K6uBEObEAwMGrDrx84boSuIE3OSmaTWF9kUFsn6q4NxNvGax7C8rDKw52t13vsbg
QPlWgZWXWJCnWIySjRaJztgxLxVl5saaWy46YHJriYOFIDepdJ7NtX1ZGcvr1mrJzMEJ7fsyC0Fq
47Wx1Qp/aM8QjIWhr5b/viJ2M7yAv9YOeT62TM+8AAbjnDcBmD9OV1R6JKaRlMZkROo1CGGmBNb/
fnzs+AB4n5tNdyRAcwM49bFF9a4XPQ2MH6DZbEqifdoituvn100qLBbXlBo6cscsnvVnUHTn4gXz
Lq6ltLMzEamsSE1fncNlkoSDHdb4ZTKuoRjqM0FAa3hlRo5ito2rslQSBFbSP9iVscCMJGe2Y+CG
kKjSDSBByF59zefYGntLjvJh7uXLZP4Gw2LSOQXVTHZ8O0qm0Nx/XhH92o6MupV+Ze4T5Jo+uR4Y
1op/kC9/tXCptttzpbYL7E/iOH9jKBBlU8LdaGxqs4jA1iFoT8f+IYLdoS98TUD+3s949Z3nDl+g
lZD7+FXNA4lsk1qC7KFbhw7Lrjy8p4t19geiC+/vgT7MWKIYGwSWjnjKJ0rdldHNCFlc9wtMSysV
ZvPLIFTJdyTEV0OXKyYftCQKtLWm7PBxG8jRRFIgMH1tHVKLjI/K3brb8JKKR6aezJm5ncOrtAMz
Pb9lCCuiVdosaPjawnSgkrsCSBKyWx9Wy0MwC9sikgNa6zKd9+eWYlKze+AJRIbrWA+Xaf/pg/65
LYb2OPzwBD4jba+Pk7z6AJdPqtaxUicAsH6LGQMTtYVlBduOV+TbyHzZoLLWSZAAbZGJfXEXAVHp
xsUPi0eQquE4CVaV2W/rEu1z8cjSY4teFof9wjnIWlRYrMbvl5CtjSH2THIyVi02NZFh67PoqdSn
hUm6qb2PZ7JdCi5/a+WlVtWGeX1TQyfBPYWawHRk0vc5Qdoa2xa91j8UAbLm+YtzCzrSc4G2+yg/
/Q9APKfJ0cC2wHMWg0e7HxynWf958kHw0o+Gh5ee8jRyDuMoriDNGrzvYB96WCGxMlmJ8yPG8yDn
gqRKwiJtAdbvzp6CfQYKc0x+AzBCmJ6W826VePQzEoz7Urk4opi+/ftiftm/ei4YlhXJKvxEINlB
aDHl8tW18Oc40v+E0IVGl705PhZeb0H/At6rjVi2JBEIfQUOGcORHnQCbJcTgr1ECgCYJyaM8Umq
FQ/IBdCznou6N63V5du9UzPVFNXibtbdHaFd+KICx1Obl/AS7qjyk7W0aYaQIBDxkpPB6Yb08mW1
KHpU1NWVaJDQnfnexoTBjUgKOHRYW1TPKTbzVvBNfBEC+PnWZPUcvqiSNmizpqW5+dg6tLb8HaxA
ojRVgVrjS6lSu1X5/h+0pkgNmFcO0wHwUpNvXTJ9UDqPSbtLOb9Vhi0zScOrYPG2+K/h2zDXRXTy
EpryEmamqxkIenvR9Rb/oHpxBixLEMQFBYYB34Mx8+W+oLgGtk1gg+AnoJNANfuLhAyWJMU1rZzB
CnK9mq0L1zoZciEyRXtEaaGyhS+A5lq2y61YkG9LOr5zKc4xB9sS8wB41dk2p6hqlJ8YoJa0Jr2K
sHg8OSn7bpbbEp7u83GXylVHVnPxldiJC/d7tvYbDhibDh1q9bhvXnBH3sGohsdOamIEg4uzqFnP
RS6Gx+3R7ObaRIha8Y0U2aa4JXxsL9Q9APqSM7LJkR7zkOvPVcCYC9WGLLr0o2tto4+HRNg9wXKo
pb2L8+DPE2FmvX89FzED1nGTgOfi0To0BVHEJ3AwDNoU+zKT7XyBjviV/Z2WO7PKK/sCYBwXQdzN
tqgoP9IJqsemw8n0ryw3vBjr9gAsv0viDcEZAu5saBa/JTwkC6USRK7Nbijgmn2lzUO1wvIJ3a8P
J0y4r70b6AhNZw1d9LrTrd4niPywONoSoeiae+9RaM8T2ta+xKHRKZw6y7pOVqncq4WCmYSDCjYY
36fzZNCMI8NsqFS2VF4XHfj2K3pp0VzTm8MjATnkJFfQWwV4sBKNYSNs0xOoRGW9znkYE4c3aDvS
WmdKMImfimkHYUvr4ig8I0ar7Jh7wVmCHXOVRniWL47qdUi55Ayn5tCeRgjvxCW1ON3xRLvAC/I3
8ij+uz/K0aQFM9hbylLWO3rOpol7/yu1PpG9VRWsFfZtZXvJVN7ffkeLRSFEAWK8FvwWVXYIefGJ
l03wyO9yHwEBURpSPqKmpWbxTbwaJpEHcnYzegilG18OGg46sFkdA+xGwBe+RJIaEyqiS3I3uoxt
EAARHHogl9Xy4TnJWd6cVVducKXcp27rLeE9j+GLy+eybe+3l53MG4ysZ7h4itZZ+JLldCpjZwuO
FbX/Lczq2XfZU1utzi87lt8tjHSqUNM0CUAzjUWUIEC+aVHNeXHdNI3pvUF0+mcYWpRRUyvh1Jbe
6y+o0ZOdGxuhsqIQ4SW6/FdUixaE4bbOzppQWOb06gVYd43O+Uzrfg1DysCklgqiVL8KTWRmp3Tb
ya0XuPLwmy7G8dhuzZqEaJMwt6SwM17KmpeU9Wa5iZj5AkyGXeuUZ71JdviJsCvl8Ad9UHnUTRzw
KB2p0SMUVePMJcXGo9vwUvlzUEJY0RMt1DGXE+3H6MlBkUYjyDiwhDTEhX0Hiz/JSxB0e24VqarI
Fz+njMzl4nbQfUrx9hp57iVddnjvLTBWIBtDrrImo6m6EbgmoZzD2rqWT4vIKvg050b82udZW4PK
l2ttx56+rKUiZZ43KX4tvTaGZh9ezKNa1r27j0Q/bhkBPGNLOakiY63TvPNmlOwrTM9BSNGXghJJ
vYk97XMFYe4HbNLdujt8HmJhiPUFI3ocJ4Qdd7F/+Ug7rOCjBoOSXUGtGEodEft/npKglXBGyw7w
uEWTfDNkegg9D7mUtNehzMiHgDvvO3IaJkRKA+JQ36xGseO4ACz7udzl0CVyZsWd7lHPIVJ6bESj
Q0EgS5apdWgiNJh2rlD7VIsmN9aTnmAhzG5NQw1ilNLGwLHgQhrjMVdQSJtK5Ubd0GOjqGswLFt+
Yys2/dFB3OVPZ144RW7UeUIjSLvT+X1A9S/xi7Z4penLzRZmRMaKwsYb8YMhDYKnq30Hq0JWOOsh
vG6QIeLI6cIuoYVV4yrxS2l7bRiuP5KzgLHIudSjiyEVZojBDXcWjCkwosLDponZLXA2PczaH+qK
daUit9p/4LlVJtixGbilq8xLr7+hhqkWYpcUts+l+H0V25h/03jZnOHGPPJb3NKO7zO1qA44Blmx
6euRDtmK8s1SFlAbJJRVhq5kdrlQgseJatholMjhdYO3R0MWzgJM4XBS4Gg6ayX+cCcuUbOvENjp
RVpmBul2aKz8E2NMPx5U8T7EU82qca2jGH6XUFH/5YfigsU6c6CUQFCp+GhZ7JAeRe2UdLl6PGSg
MfhB3HuQOvNPEWwi6UN/VDbEfBGJLyCi9SaCTRKptn6XjjaTE5z41eD6XZ+cy33HHWTxr5m/NbS6
P5T2MFf0xTnLHBxPDHcEjuxDvV/90iFWQPHrcUHt//3MyKbQhtB2upFlW/jnHmnWQ4daOH8CNRUz
bDVK/tCr5FaquyJ8rbpJENHeSnnzkxHgFBPHLpfytftToYJfrmSVYm99WRdZM3UKoV6MzMS1iGXb
M9C9YAlyAs1l5cjI8NvNdY3hsfk8gDeWMk5wEQ+0pbHvd0Vxsx1kzxv8s+5grVjzR22VruCbEpHU
L/G25Fjl68F2ppuQiTUgulipxpn7kvXpxG3FWxdKKpdtRfTB6N12j+fGmOjdt+1ksRK8gPE5ZJVv
Cl1eRN3MoYTC8mqBSt0cf4CYWGJ43d5sEdqsjvhOfU68ZzSBvdXKzDSZRwp4KDMv82yZ+GcrlbsS
ZS7tUZEiknbraFQU6UfuNTAJ3kup1qcjldf3D+Tsn7v/MIo7FJm3hAKAbT9id/RP+zNg2W0X3uMR
UIZvOvIy29fdAh+yHyQF/THVquwraBBZoVR2HQDNVGx6E0aWmXayEdPdvz2ebXEOR/OwZ0WKFXVP
qQhKbPGgW++EtKyIaXPrJ0jH7GICsfqtCf8CXFv+4FG5rC0qBXs2YXGIIfqNE3Kax3opKu7jczlJ
nlomH9W8OPZ55XkEDLRWki3UVZ3HrHngIQD8LVvXII5eEabWwGH9TrcE+tWYIg8NzQSQWQrsKjD0
camN593ZvZwARO/CLkG5aQKjRFKqEkR9ktzqAZtH1xwv8Y0WXbSoekX24p2Uts++3AYmbeg2J+GW
uYmIY7g00bqIO9tMDxBayun3Xija4jkHgZpXT9RLD1K7kMs+zYdguwbuilVMhAwp1npfvUec5LpM
3gjmJ2wZhI9h7gF1ZMctmUoddQbyN42Ij3rTFtnyOSq4uT40SHSYKhjufSU0fGE12+sfSwuKlPLj
xMJai8etYdbDUQ/NSqBF7kq6yORZttKCjIEf7FpAPa2rY1IvZXjb+A0oeclGnCGkiM0x60NhTfpO
Sxx/cEKX7GuZrkrqoLvfxoJ2v3VVjZbHPr61xDA8jbqpQxiIGSU71RQvI3bbzuojlUpMfUax5qk4
VnLzRWv8XClgGxcRfDzwhG9AGF8PsFGkWgvTqhqg7P/Vuy3vUbKSn+SRq5JBDeeI1moH9ZFvameF
HoJ6N99JVBMWEUTnNkOHERHbCWdvmu2Wvx7Xn6/pWmXESEl6vLmNRlIp4jro8UVTyyVoi+NBssWb
AXSXo8y5U7Z89TXEU23TjuuOMjyPQWxKfXIhsFSRMkw/Q51iWlAJQTQQnVG/FfG8lqYe54GZCHWF
aAmlACuyJ/ZrLPWh11uncs4666isQxCIZ2ldFLs9pyupyGEeq6wC6v7VZk6fiCNlLV2S0WfbShuv
qzc2OoEDw3W7vQq5X0gBAHuROabbER0y6u72nEL/NdZSJnc/UbDuPQ6A8gAje0pVR2fE+biyXuTl
8XwwZiaBMuh9eOePPGJiL9wOsxasrIFikm2LKcEO/02TMIUK4yJhMTpwAoI2dqXph4ON4Pfd9t6v
HJ7NjvUWR3UPTm2QmsRyQdfLCMnDuzUSA63PuvRbVMKpgd6JhNcIC1iacKz6PBvvEf8q4igZnFYp
OnGXpCthIKmDu32o774Sd0E52W+yAgKGXxb4WrBLqPUQDnxScpQXEEzWGjC+n7l7xBA2QPERo3hJ
ZGEvn07aZIz/mZQm8d9J1PfnQf46YEwduuDc/CYe7T8MzM2jJshu3gyuhyBq85qAmF5Fu6eF5UiT
wD9w+hIHCnfzQhcY1EJ3/NyRWvMmt4LpRIXp920XoVLJkd39jLJxHbuKVAUexTW0CqdGR7+c+X9D
xsvU6zQ4/xl8nD8quu3PU6VN7BlBAjSJlcQ7taHtYHm88KCzmxMGMBfBlg/tJwk5tt2nlaCGm82/
UWMAxM0UfRcsiZcQ8ogo37b2vRI2mLycZVJVIZgpQfFOEvpFZ0lN/kfuBp008iyM360ERO3LScjV
U3LoGzSnbwvYla6b+/XgQ9Otukc1Fe3ybbOuFG49HqbZYMZsOj62KUe3IuPgQPH8B2Qtg1KwlK87
wvaeShNnWX8IPaapVN0fMAfnIESD0W7DqniCCAODkcz8VZgE0pc/GtaSAFf9YYEuwwzpSb9O7Qpo
kABhX/smlc4jx+Gy4rRybXJymfyn1T1nNlSMntb852BNZn35pi3gZ9myXuNsIfDMpKJRcEmL0qIj
1Zs5GjSjSgIeGZm9spttB1tIg5su/iYXKF14fLc2F3V9wdoo/qB1r8Khz8VZlAIuAX8WPAt6mYg9
FXOS7mDjnSmE1nUk3nSw2kbDJQV5a++Zstr6jh/7z4PQE6I+17G/W5BKzJUbyyTYQZI6N60k/r8l
QviOh+SxIalcQmK5bs/Yg65Lzd9qreZ9HoT7NX37635eAQ/ha+No5GcY5J91A9woXOe7Cl5wPbDA
2+GzTdzpeG4rv9bKNYvE3z60+QVkqly0PcOlAlFEHJSpdIXUB0u72vRYO3mVMFmUz1knHg4DPtM6
ws8qrvtHXQUfSiBoUDuNdurio5DYZx+LJOZphKtvhngpKH0BUyzCFlCObPmzt807RPbVxJ7y8uC2
K5+mD9tZhPm8y+iEeMtA7YxFoH0tNU3EYkzXtLUZruldcJ1ajVbJ8b5GSR/RFniNyvxJ7GxgTqEr
RjCbR4NC1WVmPGWR32rP0uAgWel160CuyctkTfEWxkhw+K6Ygo4BOQIPtYE/x7vqg6foiS8dFrbc
E938b9rzHQR9sVpHgNhxghco4w5tXzTdAmUEINxUFCNFqAd80/i64PNxa2BOdy+IBHMnSaBDsasx
ftPynqB2o8AgIvU+phOjb2uHguh0IjetMtAxED+8r7se//yKoV1o4MsnroJfI+IVrQBTfsFzoqMA
QRadNzjaf8xEuXb7F82NM+K8158OGmGvr0+khNu6hmRM+LGF7pXF0vUX/MoBTLct3ZJl12gvwqnB
qRBZBBgqz/+YGyUz010MpeClIicDu4UhntFrYbzwNHSP5hfuxPOEsiq9g5jkDxpHde3YoAb6600H
AAnJrriLwKt7KYPs1FIgBXWu0k/GByX7aoRvvsKYxurRh1EDAI5QX9PNZmUvIbVwOVnjVRl+wv+G
fKxBC/tY0i8yiQR1LDOwpQIK65y2l6PVLhMtVnM9TUuIgOMczALki/3r4t4isVcGk4g/ZJ+WERcU
9rQuwclNYN9ePMB0H+929QxgSzzpiJ2Hc6ggqEIEEWuy6TYT595QS+g1eC5ZFyfS+ua65lZFAQWf
T10aV4dORhTLjsnM24HsDhDR+2vaRIVukAiCzgaB92Bh//dYMlSE8nh30RR08uLRG8W4COmXTDc4
q4onnf2J16XkTjsSlXb6ZzKn8HqYjlw+jyQGw0ut4AyyZ2KIyybp6NSldQBCV54ArEPge89XqCAv
+/USxWPWFDKnBqKtK5AtND7J4AyVqjvVNDybhPaeg6Hwp+7opgtKnOoO6OgVUAghWRSWkN6/2r7t
xhALvggURCNU+JqlNXYbMYn2whEx/3Uoql9P2Ng90BpbzYue19tSeGIgow+ScRdzxh00ei33W9R5
EZTCul0zJgKPnnUcwieOCbI3gqSn1kXRGzyFqXhZ/L39NYj4Y72ryy1SroAxsMKcNlWNq4ATxxYr
+wGl08Y7/5+xvZD0T5pIKqXIDjLSruAa40h03cceim8bW0eElOegiRn7vZ9ne5p9B5W3SMKudbi7
97z3rce5dMu2AL8YUKdBhgxYOjSLLiPoDmUBJSDxih1p0f5Hf5XTyCha9lx2wM3TQSx/EHGB3fjr
IdwHbfaz3K1KnnCwajlWUtw7Uwvj+arNUqG2qbjguGCTMWpk8DgpACJssEAPb0jw3Y384e976w3X
RHqW/tSyVBnsR57S3eFnfPOncrfH428IhQtDDACK2vdr1ZmhdnQu50jR0lNL6nM3lxweBNWToFnE
3MOy2J1l04NYi8uOGOxM7q7mhRnUwC7mpEJ6eabbvaooXFtCc6Hyp7Ldzstogqj1dQb3wm5LaUjm
PQ/1hTaABTYc3CQCeTwY0RQXnkss8dRFJA3O6k3tQZ9CICR8XavbGJjVX/edhPojhU0rmq72pYpg
iRoW8ULEN+LdmhhAOS1rDyqZ1r2vX551S+oovovdzCurI4Vu7GcRu4rXQOk+y9FRS3kDlyzmJXIO
+i9THZvAvVLxbaYX7oDMohVMtTNdPeN6s6s1IqJ4JzSp97IIz0qAROFr010fWJiZe6P7TaLdr1bb
mQ7Dg/SRhGssRhTEeuUNs/c0qR8+w9Kh8QEpp1ag9g8ifAOozs9ZU+wDY9ofx88WRQQ/75C1ypq1
uVjBNlVU9e43nb565Dp5RPAIU8SWc6M8IV7XZDVwE7Zx5z66GtLuGOD7LYKkfkC1XikHYfOQDZnx
Z5jZSv2j+s6NCkRUfnRIPKxTWMayLtr9iC5MKxrlpZ4pEjjKPXpFRw0l7IIWyhPHiNAl4Rv1Bb9P
CsmCwjk6ACpZjxqMxWjzqxVy/5AGCc52oHELp/Rq3opKNp9naZo8z1yc/xBxNz7K8VP2ovRuYvCj
3TFp+4H349ZxDF4KPSwm2VtQEWbl7cbJJvIL86w9hXQE1shSPDox38BjKJFQF1M2G7kLa96Lf28j
el+qjwJsUhZYoDOL0tZnQ5DQLEiUmRi8SIIYXzsg9LRyOAnGzVFvfDpHxhiN7jtTVk3hsuh0D8OH
Sq8uLaDyT6PsWrSvgNX72qUSIBW3HGm5rLAVT3i2KNVNI/sGLorw6Zcd7atCLG6rcOAf/4oPbsic
kyNdoxJPUq6X3zA+59Ry8vt4m9KYmxzijBcZAB5CLpjJ5rQwbKc9Oe8KteJ1ftorg5cxEdTHQnlr
w8atIpOJbdSBRJarrUaNmfC2K9tTGO92kMkQGHfLE4/liu+HS5ysZ/DdqSXJq/isQm9GB/7y1QLW
bsgvpmfHZcsX9KsUs8jNRKjMohKOwUwfNbvdtq9c0+Jnjk5tYwoDPkr0PBJJPTydkW0xVcdh9MJb
7xBDVbfIrt+0J5IdKiDDOz0r9LWIJfHF+NxiqscUJDFpEQhE3zyj5ph2+aKUkQi650ZTk/3MRmD+
FbkvlmcBQip7jGIFMZ9E+moLG6T2XqB+GEAV1s5HWHCImjRqJdxqtVywIoV5R1/Z8FSS0GJMgUhO
e5LnOarsYlmDINZHIndkl2mb/2STvT5jzHgwAtdl5p0aJCPoNRuGNy9FygF4KYMNGZN/oEqDEKu4
8vGQmJw5LWxrJh8EkJ5Mn7EiA5orSqvQEO3UrJ/JtOTV968F9xWF4QRqVmenj/de7VLm2iv4tCgE
gQqmlGPRMjAqxbUvwRG4LeZLB/y1V+s3IvKfVKqJEbrslzKU1yA0EJcUmZvFVsuH56Vbo6brSzIL
Rek8KZcFDupMaIsZSdMc/53kEmt1zd/xdGut6Py1QE3mxPuAQswpvjDBcLPsGZ/w5ZkLnQLT9N0r
EDk1XkooXYxKlLQq9OUkW57dBjj0uNYqUUOfv85ATR+/kZW8zWwhsp4p2UdFbbSeH2AdRffCfPo+
Q7Ya+Ypj3OF1Y8UwgNNl8HWr8chgiUI8QhF7/LSm2GqQkCBISHniZHlIcON/S74zJu2EZy+aGzJ9
Qf2SHAt9mkisKzYYh3I29drgmJMbNJ9pCfGSUcB+v/Lulf4OaNzzuF//e85YmGEgqR1lKJufPEj7
ObclvBPvZppl93IbrbJ3rRiKtJsE/0HtG8EDPqP3OkKYACjMLQo/jmFTX9Fh1r6Lzu9+jsSJ4dA9
LiD6FQXXL7M8Wp2jSMAAoPKJe54zrH5N1jTcDpX/eK34zHoyWZXU9M9kslNHnuXWMURNm/iv20HY
UjAnR1TWUKgGgh081U7GOPsaOTsR1W8DpZmkgiSrSQkM6JuK7CqkXUSVOgvHtTI2HsJ2FBZ8QR61
vQj4REiLsXY7ztpi4vE3wqPiiil9+9TgHpJjivh/XN5DRaKPfNGQMeCo3Zi2889RopZmv/CrRPlc
pMLgy6vaTkAT8vGmIrCzaONOZi2oWsJp+3dykLn1UbV90I3fM6bK4mP+7ZH5Ms013rik3Vc9b4GF
yTY1+e0aqGwy/oSZlN1Ypnf+551t2IIp6gRL+R4PkJkwZEwOei46tIMlSARlcT+7vXIMq/Yub/1H
JYX6K82BKJi+iICnBo98heHXrIWpEcs4dWPGTuizR736i1cNlhQs0b/8Kig2gwV1Cu1y4hJfyBLa
NNmy4NBrA+BHIw1oMar1DucL2sI/u+KQqJXZAaz7KTP/aX9kzgncG6M0RZjQQvI8z+Kn0o3HbEez
S4c69qTp3WWe8wKvJcVs45IOF9wl+b7ePaz2yibCSrk/XSk6F6McuUdWPBe6JA/6GauygvGNBguB
313W0HWBzc1f2blC+hBD6lSXRD8ipnsaGkfULiWMQGK8IJDKfsDRCOy8Y//+vBIOU6vhP9kuktwi
/sAurYn8EAvPqQ5WC+mMtglkHfZ0KPWPeyCZuxVnL+aQWuNKu9+V/X8yRXkHhF7wbS4FrR4ckTEo
RqUTJilR+7Oh48hOv8lQjsHUwFU57YcjnjrdHjDyKhdr+OnendEL8J84c18ae5EqJAKOKx0ck+Ow
95le6MxezY05EntEbbLrWpmCPGBkKMdQxpsLgyBLxsHgfrVLOkOCVYZiSr/ETO0VIYO/hXnSTIjh
MPKeRZIcITnKKk82OAPQ9tBkbz3sl8ty/lsicT72S0z4lh9mj7B5xLPhJfOAuH+8FHR10nXOMr2J
FPNWQv7dUHFsFAqgu4EwhAA57DB5rLOWc8uXx2BkAUsUCTfGAUqgMBH2MBOXNbCGh7WJ1VZqWLQq
3SBTam4+b76vwN/Pr7mtWsC3Rm8MWN+zzGfPgldM/r2DxRaTojnNc3VxOw+YGIYJ6qtOeI7bF1w2
4eSoASEcFRc8hjC9PpqNzQjmZKLmqzfWe1Hz4y3T8JRtxHIRsPTTvtrT+smwpqXitanp2WUSWoAD
ghujyAp+igjxIjmfUuErHW24mrTgkri2kUHCmu8SBoc4o3rs263Cn1syoS9K1XR6+d8++5i/sP4v
de8fz25p7pFZCkU9NReOB4MUHcEZY7CxYaR3b3pxqJuQURcqZM5jJosTXbx96Q3twF2QycGCWDp+
1aPlrVznFvZoYtuYJt7O+EC7zaiJAL5gEc16BZ8ZeE1h/0EsL19r3rez30/5gKmgItINCUjvcidV
jxtSu5v7UiWBm3oISy0OS5akQBX+yZKTVjS7DPX9vwi3gDQIg71gXsoeMMfc92VzCJSsmGHTBed1
d0sHRJjeXjjYIoS5z+U+p/NPzLnbbJ7uLReIKQrhJvqt/VmH9BHbEV88+Kzf8Fh9x1YOG+bZ/Utc
sgGPsIB5kp1Mba5hBN7X76AkakOatQ0Uzwh+6A3CHTUsdOmubbxLWQ5kyNJhetVaaEABvRRKGNz6
OMXV2K1MlKASECM77mE3pP3VgeA1Fwon/97WZTjItMaY7RLGQnmM4eIlPlN2ham7ySjkbgoymH0O
aqt84aVIHZ8OqFHjAG72MvYGZccKx/SM6Hy3gYnl9tlogUiYBNZKXm39MTf+o4aN4HedkEZ9udEs
xV54h2ThZzHTu/UUaiNFLQwhe+yFs/j1I9KyEC6/ILSYHOFsE4VhX4hI4xoM8vIc81V7mFyL8B4x
P4TkE6QHB8f08CHe+FbW9mFzEr45j5ZMswA/cUpVfRBNYHXyW1bCz1AlxTgk1OfIgCysZaOgQME/
0aP6MSePGfAM25OBQTuM5LATLCGzaDp6zifrrZpffdH8xpvlXB7hhRi74DIv6PB9pCNfGAytHQfl
+sR7oIEoXdyy4W6N+xTzbqwwONSaMa+sODq+AkPQpRwalGC8w0hQOZL5pIv4ZK/Gz3J40SPGQin9
jAcyLfFxeftbIUCTJLCGRSFuFnydn4YwrnsP/JdQg6g0nk/7S+bNtMBxCPnvqclMpWu9/hS6FBUg
lohawc9+D+xiMdya9z02jUBiXcTmqFxLkt+fsav3uZ80j5Gsnd41xacdoZKHUs8ERT4H9PR3D82I
lLp/s4AQGejfaJXNDwRpyQp46ko8MI4CdVEcy/rlZDx9U5n0KGlIpJpzHFxPH1pN15tiv0iE2KcH
0oLPjwtwArDuCyFieoFaonXhiKfp//4z19Wkfni5wiEC4wMFbyFSoFsAs0SWwaaSBebMQICnHsOi
BbVaqQX11EklZCHvsNWE5iF02ny1HJ7rG6HmSH1VbnHRYD8suqGpAbYBGSApLR0RyPD5uXzE92m6
9jk+nFUsfGmccphU3mWRBZX+zEXY8Cxodpb72Oa4pqqyxErx4yd5ncHwPvHe8Lgeu/W8YPETErGV
CVGWBmUMsUNrhbeNgKA1N9nab1DbjOx3AnbKvUQe/ZosHqLONUA6YgYEjxXxfVtmOls9GAkfuBZ4
Ep5yiA9AR0k3wmjb2jmW7txafigFFApaExu8z0++eTmT/hCXEp41GakoqZ5Q9oEuk1xqg1zT3i3A
BI/yS127v9P05QoW9QkobOtKtkyVZoFIAGc+IgAl0IoP69YWXBqfl8rn7jeK/Gb2DXLuefk65lNF
/F+Vytji2MNDdDF8WF0Kr+6oXcdL3CDspNc7idwFl75frabH0ndoQaBABFW70nUtSxH7p333nGlZ
SiTabRlI8ahTGATPWanAhpdDhphFKAgPjP3jwbzoQ9o53IO57UaA98a/1R0e3HRHJNANfFlvzy0p
Tpx4pMJvrw3jXtEEemd15WRG3qdyR+js5DKBP0GEyvjJGrCTXljqTwDcaEliEFLWBOsoTOYWUaue
HltsVvbJGUXvphgEQJsXuzkCb6457y7Zma95K/Hs3VvFNwpfR0AU4Gkcc4bKA3gW9Bp+elmyPFBP
vtIdOcGLAWnEUTuZCK91AhDjynoc50PR2i5/ebi+vKhZe3s/XBC/VwqF1yeQwnOjfMR/tkQS9b62
joqlU8VFPbDzM+RpYXSDmZxvUYQ1lOc3Crit3CkYq/8C6Rer7WvwEZ42mnxGduT97b3RitWJBCum
BVgV7LUO9wRdmECYf5rtAtjirVCVFXX8AZocvKBea20o1yggGt62WsM9Bz9+OQcFhAsvxtEIG9tk
LQSogvGK/dRYKiEV7bDF0KHNeHLgLenIf4YSXLFVL32WofQalYfdWDGxeEII5pE2S+fVPHGVUSdS
0frs9rZHyBJV48OETMU50xgPm3jECjny/W36BejMA8kgvUL/UevVK+QfcAljslIj1bZcZDfN/D1+
W6SyNBD5emNKyDUjRsbl+wS7kdZxf8GOWoad7jWqmSTZE4phrt7aQYsWhceCpnt3F6NwSfx5++xI
DSlc3FBRz6TiBFk0jdEJ5Ym42dNrLFRYSP4Xy2l0QBeRVz3C2ig4ERLS8MupowVihB1zb1fQJyIH
VME+D2IMmY+r7ZPAAxKEvTzE6NeW/McNDjzOZoRpDQU1plwfGYVR1XTjbTjv/4+/I4GHRs4sofIf
BD0BCUx96acIp689Wjaqu4VUOyWtrZu3C4BvPLSnlNXi7TYRjTatqzuGpSOr4IluLjjS9LUvt6bW
IRkwlCYF9SaHwulcpajWWlkD1iKSCYHPAICBdga4H3/5oYUHMMOqtuV5TaP3GAuyPFssmkWulwFC
I5+xNHI4I1ZTf9t6nc/ibCCBmvO/+PmUW36w4Fr9EWd5ZKoFZHo6yFriDQG6eGlTepJjksUYFeTJ
zz8VCnlv0DKY+pGfLngnQkzMe3Du4nrEs0+wYTg7HY6g8BVeGAxxFlHzB9u49MIEMO49Y3zXxNZL
qmbXWCFskgzbA0phS69na1PItISOgg+/GJ0sVEwAQO6JbxcVNHV03uy/PB/LZBTXCNeiXWvwUlha
AHogRXj/K8hgmZvWTNA1SEkO9bpjfhmYIBCigOimbb7gUyVHQJkFO219tBPrixww4HP6yQ73WW5C
IAvPZ+6Kyc2GqhsCXjsdQ5fyA3iQt9rFwZfPoavFs3o5iVgzmLEkBOlSvQSi/EmHoZ5ZovB/aMVK
vvAdkofG9qurOTbnGUQ0LDqEQi03mwSqcdsXsfVS3pyG6oDjPwce8RyMfHOl/0oi7CHv8Kkr/50g
jNsuVCrYgABOz6ZEkIXIczMjJDBMMQ6CdgnpePv7uk8UbpMIawxCcDXmvDsNHIJfZODA6z4HyCEP
S6zjdqQnIHepnMeb81ubmG4G9DV7LNfMdQo+B0/3QkudqNrcD7+1zJKj+dfchU+dRvk4RL+jlGU6
GH/yHPI1QLABowiWT+ceMOA9pMDpIES7R2f81PECfSq0tCmf4NWjSTkwKdS68GPXksNYJH81ohud
BYIYNqIJY/5Ye6U21nGSQVQlvtLeAZxE71nXsZjE6JCZp9OAJk6xAkWTelvcZ+tafycbUaNRhemU
avn620XQfyYxxnBZIEHyIJWqZor91CYYraahtDidwtNeddUp92+HPf1b6htD12W1lMtDDXZeX3p7
JFBNA2MjpDh4e7Mxe4Q/y3smoPrVuhK3IzsV2tB/qgGoIwUnFl6qx3JdmVB97/t5/pSmkFi2/rl0
m3qa0vs+pXfCR455J+0GehbNJDLkJvwNxCfZ7kQa82jRVVwyZzoD29LHOex7d0i2sNdAvdKfj5K5
qnciVqbz9LZgk4JUvhPxTQ9CelmmcX4blpSuEtt3uYJZkig9dQUX6sfnG+DfY9KX0KDqzv6GnJuV
YFBSot7EZqvEuRwOVZo9l61s0VO8GFBRHl6LG1fxbe7+1U//d4/gtExOFlhGm+GfDnue/rOsd9xn
muz0dxh/Skh90cAK9TuN+9cgCDwJjzLH703GqUC7WqOSLW+zEIyd/k3gOxmrDT1TzNSvqEMbNXu4
KBZZ4Vlji0LZywenbc71TD7XbN4NB5KIHcqfk+p+NxAHFPWwYVY8mAeyza9NDy26u1iWVMA/cpZF
oW1aQTUVgt/gyKwjPDLuWDcaeYpxRIVVvTFeQRquJ1VGm+mIMycw6rIJc4TOCMCw/qyvxzHf7l/b
mQOxEU9iTe7qyVPKcurpwacOk2guipHgoLJKdkAqrkUGWI8XEcoPtAKNmBFHZJZWG+nA3esy9JGD
p5LxfsaBREcYZaniCW2TRp+7iy+qgIgmjKCu4fYcEjLvWmq1tq8kUBBSZ9G39ohlqWdkucV6KqKd
tI71CMzm0ArR0PJbcHTF5keOB/0wCTRHS0Cd4hhba/Y5ZU6v/PkjaTUVzi4zuXbAplVgxXuxFnKo
zoHxBcPNijYFfJOjNRuyvx0WJozCZpdHPoYHUWJcyKkc6sGexQg8kuZEIDXZDjbLC7wDRsMFbtsa
qlNk1G2aAm6ZKKsC3v7WmJW11rPaamhd/dRnF5DdFjCuNfyK21jfQ/xZpmBfwvzqW4eI3A2GtfaZ
BmMJvOAQJnWpPsi6laYZE38FVpxDkp42gdf12eZBreOVbDgzJAKF2UMcT5p68HmkqKGLioha95YG
kz6vT/QY9imbz2fF7BG04MpMdU+edmPhB8HYMBNZnfUhlIME2pAgtBQoqWHqeBGipgCcbCtKWjvo
r7uthVA95rl2eXIiCBe7HPrfy/SXNhGBBNZR72rD+1Il7SgDDdjjqBNVDMuY7xbxwiqz1FgRxtxO
bvJZ1fVEefphcGxQcPADusa+XJzOs06WLHCA81q/nKG3/1qKBUVT7FaXJ0Qd8Xu0EP7M9xeiR5It
5cLIgU4aNtsv0ZBIX20adN4tM3p+KPOIkV5YWKG6XLUFzJk0miPhVWQ3/SC++tAWV/Bflr8wtA8p
FnU+d55HVk0wCkQRrajUP06oLo3Yag/gqW66eMApS5Tmble3rlakr1kx+VzpG0txTqADzbH3cLe+
n3BKDEOShMSfm9fUErhwFwySNY/HJf1T3rMwFLorxA4wur6m1dcEotlHSAllz1pP5KsZPqJ6WQwL
s/pJS4Ze3HO4dY6NpMROySgbTvne9+J0YRn/wsoVbrqtGApSKGC+I9Swjp/6jCy2ZYkBahoXiBdR
9MThaQi8R/QniUUh7gowK3AmS7Y2FdApln7UdYgdFGRXlqub6gy26BkxNWtiwxWpUX52wAS5czZf
o4OYvnHg3714Dw4NSTLPYaNPklvdSssom18+cnjhCVRhoo4zJuH9W9VHQ1Kx7YWudVuecGNeOvKY
1NIpEguKdXYPnzfyLSTJ+0iGGCQzsDM4Uc4oAh8n1gmwTyg7rNZYbl9fNuO0aYufEL6V3AWy1BZc
aXe9AzUglbPz2ppb892HSqPtg7S3x5myXcUlghkTGe+LhQNfVOttcHRmmHNPA2sLwnYDE6ULv3Bb
aIil2QW4z0G+I8VSeB8E9IDc3+mfUo6RFC/kiuBXFs1iQ4uciJL5vHzzB0FkiRpkUepne/xIwUzu
iiw6w1/2wK0APP5gECskG5iG0JlyCYyeI//VxnBfzoJo0shPD8rwSzKDY9V2oFK45/QXkJGKZ/6z
ZfC1FdzMfa4fr3/Lsqcla9Y2hYcSBLOnO38YWyJQUC/w8sxd0qFV8J7YPVZmqqvNHzW1DtYhW+Ks
7q2ITE3Xlx4H7W4z7kz9LCXNmSpWM4c9rhd+Wx6ZeyvJw69XIDMA4QjJEoj3zB7yLBh42+Gg4n+q
WYj1u1ee4b9rpEW7TdDjdSFl8rBC4Sfj72cGio49kc4JnCASeSeSgiU1q3M5VfZloAlLi5zC8L8q
zRT/1WlFVTJyeZ+DbcWmvsjv9bdWdP5gJXoajLQNpyyx+I0PXhWvTDX1+F90+K71lfP48/AjTnfG
ZCjEia54eyepXeHwzmWws5MwhHJ8Ws2kTMsBrcJ8FRYgX7k3J/nKPgfsM823D073oufj88bxfWmg
fLuaZkltbvL9HiL7rY9yYdiE/wSxZPV6sL3IUutxel6ytnnjJTlflAeKTs1EuvaUXQ6OBSXT33Hs
J5iVw62fKw3dlLagamXUIx0/PT3QVQ18gko5zWUpU5ALg7ntv/LJJSTy7QKzIRzfH6f6PvknvZt+
T5fOOcBHAiHzixvHcTQXnVSbYHkgCvJZgVIRwR4LH8xgCzz9MkJ+CDQvbd0Xx1ZQIIUxEBD8N9Yu
rWtUIpAvL/EHU6C6XowjjflTg8rdQvx6fPS4pBhR+jJw+C8qmz2ShxFvDlZ4JsVBiKqTBkAa7vrw
b7404z3Bh3VHruogRACInONeuwV5fZHIhniVn34NKKvICMd8mEl7LHZw5BrtJSVLNyHPrAiGO+Yd
e66PcJXliWHquukXhY339e4Z3V+E18Lg8qFwgcFhfk0FOWqlw2J+hU3pBcZTcSmnSFLIaJWfXpJo
VFSfKwharloKu+NgMSIFV1SJgZavU9EwHF4RqSxQv1GuM6iN30RpRFjjbD1iQIE4AbRoKvDio3Ls
fMTKQGzh4dVspkbhrbcC4m4rsFbRQooxMCzTZOs5lJuRZhIm99nXGzMUEGqXlAG5bdYEa0ZQu1XR
m6VEujrRbf5HiXMVHokfvArPSM4il9dLoegK6FZRcQ3BircJhbth04/k4WI79TuD7f6G+jVK7Vtq
O27za0MWvQ3dOIrPpiLBSACLXLFqIwev1hgU2OkKV8a97BxgIwvJ8DI36e0j+cogWvqIvB0d40db
GJreqa7L3yFlHqDqtzrGgar/ZuRYWk362uW1U3mqOeRfUM8zYrTtOyPJauijxuvPXNslyBpXgWhz
OxtlH6Fj9fggDuOP+TPqQO0x7p5HhHW9GYDiohBmoomvTzxDemMwd1pQxNfUangYt2ZWZNwG776d
fCaTZ7dt8de3+vVIeGIFmQkllUXAiLB5oqP3Uq3VtxttoBKAJoT3VNgcPlPHujFCy1Vmg7yMP+Oz
1TU1F8oJ1NH1rkoj8oeWkTJHy830CVlaH5fNrr7eqeVSESOjLlDKcjBvU/BxJTPSlUl3Qdf71Igc
f6v8KqYnPl8JzfNWlvWDix2NU4ob3ic6XMkPOz8VRXuj8efMgi4cF9Mj3ovUo+iQZxHSc3ncxS05
WL/akCsH7/0yxC+sS/aQFC3G6Lwz6g+ZJs6yw+qHrZXiMTJCwu4LxEoJYUeukEE/90qBO8fJ4IML
Ae70H8vo1vOlSENNh6ZT4Tl+gLFkj7zrg6uM7EQm54dxfSf5oK7MGNGj65runiTSsV4A6neT92TG
55GXfpk3i5tQUMJXY4HuTQ7Wveo7ptWiP1sdXhSda5BcktyV1z1vPsjaXo21wrVYmTa9lWTQdbC7
Zu2w7HkHR8uTz01Tq+coz/qW/cfdoXjXETbOwoEe7BPMs9l8LE2Qs3GyGMEUOWvgYReuzrAsodBH
kmNhaXvW9GkIVfurAiw/LTIF6u+v2jv6udw+NZbOofcXZ3umJ9Z44JwlX/kQ8omaZKHDCdALBi5z
JM2Rs+9+dEmJUJl+RCeTUq7XachJn8gVVyJNE38gYHEUWaW4Zd72uXxuKSg6rynb1RLYxjcnOrj1
WhBjRyC1vjAl1rXWVI8fl5t5vfWCr4bY4oVPCqf+l7LSmg5tLW7Fg44WgwN9OmYmaf/JsUtAp5nQ
ZZ3ITv8wtK/l0u1lNctBakvLmTZXk+FIgmwi+/6IXCt9m2sES8ezz5GaJd6R0drzEbXcR73DNaD5
r1XW7/g4gU3A+HgQvkGY/2KgDDuS9TGHV1bLF2JbaLNeMfGlQMOkv7atK/s0NPOQZnfygV81TKwQ
iGn6unfIPH6gns2rahWOUBHuGvGORgVHbP1bzPpoUag03FvbKyl7qpx4ypEWaapN9lAMMbMcx3E3
KVB9t8UVyJqKSbDLIMYhb8Rs5QSClyVbienokvFsfRTVhTk2LNzbCdump7Go5rtPUffNw00Tv2+m
kP6FHeSiEg57ZEWwRbczEnSs/FvPptoOraGa3tRjljZR/X/mr3rOk0cVAA+Wzw8eNbc17pmdPwFD
6NXv2PMfIwvAomj0VAFy3egY0OQ45GshHh/PMR9zGQ1lKmNHAfnqdKF2UyJowIVYMgOlPFn40QQL
eAyx3znZykjkH0A0kmCCo5H59vOwe6UkKHje5a2XbksQE76pfcPhbbFQC0ZbQWMb6y6QcttfSwhG
huhsFIf7eCSItGIZL/SyKVrvSlPVxJY9s65AU15WcOqzcA2Q72NGOuURlqxPlrLEaybsROU+WvH6
uiQChAMgEGTLOP4DzZvs3nfYbj+8x9OnlBQsl0ChnEtiUxqoXzWrnJjF/1V5Mb4ykLFiqy4ZjVJT
xb6hnlPBSMcbYaLZRNrhPE1ic0Ij7KJTqOSsWQPvie/OCPL6GP6nPXcJVDWrD+NvAro2BwYUy3UA
9NsZtoW0Jd2Z7liRxIbwLU6zoYoR0CpJdBjBu78AyyqpBGJgXuZ2BiRtYBp4jsxoHHfQwifdMWAP
mXBFqkZ720sZe5o/ZuAz59TTolg8GCiHO0tsHYM/yFwMMX6aLKwILkxE/H4jRJwb+iL8cCIe6p6p
sthfoJ0HXb46oEvc4sp6H8azXF8tt/nWwWtL/hKodY5QEnxhDHqD0XqfoEGk9eUZ01hB46aEIRAt
p4vpVkBOg8vjenNB2Z4hme5vPEb1n61wUJgoE+bKz3NOc2hl5v3q4EQTLd8jt5wCtici8HedmEev
9yX+BjoIogsPf9dZu3oqP81qCnJGImwIASn5uBloZj1n8/5OjrRTo7E/xBlnsjjxtvIU3wk0d58n
ZVns/V+siD+53QQgGu0YA2jQzTlWm9rfavEBxDKEMgUJlRDTkRvbh9cKOAbWVfn2qVqoUMXt6e/E
J8L0PSKSViecrigiP3PY3hCUGVT5fU8jth22F7CFg8rhgFEAS+WxH73IdpXgGSv1tWXoxLCrVzHn
CP7yJJQ3i5orCuIDgzxb7oT5VH7xQmP+12s7YNgMtbCHs24S4RFPEDCvGXmviaXpRIvy9ZEE+SnR
RJqx6Gluu7lHS99khImgaHLBnJPUaLeFwLV5tyDe8Wr/M75xjYpr2UWJqWFuFW8WzNQVy/gOn+Zp
m3xDgoD3LEwYl9Ddkig8sXxjTAcMHVAnCNNubk50bGIspykGNU/9Zkz7h7xeEcMSwmtjHYouQgmf
MjUczVgi8o6YaHexxZVjL34VLpRg6QQtKWifh4vqEfIa424+bxhBAahZnzjScH+QMpAPhj8gzx1T
veYsosLk0vZdHiU9f1jh3UAs6LeIKiTevcYBuMQFd54Up1fcp9MIuKnsgCPimDPbwiyha3KBpaEX
Q7tG4AM5XvkV/uBJ60Y88v7KGGWKjS1mXqUw/q68ZU0upNQOdGH5RBrCpWVH3WkFxxPfLhXehV90
5As0ft5/AVRlh1n20U7Tk6QIPxIZsQO7pnizGVwPOAA0p4poSiKkW8feIax+6BqfvlcLTkQz4Vy7
J5pwgVTD91r4VGplpSayZmQGhvFuRjWb2RlOcOzO472SKSfiXdPRCcqRwd6F4zgKAuLKfgUxOjmY
2zBlOXCdKMbA/Yws6dcinjZVLXRO0VbjaPoeycnIfEcOiGzXD0DdjZtQ2vduDYaB9tPK2q7l9967
DNNp3Zu1Lw92SX29BNEGAHwS5vwCXQIvtGsjyJaBetw6Ce3qifQgkGv3+t9PJI4emcR/2+hlu/Sp
1siBNIKFxQxBKLx8vo7w+5nIImIvQtiD/MwLX0J8cVw6TzKzGqDPslP/1XP5HurYdWCdlpA/V9iw
EO66dI52SUzKPXzX1ErT2RKctiTU18J5e0Zdhjz37Zkwgya6fYh9CBhBUvAVU/0ddV5H4QrKPiTG
j2+ly9jIPNh2Bw26+VewFbweno1xr9DB38WgbuFWJGi3Cb9G1WYv9swF2VW1K6/yhGG52hIIM4wQ
96hZ316yKMTaTfKIa0ppAZYgw51K5Ge2fhNCzT5QWCRg2LPRl0g0QAE/rkV2pjw6y66PDIegskXS
g8iDP6fKMK2nGxlFXJchHlDKJLmbCbP+82HOQWkuXawIk+dUYNnm5sMkSe03M68IzS3z6bFs3SsE
/l6sDTPwJMVePZO8vbJEEqlNuj/62pcabrkswUIsWSgzYWTIN+Q02EjBJr2xrGeZb7OM2Oqk9dUK
pKcQxpbVzTQA/YQGP2V0d+v0x13qZSw0FblBPJ/HuwrHMSZ8Ad9YWEYs0ZZCRJScqv6C3qJzBAHI
al1EWaLoc9TmfuwKgUWGEwG1AO4E1+n2nywLXNixcb4nUP6rhx5Ib3q7x6SeFN1kX+pqA7osUD2m
c6j1SfGorvxclUl+wpsdDde7ty78dYFYl/iYJ4cgh8Ca/xrJKfijG3fgsA12LADymKvQ5FDAZR+O
VEks/vW+pu2crmTP0rFDEv+muFs9kbNmTHh4VBBSkXclCG9Kip992HBbHzLjgVQzQW2CPyXbIDCN
0xdjH7ielEJDLNt+1U9iHC/HmIP+l2IPxbeWVCfq4gCrspmwoOBCX+KdUjeh4KByuVF+L0thL8Ax
AifNLDKuRyvCpoWwmdTVXR5NlbEC1Ng3PywVm7Re/ecHgB/b/KIIwtGIkMmgR4enDmE0WRIC7tjh
WBWb5UU6JeCWAGzIE8KAoxb6AbTI3EMyEWzoz/lhMyhhtXZzVYJAU4N1adGu154Ol8DhPizvM3Kk
C7TYbI5H/+GKs2lGcVfu1oSzdBb5RdYX7QUMz+g+AS7k6Wojo8o7adKSvBqgL+B2S0EXmCooUVz/
+rfSUOhstBFVUcUlkmLlreq3tvfw72laeK+dtvbbeUctOtWiiNVaaUWgoFA1l8aVEUMtAeBIRGdS
51SSGuOqlrWTdolrYNDj/HNUDHN/vxtA2ohrlIU8b6rRxiLvCLiNNCcCcLzoKuebsVpHQJmjs1x+
fbJtJbpkA0WW/r8bKsnmojpigskIEQ3/qv44m96VeY+b2V4JLz/kVkEhxvl4qU5I8JuIpoDP7uL3
fVQUgU7svWlrn8RpPFPKPve8GNWErbntvsdpcei5TuL6vBuar879b4GsM17CF3FrFBFdhPNoTjTo
06AtS70QNDQMjkzlg+rZQ8iVZH3w1P7wcaU7/NkIij6+8xW0Or+wlxL7ST7PTeBrTz0nagAw84j8
dHO2Dh41MelKAHC9NXLg6aoHnRM2AfjDuOD8Hh/hcGEAYj8A5BK0OdoHgeXWZ3rJInTZzR4qaGuT
YoGsq7qlTwHC9nxEX98+enUMsFVOtxL97dlibjKzpdP5w8y37aiMkKWatGDMZG2rNlDiIe1XZwE2
i6mLWdFOZ0hmzXoblTHsyhxHg0TVKB47EXC8iev6xdseSP/KGTYsZhzr5DVoY8baaDGk1nKYd2y7
orUtqfWXk5QAZ+Y2zecWMWvJoP6fM8pys6JVXEWhRPYvqR0jlqRUwG4mRcQ7J6R3mHXvr4PC/9YZ
d2kxkcBe+m5vZHArXvkonu9AaOmNrkR4G/X6L4e9owdwd9KP0PS4/Qwc4wsi8DE19rpeQac/Z7gr
UfAJK0lenrasf1Cz7Nx/iOJ5YxluthLt/7WThe7vpdHTGwPfhQQONmb3H/MV0gN7msT8gNWrqdGP
AZY+uGLT7cV8pfHwQiVbe8OQrXPzOO5PyTTPv/ICq4+wFPypSaZlO3c7sff8V+kbG/hHX+36rdz6
Yea7gPny38fxhMII8Lo9aAuiF0tv3ICMUZ6CBx/fqc/VHASyNNcGVp1o+h+0jwVaY85z0RXRIv9Y
heMWxWpyMj9rp9xVgYIHsSFjjCbBx4ruWurg4rXjyIaI0Jlex10SxJOa2XK4wpmMxPRFZOFCUM+j
whdyIlPwF9iNLEr70jjjlR2AGLwV+Wpsv+zW68bHuWn2FJzRPsv1cn9YIGCMRlN0wn5BKZyrKjrj
YM3Wge306uubU5eVLdls0Zr08olPFFfQS2z0D559MreqowRjFjA8FISS2b+WcubMRsfUlf08TZvj
Cy2hKBFhCJLjWTAUeMGY9VTfocC8Vz9KDymAuj6swE49dEur+hHOMAP6wxhzoiljCIdSckOWmI8Q
PPYn4vRkAAr6n8FJgtV4jHXSvHhlqBcvceGvTGAiwTb/m0YUucVvgkpCgomy4u9Am27bqeLQwv2y
DjXFXUepr/CyNsOxvAGubIHltpdJkX5S4QUevacoMelne/5NmatSMWTGJlazGBtLea2jWdhAWrnq
d2aNwjmMt/gQxlqFyTs5eRYZDSs0DhrlcELM723NBmQycgs8ABwaxJXX0xMB7ZcwGuSeyLj4QvjE
wIhXJWmbrnrSKweR0GQ4ZC+U4QwnXJuLfFUgIZZhKpTDoAFfGrEdT/3YqX+REqe2biT1NqZU0LxG
8HLbOoHV7ZobkLPzOg95CWEQ+cNBJSq677RDsKGXS08TTBJFW13+RUP4q94fhNW0bctY5XxKDLre
yvorKjRcrCvSAFMe56B2UlLdqku2mx7G1DNFhupd2kkSkhNfmknRjtu6PYu5QywFbajA1MCivD+R
eqQecEX77X4dj1Q5V8JiWSXiEoezUzRLf9tzi2dGHtBX1HaL+omTeEVmejjigk8ywmTYR3zvIVHD
+WJAtTE/iztGIwafud8cDFhP2tAREwjHJI+/ubbDzeLLHJNMH4xbQ3fhnBuVEH1cSS7jRCHbYKYw
pMaoqjjxWABy6GycJvVAIvcBYLrdqZspxTGD2iJsMNWDeAt5iKAVE1nRXmM36nuxgGvqji5sbi3i
svG8POKVjJ7G1Q/XqUekZgdMlCEtH6bGb5Z+tzsfXfu9M98rm/JXR1QUV/80HMK9JZHJJX5saFYr
hi+FUQljX7TUFQ/y9iTH7g0uxoRkmZreK1MTZefeHA3pU0xQwkAf4XMV+QBHs2IlDb5wnbkdXAYz
r0mn7cLC/RHXU14PbNdAWLckq+muW7zMtqLn4vnWD8c0AaqlRinO3wV3PYVwRpmSnaGoli2002Df
cL/YvuoIUMZpg2/SVMm/U4pWkqWevoOSW/TI/vz9A1200Xp41y10iGPjRVHvMhrlJchMQkqAy75o
s48O7928O/cGeRnFqr4x+Px/7ICqnUO70KiUtzeyG6yMWYUTa4qo3rz/jI0Fr6TozWRQqJ18X6Uy
gS7X1HRxRQVEHbNNCZUiut7NI/Sbs0BwP6HH71ZsaUzvRfpPDfau9hI/1Me5CWenEFziaMfaio8W
P/4czFg64mcSQe2m6DA4KymWDjqH1owGqza37HUkBm7wX1JFbeHXIkiVLDTQyT4cBuMI0VNVxl1q
ff+mgx7gyZp2Ja+owQTWiiWGEUBd1iZdEGBi6puY7KIGhUldmvN4j+s7VB64Ltq/Z7OSD+vclTp5
zNoIA0wghGvvw5LO7DwEm7Tx122NGEzmsoEwttfxtPjJssswp+Zuv0lKTUmDaAlxKxsuD30IRfUv
2kNSiWrvlgXb6TE9VSTAQ2IzSR0v/dqntH0W6UrOLY5xx+Z+DXUvcapK16MCb8t/v0clSrzZQ+UQ
AJVSy9Ex3SXaWVR5sW7VTVc+7qYI6KJ2tWZkmWxd1iJCzXjn1apBlw5GIXWQ9Wms+Di67xonqz8b
VRqdHPkp+1EnmUCjpKyk7uZ1L90EFoYLzSvdpQIdzzU/Awgu/bdj0KrRmF9575UXaxfuj37OzJGs
5H+CdTxLGkT5VgyUSux5aAkBiAKpB5LplGk85sZFns0f3/19GQzBQKwp4aC5QAWM+YFLU9vqVXKB
TQRFT1dZqxRunZTi1aawLiFgQjsml4U46dHIo81RgXz0rH1kFGb+Av/SZGATYuaM/YzhLbmqaiMV
lw/Nj0LmUU7eswo6pAyZaDj3cGqc6rfQ62ogYh/ZNlgDljhgn4v6sqrtbIKXPCA334DS8Tk9PQwY
VaH9+SDNA8OAgAHZGmxrI4aQgcwLJceHcgn6aZKnrWuMB8i1wdXSvI9yhwda8WPHtNCdt2K0lEnX
3qLvnGqtmZ2WWdpYerWzjrM82iKO56ADFhR37Tb93ZUV3ifwBEwJ7bkRTHRMT9dUROYK0FRrltKe
QtLGWd0LZlOT3+KfLjI2WBWWAjrC1pDwdVs+kJidIWzMk5AxR1YJHnNrLoqOkM1C0HTDCNdhLrJt
v0Y7EJEsTBsJ9OlXaetBsZRrTppVcDIKsAYkOra1Mp01iAEITBRaj/Jgv9KKa4oP1hQLh55gKAmy
S6W/wKUEtclsjujww9w6VgAxa4gy41XusgWHFf5XJ3gNZe2sedRh1mJa00IyvSEKDw25wNbul52i
Q7hX0LHyj0TvyV+8sLg1vnKv9OVLTuGpoivu6guoC6tgOcrW4QHByc33FObm9ejPLV8jblsSoo68
XrbFVSd5T0nTmXbVlk8O6IVFa/D/Ryzg7xu8h9or8P0NfIfQoW3hdCyIuDAAiR3EUHvL3gDcM/n9
m1WU5uZZhId2K8Xslqs5igo7In8ReTDVes9vEhqfKXnJAUprIiFewjhTtFCWcRmodfGdmAP3aBgZ
NVtMeOl1n/ytlB19/eDYDrwU5Zpte6l+N8sgHy1jp/iJEa9qh3q7eYyqN2wRzmCyE0qZWaclKIjt
1lzZlYQ15ZRVbJs+zlCtS+Fz9oR5hq7JDPjRf1a3mgPbuNDQ5cqlnSpjQx3kw9cxCgy+W31AH382
I6TciqNR0zhcKeEDHnzSHVyMyhXzRfCMZ3QdHBRSt7hzQmayOtXNElxmRMNyo7erLpf7bSUkdzg7
67dedsK4fcM2vEFQmUN8V3OxNYZsi6S98WcIpL34TczoHDs2lnGGhq5Jow3cAZxG0kz03VmYHWAK
SXlb2TzfovwsxM7UARSiz+BKQcenWJe/iI7x9o4R8uojEy4MsqO+p6N/UDblMNQRltbZ8ufNM59g
jW7bnzE6KgvIRFWI7+5m6HgQdEqC+FTn3zBhVl/GnbIWZEZ0oY6nuZ82xi8iLuBw86NooFtxeooG
AfZF8ZLDqZi0iWdoI8/ucwtPbhO3m0C2zxcJvTxIY1UjHG0yESt0C6edPXGjOg7V6Jigm46RhyIA
sdDpERGqSI+hJvl1/wugQmH+oI2pt7KTVva7hWaRperC2hsXzcYPSmEB2Effmymq3HUUjoVgApNO
KoKU3NB8W6rNcWo6mPN9AvAx5YOCOJx0ZFh5cI+Us2rP0ECI2W3FQ0fnfxN5AqcbI9vgketOF1kY
4oJl2GIw3uDDnQXy1yIgqjCwtoSLkinsWnDBdHfiSTQR6IGJrIKNOwQUGz/BZXKWlrpJLWuCupyv
N/QXRBPWNgntY55H4ZwygWqul2wxoehKC5utE+fjWTlEmBBLZSKFID/qExJjRJrTScEEtibLfKF+
Rt0hKdOOJrJ8CHUmj7Ekhxd65IvdItGUR+qZ56fDG4F4JVTf7gCD5sdNCwyjdDSimYhyi6kQlumA
c68+ZygsLmp4E4rZ2+5UB5cfw8mAfWjYguS2xVdN9HP2cAxG4i/q3zW44J8NZvwuv/nf4yZwpi3E
iC1I9fHNLwMrAfz8jbA9v81bJWPNO3YXPsrKsp6No6Q/KMLGB4mXAEtz9S0m6ds5ctg2FfajHQES
2cyLsXT8iF/sEXHwwJUbtoMSWzj1/ZzLBAgxU6A+urie3KzwCPwizut1kEWOUgJlcay6kiTGilF3
5/PJqSoOvqDyuPTibZzaRV2shWCmq4zR9k1+yuxU+CLPViSg/oAXMSINSD1hlQ0KKCE9uk1ZzSda
sAwFIAUWRgRvtPPKFNBCGB5lZNUsmKrD3iK5gKPsMHxsRCGSkojOlSI92MFt/0Q3FSPZtv3u3TED
AhDXolnYiMEpv7zpQbgmHns34BwpgLzf6CoSYnwYGxTGQyJ0Rym3ZwOk2IQmqrQ225S7cvPTs41D
87wgvBMiUkCqj9DujZGpCSG08ygQQH3V4EJfHMZYPMjsxyT0yrf5hfl3gj7N550u+mEKTblrr8O0
NGoGHrkK0IZ9IuWHcMIj9w7MfDub63Xab4eJXAIpx+LM9xM2svSdpqDJ8LglXFehkjdUdHt4xb5A
WmfCDT6qFzfW14p1uoMdIg3XNHgLASdeXqROV7sES5ZRZxCL2mbFetSK+kTwRhRQTxTdElpJ3TL0
51Dm1Tu1HVF4SsQ2SoTawUP5G35bIA8RPkQ08R4uHtak6UrCfxppLUnGzqIZs2DhpDzzhwmzp1R7
+0Maj93Dhxm1D1b5LpoQEGIOq4AnbY1Bl1uj3DRmQ/+eUw0fCy2xhsFH5a5KfiSI2QbCO+HUesty
/HH8o+MNthBl/jvyHprM+q7GQ5kPs+UMrJQJfcHIT+aR29KfphxvmwTfpe6ac/X5S7Smz7pRd/Qp
alRs/o2WzeMQwUDtIB5Qx7TKI/litSB5WcP4XPATrm7USVR9c+QJSQpN4hi+TCgaAHpi4YBrd9cg
mSeGeub2TK6HdbK3/l893Y6N8FqcGJVaLf+Yp6xkG3tkO+Zi9OLvR/0BY6ciwYYZ0qgwUxZHMuOQ
V66f+zSsp2S3swRuWy//KSycvqomCpdPo0qtulLemFy/FtVirRDY60Dmc9WlZ5wKYCmqfaLDboGL
7Os3c9wJLWqMXGVa8wdC6Fg6QWS02uRKaC1KgZWYabdrro9dA9chDKE91Ln/kgGuWmkaQXYl2Fur
300Zl9qV98Ni7ZNrpa1nwY8XGedKnEm6JzK8ieqc7fh4gA8e6yYOA46buat1+mFIqYSlSxM3lVRi
j4Ur+qHkFyueG1v2ijrQSafmt/jNMEbxFlES2/fCg9LcBo+9TgecNN0RfJDG7YDTnniOid2FbzMN
ezmCzOO6ZDYD3QUGuBbNwEWZ1OiASo3VA5zg4A+6OIzhF8myzi+XdLaOvcjdxj4qQa+iiYUP/odG
PYIqEwAO3UziaTEeXTjRBGZjtYMoA0m9JknyUXoPNTzys8N1kD2+1oh/fchRAfV81JrADh1YC231
AGCkcgkPeDA12u/SH9hoE1fE+diIjsZFOZSHQgzIm3diB+/AND4EupKR6P3jmu6tfxEt7hpWxGIf
GNJrRpbyxOPb4AyAKoGJlHQV8ySW6WJR/q+OgzcENspdYsWXba/ASyNDwlDPuOtIEkIX9gynW+x1
7SvlFZHutVZLalgdOvHp6Do0lXn+GKyuoQ+wTs1+SHIlN2KQo/WFXreJyGhShx5mgLuIY5eY97qf
YIbYtuwCIw+QRLkV48b7i2opUzArzb04GrEu72u4Z7iFIcl7ETLlhdiAuBn8a73FUS3hr3Wkdc80
by95aKYEyqDhXhNZGG/eaiAaMntaKce5EZ4WFo40FP4RIlZwUWW0/SZxwsNt1oNiheKOj3dhG+Wr
rnJltbROhAno9IfIkapWK6rD/qj2lDhBLEbIbtBff9JAUzfLe3UehTuY5MDaJLWrTl4sZx8+nGNZ
UEeh5mDih5Biy+8obvovUwhW4/CFuA2Htc62hgnJBpElgY+nx4wyrhR6cByrC6VhlSsecz6Zo5OL
euyjNrbqpMD6irHCs32X14ewOadDGLd/tfUUFzAb8I8DDb+8eIkixeSpjYGeKUzStZHEBOWUGtVY
5BMSI3L18fkvBedfDIWezvpXJoH8q4/6PcCYfEPuMuvUDn+pI2+GLxBhMQK24YbHJ+tF3DWNk+tN
5uuSz3s4vO1as7lTFBI0fMvMi8hiZ4RX+YZDG/FURgtDEwmioOno+DBOJdHoFnpgmH9kMkEqnyg1
afpyZ76vZuUeoeDDLjqWlrPMkVrjigJau/OH6fdrHu/sheotsspK/iwbKOpFXNvhmVkACK5UA2l+
vx+uHztPNwCx+n1xCel2vJ2JrEGoFVIYO+c2TqMbyJFej03rWnYfkESIBtWlkwgmNwijExc1tOna
5HtiKExWmS/gQeR01DzycbGNFWzpd/vdzXkdpm0dEIPxlA0uLru31QCfKciPFLUxnJaHOJo9S3CR
HIf6Ks8O3PjN2C0WhJAmTdDlMGs4UOo22VIRVfonvv4ag5mLbkD/q/toDza0PN3bw1/GPPq+i8Mt
kn9Olj4Jcxxs2i/6+qO1pASWjTNEyw7BHyyxmmK+5fP6dZHoDHJtnxQEePXwrfJu3WXDzg1/2YaU
IrEL3DNsj6bBRUvTdYH+Avxq8Shgw2cY6yZoUufN3isUItuMcQFxjn3JiCh02Kdnioo5rdg0/Xvb
7xB5Flly2uJESIlwo5/WWPvTwvfibfv3U47O3v5uq6YY87vumvwQhNwyYqQ99lIfvCSK4pE3z27+
4d7dm8tP9rI3ny7VZ23JM3OiP7oKhEJoVopyNJpll+qVYvYtK13RI+lKHmVJhIvdxqJ780S0dqy3
BRVaEx0J8Yc5ULCPtCnA3a9KZqihxAr4hz+mksNbAVn7Qn47kuuTti9sXm/l0dIRHWi2I3/R9T2b
K/cA/geP+ynGGE0uVu2aCV/yVBH4GBTIsNpKBiZJvK0GOLJe5k07/BaNfCDgBcQJ29zjm5Egn17h
ux6NBkHvu+dHicygkXUyn/8tcELeePsnCMJsPcpi20eB4EKAj36cDAJ2Z4nd3H642ZqPC9GmchQO
AgjsgUhKgc01kztE4jweEs0dMmm2oKCs1JXi1A9ltCXJv6H/XNgV/a7rb8KciVe2ibfFEXtEHkIC
i87RbB08Y7R78LcH5/fRH4cFUgjNCT4RU+bzHYGPd8qkYnCJF0uFlhJboRWxfQC34gD6Qzai3T0N
8pdch+pAZiURMkI68/7s5jLhg9wLQlW8UWs4eYQGrwYi1KQ+C6hboywufPn6lxdbvP/txnr8okpQ
IkGJjHRPxPqvx0lHbueeo1TMfcAfgfHGeiPxUT/ysb2/K596aKUzj+hqRgcrsQch6hx6/Ic2VhEY
jwsaBaryOJdW7V2YHB8Q/aM1FZZo5mPYx3UeEn4+zB8UdaQltyFvsiB9yQKoMWsY01aYOgI/cRzk
lFcjqkgrsoemHeVX8BBW3dtXwwyuT5oMjh1yGFTJWmcjBhBJg5QtFhXhDxn57JfGo5Y/7JN3XKr8
eb72s9Zh3Jt+jfCKMMhfXR6p2a3Rqx2VwLlG4YhOg1XVmyjVIOCq44UaV+aylNmhpmBBUWpAlmMO
zZUIH22ff/7Uva/z4o6lIBt7QnAiFAT7lHFDnocflIi/GR6bV6SDsIaUdCzACfoEW+Y7yAY+rZ1Y
juPefPrL+tHedb7UGtdikxfDY+Hg1hQK7zphSKrKQjPYo04bfurxIQn+iG++wdV/4dxVvAwqNeuv
yoT8wgD3dv+4JsTVp1JQv8C+brAWFfCn99hZMITKdyJ4AzzmdXKQOh9UBxKNQEaMItOF9ZG1JrvT
QSy6gm6bBtCT5P78dhdEnKsUpW7JPkZt9ayf6zQZ1SfiqOD52joqVZ2myijS3+BIHjku4fJoIbzF
DUXN1uYoq3+aV4Jq/ziHDEUs6803SORi2+uPKPpfEDFXspY/zuLZVcQ3ZmoVFwTgsIc4K+oaM5GO
bPwD97J+Rlvg/PiOl2k73KnY5TQeZZIY2tGJHKpmq/wsL6NC8UX4diSzWShY05QIOi2RPb57LGss
Zkjm3hAxBTc1hv6QN/e4WTC+7uFO/5DnjQWIZyIxixKau8GeDSavnAD1xzyZ5YtUZ3tVmmNlCMDd
DOZg2tj6QiMKrVydCh0XBOYOESoSeQkUKGHtwIajb7X/g502GIZ8wJjn35WOgh1c5LoCzgK1YMSx
GADHgny2vjslpv69oN1q+LT+9LrGLa+ZeV+mauxN3U52Q6m4DgJQXcXvWGTz7EnJqPeZJAliyy4X
dPGpL6Q3PO/q39yBwIauDZrJ733eGDaMDOGnByMADM9mEU1aC19umrP1PM1H+FEuySlQ1PUgH4mi
dqHu5gtP0/0RnWqZYQc3w24Vo6tUeMwyqLRujizVpa/LPk7Znn969bX+kHX4UymilRdnQBQaOF84
CDvtbTUflSDuniQhjogFdIySDywmGQBiXOsQYxSCMmtUiRrRO+xE4cKc63TxzUGbxXlibGjaW+rV
lXRXFYZmz7aqnT2ayFGuJcc07Yqt+ZDdDzU55eq6ULc7t/O4OifqClvTmzmDVkYUZv44m6tW/vQg
LWOgRh/fYs3/FsBol0lycq3jRu9iQe4NLwILxy595NtYzV6j0qUqjFPGL0pKE9nBP1Crl6CVPlsB
KCHDu7iaydDc9xUeSwu49/3TW8d61S+txFjdyEhMQHCLZkNcNnS2V8XKH2JJ+mAr2Ni5E/sQBtVz
xpiogP/AV7ueT3irdcW51AAHilpoSYcMYUJL1cSzvdU5Yphg+F+FgoWnEMMnDQjd2MEbx7zPBSkW
LjLECNw6081MPC1yLJ4ssxWS2ZCG1zCjqt7zC4qQN7JbT7zRA68NZroPXIpR5/23b1j4R1vaVFtI
Tf74snD818+77S7UlVNsulH6hjtXlB7JggK/xRGfo9u54s6ohAcqgxcwDNPK4hlp8ckHgFQOTgsS
p+A2uDSuSgslJiLESbLnCxqbtPidrCb5deNCPXhfRoGW6tJpAfqm+nSu1LnKzwlxcq/nBUwLA8XF
t1GfG6ZHIz/VnvVilQ/YsH8xGqXL6Uj6isJMlQjYNDb3jWzwdQsBFYdJ7g3VwND7uBzEXM0s0ASd
rXVvW+MV6+IpmjNeCO80C9rl1Dh5eDnXUFaCODMPcz/UrThE/rIU/bV7Y5Bf0JqFl+ywWfI+pdqH
juFgXjR486vCfaadlyFdY8MLtP+otZyAhouUoBbCnlUXOOdr64yxD5hIu6oe9RstMMA0dmQYy/jL
plzGncjJ3wb7KH4iaVfEaYH6FGSQzPbWNrKriEhNYJyPWXWDYCY4pYt3taunNS/BgjyNDMdG+e4I
YL0SiTGTn2+tikx5qeaf4a3sIFs6tJHt9fTaujqS2bFiFZqMOYQBRN6Bok+cER+1BjQyYE2PYpDD
jv5Nr0Vbp4U1XZUfyGzl81LdgaM0uNvMcI4nxZgdCKjUTnwbN5kuSvuWL+QXX41GaUA0LTbW+WvH
f83AQDKV0ZKYAE/JFeg2J6U0s/k2QXPE55JgUMuTvBKmQ0QhD40Nquv9lrKpZG0UAhrqAFzCWQ/C
n+UG7XWDIvgqGI7StonfgLMtEEu5LZQtGjtovhzLYQNWsYOrw+2BRkygoci4pW7INw2SXQ1K3avm
lNU/MxtTmcG3pej5m8fad8RsFjzDJuEDs0MJUIP0iyWWCRL/IQ2zUJX+MxTaCwvgHhVT2qitw762
xGruXJY85URT5sPIWAUZ1bXR86jpyoEj5WHav6DJ7zSDmhK/C+NZkEsMYKuNZH3Ky9EQn2/vmi/T
M+FGiHtdJH8jJ9z9NECmM11eYCVVqBzzPShQc6s0GyzkxwbWOufKL9KyVB0txh48cDgQwY6906nO
6oxiVk78ezYxeSdJMVGgagLRW1gKrd+xU3UxOA3JP3oMrNamR7gOSM3BPc6Emn+2AQTPaQrngskT
lLuOHysmPvfbXyHiMDBmWten82GsFG95F+SHnqgEuwwKBHRUWDo3q75b4Qa+cj2nMJfy5Y2X7NSY
YDdtB0unj2FH5vqQIyEnYRfDGgnphHWlvxPIJ71w5pRoitXVljMAjre5TuBgJW5P3UW+75kuXJDW
Qn1Nl2gtHiWhP3WBf9FvNqCHTh+vA4rCyaJXBa9qqBvjTmFRLh8T00EvPR4b7h+JA7Jfc0HmHk+g
Uxri10uk8EfMEJYjQ5ZdH1WmQ1P3r31MIl97Gds0CDflBpvo8+7ya8li7ph5d6lVETlv8RkZ05sg
z+76SxoowRtB9pHoCTFjyGh6EYC/IUrxOIGmjObdLGmaEo3pVm9MAUrm8HuWKzR/QA2QMo5UX6r+
hERQMVAXfpYSFWO/MNI2w3PO7EPBe5N/F9W0KOFQUu5rghC7fAmu6XQ6FqVos3BZi72OnkTs4/PX
b+sX1wWGrWcUIWpTUdypofa6NeYHAjQDPuALzrupYLbXK0VJ+ONDfhlFPUCfrQxIHvdCXup7YxC9
hBvzsYxHiGPtzCebu4nCExr+Z82UkQkRiNDdSmOlKTrXlnAUoRvwJRCVtOqNRav1bT3N8QijFfMs
OX5ulTZD6zZDW+RtwlDPdBzXq5W+HuyZsgHaG2lRHRlGZkKZt1c1wqoahti5HWBev306obpOtSpm
AaamTDLZJ5zAU1vb0lMRjXkS6scTbZOdSdvh9wgGmTuUohqtU82xIN9bdy9CT3KFEDHK0vf0c7UE
MijvSirix3tclZZMkYApgg44Vb3SH9Y1hOJ51EQrS7f0rhkX0Mzl751hWdVZvZqqCyCL5hlRPsT8
h39WZ6b/nbiXAeC3QujGaBbW8jWurVG9VufTCB6qTWEaoMbkzvllTN73VNeR80ac44mS2/lCuq0s
fBg1cwJhRrsW+taENjK0FDeALxD5MrJDW0Z2M4ok8shWy0FRHq0XWNy/uKN3n8VZ2FdeD8l1ROLQ
WDHJrf3D0jZpvO3AI0YljDqrPOQP/964R8Y1ncgEbXljblIW/gnUlfiOl4HPpfVg5Mg6WR1ypi91
InTCvBw4W8SCVYaAbru1SugNbpXFTtKAvWf/ybd0Fu3phJmQ11iEimsHP0Drb7KvtxyZxsmiqRHf
geNKLJDaao+Zeb16aKBMhRPpp8YJOIVX0DSLBh2LQzbaXIVunW2wzR95+tTovsP36m5KLQxPKZz/
uP1G8Sjsnyng1Y4sI/CELc77WawgMvQ7/6mKpt9qJKZIyOEzUERGr9sls9fgqQFKSl3H6Bo8ZxSB
EEEM7UbfSqq3vzPJV9Te+1UkOVqkhHmxeVVdwAvRTD+/HcmmF8b+QUlRCTRiL/E6mZ8G5LrXIBZe
iGO0qA7U3B4ImGOaz595SHK8NUBq10l8nbCCsN97oncc2jyErZ1rce1JPJek8WaRdNC1U2x3+dGk
AT3/+blJvobD1WIeNpglZm8Vlo/xTmS4SaOixxDmOXp5dqEhEjpCAILDRP7zrrH3C0O4lGlzk5nD
R7KJNW80CNfmEdArz/9afpBug0lRSawcj9d5pm3Vch+xKu96aN0B3duTMCY6UGv4VCUxCN9nrx+M
+wkCT8zMLOhFAZOIXhHFfQtshAOCjj21mUWSYWzJI483Ss6kJVQKfBYSZ2vKq0b7If5bCa8MUA1b
8YmLcNu/yfJTF2jOvB5PakpQrtu3O2UOORyBK2l1Rrib2dOWn0RTChizGrApWWZTIm68sS+4GsdS
e9NvW/PELc1drIr8HYDRticU/OrBYYbrZWz0ipml4G3k/Z+IWnYL4WbC4W18LAtBV2xw0lAcMIDu
wq3SzgZR7gvdksBEwI0ysxfyX4GNqCmZr+TaXt1clqbhavLbzF9r4o8R6cp8J3ND3jEUjW8oedmZ
q8ihVt2cw7Kw9Zs+EliqfHdYQwBeN+UaMXsYvYthlz4sJHJKYlHJNqyTbaEIYhng1IJxVxfDCQIs
w8J8vmWPS9myhzIyXbK7NWYQciEfGuxtErQeGzNSK0Sy9KjSNXn/DN9g0/FLI8fb/60CXwa/pv3X
wV7jsHGTsCD926EnV7X+iNO/dwrE/7YvofHt6LH9X0swU+K0KIzFz6NoYQz9T7Bm6e/6Xcge4l9o
eDoos5OogeTfcxi9p3wNyNMvmlLTaSkNoxf5ylWVy9TQXfTUr/UzHi0u/p7GQkNNsVyp/yIGl1BG
4G7zxaVjony2vK1CCK7PUYiMTbu891B66mqh0SCUrbd0ANmAR+iuSYfEcxaZTGvSmo3LHYWpUNku
Ne45M6WmKxWdspfQ+M6tntvFuLyHpMy/2v5OvG7Dya+EJDr/F/jWhPFKI911s7Qk/X2VIIAua7TK
Ola0uhdoDtJySfwtuT9UIksL1NHEYhAwGxCSjkT1XP39oH0279/o/PPAFGI/z15kVEaulTO/qUG5
1fQHW9kWtKt5kt3jZkhbmgGBEe45bWcpgGfIXMY9UASiiZqbaVuTryHEKC5BUzPF8OUr1oWP9Tzt
SOSBLo/dKYltlFqLapZ0YCGAG+O7fyFvGR/NXvEqx2MFvlO878u3BakddqZwsJAe4S2v6z6JMTMd
D9+pbNa7VaxhspJUjr+RWKQYjh089OzkesC+TSA8OTkpwp8kKjy5Bwto0k2dgpAg37g02S3jVar0
HRcscb+Rdq1JviwMy1u4Lb8nXnNgfePeYUiewgKALoghWWw2LaAvMUG+ljzMjEEloPXXhw03tOe2
Y0auMH+Kzv7LiffrHp8yCuRdUHach8Bkg8xcWP7f4jC2SNgfqtdmcxcbyvkCrCOEWCSUOU1WIGIV
LJpeeWi9jh8N/ocTxDcqeRgIFn7YVaDEhJMpmm9MWu35aG76uxKDsBRAd4gM6T9T+ag9+nPwRsQk
zRJG0Nh7hVcOUvcwylTVYDYsQa5pbl8ySL7UOKvV18ANxwWnq0rLtFVMUq/s3XP9EsraHGBpYcdg
EKn0zJwmSMiTyvGV1CmP7rKEkJGxW8ymNjoqxkFePRfYfblSW9SlNQOclu1nqFWdc7v38m86LhPa
T65oncPxWVk5AI5kDswCxb2c7mYcJh/GrZpFzdjWgCxhxBKbzlvI8rn7MfXehG9VylUF4gKa+TD3
gd6tgofb27y3XfKUfZ9nL7nUnGKF6EwMbukou1ynfj21nuABt7tfHdV/jcURcxcEjPZYQexLhLje
cZCnxmHPAtDbH+scOg7T0ZTwUgOPx1887q8Va89kTY5kF3NzN0NvsxbefCU8/upCJvoa9M+t2OXG
2T7s/kxey6fe0MQFktdvkBSSQA7OcK8KS+sLr0+QjCdgnxrJnkoNR7OYMGYhkbT5oBhEsFHQVAvj
lFWsRwt89M8WjXOQkbfwXM/+Jju2Ge8AAYeS00VUPxuplkzk2/6a4ilX+DgHKlg1IQvmKW+xjWrL
ViY8D+ZMmThwnFfA7eUImLpaH3D5NkLQhA2yoLlykj2W3LO8pW8W2JVjG+CO17DwrkER+IgM4KFG
Ha8Zm094m/vjkfLyEWrlK5OBkdc4sCrFIduC0WAuTqFMJoanrcqaSwcrlgbSbF6cNBo2uUVWBYgN
etYQe8PHhm95SSR6JcrcDA0OjVVCwZSTfK5hw+5UP4KxPTml42h8XGPaI03YTMjfnfuGVNqcE/mj
+uEBlQgK1FtrT8yy0Q1iBHetbZS1INU/rFDqUHKi4zbW/rpeB6eHWhbsitJuu9AdCYzs9gij96Vu
KYF2bXXGxIbja2c4BMkbrIIJ/2kyvsILcV6Syt71RyRCloUKZemcgef6OrjS6pmnZMZoRPSnzD9L
URdrbgcoWc+RX7acoyfw4yzUukqzHeTQrYbVi+WseGwFkAElU0ZJIAwA8M11v1s9J09Kpw4mLDJw
mtPXGn5fabsB4woDneOXVF+tKwlyi4nEXb/3mgnmqEtWWd+0rzOj9MALwwhTqM9kfiJjlfpSNPQc
m73fW9BhzgB7bV+4X7wXCqNi/CyQ7ecb+hayTBGDYIIbq2sB4nEbhM80vKs/7xgp0IJ+xwyfbZaC
VM+DR4788ajAvrcQTSzAzibY6qhT70odFP8q9UW+tL8ZkxWzz1SII3ucK5VkKxSZVocTcDOHpim/
d+mq1vQpGMINUtvcqn1bQjdHvLaYdvF0iR1o/cpSjELsqhLao3IfjFocWpGHdFrGQiuNfe60AahG
2vKNtlzfRbFk4lQkU0PLsmq29Zl01M+839lD/A6bdhCAT6E+/Tb5BaTiWDT/tI+wk7vv1CLRLu39
Cixfwnafis80Eh/vMg1bOky0xAh0Z8n0OroWgu4Zzd/LXyF09Wads7lNRmQZDxty56E+kaAAGbu1
FC2MbIeG+oN4YheluOReSbBulPSoejJgN/L4tnEsMIOim95MjkOJ8rpn5L7gjU763bcFVCLhm4mU
zF6ov2adEWvHenYQioLEonA7GTapUYWaZ7zPPvwjepOu0ON9zFWqwhRdDeRp3MpFcLhsilA05etJ
DZylqRJ2eBTYbpjJmNSbH0r1mSKrVUXdflXq0jESS05Qj2LKVG87HhET9oXGtxEZ4E8Bbc6OGYmv
OgbRD8W6s66J/Z+PmL+w57vgC2gGTrZkDzJ00YiQaJQMNTQsuRsy86ozpBguWQFwzDG5qZkq7L2W
rhSLrewp8jZtHR+NMFIn1DqNK6yYZwk38IvT8dJtmFHDbEU52xACdrMfjOPf0hDfXzwZJtGc2RFa
QDtRxkUOA2ZLtpEWLCyim/W7Z5tIVwpugaGaMk0I+/fMIdPssjqvGh00c5dtWYYHaWwk/66CK7FR
jTmlZhB68EuXMpXWLbR1ne8sQPWVXEuomPkpc3AGtpGL+u9BI6Hq0lhRlwpx1KJtqfi8I3gN7g6/
O7mmVHbCNyGEdLA/rukrMTFuZT1MenH5JWbXs6/YYLpXfh2+j5f6ZW/PxmevwRWhudXeGhE8fkmw
ME+TswG6VJYLmleUYgB+prdkzyWvfhZsNM94BC8q+JdaTp5KwDjwPgx+BndofiyZ/zrNb59ZXz94
tNgWkUTORrVUupQreaAW93VJ1n7PTPwaBEp5lxjkvcl3e4eDaVBwoaYZPrhQ+JFRdaKk5MTKJG2b
BxpLu4o9TH89Dh7nwB9D9ETJU9rFpeI401z3we37e5h5zR7phR5scdwPvkxL0x7OfskGDKzsW62Q
0XysdGlVGRBtS0ooVbZN0NRPN0eVegbaAvtrhd4qGv5n/zFM56lC1KwQijpWnWyaviGEJaeqi2th
eMG437KhWDJhs5aYHvCockWjzN/3SqsSoQiUUiOf1i8PngjcyGP6cWu4Bc+lT97dPKTSj5cUzHOl
uFNRNc97u8/lOaixRFwhgWafY8m5ntKhkC6h0DH/icVzP+hb1fjVR7hX8jaMO/7b2fPlDXv1x0Zg
d1ATHyvMRVrrtumADU/9XxtGzHv6VP/aiT7mK3/n+f0dR4KxIkDUf+ypHfKhRJ1r/repXFn8oIf2
nYlS8v4QGsP6vf5fV/16wuuc9OB21BS/wX8zxRkZHbsd5Fz4CqZYfBJLe5PgcPVadfeYdp7LzM1c
Mc3Fw/SNnzDfUArd4eWwODRNSEfDGrOqmUHjvFJe+aWnurDWKTuQpIpP/yg6BXS7PEgRWO2VEC/F
+emvKF42WYlw0t6g+gCGU2H1sjGxCwkwDyGsmy0DXb/TTdmiDuhx7eprtEPSnnfuCLC+9/fzQamF
tbAF9/V0bJvScu/SaX8kPO8T25EZ3FNBd2lyZj5ls2iKnDmKbi7iajGvLVxnVXJAd3u0TAc7kh+P
2Vx1jshXObYqkBn10a8NutlAOLJBkwKS1LqnDBNDac8fKchzm4Vfjlkf1DDb34LE5CJ/5Pd0lX8v
mE1PheUj5CHSn95zfdKQ4mUJ+QoM49FrTH2k6dj4DwHWuAWinoWG6raIITwHBUwySkVu5ieBrTNS
3+B23R5Pzyw2uRAoEe/s32rbVXY73SJU93ExNu1nypo6j5HhmVfxR8uOMDqxFilv00n6hfw5WkeN
UTzzCiNoaZ39sGc6g2xP+uv3oIhTyFymPirUo2RM9dnjIBG2gGESx8dse1tujYfsiWIPnBq67hnE
h2fbhT/iUEdAW73G/mk+7Wv9NfGNx4PspqOHpgwCLA0G6rxpvm5pZXEgUaYw9OUsh+goF0dqUfof
VUsHSHof8yz0QrG3VXn/mzWzo6cewIFHuVrMIWcBMdv3R6yXIzCkuM9kRDgHSEjcvrR1rntyeZez
L/Si+pfWA960DZ7cvshufWMLQ01CD/TEet996+iY0MnYS7qKAug9qOjarOMpPvJPiJoQZHFYr7Lj
HmmpWbwJKy61UEoSwHxp8e5QLm1D/35N8uC9A/K0R5MssL2zjoicjGIiyJD3+BCaA4dMhlZ9yc8t
UsVssUJQFZmK4y4JgQ+0uWTgzifNjaHHWVQZ4+Ky+tb5saQKsg3u+dvmExOmo349sa2GXhyvca6B
lA==
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WiwaPPbP690v2k8HaZcFMQliXY6pkeAfCs+r/QMQapR1pb3R5P4tVaK9ZdCYfgg/3d8PFQOpuHGm
1dPiqOhQMh08kE/y4wBeLcxDdvtt8hHA14xL0036NWeaKl6f0qO43B4snMe7BA9bbiquMKxtrQz1
5TKqWg5I8f+VXgGjfYHEtl+53N3Aj2dWJM0zxeYqieI6rV+lcrZiZS7Oon85B26Tp5JCzK6TdBKv
lzB5NLrgt6EDR8Ds+DlHPybLgBNpnqNekFHXK/oUC+6jepFYVEP0caggxx2z+s5BXiyTCg/ncTBq
jd9R5f4nYHh3ueNxMtcEgjIoetW0Q/TxdBNklA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 124960)
`protect data_block
qsU/RQDlCD9+S6XyPJeGZaX2wt6+k1G4J5lNqIf/pa4pr/Ia4GXIyz5y8CNvFNCba4+TuRFtyyv0
l9WiQHXNDgN9Rg0ElxGQ7rBrwyJ21hAAJELdZS1Q7H2ItzOIrkfCxQ/fhKBGpkmALRdWIODBCLOu
S5LUeMxFHMGvzI83yuZREWV/ANd8x4dzp+jXnq/pLqMd86e1nXwVDwOzTDh3XY7PXE4yZn8lNbgf
x0SAoRLb8vedMhxOkFYBV8iY5c3BG+Pi57j8TSVu7YhOkRiUpCsspjWlNLv7rQQz5KYBHvXT0yBq
rTDhV6jRJUuvrOV/Ul9V0nbiimtaf6W3Ez0JRMsITicQWkQ+iLV/yyvlbiqYkNa9dCxjSPbksn9E
SsZreaCE+iIGYim47fOKy2MkZcTtpXimnDylBhc4R3JgQtotGHM7WMGXnnlLb9QORUzGrbOTmU7F
D3/cm6guks0AUC3RPdA8nZinHIiqp4qZSQfj5DEHYVZc/xMDgMZjHbxp1BiU0lFcMGt9vzOk2m8t
RtQ4qZASugIaW1YIIok9v2ZVpaXuDExGNHuDIgvtLVH44RvhUCS4Za1b9Egl6RUlfRVxAceHc7UH
SsEKLKPJWUMIX/Ec5Y4nfI2K9XAJmmwYgjfRp2yvjcEee1tho5lOt1x2k9udlzkba10eUTqF150q
EtW99XLNe/kw+sPJaMUHtnM87wQG0dp8xsXD4KBZ5LtJDzHnYq+TLmmrkiuML6pHX44lwct9ez9g
1l5upE3yzGDqMo1FPJLC4EilAT563C1KR/PDQQ3otpX/HDRTzmNZdrJrjfzG/TeXrQP4WlCNG9aC
P+0xOu6eRPstpSdL6A5U7TsoIdpgVoorPOPvEs4fQAJok7LfYezhrHjxTbSZ7GMlnRO3v378Y2QV
CneVBsrij2S1fjLsipyitspmyDdRmVUcEihYsCE6I5Uepifyz/GU1TinzdrtC1cRt6YTW7hDaRZK
ZcJYzx+xfoNUEgIkkwEZZJrKr9KK9+SfXMxP8Lh73M8mse2dB2ZcLj94RlDTFO40IKqpxxnrXM/F
oBGIbdvU8JmSlLyhvrD5ZqARxaSqXLMgVDqOZeE8IX/xqZCi4GvBMYgntaf1LrSRFkRRlmr5FVyA
drI3UA7JrNHZV9gI+tgW7W6zjWOlUvdE94h9tSwtzGsWlols1MbsbgWxDTplfipzL4sn2IrkJbzR
HXCyYcxUsKS2EzKoABL4rRRFtG72w/XPLgLw/dHU400UPrvgfZZr/5FrXwfnoWuo9w4viojiyRYw
21shfEIvQZQphUeisrdddA4xFNmzTde2f7H8ajRnzuuJA2/q79fwcKbMxZUKSlIOVrnFrG7GCdkY
h0zs7YcFM/5FuOvMBxiGtzVawapmPDnIJBgUWijrwKnnm25SKDBSkccWnVj2ui5tXW3fEKK9dak5
+EUDHnSvBbfORAIyQN39JNCGOx5CZaElv0YMw8wKmRQWhPdWEUmRc4PD63srAivwZV5rAfXw4l4z
ucQYIruO5ep4Ri3LNIuJEaKUCjB8gG9gtxwAv1pY+PNlL1lU7TnBoxBRxv+v8rWT8F/lfuSb/9Ap
LYKU9WwLs0dS+H8mAnGy4/b6smu7cZRsu08e+ldpPQyZoimnVpOODObeN0zvZYvo1ApC4PTDUwAE
Exw2U5etsLfA9jG8Hce6dz56Mua51q0Cp8RnCGsHNdsMoNEFzNAT7HJTZ517/aeSEAYaMegwppwt
kNhfoYIFfA6bNGS/aB0Zk5PcI/IBfEAQMoHk5V7+BetgCBr0R+8wqX1dC5udjJJz6ls+GAG5U8Uq
omWTqGjP0vzo4HiCZ5HUt2VBC8PkKHnr+nUiORsJI8zksaNgdPYtFDAZyrFhGINbay/kuIqMheYs
ax1/TDgl2vIUXbcfFECu23/bL+Ut0YQzf0djlk+qc383Wtjj0r3Z9zPBumjCN2f2B1aZqnoaGqiF
b1b8kQW44bTNwLjXm5VeWV9bxYFitwMRYG6gvh94i8qSTdLKcycTvR9DevyZwqxNhFINpLJtoEum
nN8nmYysFYP/Pl10/VhzGSoa+ADe66vLf5yCUaj30hSaIpGiFOpbPSp63N+4k1UWUVFohG034S4v
vzq6ex7wc6w5O34fhxp2XERYLdw2h2yq0DPS8KywwjOJCbGaBED+dwWCGRacw+VBYM5pbtbP2VJ0
PoY8L0WlZArP30QaZVpDzjAr1rrL4IxIyRZdXf5dKAvkPM1fx0DBAVyk/ELLBHakb6ZGjZtgvV0D
9tJ0++nDnbw6DxrNhBlMSP5wyw0ZDRXM9E1B4GHbM8HsjzsVGoM0MYTbPSiLzDiWzIWWiRmF6FIw
blxHbLxrGr8I+LSs0Ka3jTbn6QhbmsH70UPcaDdB/DptcxqJG8j3AF0QuJiW2hTcQJXghLH4AmxV
s6mu2tkrjs3sbmjSpPHDWMDzdStZVpAPi6ctU5iBfL+B8gB3emo+aKQHAKpJWFSSQYGjgW2oRmFZ
e8PobeTouWFLJeOXWi3ynhTLnU057vai7kL0S2tC4rdJE9P8EWrPk4CDu4HBuTE+6RwLLdr7mupE
jfs8OeCphy+K0ryRkB6XGcwZwtibP6i0fJHlDE9onEakPk0n0eMTgQLI5wjeVXauymlD7ABaeMfu
CGOYZUVoz1+lVD6RRh1Bqlp80yCikSqL2QCXaBAYfzEfihKuOD/Xd3zJHBcuUng4X/o3SlfA20lz
KI3CB2ogpEseb9n45Pzk6Lzm+QEj5PrN6XryvvoOxAPUETDG5a0x4mth9sLtM9/kJNb0Njc58L+M
/3owmrd3MdfgeWNhaxjdT4TFmO/+S2CI4nI9GhjrxDCXpwk7Ce218M8n/B4CcruRPW5MXw2L6dZy
5Y7VFeEDWz4lKuTMJm6cMeRO8Mt+RVyowaZTezVUODivIjMsqj/CA0mcRkNhdHE8XtFsPA/nUTNP
2O8KpeBettWDIRcSVQQDpL4pbOjMNITVSaCJRvZ9ZMv+3T4S8RiGDRxXQqA5j6p4WQMZ9xWVfpqN
9ve46BO+aFbz1kfgsYqyqY7TAdKBfPafv4dIYil5sHwBG2+/VcQ32WdXASiOI8A+2ffabwKREykc
W7hohdKWpqpVr7v4AxuPx8e3re+rAqs+zvmfd6drxtT3HyIc88WmTtD8V7t5sPMUt3l5AdyW9M35
PnYz4IqQvm68t52ekJZOw8aZ8B8U3FLh353l7Q/o777x0o6/Z+mPyNUw36kbYCirO7Hgh5keLiWP
sNMqMwOfCiVw0pOBqiQFQsPaqLc8f2rz491M1GUawiOk2eHi5ZniH5TC6PZOMOXTd7Ds9eO+H1nh
L5+ZmfRAFy4ocq3h+Ilj8LZjLNMChjjLCzOMjk1rRB3RKiRZfmBI/3MfnfcYus1lHlJk+pwHBZrp
/weoIiP8nrXUVqU+9WTe0g90hN/rrz1OcuGmjjc8SGkby23F07d4qC02gtmErSyXiedMPOpBb5Q+
uaIHTB5hz7yl2OZAB2uZsld2glQxBA+lXaoUM8HahWjmJppMQhrG+7qcU5fYg5ZRXG4vohIYjh+U
rIz7dwE5U//YhczZRpcl82d11PRpENulHxR/6Qcvz/F1uh8lyzQuyp++CezTIEcDkeS0UDbH3NRF
ODsfkQtlv0KOZIbWeFR/dgblzRz0iKXws/PShJrfMH9fbVdBOsK+pcGudbpbH0Qg4ODBcxQXq0Z7
V5XyH2l3Yij5JqYGYt7NgAA+H/sUgZKnVI3Qz3gmC2x9QWLcN2VtNCtGztnOYzC/7rZMM4VrwIgR
iJMN9JW2ZSwv2NzdHHKd31f0NZ6U8aRBsZ3r5wIU1Wp2fwj3Cy4WGK3rDGBoezdJMI+GuNBnYVcS
NgnFAxyVUhjdBe4RLV5CddJ5LNmRSPE1y/Dlov6AE3VTa1WpL8BxWTVWfdHaPT6gyk13Z2cW342U
AcCIDaNyoqr1vyR5Ke2f/12NvwExX/UlAsLZ/wgBFhAsT1Lip1TyJVCE5todldY83EKUuu3EXwHC
lcmMcmBH4CWbeIME6e+14czZz5bAL0LmIqKKmYuUFMgzXTtRjhYEFQ+4e2P4bEfqLIIuF+RaID4m
2/XOkt4Sww5/2c5g535ny3EOld7CNxjlCXp0W6nNeFn0Q1+t7AdKNH5zDd8F8wCd69IFuIsqoxBf
GNEEZRg4tY7r8brSvR8J/NM+vRAGo/AMNfLHR7MKBlbVsiHn2NgNjuRl+H5nOEglId8pWZpfbtRr
GD55UXWgDxfjycXS5raWH2FmYnr7XxkE12faGPFN9ZITNzW227qhkw2aOChucoOqtMgye2gqLORf
2a+J//FepZeAoEJxg0lLMJH/oOK6JGYpA7PBG+JzHBWHOUOeeX1uxbMLqsNBJyVgfa/dqfnc4O/R
BGP9ONVxADyGhqq/rOqXP6tx+ghWVcadUuXziYF/KMTtjVgxqNyRQqPRnRSdEwN6Dx3I/YwEv1W4
iBGENR18WKPMJTPBvDXTlxQcqHuCpdA0uhfynfiWe3M0JID0J4oJxCQGvntLEZ0/fif4fYJDqpg+
7xvaWSPEAqkFWfPDRRuy+Iuipj+CKXvYvJ+5FyCHZGsfdFAbCiRE/vYnJ2stIaVIJ3/GyulkCsNq
Lh97MkVZ+xF2yEgNPEIfFYDuvZwvGERWN9jPMeXXzVPESxuYvm65ZfJuGJX32HvVecXPNXqYo4Be
JDmGPFP1WuHU+lhbp8/aHsWmOdciNSb546ZqwJuKwoBeDJ7gCBpJQycHBJEqDSlVwoCL2zDKbk9J
o9y1tlJNwBwerFq2AzTho8IEWYZOxW7Y7jp08HZgE2UhxAYEFSwZNX9zXhzrAYYrro7WWz2HyqBX
wX8jfneevRoDdsEqi8DKDzOfeBubdPkFsPbuzkJJYWMJSj9gWxL78bDIpFMBEk1mF40ykNwHSWxG
vXR9C5XC59AeljZtMzBKRR4jWq0s89AX6GRQ8vdFNh6fF0fIJPCOjjQsPHqOGz3Wa8RB5Z7S3tWt
uBwBMw9Eqra+jJeJh2Fw7NEs2wsjE9+U9DpxZqeSPN04CipNOVXUSvsVrbYwu3CTLm0RGZTGc+iV
vCfhFd8M9GgKzF2PR8ZkkmFu7FfDQLk9xmDNa9JRiT1SqUyDywqiWoybmxMI4usHuaaVR8n7B5k2
TvrCPyICiHEiVNTKUCeAAyhK2osTjJ01AX68w6+Ys/f9pJWocjoi0oDPU1X0BaY7ExIvXrQJeB7R
LSVT1iFR8AFl5XvsRjrUoR/RSE8qTcrxgab1N1iqVtz7TozV8SlgFQJ1hVlKikXLKQ6Ec0m3tgPx
1FCC1ZQMpWmKV7nqX46AvgsPBzioSeF4VQcAXnJ59LMUDt6589AwFdotepY4LdvTwgMiTNg8N/L3
YfHTHhrlYt9j8AJBLMdE1yTR0yn3mr4PEcdTyDGBmuJAq6mivxCzbMr90aIPvqYmzSwSw/F2ixJA
he+c1s1Ii4MPiT9DhQPHbilfdJI1wToHfha12xb1FBqebwHRblFXcTiwr7d7NCDd1OKjsoCotv/9
8eOVWBJOFPrimWJHgK6i31EDC8o7bslPEsZzaA+rUsbjFKxc208boD1LQoXn3SuHnU/PddKiQzAk
dVN1WhvP0xjqGTjx/WVO2Cv8nrvpuw36SyzLUMOaYQB90juIbdtXZRNCk5Nbg3WimQna/CSW4bvY
ZGwjcJJRSad50Jp5IJPVnsv1PjGZrk+T/4sCewi6SPVPJGP7Eu7rlsd5obh8sZ0POSAiVZKo+/Qz
Y8XX0IZukY1ajfrhfGFfz3+zXThjG1SYlGyBrdAtR9KnNa+TWBM4FQaBizYPFBN1XsLkRaogmTES
iBDjyT2Yr7ad2g6QS1g+LjRZA6fj/m5/qIOp1UppUjwtEJ7cfikSxZzdUMVQBfBWmehDxXl3XKoi
caQOfqm4l4h2jV+IqkSUjaciXCrjMbAdTBI1TJKzmrtIkt4aEPwfenbr0Y9RW0Sb9t/mAfSJQh4z
NnERVr7QPx5h6GNAFpSiZthfuZhETFRQrQemo14LIaFfxrhKEEPBGKSEW1czjPJal2faWUH4GRx0
L5yRZubo45lctKoCEiY12lZk2KTPlPs0tzmbWMm2zfNCK9XfDvkW3667h1xY19F1FackMgLA0J/W
6ltV486Klthd2kN4jtmUTDEMohqw4g+ybPw0QscMrBczoUVp+vNFa8sVCRmeJSA9jdGoYDVK5QCG
TRuag5zY9UfIrqsPiQWxkSWe9dVgIwOnsktKyuGY6Sia098pvYnQdDK97S7cuBlBYNhcIYRdZZZQ
yU/4kxDS+KWkLDECx6HnUUowlyhER7uSmn3yQWnPfHv8SJxkoRzcqCLAF7P5urvQNrGNhrqBOKr7
ZDQtx8LtJqOHM2TKU6ISwODl22vx5q+iNszz6MHcpc51EimBDp/i8z3NEL4Yu9WNrh+fhDVALjb/
dJiNWntqXRcTzOxv5swWPnUCxkEp37KZkRsG06l1R5uEaamaSdXMyUY+WC9WKlKA1g9VW+j9aHn2
0iX0y/hsqpzcrcZ9YrNKyRgnSY8ea4mNCxMv8sKFMNAjYpg16/ZxjNLk5i2E2bNXlER411j2V1oX
e9maQhn1W+VJnDoonD+xqZsZ9dRr566QclpWsWqYvompa+ri67p5RzBoX7ZJDMGZ0bxM+lngwFo5
/QGZ6rdBlGY8ovam0rk6JbclkoXbr/Ou7nDa+HphE7BDWpAnr+RKwOYeTVHR1O9UMK9I7Tpcd47F
SbvxKGcb3DUGi9OQ7NRmEaP2TZ9yk6BABSaWx6+R70YH8WK88rZRZTgShsfbSBAGb3ms1cvX0HWc
G4xIjzxQ0kB56LmgA1fHCJta3YHqvd8XP7xR6VEf7kLTf8xiLnVJK9bXRjOv7T0j4INWnwRMZqpN
SCK/yHQP+DzlZAinkwNXiSKldaQ/xKH/ZHq8FFDzvjK637T/ue6DpmbJqZLWvJ6w9WDMUtGd42vt
t31UGjVpqA2C9H8gbgWgkp20pe4bJqP5+61JBFWpmHr7buCo6Z80qgWbhp6YRel6DkdiU14qwOG3
gkIKJpM/s0XXgkufvZh3zPovOxcFDKAaF8ou/mFV9BTRYVxF2S3SJFr++BsfyBHi9wtN3XeUukFo
Bt3JN7zO45qakCEAJYnS407DtIQoswyUg6c8tqgm6gbphcjOQZ6jpx4x3IoD5eNhAPmBLl1yIuie
S43oucj8+05IeE8380z7ek4z7LMo6+X92BcQS4o0f6oCnOPi8URIZqzp9PsoPgBd62ACFRgzZd/s
6vPSjQrBrY4Hl2oNkDapOimzA1TjLPcAxbVM6QDVuaZY+HpNjQ88Y8UBM6J2PMRnZcLzkllqftgI
eVTJ99JupffelNpxAULG1mFayhtTFNsrA+5B6w7dlYmeXF1MqBSTZaRMhtekG+BbgbGmLdRBJ7/W
/QSKengN1ziZXHTn+mxBtiWixvOcldh/RVtsgexET7ynYJuXvX+IIA6F0e0m0Vey4BOM7gNUbxMq
f0CAmT46guljoF5+W5YOemuELCHuze5mrm3pQE498oo1YEH+fJ5of1YtX/M9vhCl/jpp/cXKqb1g
RC1BxHDZ5cy/ODRzwq+qQEf6jw6N2bAmxSVgJ8XBcxvadyIMFPP7Gy1wwOVFrY/gdRvpAWIJ8lcB
MaahFN6kuWiiQJa5J1+c5pBPb9XpnRSOovJ6OHHujVH1hDMndGS2DOSpyG7zU+SzhhQ4RsbwVuXs
Rr3/Jt+n+lXF27E22SGetKjUXCaWIAeWOX6UabwGWlyOT8OioA2hlSbBMVAEA5ncozDMSMFErKPg
k4i7sdjCjy5/my5QkyngcRCVvvYxeYrW2ybdMDExi8H0mhBmfMafYQlAi1d+s4c6tS6HbQIgzB9v
aJQgxVGPravB3LmBfPjmhsfN/UfZCKqw2FhDpHnHTOFYnWONAZncdq+7QwYShSkONeoNYcA3eJ3c
96DtctqEGaRKSyRHtVjv0D+weS42Sh3KN+ESTRkUE+2cD6NWSOgMGV22Ccez9OThkPY7rb63JtKe
hfMHqkojT6EwGpvSbTRmKm8Gexp6LVJdQkjyWZmfRrK2BFmFKGgZYLdz1HoImkyUX3wgIO23pv1V
4lFDzJMCru7TLGJqGbzd8TTV4fmOmaRueecrLnTBpTkBA+TwWWdDunbDvZAmzu2jgG77lAnhIC81
DTQOF+jqnxwedJypZwen2n3p1jbmcRdxWyhmj2NrZM9CBFNFmyR/mctq3hapPX/9Mg0vrOfeOxC3
e4pmWuBVhg35kRzAf9WIaFvHItLjU8bAoSI8shRcYl+ybyO5Y3VA52zo8lDdimzySWDJl8Cw6Smt
2Z/A3x7mWZFKHhsz0PvEsZ62ejdJLpZEq8JGmIyIKR2p1K8F6uOFhxNAvIHTIP07TpuioO7Xpvs8
2X6cvF0ddyq/1Jm57bt+Ftet5woBRPFsIlCg7C/khuVRA5aO1wxt8M6kwIfhfH3osfBPiRo2qcHj
a1mWwa9Q7LK/CveaUNKJfEIzYdb7fSumxAVhA/+De2wXZIhgftddD09SLeEC3PiHF5+z9yOb3agS
HXu5a0rppkLT8fd6VT2XXNzPbMJIQkoZqpfg5xgZ0spKkqA0WgY19707x7X9gm8C6D49D2056p7D
Yv29a6rrmRBp34iuzQ3riOfDsWroUS26AzPZS+FnELoOcK44NdkDnKvQTqzvLJaA2XF5wOKU/aM7
A6cXn2Eow9EjO4DaGPZMyAMiknpKSSVZo4ERpmZcEH/zzmOurc4YYO+eYfS/EV9miI2hv2M3Z2eE
fD1rVhwY+L278JESusuKPAXmbSBDonqHVnmOs0HOF3ac9tJEiaXLW/pUbyEKl4Eo5Upt0pFMTkR9
doQisECUKlT4gknUvuBkq4lpFk9PZbEvXkMpJS8pnvRVR8AvDQ7FA+Wuj1cwd//RD9dgAXu+WMTb
rc96uM9yJ8O5nFODt5a7K/9zbosQDlMC3R6wiyi8krwf7A79KPw+loNRyktscrnNk5h/IU6u2MZw
5qkwge6AKFVNag4gkTMq/kADPb8RVtd92flNPBBzRu2fRZaJj+57C91QNpy0AzPM1Dit/xb3dr9M
twyaV39w2MULTABAuLSbOSxwV1q0fXGOHgysK04yYCAMH6n077txBT4B6ut86hek4oMUNA7zbYMG
UNaDZ3rYrk75FU5iJ0sbS4Ju0JXrRXEVWOx4kDDYqXP2hOOLcL9+ZjGFOO8gOlVEdtTDBp/Uxb2S
A+fqD3fnGBAdpdRrigYZJ0AOQV+D/JyS0e6Hm9rBJZCVQ4I21cpA8IzlPs5k9UuQOoTTIKnU1EI/
d7ntfSwZcouYRkfE9q3YxcsGhHPhayGZRBkMwn6mDQ9yUNtVBrYzbW6YaFn2bfhxdsQOY9mdLYq6
aTAZy6CmyYroRtUGJEMzrGBMcmnKyOSpbO+qjAy5VUGgLk+vK8UrboW48bsbSC1o7WpgDXppwRkO
KQQrBxudT/ChwvxW/+RyfT8EBuv2QQNcrqXR2XEInLRGDAuXPkmr9PsxfPiXVJGve7tmNAOFwKuq
SiJNUKbmDjSlU+H3PoxsdZEZ7r27tmPcc0CUjddQEoKpbDer9pIUDM/8bScpArbp86oXSK5X8mjL
/iuImOoynrbzj0TLnE3dby53VR/dVfFz+v9KuQzeXEVW2IfPA7BU3g/3AZ9yJN0DKXBhIoK2IIa6
0qAl0pzQvRfiBz/KO/UFmEKBV5JncLRVgqFATDYAF13SKKPZMTpvR3DB+fK0BYx+DEFsvhvM7O1X
LNwWa7XmsN3RlU05XoT3SThWFHZrqLuvP5rCrjBaQhSv6eTJo71LyP6b23gTEw+IxdG7wnAU2Ro2
qABpScP1mB98FHX6ZR0vCIcpIgUaKi561DkQtDoRTqdlyy72fqYSzg+7Z3P4ZH0/2l4XL3V6nFsb
wtv436O+AG+k6zLh/PAO/f/+J7PpvgCAE+3E8Sp5exvZy1ebfi7vDhJp/GMvnlRxXv7LaOifC6Dg
ASaPWK3arXz9Eo+6k/PwenYsuzJChIeeLTwiHJBeKX+bEArWeZzxmjjBZedctHmNg3hBipBKivy1
mvsBZBUa2rxJCMSx/ycBK890WP7WXYEQU+ZEO3uZXR5o/XXIMc9/Q+6hiOefG85hHl0H5stxjuai
5nepeqI+Qxm+KjGRu7QRc7X679eLvvdBCOVjSdcPRobaE5QDn4RkYXyTA/ndkFfvFRGLF73a5ohI
hG6ey9gQceoIsFo35Sv7t+GA2Ktbuc9Z+Is6VPXUisrPzCNylhQpVeCS7zVR1qrrHYrA/1pcRi7R
8OD92RqyoLG0cXd24AiEznoCSZIMze+kqW5207kDbHU0eljPsY29DkOSdsFS4i9h3yde/Znh9lGv
HHQRLej1MHxwrmvskCDiFWq9/dSxKf9mH0yBXnIYoVIW6oRFI6rbBk3VZh6e4DP26ZM+R5C5fnpz
DkhT9b+vE1T3D/vR5o5uALhxsG12Ah367CBpUjTVbFMTK50nQ9ucHcq7ScMi8uLh92O8iG1j4Vg3
/eA4zuQDMyOAKkYYqDrHk030vzw53hGzEAERvxwXvdM1Wx7xBIrex5w+ho6jmTA7kfDaq9Ck8dTi
Mz0Dmc2NHVZRizqVY5M4DYZcm4PVZsU1S+5LIxL3+IFs8rA6Z9Uxkq7Ao9c5bbP6URgcUpdpwkx5
XosY0VxhsLm+S7nbSaW/hvVF5EzbP5RNHL1s2j9gG8iZhY1CDTgtD7DIGIjx+lSN0/bhIv5PYvNv
H5uvfiwuzWZHgyzw3aupT88BsB27iMoYwym42HYsGKEH99xCaxcR5zq4aSW95ZxR3UZtT4DjeGwI
GoQHQ31iGW3CtCyS8/kx/RcO2+yeGLlNl1121MXmwg8I7tfZODcmWxd036b9nyiqeszevcnxJjQH
5LjVivivREO10TpI+OJxf0qsGpsO+yVCn3C1b8jCVk2+h8MPFQULbc4h7YWRDpxLCelFdrgT+ZGW
MGlllGOzWYbPrGKpdX1DZc0HUzUZ6VJVFIB4Mc1ROQ6t3A1Bm7Fu6My07PEqsD6KSYW35PuopQ6y
QNcaPDSSboWgxlzWiZ5X+9y/mfxcbm2Om4XLRuADXxraZv8j/Tpe8sMbZyo7G5GvooBgjzWiWaSQ
GWkWZmtZPEJhpAuKOqiN5yojY5Bzrdpa2I8+15RfMm8+W1Uy6f9oiy03vMcHQRe3wDfrfdAkkdim
v4f1h0o1kulSgCaUKMqsKmjjHJUBoQCEJLWd0mQSokA3wm1m8tLrTfn9oRdWCUPlq6vkZUCplJsi
S9GNUZtH9U4uCjrHsmcktGVclcMWh5Sb8qOjBoZe/02jzby89oSZX964RX9OdOgLAQ5croK3wiBH
4DpI6Q6Dt6e5rXPkJ73i2n9gL9walRJlneZ5KBdjCDmjqZt1BqcDm7BXWW/Iq7COK43Pi45Y1g7n
GivZf57qiOXdeBTbiF9WK4GtLP9tXU8MYFvSAbkJT4Lv6TxCXOOFBryySZKaWQDgZ8G/jEbANPTt
UOyCbxq0hC0LrVQrR2uySIkgWRnQbJn9Tu53VJFCQGtHuxT4n2QEiOmF7OqgfKrFRfqSX1hbibnr
6QTW1nhwjMbm6qcUyGV4uyjuL73LZKLKsKfYEJ1GpXCuPZ6cxEkGJL6lZ5JVc/tiBRzUxkQ/6KOX
VRgo4Z4gQwZeruufMsGiw1EWUg75FpZbXOBDReD2K+MiIUyT35fvynbTBaUvh5OsFFGGSY0hTA6c
TV1j3fOEjikyRFZ24onRXve8BF4Jnt0gUm5Chh7+c2W/5r9yjbJEeYZ0zfLjbY+uz+RUqeoaAbUf
WsYhYwe7Zt9ZqEVRQ4SGLX1fMNs7hhWrth48ipvRZIzddOMyUkpE3a+SVUk+YgJlJi8fPUsuukvp
RgYSCCkNqRDFE9Dgoka6e0eKn6o3+cyAJodtjkVjHXeakJqqXmN1GrhfLY2ADULEBiFuboA3Pt4S
9ldj02G9hqwGioo9h5xvNTRosy49f9yCe0IsM3IK7p39ZymZdHDBZq8zUwSwHPz9hYo+2QTLkbgK
IGz4GAyJDg2tEdDOaV2LakSqlRHiQHm+VVaqodOKbZnV9331Tz+dc5TgOxt681m6VdnO3zT5eZgH
WRBSJTrXGfxGoagHeKdjZXz5+4jOQAOcfIaCUOqzVpyDpnvc/G9u5BjoTpdcF5fKHQF0rXkzhFZV
QVfd+2NrdieFB2blV0BSL6nboXgEaUeN+BdnRTyjnedE+019oS855SM/cf0KTRQwU6+cC6gM7c42
RMoCRqLYLIxTDmfuvBWFQyYf7B9zAImzbxqjEEPG01WFESPRYhNcseMadmtfziv/yGj68Q3t+m7B
Ryn1gcDNZp5bsEHrlECXlMGApwYpsnNDXYyauJbIUWrLNq1ELbgBrhE5DxNDoaToxVAJv/FgKftT
ls4oyGQ7BsbegYrQYhsxl+m5t8DPywYg5cxfLytKMNsAZDzcJpoG5NER4xU8up1eaak2CsIO4P4q
chZFQCHThWIVq7e9hbDi/Y/9MDax3lhnZUmcCSRUxCVF23l21YUMYQbqxwYG9ZvEsjWw6oaNCWFe
PwQtzebUTBGxHfKVb5MjKt/0vSD12BculXkNxkzprGqwC6tBRSYaK/XIj48+XksEdvpam3kX5ZGv
/cYE533/y8GW6/BGoTSGh9g/zejuOan0RTyC5AIBKnw9/k5YcU0PEC2ZC+4NhuNkee9iOayhQvB0
ZzKgs5RnPs4VzpRUERYwnok0mxqU10Ju3Q1JSYOssxVLKkso0Xeh3tMMauNHHl5q8/DGk31FFWLK
qtKsN7oWOCPHXtkvSuwRxhvUpqfncct+/NnKLHtsOwxvFgWEnlj3JAtf7+Po4xScoW0A7sIObzd0
5A+2buLTby2Di1IFS/HImIAs2zDT+DAWIXFnaCBfc3BHJGti/3Ce4o8ecHc7tTX908BRIkgjTc/g
GuYZRXmJ+SBiBwkGHoX3fBCK8hUvC3q3piezY2vcJ2XdDWYHCf57iVh78MoReqbccPQnjULUTiKc
DR6sbhZlyWnnYPkmDDxjw0Mhm8M6+j3IZYyMakPf9xHazn+slciM/CpMTxd/sEkgOeXpYoYQsh33
/f2DqYSuBEhtwoj0DvCj/6AHswdIEmQCmpDCopAX2MUjCZHRAye6wdp1NQekOxYFmvCZSR7ovani
qR2Toql7C6QXAOkaGx/oUbVtgK4SKyAf5KnwyL/AkcnHHWhF1F2YjsDm6lRzTBbpyt1F28vjG4y2
fQcMiqne7wkY77qjrddyWt9cPYBO06G1pbPMP7O1t5Jo+Rs0NJ1Cp7VELKXRcPOzkWxJHFJF94kA
hoc7ZbUQJW29ZjU40i0/ykcgvMONJA1N2PyfbVrADcBLTHCLYBU4+1NA2A3b9gbisAicUE+dIOt2
XJW99QZJdvupnvpR9PKhMCihjWpxP6QR/Me1GjodF8p7HHS6jH+2btcTLp/4b1kvApOtOost4nV2
oby0bYmhQFwQHhgRc1rl15epiRc2GTpzYI9TEVgAQrRGTyuJb31tuFbiE6qyrI1bFygfO4VYdOJg
veBjq4WJh2S4TxwojUpppKDojMzv3iGbdrTaFztLCPkJtC3hcczVzKBgSLQh1ZcJeiLtbK0k9y1V
rPYL/KAbgMsEuoeKjPsKVMeRb+8zMkRFmKacxG4E6ImVMqOiZtLTnmEc8KRqUVcx3BtvJ4ZNotCF
6xzCmF1l/V2V8TMlEOAmtyLNM5OUMUe4Totdm4Yx5Ojd1XEMY0dUDlALDWveeG0Ph8xAKug68H4D
Hiumea1BVXQ+kwUc/PiPsMPoIqh8ez7yfL5k/Z0DQsfhz3RcYu3OMJYzQPkATQ+n1UmkrpUJYB+e
A/VTvVUGNFIg+WlaXdfF28rUh42C/jym6eMdbgGkDnvwduT4qURA9vaWkIfMcdlsWVo4gIjlNoTZ
s0Pf0PO+xN0vCsE8sdY5d/GJYc7u8MhAK+G7n0vn/NcWNIpXDczan2izlI2SMfLVzJ3J8U/TDWbL
jwiveAbt63LyZ3cTIEuCgOl/h63BQHEtdXFJWkwFiPn6XoKphWn74E9YqrLLSOH8b9uwonniTlse
R39fhvaIQOmvZ/XKV6PxRW9Y4IBAn5/2oY5jtu/nwFTZftKbYJpl0WB88vs6tGoOl0FwbrQany5T
GjPLQ08gspBJgxCNjGhPCFnzxwGnN8U5sn8AnI4loN180NBm+audwEH2xAKo96lX52CpR99/gKPc
tKKV0MsyhzVY1XMwvM4uDZOCgSHZcxYpKA+MtM1aRdo7bTDx8S0iRLsGKbYwtQtPVZNhaV0Zcr5y
h2LKvBeSGmaKWT35/QzIO1LOruY+3RUXrHtSsEHSo5zqQM5DbeB+cqddNSj4S/hBCG7oSRRVcgxx
hUbEqJ2u6X/bZ5na2DzFU6LE86XgB8EObAzahzGVQMAQm+YVby65z0c2I6fyqsE2JerIjYmYCnSP
YgtWVDzMvVn5wDG3ZTAVt9FXQfrAXaDunpEBmv7s21pt4EQS4zXa4Ij/J6B3Q/PE8nLKNrDqPuOG
RMcvNjaU9pGUf3dgOkUB6x5YPZ+BvD4Mg5UD5/Mpq2mWo1SZs+hwRCKoCSi8kTjMytvkA3k9ihiz
XjtuyDM5gVa77dwSkg+ux5iCvZp9Z0IvWRfKN17G7il6QNUjqlJWnIpo5wVCfig04os41JpglQz6
gHcArIId1hXFIu8BQaJ95f7H4QU8Gm+1h+ty3zZFAyEYMs6rB7IJR+R/HrynzK++tLpZLz4ozIk7
nMKs1qXLY3pGBvstSBS3ujWnCS4L2Ag2v0b2wHXPtNiSLtIIJMjjSRl9tO7OIOSDLRGwUwsF1J3b
jOED7Vt2iVUAmG6MCBr7bOBTCaqQSrn8vlfvsveE75K0NdoNJsLvadpW3wQ5kFJDW4fbggqt8S6A
U+81Drb/b11eZS2daS6R1O/NVNUBwyESJdfm/aYu+awFzr9iizv5oE5/kdHkynjoQ8SAcbxuRTMi
7ZcOEDrg5pjKa88GSn3jkhxa7vjvnR9Xq9jzbGNMmk09GfJlr7KShTyXg8868/t3Y090d9mk16ZK
xcRSC40KpvUieQWJgNI0XPCmrVTlFywELlQ9mHNts1LGojUZvbR1zaBRjkl/ysdtJvdA2cJHwh0m
z8R+vPDmP/KaLEcPnq06AtSDB2XeYHxTVzo8RwjKLjWgJX1zUfsqH4tkeQ30fcND6ehcnThQrLMI
3i4CWjJsgr+h7IBHpv6yd6o+1LAlF3i74STFtgjYjxrJt02vAlM26v7578PZXc4ha2ZNMGSMQNMC
wmF8MUU5+Cdl3bdjCi//9xWx76M9fGwUSXrbRqN16S0sPQ4msfMcwl6THV/lw5eTXOX7LcicNQe4
Pd0CTJVH/NMQp1zs47Rr5avvdi2ysU+eOq+zhU5ohPDV9lSQlBGinGQ0mQXEW5P54+Wt7UEWbBh5
2G2dtc3GJmFPG+To31zryXHJd3wB37Lr+SflKQ89+ReyFj0kzdqTTRguxVpSYgRFIPBaev+3e7Ab
h5731kU1qlTFX3BP3Jgs/oVgCX3eWJRudI9yAkZto3N6XKBc1bf7byI8y4uCFo7RMjygRLEXPjdt
qjW9+GYPn/9GeLDwoGulB1U2OZ1nM+0JDtVn8vnj/1Om+nsS35jtzrnl6V/jfuYAuigfhWU2TLML
pfUVBQjrcUfRtBmmL6iRJFrutlxj6IUZdQbHGn+zHv9hZbZAW8/8hSh40MAcJGUVToI06AWmlk1b
w2p5rgQGm94PPPJoANZ6/UVdmbzGT96t4TQPk5jP66KRhdD0bR72m1oaudmHJ8LuTnexCIk53LH5
T+btHsiWuvjMiv1G1wV0xJbbZAK4uQfiSDEZiw+cMCLnsRs+Dc3ebYofa3BiR7TLvqQNUOUTPR7z
pfdeHOxJBsnVIalG1lcbLtLC0VgXcBksh8kyObY1yofBRAKzpjU/x1HQka+aYfIREiII0ZUm7Yar
ueV5Qra9b2Q6W/i4+I8QGKnvn5n97LyzCMr9N6qqPZliHm3mxMbfYQc66VvoYcFUoTma3JnAdy9A
9/paf960yLSrBG35wgV71ZWXaPkb79EGNaKhyfjhC6QtOOf0QNemzFs1IDfWrP6RmQNaI/P1MTPi
o2KPyWnMj02hJ6II/FI8AMYAHQIMX5HP66VxTnAShF7N7Q74Rjd23dms/vKVyPbx+Ry+SsHG1x5K
20khQLlWsU9Y72Xnmajf2C7uggyf7Jq54PB768aGfYeuOicvr/etB9tHpjVesmkdcrMnGeUBbpm1
azphnORQK4D6hYJcOWOoZ+/kJqZa3FNApoI40chvciWCLN/9IC9LwFwTYTM2RGGsv+FKIlK9/Gjv
ZMY3DkPCla+6tkLMWEMK/Js9yyLWX84hjEN59b0Bfg/dSDeMBmOxA5BzK2Qnp6KG8Zc4sfHnwT5I
em+Xay2nvuPvmHk0jPFLydEclUzNqvi4d6fq6x5LJL5BBkxYF5sEW6fSbji4om3UhjnjHiH2l3Oa
0/ZZPQvLi6/YLYnX1DJNS8q+cp6BkImTgCUtDn85tQt4JUGOTkN0GfPH2j7lX2Yv4/Tq/fLDzsMs
N/WUBhg1k3n3K+eoAFyu7vtn+44D7i15VrZF5I9dgCE5/UeD4Q8UtKPMzPbLvtpZsE+X2NfHdf4e
rNdW3Wi7eVBeys+qzvip2nBBggG5GEsgWvDrrjwM70KTu3t8LdMf8uT+4QNyUk+CEWOdGtgRtGvm
hGYeI2V7Sm3lwmPozcZm+M5FSk+hLouGm2U/9T9eBOXx3XVRgKb87FxFDwltsIjdBiGtduD9L3Te
ny9Ro8wt9JKp3dA2T5kcVWJwyKUc9HMdbb70r+zdqxQSbaK3WrZ2JKVgE14QA4yRApAlDu7zhzIy
v/dYwvvge3s3JdhM131vAvMmyAoYEtOD/wFLeT1u2/m7V56v4Avl386kvjFPIS1nArTSpeZIPERL
ehraoTBqxWYbQqGntyhcwHhD1iJ5g34FRfXFJwNQ9Jh2atpSl4JtdYmVwzxNZoUJxKyq4khsh9r9
Lb+KejD95PYy75rrdQZP+bsg7NNm8plANtUJlaVDWx1rxFBxGvx+XaEwEav+3lIxpCghglE19a1f
uS4YoHS64O5Bh1NGKeNPHxEvGBwdiZ/aBLe1Ka30uyOoY5fSEPhACfjtU0nr2c40/G/hxVRHyqog
ucqH74MhEwnCEYwH6JzNrhdGz07cFgQePnrPwdJ7a0zrzAsGrkoSnPqGFYopck+YEZCGgNu3exDD
O1yj9BSryGjqeM8dE+6aXeUw1C+8Y9ZQrXwJ0siBUkYVE4aYPKsc+Az3BZzlRVDr9sfh5GOQL5CD
kSpcn7F2/vZMUpgsfLYAOzIPXCY15unETXM0ONA09hzgToFYCGDYoeLhgkXuw0dgJlx0+h/M/66i
woZXPje2n6bYRyarFx6pO3one4wzyMjkUKsDYWEWNPaC3x2pBjr5wn8lBFtOh5rafPLvWrBMM6vc
8QpWiia7ajl9XjF11GB7AevXOxlWjvIdCDQ4XFy7ve7A8MvxzzjMkd8dKMkpYT2ynxBW7HT+p3iO
RKvo40JiP6cx4ApYaiS/Ygvw0z/thf5fbL7WpIhXMMCbFzFr8TRJBbwRPyN8zMht8qV/O478kbIf
m+435S4uAmVOJCkyI+mn34LRQeCFLpmKxpVU7fVBp9HT9rAixWgq9Hdebe0esOIc0YR/L/L9lskc
qiuNfLqoHtvzVNvSqV+pvV34vgQ5KyXZ8v6aidJkVYuC/yJ0LyAdkb6NmBueXLLBkG+GAwzTNdbD
Vsds7SPWGZTW0Uqwf8r6ZxDsbNell1/+1OkbmIQrV8k7Yu6aLiqCQuNE5g+Ydt80oppFdwkv6m4y
SVaRnIahiIAFhYSXQefAs176IAl52s6OUjTqn2EmU6a5lfy3XNouv7FGngGodrrSxr2C9SHOMa5H
iI8DtuY0MCfV1rYYhLEZfCveosr6nvcF50eGIWZ9UR1g8FjVy6WITwhgm/t4AEZT5PYMggOXUhm2
UHOLIUpbhfkqMFbJ3iFcoO/G81PIZoSqVcl1pkozdeBDpRgxQQBILHCk95CaM8rVB4v5UjonR0hs
XG9J1K9R1K1mHvDz9b8cJ2sWtT9U2CRUbWOSSDZYZsujKYXByTUNNeoehW9eyg9Vm8CAY1BrWeH6
2aJkrOi6+XTDghya1bbyffZgZDQBuTyEq4DwEu4czkagVLRx8Jb9f9fFNvB1twHYNxIQfBLRbkZr
xPDkGxGy68X5s4eQtEfyTE6nCxctN5nrrkeN1pCvxwwKgJKHeqkBlWGFlgZfsF0QoKLipTSiAZfF
0ZUW56vYfl9SGd7dH38qRZYc8Ilr66URoPmn8Ky6q/0/8Msp/XiUETFZaDKi8es+eyIfIDgkM765
wCDmneHUMZ6kCW33b5djWuBkR+t+U07rANvyza/MgzX13gnYuv7/E+IWaoJRPd4NP9DqwATDUxGF
ZQzCv0KoWoSoxsYFjVQTJugfLmbFITgXB8vKeWppzOgwvYS36VRz+sgoSnUmizfnGGV8S8QlCac1
rX/6viAZpApai3IGCTZ1+0quXrt3HFen2rIaO/Ay2hsFBw/nSBaJkJ2B1TGWTPuxE3ngjukykkiP
3+60IdaXFTkHdYZianuYorbWG7lDDlGjtEibTw/+CNyOgH6onzAVdPu0wN7NwHlTSd0ZQC4GuF6w
iEm9nmRk445iMyeKX/MeJuT7Rll1uEv08zcdqIWVERKXeK+qv8lr3wWgDto9i7IVhgYKkqB2EBmL
6HfsOv6bByKygyX6JgSqt2QQz62lZ6RwSyzHmk2NPnVW1VH5UB/qKmsxip4OkysTq3gOWp8qtL8z
rF6WQ0uOvoELD8tHzV5vYDgRDN5RNgOzcfZlkzMKdLrD7JUisFk09s2xkncQiXe62UCK0cRToeKh
rSc/6nSJ8ZmRbIbdQZOj25chj7EDgfLx/9D8vGXm3ylbXb0EoKkgE9IFFsch4Vm1YRYnHcEKIv1U
35UFtRUrTeskZkhAeCTAiBxj6TAsihmsSt2Ky+P8Q1c12fecEvJRNPFvqK2ia4bNvYMbcTnD/46/
2BJsNYWY+JdjE/bDHldb8xEJTAgk5fFZoWxGJxbbZ7UpOcGUQD4dU8SSc7McliotBtV9+KzUPxxE
Y+jTmDxT/UzL6dHbc+Kf+BDr+LC0mEU09tnsgWdSSZGzCgxkJ6skrPRi66D2gOBDYLcEDiXRngWX
gjUDNDWEljEwdb8Tds2SBXjlIlI3+5RgMqHneZfCNQqTeEtM0nGIY4lcHsNCvKNnuLcYbgg5iWsU
lWWuhaSze9oIbO11exbwCOgbF2Wqk7UPfvPz1nwmxHQ5nPFrkB1L6zQPo3gCU9OHOjvxARymLpgr
NcXzG3Rq92eHwLqSvuE8jhgtCKOLIi4qw/bVzVB1ftlk4WUuLHfgIQP0wgdrrnmO/NjIV+cqHt3t
PSmuWhtSedNHne5du3jsTnFOJVwDzcZUSnbPjsKX7pOBLhRWxhKyn0oRpzLP06tYQAUbVUZbsmhh
O3qs8CCYHGwHRIWcUIeN8lU2mya/JmUi0e5AuVgSxzrIPIlQSLcz2jch1/qx6v+pJB6tMEn7aRyQ
dHInoUXBnxY2ABvIfXIx+q/HY+f6WHArvLaHUKCtPREK4woCIw2zqWrmBmvSUs0k9UL/YzKV3luL
IWXYKx3HJdBK4VFHc1oAUZwSw2a137KfiPWLKqe+ER+8r11lTXMDPmhDn+bmlC2ADg2S9Coi8s94
H0ZvH+wh7TDkYu/yd/fG5bQPM6dlhaN0/QzNh7qVKhm+wZByy2sr1l3jNI0WpdmAE0E+hNcN0qeW
YHsi5yE4sHa457x3bvu6aeY68cG283R416O8KPCNNQ56hkFMfVve1G9tT90QqmIMmoXJ2RE0sfEQ
qLFAl0BvaEAMkHiD1piji5eXjDXDLYvczPH8ZI5WZeS7QYh3Hl17ovpqq7ehrZ+P4mLXdTyHe1ha
xVugSBeo8JfQ+tpU5tu0fDM4vUcpk2qS0shFIraMPgYa66rO82mFyDYIeED68V0lRsHQmO/Vn568
oH0szqHw2KidvXk7XAp1sK6cP44hvfVKalc7FJmubuaHpZC3kJkKg57nAF8qiE8Ra41lGWvwweUs
flhEIzfG9O6VRZYXXg1w7L3eIOAoDDrsG68ZoiOz+U86GsV7zJClgGz3mRhlcuCKczNn67NG8yUD
skyWtV0AKG5yUnMNNuZgnma8+rVObwJk6j5M9iWl2XVyvN0C2rJZ0PCop7P9h4kBA+gXwKM8phXw
QHwZvKxCzMigfS86GHpWhPMzmscdr8Zf1cUYVrIcwytftWJ8VlMSRQBbXUMYGk0WqUN0hlixRqzU
e/lSM4vQGbKWc3buOSjcvYxdHPKTMqC4Z0BzWCO8axH1RzNJ+UWfmzg7uwqs9eRAG/m2UL0CgmYg
H7/Fc/cA0mjoCUNBKTaSQsYPn3z/fhTlZxqoAvFSE2OB/bp+XTnHCBI/fbVLYSZlQ8rNJ+Fsj/l+
Y5jlO9M0WiVdRvqbINydtPM9rEhQlZSLMBc4Ac7hb3Rg0P76YOn1fWIJuvcEhVifbk6Ph1f8E0XN
M23td1/g5UYZzjyoTY6nq4U32ygwd1xmMFGZw4srYvoU0q+iwLOtm7cT3YxChBaSJ5Ft8sDw6R09
xq46tYDeM8/acSMvaqxsHoYDMzQvV6K5rymUt5iN2+mqvfyG0ltF0K73QhF3Sds7vdwg1ark4ZxF
PYTWgw4Xu9AnpcneslStO3EJrqQjRFOiuhFaoBBKmvNReC02ZlJw3Kf3yZNqwBqxzq8bWJ3T3DeW
rHepL91Qu3OUjIwuuH9fhmpnkuX6/q5Z98sXhkAqByE8PjQk8aXZHBcNO+ZethHl5uW6U70Xt3UL
/Kbpt1dR5Gz2LtMUBOF1lZ35hWXp/nqZFK0xbd8QJBeIZfpwJr4Etq36vBPaIkkTHQyFnCcE4JKq
xo/fiVzmXx13kePYnd66OumRM2z8/uRc4DQSHujnw5BCXHwOJjq4bLrfQEE3XnzeFVE4ZHk7lu5o
I7cI2YY7sLhM+pZSK1KcElQD6+bgXgsMp08sPslJpIH0e2n+Hgw2O8UxCY3aqTVrTKhPuBC8bm/b
VwXJ8h5w5ocm+6QZ5K6bhUZxgTgOmrLK7o8SRyTruwy6xZ4aHVNSKBlujQg1+xsvJT3RoOfQQrgD
N+v4/bN2DpX6KwW8ULiaYfacDoCCJAJ5BC3Yj3pRsoUyH1Nud3LCxV7+TQVkuFHhIvo/IKeJlmQ8
TGufz2ml+8+51T0QTh4IG5znVR9YLUe4o8fq5xNCLpCtsDcznS1IiL8lMympd/515LTfVuDIy0O1
erw4rND0El3JE7CSNM8tqOVMTKLtxLaSTiqb8iMyDCFJorS30mldUQtr5i3z0GwHX5kwtbXsySC4
Q/YNHhvAYAFUM+9KCuELgP1JfIXMOSlMAA+T905CQ4rZ2MVXEVX53Bybh4oiwvUAnceINl4wTBnH
N4Hw7ppa344NKxSrHlU7NyTAtCcmzmBv+4Uy0FfU7jkOWYzsr+lDLNVMPPPF03nwLKedTZAvc9qI
jJMg0tkEALjRAwB1rxqUeH7AmLTkq5lrP3Xk6QF6if4kLLFeh328rjSD7GxznBY7WBBpwaQC57c/
In6nqgtSKyOg7kZQkZqQBWAL4tQf/69tWHCT/qTEhRShkauPET1pgWNdfyMbBoifjn1HSLTws79p
zhNuJy5cPHRuatP5RAutL5jZp9qwwtSbJ6ahTL6EZhUqGbHEqy5aZZ8U1QYer0+4Xg7JHtNvg6xV
WWA+l+BpK05zYLcQGGv5+DTaRJ9OFj9UhJpPQw3JH2F0os7pBQSAk4hWSV/Haji6Ixo3qLrS0yeN
+C5biS7uKhXa2VMJe6jG/nxX2QxYDWQNto3XGNggB85J8OKial2GF+ztfgvghVPtuH9NjxkyF4ES
gpi8uWRrdPESU2lANrWWX9IUIN7itLrnvHUNjqnGpMYJ3czX7TUZ0ACF/htPD/t7m5BDRibvujsE
wHET1P4nP4yKFyy6uheH8MjjI+k5NXy3dvRu7z7joPsosU3OtBsrfBC6UF0I4YzKCziSURoDr/fJ
MUAdwLRs1gsF416sN+9dwDNHfT2JdWm5ZIPlGwn1K5nnX7PDDZLBSr8gMJIf96K/u2qFZW9ArFDW
yJcF6L/kqs7dwOR8btgvQXXtErCJ1HcUCMyU8j+TFkXzgzExS8jw1ZqrFCPo6c3PjwTVW0SqejT4
JYA5Nd+pnDZUIUJq+K9UzjE1/T3LqzntdeayPVvH0quSaNGeYunMKjUlj9iUpiCUhmhpyyeBzTsv
kZTRkXFIvOwvYu+v83x0vy+7WerFXgNFtApeyagibDkLohmiwUTq9Dr61X6hVNu9YEN8Ht2aB4Yq
9bHW396iwZpcV+zE/0o03MMr1qxixls3PpC08wWoNuMYraLHanulQQvnago3dGtGGlEosUstHwtv
1+cqO2eCCBUYZLGbWTbnBF+ZMUvBVpywFXb39+DLclFOhp4y+043kCFRrUw3bTSQm02Wz/d/TJpY
8PqPlDkjqAVBqXB/GGjaf0kes40B9wZO4vjBd28zs112LQ5jwSNhGum2b7xAP8Nvxp9FNwkSjW+L
jFfqXC5KLx2DuOtYWqxV2YMrZzIRBE5aq/LsHaUBZWOlTMHdd4O7BB55eDAau5et5c7AlafhGoTS
DR522FCKSIIsM2oCCnaxHHg0YM+fM36cAq8qwqsYCaCZLk+PeDkq8dCjOnaoM9EdIRlLGhnyNbEO
qMsgDI+CO6BFlJqMHTABMjb4Iwdd0T6MeMU95hUy2iBCj8aUXRhZ/mNtxity4F4jWKixJPvq7uXm
PJkdIXRlyZ0eoVI1sQMBRruE2LvYGOshZpTpiBrawdCp6/0gooFtWHy7+I2x823CRPW6xgu5asWM
VzVtWMUzIHOyYEnEKFGQ+AA4UI2tUK5IeEt16umXrsCINaFkp7TeRRjoR58GNnCz6kwi5eMZFuN3
mH54WwvrkFFt5RmM5mZVz4ysfs1er53G9i1W7RKKRfsohQeJYfCDY4kSUdh1xUx4mgwU8EMnvncL
XhBofiC+CzWpI4BuXys691OopYGOZMDs5L59dSvn7cinwDBgcr/sLngcj6GDz+juG2mdWF8pfCbL
ujLdmlCtxIMF5JriP4WMiTMzsDkEV0bBEwrd7b0n6ucKg6fFhaSlOUI4snhqfzxCbKWEz/gvsq0u
KSW14wOAqcluFxUiGrf52dsJZf0a8cgNcUdGy50xMp3enmWgnIYcVK80o+kTfEf27IlY8r+y0P05
BV/AUsmvbAbnnbIejdXQ4JnXZZTzxX+3xg+m6z7WI0nepHF8UKLTk1AF+w/vHDeHuU9ZpQsunOG3
5j9ilJGbqCsqrYNctoIyIMFOarGTsXF/Q+XMaEW2vXWDSgeD2QBnz+2/Hb8xBLJx6YuOL+fm7YAK
y/Pr7ElsKJKDQ1T+wv5eMFjW35RzDX8SFfkzhCur5vBmF2hTWQxcRs94UZ0xijOsQZxiuP0yGDCC
eRgoaA0HoTLHWyX1cud2vXyEpX+Nvxb4Qv3h5NjEJiv7w1V1QXaIheIfdbuGLPuNL3LGXUovN/S7
ZXRAgR0PLzbvbeZPr42cZmk31X/wokP9rKLKwH+JWuUvQ0uFADoYB2hdixzslNvDuHgVVCrMy8KZ
lIcfErARA/rdFYD7Axc6Zl8RBiIDlusrF565hdVfMV3578ib6MLh0WmtvWHXSDCQZahCOSW3eBEc
yIIFPZOxk5BIyD1+1sa02nNr6FAVgELsRu/kb8WO/80yLunlXnzdXi+8PJU1K1eft3mdmHF8zdWs
A0kWht9OUenN2Ot/7JfGUftUBudXdHF2u4fBbnAFKdmSSjzXeT1MJqHAMfVsZzi80tGBWfQCd1U/
l49lr0yueTJ0RuDOMwhIdjEiLf6eaXWq1C+et+t6D7ObnskePxxshrJ6LkjUirN3Q0bj1jxY5RCG
6X2+N0+fghOur4lXh0SLQl0qm+fluZzluXTITpwljjROOOEHwBBPyBtHRMw4q9S3Qyf5qSAheh7L
zIMmi8OY5MOY1kvlIIAkGNUETU/mwraky7R/4pwQoSVUV8VnRE1XC1WIiI6w9P3AFtSm3tBzJFYw
EehvNPQFSD6+mH8RcikbVfjpbqjQJdzsg+DlpbG+Oe2QZBL4SxAiTU3+/J1A3NHd7jwagOy1pKEb
+y5WHfbuAxrDdtFoOY4JrG2DFD3seHJgiYj8yQzkJVFUtS38g/8di/E6X6njtoCd3Q2qGDS9QjzV
R7z3e25UxESVUsUqoUAB3OOOZJQk8MVKTcqaVw4peGzITHxTJVn5Neggn9nmXKQ6J6oA73o7v3lz
kWdMXwub42frixS9qEjrBmEBLvumKmcCFDLC2wuXql+nvE+evvUMBfavw9tBdrYKkjA3b4lEF7Nj
pzN2K652ynurFxpyyjYxLcXIp3YePerkbi1R5+5U//8OfzVX9EVoqUGFcZnjxh8qlrThWU0Gt8Fy
jKAFhU4tMoYndw66hQGyG2TAt2ggo8caYyVaZ9GT0eN1Luxtb5Fl8vnZat5oTN2ES2WmTv2U0eMb
OoR8Xg3f3mZDGTPXXTGY40vxgj77Phy+TBpQbOynKTAOTikSbUiHHpMb63pfkTOZ8gvrFP8/O9RD
TY6mAozpPdOEAjJ4zu+xSIOhG6TQJH4xU29TBtYqMrhUZ2D+bUFS4ahFaITcUbgLUJ23ETAwH2CQ
rS9AcR0wsKxjYkHqr8t0qIDNgneGKRcXqIhk5W6Zana8AN4SbHcBYaYzX1i0bv+yiv9giKrr68/V
d/Oa2DDUdqOfPeZpT9QxI0ygwH9VCMCGIfvGMudTEviXxrMi0iPHhHaBtqDUJ3hfkLyMp5w665J6
19gMNMiyv1MFKi5VvIucSGxeGJDuL3p68oDe1/JFo3aoTu3knjpe9GCV1ZmN1/AT6BYjZW6WZQqX
ApePwY3TbK110XmwWuBSL++lLBTtFiLDd1ZQa4VCxnEqOiXeRhkQ+CduCX5lFc/cWKh7wK5TWg+n
PKmCYWPuzUCMLPOMFxqceXCRpUe36xQGphZaD2Wtbj3WYkTko95k5fO0h82NdL+HDJa8DqwA1YY0
jhyr4ZxqxkepK7HE0XTBDZ1ob5nW2KRKbAXzPFzHwNll805NoLwXqVwbUE0UgKTYRQCAjbWOAwub
OwN0/hs5s0WYUKtYPP9iA0OOPxBtB8WH+A+jC51p7M4MbC6UvBecXPmiuvMF4+50k+WYtMu2ddnb
q5katEzCMmsJyCyJ0FS7RHxJp7JtqnZ62tb2utvZrdchJM8DXkIVn9tOD6hu+KPbFndw8kljNVL2
LujU/AZO9lG3Snzz8ImlJuPeHjEc/c1ZN+ODLnap5G7qM43XIoNCgQynH8x+7rKf2ROAOiJarcPi
6LJNXDXvUQynWb+JfbCO9bdBQv9jwBH5aX/45KAi2L25ZevZcanpx14wN+9L76T8w4BCjVQr52UO
5unTC4hjj5ATKOfs/bCFAufi8dJ7uAReFHEHLd+gcBWf7rEducCt/wEQJP7UL5B3P2CPLRVnDDpI
LhFiO4TfcjjNfIig0ZhYQr226w1xDNbXBS17UasfmOzyy4oPvd8yfskmStFVuhbxnletFCIovaei
6B2HHsgDJMGCFPXWahB64T6hJzsx9B/5Lcne7nKP7F5BRRIeDxE3UOxa/MIWGq2tYIRMkclnqVMJ
4lO8KZ84oQvp03+C6qg34xQUSmX9TbmFyfHVKZL3DSxYPuSHijVLXcsRk9gzI5YdnOvcrGjxQlWv
XYvDYSVzsEea3zrazETNSxdScsNnL69b3QX8GBUOWpG4N6AEdT8beSIz8fYBOJPgoBSrR6Sulp4L
9qJdVLdl5ui7X5LWPb6hhLO35S0vdI9r6z5gu8t/RUlR1ojvKuPOfFmLWTvwQBwtvL6REuOFWCpD
MQfZtQcF+DRa2xxYgxtRzRS93Dd/40uSKEYDR3QMudM+81w9iCmhLaOzlDjIBk9QbTpD2yHx21Ya
7NEbiA4DvtBqGEu4qFcP+Bcp6Hx5R8gzdL7yCyZhUKU9aPJ01qJOsRMRiztgyIeJovv/1Fpbc47C
zkC0p32mP5TS+GjvjTjchn5/2XWGU1xhYJati/5fQ9eoqVumK/tp8omCloyDieR+NOmnmmdqf0kR
93B6oRuCd2PACtN1bcQgwHbZh55YLvZYUmBNlPJKn+eXS/dIp2Jyq6i79/soV90e0w4ysE2A8tYJ
n4Sl4j4yVj+ZhHAcwvayz92M84GrwsOpe8Zr9qSCn2e58mi5AHq1XVm12tZkZdBsRa2xRSN2Q4wp
YSa8dZPNxgwRfklKL5yepTi72ntldAVgO9aunn2H1qfbD4WYfIMXOtAu+UzbqHcZp34tgHF3dACn
9VkDzzCtm0OAbIOhYvBv0+WWmqsbgUPWLDv7Hv/Gwc4AZFYdlc0Px8FDLY77UMGRJtrI92FFFH65
g1tAqEosbz3MDfpQSgkQTK6KmEC12J+BlvAFohXO3VaO0hdS3E/vIgLcY3J7bPtnftEsjCejCR0z
eOEHL12/sRzBMwasPwKCL1u1fwMLfhKi6RYHN7Sba8Dl1hZFL7Qxs3nEyTeLwwg8WwQGih+6ZV4Q
MaUFpZvMCt+tIDG72SPp60CDoA2XYEEMKaGrukVdLuSJdzUdOex4afNdWe/orx/hZnEoCq18GdAh
yCLf7Psa7jD47g+UAg4ZEQgW01ar2KVXbxpckc1/MS0wdMkx8z5ZB8KpUVBUokkNmKu5zuJ/3mop
0FE08sAZlv1aQIkgX4AcCd/dU8jHuq8+DpawwKtj7bTrgxFQ6JtaWmNPg8XDMhX/ARk1+Dv7i/5C
grZm8qP3lvUiAKibW0mFbiXKzdl7yG0YIXKktGhiPfZltS9OJZKiodp90HBpolpOEf96rWETpAHs
4yD3zZSI6wZxz5ib1Gafmh+LA7F6dG9RCAPL92vHhT5dsWXf+ylczmbCOCwgThMXeEEluRdnf0+O
WIbozP/Hv3YJGaP1VfsQlnTz8zPIMCXsRXbciwO3HVxO8CbZyoQNHomh8U6/xQ/qpIWTNR6fmags
NYtM40QN6kFhB2Afbeh9ZCokGV7izaGxhn7boSK1Mv4osEWyuTScGYY0KQpjdcdKkIILX7G6hRle
24RtHY9eXP+v4YgsLIYVSxCqsf2m29JLjVgmhGbVze15ijenVBMfwOYMyO1hokbzfhilOzt6JM+N
yBsVakbosWkWLMPI19n+l1u33mMUzZ3TOdAHvYsNLTNqKcKWJW9tFxU9fW5rHKX8+ATOPISR2qX6
eysZOoTT0W1nUhqQonBBHgJ6mt4h1iIO84XWPgMSM2GcwuJBWS6J7bZ67y03NqgUgdWz56znF4/S
fr47D8OfRdtnGEeNeNWSGLKAyThMb59BT23vFvjrhF4bBrIEk38QoQ1NMnoOHVPbZv+PDyYmJraX
BLaLJSOM4j77D7ksD/rqdfFLED9xE3mj5HzMEknGQ1kp4pSqpjvhHKklYZzj34KD6kDE5f7MJJh9
NsSuJhJUXojCo2EbiFfS86arIxUSyd5mME0VStl2aSDSW0J2YoV/x/0GAKRpBoSrsj1bxinYhR4T
WGYR0DjtTND4zemORDJhFkxXIpaqTKA/rgCYgZuXM3Z41ImicF1WjflkRjD8eJXwY0TxpE7xOnad
ECI3Jn5vDJDXfWS//2stsxv5SOlCdqiikzdsIKLz5u8WsBeYxEEeg4bguk8AZM/RCBHWKExQSVnw
VxawZZhZf8B41ZvB2nDUPNFs28/fZXA6sg1/Tx/sJxqxe63RCAZKpA671U8XVhJG66ivAOWPc0mq
uSzCbxO6pWKNkv6VKe7u0OvVZUthG9FZnt7jTvrkN/0IU92wKSVJ+cak3l0mS8qq99T5D7wTR4ug
7oMRacwccocp+XO09tFZlyJ/8IJQVPtOhmwH2Qv6sDAWVM+4h13NhXELKhd0LZCOfbFxqDJiix//
VzKp4QSin6EEilQ5taXq0G+VHlb6w/IAHT+MYMFlOvI89Mz+lQBsN7sMKdjCjLoUEPl7hjPgO+4e
3lfZWyrHpFisDc45WgD8nnp8azSoLVNsBOgFUhq8zBTDrCw0M12Wg1HWbtwMwuK85KJEJhUU6SoK
IXzVrhXtF3YnL+GZgSZlxDtieLtOFNqPBmu1Y3fQwCoi4Nz2bU34acJxAFUjWYktHzP6xWM0ffkV
VeJDg5YUIxH5p7S4fRSDZfsZggyKIBKFU9wDeRef2AMFdvIbvOMSdhybwK1bEu8nL2hfhhA8/A6g
lNFzMdw68cuP9kpF5AsllHZVJZwlbRAGO+F0UpHk9sc8GA9W2L2hOt0IpHTDwjSDqpNgjNks4IcP
E20vHFA38eRdtt6m4pczUWUD0vreKTWAy9id/UfIeC8TgVb/WtsAYLXFVh6fuDxzHPgXkRRqOX1d
slIvP15i9ya2QFinlI5DKh2H6gytr6IVMaevbpan7FjCAiivjzY8kAzi/ZxkprZTmaRPMmmtGHKU
qR/mno51xSaV3DO8IwwbgXrwC2stp2RylZmdJSvk5oU9L6soUbS50DaB5yMlEokyEqio9NwziPAy
xrHDYk5RvBk/7WIQJcQM6nlHcB6MY7k0T6HLzDREOAajEipD6YHVZ3dp3KN1aOkOmVBUM12sKieh
qBkHMryXxWWq84/Tkp2GnPfkGFRyi5ixL+j+bChQUC5+1yvQMQcM5MvTVKr62Ti9xqdcc+DI8km0
fsEcqafzNH9DVE6k80Rl1xwV0odVCmeWfQeWfzo01EHEFNrcNwPZDCGAlSM+nmI5mwRNs2Kk2XXc
mZiJcyOHc9HKVYC7doQqUFGCMcz5HsyC2gYIPmiiJ06f0h95jvWl3OM9YsCu5QVrXrvz2wt3Q/Pr
DL9h/KpG07htF9Ch5IRg+vLlyZWlPnsZ6A/uuEUTj4G1ADYg60oNbfPgKYROs+QkW+vEUov3C3Pu
8ttt3Upv8SpRxKx/+isZFKD3F47/L4mGDtnQdB0K16N0EkY/tNpR4ASNAf9AHgLh6XSeFOSowNlG
ywOQDtWO3koDlBYbYX9j0//wL8OIph6vVq0STFUlghpJyEEha7YKnygwrzajQMSGuUAXguvPClsR
W4QgLlmEVtZPCYpxq4426yp5x3WbfsCcXYyByX273XBgmapM7l0jWV/yQm3E+ennNU9WIIenvueK
i4Nie7bELFRXhxSTk61ET3xeQn5HT4e2UxIsKFiuxr+kwTJvySriAldKYWTURBGAaYMr2LYqoP1Q
bMztYcNKGbUsMOrg0wjuSMjr/Ptu2wYX2eR8iuP39urYc7WLRYRNXtxgsQI4ZNaLQAxtwonCWdcS
M+me2SASAISpA4KiozIz0uWC9HANAzDGy+WA5e0FzFPuaKjeQtSjI3Q02jw4YCiLJbkeecspnfP6
CcSR0pvpSHyCKLd9soEUD5619ITQZtyr1Gm2mGAu5beobypBikY7Ai1gtIP5yHjzINTCEDXKg/o3
I3lFPigWjSp5HW8uLKwhn1o2GQZA+28BilAa4Z9tai1itrBTPsU9FI8IayHNiEon8FCQyGPqDzcJ
quUBKJcj4K2yQt5ohleXZrWRUoj1lkAoxZL5RtCj38OUpklctlp+ipqD7SVNEuI05dPOPY7Qg4MF
+7ru6zQkrm9MeTof6j1Bx0p89MBoS+ooguPsgxmLJUjaosGV/hFTtboo0P8EBeLvRQSSQEu89BJD
8kRncUq3Vn3VSzpJIesaqwHKng50MQMbC3a+o/YOZs96ML1YueZEDBzocdmJrHvXHroZ9x+xLmVQ
fCd9i8XcS/r9OhUycrQ1DeT3Qk8qLS5zaZIq616u+xG7qZu8GLQxuB/7vMscEmByaH7xT7qoca8o
pJ94iJdr+8eYwHNSmv9lLduSTLeDJybe81MCzDBkPAHb9ygLmpJ8Dp2ZJBCeha4VrSbQP+QVay9W
EQ61DaNsV/07m+1HlQ15v56Wo18ZWdo5NC8ojIJJGcgkTuwxuVypugyeWsyKcTMWl6wUL0P32A/x
BdQkUea+vM9Zv7o8jeawbmsOkqru+KuPbBanVmboEhdf257JpIZxR/26pKLUJ/ctmd8fZd3lpM0G
BI16mMWILyqwJ/5aKvQjFcSlAgWPB2sQVYo1+Ro01nsvNyLsCOovwTpHPAwk5HehUeFDj1UQ/Ums
gqMWodcSsJcdkGwNaRaaS3n3PTF2w+Eryat4Zt9593wr8OAV7Lef4aq7Rc+0wNtnnXW4HQUWbh8S
+d0tCHU9bNflH3INJ0rXuUV1wlD6IcTaeX+3c+grzfD1QGMxFFOGqDFXcOWtCW0TKWeyjlkxxQ++
XX7W+BM5AoTHAvjxP48FAy2vsL9aZGTpalOPoQMfoDgicHQ9fzKy18TwsHkFq+imKLxFLp9dHek0
ieE4T6cjkZrCnCESHroHS39LP6fT97C/K/NVuSUsARux1jLpN9i3T2FJ8V4IS70VqnAFHFCX42IF
5+t7c/vqyZEGm89rpk2H+FVjFFG+DjL1MLRlTW1x5fD3SZowZu4/P7oRiPlNw19or1ERovqQYP5N
viL5fnbpFCdU+AKWx5JjWgxYjUKJaHbd5ex9nCbRobJNjccFtyz6zm2DGq3rT0BplT9yWA5WNgzt
XqBLYA1kEIm5M8tsn6aKPFg5QdYadqGQBz9ky69ICaDl5c56bmZv7MOp3dQ3Gsps7ggWDaWjTp8g
yxuCmBSLbcvZPmOtJhiv3/3aRscQ2wYliMxt3+UWve9j/X1RZlq3e7hklp3sHtGbZXLIAxctxzNV
NaV3TArXD+jfbOGH03ycOUr+E9GxUrpCnQMGq1MCaBpIYZPru/+1shreSewZfEUlF7G7EzVF3tEb
YL0mPNEv7bL2rJOO7vwtPu3lubtFPTCPjmCGWOha2ydJHlR4LnXuClEaPlOFZIMULypALQSkitJP
csejEL2UehKHnOQtRwffvPw2lctsKF26kr1QUVSjzbICluCh1MXJ9dAXBAY0YVdUi2tfRftY9Bn0
Uf4iTxRBkK836iJQGOUx/qnsmuH0Afo6V03sGzQGj5cgnTUnGTc7AI0xtTMS8ENW+dH6yIPTw9g9
JcVnEEo426pchMKHqboyKhFxVH2XfMqMxVA96HytnJPqsxWhPCgh7H2AYbOSmop7VpfC/geqIZPu
I3ZAwEy5anJK8tRSYgn7L3epJiZL3u7QSw67M1aMQ6UY9pzv93eqrxcY6AxNr9FtEwyyD6InMcsH
Ui3JcuVejPJLZRRDn1cOfx6ZSxwc1zj0Z1Q/1Iw1bLwF5sYlLd9zMr9Zb0BcKF8Lk3lkP3zWjmE3
M34wrVllC1nMYJvkYdAFK5ZSuzgIJHa0/PWtdwWlo4xsIvrtw7CqB+9FGuf6eevZO+CgOm6/pXmu
IUp5azDhINM3XPTbUpcYbVTQbbUThTU9HgV3gqsKjO5pny4xhR1iJ48ixcqAZaNVRppwXkYQMaB3
snct+TSuFUZcFVewwpGhtYUfHIPLfHdCesPNdJUC6gF2WqUTU2AfQpcy4/FL0SPn/ZdaOiWbiW1j
bc1Mdft0bSBwQzwywsZsCxJbpb3nE8SNVbZSv9vl94E32hoWmiuJwF3ZlqAGRNHcBTcGAu9v4sIj
ETKMuVooM3N+qpgGPeeZTgmfnKDdrdaVd5Kh5VVg0Eep3WqEwjD6f4G1Smi8wbPXj7Rwn4GhQ2CW
N939fDtDAmTyCs/FWYZjuvygFdej1xfobRolofPPwCL44WEsVnuCTuevWpIqBMVWK3ipKGSo30Tw
1DP6TOkqHQL3mx7wEA1XjXldJcqjhZdM5/39xIQzOWxQd5K32+f2Wn0Mh1z2s2AUsVZSduSp1i6t
PyCMSIftGEzqq6KTwXAN7dyLwjyqEshYfiowjP5PsWnk8VYmKIf3ZWQrRxFrFoxl8U3fFTk+gxQ9
TeE6LCdBVRufJNxsHC59C3ROgBIRCJuDhAlEr/2lsxyE8vPfvrin1UJvskdT/m4+R/klGbr2RG7N
Uet87DtDAx4qKrglq6cXu+GPLFjxZXN6kgGz61Vp10MMXsJVnq1CP0shF8uZAou+dhDAou+qPa3v
nZpVOJMzUQ+X3LPcPWQ6yrcxgF+iQSYAYIZB1M7atxmyVxZfKCH2bQ0ZYDEeF/cdU5ix4qHMTErj
yb5Co52msVnF7eZov0YTNNoYqz4k3FwkXaK1F71W1JPvYB6Qdfl7Ki3dvCn7SYodwcRNoq7Q4LTL
1/aSAMpBVJhoSV19vrI2LriloYazqqbGhjiE673dfUCDPQ72MiNiLkqRnSjL6ISoP4v6/dhsBn4f
N3v50gIC3TWULz9XtIDTo0hFmIp8ljO8Sp2kRDFdAhjzww/B46LjB7yLYTwvukZB4gvcNigzlJbQ
i70ldDlCKkP+wUGxVHCMV2dJuX0EStd3Tar6YdCCFTCeUZ7mwNoirleJEWcGi3aa1JsdzwXmqmCj
NHaGc5GfMyBXGYW16QpCdvgMVlsfz7HH4l5BXl04nyzglfutAO1q5rtVbtULpSbwGPicg7jH7FH4
ruweSowVUObHdx35z02UPtEMU9lkMI8bavdVjsdhU7St+9QK9uZBScNX3+7f6XxaKL0PeKJCl2zz
pqcXig3jL10lUgd99j7nIQwaBLWTVGkIneYhIdaFQRKKXtHJZo6YlJ/WaqwIwGJWQMsfnetzdt7x
QK9EgnWXLka1YHeeF/+wqPRZvFWRGhbKGbuSan6+sYH/EKOnfiPfiLlG5R5WdFYq5J3a1B4cSQhl
Q+n6/E6MyjUM485Y+5Yp0ItGhrsTsfWb45RwUxllNKV500smDUihDefTo4Pbz8HtAGyR9XA/9zKt
+7NTlbijpMhd5rCn0PPLRFn81Tjq6qUWL9ueGAPXtKjTmaImIgTl43orN70Mkjq+ZaYcOjxb2ER5
1UdFZtYSM+v0be21Ekj5J7AhC7X8ViZnwCN81khxN+LXcUti/7L08uV9wvdPOVjdAJZPeeXso6Ju
wiABPT8o8xEeZs/f+TicVFJlcnmu4Q7FfFc/29ZYc4OEHJC1JyVCKNaLQwPpzemQ3OLsk+rp+m0o
tJdgp4776KuSXbka4rgiOJAgv3YwdSPnsnPyf7DDguJ+qXsRsiZkG6Q7zvyT8fSpPqt1v0vle/ca
mIZsT7h5yRZQNTXj5zRT/ZP0Xw+Kk4tZgX/fTN3omAp5BklMCSAqaWlLFzszzrSh9wVUtVWF16FH
ycYBGwea6SsQq7yQsZ2TOmm1nzEeLXbxHIJDyryqivw3xYpt7iUdYYlMhuGRb/1++n207lCh08KZ
4BB5cVjolSaBxfwHYexKineOU5QE8PWaJjgVulnBKavR1KP99WMutq8C0nU+VrfVCp2QLKzxft9Q
wTK2CCrQI1m6Qd7K/reer+LgizHZNbuiL15qHNAMlojDi14B0RZ/AQvY2je1fKaUtBOlrKGFk3WI
quViFThw4ZRERQskhJyVDsuONJCpiNAH62anMWvAGyjUoecQUc6ACp9ueZa+Pda2mmtwM6M3tZM/
nwtgJoWfW7ukcDX8M56t2Gd0mqLxw3pQED55nBXMGxyVPz2R+PV55e3x34iKVNrp/0Iqharmd5s7
Dxotk7xdi/NABVhc6YjM68ES+tRm2NsVLJAYNjmPbtyN8hXvHLBhzmhYAMTxQsPLfS+Nm3ytW94A
tkygLrlvY79HDuTqL5R/5N8xd+hzcf+LM3Z1PWp6W+yiWuokdDxaA4RN+Bi0C0dgkz9NvVEIm6Cw
VSeIltbaJPP60OK6N7I0Lws4cDn/XvJQk7HbMyQnHFdnWiubc9Wbq1mT62l7GFl9kbnnqbbseedw
hf3Us4ZfxGvSzJ7MY7kRzhuEHM0Ch+8+7Lc7hijBUrrlbqvNKLBRHwdrK6471xVVcKT85Rk/sGmJ
WStM3GRRGXIZr23iRFPmWuAWq7S+TccLE4K3uE7F1ThxLIaiM1GH03tnUS2i3b+yR3lmhMJTPWRQ
mjqa4Ybpi7WzQOhROP4fNqF+wdprJPB53uWCzXabW6Cq4S8gAdK3IJtDbtKYS/n297QQl9buOqRZ
n0jTC0Y5/lE1R9Aq/0Bfe8dK+H4DweYtCwSL0o6iHVFNnCskZPXRw65OkB8umppFetlK3QQILRK8
fyLgyDmS2kDUoCKsFzBsjaYPwcYnpiDQ4ZqF5Zn0F+haC2KLiGI7gKvPSa2v1uVZd2usTUA9gcuz
Jnkt1ySmanczH6iYwtkbZnMd6oYSGDUJ4zSZPDQuPngMjE2kNhV7JC22Vhidx1gJ83BEdmZRl0pZ
+woE8Dr9sLxuVHHJ5RdkGxXKLaJOfOgx3FKL+ojEko/rFWuedJ0CLLp+RNeZZNqEzrny3xux3TVk
3ZamROE8b7e2VWyUGqY/ufWKGom7dACZ/k14Ug7b1xgZGKzuOjPfle8e6DsCZQ+EBYsORMJEPtps
pA85T92rG/1RcJFM1aS2Uvhbq5JdMbl7sgUDLJM7nGHXAy7ovGAtRippiE8Zx7HISgWDCunE2CKS
KCWWGHs7khK4RFmAsUNlZ+abXmeHBhyWP8yyF6FTx4qsCRz4Gjvtssnu47QWexPx6FSUcVsfz5Y/
IyPdc5b0+Glvvj4LAIpbl5iCdWh8O/hOusuOZh+VYyfEYFf3aF1vcydr6LrMF3L552/3yL3T4mzm
1IDVBUOYyQuagI9DNkHAOrsGwkcVm8pwZfeJHA3f5tuy2F4Obb/xu3yxjgseXmJ7yVIdE6BQYlr+
RJJV2dIPXABCl4rBtmGBTZSx5mAKPTvHvl8Tp9QMVih3Kka3f1Zn88SYU5PAgDynJSg1wuydgru2
Y6SLxbe5PfYw9wRpH60jfkc9GBI/WsC+4ONWeVOynD8tkxR9b7sjDoQznnK5RbGwgsu6wg1DD2ky
GkaNyj6Genp5kFbwEXzjBeU5lvG65Y846sf/RntZASUNNh/Rj6A8VDOlCb3NL8LTO5yFMu6Esn/6
Q2xA7ZKUGUiEg7BruuN832n15rPmhxNFyimRl1e5aGQW1R7uh2qO2rkwGMR6B0xpBUzuyYQwS/1+
h7Y5iTZp/AaEHk3go1OtdzifQSCccJH4jFkvRM0/IWMFipqD0cOWEO0/+Hbm8676EAMlBj93P//q
zKdwIUPvqU9k+qxAKdptasMCfFcKlVs1hFvNuL+qO+wfIGe7G7/UPmplASnup4T47efe+9jMEEDk
ogTi/xk5ljyvSM/ulI0h7lIvhTWbtcZPPFLQA1+gE2S+QjejnXLQKPwl2gK4KYDY6PPiNS7Dq4Sh
bbayaakm9R+fqSTa8LdYcBDLrLVDePhgkPsNN7L8pe/dDIyRlg9Qr5RjFagBRXlT5qAkHcU9E3of
NMCGo8OrZFro32wLlsIBeqnjHwJJSmrnwGBNv5cLDO+S6b7BO00KOCcv1fVrdcPrG9MtIGyp90L0
pMDn2AkeWMPYqcIJEhqPVGP0wvnn6IyqanadYyaBOPmxXNpzjttWoS659ypI6R0qzANdvOtQihMU
sE3mqhM32vGWms+1n07VQIJQK+05P3lIVnY5ire28D2RCV/XuWaNf0qQ7c9vs0Gf8g3PEmzqdWxp
+XLqNRtyxE8mvIwSAvpIY0Ouu/mCU9k9FNMiPGdF+y1C9uctKXcBI5EABSzpf7CEuognm8pXyN/X
8txuBWvebilb0elpNY4/XtF0XH0qGvdQLmI0mquCEaIouczMDfMWoZk95PTUcWHwioLkMo4YYeip
LQYkIC8AhG4+zGKpx8wmEMLkhz8v3rHDw6MYSpklt7QD1qxeNt5e34qRprsdUePAilkBcj/gple5
z1LiNaIAxBzUclcsJQxEyRHxRn3JEuvN/Nhj16qnN/nsSgAeFLCD3m6LHNPdlwFHZpNfRqRvCDvg
ccpvGqfgZ+ePbNuyqOC17j6H4Faj0Ma96TxuUkP2Na69tR5agLkp8HJmZMe9Q39OVOtsUpgm+BZj
s82dOvQzhyRHeuGSGr9Y/Mt2n5cLOBF/0cQ15zLk14AYgWibn2pC9veveiXM1jdMxTDIKQhCcIEL
j7PDTkCYcoPDhl+MBMipDr6EqbWx1myuTA1T3ODMcQRIv9vad/ExdzkHIpeZdjv2Kz2/fj88cheg
AXHGtNyVsXS+wT2HQKeZr6yKunD5XkgmRpnS1Wem4P1ZxG8R68F+2Lw/LhbyB3nhtzfyWSLcTUoO
h42GiijyCJrWN76EctIsLjfSyHf5Tf7v9aoWUlFUhjUjoDz76V/ivFFxb2AHIFsLvx5Cg4YXKNyR
19NsFGvVeZrFRi0MDB+xlTmgL0+tTCK1ILsoBh2flXvxFYd3BJ7EHSjctLYYDfHd9S1HUpiC6fup
TbKUwjRfOEuWv1LRP+YlwDbEvuLeg39MmsGDLKyrn1gYuO6fxi5q7EJhuvE14la71z1HUVAld06G
HqLK5CNbM1MoD3urmPNKy7QaFmLT30Wh4GuV8Q21jcLfB5DdP/MBEno4Aeiqe47zj1zA1ydWmDkM
lX2vcGj6qQx7gyeFGHZ35q1+fYNhFKQRGUz9YHCfEz3jt9FnH73uXT1nrWQvtBYnZVujwPEfXMr2
7g8J31Wwlebgzy6P6LD+DeC+JTvbwiXHvct25lh/c3+OJCXvBzZxJdWQ90XFUjLvs9hi6LKyx7jm
zK8BNiHAjirg6xt8uGjkw6XyXH4aV7baDa2RZ0HfoRLeuLB3vhoCMxNoItwcX33kIdhca6mJR9kn
R7wv7AAVxXTI8frvDX+edrka2aL+L5s7n8CurHIwrfjGFKBF5fucu0zKNiKtG5tCI3TVU9isBwqw
Q27EYVVQV8UR5Tn0KCvCRndEVch+0bKKu2q8PcDtcwgaM640YOB95sncnZT3cN/d95Hu+T/LyvY3
/dhKHqm0iTSKAixLXYqnaBOiWZYnqO92uopgSBI9i5Tk8LcBTMdrSewEqR8A67J3aT68UWeoODJZ
7DyCCsdUkabQgHHQD+UIq3H5vkUcn7XNv+yFx6dNq/nR3rBYp+DJtdaViFyvoYC89ErzZfYvJVb0
NXWSPfVkGLpZbF6+s3W0IembiBYjNj68nl/fqCrTTHb/Wxunzp7VvsOtv/Lp8oQNb6VrPYjZB1EP
Igvkwoo/s1PDYF/FBFZC0PwFDAX+fE0KYuH2UK2yV1Tv0woh6WYsAY+7p9n/dVH+TRLUz9t57xEg
hWQ4xNA8dBgJ2tw6679P/Gd5/tUc1xRPnqP4ta1KAi+YA1g6qCin7H8Z7716ML++E4Wt7ESNyvoL
aHwlApDeARc4KSpvc1wj1lU9sNpEgOtiGohF2YdT/mPCvGOfalNxu+sYeIRiiFrSr2JXNDSW6sIB
O0Lk7+di4tLSqfWEl5l/Af0Er/UbOCmuU9NbfXh9pJtPz5vZzqPryIHdsltTk2KwPorJAKj6HWVT
ZSQ+HL6nw9fUlo02byTONF4tuUl3829vP6VCdAIBhqN7KiykbQPuJzfYKSrhwR9DHWVuLKO25i5u
UpaUXwq9ZcPtOKnBe0TUiRhd69EdDcoxFoV5ecMjSyP8feqZ7u1NC+V4Tyx7gPyGQMg9LekztAAY
0sE/wu7pONRSmiGGI12KEZLOdYW8nGIF4Onf2iy43Oq/eQzXMMU0l0OeADsRX7p6hvPyXoNSkdlj
YAu4yMhGUCslxArib3FYUGL2WXSedS0uexCdIEk065KRMyf/SM83WAtmuY0qJbkxScdsK6JU3rIl
87IHpQ4DkzPCFcUdxLjI3pU3fg47sWiHZwJ3ScLtbzXjWsfsFPipE0AD62SQzFCwD1Z0Ywd3skly
EUxotIM+ls0LGbEKwtDUiscGhqAp1FxhGRtlFMvLbraukop5VUuqFLdaUIvRT4NpGaxvKNWfWqxQ
k59C1F+jk7m2da4Hxwl+jP4COh5OewvnIdsiWQVMdoTILS7pYBq6s9wxfEpYmJH/St9rtTyDUbLJ
sEsFNWYHI5JnDozlPAYT6mIZM2W35U4kM6zboQdL9WFSgdiqI8aYAMfIQwmF9wy5/EPZCKN7w28Y
hCaQHLzXeaBDZEQs1o+y6Hb/qJDJOORMSP00EjjOUEKE8TnOOODkDR+HhX5TDWXNuVY1wQMgyhRC
9dCtnWohgEhgy4z60FTMfO11PlraAXYD6v/DhIst0rd6FfdO9OkNTAPPlTIvkjU6Ogie0T5+Q0/i
AFTSM+2GENG36Bgc9gJZELelIyTabS/3j21E2JSvy7DPe4BlKv2Wr4aKiyCeP91DTCJgHMKGKDZ9
vW2K11Gq/2M/e/997Nhn5Tg8TABuW+77POto52DKxmCZZxUA22tbsQfte864jeVGQbx2Hz9ns4X0
8NvzfyEh/hyLCXJX4f7ixLYoLTPvlccahTN+fobLTGU3ZYpEf8c3Mf9KnforgJQ1MUIP5bO1bgDy
rlLQsHzYeRTzFxQZPFjaHZ+/ZcrLYeketiywR348ic+aiMcaN4dRM+n28L7ApPsPxXLNTb6zE+Ko
g8Jsz/7hbmuCwxDG6YfFSEBDagylIQnK2LIUcIDqT3rCbNx2RkMNXlsTo1NPJVn00YNw4TMNqWo+
UlSJ+j19INi3tYkSc9upC11WkhFnWSpTReviX0bJ4f/Fy17jQlN0Vg/aQUNLlPUqaPOrLSPURBf1
gdQSZgJKNmooTYYp7QoblARXvVJOcb40jhGCITFQfwz5BMeQ5GeH9bD6dQ6ggccUiyWp/HMQtdXe
UvKO6mR42WeiiwE8wSMyf4DuauukdOt4eP+5C0CzXS4DPDjBosp3qUHjztljUG6xUOS9/2LpNrJo
yLVC1Df1ndwnNfxxM5yAuY7DHIuAIy1NGLa0144FG8AUBmW8Dc/LmHI29lTQgOYHpz6gGEDA1ijM
+qT2KsZ8A7hu6Vc1ayUqQq5i33wZi823N6Zjltmzo8mjx8QtTeD9wCtobdCPSCqjnOKL1rjC0Dv2
QqThUPZqE+X15X4JLrmHZ2dL54bP+2ywslSfW/d/+JFdGFGr9iNBpewnQa845j7KN+bnICKfQUNp
GK0k69rSzgm4XW0EgedRE72lg0jr/dPIXTmAfS5L93KzYSB9keBUq7WpvXjo0pDH5MfOKEeoNyeV
iVpqunjjeYek7Kk4iqQjUxFaMqxxXeavYtuNMxFr3KSGThHjMe/dQn5w9H4TaZWpwPcRbNfuhp5x
Fkr5ZJqLesRL4HlsiefJ4m7CZYiYArSKr5j5fY7PZWsNCKXqhND0o/b7eeXddRBO4sMS/PQMjBJ1
Hx4y9+wpghFKuMqqnpN+JUNetkcCFhwMa2eUfSGEf+L9LEtUXdMQdQ0bI9xTipFvUsY+M7JVgnC3
93UL2gUoxW1zQGxLraE536PS0qUoQJjKbldRLaXpXT1loPRkV7U+OR2rZ6h9ro/vVkyuN+cCxt29
SXsm1NjYPNDQuwhjNhblKewh1FqjNm8Uf66BoNHW1SnCWL0D76266RZz662/cyd2OIndCOkT5H7q
D8iqFtnanFACpfcMJ/xQZNwZMbnS1NyO+xGYXuQ0x3mc+vAV7dS/R3nyrA/DGVUn+hq9Hw9XU3ct
VYvln4XwxFmbSxToMTtYBtOywfkN7R7SJcEEKmeqY0eAfcGhclUdPWzHWjnFtJCiuy09B+X10fBx
B96zjxhf/cVOVtD3/9vec677gHA4dimBoGCwxH+/eH2f4+I3kjjTHdGkOOWgWMoMFdHsLXVQ7fgd
on67jQKyM/o90jaXiwAVpJzDYHTXF4XOxD9ehiysTGpVwTLDk5iIPNPCs7Cdn/lAUBBOPMqfGpxw
aiEexOcSLG6TeswMB+shCn7wgmMwCV1XaPf1g/8jHrRDlv0QBYMERTC//Vopx0heBiTjSUuPMmav
IzRuxRR+lge61+RplFv5dPfvsykI6AtKD7LJCbm/AQp+cV+isjaPlTpYnv73FeZWkNFReVZdbcNy
5CY5BClIqzAJLsTmH/nODiV5U2Zv1SaDqxX+HkaQ7Nx16popRY+mKt3MAZEvXQkEA2vesM+tlWOd
m/iX4hc1FjTQ6gsFRMGgjdRzSSPZzdbWQbovmD/zR0ufTnjD6tXBYnRa6lyoKyyBHCiMIcSSxHmz
5SCcNZ6nHSooBYMt3pAwZcHov8zLH9y4/fpypjDzf1pbvbeQqOi6xWwOCItfQAoY+2Rcp6m6hOF9
zUoTUbvpRyfIWkt5QRG5UTkG3bKr0IqC4OSPPtnM49Ujs3i7VlNNkH0d8kpyuudS9//SJFgR1ZY9
thxsK47d48Lo8/ceE0r5I8CpvMMvGe2ylEiZx9VmpCjfYMX/dbJI0LBoK96+iXh9j8ySRjaRq/8J
UZl+CTNuuKRDPNTNb/4zXtV99+sgGgA/ztrFa0cCOZL3sLfmzwmgPuZpVgicO1nsvbX36Zzxf6eU
Wri+BpG+hqUgXxxPLQvfziXPhhz+N7ktpJy8ZIOUTLae84o6ipPjN/uhA3qUw6QUFrfl9pRS/vOu
5c5ORB1Xl6nfepxkE8/BcZp3fQBkV/KgUjiJHW2Fv1GHAq1wsjxQROsUpfxmdiftlBWm46ln5jAc
ffmZG7Bkq+ZKoR0pkLprPfapRS2bsOlTJvUnNp+UkPS/Gl02SdTvZKqYvtLIYfqnx/9wxIeOtyxO
UT0+N6aLoDYJk4OLDjQU5QI818k1eDeOBKsVdvGm4egO7xh3wOKSwR/23bPjZ6R5huYPMPHzFP6o
mprBuBVH8a1w9JOjQvtGPdQWXebT1s1/zkztqjV1FpKRMb60ZEMP6UFg+tYiuZxD8lG+e4t2xWSp
Z7AK/z0BW6YWU1H5XFEz2hchBGPcEDOthLbTdmT+C8A/5YS3fKxG268b9pyb50g2gw2cw0m/p6Mr
XzSWzlD/RpfB/x/p187gZbsVEwc7VpXHZ0R/EIp2xIYMOGvhBMn/exQ+fo6TnKnYNHi6ffTFazPl
5Yqx2cJ5UMQ0JmjXQ8L8IdNsUR3W6aBHriwcZUbhVE25M0cyi6OZ0FjOD+QvV6T3IHLijNjK15QP
+HlFR0+uhdnAxtvWgUcly9S1IGLOUKSh3IECfANUM+q3h3qf7ubSKX1Nxt+sG+ENa9oa04VkVXaX
UDghmmvjiPNe7YEAHTM6AEHoTsnP6sqIkE41LhgHohk1TXU0K+7gp1076cVndVzhsCWPjLEDoKPx
L+0l1XeiI10YRHj3VupiSYz+/LUqeupsJb8YAFlDZr9rCBmii19aaQlz9Ls9JmjOfoVXRMJsxUO7
gSqmr/6UTcCKYNh9D9XIB8yJJyd3dZ4ldxGj4wycCQMfqk3a8t3f4EB7GtyAn09fwr/ve+mT85ka
MhAy0CS4ufzIcOqkH5Ic1+Gv9hHk6hZXRn9LN/c2cUiYIZSKhQ+6bNL4uXGieLlqRfLT+fCyqTJq
To0Ef0JDKRTrhwEC33pTMLbQgvUGUPm4Pe1LeVn+SeOtJJDzKeztHOOUABM2GtQeWDY/PuKD2wGv
w5oump7B+tRozEa5Tgej97d04mUEGxZi58/0jrtgvWEW0MYAL8VZfbuyuSVgBXhTzliR+lWnQbm3
i0QkdDQWIu73h1K3y+IonYTVhQoxUPFa6ewbsXsPKfyJtDEiPAyo4c4JAGwnck4oKZ3NqcoKkU/y
vXnHJLBTi6AItOhtbvivvVn5N7jhIq1qNypQK7Ck2AmsqIfZDLDxJmkr0YjClOtoXmdiYR24A4pW
uPRldFTZyY8qcLSbHeg0y1pbA5Mj5U/3y+lQ6gWaxBjSQiNNnTyQibDfreMGHC/6t3wFnVY8nG0h
G5V3iAAP4Bge3qO0+HJr9abBAoh9lods4+3rx7pcX2yXupKNamQqxlndsIbzRvcj62qV+iJLyjh8
6Q81GxIAJPM+I4OwNRdMneDfdaklJNz2PbNTX2QzCirvW5etARUZvtZL/41X/NM2XtWgIQn74KkR
zsb6UwvRxXjBb2PxAaSpmFiAPO61PwTwC7RJJsa2Km2Eqcj94LFL6xqSZ2hgL9xhISqxvILnhou4
aLPjHA/99SsMGvr8Z1bx8Zmd5MlkHdBLZKyMeY44KC3IH5A6JlEdqDyC3LRwyVOXi/nWr/ctCzPQ
iScLk3Da5bCf8I49fAHvEWZ9T6XjAJyrKj3F3afKeFLL+OObOULpTikLn6uxw5zIcJm2LCdi7C03
4bPecNkJ3xjVI4VFD1LcJwol7cMIAmi12cmbzjEjGq5IX9qGX3Rd+NprOYHCQCaD/ccfL9SpvS6Q
NRgkKsWrVP+6vvjEFblQG8bZRAIH3LsLXwqC/Dx6vdHH9tN0Mwpo8dZw6DOwgVkYvbMEk2Nie6Bw
sgoDPbgm2SxYu8liltl//QUtw7/80/HUM0w4vO5188x5ywTYmwcVCJCKPM3V5PqdwbYHXCzsTwEj
1wRbHoSR8WdJ4yXu0w+wpI+h1iDxYy7OQMKJbccR121tdZsQGzKUGULdY29m99KRa2CVJU7fd2IG
pih9+1HLJBlwnTyxaLdy9t3I6GyMk9PP8W5B8hqRAjX2z+Dz2hh8x4wPj/tjNhtntNe4YPKn1khY
P2X0atoW4YRFjPBYDN9YaSu3FVO+SQ/V5yr72Wy1NcJs0ehElqlp4+RIqZjog2vr2PWjpI/gRM15
XjtaTWTZsC/s4L/+tEtC/lcrnqtQeybMZKh7GR+X5C8v9F2kIVmOSMkp6PGA9hhk3N16kmK8mN7n
GhyazLG6jp8K4iM5pa3f6bOURO+8/5J/91+qlAb5lL38kFamgxZOKyD/pgNul1n6cg4Q90t6ann9
kdTL8e3oNRlsphtmKfKM8WAziSvIWx3w3wefF3zFzcS50tsxkgwigzqcDM9fNu8TMYQMicB0Y3Ij
sulJk7ez2e9URHSz2T7zTsEmpE9h0DaYmMg3xWlMb3DdATqBxWsF0nZFo+PGry1huNI6fa6q5ppW
LykkHrWQeWMspVFpmJrHXirxo72nn2fZGXNQrlJSWMYSB7/bW50eUbUEmjnyT/00E0XWOzY5Zf6B
3dTEaL9O3qC+sL8iXYKyR4MU5iKxLrmF82xACOnoQuqjPPq1XmhHbE+j9js3XIIVlAxb8VmVeYYZ
QZrhZzUzVGzrcD9FuUnZeoeBaNGHqEyfDBusYd4Llhu0sZqDMcM552In/5dbc2zm4emmcv6AptYs
QR+Do4l6KQART1Y8VYq37hQ28AINlwfVeEm61G8jOrdKqyTFeOcdjlqne5LyT9zwlnwhqAsnyvmY
Qn7hWNaUGZ7ab9tO+VmJ/WwTiDoI4V0WjPXLfNM52kRDzNm0w+LhLASC16xrlcUE3mFFbG02WqhD
l/9GOl6lm6ZU2XpAn16uVy9OdqRZ9ilEYNiPo0dJaTYiYGUf2Vlqwd0662Eunx5b2UxjYQtmh7wW
Gx5Zge1YmnHJnjjV7KFxCFEoQJcDP8nU2lrBCxAHU4896m42wN3z7hD/QPkmo2DSgKuOuSH9BXmh
onnDPkvRvdQppVudRqH8pw7NjNbFv6sHRPpVkHo/EgAhwx9rng7tINa8gYrn9T769xWTfKFWfLwb
7Gx0oVE1fpCq6S73ikgtI6big2NDZiXQYQlv13M6tTMtKRxerLNsafUu7/JoDp/o9Wv+ojoZYxig
FTUsvZ0GIh+6+YHC23sAjt0X7H1gFXD7d8RcGBYileJSBOpXCnfKRY3s+uu6/G9L0bqQTEXtAP4n
hW4PmVT3pf6IC0QDM1Y4A9gra9HdADVWOy1uuYuOKhcZ1JZxa9L0Y0wdblJpKvchr2LMIY9cZ8/0
jxNaVEHHyO+yPb3UeygM5la0lCohQpInZE3vH4rFVLGGcnRUcrlXum5bElobf1KGf2i75U8j9Mbb
qLQYumoAxgzlt00BMOHq4zaRgt+/51fUsNWKMPEJQuryEGQOZKD6iMniXkSijbnKPv+mZYyQxa8z
C7VLFNBdo8omykDHpLreFnEhDV5BQtzXOGtuFxAwlk2FV2erN1wRElI1kGpAYhCNRTkImxzE2Wy4
K0iShoO/EPv/Nanaq12C135EEgV0pUgLIzxn/Ilw/SWmOUmLoGAmejiWE9nfT3P0RjvGFb7wEl8/
HA4alX6S43svjkCCew5PJGyngpmjNkALfgiD85u4Yp/M/EPr88J2s+wFAabCCcfmb9mSxfFCPZyw
sLjq9OF9kkBn4F0LO8Dd7gdPKmUzT7GPRkPvMna2XvpRb1uWvcuonCvF0wauk3xyb5ewcAsudkO0
toV7iLgvQdY2fJO1/zPOaqQ1Tgcl00UMOjbnMg5Qz9ojABeJEDUz7jTNBdz8asK7Z98PG5oafZOO
ZnWpAgcgb6Q7ekxwf6arkMIAaBce1oPrPP4Sl5EqbDpBWzkN2Mn7hqL8vdmGQOjclzeLFvXoq39R
77pBxuokfOZAZOxlVSDBDLlN8j3s83LRjmDrQXMBSP2kC8GjaMyBR18VNAasJAnRm8AlbKy8lkZ2
1V4rNI4XFJ52sN+bwTyoWSuExQpFFDUMDSQBT/YVjy57CDNpU3N+Dh6+fLBWHVD983ScozirG5JU
bXZmFyyywXwvCzI0KTeIb4Tr/RgRdvQRizGxqByogrD6SlB4PLXE7p4ceUYhmxiJ7ozpCV+XsP67
viI71vHci366JKRcYxk2EEITmAqxCuR+4Hk6/9S29gB31fOTxAtE5f/JVFkpQ3LETY42abaYKnNS
bJH6cnXRhHC4sWz0+b/yTX2pHy0nmNBhF6mXaqCW4VbX7bRN2LCSzHr+ugdrGDiAobARmdBzgqx6
TVUQaWv1m3/aKfbiYHPjcvK0fZm7wm7+yFmZi5pF0PcPTVUtW7RV08B9gxxEz+2DF28ET6y+XFvx
1xguLijBatPvIcnsMLcOpC4jPlDkMe8iA5VMXDD8LRd/c4SmVPQi3+sDm0iwV6CoQ8NPTUrWX3f0
CZr6aFj8PFAv5wUH+7+oaeweTk+mlP70IqhoxxmZAaExJkOK12hEuqyhiADLWFHkJIor0iithFb1
D0fHhapAbmFshMXDeS9oJzoQtS73naIzIgetxCRVneSvJrmPjpjhP7TsKWEfkw/URUjPpBSSawjW
bR2ru7pDbVNJAx1PzvJ/ScJF3FJNmtug+BJE9dczzUw6Vw6xExpto2tD1bb+Vi2Ptrt36zlfXIyP
EsZu1+MYWkjDhqBjdEh7QvyNyu/EkLO4lslpBcrPM0Rwj6EpBHGCXmuo+JpZGdLe3cGLyN6n+FCB
GMrJIL7MRn3fZq3e2CtbWccA50gduN/Zxy15sRwN9eF98ovg1QEWa4vVnLYxCIrruKczlbgYQ6Ws
msCoREsv41RfAddTSA8seuz+mHlhiwOSYeqSuD2L0dxsnLO4oT3glO9OLTjYrTZjKGgfqxf95RCW
LmhgVp2d/bHPogf4EQWIaJano/duPq49MsxlqsI1jXLEbj0/dlpYGwgotghFprVwZxI23+9Gj7PN
nfQNqL1WJoCaSyeWbs/Wn+3zOE+KjS38eJlhBjZ1HP6qslnoUvQc8s5AG0ASZc0CZOjX9EQO7V8l
iCOOiJc8qMfGZpeF4uL09139J04CAnsODvWHEt6Yhjmj+TiLnc7NqLK8NNuUl0brAihsxPk6qZLo
4eWIik1Be6iRp+xeNwrbH3knHfPGQz8qb8wCbG3z/7QxpovqV02V8m081XrGkZrDCd0m1jKx8jtV
fA0W5CA7tgsZwZGR2C+HJ/YWSwaqYXuIxq6KV3d6yJw++uaM8uYCxNhdKsoH+uXWXNR9NoP1S4R9
7X0lrKQy8Ndm7HtgdUuZ5bWs4g81TfIy6tYCiC7Jf7JOjfw3DbMv8anIKoHAHxDTy7+kFpd93nx/
9Bi4zaVSW+wqgFMJDxaBXFkOOkqCU1bRgk+cAG1i/u5kDwaeEKq3cYtyVYE+oBIst/RNStaRAKWK
6hmYJ8D8xgGKkARhiKxME4xjxDSLTE/2Jek859haE+d723A3uyMtH06TL1J8qJhLa2TndHrjMjyV
wrSzknE4RhGp8rORsrw6/CtAmO761gIr2N7Dz9nqoOBZxgmyZR844AuJG3apMwpqZ25kBkHKc1k7
EBwH92nU/tNZL7YX03yyxFWndoA5CKvAe3kOCFPk9mtCQiY3wbW/mt7C4ahV1GP0jO0WzEKh6qoa
Ikt3qaR1BdbhsJKZRlxh4RJM6LAg1IinKMuc6r4SeNNFbdnLgOfymX+o+EewdY0E/g11/1FRj9V/
mHgIs+vWVLIyGtI5GY06WC5YS4cDWzkcxCmj5QojTbZ8Tn2Jvgg33neYZf+6UoYXyIYk5bTnMBWM
6D4M5SoBBL4YhsW9UCuFFx29MYQZwfc0/jcZ5TfKW0IUHNzMnV3+m5nkOaTGuFgS86MvgWv+HdY+
OvTCXmWk/VONYF6XVwifXt5SNsiqAv6pelk1qvPjPEhkWeVrgRfqb9WSqzeVuVogkDHdbFwgj9iU
KNulAQiaY19PDUIbpIZpp3k+zZKIClYdKoby3euwmTmy1ziphUHQvZL1jxImLNUCOYOL1eJkYdA+
zKQ2Ep1tpVK0CWmqek71O9Cl2NWRxWNTrR6NX3+w4IPVqQrf62yWTQYLhLd+O8zd+H5B8gJp3PWB
zJt3Gdy7S2BKVe35kcZhAmaB05xu1N4PTfD+2QQA0oh2Kj4VBIGpDKIYFP46RmNgHTyX6lnY9evb
jahQs1KNJgAAS8fUBPH6Bne0eqeOXAoTtvo6ncZoqH/LLbLAH3KJRvKxcjY4WmNHhD3x1jMT7ift
X1TBiO8qQs9F/Sbl0CjLUN838+lLJA8eBlavNe1ht9+Ar6xuY/rkm2qFSzDFbyeNuwXYAYpSsQsr
EF2keQVwJckV9dEAPhhliLxEhaAOCq3y/dfaT++rEXIcMqtDBkXg+2oxrRbbGdlbMKIsQf5tkC7o
8oJuZDNL0j3zB4xM0j0kF73ECAAChTM5B0WYbIpCvujxJSi8SQmoEtttah4fvC7V7oLtd9Tbd3yL
jA/2UCSsevr82OuTTvJuIrMciEalzDKMvSfVL2D9zKPqUSq4ityMoH0vuu2REHYBxQPpNuPl6vF6
ay7fHA/tCI4az8S25a/NROlcy+4xdbX3Y6e4FLXMFNQnT1Ux9MxBMxT3DiBJ18C7mkzd94OVzhEB
gtms4gwQ7C+Hm082Ok0hRImmt3l9C2ZZh0efiosu4yW9tbMp372oMM6ZFAp1PNyivz8wURlC6Xo2
55gp4zvJXuZp3ViXrgbATk4rDzqV4IUQXuAteZYOZT/NgwIN2bkt0AUMmsZ76cAYo9LNeammM6RK
fjJpHh1knWaMAmqBbVHHxhh8P7QekwWGgnkJskl2OwbxRRzAjsW0+TQLwAm4B5CD55y/X7HUNXfn
hlxVybh0a9bZRu2dTZzuD/ALwN8TGEhOcZY0+I075Do8ItfHa7rwAV5a+/6w5mi3jlbgL/B6iagf
bvkPUAGerpzPRt/IomjvosQNm85LPE2HEbSNhlE3XUssaVoMyw9vDTzTvM28k9/rOk4bhuVGlfCx
PPq7trqWGkXo7/n6KQbO1i0w6R4Ezvmw/YMoZzuFnMcOEJbQLE+b3lCjb5PyKbLP+MOeXC+G+y1a
Hfzun06odC969Z0XSuKQ302UFj/9hSuQcT34VE6vgIPVFZHJdnsSQXbmL+OnFbyBMswHY7xSpsrE
Ux9u8IwGLnBuD/Va4lNckXHGmcaw6QHCkxx37rUn82poaY1yvgZHg4oc3vt56nk5NgXY/1hqVgLr
M7irlFCGm/94HjOpJgevfeR2lu5zH1pwNxfcpg0dCI+BEJ/eN6zu7PUSOoLy51hELxGZsyYYWTKy
5IyoCyBTrHgEOK9GAovyB1/yg3Nz+PLgQgEO9GqgTWZYHwEz2Rpta9ENDKBK9iVGaP81hZn3DJr+
hB4SUhDUdTnpC6oWsE16mDQDZQSYBPE7NwXVgLw7YyKMlbL2UCdpVo4pXsd8FFu/8vdG6TzxwT7q
931ir3xbkrFXTODcBh40Kd7oM7IF8gZX+KFkiAM2SWXY7v+x6cZx4aK7Cc9xw4Kozco8Kr8dyltL
Rg2Cj0AjC+qXTV5q2X6hM52RbadQ6B8XdwNa1RpgNL8jPaVepn8aJMvZACK9yOig4HVyokpwdGLz
xeoaXp69VftS6Rxr2VYOfwQWcXf8++fTKu94z+NqS+p9HPMmbUvE0JkgxynFyJO1GKGaurYcgUKZ
DKm/033RSVDHNHpBqArPopfmq+/MdzaGBZyEL+iXZyVZsThHMOoJ3BOl1EbLjftvWDgShGa+Mv5l
dJr8n1V9ZzfXorum0lZ2F5Zd3hu+ywQwNB4HHepy9FN++eYPClTu5LiWN2TNfhaK3Z/eDbxfxNfc
j5rmOWGYfneafSoqhIsIeQ0CrynXZJE4xs85vB/XY80dyHiV+fLyz6InEiukW96iPr9PGIEj1REf
oFMBj9dlewOl3cfxxXtr1ssRzb0afC1VKJXlJ+CC4nLkTdRtgygEXbFtxqEfykzR5NDIAJB18vdy
UMeDnzj9lZYx2Ks92CR7m8gGyhovFn6oCaFADd0A+z43SicdbOxSklQEIbaWWDK5xwR+1AQfORZc
YEiOrIisNCr4+zdmWZk4EAveoeHB1f0mR9FcU5/5HNlESsdDZrwuWhNyPNkr5zzA3pjdb50FEGjn
A54yjJmYIDFlfgVilFv+9PBBJs3Q9lZ6cGGYdGsEUIg7xK6PFR171VQg9cYwGFgIiBfodLSMjoQ+
ADmj1+lUx5Awyyo60nspTrA7bcc1X7ElQXDxiz2ZWeGW/RqBdhJACXjeXSmQfsK949hmbDafX6R2
WSihdVqpW10x1CT2r3YumMccn+Nv8z86SbaK71x/vh14qLOHjFOS6pFM0sYXe3U9s/e6kW3FRIOM
9XLLrLRnbhRI0obkLm69Lz9leRN/ZAic5CParW06YDV+45AhqG5tt0EgAh3rGr8vyMUDbMkpmAuX
vXmdTocsxF3pOWmvrRt9gXoFPnVMwJFtI3YRtt+FCNsR6/1UAtfnr40nVLhLLYENHqCPV7JL1S42
o5mIcEGnWhxck0YyAEbzOeCNKJpVNEnQ1jDRHx/jC2LZwAAS+89v5GY3f07LbHg/TE2F/jEC+6R0
JDTneWjSD4iIW4TtuMpbxwCyuqIkrJDe1Bkq9w9giFvpQnSRPGjmyCrxjcJI35KtYO5RBhK0fdkT
krw8NUs4agpS1o7iDySsohsrKHAibjcabXXeiPKE03S/7FtMk+UD6TCWgsBiNQh8pvPkwFCobywB
CvC05NnBld7QnJLMDqrRfNIGmbi09gWXgt0zhRG7szcbQ0cNgK0gjAz0UfYaGE4Y1DPXYz6HI4P7
KJ9bkIs4MUUzZpUwu4R+T3QjXm2QIKVT/5xstBd0gtZ1DhTC/11VjlETdqIK24s3bziPVir9PDT9
ECMiPdxWNa66Wj0Tf2BlZXWo2nO6OkQr9yasH4p7wsj9PW3b3FW+2Y/HJyybQTFwADSTJeNkBzor
2jGOWkV+obNA8ei+/7TNd6LM7N4OXz9s0m46EnqUDj6fg+HjmS13dtNA2A7s23vDWsSKdt2RlIQF
Dh1bukmp+CW7WQrlAzB/EMWETRoQuaUyb0B1NQQTJopAaCDCDZuWTPZLy3j3CsZyP0FVCVWaZXw7
Jaw/9jlkIVzuk56lmnZW+u6f2UQuBPfWVX1lgrJ9Cc/5xj0l9/Yen10QsbaEJxZ0IlP3yiK1GL/h
fRhsi+573BCRqXv0ugh8hQB9HGMtDeFV2rqoB3CNonj/tsGEOVXYwUdnTu8OAbRrtYeFAGMGC2QH
KPz1hlMrSEbGXO3NYqtIfcWI0iQ1LxpPi6vWHcsrpJWE/aSJYr/J68TAeEIAJ75Ggyx871xpduSL
flvgBQtPNlTjLEMdMEO4+7YhB6Lr1b6mnKJrDzkWITY83eX38DUbNc25RWk6ZufvgQvK0vAAT6vX
fz8NB5ya3Qjr7VVoypMjCH3CzcHUaGGOK4ajakcyK6u8z5A3sfCx2Qf+46VB6nyG+KZGwzh0QVNX
zoPNQ0gPX8xnbGTvWGSYIl12q23LJVmkU6aaY4JtI90oaBa8TpRiW9Xuml7Z9upM68k4h84zBiMa
rDGds84VK/1bSwG9edstwimAgen/G8d3CSw+cjfk2OqCMg/SukyOFAIo1PeH40LJ0qEYUix1jpks
eSFatLk/LscTVFbaCG/ayr6qGRQt4DcAkP1mve6WZjzWw31cmBOtmYLkcb+K2O4d8i/a6mTGUYyQ
qvi2/qY7ixP94P4mXi+XTXIx90RuJRfDs19qbtU3tYQxFMV/BmTXnYvgtNL682nw8lrC6+ws5Kbh
lrM8s7G8Hg0T4NcllhziGXkmlfV2HKho3oBQATG/UhSv8GZ4G4UuUqZ4Gz6FZDNVE6v+nZxhnCUl
fkTs/YXo0xOJOJlkiVEYP8u1HTGeZ1GQ8YWhVo+3MUDRZPw2qLdhAU6MyVXYpYiC6v4xbpEJO0IH
yB0HNxLgS61rb1FvQIkTWplboZgEE7xwa9jvpwySWea1Qj1LzObR8od6Db2c6Spyk9mC0czPDz1w
MZdAMnAj/Q7PBf7sK0qmEiWAmNrj7IHiJgYaJ9RFQTtVLp1jUI2vQNP+vl4FCQx3FPfLMAMtOYJt
XsLftwY8cruFwJGfUQQzMrysk+/ctcOsfo58DhQ8r64vEuk58ldldNRfmxwqbDsmbIIxctsU+7DZ
Jzy+KIdbTmm0mIPw9Onuc0peL9zh5E7Gvnrdh7qUy9ZYs2HHHvN7+kb21DXJJYh5pda0oMM6RyI5
le8OmqDvxojXUtBx6uCMzZkCPOdDqjlqVBMTp+LFjza2GCH9XzgIXy6M4Yr9GJBLIhQK7qJm5zf/
d8sSYim3+vCUvkeujvrepcKw5g66TUbXbohvPSL+xR5eVq5oh/osg5fbT/OTKq1x5OG1Kv9LXVZ0
4LKPqLJE9WR8vIVuOlhq/OkPcsbZOky6XsYu3OSmhUsgrPGPyZx1es/Co6gYVXu1DHfLer4/3aiM
/AiAcVqotAVZSvdOV4cHrCWTiq0iUwivHicb1REavZ9Ske9//0yqJ6LL7gU9/JNJU0hPhiu6Z0j0
wm4yrO9+9ylyatoS1X/gUX80lr8M1rax0FP34R9dGLvGnOSO6RrwNbSSBuC8sIoRWmILSg3aKqCL
eobHyLd+D4BS/blhHVu8SZCk2dTKH+iuiEELG5RoMNWjp/bvg1BozfFTcf/VdTx9m/eXXEOyhf8A
towE8i1oO4hCtCTsmSxfLikc+bkIoZJDVfYqR3vBV5Dm2b2SjtDpNfFfiq4AwyaX7k0+XfPxjnWs
A62Q137fMUUFETf4X13XcHdzhXlWTZ9JSewjvFJ3j7b8PH/j2Vg+lVe1gi4MeRHOJwaOm2yEwCVp
H2OvXAvwj+EIYFnSc+SkP9xlKc/SyWRM+8O9Ei4mIaFAv9t5+qSZeMD2k5IsfzhaTvjaHdM30PM5
s8TTMXDQt/dZu2hnCOauA9TS6arkrIutdWKfwHRpu3N60UXvqMsF+4RpG3hLUCJGneLbfxQf5muB
PVfLc36ikIm/cb/shXBxsMdSkuGe/7s0psGIvAI738IW5F6AZQCbsX6e3knM0vGLdm7uIffy0dnT
Maf4l6urdBuldRPHRW+QoomhvbG34dgx71XyyksJROhORB+G6ensG1KjmfbJCLnNwtf+hPVFnh14
t8o7Ac25B4KznlWVP+YK4JJw3GPurgDMW3H1Y+WKa6TOGGuyEv/k7ojtBmaf/+2U1ju7vZH6I3fe
ET72pniNSHw6+mRedZAsyrzmM748zaEwE0Pz40Gwm8iIW5Ixr1roBFTte7be1xwARcX10iH1Qxki
lLhYpAoxPDY7YpNuv0kPJlrdr35N04CsuTPEZiSu4YYrplyEmLz55l/KfLT8lk3lL9diqEyRaNqK
zKTG8+ldWAh1cEslfbtgkSIByfLB62OWGLYdYX35fUXOMwK7XB0qMBtSNyEQrCDoYeNMexwrlRkX
MAQUEHBJ+8rrFO5A8dCCXdkY+xgIBkN0BpzzdZBA70S7plVRQhaOZLpHJMSkKlPtKKGhF1skrxrP
O59ol1jM3xHtWRx+iIPrgyv4jRBqsk4oQJuJhUJlnQvZYSbZNAA0Fj+qf85EnHv714qGa4ok1RpE
/Re7xqxCZoZJBbo/EZD7rqdPIoRTjdFayEkQK6lrwyDGw1+irGEbRy8hYde121AqvKmdwjsNYNQu
ohsWax6SQoXdVqcaH5ftltaWcmCRwf+CHye1E6N6A9xZKxgkSHhA0hTWFGG9/BlnjOGwhEWaHpCh
ahUm8eIJXOY50JYhhhg4Ir0Ccyai2zgFSLPskG/WjG7M6GNhME9m3s2/YKZh3scVbm4qrhYBpSOC
llLGAwIuHrMxvC/prwz453o5bPqGEfZ2vXkJaRh+7m+twKbd0MhRwPmBicoAT6OUr254D68KxwoF
JvaCFCIEm2YTw6RsZuFPwHzB7BkiWKxtr42wpJfk4u4RUbdSH7E4fLWAd2aBLiQBXdw2ahHoedAk
5JFV2uZV/YRtprdAGIJq/pCzZbwbi8EmHCmebQIGucnyFhlFVgt+Helw1s+NsSraiCD9l4dKGFDm
MXlvP9DRVqhmzDqAICkYm7RwwDJcz9XjcDiHGp/8E2CCWej8gUW17sQiC+/3fhblT8cPxkr6R6oG
VTGeW2tUqterP712FrbC6mLOm7NTbSsDM9iCV7Tf6HygPNZNFw3RKrKAirWpZa/siMhboDEn4wrD
UacnI8S7u27i1wKGdn7uGNZiM4tIjFIQoP7DnYB2+EC0uEEiTLp+NZGxXOYOMmL46ToZ+UaZbft1
B3xa+8NesS/jfNlXKMH2T50WE/STmZwjNj7Die8hANP4CmhOg3JC0yqMP6UKRN2mwMjWVHCDKyHL
RETcn8iz5UG2I5opV48nCT3V4EDkb9sPqIFDmuNOghZLjxWR4HE2pifzxfWPieQsn6xbHQYnTu/l
LuoJ/WesZnnPHHuvTrAkdib317z8VYyY9aEF7nQtmjfzRw2SyQsjdRW4OGhdztxN/ANfGN82jPoL
lcpJ5Os1bA71zLaiSwumtb6eb4r344/+kK0cOlsJnZHzs+ZpXP2mFq6N68fAftCafVwfTCxY+Aph
YyKXFCJjseZ6sZyvYYKh7YXQbFbIk613prD91DCz3AME5LjWoGm9mXfYuzWKJigz8xx/aChkxcCs
/E7n7pEIi6j8/UljSqWkyh9QTucdqSWTpox1YHwEBWyKh7rMWmaB4s41W8BsleTrN9x+MDWeOEV+
FPiaJVOwPCM6ZuZoiP4rJuEQ1fXjvJq3m/vDM1+lzINCOjEi6IYabSAs4Y2YIL3PCzHdNhwLWidx
KfyGkqM41R2rY1tTgw0wTnjFmonU8iF4EN1QA/+1bpTkHz2qoXit+Qa3X7tUSD788TjeN5NLviWq
2EfM8Zi57iEFV/LmFf3QRHaLTDNo0xhzwdovW0Xgt1M9tgR21GmF5ALlUSeeqpVfPGIX/EKy3YPO
c8TtLUIZ1cJVAtpi5ah+5Mu2IMoF1avvv5XGldGC0lv3gRPk9vOjQqO9ujqmGjFgE9TZjPEs/Ucl
/UJFf2waJkw6Oc28pSmzwsePEejncBkPFtV2/aVoGiu2QKVr+I9ng3oun1s42EkCzJge1XSraEZn
gKCqInLVaCnGnewa+2483jM2b6HA9x1Yy29TUGOOwM/b/v0f6Xh9ljwG7/QFr4CmMTpPE8ojTXJq
otJKLZf3pyUm1np70EU2EdtLtI/Zb1Mc/CXuiIeX4sqPInYYT3UGFXcy6p5bi6rX62+f1nCtcaAN
yCQI2nUP7OmtAV27gh5DyC03dU+0Hl8bSr6dtTNqJnrgbabpwLKl1hP4A/tvBMBH7DG6unZZHHY4
hGUx777nS5A5P11nvXuNVec4i45R6K90QN5g3NOVCMS7sc+R49993HNElZ+iNcpSwaMQYC6mdA33
faZvQwouuCCL/BfzicmvU+2DTq1q+It9bwfRLcfK0bbdgAfjQbjpCN0S6GNbnnuuYVm7aRseXx3z
7/53ZDhDRsjMYtLPRN0A3DRnv4y9AlaEC/l/Jcuo4xn9G6JLvxdmYeVkDWqB8WWaHIxTMWQLJCA5
7n+lR1h5+M6aIQOcXzPuDfEy7HIlvdvFckcbmqkNI3MG0rEM2BdA9IjWT0i4AaGhzBrGFzTKeAGO
RgvHm0Gm20bcUpekn1B0JmuCSi06DT8Hw9OMJpfvFNkJ50Wbas+qG36Xvo1bdvjLoGPlncz0X7o6
hVqwTXGE08eaG5zebUz5LjxTflZtO1dGLaOksQi6LelbVeBaE9KvgVK/jZ5lxZov7SiYre5Pp2+3
D2XEhjvZ3xz9NZQ+43XcqUrUCw0BpWBQj1RnlwtVdTgagCFqXVLsfyegUUeXShrs8CjSWYa57kF0
LYX/N9VvI6maAiBytMk24rLPCjOmHVLy+FaynijtMypT8kjxag2Cie8+OzNl0U+rv29mS9RuAPPF
I7mWJiCILsbe2I4OLpV6C9rm1W6AlDYvQftUnBlRYYb5cXUlwPajzMd0Sl7NFUFJbz0i2itU+SJo
7B+EfiypL/8/iVIp4aiG4tMojU3TM1Wuw3fxCjS6biAbwyvNRWXxIs4hQYBUqKao1IgPVX4JJyjL
A2qvvSu4/snj5bki6KpFyzFu9by3mcvhOw2gADK5FTmVqy9p5EQYNV23+GFMiW0j2JPkRVQkdfIf
ejn5JQN4lWsYOz1i5RMe5PZ97n2HtvV9iL44geDbGc/n221l8vpnNO3crfDC060HD6/lgWFVM5n7
jk2KQYCcwqKnVBcckLuiHIDzetjggC62daM5mXs7pkbCtlCZWebdvkuifRVIGMdblYeT63HOXvlY
fyBQBRlEl/e+1jd0003xyh0HcTDi1CSQJTJzI7fuAEWljtYUxDaYwXIGJxkxNNb4yKVZUc+Dn48E
gPc8X5sSjcIrgPubEFCFvX+RtAY/dhJsvNefuuI42cXb1EMpgB3XnBFXwO7okEI0Tnn8Ulz/RIob
sCz0SL8mdqPkg5pj3KpQP8C8DKP5qXUCNnjBYkH1mT2KkK7AnjHKL+EOjf0I4kkw9YZf19oZr8WC
LOlXd6hvigtmMooOGK3N/uuIhB1u6sXg+o1qic0tNqys/ZNHIjfCFWEGCq9bLzzvAh+EvB4Tu/mi
JUgFIkeIdUaTl5Vobj0G6e72Ex7aUF5toujYsL6J82M0CC6NQjdEJQx36xWfO+RDGY5PuhPtS402
RER24nKJMbKt4hpKha/E6NZ5QTAyzVRL+ynMTnevtyUQ7dGo2UoiLdZb35lOoNCoPkeqq7+Z9ads
kliJFHbHUUgc57W5Jmevq0xd4h0G4kpeJ6nrxjn+lsdEHG1lwYufEIJmFRsNiCTsUe0UFy/JwQTK
19lqtOzxAeg5nZZSbKRSNaBtgYbKgALIimXO+LvvfyojmKYCmWxxB2Yh7l3z0UV5AbB31UOY8Bdl
/WeqEPAHRs3IYipfoZSE7lyIU21P4Pu8tJGplHN7pIm2D2NsNtGtX7WehtPZ8DlcyCkZWzikX4Lp
3z7jWwg3YaBuixWFeK+CTPvEyQ1U6dD2DI5HAmXmR+TtNZHGHskX/55NnsHyG5/at+UV02WDhZoy
IpcP401bq7EE9UGCTfVIFHuJjKerxjrmrR05BVO3e8R9YjFKrw3ZAF5oJiiY6yFplUcv0mQV4TPK
KwFGOy/nJ/Yv4gyRVgADckeLL7Ggj9pHHi+jhjVQZY8pIp239AXZlGo5XzonyiLv3Xq+TUqLaZd9
KyIoBkPJe/PMbhB7+N9KhCBhWIf23nLApLCLE5BZkRyyRPyBJALAw5PO3DiYKyqQnG3h4zsdSi5n
7BHvdOHA0IEq7Eu91a7cXXtWBjc/mSIIjXzSnGWDWDnBnJvFw3AD1Equ+Xys6sCZLY1CPapz+LkU
nh0/Di1qRKjMFTg/2Lp9UoAFFdvifPLSwejMTqeAPGJNr9AMN3Ba3uSuyrrTq1VB9wmXqFBe0s/f
G5wVuoEi6U8uzujH++y0ELGDXtTxt+Lo8nh/gaqfLDikuzalbILGPNLJxFFRvx3qhrVFA4EjITa/
Qibjq0vhoSk0VN7YNLc7votTnV7UIy01trxUvTm8E36R5de1t80+64Zi/WTews4qyJKXzu1tnmwg
ZfEFVIkoNemTkEkcdUW10LYv2gBRNctxkjgd9AQRbl6Pvmcft8GrM8RKSfHzDHW24zbOp6hY20Qf
fO2kkqdVxqcE2GWjk7Cu9sYb6QeDTkhRvsEVaXqJFsKYqoluCbFDM04JRp6vcjDhg+RE4jq/uys3
uEAnzAZaZ3K3emqmkhAH7MaNkha20I+/hnaiaPRhvrUkpG4xZtxurC0u0AgwFC6S1/ztTqODKZh1
qMCbPtHHPkpeHYLz+X76EhK8jaLmBOBGCGSF1By4JB4lCu/Ag44lkFJaM0hFJ5B25UoeirsxD78N
5yZhLN0JFzkFvsGwwGJEwGbS8oUv56JaZ+KVhyerFF2ooCarU5pkLpmZAs3vqEaWuU5k8AjMPc+/
oagBTJsxvOPc7+fX20nvPG+jwnJ/ZY74ShIxQIHZbkbY2y0Ryjq0SRrCrqDcK+FKLK0phtUh1WVn
oSucNL+7lhGAxVJDyVLPl1/QUQ8/EFidVXQJ23YvNLNYs3vpI4ENW94/GpjLLeZuNsgTjWdtNBlA
xk9mxl0y5k8Z5UDG5gmld9hRaZsf/zydxNvm7Cz3JPKz3yGLOUR8fQwDtFzNhRtKcH2d/wOIqyGe
WxtfLgvMsi5XHHtCZx6VQPXiG0IFEjqF4hiQhBJ0GOxud+bFOzrSn4xPOsqVdpEeQ9EuOa2lZgd3
3FPmnE1suWJ9pybyS34DCa2nPaodH12pAIJQUEiaqKvdHRxQOsx8ft7OvEPURA9W00zBQvEPDEic
QGfcfYuYygKVqvTCGrQ+PGrPt3yBJmjc2wlTDpFbFvSppvO+lAwKVlGl7qULgMJLvc8atQTEAUYM
FUCUdCSImVyvJsLpok15eot0wBEY8xPDx55lxQo/XYNtHIihJ4Su7t01kWPjevFhLYTEjtuI919s
oFRFUJLMJfZZQyuzdYT+k4NRHSXN3eqaQGBZFmSh37fvs5rdRppnPU8YNvG6mvGnU7+tKhX15oIo
8IE5w60Q2RVvjaNaCVD41/vdebs/iA5IvUL+dbhsM3i2dFD223CgomP9f1jlnino0LUFrEDbIh93
uf2QXaCnybwhgRDkn6v/V+tmpIaRF1ifDE4Lq+u7dq2jRS2m8eaAg2e2vESH5HPticS+UzS6Da2p
HYVFtRNumJEJBuc3mMsk0W2Ut3HRXTqXajZEdEpNhvNVxiH2dXKQCnm6xjjEud60Csj1QbxRVCiY
apT7NSEWAclMJ3gIJy1WSQIGiFbYfSE8MMP6fbCaf0m6ww+O1oPAFpSG4FkovnV8F2NPzZKAiNqJ
4DXmz5XUs4+I7je3z/2VEBvdl9sTnrgv31i/h1ClA+l2ikesat+CTjSgXIHwnyBL1LfsGBC7QYKM
kMTspff9vQrBQ+Es2ppNFe4aCbpWVgy1/dbrBtGqSJLFUh+9+8V9Dn5nGZcEIKbM9xqxEwo+0qQ5
sNHGXo3MLw8UUtsNo3Z4fIPlUbY/XUwcpdCyKuMFWEifE+jnaiWme8o7prTUGUNGiTgSzB9+xvZB
MRiIn1AQuVjvZVKVr9XaDnN0z+be85jL+r7E/o3vyJav3Rj6pk/LEWf1CF7+0L0E/fFTbMQExrkz
HEyb9LDkQ5hf5mfawNRxubKWt7KXjuuxwKj7zFDCGsPaCoPwPBUbEBUBdAE3xd1oJww979iChMwo
RFHL1T8FiSPusv6V+I1DY0ZdjXLsjKGSyiHvnytPDa+UnK//ZQrnbTcN/fAiLuKXVCGtA3zzpqzk
ZR5Dz4mHnKCV0t67Gvc5BBSjHoaht9VxEQFVVWhNun7LOTqf7gcZ7XGniTBElexLEs0BQxGNS1xM
hedQjny8LlOat+Emdr+SI0lCL2/whIFghsJ7yAd3N7vdaVi0wdtArnDQaiDwky56siZkLC//CDfO
A+LwpJWp8KYxGMK5MChFUlbLm0frPkTPZSFjufvGCHsyCSmyYds1WTLkQtbA73EhE0g4LkNgcmpe
dbNyrOjiPaMD2k0NGNSviAoozIRUJEQBUh/sWnA7DzYtNSIKstGFgT+Mr5wFGw92extZIRDu/SbS
/6HbO2oZPVxq0fAhqlxEgMxdY9ZpaHJ0QOk2NceIoqMiQsfcdb5e1VWBDugVdBWfHnL/rk0DpLjz
2xslB0zcvzoiYPqbYfhA+Flk5SgLx/dL33KsuS62Pvzfs2Ki3geBy0KjvmYV1tznHSOULNrI82VY
FakAn0Iil3Fed0OVnyf9d9/YlsiYyFDRsI/M/UmXkvIBZXz3Ig+A5sm9SJTEQy+Nnjb3qBtDRfeM
FK6Sh/5XC2vjEwsAgzGkGMZTyDPcdQ1BkcpVJJcBtH6uBrcDQIO+RxltMQsbikk+/DkR8zRPo9Mv
bmePIGeDp1Hj4Lh/PnFWN8SZvbn9vkUOoOpTLEP5Fg3Lz6+5Z7W8gdYupjdzUpv6/0D/rfBdtBDz
PwmHoh00j3upcy76XHtSFVijtC0JsSYNYtFk7vQ6FMmeTJFsOkQiSWZvNJPrd7G9ulb4AffKOHvo
t12qM9ELlP+xq2DHgMNjtVUWW6WTg3xiE3yq5Q+tdKRptpMK7pwHL5DItNqr35aF+JcrF+q+Cqtb
z9M7N+1vR1zf6w6/mMQ4ACLEFAp1yY07vHB4lG79gynSoP7Y9Z1I+AxT4zsuVHKdrcllbcxvzLf9
K7qZeIK+he2vKIb8ei9ZapBsl/xkGwGwLQOFM+mmLOj5SgLC3mXTIOuStNrY+3e18QaDdclfcoPk
Mb3c+pvs7lM8MIwy25F42vV8lhqDnmVWlcxO5wFjpiGYHYmaE2ymvad9YcHpVSFnI4OBdcVJI5B3
RPWdD96O1czTa27zFga7jPUZRu1NB+AVMg5uLk9cxeNYc5eMr8YlQhvjPRl6WQlsIzbOOjqwNxRZ
MJPliI3tHsjKam7ceDDrBatltdP7hU1Cekx71d4B3p8tCyAKYtBAN8OBrep/rEdqwh/nTWUn+lYx
fKryL/QqZNQgbVWNrai2EVwzKjSMKSBCRuWbOIqKePRX3tZYJRy2rOl4E56VhiQw/tmCkLvfotn8
OrqZp9c8x1vqousNyLn0fDKPkVN0bv5Ezl4tYNIKCl3O4f7Shcmftv1rhTURhxW1p/SRd7ir0kz8
TTF4OGeW9LFxRIJA1/BI0sa7IR6sLJrLtZ4ydd2o6QD54UyQ7Rj4hBiTTYgXfEuB8lO7dqoOwMrZ
gcJ3pzrEcYRzsGHiRbJ3R26VHV9X1sYc30sDAHKoUmEzJE3BJrr2Oc72+mRBtaax6Fuj89fm+3CS
vXW3R0UNSqWErIjbJ7JNFYDmHh7GO6pAgCOClt4XQSGmkukAIuMAljMOjtsn9hLI4VH7YrBe1KOJ
6yhF1TU219gceobCNrqUvH9LaTleypcXE8J272fVPzxEcGb7GUMnhzbVzuLhSlbEY09Ik6XXg/Za
Xe4t6inyY8JNqyAZunML8w2r8IOnJCgQHcnO9aVSsRWmc2f08P2NJswvfDmdxddyLEL9Nfafl/tK
18i/SM79kaKt/1XLoGJWMNb+ex4M84f8nGiEKG9s1+OzjN3L2fNRtnGwdsscd/zcT/F7dDdCPrDD
ahrhZkKNIdDQRyDj8MwTb3LHw0dJuEEVXZLJb40wBYR6E02Vmwj0Ia778o3d4Unmb/OUYWwdeMzH
QaMka+7DPKM/BieF2TKNOCT87u9mtumsXEf3W+DJivalAnNQGjJEtLCvwiZthH2iT4hxEtBX2Unr
NDxZ0HL1QV/2gsDrK2fJPLmtorJybVnVkWGD8H0h+FBuocz3NDoLE6IQaSIw/CCsf/wqYLg3BseQ
LBN8FqjSyctGfRf/cUqzx1IKFgeHpqGNxlXap8VOijRbCzEtw11K6FZwcZ6+ibihT9s4HoXOYw50
NiESygACuJdeJ7+v8vw3nfKamhUzag2/MYxP5DQe75r33Z9O9b4/8v+psITUtwd9G5GZ++ePpWZ6
VJ/ZIw+jVy3pNa1u5yx75GbrtDnr252GF+4CNvmgIELro3DuqU7A0ok6w3puAluYcJEW5SwoEKRi
p7tVMMIWrxt/FHtX0Z/fpd4jm9vzINbhOiBa/ujryBwPiC3lCVzY/HnRmxaCBbMmieR0gzqjIKBe
Ewp+5jSxe6aoNGgo3aC80k12Ua/Fy3tv/jukAfQv+IfZ+GIm0EGwndVPWMkEpb0qlwVdIfwT27hD
VPXlRM04gU0q0zARzIvfHwns74rUR12mti9OewBkxqBjuL7UuYIDuzccqtOTSJEaclHixZG2uG6W
6YyhoP+cEgYqeD3ADfk7QQ3f3kMjJ2Rtb1ZlbdGSl22M1v0u0u9tG6fwGgmZPCQr/fVHODspj87z
g2B3hsnfiKej4zp2Uqja74Tv6LTIT8ZW2qyqIRU9GFt0BaZ0AE2498V0Acjvf0WQ5IyANO+2frVN
KnGOJb7ifv/SiEQVLRc+9GC/l5jB6UtA9jPZNETmU+A7BHFQucG/iB793fFXSP9wGK2YH5nk6xYM
km+RwPqaFmGdFPBd+XVMnWPRFv+vJwB3BcGDbr8RNNbRgIJePj89feKB5C9U+2wFPqnYEYX2N8gj
9GmbNdNNnX5mcRt6Q1gSoEDovZUdNGbSbByntXrPt487qP6Xa1ln78wMP5Ykym+3FqmqhUn8Ghq9
1auBgieLhGzDHeTN5HMpWxjYnFYpzo1IVVzA9xyEd9+cF0vznBy0gVdWiez/Qhzc608Hdrcjcfv3
bxbxBBcDNDI4VjV8kBy8Ep3Aezn/304paYpSRxY14sDBSissosyFKt6Btc6TltkA43XaruuWolAZ
PL/ismB7kOqzx8Sl5e6Wonl+aqo8fLxPgiZMHrYAxL368QnmS5sOWUkRhBUdSVe1NltLVOKo6+Il
peyPmR5IB0BfmIK9of0k1BhCvC21LeX+rZyPeViabsVzbiZPTu8NhDcxl3n37vwrEogNKTmhy3dP
Aaq/EqY9HLYfSnyI6DcV4IWUs6oJQN3PDYrVlxPyn2UkRsKpDWWPFWr5U20tNaF4ZdmISX4/49Dn
cGFnmMdg2VN5uoQI4v/dLlOKh+rkdv5GybxkRGOWm3tnhAsmVcqi4BV6Ahk2u8911LM98ubvXlos
Dm/If3LQdEOCyp2erh0OfpVlRuB+nSP6z+fRLI6JdkW2znWD+Zhh/4ijSRsbw3FIj8aK4b7WUvte
HKYVSD4XJpCBsQcOLrEfwyg7jV+ovjCgcSB2OO8aIx0+O/qqd3CVVSN/jmRZ0r6AHUfDvkdb/y2q
bJZjeMordWZ03u8o0ZCUAo2yiC2BpuT8Av4F4DTvp+HruWlIPpBtCSbhRlzNOKAGtl6sgXb718JD
/tOVqhwp8i6Y7TykEsj1co0MmwJE2JrpC8TOq6n7Udjhp0fYACtjpAG4S0r5ROLB67cgHrqV3Z0m
z0WymBc9gxqb+oaALg63j4fK7lSVjm7iSU8bduS+2MipysojAPAwu/n0c/zCl6bom0mJMsn2Z/qz
KEESoAgRbaAU8sgwarwqJ2bXL4uv6YJR2/BKw1jIsQDewvxyW0M0DitdyNVr3Sr4Dj3QQAhpZRTR
AZYFJyLXlY/bUnkI+Gd9tQ+xPn8FvKYA9gNKNssB/W0A8LNI0p2zH4ivb6IRvpjt1633dpM5uFRC
FgVtYaDcVwJKTsy9gDpAneVvLH1MAfIFrda91CXdXJ5qRMhHjAkqsbn4V806gCXF9B8XeRu14tuY
Nu+Zcw0nR8GlH6ZtcKDxJobtic31GbNOCSQPophWDop5PDXM7bT89oraK88tUhQsBFXqdayU+psJ
tdZejqzYYLa2iGuaCflymqm95DFAG1WLE2WQUtq0qPLkhWOVkjqhByOXULdJXD7Ds72wJH4+57f2
xOAwzwjd+PW0fNQl3/bgTqCfR2QNtL4QmNM694iqG6g69y3I8pn9cFWr3JBmdH+0j1RHH3/FpulV
DS/+G7/MI11IYPYESF96/xmIDcscQQ3KUumIALqdVFhitCCV8gQWM3INj9sPgoiKWZBdYwbSWjZ5
Bpo/T6N24aI5wxZsR9XnZnt6eWxBrtYz99Oini0RPiY3N5TTVugZwzJ/ry9j02WX+w+ly1hQZpzx
hyXv610k5bzXCW28N+pFOOkPetJmj6I1UxQ3o+5SKh1W46ChID7/ZPXM22KD0vqPWCR2Vrg44d6b
vy8GDKKgZwsELsNo8VPiJr5mJqKz5FEJn7XyxWwvgVw5+heYjrU9psxcriQPKvhrNnbcLBq+/Gze
tRuSkxzewXg222XXm/NHYSEvNCsMPbDyBLIA5pIVLtoQYdKiBArH0TNtVUSOYp8Fla5H6wSUWkv3
QF+On0SXX0QS9BYdcvk2OJRW7D22Y7o3ef5ctCsIg7cfKKFdGKvtSIL+e2+dOfOLPQfEJYHJgryv
v0lTOGkpzhbAqxwlCWdu2W7IQfkrE4Jd3qhWgc7eSi59bN69U4VmDmULEQjS54uigIlM3UsuLQMc
scTpZihS+KdE8KEH5Y0kklZoEVB9peB1uJFlXOsdrifSpWlUm63kNZclIJOci/WcNMPZjDdRiHdc
/BuxfITvrXTDSL6IYaAv73+Pnc+zkxLxWJUl+3a/tRNtwzTyNZA3vMJRAWwatgNlnrBR1vCU9IYq
7eG+ORFsh6j6ullEEK2DeAkje4r1Z7gclHKG3hgi5+LTUsM4hXHKis8Lr24MQzPFTap7BTLmDgFp
376U1+23Q1lAYb5Z9t9RwccK2ShmpOLnqiqIGdfQuaqFxzE27nA8c1vUIw+2tkE4Jbt5G0x1ws92
m/q+GqvBfMGs/0Vjy4s39MndpyWwgyYbUhbcB2Zcc8uNPY7WbRX9adsAk2AfOjVxNNG5fHvjg8bR
+0+e9e6sV5tlNibWn3gO86F5EcXhQKSbZBnCnCX9WGfSaGoloEthA8ns9C+aiRWhIdSyKv43e/VY
dib2Pe7mKwywzaOKBSxOFT8iD8ZQBb6FC+voVRpR7OzSEKGeDTBLYjbd6M8HQXT7mNCogpjlER2C
hPSYvRJSI6zMQP7M0TFvwHUUD8OpQ3Hekt5LFDrracljk5yQ4QsQG8aeUzIuS7URQjcBRBog2Jn3
gh4h5DPbOmsd0nRz7J1aAvvpdYFloj//HAdkW/UCWydeIqgHdOw7I6wO8wN4C4a/GaL7VnviQSoH
EnGVPur4Dr505gCaCFE6VcQUcX9M6TrP0HcVaCSQs5IoitOYD8vV3bySv/1kyzA5LpuiDk78t2am
Yy/RWsfiOCz+f0evRhfEpoAE/XFmBmzHr/Pi9w+K2eqBdve+B091fbPP0lJkS2poJ/5YgOBQMUWc
XJ0cLBls6YnCSpBXc8ZbChbEu8nu9SJgMHjY6w59/8/EO3JNI1i0vXhwsgStH03cxt49G/FPNGIk
C5826XwWJauYZ5Vhw2SogHBRqe4R9Rgm1a/zIqASz+6Fex6EU9LPpMQNDIytiCv4gi3dysvCaRmD
cM8HCD/fWZ7u+/MsN/5sxK1fGIAsCSquk2GvpIv8TAyCehr2NNtCscSbE3CTfAEffirjh3YTvA/I
uREjzFjvcEgaI851q121Icj7y7pxT4NjHy9PjMEZ7yTqTGsS8CPwr0zPbCjDCDDSlPg4c/TxQcmn
e2fGD+UtC7Un9UySNehRdff7jRcM44WsolQsm5rFH80e1rQQ5Vk2QGtClh//xOdlXgzL6gmpXUsj
Fs+Ku+elOq1r8Q0MW1muapevo8l4oCCL4vRrDJw6CW7vDHa3IdxHT3Q9tk56+Knjk5gMQ98meiHf
z9EDI1LoInqRki47zbMdPfYke6/W7Ar/0mTy4dRsJlB1VjWfMYYcQo3Wv9GhXy4QTXkUi9d3wR+S
uvF8Ji3YJ6Y24Y3KMndtW69zNu/VRD1Wqq1b0bnJu0FDtqL+/sYxWIoH8ZNKe6YYBR9xYY7wyK7E
nhRgnXlgQ7K4+yAKQwOvL1TfTrza6sl8PstB4XTQ0Vf4iLqLrbmvvlANjUfX/TL/bUq+xcWpCd9s
sp28o4um7UH8kCFtT7V7gvvoQ+VtCJnONvpMK1o2hZhG4OAS/KCUZXXQ+FLrNEAPvsIAL5B9PTPP
fuUuOa7R4uP15mJsH5iw5i9iJ7y6TneU85UUyHIGnOyl/Pcsu12i6pJaMjRKi09nV9GvMoCpUnDN
P8p9jy/y3Mp1MSV1mdN49QLbib+/5vqlZo5pDFCYCCvCU88fWMmlJHCCTMM3R9x9u5SYlVwgvzbf
KeLBIe6Pxk/Z0l4tfSYSaECJRsaXRYXrPYxn4xcGtpgUbYetj4o/YK5xkRRK4+QsoHcZmAJSgkbE
w/cE/D8OZJjqbuE5m+dqAuq/rkB7YXzu81OiUQMmD4k5ugF7jqedEPdf/QSlg0AHP2lWVZ2LN8ez
5NAutJ0+WW2PFbtC0Qvp4lxlfcF9lkRQOInVC6sHetNLyX0ouqjCXvXoMEW+zJrpevdyvj1Qyzun
h9J5dm8ufEPgyNxnnfeFfTwCztiD+5TaUuDfo5BCSMbt6cYZwKcdcIMtI2HmXDdS1Qk7pzt+VW3h
MMqSPeb+3RJkEsnY0zyw+Aajjy3G51Vv87GVgpNI2Yc+IQDG3Szugns+4GSQAyXuHCPrSh+ChliU
s47Hcjo8LO500fIgm51k/fYdb2jjz10WixVTHuqBA5mX5U9XUJzBd3L9+wIbwI3PYVF9ysCyM5l7
PQDCAtRsgmwWxvuh8HRY6BERpWIKITFD0hdFORw+DSZnWf7JPx86uysHK/55UewVN9lKT38KCtG1
cUgVSb79dfiV4MttIOCktYmQpvH0qDxBlyesGPClJP1AGhWCLc/iv3umy0XMr7S901VRwckdRjmK
wbQCYRCoD/9dfmpAmF8F7+UbGxI+KGAPRPkB7vBiVhTn+ceC7j5pWJ3bhTZ7GaPhp8xacQdMayAs
FfcRmTGxr3bq0BkKlrgnjjRy8/366UPTg3yuh7TydppljIF9K7jP2Zj3w1Pow8jYDWS/ab/G+18S
eDxbz3vVwdvhLJ+kAslXJ/WMuEiTwi+BvdFFUeWnxtekMhjpVOgNWaE9QWAOYDai1SGabfCFi1DY
QeTpX197pfsVPFSIwEU8Tf1gmud/uEqqf4qC6y+i6oJqvHdMZM76sLIRKlXv/SxMlYUlLpypUC0W
8qR3hcC5TCqfpboL4J04feieK1+iWYS3f3RwST5KjeITeDqhKJLWk8D4gk1lpFLYf3QtGRrksHxK
eK1AQH2hDxb6BL7o0iKto2hK60nRc2ZHGxQvgh5McqI5oLIeBzxRYrypcWl9yFzfsbTCTC9wHe8t
xYPzt/O473UrNGnOWjx0orCwoOJbYfkd0h6uiMc0oYuHnbyV4dEFztF7I/57aMSXEqrWlgc2iiDV
SMffY4Ca7Jsgl26i24KMuUVID+Po34nsibhxdGesqh/TEU0FzMAkMpbsP0yKC/NHLhCan3hniUlK
buJnryUjezKzp17hbmdczLuX9slZbMKuipoGxMmBpUvC46vA9ImFrzprXs1A1BWagfOGYI8mdT1s
jrtkCOA+56cJoKbmnC7lTiNM3WZqGFhd5j6cjwyrkWqb9ZlpZI5cZxyaX2xgiUKq+ckZjL71Sz6W
gf1XOIZkkO1uDowsFkEMcsPaOwljw3+dcCsfBqUxkN0l/HH14Soj/4XKLOChGlZkQRIm1IGZ46zB
J76kDJ0ztduV5YWKJcXL/IrDfTmK1JZTxjX2ao54Z4opZSE08L9tvg3iZsohYADPf8VAPh7lKeRg
iq3nIqSQbyOT9JvJ4mXkEABsNge+vIeU6P7MkuMkajRe0yCK9DlrbsOsuSdUyAUE4MFi2Cq2f94M
64Sp6IJWWljAgC1aVTN/XIWyGEIp4S3p/Fxaqp0BCGDZ0yzhQYRYgTSnfypBSUASO2Plaw0IGGpG
th1qtf75OCNvAqHLFSR48NawPklVERH4X/McVKS5CO6sfba/ZPd+j/7aEKJ29h2mAmuSY0b50Caw
/grUNbVJJL9cYHTSu0AenR/sHeZE6pS6HNUaZsW5ucBQi8DY8EMwNn8LisAuGMrgNAwgBn11NP2+
q8EWcjLkuEgJCsjW2y+l6xO25PVKsG25yFepi662YVXAHKdxL9tDALx7jCiBBb1cvCUkZQ1M/ZXh
8n9TSG/2syT5lwdIaAWuNmcJw3ZYc0UDt/6YncezphXiECtp8U6oo5nsdpABy6UFdXMsh3ZymyK7
M3iod/pYTFh+X/iBkMABugdpd2Zo6KBh3iXKRUtM6+OXCaEsTwjThhhMUPtq6RAyQeGJ2+h/qy8N
zx5TjrrgUFNzu/DY/2PS+FHBIAu5kSmzSYI6l9YpYBeY52mkLjGAIBkS2aYVEfbg7fIr3h5LuMhQ
TR3YKEZqkYKdqdb3JAMMtwD3NfqcmJD5SIbcKUZDhWxfSX/YXjgbD/O5yZb7b2d6ja/yB4KF/ogC
aekSLVg3oAniKG1TrdPHQ6pPLkuTDLJwSzLZqSVml/+0ajianu8UmiFGKML1AmWr/ptuDB3tKqH1
XNDHLG/bCjA6jikWfNC26LqJGGClKF7f6+FlfAR7Ve9nvplL/viJecLNOvQ1BDWjVGfhCMRH3Uk5
YaL3uz242qS2VuJsXypJjTHp7/d9+z7tRQD6yAiy/bNPhhnkIc7NbQ/A25lfNQSQbQq52jxf1F1Z
8tDqy+irgIt4wSAXXnAxCcuIYM+ovGY957NpIYDa7eO53buUdQfJ4BbGLmhhfa+gTiq8l3GxupCc
54ssebbLbq6kwX/FOp1GeVBCpz7w8R/TB5v0wfXW9+LC3hJHKQZC1LlGZJiWBGgYI/yS7FasnqqW
4b8FiFNSmpxwWUASifHbhDxo6hyqL5BZuXzqzFxgm87A9BV+Mak4KY3dQCpBOSGZlivWr3UlFsul
hUnEanVx4zj1xVEdE7beP9mb+n+w3qSGWzsb0nDhzT+Ys1bfuQ2kaDJ/rXA8i/PSYi+5OJrms6Gi
yz1xUUOOAEqUANHQjYJ31FFa3ko1xp2DzdP2pg/q7OH6RTMOEgAdZt511RG3Ij04MPUkycayMJIb
M2LYl67wUx4vMjm8QoGsSePHp1PKo6SL078uv9NuDnVRb9Dib2GP4EdkNTnZPRz/WtiKu1/azY8g
0/dnuEy4KlC8knO0o9dTJe+48G5CshRPM0N7MLIfu1j8as2kDNCk173mdz9ngA6QDlODtOly0DnX
mCcO0VyRZm9f92OJiT50rAPQg2nUBrqNQY7p0pf+5+CwrS1JOcBXs3V6W7XqXNoOSs516m0mqTHi
+BBEIcVi3eIyFoJKcorTZn8ql3j7aqaSwCJJy3C6sELRKPlWNwk2ENlFIZ6ODctgzO0rCCugbLHp
+n0MNsb2GbHgEJu1cw8W5kExIvzatwlh29BQng6e1z457xHK1g+A6h1IOB0L8hWGxaXOOzIUReDI
Nxt3cOEFLXbU1h/tLzNTNJORrPug0jFttgGku2q3bKw1H0F+txx2KfdBg2a1EtI3j/YKBJEJK9sb
nzhnAQax1vTp5hLqvfpjCS2PmL6zAsRMMmKMnWlVygZJ/zde/ng07DSS7VrtWWKJDNGEBrp8imFW
kxp0zjcQKYnVoeqzUgQXw38GFW9KTN2NR9EuyQ/vLpQD587KZbS2Hgw4oQxZFYuClR5i3kjEi/0D
h9c482IsTYHcBXMKp8OcmznV/9nPhyxBfHj8+to7GZtMrPUYX+3IBuAOdfkudOX4RV28cYv5N96P
mkKMEi0vyf97DghCnnd6gA9ZvxgeXTwbsl96pzP049YLzs9fo2BjSjF9HzSh9+lUF0spL7vLsIEN
aX0hKdKL8+k4phknONzQ3qloXnBj4dDQOgjSfLxclL8wRTn+ZlLdz2tdaVUd51qdb8Xk2Bwjiejh
a+AN5eIXPRNC6TzWCsqBdA6pfXfoB0U0ffrl0R4F4eqLGJhQYPwXOzJnVhwNC3GrhKmkL7bFAOhj
crRl4u6Njie4b0tTE1Ml0APZQPupnv450vO9hn6EwMZuXVBBbmnBVB3WOOocaA6t/w0JO8Cxs4jB
TRhNSogmPq1TwyDBML5reuDxuAPU/cXIaZRb3cgPSx5ITvZ2za+eR8TOkugaFNv7gaqdC5yiERPJ
zsVRwk3Fz8zeSCGKkVyCExvvoc4DvDXuWlXD79beDjqKEkutEHPo4V/Gh/hwYAVYjsf4MCpXRn/z
RnsNJmch01UnZEspl+IxsJB9HjDVlWDLqzy9kMSCE2CtB1JUUuZf0K5znZH/Lg656U3xxon6BuSO
l2LhZko+jscsN9a/31tSHVOcD4RoDcmtuYVoT4xxh1XEoqvZyknjdDIkRnzX5Z67Y1Pe3ig60BIa
UWWVDWMGp55eGZlR2xajKygdxBc4LM6nZZbYWVkOFmIYZM4HF7tauLNNN+mtbbhZlhr269SFuFh6
JFMfhw+Zk0j/TbodyQVD6bqj8S2ZzflGlZonaERTXVUOdRwrOGLMN3g5sPlUIlYnbq0u0lXFAqHA
3qJO914jCICKZ6sjLGSQ4oHbmR3Z0kcxdSJcP6B0wUkxtJJBsOjiZW9TvzkcOah7Hfye1RvE5z+2
Z8dS3ALnr4GRk2n+Urix9Hhn5iDCudbDMqyXPtjZq8s4rn7vRsYqRoyStMyDzNbzqD7o/IPeDSqG
V5m3XASSg9zLiZx20owbm82wVgMtPEwAHT1EpbVqSkRZN3A5iqMvhk3Ox4v0mIdSV9xF+z1GBs2J
DyV2XZ1P6TV2p+K/8sJyjeSOR6Q85vlspnPt7rqvHzgCo8g7c+L7yjqZ/mnoPZUrM4laD4KQ8Dma
AhTPBMkrA9XrvpbL7+5B2smEi76dqgtmFj1N4arZiukZO1IM8S3zJ6TC56Q6NycTEoaSMLWD3lLT
4YP0UH2kitd6WWxJYNlrBpyqHd3E36PAfWrJ6SetqS9C0/UH/SzBIjGs+zKTq71+VMoK3euDtvxx
SXanXpFv/rXnG1M4kXMjJq41dbxWQBjPA6beBZbqiOMmWWzxUrFboMDTptB8VukUkC0PM3kTkXrM
pQqDaCpa77jY88J1Ps8ZdLzCTCmvzEE3KFULuxoqctg+wDQHBy29p9IevM455BnNuClZfZmVAors
+yTO0/pP6gfPcNojkWkw9x8KHKynTkWuucqD1Nq2puudsjkzrzRq03bmSRrvRiU7m0dYO6bOPRt1
MItc1oViIJVRa4e4X+HhPuRpV86+QIOkMgo0jCqvkZl5+RIDWi44+1kItBQy18dl4s+fcaf3Pj25
wX2ERSQpKP1YXW6vCjK2P1MoKefaOpSjAkvdiiiqmN2Vcftc6Lo2x2Z7YPs/4iA/8Lh8BU0j0aV+
K10PaP69/izpf6auFRj8nDVWtsHQ5rRsS2mJkbIib/vBnlxvwC74D2zYEfz/e8Cl8JJGSmPR4Eb9
hYPrQfO/S6D2UdSGwwHWIexcRcP6mhYBXVGifO8a6dzoN9Cecg+KPeU/gwvypnYPDsLeZBZ4Shp/
gSxOMH+a+KTRV9s2lxi0BAFtKH+pJVErqm2ZakFb62uQH2YQHpOrcfjivvU4fRYctrRe0vbAb94S
+LgNvwLTulPPJSc/Tvyz7AhmiBBy0s2ef5aRv/NyAP+UDyKvnHZZUFKiSEtLInkqD8YkbWtqEja8
DOu/vyri8ORsAZumvvVhmg0QC2gKIzHLtPhkRVAsGC15kQvh+5hAO6ehtpY8EtGpujzTypVBOGCV
m0UAQI7WawRfK8Rnu6I+S9SHY9RkMfHfcSJTDPe3AMNHQvvlJflKxT8MTrtTRdvVBo+5PKHrqXLW
V5MnY7swzRlDwDCWnGG60Yw0mxYVBcZ6S6w5Nb2QmEPTU4XgszQO3t8hKrOSHQTI8D/An/lCLbOM
6L3K+odKYMSbRyuVWVMCkXqbKFCHIbWjIka/5Oza4XO8FJH667uC0yLz0+Jo1R8YlCFrHnUeyjOy
r8xZxXxzCQU6bE2x1og2fhIpjmyFCDL1tWz95rBp4SOpAZW5WCPC3DdaVTf+ZzlJfb/v6aIv/Nn9
XFt7/SXjd9P18M6pardVYkCsgY9/AeRu8+TlFRQDpNaQgUKgFaIdGNbQ74yirfNHfTdmY7j1IPZo
hw2YG+hd5gswwzvqOg+z871zhshekmw2bYTtp9ILz2j/o/JqeukQHLnk7nCGpIfGsyO+CDdr2w0r
2PY7frfAH/It+4Je2yXJAEVb4HTjmaz8udENeTgxSlOG0LodzjJ4j20+CRywyAHIDf5oQPKPm9Jp
CETkEhjeBOY+Ewt2kb2Z/kfcrzF284EIqw5ZH4kBbvLqJiR+P+oWh9Y33ic46NuRlNPh+78G0z6d
hw3/i9t+JRoo736/yrRObUyjxihxQTaUY1xN30n2zHdH4XddoW12RTT3VnC+GxnfLVMG9MZ9j/1H
t1z/r+br/hGeV51XcvlHRJlXM+mZxbdR9W5HB93SEs/QZ+BVVkQwBaTaJFieYnxELG74mY06zqlw
eLgsQ/Q5N8f97JJa/cKAKTI4DkmQ0lWynqJ7OHcm/QMhydNcXMWt3M+akEUiJwGOxJvyq/XqgXkj
CPq6X5JHn/bVbwQsuxIfUVKFVAFBz4Mj1jOmWXoTBAelZUToII0WURNcni2PUWY9xb1oC0GhAaV0
kZ4sZrFmrXeJIrvwoHRF6PJ6x7GAt+DIH2D0XSA5eBcJt83deTB9E2gAEEqqiRmIBa8IIganym9w
x4a3tF/gktbAm3+b//sw4fYrimOR/Ek8urVEj0YtJAeXCt4I5OVB3KdhxFkZgeg97oAqDH0pSisu
4QV6IZ3lSgbS0GpE0oUMxE+JxkAAJykXHBdE7C7xqlNt0ypmPznu264AjK6fiBJbrIygKWVLbks3
0TuTTGjBH5ONsZfjhWKXAHJzyoyHYwC+hfw2wwCjFOBwQN1O1EL55obN5dbGYqp3mRv02Y+AY93Q
1rYO6keQcPvMlLvH/iwtlBnO8WBCphKBj5RdnThiNOfFqDBsirzt5kr5k+YxAMNm1DPQ9wqrFmdm
f0RC2wSqhLCc15SKvMHfULWgv64pF7BBBnKUTRAoFX25PswmPxswuyCJ5sZhQxWSN/QqgdAPhjq8
D5cy89IGfGrJoLJ/JuBInElljeEmb6i/VErxM93cXWke2dz34NUOtJb9RQZBeFA3rEqclWtAcuhf
xyp9h2ob+8S8ynPv/Mo1213WTdkfH6OtaTFAqbfNSnrERVxTee370Gi9Wc8S8sKi1TRWMo2w2WLT
HqyPQmqg5Q2jsepG+K1IGzkK+2Ek1I6LavMUaG+gTEsiZjDEwr5OArz4eOcuqNrZ86Ya4p/i8Nq8
PexXGUSQCjIJwfY3W3L45/BET57PFlJowFUSjqRhTVCDtc/K7GTqGoklAt4shfj2c6fc9BSZ5dus
El7I8v7LAWSJCyoZtyiW9LpNqKRqeMaf6WigY1WWQBC0yCK/W09tjvv7WSL0BNm/SwCzSClHnSmi
gIe9SBSpyX93cKrg3YbP/3vSmWkChGH5p0OhJodP6eDRnKBlsIEEKiFTLRgcnKk6XGvSZFiiiMJN
ON1gopoqj7jXKHTq1eKHtdrGIuvCDRdMCOBqBSlR09XSJApJ7CpLrMoRb0uwjZb7micZLOKjW3JJ
KnxmrTijxkxajLtppgvA1BZKFSu8Vt9AxiFGQZOwVFlk13wh9gyXKE04+hBrJ2NLJCuOA6QuY+Cy
mSInxqXNBd2xNLnosERLGaF3YS2WSMnW4Ec30z9ZHevMbBGQbLUv1ZlvOFl3h/nfSyPI7IX70UP+
nXMM0JSh9BPM/S9KEDbG6UBP5V4alcMWxs8gNH0fI1hY0mnD/HNfMxmD03BaXDBC9IYt2PKQJBNv
n7d8Mb+Lh7BXOf3kXYM/it6TMMh5mn880u+sC2hvyEICf8fgFwq3G/hBH01JegZ3wZLezTZyPnTC
A4dLAF/7lV8cEoEG5TxOXe952ew0ha4j2bu5Azxb3RqNTRjY1PnClnF4qZ79+UUsyFGjzOxtBqHK
CEQAt4kg0gb+G2JGDCnF4RFAvWpY82Sz+YoqeDygVKtr9Jaag5yP8nQ6wkma4TvYF/FmOUr/Exop
smp79aeILaHuPbodRLxycX8+rK21MQhYnpIXqRnSFhtWSKnBvT/ItMovi0NsZAiiqsfGT1qtquqo
MYw3I5GsI6yE6lxaMWPLdEeKu1HQ5ydfnK5N0S+HbNMfSjzl6zF7UhU2NDLExDn0+LFZPrJbOKvJ
Q1j2JC6DtPZwKRlE1kwT9bY8G/Meagb3Qn5cgriAfnnr+3eX6pDUKMhK+XTTa8ZuLHIwSB/rkXNy
SdaEcQz0H59fRzjn90J60pKDlcaiciK+reSQaHgNQuPU8lk+SLJOdCwF/HWe2eFq1gV01MwLDpv6
NnNlsCua42WM9eRwoEDbAnFT7vIrhz9EhMFyt9cMNzitfMLS3XI9D2DTVSBjROJ8eQCaDu41ANj5
xbzHQkk5ewdbykpT4PDrJuXC/B+VA84uU14bGYXL8iS/EkOJY4LDE3UJYCGB2n2InJ8vyKbZ8GZv
Ot+3XGavsgsd+zfAzYHzM4Q2l5i58aKqiCy+TVaV/VH4ozRe6TzGoWNtsGgNY5eIt61XWZaRl4CS
vAR+xusaeOxuFAgL8uOey+R/RialDjYR3I7k0Je52npc6r4hkVaPNf0vbFb28clF28kTfuHDd2r/
VGo2A/DAf7sASJhbrWtGrLSiQFXg1DyXV+gDHaif6etrlr2zzQaqDt1HCHvo8NCxkhZ4en9wfd9Q
bPxQJvKPEEqaREsKGmPCexilvWDZ88gqLjiVHBc8KgbAnIsMbUFBUUVIhyfzjH9G/rPokOysKz0T
3gGuO2Vbs9uuzxEgR4+SmZaDyokNxeNksAsYGIjN+3Kmo4vnmCXZT5q29vwnR5GaM2+u6n1N/j0P
U2/G1LIgENk19EpuMRE8STnveVjYU+GhlBIIJg1xmkWodDpK0ZpwBRn5wFHg+5IiRUj4MOSY9NYs
t1qBhINcCis3SvR3SbQUy7sbtaWXQXvk9eudNaVrYdrPJfMEemnJEsWesxBeLrbDTBXCkL2DcEMb
RDWgAKOG2LIbXRxP5Mk5OfUJPV6JObb/7wZcgCuFzwUagJFeknDBdhLPqggsTpacy+nKashAAc8K
E7U17G0pfzKe400fVX22eGo7A6C+hBIRCtE2QBbkVnHhaKifCBKpYgQgifDMYQ+7Z4dsVZ5LUYnL
C5ktBnIGbAZi/GT8Q8Yiwu0chQqSvkqGCwuk+PFguc1o7bTHRxfWf6eSg2cu2wCviHzeTjfexM3H
19wV5O25B0qMzYmO+wx5xudlvfem2N+MsMrJiPt/qnaRXTkVnGhgUGpdQb+EDxppNd0WTdETfFH5
FZxzCsrVwiu/DKg8QxgVRLYQQRrz9t54D/hRD6Or6ejqy/9jlnMIY93aa9GtrhEtsrBpQugiQ58P
1ljlX2rvK3YizCbPJrXK5whM3jdjj/1wxPqiCqEI3wHltzmjRkvmNUXxb1qQNCBA5fr84k0Ar363
rZtIX/fOc2pH8Aq3paWdibX8hr/mmHze1jAqrBovUh0RyYMWykv8vu9L/JTysarFVfSHFTitCzyj
CPGBahHYuHQeZzdrnI5bx0ycjQqOrjexVaRuTqTUUGboqawXDibq/+9y5tSyzVC1aYT8fPFmcxDC
PQz24dzTnDr4Ch+eHTVMcGkNGwHdcXLtJk9ZLGl5+gkpY6XPu61/dKXXuH+QGzHBb5/a7PUm55tV
/7m1QZ5XSqQ7pBqm5BF/MY4h/lNVzXuDd5pMrqXDgX5Ge4QBpU7Hfm0WMoyeL5FN8uw9V3fPlZih
jZiqEjQyQjkKkiV5L/5rMolHwOoX6pgoT1UzIbhs+QGTOU32mCdxqh1NFSUTXHLr1dut7lRZDe7H
OGQ9BKRdZyhN2KL3qNhSLpZt7jixcxjmWYbrq3fxw57foDS9tpkLPsleGG1N8AJHbxPzjz8Dp/PL
8XkolN581RHBsTbvnSSHYwmEmflSVs+6KqZU7COfiLlhdyJNieM3nRnkCtSwIs5J+DmFmykFbi7F
upimQKInnH80RV9x0b5nzS8HkFtzZb0Z9dHa0GlPvVcED+Vstt/B3xTgCSDGRrd+e76MJH8lRX/P
UvWuBTJixpS3xcTP3NFrV9Pp+tT+TCtNOI5zyvxOYFYscUAxfm+wEyrJEg0J4zPcC9geLvdp0Po+
d+LxrAmS73T5tEzBs1xHPvE/b8Y9AY9X/0o/jzOAvUJUSNwE2rx1dnrjGttef4DUsi4F81Fcw8Ca
rWxfoTBbpWAqBXCd/s7bIXMc2+SLGX8qisIdEReejMOBehjQL8LIURlupEFsbMnKfvRHMDsXred3
Gms1fk9dkIPXEIlLKXI7BS0gmLwaY2lySnJcnAlDSjrh8Z+8EX5zE+mSIOxwx753l72CVtBtW81f
LK2j1o/y7vv45ks4/PLMcoNZDPvEY2GcMYGnqWUvgcUwFUgEIkCOd8JSfxNGUiK12pByQrVIQDMT
vo13DCSVQgCWOhrAFyPrp6XFB4J8ckP0r00rkTJR504j8+eV4LR/kfuzNIO2EcRc2C/VdbMAREfs
WQDzsQT1rpeYd6s/jdwIZeEXD8dQp5veSCcgndtarLPgeiI3+9YdiupdAqkn9XjeWdctwQ62SXIi
1NBiO0o1miDzdwGmrJZCp24u4C7FZrLo9gERUeOoQ98xOPTFWRLgjC5MD5z4Vi3ySQJ5w5lfPd9K
eNkEiDZIEfzexpGen5eCpWg+Bp0SEszQb13QNjWV94YfevnCVXiajhHhJPxCOqZRJPgOAJKF3xKW
hYlDRnVLFh4pGV2X2kT1NYxTsvPEj9hymp9jSW1QS1ghyC0qkf4nnkIZ8//fmfA8CP24YyU1ZOde
sxE4RBHlflvPSFJdsB6k1ewWUAEZR/JM9BSIUxgWZ3twRHwt4reiozLc7eWt50C6Eq0yN/B3LZTi
1fy5NwhIjYrB7gLihsBUU6MvFIM94KDiY+96TLs3QKekind+3kuk4bSXYwEJf+K+lBm7BghZwK6E
E8aeP2JrvhDhNrFfnt3kRHqAtVygTk0N81IXgMVyrXgdr3Jnw1I5T3qfDt3cmRo/2MlgZoH/B/6s
+B6wAk3qaa2T4uTDzE4Uxz+cbHuGSNieNeCFXR+KKdW1srV6WaUNm1k7OVJO8ujzDIAw/ZlnLBhN
HClQPvHwx4VYYFASE0du+D/f6fIUykTtk7QS0KCu3AZ9GxplVxKxGTKXY0fdlZthA8qil5HsziSf
JykHVnOtZN5QAiOXsztpFfMont3oe4SD4tTTUecSMT8DIt0ebEhCWPsA0up/v3dp9XaRDAUltK3E
LCfrXmIw8CnshjzBcsy8phK36FY+68AavF6zz+i7ADMaZawLiKKzrxbtY1fFCOaUftBdyAKfqXR1
7rE0GrPr11OZEXfQUr22wK96DoZ+cpeQbc1iYGSli3ilxJOyoSlCtdRhKXd43CF7zWZ1n4yiGDXd
g9CO7bokLf33qj7Zc8hyZpqSDxCgIB7ZdNDwsP3lORgXaPQyFutYm7s8RMZlJqfjSq4Rxqb8YB3a
y9MY9jVZoh+m6OqWX1+gPhMdrANz7fPsb4l+d+WSgDCuJpCowhPEIbUqYeD0T5cbhxBgqGAJO4V9
iINrTANTz5x0pUMEInhF6Gjy3Z8AdwZPu2/XKZkrbhbtPHx734IkpNoEULov08fax2J1lhFqIzzm
T+WszwEHZQzcHtq8tQcHuohav+gpBEgd9Zvw1mTn6RBnTzOX47l6VFFQ1oEVUFtX7j7tvBxgDLj/
qy3ul7PxuaREyEptQUXZ1zTBlxmk6IufGJGKirIjljnlnfhFRDAy9DLaEjCK5gLPLvazbCyg/Gau
d9KqLjwuCU022mrZqwgufKQyGd36Qvzx+BLXsj8KrWAzRm0aj+wyiVE3iPq2muyK8ZnAD+9IX9qF
/nu+cZUxnSsJSCLR93RgNB/KHff5fZHoXVxEBMTPHqHPtVFlIIcgTkRheTt8R0etAMvdAet/G3lu
Zg5NG3ZbdiKELt94Icshom/1/iBaOgYu8Vfj/tHKAy+nRwWSRidhashZNOLkF6afzSY5PFNCkZht
6i/I67a8/FfGYIfpud2DY9PRvCbHHS/4U2SBwjnkCsjC6cGy0GK3rhaMZrSqGcjl9rcOPH0KD9w/
HAvGXh0X6Gux0kBHSRIZn0K5sYMSSvaHZZvZb44xg7FfyTWFTV0oaQ8kFvaUkc98fXF4QVb+NY4c
IySL3JWssq1Hy/I82rtYBP9VSqirD5+0F5Drd5wV1AVNclBM/ZhA0gbFumEql/qds2PW4zj2KYcZ
eKWiBxyGW4nJGDAYZjoPVk1ajkQbPQCHaP1+f5Gc21NPvvoHJ1GI+QqgAYOrRML9LIrQ+3gVuTeZ
836bp3TA7nxZ045bXcaWzKUG9t5/zy3pTrfuS/l1PSNztAwlogxiIDOzcyNbdXPvQKkf6ntJ9W8G
kS97bZkmDLqxj2BgE8imr9c+iyZN9rpwJTBsZeQq1a2q8ebn5ZTHgvBjkdx8GIfsDGX+p45A4Hgk
fX/m0cYy7/wQIFh0iKepCNTvraWb8GBDEAd2sD8pLz+BH06SSh67/vka+xNfq+m0lbBV3ETmI6Jq
uofoIsOa1yPUG4MmYo/nbLyGAnLXwy8Qc3iZXZDj8GEKaN3GjmRZKevc3KtO55PZwcat9XbmJexz
AtoKgihukxIAsICiCo+D2djZphiUfuf1SCXzm9QedCfDSlmZG4iVijZwIhF70OUVaJAaoqTzqjBA
7tcp6Qv1ZKkmNMoH5V0tWNIcjJ+nDPzYj0NJ+v0dTacbUiDZTU9M+2UctutKWVG9uf19tP55kLJh
ET2NlEgOdIangjc7zS2TspIcP1H3AY5Ncx73ncMwsHLYiUwjyCk8PcrhuG9/jf/k3ITR743mW7/4
GNesJUquxf8Rt8nrgLZbfpf1dh4YEVyjfWayfr0/OwoXWcVEDQ5HE8QYCDCHLXDH5++owhBNW4Lo
GsbopBI3I9Y+O4Nh4p1hw+bHfZfrP8NSFS+b2EiDr4aXtt9TXwx6YHnNPtoe7TatOfT9Gcz4zLTh
lHvx3wAwyZY66OkCnwVvXzHc1wEj4XctAdPXYTyYr0xHWU26bvIVGUrk9ndx3LacBJ8EEBjNiyif
H/7j7QMESyxEViy0v+kMExIQ5Zr59Bh9Kn7t+EwxSb+YPfgDTNXguSyn9wshNvzMk1LfWv6Z556g
bj+r+SlDIiga8S6vIxMwJeX62KCCj1Y/BhCH+mQiSG0Ake4g6fwbkX/eP8EoGkKP5WjUqeUS4mnT
KCQodQVwH7CarspiO9NYZQOkLxMK+9zf3JqyaMbX/46rNnSnZv7mSDqqxb7kqLkULzfVahVCtqcz
6/WF1ATqHTEhxfzGnErF4XHZVBoRnaBe7vcGAJrcTxsbLs/j7VsTfNeDTeVP6v39nCNi2MthCpwS
9j7nEJRwQ1ETVG2EVxuy6EzaFeZEp1cVHiG3GtMPUC04Hqx/FcOI1dMC2KEhxPp6t8lxlxRbkMSe
fxi2MLYz2TrLw+BIEJsyBLS9UTPEt7oq+/rkArSai6lC3/nqNKSHYO5SNBFjhuNSFqNLLLW633ys
jvA71PU6xaVbL92fCvADWxudRU03Pt1WA0l002U5/ipnifMnIK7L4jfJhRBbLCHunmiUokihhPqP
6JkFPuuUD0DjEmNilsmCMLRp6TTgfGYfbOxj4bRu6C+HxgGroCdcygLnwvyflShjU/iQkYajBjSh
5QC+JkMPtk5+w28/ysnwiyw7PovS3ixJqa7JP2/TL87Xc85rvNidhmPn/62ZZ72LrM9ED+oQMx/O
kMz/i+MTU8XuuVmoJVHNhIdSxteHlwIBzU+ljRvoZn6J1GlWBxkSCVQD9kvnqOE9SJTOa2lLnDHx
fGVzZheQlUzoPzIvkOBWPNMyr9FUEdkOUkgMe/mRfH4wDn4WkHuJZBSAfhhsPLHGwjxNgRAH0xS3
F5EvetewNDOdd5UceCvUrYvrgpjVgFNtF2rY/xMD5m96dbemg/tekiGjOeWYpzyuEsvsMlBEE9H4
xzSPCLnjRyZOFH2LVGP9bkDk0EPeoj53UST+01d+pIUSOtJbONwzJjaLsL0k6SZX4E+imOUEerB4
K8dZAVDNDo+JEKsbPCtw/E3b7gT5vwUZeGk/30nPrr6WtABTTWCHG1VV3h04609DFePR7ezzx+Hf
Oiq6JxhEQx/OOIoGAD16qEejFnv7dqhjNj38UVB0mDpB9A056u+OmTA/f1yCOJgIiWKTXliPnShb
Ch4fPhkCjmV24ym7XQy/xeVksWCMrH1N74vNhVnlbRUwxEPv3FZpiSXPBPVwKF9p2Mg7KY7CY2Vi
dUGHkeGj7jdPyY5GW1oKfU8yGK7vqECYqSTEjDTZemT2gK5cm6PIYDbsqYfRnob0PZLq5MoRjBo2
kXWuBWvLcoPRkHZSQwvbvPCSvTwbLWyFff8cJ+O0l5dSmpn1aJdv4/FJM0zJGFP5nfSc72KG6iIF
I5VthzpWZFlBhXWs36INd7hAaZ/jqWpZz285cwHcZZGdVEQlLevoIROOYeFvyy+CjOZUDtaHQfhS
1gJyJYyQEVBiHpUNQ+gj877p7tiK7X0NROK7yaaF5fffE49it6ZsKvMdYRsvjMEpUV4hBt03VfVM
uV2R++q6UQuo4qd/tMjMdm2rXIXXykJ4KTMP4l5WzBcibRS7BRm2ESklwPg1ZqpUwA1pPD1Sabem
5338XiEC5GdcLr/UJ8ennqMg97ndM/07HZ+j6Goooa4QbgJaw7BQUhvDfotsPhhUdls5GKiOOMb8
fMIuwIElfvRF/9KutOjRY58JwXp5SUyETaHSpHa32NSoOfpGgiSixCytweCkphar348QZg1u+ryC
2ooke0w5uE8FHTfaKpQ9+afeYyI3VktM6XlKGbNzAU5okRrYoGys9IEXvnuIpoRZSnl5DAMddYxv
uuPPeHKm4OYl8K4G1Dkqfr5e01kUcZR4IDAjJ/U4MlD7MuVbcnCmP14LGznAC/575XWJy6XgrBmb
q83amBuKGdNiWnbhexsaCCajspKGKCs87cEvX/9PtU9tYGE45VzK7P1Eq1ovgTBB/3a6vZOF2IUT
Q3VaFd4uD4o7NfXkAOizjHk2uMtil2F5YhyIpXFzQ8S1IJsOYeOUWwqSU6jgtdCTzRBQGVVdjGzO
9ZKcd2SyG2lGVlMUT3P0D0QkrSfiEIYZGrPiAiBYHAkiblTFzE2QLOGqlbKECas/bxAJ06QLVfr5
ygALtQzXwPjJhbuiIDFUyRY20e9yi0dwMvRHq4Cuo/v0D4FrwLzPPcEArHvN1KbMFdx/SKyRqLzv
XA012ruwwGr87TzORhPhEtJhRZH3WhPqPEueURqvlE3bW/d4QaeTwk0kozxx2QhHUco7XxKBxMbT
UIAZR8Z2DsolPpOOB/WzWDh9iRrt2PMyZ5ATOLUK1NRu+aBneNVU7W7qFpIIcn3r3aotuSbeJ28Z
6x+5USOod7cqwVhkfQq9Nh3L9RBHYuQoRaqOxjFnsYMUMKJ3k+wY4jEZFrHro/AyHUhPR62QEWey
WaYN7YEMfnClPjN565KbT09gCaZgYUnzZzIKQ3Mf6L0bd9yccRNmAlW1JJC9g9YY3wB/omiQYJGa
+tjlcrhvw0G63wB5M5hUAvqnYnJacn/T5Z7fLdrtoomNBaK1tT61ZJg7VyaLNm3GZppuErIsnhLI
K1E4toanSTRz19hsCJzCH0VnVXLCUisMgTWkPLkIITtn9ABt23zjh2Km9RXvZMOIS6rwQ/cMQRXS
oA/MYgM2hOr7V8CVPhZtVWVX+RWFFQRAqvXUXZREMqJ5s8Ftb0DMMJoY1OJSd76McODgI7Nz5ihb
UTs4lM1h1uSdWaXLlKQeO3H6QcWSDyu8n+0fuSelc8ZiiodYkH5sWhTCnIuyw9VgRwmbc6n15TmE
yjXDC1LO24Ug9hI8ULPqHNLqPxZ/xrMndqbRp0VVP0cs5D301xo/m2kdc1hibG66JWZEy1o6hm75
iAYnz5sk1AWdMXUN9Dw5gLk+HSnu1OC5IBxHbJ59LYmNYhvWlDSiWYKTbymmx5gCHv6JCGU34e1r
3Si76TrtA5+VyL0wUYBBtas1mJtkmmbuaQjdFaxwaXGzBn5OumX0XCZgcLijmkV743696MqsCvOi
MU1uzI5iOi6yx8Ym9l5n2IqR+a5faatIkUMQ0PG2RzgWv9zaNEWSpd7cHnPG1OlUuo4uoEK//MUO
iB+Ric1TNWo6I0SvKYH8IuyXbHXvWyjZ3/vF1cAbxGLyiwhTvNKBWqTTtjfPISiPq1Rvqs1z8hxe
uxULPuSmiPJ3lZVt0OS1jC9TR9QLHnWM6pbcG4dkjhcYVH05c0Bg+Av8K+gvQLRMpvho1aWBsw3o
Vxt2OCxVRQwa89ExzuXLKGTyX+aqei+FKe6wCf3KPBv6KXYqnflPt5iubawmzNgDJ9fhzEoI/oqZ
Ge7pmQO5Ln3Q7iGcbb8rHAFcChNxxCEjOecikOCKmeHOG8l65uXGBDgjXnPRi9JmdEIyop64YEwk
yCdkZTq0YbnADUAdP2D+gZRHMHmySRZ7eY5IWSgpjcQATKbFPcEud7Mv1/1ixI9HS6HPPOepf0wR
NKpxsrWtzRfxH/OUDY6CACt1uejhl2vIXyoWG1s3Rw/GQvYD4Uaep8D4afyjRG6t0f4rxxE6u91F
yExvRp9xLugD0oZPr1hZ+xsHmCzRu6CMDkQM/Zhct4k66NdkpSvFp1RggFvYKR4og8aNjYIPBGs5
1aaZ6ConMrrB/cFEGfrEUcAY+zznj9fPFQ/xPehX0v26XJFNtTbtYLC/BHYrDARdbBqJPnFTo9q7
qRcJSuVGsEAR6y3Nut3qhBKRPoXGJujX1hTel+cgGiq7UaEtzU6+C6k80t2LbycWuWWrwPWMMgyC
M0RDhvRnMZ00uTK1wXC8xdGHaqX9Z5xm9dogqpLm6zA57ja6yoQrvjmuBZfU8VIY2DkhmsoETD/a
BvmHEIdVdzynf2tW+f/GQU73mCL8EHeiV5em3L/7o9YbD/xabSlQPBiXkwyyIeAGpXJFHAuVgeqN
mwbNTQAiBb5PSjdfem9LaPiOnBGz4/oKKB5yzgaZtnhvGt9VyPHNOF7bWCl/m9gi1Xi0oxM/eivc
KVnc9PRrITLVgp3iTpBFD6pOjYyqKvKG2g2AaCMfiSHCGzvD1y57OWabzj3w/oU49OwuC+gByknl
07A5PpD3Hc3MDmzTYjqZp/XT0EaKXpVDUpH/uZJzLgoAwLI8U++VPA7rpjoCP251noUCiYwkG4YV
zeHZ0GxNSFQND1f7YSV2up10MBkyX28BXyRvRhRiuGt0LU9Ekz7Sh/s5ba72xGcGjX0jQOXkkXRZ
LV4n4cwVFVD+6M9BfjXHbKYDvuujd3FulRUnR9dJUAvNPM/RQiXoV15gDOsKwe6PFERUenB89U0N
w1lXCS9YoOz3k6DGNRb/Omx0BZHQ9yWcWrHsiVI/SUDBnwRxXWa/Q64HOkth9Rgm/sL8oDqEfUC4
RSfrUSBU77wW5+PlFB0pbrqfIKMoUpBgAvXnbKcKPw8kC48A76FKAH5lmH10qKccVAvUhLv8o355
HRqjjzboAUthHz/zdn36WjRrHrnrKIg4b85yimmlmAdx8nCWc64Lmm70WMI9c+LpDftthJE1EJvX
B8I96R8w4gl6qFttbZ/60aaf5WZU1l93Q190e5clRW7HsdJPBcKtpNcFW9QyMS1AUXO+RRNGN8Uz
wLf6IlcmhMdTI6LwdqtbJwU/KHPMqXP5qyDABwqfZXclS2LjatnZlzQpG70NgHj9F5BQoqrsKmfQ
RydqTkiN4idVLNJLm5pTn4QNeiclyuYMnNuCmRsxS8vk0k6Kgl2F3Eq0UmnHbfOGMi8ijh+/cXZg
KRSU+E1kvDB9kTI3p2piFYt5soJMdiiAyAh2hBUO9HT+G76HfOXSAl3DzDgiuDdpr1QWf7LZ5JSa
FJyoAJH1T+nzG1DRaA9UoNpdl951L0zMYi2SmamKJalSYLNZ73xkMmo/vynX3kRcfp/McqDIMPjK
/TNIgBSVoyBOKqfHeETKtdVPeWeryI2VreQbpoiyP/wiWySAMukI5sKLnMP5gokZs0ztqMxwvTX6
U9/RLpScFqlQYfJOqirsjE5duThZ57S3aCtBDK+Nt5axPd7+AjHRAW5R+xFSNzEao8trzKv/LGIn
bt11Q0KmhjV6JiHG39HMghpgKurDMsZk5N425oHIkMw6w3ez0p1WVvmze6WZokNfU5XMOPlsm5FH
eM2WjncUcRUH5etFJrK2nHBn5VNcxTVav6ddfLbsKl+jRLg/4wqxsNC5bW47qGeG/9mxc8AqzM3J
RBXwEQgOxejk49CqQLkpOsnqPy6t25tsHTtwQKR6qd3UdQuMMcFh3y1Zifr1xSQ/bPXCi9ma4FML
vZfQ8CPogY/xRX/Uz88RCB5zSRMuK+JFHVXeKiesnSd7orCSS3e1ICRz6ZiV4kveGAv7P/sGkrAb
1BroWCsFNKK591UzoEaTkGAMsVfE8qBtIYwS2xee1PSQf23ykQC2ZtNIghrFi8Z+XEFH/kR6WwFf
essxMqAjBOc4OR5A7abzVLNnfYWMJTMyRhZiCkwR6Ox1pTVO7whruTWSs/e216m2kI83uaztNWBc
6c4hkASvXn5YOc6H89RjnsCJOZpGvIutHw/KSvDsfp6FZvnE+lfV3vIIuapRCvOLtaC0UyvXhbJW
pAdRyNLqHQEFYg4ENBxsvNTZP2vju4IeCjydx+YrCrpMVKaF4P2WI3m0s2s+5n7eYfjf4kkAb1V+
6FyMo8JsAWoXgKXlM3450tGfx1FvdQ8xzeUAEpbO+r3ugfQJvCWyyuAY6m/SA/P00FzAc4gyWfKm
qaQ0hL8bBCjDYUEYcc3IP3huunXbSaRkz07dL/FCJtlcrK0NwJW9nZCD+KOIG8VRl+usA7Zt3Vsd
n5Sbrqv1aADLNPKmvBXYD0nxHf8uJ6/LBMHgjRzb9bo2MuxN+kaMlhBR/fXNnU9a1l22j5yo/TDR
qJAojwUeD1VWBhf4ys3kV6zpLVzehCSagZX/5N0pU3mKUW/zTZjv2lMi19O2ygw9it+5xLzyvrC9
w0IHzhNJfhxcvMIY75XZPsG8ysdcsE3KpwRYCf9TToZHtQ0C3VRpPLLbLtGQi0w7xOMFTXHRJXGu
VnComDvxmUwLgrhjLmFL4LMtNz7wHBpnTLVGjRLlb7nnqZnnObsutOu3yeZT92ZvjD9CTzSUPRap
MQNnJHZKQVRLN8BZcol3VJkF4uqYyrbCjL59a3BKAAzd4s7ae6a9vjpMSasUNocmWpuF9P56dD5S
KADNaWK58gCfLBhwyBuj6xJljPj60OuWqEUGpqRza5C9BXaVLQiBvlkEN5BN5Hm3oie8y5I7jyBe
PlsQhODP0qPQJTMssH3umcAG7Hry2x706pIvxmrr/CCRM8II45LaV/SnzBCEghD3fuSatAOXA30Z
hojJB3d1FiT1v/CDuW/pqkmttyBD7TLfPPafmaH/Tgta54ICd74DZlY//Ocf0qWoiup7A+u5da7P
FD5aELhcbhrvWGYWNSGzOq332m4Q25pxGPGgNGG+SwCDWNi9xmMIqmw3BCQU3n6bYTU4MyEB+aLT
RQvD6f5iiKfzLiIzMPjWfKF/PIz1SuTj58vJGUUhYK6ahI/IV8DU1UZrvGFFldoXPEaJlGmyO3B2
kD4iwQ7K7EYJHCCHrS+U95qv9jTehYWcZWCRTnfvz3+Qg7/PZBHZ1RuDVYA9h5dLbwB80slseh5a
ffSSWuodd/OY4L1L7XvyUrtPjeGheqEX2kMoCER4cclJKwjPiVvVCbiK+Yzm4uCY88RCT6VBDXDI
D+6qNhg2V/Uq7bxTnaf+Xl0HLT69Is1LbUfVpLm9yfmD7nw5bKayOndJrs3YDKLQoMvp1wi/YOaO
rhrmml3ivltTjdye4MmophJI+cWwnT50Bv8ecZcXf10oVgctNKOafFGkVArHO42NpmuDXb4LtlQl
pL84gzrzBuGNLbpQe9SU0L4Azdqe4T4ZJlhkAeN0PAA195dJ0YGD85UmcY1lgXFKPx0ZvGY39W2V
9CQfDznFeMXeJOjE2sicyMpfb5ITsmbb8r2mgc63/cTtXdfDvc2K8ErBwRCPreTxrO3/9z4TMcwX
cWcCcxRB+dkpndpxLzq7q6OHcjtZQZgZNyEZ7BQSm/P1l292oc9nCOWwToByipNxdj1vu3AAjGGo
UN2wkz8/Y/R4fH5Hj7UyimMGXfOCDk0aPbQcj0q+fs1lKOGyfmFkAwSzrlI9wtUjVp1dzFidzIYU
Hp7sd+cg6zJ8pZ1lzn4PmAhlJflAtX8sJkWm2WpeXFovcL9rfbZuTHvOchIDknSDTxXMBvRvNHnW
nPWTTixQEU4QNrl8UY4tRPu7dzSCpF2+UZiQXedKxICGM55iZFUgg1bYu7WCRnkZIl7vpGvAZiWl
+k6C5qVgBNC1PIYTYFDP7vrqNipTxs5ujO1mtV7W8P+Tr5oMRqJnxkXlFxcLxzFMwFTSIITB6HWr
u0TShPX+Ed/GOboutrCOp/7zf+Ow+tGwP5JLEMJulMY/83h8TEiGuHyQWXpeHRFHFyzLyAF8TOP1
3EurDdK6N7WxrAxWNQAF49VcqEEBSt6I5IwG3TYCtFz0wD/ZjiagHma/tUT4i6+awo7TfmtBnVuP
VUGb415ZwkyufE1I3VJznarSSl4+wiTx9QRezvHHAFBsNMeyAsIKtQ9Ni/C/ezO+piuFTHqIdz3R
oPWK7TX0tXKTNMQ0S8OEQdSSXYwhbu8wYH9llSYYuIiGr2KA1xS0fvMlX0XaJttqj3zWd6eMXZrl
co7Q74cWU9hPnhZgnCS9cXEz4doau9Y/HG4KN/qJEC69+H/YSTvf7avbNknKMaTpdWKYb6gt4E6w
nbX8v7yYOYp6w1gwgFMqPOi2kZCZqdtoUXnu768WZLNvsIIeBWEnXvMyYCxWf/0lJfxkejGeDHvd
RaRLFehlOg8ZnHS7YAOm/Y626n6ClACXZRQvbUe4Y9uo1L5iZ5DlIE+EnqyFN3hQF4K1eTpSrvYq
mN4WMmn782Q3ISkkUSoJeRPMtHBzQ7UCD3pdakHtNGHHPjO8Lsue/f+wM20htIhMEZCP4a/SlNQX
Jel0meHnN3JlxJ5xFUSMP4GzBzDVSEJ9FToSBzLkWuC/NqSvVE4IVZqyd+e2/o6jS7vepa0mkLD8
5XcM91E1nd1pjff9CYGND/x7yPHGCvv4LFbD8LJjstJ2UTYAj1aacrEo+Z73AaAP6SpLVUAM6K0H
auGe78Oe9ms5kz1h+rQNO1rpbnc8F+fuRO5YNIWCYMqEP5VybDfWaufyyVsbTMw6PddJpO9aROrj
0lLbFAkf5JyvEzPFIajr/upCUWL3C3Yn3VgFpbFhgAdqVWy+6/W97gmtxbwEPXcQo4tl2MREMO+V
ORb2YD+VHsh65y5soB5D1HElFxshKSqEcwXu1qyI8tQLRKsQZ+V6vQ5yzBhw/dmA6AZjEAc07bDO
FYhOQWMipQj1q5ck/78dDfbw8qEs7odGG4vRf0TiM/n4hOCdBatDqkQJIbG7pMzFV/LVa3PfIDc2
PkW5EdZzseN1AB3l72BYQTUyWbMv5FPF7KgMZemdhHQvHAJBuQFrqisttoAJAY4T/+nLGPlEucS7
Amx0HZ7Dt5cj6FiNsARFys1UqwM6CzDNh7QuL3E1x97kdN8crcEMLEU3AzYUN+7kKA4gfW+RQEdQ
8jn5d/dS5KHzsajIZUQVeI7gcgsXhUFrhUZlKN05HGH2N57IYtwhxiyEEpFyPsOsXkjqwB7w6a+Q
ysruu7lxxkWJU9ZzI4lWQhveM/EmYYgqseTMb//2GFJu8L7zzEMaTbY9x1KzQEIuB8GgoRaYk9TY
OWl6OVgHfvnUxytnjvX4jyANbhZqZ4wlBGgZ47rzj1FtLAdRW/jcQozimUYXhu23n8/JtPhblZws
haMosQ3lXWgavPpoeyVlmYcmdVJutYGAsx532+aKEu0biWf8bCUtDLhcYVeAEV4TBWRfu6+NpQ49
ONJXDVZ34rD+zVHX4ZgDEGz6BL1V1js8pQ/g8FHmmneTCUEFf6g/hYqMj32SnQyiQAXZaJ1r8FqH
zghYRRmAqfWfaiTSiwhxPZL6Knm1M9b51blolLRiCCipWKlikJFX56FZorP99cMOuy7KhXo6bk7Y
vh0QAytDk1QuLNlI29M+qMYF4OW+YmEtj0NqNtxQh8SzzCQlNG+S3LVsWWP2ufBtRzqnoj42p8BH
g94T2aTMwyhxl4674pENd1ucfgvyTGsilwu5YyROciE5aIelFblvDxGKIxXultYZc0zMz9CvtSNH
xeEcXD4AfgKU6Ys+aZVvHGe66HTGFRke0j/EmZxaZQRkxW11lZvqQIPPgMtzcZPJUpF5G82mizvl
tFYi6aEtMbfZQCoKhgVe4MiPFR3Hvg92Odu58AeSf5+2nOWN8xwR0EjHFi/RuRaTcSPDETxWhTI/
BeNpilWVl8Ivi6OXPGb/pcoSNPqUtUsNWejjZyadmP6NAYAKEuBDipXfBS220VZZ9K8VegcRZ6AV
Yub9io0bQeDBdNYR/gatCK1BK2YcgLHXgqOS0M4HzwwnFBiFDwS9O3tCuO7QRyzexKet0SIBDwbz
GbIwdA7hf6H0DalyspjX6ouJVmwLzPh+Pmi0aZ01DZTbdy/xnhTVPYWtVyKTfW5By4QvE80zCkd8
7oFXi0PX1OVX9WmcPBeXvmz+RQut+YzjmqXMaFjOTDco1ujzLhXUbJXTkIPMhaze7sqAu2sSgIll
Utjh6+GiKMyGmjWeVFqaSNGSyFj7ed8hDRhoqe3YcYjPGRSu/88OvEVWNevoxEQVx7EuUoWgvy1g
MF9xfYI/fpV/Jg8lnBgya9bRg5vnp1AJgAZvElnf0caHj4w5bl9sxMrbJGBUwj5z4UgcNTlqli3d
tKh3EixdfJYt7/XapyysfostTavfMgAORo5Hbab1NoM5WixUNVhUTHyoBnnCbCsFOG8DeqUm9eSY
WmEJQN6MjHBNcrXY8ZHAo4JQAz4BXdCgHicPPELpTm/mtaH63Vbp3dVqrkB+Yk/qymoOz0jt+YoV
SZe/jeUiqAsAN7iBXWsvo91Z3s06z5JH2eHaDTFASw20NOm3e3E1aP3lLxJqXsaOUbM+TKotCXur
ChSeLoAtl2p3VPv7ToJdO2fC5DFtcZ5vTNQZIYsTldOaHD4xJtHSdeyQHbvS5gyLj3FrDh73vqFX
VLXZ9gJmbowjgaBFRE5YIWvZMvFAsQ5PZ4bF0tf2XsYmJTNzfrnZA9W0r68u/szbWHNG6x7OJGJE
6ygt6NTNGvpte3mA7cd1BMbZ7b+Jd0bYaHe3YENd8twR4WhJ/9/O6s2nO/CU9BHy5Ybw9yJ2AZqq
oBqozx2fqY7PH96a+wD1xGrYRtsg+sTFR3PcoHsxasweZUqeyFtpsCfK/VyEGqP2+tbawR9hzJfn
wMyLpHaZZ4grgieBxREIlg6rK1l/8u9zgNnOIyKxlT8X2i+56zOK5WDP5/QOjnfChRi25ReAzujv
MdJA551IHDspggm/FGef8cl7spTlDpKCijkcnq/F6lP39EFy78TbvIPbgfz37hkVUkRplJPVmRY6
XpL6JEODmNDaYLcO43mb0oUVCbYEDjCkbCMKBxTaxNXVe9PLOAei2FvbZAKzGVKyej8/Pi6ICluO
vbdbOmQpKzoCNHyIXRnlojuvurVGUy6kkPadYvbQ35R+xImgHX2i1jmbKaAe5lloi6+RDmo49uIs
wAQ1VA/FlcTQTnSseysqbZeFelEcUf69fMde2urj+lvBSVSWdZSF3FNmTf66qMkmvTE/l3q0l5kp
zk/9qWu894stG6vkqaUU8eJe6kL1d92WZ51IGkHVjkFxMpWPbwo3+P9LLtUB0cQCICtP8gaqQGdx
K4ar+PmhOIzFNzNw1xwMHgyvNv1neVPk0McNyofpj/qaCr65294y479UJanz+oEw1JOOr+5u6O77
ZSfyTkSvKLXLjYUYvJSeAb/Uy9F+7CHe4i3X0EN6oRQlVnr791MZtWj2Ey53KkWyum6oCZYOmkIp
jCfkaP0sWEAClfgpgRS+HJW50CM8iT9iVnFc00nzUZf2xLRU2m1lDbLAH/y7HRGymbs+ECWYFLWn
KwtlAdXqdUEAgmn4XCn2a4q7eVx255cqarBLsTplINjb4Rq4EQlY/m+E1sFjPMhIjTzPYXRb7sXi
lIUR1Btw839Ivo9QsColZ7u38eohgzeQwz3q2tVQ6+nTJxoiwD1Ge+wa+9keeYkRfW5D0tVzTjYH
lXIK0BxL9Yq2gSH3BYkqWuYI/YQthyq2ubD54cvQqrASKBPxdobH+DrzOmedBZg8FAM3yATBc6VJ
24z60dND3NtdlVc6SMdRUz/61ag6wKFcmie1CQKKI5iHk5IxHiCNxBRsM4n4sR7ZSSEsX4x8+ggp
WG7s3WhxEL0VHKaC1qjb2efbbgQkXvNIGLHVyUwKOmUO2EqsS6cV/nPqF4lUclESelqsYhPOMBfY
liGxVfCpWQMRukUjKntEUIRSYRviiSniDveEXxDMVExUvHHehKnOl4HM95IBfL0U3c+b2B9ofS3p
8bgZhT1rWE6zaWpPm5JdGym9TRAQ4QdWVBwpESZ7zz+dSXoLBstjd3UWZB0YgFMWpL1nfcW9Wfx5
nSnDRV7PCg2OiGDKKpBneQOOf98nTW9jpYewTtPpdEolaKZuSQDUR2f9LJT+pdzDkiUPdyFG5LlN
NeT65qUAM/osSDxaEEqO9/+qc53rFBMfJ02I5PzB6LbqnzFnvlMZT3kn+nNxx7hYP0q0kOl8+KQm
pxwFiT74xNI+nlqqPCWp1iq3VnfFp/m3P3v2akqZDaZtpKKkK/ripqZBSvA14EE2sCusgeSgzMdp
WNQQjnp3nsP1fMeEEE2ZTHSWW90RArqSZuIj6yJcwT3Cz+wNjeh8CLL4UxDbGoPk7QxAFH5yKIw9
gOOoHbjDeFXMXUXZD1c+fOgxR8GItu6bNFt7km9u1Hyg+w/JEFvf8c6Og0qRaRHee07I0HuvGM9U
uPKkHmSsuH9D8A5A42JOPOyadxlRxBu3gEAHLGDUrqSbIIHaog+efTzW3zkQ+3SM1m1hNjZxFrNa
ui/H+xDtnAS8Csr5XtATKN7yaCxHNCKEcAPugDxhLb0xdqOHXL48Ok9mAgO7KlI9spNXdT4JH7GU
OQCe5Q278qRA2SUmQNOYFKAyEtt9wVRJphp4ch46qQdf6vBrZ8coCUZA59mPi83acMUSnXW5hK6k
uD8XFVH5v00Udd/7hMWEPAsy6/bHsNQcSlFuFEP5T1TTnhpFQIBK3BQdAE+yIRTjilLGd+foW+NU
+/HpjPYVjuGilsJK4h3s1lP/YV3v729Td18hgcXdHkf7MWsX/iy53puNEBbJNhYp6W3u4D4nUrIK
08Vlo1GRbS6yFjTaY/sGGxSfDKAAZi0fCw7fs41ETGFz18IgC1XrAjCezZfMFUVCDg8TrJGM4v23
8EpsoJwuETL0hTDnACp02azizVUHfyNvCc0QpUTMONLTof58lP9v2lJKmE1QDK7sfPCZvCgn3mjU
CgPtg+tr0UThrqRBd0oy5jV20lWkp93fJbLBtGkPgPAtrQn5t8A+Zacq2631nXvRHFL1dUbJgH6R
35eM5cEbtAGsM3VxYEDX443qbNj3fs6UZPlv+dF9488dfvzKCto60YTi6Tsm7FrfVV2fzz56M0Xu
uDeYklGvKO3HcNYydwh4pbXPWglChZZwKsT4xLo141/qbaZ9/6Qr+dwMEq8fWt7c//SXQXEMLu0G
XW5xVjQMpAd1PXxFBAY8zbzypTqHRzNOrHKLjaJHX9VxZDSFdxs8nkWtqPfJ979O+fN8cuntRM2+
b77UI02pYsOX0khqMVhvl6sIzxuFUBhyDrKU06hc3EALWAZHu9pMDcFIvwxp+w1mcGl15T3Ob2iN
4Ik9a3A726Gqz/cvH0VyNOrHsMn6DQYuaROkfhMbxmK8RyQqie7N78yNA6Ejgdn8jXvqjuSEfTYV
YoR82XbpvfqZucYT0MWcVdbxcTVmcxY7Z9WHsp4ERV9NCQ/HUjH2OVAHkofUsXGlDzn3KztMp9ah
FOrRCl4a+DFTA/wtCCtSfC6MUnHscv04q/G+wPrM3A75oJkG/8LM5Na6bTegzyvjs2DehdZpfsB7
x75yLu2cl52Hxs2QcFS72bdUySc26TT1xtJdchKDQ8JIlri4HMjZCdiqDD0rf3OrJSfMYxM4EzFq
LokxpB+f2ETg13KsHNhiFEnfVzF7LS7I1a2RUdQ40G4XbMo4K42e5piMnooCijSm5QlbNfOSj/eI
JzVROt9/2Nb/qxNw7e2hnIjwZmEnqiF3pzqgsWJoFaKRMBc+o8tOrvZ/0G4q9rP5TZvr281c4bTV
xIUtU5+2B2twuey2mmVXpLrERpn243Pzb0ZJx56j5VxtMIMiLnAr3EyaY+of2abJi/iRv/HFnak5
JkbLUGye7XiNiZxE+28iUv7YNKpMpSqTFZ33dMBXrl8Y7ZMeTrcGLPlyniM8+/ZBPMTnvWd9QuZY
l2bd/9PdurBbv+nE3Ln8o5X1iCpr/X6eyeXG23OxzKMAc60YddA8nfMoWr2CCkhAYy75GI65giAX
ut1GxdvPaf+KKzE+vLfYT14h+DlGDSeQooB8MWBN2J6RA/OeZvBtq1ezikma4JFQoadf3ZgDePrS
RqygvnMRYuDwJuzVBBbhJ8FL2Gjfi+DmQNRJNlF2IMp2yQ/IsJvaMFnMcyijm2b9ov9+rxAHvt6f
g74+VlxPcHfGazOMZSDmFh9eRMDY1kkt046fKN90EtJXPGkceAUW/u7tqp+dCURMUpq70gB1z+Qt
wjjaVP3vw8ZTUzRW6ukym3xRQLyAHizBtCNfSFaThOVB4k/U+5XIgDNXeWKhJz2koCC3QYSZ4BRG
6bO3dDD6rKVWXJJIRzwyByN8NrWqNJgbqac0dfWo8W06NwBwEbYNDToB+bnKiZZuMxAXvvx/OXpt
RHek+mObHuieu2+tmmVTwQ+hizg7gFIPJLMfKQq1o71yCialPrUtiI9ZJ8hMKz/em6B1QdSYQxAE
0JNWB4LtCduzjqlQYRLvO200Z3627Eng9eWE5PqYZp1AR5/IIFdaWfMgL7OPyIUpVM+kTmXkkES/
LB5xs7/oLiNO73wLSu6EvNRJCphQRKmXfyHKALxkkc6sbGH8dMVsS0uP14mjB6RzwVjjjTRVt6V1
md7/HjTV5hsAkchAM6eAMENkrB+rurFoxFWkn8BcZEn26ngQHu1dLQZjWHbErvwvFhrxetUgh5aS
EI7rQLlf5WH/pojabfwRbt4H9v7R7v8irjQkqSb8aXUbQ3tPYlY7z5vRPfEYxDDULAjkOzfJAHWw
U9Fwsujw7p+YZ8I6RwirzJZ6AFdFZgu2nA6j41EgkOnPzhz0+afhBT5qbYv5GX2So56nkBcy8Bsb
y1vv8r3lyjdph37dPgUmJlVxppYn4FuvVCNgw/H1I/F0zFmi6bdVNvbXHCj6GGb/afOqIsw3D3qV
TWsGZQtWbVS0vWtNm9oTFT5yJN45GYORhq3ovw/Ln+2Jh51FKWTVA0K2YQNUP52ozZIIZGsvVD/f
mZ/JKFjuSXDJfdaH5hHvIPD1Y+Z1MqeLmPvj8M1Ma5dK3qchUdLjTDM2Xj7mcEFnhzrZtzdic7ZM
1jeVJmuxIHJiz68p9sya8Qw1QinFfQU5D5Gk2BKatsfz8lRbh9EKnyvvC20Pn7kF+7HTGNTPdADS
0SBIS77WlRkJjRw5YWcTNh42sGOcqtV0uSNl6xmZJBXO0wHCIeU673sPqI/NIZ72eqjDeHv72nXN
oXLAS0XmWXxoG5XmjgcyIC3fx4tiSc00YP8M+T32EVRRmBBJkg+5fIEwa6NE5k+DJkDDZYAbm4wD
aHTfo5vrqNG49lhUafweRR8PjgC07wJSWW/VFszYR4XcazBQ7i6vfGSW/c7+WPYlsWmym8YdUPA2
5tX0ud+0dvZNrpsJqBM1/gruF9QGOyex8tj/ZdEHfWLI7T/iBhfONC0EcmsO9BZ1s+J6uSjltUpb
oFtJc1ecpkOwa4iQsOwDNyrecy2vg8ztKAnArrM0R7+UzddD9KAEjCMg7kPc86x5ILx8BCQGGCNT
uTaWJluExJ6B1uQSuWM2sSzwP6ZbnXjST9/xobnydcvgwE86HvysQ9UduEP/bvA619kqlnnKCGGx
ioxOrvhyb6NwUtAQR42PrkKruCrIQ8R5y642ceo5MPaMd3/K4oFnq8zyqm/6eT+P/GmIARXoz96X
TN0I9URs2z/qm2naIROjXn7wKTyA63ksfwmMPLB7qkSJ5Ltb9vQ69AGbIAQC1Yjaq7+xkXFux0IK
8LwwZ1ftEnqKjW/+C2elNmgYkdLBroBrcguhYJyNfTyNocZ5YvYIVTzxEKpPXETJPdfWNGvpXFib
9r9PnKZngblQDRv00wtkut0AlREJ0pCrDYDUOyQE1qSfnneozm636+BO89iadfOAhh8g9WMbpdZ/
pTbnradiujoblTYkEt7t0O9bS9gN+k1l7RcuEdAuzHAUj9Xd2a9O/nx5ACRui7R+XTue18bIDfM7
RWbgyIjesLRz8rIbDXOZ9v1hB1ld9qk7yKOGz1jYVYESF2rF5IoW3a+tIcBZn3+nYF2NUZsheUOb
tgOZYTtiCkbcLyyzcXhOUSHNbUufLrZ50exkh7BQw2fV2+fSi0JL/xkG2uBnOpdrdMQlVzIAqXr8
5CT1tqb8UjTdsBVgNsIDV1pCIK70ew419wvQPgwCEy2HAFCSmprA/3pZIlpyKe92CDaZbyakexRX
9S7m5buejND/XPcHAM1Al0ki/iBlsx83L+FfBNid4Ehwvo9T8kIf21NJbEEcRvl1wuVNWf0Yy3va
PC7ZAswWHQinRjN//riTcboRDkBQYGXJ5ADqwOJY9qjPQi03+RTZmX3+Qiy/3VgySJ1Knj3bczeF
7XBPJhi7tuaAHHiiUafDhLdeBr62hHQ7YGXhgQtwuhL0HuP9a/vET1UdWy2zuSazGFf5/UJ6dyy0
9HyW+fJcbwlxDsL96uGawEVNUDS20JFRBXf5d4teNlsyOeghKAWVFhF67jnwEQKHjs7Qgc1mOEAS
tBfS6VZeXx69IfUhyZWJoak+lK+aMGfQjBgYduK0sAWlATEsifFonU+yVIV6OobCTPhUB6t/wwWE
zMPsyhaaOK66LMRgsao+wlDmCtEgy4tc+NdT0By9MI1Syi2fsmcU+Wt062Xgqf1MBwKewSj2z6hd
AYGyQ1bDHOau1jRO9Qa6Tyx+zVd1LLktBNkN/pAVtWim55qtsZf+gshJ6oodt0WjBP7t+tBGH3ng
IzJOnAVE0Az81BDBRjAI16PUTiA3vU1G7yi3x2pBhnCWHw9FFX1gCvwaS1DCoMpjwY9jNPpEVr4B
bZRGHOPwK8ftTvLWD+D6LZFCVgIanC8OLynvztklGljkLpP3gXi2youMWj1ac/ShALcqUH1ccS5o
tLdVc+3g7mQdM64YPI5gmsp7nGi7L68I0kh3/emCMuP855LiHpQ8LccbMY/lX7eo2Xb3cbozjLH6
ZmYrJ8Hsju6MePQwPHUrv/YqnjUy0Ig6KDi3/nj7SUVQcm4jZa07R9961IK51BZLQjguqIMptYVG
Qm5pOWOB/z+he1U5plb2BBJrD1LmsOlw0tzFh0Y8vroLShP8S8CEU86WZFuHd+M0/4SZ11iEnbzq
96s8HThmd/y5nKGfrlMbohkEoNy7Z/nsrUB9CvN4HGYSZXGlhAo6r76J1f1MENJRo5TMsy0Qb3lp
zqP0b8o+mC8JHuAlxd5oBMkwVTmg5/U9QRjeobIs8wvJ5aJVHeDzKKCWQuQU9xMgZe5RbvBZM6Jz
t3tCgxsdDnTkkDQDqQ9idaCiux+c4Klvq8cHriJfgCfpolEX6Dwb1AFtdpKCpDPPLxx86/jEltRi
p9dVmcvCVa/yi3zyY9/OrqDm2pPymQheDABJYWJmK+JQV60pfyE+E5htQBnX2LG8dpahXwEBFqMu
n5tFBHJYyuFCbatEApF2NUwI5upZF0fuEcCO97b1McUPpZLTyC2KRUU0OBbCd9kLtl4vHnAcAbK+
GhU7K+FBow/0SvROf0XYftDgCm6pQ9SFuncNgnNdc1YdfymYe9o+MufKMQ7Dw+meU8rPNxRM6fdr
/BQOvktpARSBwQ38SrAMRVIHy4SS747jnYmueNHZMGjwdRcq3ayYTU9aw9Xe1+GmovO/4WX/log2
ZLSSb8TSgR9beg+zAhMUfIzyDIh76QHrY6+9g+ZZV1Nnvg6/mj5xvDheJvIHShbyJuZQUC/M0M3i
FWpiUCTDRMHqbVs3tKUGdCD/fkuapIe/UU8uwlp5ppJ84Mx1uzM6RSIvH4hcz15UaWEyd01ZUAhL
gx/+QPGJJ1879FffsQ316b1AnFbXmkFcYaxxvhIBHsRLdCbJ+JTjTxRAHGXjxmY7pAIQdY2SF6Eo
7kwx98m/zWIVpkncWAPb9LrBUg0mjFQ9vGxo9eGa/YSnbyDm/+DxwIP1t9Qyf+LLtq4x1Hg27eul
yJjijh4PqA4kfrehIFA/oyc7knDlLUCoErP2J1V+CsSPC60IYMHtGqwIO71eD2aLATPr6LQJ61u+
hYhUxEajdT12NZBkaVrETSVlgdgo4SnLJInFFU1G8rJi4VPPZsmhLnK1N8uBcdV1Z89vhmfM4/5g
x7D28as1XPXl3IGaG4bDkHfiVCgZ2CCavnO4dP9B7x0/JBBgZWMRO3n6xz067T6IyfCwF5vatULh
sYVVTq4CFslFWaOqc/k/8e7ralPmIvUIYgoM03dgA1/AfbNqCxl29AT8JqIFzUYZvL9b1do858bk
rCZvzYs40Cv/9PUSYYCyCE7tTHW4oupEmXYHYjxSKoIVXGBpIYg/39czLssso7vWY43FuRLSZAIv
0K9k0Heh3H17x+nElUrX0g+tvqMEzNL5YxNS44RPRgO0X7G5UZR5CsTLPutI5zekFRxSCNo+4t0j
FIp37aTXlAcBzZXUtKwWmsmvhxkejdEJ9RGq/YP3o5wejcsz0jV8jfzboCLV6EaKpzT+EtmDatoo
CHJYuh+XppDpdEuhWIiA1Q0Zd5gHEY7haXSM4qXWHHmTQ2viDDL31z5GajOargl36rWEZfsekUqF
93Vp1fUtsvBDq6Ks/ix7mUWijIN5EU2l0DwqR702RhBOD1GNXCMToNbczLWP7nEMFE2+0fs4gAaS
i4jx3tuuJu5ZbROoSX2K7afjwGUDhdXVRs9cDuaLqdRQQvbUSux2b4EDyTF23TV5g6X1kqWfHwZy
TZydI1G7gKBeu4PwPqAMudCIJtypGKXXCr9bHZLuQM410S5TEKK73cEMH9G2C+PQ2xBSxit5MfcY
Hlg+9Gf6KE19QfbZK2vBPR+yVFbXk5KllLynsX/T+FBFECNpgb5vBhqMz/b73io+PfHcS7BmFgPJ
lpEJSAAEbRZXmfnr/6xDjzOW9aZvwhZUqbUT0qKXA2QN/NHdrZmKSAPkMCz83ngibxfEAL77HTI0
fTmYCuT7miCDQUG606qvG7XYkHJGAUz9WQt/9FwBlHqr4KY5rRaOb+U90/FlCWFhzcY1iufs6RkA
nKlshto7PDnujetnj1+CXXXLsbxsJ32tXK87vaBJ6zdUOcseW5adCRvhEC0S+0B6dV0eMB7Y7fUU
dsezdlPhDzeMV32ejZK6T6c8NXHNcgSVy7udXt8SF6zjgEAI+N5nTmewI9eO7O9rBFx86uNnZ6U3
5Lats5T3bJweMFpl608lXdNsbSRxpQRepSsvNx2otRWuVzFPYTArkqx4QYaw/g8Tnh0tI5y2PYkm
5jmVBtFyOAngC4qvOAe1Hn51fq2ycFraJILNtPimii4n4h24znFGh79wUz7gxGJIeY7gPML5neek
bKiHrZdnB2ffgKI5hSaYyA69LS+8lz+XsWW3j2lDvLvIQv6Vw3af/bjzKfJSlHrpZpoZyGeZFX/1
a5WnViHR688CwWGrUr7TXhl2aqdweMOokPTpZS19twtiGi47IRcA+UMiDHPAv3VDlv0CUPsD6+WN
bCa51o+hd3iYo7RvGvcMLHhuyK2s7tklFS4RmnfbjyCpQw5nqhrTwa3rUCaIiG+IvVAikKS7V/9a
HmFtyzNac53kR5xxzTNPZHkGPsyp2JwqARp62uJPepidPcPendwqMXaDdJDlG1Izlabu4z09dkY3
rPq2OTL4j9CY7AX/7RGGAsVTjwNNgdr1ADQAQ1hwQENDF5iI9l7VYF9GBOpB1ckGwUL4qsUC0aCH
86NwwVpJZY8xTOU316Sn/AOyFG58cMo9XcG08s0z783OMPfbjOdi2iys4Tu40UZj5tCinEQ1+VvG
tvHRfAqrSbkpkq3IIFes1hfjEFEEXb37NA2yXadDyu9ukvFTlOa4fKMWps6UeVwHCbJP9mtYLjPq
0shG4zlH/lk6Zg6t722lw13ecYax1yZp+KIjxfz7595B/nKRzOpu0q4qAoudUuXzWD3RN3HcrmL8
RfdaVmGo1w6+/GCKlVtCuspks6lS7IBmFxDQXICtzHs9T2JeplYu6r6Govw5VYx2ka7EwEx59gsD
/dTSOjUKuzQuCBDkcqg4vEQI7WTc/BpMZmfJ9lwDU17Gpbl9KV0N+Pqn7PMbjRT4GOuJLQXwKKNP
n3El7Qw18nmDgNIo1bLjFRpIqQVJ5XpS7fQCjMb897GTDhorQ3INGwOaQ44eMsCVX473Mc+pcxFg
4tV9I5xmTYiHs2P98tbc1rP+veK2kNfa9BYgsQvz54XV6Vc0AMNTrE/iwIS1AZwl/ZyqUvZ+MRls
4GbK5/mxXfEIaYuqvL5tvPKhjXfniNipc9ffhAw1wNx/fzKfbDd3xrUElfb2zXCgvJcRXfVpcfb9
h/ms9RU8WXhDQEL8z9G2MgOoaSXtL7Il52rhP2ixeP1RlPADCO9WhPf6aTugNvDetWdCJxT4qz+k
ILLM3AybztikrjAadKFpbUmeI+Y8Nz6aLIKRyeARcUc0Kb8caXp1r4AjDMBMHiHFkwfzhWDfHUOY
YAqTU+lncI5LuwzgUobpPY8wU7fvILXVR/Z+ux9EA77YcvUUHGng5ELvvgqkjB9t/VKP1m/XFInl
pmmtz+9MOOFB8OrqLdtcRBr46vG9rYnWVY9IL5PUJqAsKPjK+9bbxqNe3tOq0ZSfoUmKAaF5ZfDL
CfIKRzQjqXq0PfVkCvDae9h49wrylvsNSag8yhfSAq0wWr4q//BBu43HLOQWpXvP649Zj8+shY8P
lumUFM0SeZDBVurDjAUKD3+xKKvIjrb4zHSr00yZJ1ikhaxZqgZLQUkYH5HZafmcpD1RCbXy3QUR
hWwz4OnBUKDc/dfhJ1DgJNfstKAUKimpph8SWPZUziVbLrysnFH+GE8Q/VeWNSdsNivflKXjxIcW
T0qAygEL3Mh8T8DC8pQgUYwEOjosLW/B0qczqQRfzVwC6fnSran+5QBFkqvp222wOvPzizdU8bmh
04Ya4M5dJIBGFtw4mKb9sGAgCsnkmNxDrUCKu5RlKJsB57Gsq52RY5OTIgr50PJBWEvM/u7akxul
k+UvkA/bN/kdSjTZRj+fTGa4mHAyLYP60HZ4kw+JOkuER0EaXn9hq+6rp4z7K6J3gKwHJCT5/en5
4xJGyZegXDjb4LtStnrVyOkXWfGHT8imoUyikycdBG95UccPIaWWJSip20WGnyUIZZIRh+n8V8LF
L6A0IThnvvWIEhly6wBmNO/IsELQ3ZQskwpk2TQN0Wqo4tDE2ms/pu8BWjmVuh/W+oZE5Hr0Mpjc
Ah9WQwRcghFUbNUHRGdQOVC1CONf+o4gwfVmajjuWAvAMSKh/c6e9cquJYfOlG9Mt16qwNrQNjXO
GRHDWOq4dX2twmEczvA1eEsp/UnB/8BCeLwzVHBW2I3i57SWC+ZjyD4bphnCWRA+TCs6A/ZaLYtq
8bLnIM2ZKXEKS8lCqv5oWzkkXUKrHdjASjH1bs0OctKRduTitQEDTIRjj2SZhm8v4IewBvRj8cFu
z9y8WUmwRr9PzRQuumu+KaliVKCA+gEmzRxhYH/Odp6kR2psD1qWgQK7Tow/cnHEh+RIKMMZQ4v9
2ItA+3VXmKvlQF56mLskptttPLqwF/Vsm+8Lzed/RLDjEwksPla8g5uVrUzM0EZiBNQQUWX4z3kH
pXP1PtMauDWRA22Vto+3KdmE5yXWZjn1CVx+aPznYiFE/FZe7C7iktWgEKYtbkCRolT3u7ZAXMF5
8Cl+hySEAi+9nIViRYKwIeW4HNHdGOSTZWobOxAz0rBw6EVdcxKlq7CVTyvS2mxFje/4Vze9V7iM
fXWP7gH7NE5BGk1b+vYWQgYtv1uu5e75tDsVY2svftpDVHI+QUYHYArCUV5cNg0uF3wTozGQvV7E
0Iroyj2qVpncvTyyoM58nrW5MsCaNyQMPHafIk6IKAQ/NOQ5Mn8LDq0Ap1QKAdeg83RyGmohJaw8
01i2bXlyB4d5MF9jHtsLbdp/1ffWF5hVx+y1yozW1e11pTUyOXQGqoo8QrOI3T5Aq7QWSvYJflBn
epmplUOMdRGeepugxEDT07koB7HV5sBom60cy/odRX5knRmrp74xfdjDv84G73D3LAmEFmwO0/O5
gXXbafKXYG0XJU6nK7TArsUJ4HihxlCcmM/MzNxPE7Oco//DmyvdBoZ4om0vjNfdGhYhhKJzvL2P
4ltXeTVQ1Bvj/A/FZVc5AeEhKPL2X9F+3EaIThqH7bzOMVhBbRsfSDz5ux7mU3aqVJYzFEp+k+Oc
UbMuaQNshMgrL3PK3pKUG7lUkiU3YQiBPaifmQr4oZyik5rqww5hZA1+BC+TlPy5cx/AkXCj0tBr
TuGWxyBQ8l97A2fEvAqX2GS7r62dnGD6pWTUzUd4DOE7q3/VhKaFGuGXS4cxSOs3m1miclY+RSHa
C9apbd0MokhAF58pilxmq0kexCoUPE8TCvmdM8YIuEDs3BvS1w4PjtkkoF4F1wtFhhmuqPT4/jhU
wdbLDaHgDE1NUlo502sZxHPxa+5QtbSNpUcrgs5E25f3JTeJAK1nt5fqv18A3u93e+QkAJ/6Zkja
KKlNMt/fLI2NoaOz0MgcPkabuA589+8o3EQ8hihgSP6N4T/9etsy4bg2vNqy3ioMODn51+ZZVmpB
e3wldwtL17UBIoeCwjOjjYDOkSEBefHIKcpcLC/y6qSd35OsWNMVc6x42yE8YC3r9Gbfe/3grZUo
EoRNCLVG8tIEh35aF+qnKreZ5k6egG3eJhf5XG9wwih8B7x88x8tkTYuk+UaYn9Wi1Lys+TphB7P
izRL+QZH8wXL4LFdHKF1nKXFN2b9vnIrU9XKDAQBBGR/zzmU0unbrC5nm++BCP3nayrBOYMCuCCb
jf36Ds7Fltv/McbxOokpQ1RhfSRNijtAYxhw2RjyY0jeOqy+Vr65817KmSR+jnsjuydMg7U9MMQd
LMb3h1/F4zfnvBOs5HRFESTHlLvZE2eqtwR+Suq31Cx3s5Fv18uGfYGKQOQf7QLPqExb+pMTWtwn
g5L/LAYZZ2jWOtXOQX/JNbywNXX29gyrSFjBLy0lYgiSL7hLD5ELML2Zr7wsLWrhO+d/qcFScbz2
meEqIeFXfRZwpauum+qZYeTnr4dMXXhNbGxljbaOp6kZl9zgY3xACrzObrtRi0aYvraTsz/LEJAe
FraR4qlml8MzCAAR15A3wOwqHoKb5g0SiAKEXIJV1EfSuCXWE7V5MFZWWsk9lMRiS5czwmBgA7eW
dOOwG8xDNjxzABVXFcjSxPAlNU+YxcSbi9VuWutNj+wwiBNacOL9byNbwcrbGhuTaqw2kYeoUWFK
zSZsCoeQ16DsXIqiNR50t3rRjKAuoRgSDF9KuhLAxRUt32IwmELqU7WiD1JCZBqLMvM61/1TyPCf
XPGjomQSg1v6LIK8ZNkNPfNExa/2mIZoC9uZq5vMGyOSvy3VXFBRrgZMTJN/CNjkvfi7UtMuW6Uz
wc6IttQjg8fEg/tGOlUZYByEoBgNYpb8aH0UodFYCGTgolS59p5baHrSyZYZm5cOuVZs/sazf3u6
zxNFwdjl9YH9ZjOcyNm/hTrkHWQt4prqTvYPnBrmkVpM6qU8lTs8bj0SturYhTzqrdr5WfWDj/8m
ei1ogT9wIujQmafI4L8o6/XQI5se4SWdt4iI2YV4Zx0FLlYUF97tMuMBW3tBxX8gi2Iu65ILWaVx
HChVctlu/vJbkzvJ6qbv6oHM70o5bJfMA7bnjIdAsMlwjJQ+R1AyoykJGFYyOCgJOoYz5ZREGPgJ
OAm5LWB0scgVKRSMjX0MMmbxIXs0svKQEjdnoAAdSQs00pZjR+h44B+xsF7c0GincdfP32fdX8jo
t6Fk1rcV4RWdVOPmknv0l4JhBMKB9rrX9wDU6dg7wmj9uJJZz4bUdmhexj0YdV2jmR9bTchyDgZQ
e806IqbN6qTFi1JWmkSzYPYsbxF9Ye4CdrzhxSfBOoLD6mhKxTDFR/dA0EBQVqdT+i7HxEYGgWgj
mnW6tJFhN4dKOpbC238v5Pt2fe/4Mu2qne4dq8hL0fnVkacq5Z0KOBqDl3MZsDgU8lglMvZ6n7zB
s5PaZlElNByjNvyBGCNRDMrCOReVnCp+tyyO2his1E4OO+5E8IxCMy0FCFJNA1w4yge5dX0XCgi/
+OBtQda4GKPNi3syEJIN0llb0p3sJe827HiBkE+TWBB8lAJGYMprZEDpc4Jt3W7goqLcanPPDvxf
q7OpNXoEv+DqeQfOzjLIfm1sLQAOCFU3908hFDrKQoGzV+2M5zEFihYZteUap0sqqhg1NkZYHvK3
P0RRBYb9JHwQ9w4hD0VHi5bzDHS5sXauTQTgZ0yQLhoSvUi25kmfkDIRk3s+ouWixB/J2AQng+Zn
mYNpZ4ZeB2lZOGzzYDi64JU+O0FMX0CbxDJkIJwcY1hssA3u1zbo6nezvQ09L6oh19Dp2bo2iwVu
sT7dU4Z2PfUgTNqgmV1EVbeQIy8+tyLweGEol3af8vS6GzL8KeKJaGm7zwijmRM7N72D41/4UB32
VmenguLzyJrbRZtSSCAq3GAymSoVEVdCBLEuUQyoa5Cogj9oCxwB0yX6T9My48WoqIZOV8EVNbmC
yh9c1DCLR6fHPZ8XgK3KMtPIerIj5DvRwBhOPDd3/tch65gMsJCletVy6ZTQwaVVGzoAApzBd0wa
nLysxMLGHhgzeIkbUXU/AsRO9ri7gEU3rvDIsFucU6ukJ+ijNF2t9fWCVMUMbc/cZyETSiHPFLo+
HVpZWVSEPTQ6LUVqiO7lZfbL3t9M5hFhwSi1+SJIXUctNrYqCyQutRsn7OSiYXzYOQ7+wn7/37h5
XP3jCjz1nJZgd4gVB984SQ6A2EoyXibn+CoS2XzGXQSKy6NNBZ+vYgTaBfUZTxzYb3MRnR4PkNjc
9imcb63WmuUxZXGqR7FQ/ra0iGlfRJ8qww3OwU/5LnyaRhl6drQnvDxmz6LbCYyclzjkC3wg9j2X
1U7beJnpKfTMy/I1fglk0sF8k/ceK+33HKh0y/fpGSuvkDahiBNBqJTxe1CmQ5txnUtU/GKLgsBa
CpCL6Fbop2kPjd83Pgrb2JiJmnB33rFV9E4wFbLSuUMVDJVwYMetR7bOMqTY//0fa1DZDznOGGTk
0gto+O71jl9zxRK/Y6szOrZd5xu/tXHMoBn+KrrfX/8CE/wcID/RjMGTfd5cLOG20xuFrg0TuY9I
7SwMbYqULl0onuAgKyFRtsIBt4JNZ7n63b3hXiThkZfn89Jik4F3WbhgNHEzfnumE5x8yu4af2no
iTGYl6aKDDqDV34et8JYXhvRxqNSodDEXxgzhF2QnqmgkRv+zDIie8sWVBFYUYvfEwW7ghL2oV78
zUrCyvn/5CPRjbzF9VD3yyLX8WuhCy6I4K68+6KQF9eEJw95wWQS5zng+wnHVvLLk7ER9H8SXgcX
yG7eD5Gb+G+DC65D8+7KQCy0xLzAEeWNSYeGe7yeDA/skQw0anPAUZciYqoOcb9gdOEdoIKhOwzV
nrQGu1Plcq4u+IZk1xpwB83JPIuGK2B7jOCWc0FutPDgiIXJjcc3F1KrgkX0eVrbtEyPbUi6gBRF
LPxrXz0VyIdo2UD9BLYdKg9UK+DGbNwCIWpeBXoQHq9ojBqZxZ+HRU1tTBzc/MhCE/TWU9teS3bK
cKNxnDaXx/nz5+R0aJ7iuacDEQq7P04Res5/y6jkvwXEVmLhQnFtTJIreaJqcGUT5drCrUwIEncH
3UVRXhnyr3KegiiiU+H1M39rmSfXuFuGkiUKZv+62oKSSr4VsDT5irIe6Xg+f0gWSkrMpNxUZvAt
PmCtKSDtIgKxVub+L+lk0V18jwOCLmhNGfj8B3ZM7h6IhXk0nrvb5Pc6ad6jcTel0J0Lmm1u45jA
+boIpIj5khyEITDxfhfKyi23px9lrhwu2xskErxeTuANfWv6OCNbLLnt0Gogm7MlUth9r5Sw33NH
3EgMsWHEMJR+OkaO3H7naQZEVv50QNX42MrjjU+qRRfnTaNzW76LX+OIr0nnjN82B56tqB1uQmXU
xcWB/hyE6gMO+WF69fUNrClFdSY0rz6fpRcgb+I7chVFWJ5NGhKPCygBQ11meYNLlOTzdSDQ6SAE
QgNL/rF8Z75DIZawk4rqGfD6cj3agrt4MPmj70h9c8DKuZ5EUusxVoGJLIkgV0HtWgwFrSsHYIod
qz71IWiUErrX7S1kKNoa3V7K7Yn15/uNYIh0O42tRN8AgzzVFS+7Nz4mf/QgmCazlOv7bQIuAY7z
QvUWyRTNlQznBjlTwmqw38Xi+vU7VPweSYJWys3OkwrXDoYUMjHEQR3Vhm7PW815P+aL9liSe3jE
edy879/a1NC12Vy3UUx4NiFjOzondig6XohbQjlX9Qx0NdqEOdtNcwpxEcmn5K9OHomLIXoifsVJ
xO3nEcM6kIuud6ac3/5uUiUbeZGGDHiG7CBpNl/tHlP4uXLH6lf1ZiMPeDN7d2chqaea5MwXXl7Q
RN8Fe39sp3B7/hvl0NllTwFrQvmsuPSAEa43/D1oBAMzPjojL94xg0BS0o18zs+7pVunBoq1Lr7g
JZ2iHBKZsJPlxHAOmn54mYYWmBHIN07KruZHjf/xhCPwJrxmjn3VUFNOlX9MHFiXImmHiAqgstiH
oPxlXl2s6Cnz+FLmzkg1Ti7KcIasE4l9T2DIgDIPZ7B4+0+yhy81nF++lcJTdguETkGrsS8E8oWG
M+C/RMWQllplPoYCAlwwg/q+BkLQpw+sgvIwTA28X9NZXBJtWKHF/+cbeOfcPNMEArlmceEGhmFM
mxj0STSkAYew6RkIcYx3TeeZ74kfy3HcfXOMvWrBk9+nmWCK7BogCKNZyy7TzZWzJ8IkEtb/gL2W
3QbtioPe5Yup6rFk0DgRfD6CAPp2ENK75EQMqAIWEUtzNdb9rv1fhf2as41ltr4xcBiEc2lnh+Ua
GT8Wq7R+Yt9lWQPqWder6CP/n3XBTWbwtPQGK8BvrX+SVFvPuJ6Pgl/+QKNLlp5YJPGx1BIN6cre
rFJGGM7AutXNLEzfcm5Qzu59UYT5KymfMg8jPF4dAGJzMX7ts+LoI6TJ4cc+KgNBxqTetb1bebEh
sTX4440ovIPD5eiWkJfvyCb2UgwznQWNPkaL1gKkDJ98erMk4l5GzNKhLWPNtTZ49ZU817xzKBjN
gReZVYeHZHR9ZCvqrvUhmBieFxGU6F1f0JCWZtzwCV6beMYGyYBq1tbmkFx+I4v9ACD03I07jEvR
ChS8JrPiL1M4dr2iY6ADkedYhqdhAOd73Y+USVqzoiIppfxnn/dy4mhxd0/LgTU5GAZeLDmHXCft
0DaXfCbmLlaSbkHsXUI3/s1b3nqqBhh50Ty0Wq0VTDQKIE7pmgyJ/nTScKii1iuO9hOpu2Sy/Vdi
I1jtWdIMNlIupp+VmcDn6DAZs6b1LfBckfu/WmYAoeznkonIEpomVavvPDDVH6A8vTkg72qpx5i4
e6FTyugXb4ANve9RStzNWqabHc9TQHA0gg3ujTV4LfBYJZORdX+5u4kmSnwEEPhgVeplx8zk+gC8
R6vuTadi3wYzs41636DsKiU948kVf4HBGBJkcsbmisapyCe+OntoqDdxBfm2ZYjmexXIOpVrVx8x
bRgYHv0Qvs8e3Shx/cEcm4yVqcIpndImUWhW4XcchZ1jN50+gN6j01Lx9BHo1DbnY3G8/4BA41UM
0bGsU+8Qt9j05fnDTlVga/XRhIm1lS+/lhHH0J0TCorxZ1fqjf1mhaDmzqWyooftbOvInvb+xgq+
qq2sFJrS8mIeHbBRdO89s0g2524A+c09aoNbn5tL0Cd6Me1sm13bxgXlmpsvgP/EptGobI5zfgaO
EtY6uAFRngSml1yMiDHbErC92f7WlDJ+1SD1Y+X3XIEZ+1ijw7jFqN+PvDA7kpbX5c7fNuwlox4r
v0w+WHBQHNzTIBCE1JKWLM675+WJZyZ6SPl1Q0dS4AlF8/F72AxoVnOOUO1QMzhUBXMUjCpAUMvI
2xh7J5sND0AG3nmrPbAQUs7SeVmw74OahvYNExsjLX+Y6+9OHnqerbHVejygJWd1ipGt78+l6Wz7
hlUd94lTnm3PlakKnfwpb1Ta69G5PjBvzOV/GeeTfyBldl6HImoIDMKI+48Wv7VQ4GbpWwDJ/ehW
uPjrXzXDUZp86haBaXmkTEjglavxIhKyNt3VIKf4O8BynXbHY/qbzJdug5AXqeDyDRX2g905ZloO
MkwExpX8GPAuqVseoTsZ2Jvdi6ZLLZCTXqlG8vkMzUp2h+I6KwcR9EdxhD7ZkVLpeGqFrSl98h/t
5fONYx530SwIpQumXE27xQgimqyKGY4dOUqx1aR7VMHJGF61+14jFQJLFj/vHL4PSO2bAePZqKzz
tshNlsMF8aPkEZJ823bld/ZelAztko18ymoChooWBP+KCFvEBP7d1ZQtQ2EdioStwYbLC9Ud/J8a
+SSb3uNoTp4DEVLk1231P+KG8yOtoIzHvYesg50CZsWgCxXOkQF/ABekxvhwSV/91HD/y0/2FNyS
imF2S3GjZPsuvKPnmX3laCdz0vsa32K3Yr3Pq/vMbBWFvXTsRoxuyzFqFDHgfs20lgueauDrfh3F
aCqPsTcZBF/jriwA5HfTATxiwLAaYTjLHgpJJV/QU7XklL8OV2mq7cWmQnZtZUEY5Lw5JyCGZPjX
7oqeLsgyAPPyCUODFVp0SpY2gSk/vFkRRPI1lcGj5yXU8oxPtXvztli83oTeHRjnCYhoEOUIUX2G
YlvBwAmMABJcVIqfUz68EtiKSFp2f1NeS8uF5bfnurM4+ksyD3PMvMExZzVycEsG/YhCvQ27UxOk
jmi+T9RU2v1ItZdi64m/CFaQqt8ySpdaYODaR0AaYp3ylXPo0ZSLfOWD9k3aFQKvP8TuusLVRbf6
m9xa6lNrcWlfhtTei1mMxgXRindf3EALj61+CrGlWPDqPghYwW5Z3CCVmsnjLRh04IFEEsIJr/eM
MKgIxF1YO0e8ZI/7LA2nuWVg2W7kWrMtwCoOPACgp8FIE0oU+ExyL6ADID1AtBU4rjDY1N5PQgfg
70Au3YDCpQONvw/E4WJ1RS5xTQnONmSpSahS6L8IhEJbTs+DbCFg20wMNDaXeZRhkdR/W6I8XHi1
JsulFblFMoaplEZTPojJAdVEu1MVdSAoBlla5Hn3Em/um6wTYdN6dPcHNpTV6t8gStF2GtaDGRnr
xK8EOHAcWa8FmkNI0x1Q+O0u9QGB1Y5QTk3msSZx7M1SvIdY6tvRQrEL1rNSkzd6M9dA9+YJoi35
nsWv1eg1mpZpG/irF2KRGN0WkxBEwyq9HtJCmt+rFcD9w+RYitzMmE+RsmDzkQOXdp1Y/7cLuWGy
M/vIEZhKA4RNK3fEevzq1XMxR7WNQ1I8qwgbV/ZMxg2r7KCO6qm5SGx8MluHTzLtVo+N5T4RReVx
LWqfvq1TWImPZCLcysRvx+s2g2F7tMgMPPhTXS02UVqHFkNpdRJPV7HjNo93rwEQSCnpPZBPHZci
xkKwiEd4Oe7AL9I66St0NcN+MuolnVqRHfvuTlu4642JmI1n8qgpJNbM9+LI5QtSU+pEzgTlyclp
fWq/fXnXkHsuAkqJnYDq/L8PPGfe9N51IltlAz+WBnh3e+XefxrKX3pqoJ48QSAvxDMvwfZlhI/0
xWwvFV3csCbstIIvGOshBaDMxGvGVGm7Po3rR6luEvRuiPZoFiXXLQoJgkVQflBlagC54SAYT/xp
GTmFWak366A3QKDj3X4tRXFXGaBF1PiWOUPR3BlUUvcH3En7j0GKnoeBoMWQ+HPSxh5povqAYgSF
2bucpxaGAY+Di0BREwHBg1WIe1PlsNhZncKWoIJI2FaYGNGnhneUTwGi0aWaf1h+AFmPW4VLG39c
NPS3EF5r8lYqqGgMABTOnR711+pzhyr5iyIeXU+ZJHSOeOynEE9qC0OEZQB5NQ2IiESfcHP95s81
fawcl8Prt5qdnLm8shn+f7bo6X1aM1N6OahoLcj0xzUHX0Z4XcIyG2XUHwU0EB0gnkpXp7GIxWpa
NZWXSZBcKfA33b6RpSEYv6Un8u6P4W1+AnyqG/j9CqlDArB5NUSP4/hMFKRcZUuyAhA1ZUdrIdXy
/9LD2my+t1hoe13/IXD+9SMyJeMxd+7Up8Kp0jEtPOK3o3pqkVUZWoHD5LIXjsVVpk+ErcyREPhc
Fa5jt6i+5cz/24rThY5iVhj4iJYnkLpo3lO1mGtm2znBA7IUvtt9IkCsw0WiFhPdqW1bVhP20225
tIEZhbmCmcOhtgFTk3pYsPP8KONVVu7colqOQ+gvEvn8bYRUrtRnX2OwMJfJdVy+pPBdyQHgSl5n
uWw+jE+A1CA8BA85Y9FlQPc61WXmUvhlYeUV2AS4BRDO6yNhhDKOJ0XIuIe7ekwrn76ppkDB3Q8I
7L0x23ark+IPIbR7kSGm8HTWMrv6CZoDxGswX0IcdFBK836QaWi9qUtNVWIu3Dmug8n6NbPiV+A8
wT5xDA4KOptAu8HGC/AfokODiKuMpEf3xo0973UIo0nzgWxsz0TKbDu/bH0oaby2O1G8hYq8QaH/
sIone0bsDDQ/i4ssqYDWCoyhxjY1BL+vwiyatT7qgVmPSzbt+RkhrEG0ZY2H/AC4RdKVFO/PEf7D
sHlbLSIupfVQfJV0rKcrxr5B0k2Lf5hawm2LIZfdcEo1a5DDIHSDFp21FtPRDl1xKZZu8OHfZHyJ
eA6/zvlABUuaojIhmgx6v+AOjTKBSoA7N7hbdFLl0zyed+FGKm2reR9XKhIYdqu4ZS7aOMLBMwEP
u/yIhIzONonUksyfv1Wn5y5Hxzzp9eS1OAXzL78fm9eL9J89uBnTmg2Z0klDYRA9je1QcUmtwBQo
hQ9V1lZVJ4sPBwEhMzh6rVDNmwqafGt8VibKig+Vq2yz37UI6DMSSKqfooFEvbRcqRDu32Nymqnb
ftDherFlwogNlkncUvF6h1gaAnH6XLJgacTW+kpgNgn1BsQXgFbTts6/e0p7ZY6V1GY4iKvQ5UrQ
1hNMydwzPVl25Q4GEV5h+fdGTebke41rcRSKY9/4kcq9v9xoRDVBbPr1V4FNxNYg0vGVmVCV3O8z
fZU/E390Lr76UofuFGSOpT3L1C5+o/WXn/dYKjDTLxOqygwcupduvukuCtwyJvL9gls1NkJaf5jJ
2ZkrrQGucvheNVVVF//T9pSJbcij+qiIcnZSxx6nIsVNmd15uPps9ZliIHFb8ue3tSw23yzx7Ob3
XRWntjkJmKkBjovjb5m58YehJcewjQk7EjDBh9emfcGIVpC+bBphERqAzR3oyL6FBqaND7VQ1KEt
gAneXvWLwrHtFimymxV/Zbwp2v6gB/PP5yMhLVWFX5DlRch7i2pJwAYNUtu2wzEgAVOH8wYqbat4
aIalEijweWEWieiGfo1K+wMN96llYsIPKOcU7VgEDXF7megfqnroYdmuD7QEVhqlJwZxMA0YUExy
444CJnv9Wk3+hGnrIQPtLQbKoNLXo/eQY28j2Rq3XUG4jnZS1oXUVqZSDJq1lAC4d7ypAryOP1Ix
VrfoOYlZ1z5ivaIZjMrla5FX9NkR4KGtypGJk01h+56Adx1NFqu7X6tEslV54WuPOiKQDpS/8WvZ
+OIc6zlsLv7xl75xZfmH1iGlp1ptv0hazfD4XrOKBtJEGlXbqODwHHe0Ey1nlZ984UxT13NRwsaO
IQeFKLYtxu+eb1YxWMGytWca6KqsRoRyh2YqtJs1UmukdiH8dTcnjRmusX5jgXt/AX4gohaJUJ6o
VMKEp2PMVACDh/g4HkxzCL9acBbJcZoZjYqEwCnAC8mWJlu2XYBahNaH9M8tZ5gAHAhJFCeR4paQ
fGQBK2wLZmPvLKbOGTDO8ovVriErY4O0v5KpihIh6bM8+CcApIphHQkrFU1u/dF6Wqhgre2IZHod
FP6ifoH5qx3Ptdece9TsUC4mYdi627LJnCZQQu48PSx0OJkjVQ+I5matJug3HjrZ/erQQCUd6Crb
jo9WrvIsJCgw7oXYJwNxBmtVypQRvDiomJd41KYZMyeA1Y7OljlFieYRXGwd+In/NC232OL+nJu1
55eBLoXeHWXxaIvPj5oM+6Ny4wIp4p26FZHXhYfR6sluEpJqmCK5Tk7macgvpOIDxMOVjdigzpZJ
jN2zhiqR355NDFaDE5M6ogXd3dF61T77arAUGt5IfOINDrLvwTM/15TLzY52Qr3NtGN1whMvj/93
qofcJIS6dKioDPHWLPTy3+DobsqnaFpXIWzc6gydPmttoXwmXOiedSFOaSkEvR7TbjqQrn/q7t0K
tVHPTXynWlaEqUOSdUw1Hpast7Fku3Ag138mvzrb/cQ6GJSH1lh83mSnTTYa+yrbdM3zUcPK+qgq
kl+jYtIPEaecpfcKiudaGBSbvVgLdJ+rJdCjQjyRUS7mdJ/X1VqOOiAmMhZQdf+IbyHiSs/uZ3oG
zZwE1vL6GPHDJ+1u7Z59QX5NOpp8IkUh7YRN4loIF88XjZl+0QfjBX1QU7uDZzt88rQtxUzCIjKt
hGSemskC+OFVsREPeGEoodcuDdI2g8LabK6ej9/EWyR6LJOlYDdyV+iTs1VYWVhnHIneJqcmeLA4
kReUf2qnmY3Mibmr8/D0GuurHkPJyTdPTeAUcuWW/hK1XkWZsSId6hm60mf/3HSm6zzVT1oQ1Wyw
wZtHLtn35bYzVJoWxjBV/rmCEaKX7YaT6f7P4P44gHgSMSRZuemcG+tZbXx5yRq6NWqlGaAbOMTe
ct7hkQARSIlVyz6YX3AR55fegnFvnGlhnW+eiwA4nOGvwMCBppkKtZscx/bu8Ouc0d1D3Aw/ZziJ
2RoJp7n/yTCOZdKD8hODzgd5GarmzMNIWqDGW0kqh8+K1NGy56KtVrd7Jkwht+C5g/nzaICh2UBf
fC8iqnNx5UiZA/eBaMJj6xIgha5X44YgZzS5SG26HVFsJEa8NtxMjNF49iyIXIDBbdNdePl8affg
xEXYqvyxzh9z1u+wbHX+AoSzBfYuFwL6HI6VcxGKcPlVVlnwx7Fu2h8n66najHBpZHe89WFvKhBA
IvZsmXiXCESdt8crJzoJIq4t9jvqcumx7nSH8xHvCWEfPdtFe6CPULdUMQuukQuzXHPoAnAnjc6F
aQCy6z37GR+TDluyQPZlelvTGobMPfTWO8pBkkGG/FdFS+tyMviZfjA66AEMa0WnMCO10LzH0tO3
Lx6lLlsF+Kx9a6VmXs4PKeiNE3J08NeCpuf9rzS8iSOfoYgEtWDHp/OWpcXCzdtrDE7g9NzOPmWV
UMgE/by6rNuIDGgmYj8praI44LKi5RT9NpZGK7d6Ns3y5aO2S2DpqTKwkXEKz8C7a0wrXj8CErQ/
UUc3IZP25L7Y6EXUefwzImj+ImXTSaUB62qI1l4ZI/q+cqnPEWRSvZx2a/sorcAqNCnMwkwA1euo
rBeFJcollk4BH8ZNQhhLDb+JhdHJSwm1TL8Ie9qWoyQsyU/t4hHYz44ThmOpqMugg0RiwFgW1Ll4
fstqKlIiNLOw/huXsW61qvzE/7dpTRlWP6xfzn/ClH7Q2g4B9+wSIfuZJQVpDTcqUN8+ttu9CoP8
TDXOn1Au7NZ6yotUEOy4pk2SFO0nhz8n45DICoKzbzKAhrgNz+lAdAiFp1Tg4LhpN1tHItlXFccd
NpseRVCJIb1JIp/d8vxdinf8A/jr96yK+9wQ9ENEXa3Vu+8VSzyfqL0fAqkiL3XNQAm98+lCl9Ul
22xntYmdNAj9c++xTKyIXVbWc5U8M7Z2DxSS4WXdz2RNNQ903iUNKAF1DHnmuduiZHDqLvMDaOn4
y9tVsV7x3dza4RsXhvNKWtf+R4s4amz8fSVN0j4jtPxYunGwELW8LkNnVlPly2VfpMpB2Ksg6/Xh
W6mu6KIPvroVsJlLXt9m4YDbQIgu/sRcevyNz5yHfTKHIoI5gofJ7mwcdTnhOvDRa+GadgyHgtl2
IXYErls/eDVCOEsuDNVZlJT1Ign+HUTxocwQXXLfWLjeDcmjxHV1rY7hc+N7vsxjASn1vuK6D08p
xmJPMWgPnzH+k7Lq6YGMI7w/anKePa9h5zU5F+u2yZvChIcoO3Pa9F/VqteDI+KhBJ2e5lV4JNcG
lwAOZ5EZOEsvPG+GpI+tojqpd3KWvtfc+mYmekV42FBRshBkkJGVKRobMn8d7cLexZeJ7n0C1V+w
v9OJFwblS44JFcTO1niqjgzckff7J+Kdw1UbxYBj0IvCSS3DkXsfhW4eyC2h7tn0V9nfMxz2EqAv
sEdVtHyCOrpNMR9qDMoPUVXQa4WdSh/4IOjqsA0zKH+DVwzAsxiNfzuahSVk+ZAIcpxnWHgSzjwj
w8/qKYl95UmGdzIXcbl9dbKc1olNpWJ/ALwC39HoZnFTqIUJVY718Os2pFxAmrNihGInNlR21zR/
O/TlUZe1Fdyb5EBoOp1dvT3UXpqoFPbMDkcVhreM1c5n68tPis0YnUPbwUntsjCC6onuGwdmLdBH
kY9B+nd8PRVM9qPVNZr+7OX34INrV6juQrzrLLvvzelOBS1T3agbAUFQJyo2D38/ZqM9Zu1JDeNp
MzeKv+dPFuEPoa13blYHW/AzKkqqjUn/jP2tAZIE263AMNAT/OrxOOPMpsNwn5/1kBrGzCTp2dG0
m4atDFYrGhVQCDTFYU2ifbnRZhuhicEH+ci1lhjqN0TAb9K5Cc+chuAfbfXnBPd+RsgYtrQ1o9oD
Kk+rfaKb8J8MekzGzH3K4ThphvqNjYyU7jf9uhBtV+qa6ZOodP87/dogtmcL+n6QIzA0kBYpd4N3
r8eZczhZNxIAMEcDJ+MW2IHiWdzutWO/LX5D9WEyaPLTqDstLw06WUFMrArSjzN8Jxt20hk2c6kZ
Q1kouaJpYnL60EfBabrYlrQz5W3nXKX5He/ht1SqT/cgvS0xptFWC1WNvseAOZjTuSVEm4D1u3XA
lyfOq6eft4gq39PjcWfia3I9POAYJUeCdQFLYijwd7bitpGVMZO0hrVnkerzX7cMUCH/1OPMeIX6
M7MwBKbdSSb2BC6kuFpl16F4TNWW7J9fiMH1MnsuiWVRXJC62m6Ka5M0QSYATqlhwHFszuMrkQnc
3ZBjTkSUlD5skquQP6AxSlJ2D4uLsFO6IHzbuGTembJJB12VIzI0CznyQse+KZrQyPoY5nI8RALL
KQop2Kb6p0ZjtYzALtNsVOv6pL1lRIUQwQo98jfWDnV0RicJXaVCjF+NlnDAFnSB38uVL1PNRE7a
9EfS1n2O+XFt8cpbcO9dk3VoFCE11VCpOvbebm1i/e7q6E8vLe1HTYO6G+PHSFY1woVemkK97ogl
gs46FLoitG1ucaGMTMKMfwpuli+EV7GY+wK/BnRO08hBKEeKnUEQUpiWMDl/6i3NlGs07/EgWx8m
bnJQ91fY7GhrRPHmLxSQS5lE7jan5MknEX2ZG3uM1B48/U8Pt5vm4aO0WnK/ant6kzCV5UFRVd05
eyXUo2pbiaof/X+EDrFhEZbZqntlleBMyYaRGSwYtb+W5JfMSMm+FWf8mHc7Ihg2QEV2sH8x9rft
JMhem8e5RIjlJHHgZB2uOb/RP8EathCA8AqeNJpj6KMPwbSdRkythR4i2tzAr8eVG7EQG0tASXFo
SNncYrmPWwjUJCs2Uk8PmYHlezTR1FW9nlzgegNU+92qi76/7sVeOh73687f7hJgshnBVk/nF0/H
TmIAsPnxxjRCB/Cqjp8F4MTaL68b9uzow9I8zmAHW5yIEnD86vAk5++rPVZJq9XUPzRr7qh7gkXH
//LzybQj+60AbXsDruXKwrBAwNhjxELrz7hDHft9xpHmdGcs4LsuXkhFyy7C/JTSdl5Fvz3I3M4M
+/oBVOIq3rRmfkyJO60j3ttlsIAz9r694aJ4/92mGs67KesDfsDqoM8mS/rJELrZda9w04XD6TuB
QNqbkVCXh33b887PgirAurcuXWJYVXXtOE51E0V+06u9UzkErNQ5gMUR2eQxXqzd24+abLdz1lwo
wtmHME8vPCXx9cC5DGlzxx+E2dLJVkkokJpwAni6Jd1NB49LYlLG3I8yyqLuyTtSdNldzRmycVYs
px9hHe2EOBHLIIlbAhhW9OomPWFwLTNRJ07bIT3jO7CoaTBRJkpYm0GlZ4L+I8UmVW5DIzdakZOE
Z6Kf0lbKZnQ/aQAG342js4ETFkvmMBeciX7MEy/48Rz896yWu3J/sifej1HlFiN2eWN7BYzfzx8R
LV+Lrl/UveOadCdrjKK8RUV1I3JEkrAjno74Thm0NOX0Xz+8bVmDbLp2QomkjvEB5vktFZMmFuIs
5uJGQ5Y9ZE3uYnkYst3Fu69GD+LtNF1p6PzFzCb2pDpznQ8fNfH39E1OfvQqq4FxCsZ6UTWC2CNy
XqmgqHqjvd3iHh1nTY/yFCPEpJHq1tNenPyRd+ypO+MhxGqz0GlF27YLpuzG9IhEA35DIox2Us2T
0gVnpjK8dHX1Lp0ks9GBh+EXbcQr7zPL05XWIAczwO0mE6UelIb2ocPMvauphTNIB00k5T8HtRS2
utaSeVLk3gV4EQoz6O0XJRvVk2JcwNknOkJxUr+JpxoIRHYuHBIgabxEYLGNJ8/LHW/gLQ8FBpen
Qnpf6L0FMr4ECApnKa2e28MhmSmX7TaPvxYYCagAeFonPkVb8BBHtHxpn+QQAcGCKgEJ3W8f03CV
KE2DYF3Y4Rh0X1fjfIr26kRBB3TKOXG+ShnxnzwVTYJwZOrdBIvVcYHLrIGKZnRKOjjWS0OHqLG+
6QSP+bRFp4c2YlHynAirbmY/WWTm26T9FwU0T0ZtYLuvkpH+MCtAQciV4d3sEF9vrLfWvIJDjEao
XncoL55lfp8Mn7YD6fuRw+/NOii1+ubuDhxGGolcCoNxByK77EK4Zd7TpxTRJjBLjCBipO96tKmR
5LWFJbxsMSRJzxEnX3VOxRqBwW8/xIESqdDUVLV6YOD2UolVAvagpKFGk5NXzBHxthtJMCSAzrtV
eR1jjhQzH7wYSukbPUUCUUgakQ0uHIIz1tIZ2d4a6qRUecLW0rNNl0qkkBzJ07mUBGI9EuhHj5Rp
wHCXMYkkzXLgSzm+0s3v9Qyoob5ccIBycAyOyn9+MHQwFusRx4RmTwrt5c4iOneCHfDht3rJxXB8
oQRH9NkQMawLXAgkrQbFZrjhLwFd6Ai85+Cr65XR8FkOypgJUFvz66KenXplHD9SAoeNl+0GGtnW
NAsIIhoqJN72vcWW9ltbKTuYi96qFo4hWOW8XF/QmVfKVVOqJUqmjMimHqjnc5FL06/tXBt8mNpI
FGpyEWnTzwOA/81QoMRiRqeji12kgS5edHaSw33W5+5yPMYLMsldHaIcCaeP6FJ6IPrB1SfarUbx
2S9w9BRmMeA+jMKwA7zgJciASQ6ZCFmlDCs5eZuoRU4RtSAV+8aOOAlm3pmgDQ2N9S/uELYlEy35
NUtbS6tfpR598Z9eHxaffv13bn3EmMAaACXz62FtUgz9ZjGIqY09KfgplDu5olUaC9IYAe1cytny
MGatwX8tR31RxAI8eeGmmAO+dAqXRhugjtNCKrSMawMELITJg6tfOH+OC4EFaV9Pra53ZFBqEjih
3NW0oKP9ZXJIHrnT0M1EeJcA581/2ROOJMjQyDZ59+Ie7FtvBwhcYNysvgP6LVw/A0I2YdeGYTTt
x/uGxZlTx44yffY5FmQ87ITs37mAShmEQvaagWc0gi1uoXTIHGY6og1z3tQ1LlCdLsuJXcEoZ4qg
S0XZ3Pmso7hRlhJ2nnMnLgPcP2oyNfJFX809yeIJAccOcw2EidgZoF7PNclulq9zpSFirBmGAXGz
gpa9k9T6UGoFvc+SK4A6mxrvYtOefSbPIvRt2Ao98CzEbIdL899eCV68nIxaOgR+vdYVSgKQRkTr
flvurqYUoagAdTrn45I2GBRRZeRwRoOpolWrOaXIfHo3yTiHmgDhNx8uSPS6YeMQSPL5RBik2eOx
Q+bw7HrB/X89+TStvibvS+Nb0CvUsNfexti168pZf/b+ELwtVxhG0a6qc59qyNVSDeQEQy8r09uK
nHliuNH/KOEyaOMir1CVCLmlU1itLYTMrImB4w6DXr/XDiqbeCxiB9woYQLP4WgPjXKejReVQgnD
5QYdI0bkgjPOcXBtyu5OrZ+Fpx1qUf3s2/7nhsyjdVRfx7A8xxiPdukQ3o4WsS5NkOlYRMOHezM+
xVO2eYANuhZX0IvAlzvMbXIHwbz6tjh+31CcUoAmJHY9v4BnyBgsh0TdiTrZR4Xhe/GrVlNQmBYj
BEA3FmJfxMiLgBT8M+VVaWsoJPKq3MSN9SwTxbEqy4hH92oN8dfldNhdHzCIsbnBH8gtMFXRF9gK
TjK/zPENEhtCZPFZGE/l7PRYCjoCtBv0QhY1mr+J1hirp7xcBmqB5ye1WwzPRLBy49s6Lz1pj/PQ
gHyE2DKlNKX4bNPY6ERU/sM022o8d+CAQEOXPZ81DO6xLpFLsxwq4PS7MkiHZv/6vIP1dgChOd9H
PjWOE2s3QXH5ec+NWNLd9kgSgRe38VfCauTIoICQGvancxmI6fN+VSOvZDwxRJKUEjZjR292byF+
yYk/0v4boWylAvnAVyc3swOQwSP+IhQmWf7aoeVd0seD92cU2HkETTfK5gTtz6qZ8W+EJXneObwm
E4LXz8h2k1HNpH0HvifynV347+S9mwahWlcbl1v+J0nS1quz/PxqnyJBfx26dDbrajtjh7sBAYDZ
0Zc7AkcIXntioPCY6Ob13p0iTZthcr7rMEiteqZK/larXgaEXnWQoZBZ3O5BJQxUQgfxrA8Q7fCV
/+9LBF1dTnCbNM3Qf3lPxnTmgiIQyo7aG21H7mHmHnxp8um5idw8GVyZz8eoEbO8kb+8iDDR4jUE
faN0GhkXT6GzY62XoSQPk0ZHpDlf0RB3yCIhQARICcY6ohUWIuMhwtN3C0z23J9TJMqvxYi4J+T6
XVy8aXcB6v4Bu8XdqtkzJL+2P1P2sN32M8s2CItnQz7rCqjAIntOJXk8Has9w1wEECBrMFbX4u8G
OsTbXa9g0butiwuxYGMOhmuQRuIgAn+T9odck/9b5aJOIvMec5u6Fo4TkjRoA2d/uxZivQJxkJMH
Rk/NaPuCTeZb+n4yKkx3eAsULhgSSx+74O0acl18grOss24t0xC5YWh79I2tm6M9vazU7ilEyxJL
pMXJxp+3EsQosBxltYZGH+kld6zM+ot3hy1GOyzq0e9U6zyEhv1Q9zkH+Z38YkWe3Xg2oxXg3gUc
i3okMoD3dRVBTjXuv5ouPQQiPO5ysD+px+uf7uJfwduulwnz7nxOihCxA/FsrCOcMT4zQi/FFvgf
NKs/nllVbJHMow58tIptF808twhjQML+1nWWEinNvPo44HS5aqYVO1eE/7zLoluL9J8QW3mjBVWc
0292oknEgstFRfudh7e6sLFQF4iCWRa2XN9fn+zJfkjbEy26iX+S0ERhxZqrbV8M54idDIRruLBA
7zWqC/q12ItI22wp1zcLIh8Wd84ju4A4WGmfhz5ahz8vzHspukFWNAtsp8At0ZVeKthCH1/MQcO0
w7l8aJ7C+wdf+kChUVDtbBrRTUfvdKXSsVZ8+9j0r5Djlm8utNx0v/CR7q1DbNQdH+4ZKhiggqgj
/jqi7sNA/EiKLzssbCc/z8oN4Bl9ugG43lAZ5XLKktI/SGzw50dpJ2Z1lbWnaXEjtHFWfLK/WhQi
d1OLFqpgUOr8DDrZGp10fa5+WjhCskhz05h/ZfuPhc6sOLjC1bMoie5u6B7l7xxXTiiWGNeM95Ja
EE7mUUVkjHUgBAwk58nwHSguPiaYhIFlo9d6jxtNjqrF2GqUdStAnMfW+xfGiktcw45SVlu88Jg8
Mplz5UtFevwr1kNHRZVqumPdHaHuh5TTDYBr7gRZO3rrihinzw1M570KmXAXZnOiavWcSV45KpF9
lkRcx6llwpjfK+LC3kTkveM7A3OOf/ULkDI4+wXUst/KWjc6/F5VcVE+2xS01gx8Id4s5KAvDy8/
Qwe1pt/eTr71pf98P2qPDydIns12VnEjXRs721E+20W0+V4zkE3BYUqU/Q0sNGSuTXXXalp9MNYI
KhORiu6A1JnJrNaz+6SYMfz7oQBfMV+g9Zjuhdw1LLkGpp6OJmz9FtZFabblbkI/qqaiTzVUN+oV
rHqRwjz005zjoSrnx481hVuVa2X+FEUUW6kVJcvn1XRsIRaAq8F0UiIQn9EJp6BMTsZHWC7ZM3sj
0EF0Bhy9S5P580Psj53xo16KqQFCFTVGsrNBnkJjf+mC3U+gaV5zxiUi6Yb+ZKuHnCY/0LDTiZf+
K0Z98H7o/7W5AtK/RqSV5PbIBHMBiGl4POJROzmF9fI6b4CEW8SlqUoeHxUQhd/Y7Kez6nB4Km6i
Ef3v01BWOXDRAW4uphncxWVGlEkU2Df+cgr+FoNeGk4l7id4S26AhoaFdHOhje0y/Kn+LtRZAKXo
zRbwNo+yCxw+me+1O+trhKDu2chNBgwQmfzjyvvlwlNVhSAx1vdHrjIFnCspk/wvYhmbx2/L0eDL
mrV0Rfks2zD8m8tX1n9ZCPniA+T4W9ULCoKEME3wFxPSR3mcnr4VpYo2MMZ+6ZQEM23Oq6bJzUuT
WyUtYqAa5q3zcAvn52q6xdqV2nSIkE2bWqqkY9o/wlfh3Pi5prg5YzrEtONxqbZtegZ4EOQF/mew
I1Zkd7jF2D5V/D4CEcYAFGEKqr/PlfddIwzUfURf/EZ7hXXNGRUK2WeZsOMvuaT/OFwsnuzYjOLK
5CJmwB5pyFBKgFlYdtXbVpOUieLmHpzC3yts/V+J+WruxpTdPgrj4UcPEB+ivAG/63diiHPr/ESP
JCfetMEv5nK5KJWC7mpPYc4rk67fxkZvb7rkS/cDhUfQQjze3GCZdjG9MPueu/oFIPYQyeg7JENF
zvYkPC1ciEq05APnT1jMXLEhZ5TiYuVR34xdBbllN9FRnTozaMVW+NkKZ8dcdFFcE10MIxbYs+OP
3N4Ksm7a8p3FQiMPISANIe2zJ7PLJNzT6tBtYf327bUy9GQSa3UypGz6XHRVlas8sYeRSlAl76Aj
t2a7fHkQuq0looNYZa71ZBmHLsgQpcjw9k+kyRAwmYJxjfibSZ3mmMPjL/qjIpU9qjtMtdFHoLex
mGfsCcTy62EQyfIxalVstBQb7O5XNNF0+Ut/fzuVvR0HAcJ4fXwjJgUw3UPFb7P7RU8Jl6X47dvh
MdUpHUQzycoW6HSaH7jFHqhK3m8MPIfVIP6VEVU0l+WRENw072bOzLs11pWAnsryYthac5FLi1XR
94si55xZGxhLeBcj0NMSntzSqXQavWSeo48TzYAnc5fiju3N/yjtTV6DhCuldTSBE16O6kRHQNku
KaKjD3Ktas5VO5n8uB88GUd/KUDRFzoaPsmhCmkvMZxLHQa8npz1PVEozitvNMK8uZ3jRwMauAJu
Lyd3VuF/dKC7kD7LdyC8cDXzX1ATFUgs30MugJoHbkIlizGHAEJq05WVYhesPdaGbMYVM6wsSjM8
jGekxwDD98y0Fu9ECa7/G0RbX6WMQ94Y3DPOGb9LPndyPv4FaENcG99kgic7h51+IZnfl1/KmL6F
9jM1lsbHc+yjeakaB80CWQM4s3fRgLaiVGwG8YimJxxmi6cA3u3xuUwgVrD2RnQNKgk5fYNmiytI
SIsdP267vNZnnNX6kP5q3/5zIe83vts1C30SgSKxu7vIZZB+RY2a5i08Rnd1798Bjsawa9k/Rcp6
eF22/P2B5N1TJEU0TUF+NDbOG7wYjb0bbZdm3m23ctybj68q1q3q8orjYeX1xjkfw20Dhbp+a3+e
hdilB73A1fWowLKDnyUlHuvRe2KGCnMOS8a2aUbBpXjeKqPKzFUvBcMwTGdXYQs873r6Stww2jVz
fr7wKf+DWC1H8OW/Q4WgQ3o2xkVxcxwojta053zUtXTwnK4VDkBAV/IxoKE800+T3M0MD8t28q68
HaPHd1X/w0JAJjWliMiZKM+YY2fcAnncDnT6l+3kZ/N+wQYrFSMUdYtE38ZMkxb5mOmEiEQ4JuIL
XQxFkd/uJlON7jHpC/Fc6J9g/ev2E2q1dDGBkfK24yLFrwUyLi4FBWUqQJN+FXV7+dwF4vnV49mI
XdJu48xg/VKBHIyVrw7uXVJ/g/qfMISH5fCKvABFOEPX24WFNHmCHn3FZHH+f9u7Sjk1OzQoslhV
oG6uiDavhcQR/ZOzcNZ+MPQ8Dq6VpKKvHz2kMJKCI9mHuiqEL4S6Uj8C30dHv7WP5WMjpS9i4OgK
ElXubvspIrs3ET9l7l0ac8No06KIt7VdDUHFlSasFSQ/eCYpbCDIuw9rcIhHE05YIW7rCXVIpP1e
zxYxFdb30sXegw/1I1QMzExs+aG2FLYNNE2g6EakT+7BLfmrByR290KyiKvnR4We+fMMUsoZFk+K
xNpl+OZ8S3ImHAm5LXa2hjvs6logn6IP0SHUNubyjwyFlU5NkcK7zzR7s6PXrleDTYNeNqPCh14z
PDqOlECch3REEj0/b6nAmxFOuZUnR/tK8M6+Z49RcaVVz0OZ9f3nyvns8zw6GzeLkOgeRAcwpOHO
s63S7+cKj8NGS93TvhWE8cVNw4OgRo7VIU01ftBKpvIA1ac2V9qT5XKNZnGs4sxNkHs3AVxFPS0g
a1Rv+i3J9YkyPvDI6hiPmLtLnQEmEXGvm9Va9oujAiKsBGH+NpNGiGT7d5G59DwxdgiNuH7xeq6K
Zwwnaf9wuSBKqyKwvB5jPBpwPav/bopJl5nB1fLVIOksj/e+NsJL0nVxxt6atLWRxqh4lAYPLlWR
PnO2Q0rxvoc/hdSbB4CYbr9yVMCBb2TGz7px7vUBFHDn6T46OYgF5s9gbaiihcFvXeGYzCYsWjJs
Io/hJlLs2b/rkeLIvEdDAfTvBzhj3rRhj6lBMaibECyvLn5zn28Vv6JSKHSlAAx9pb5vk62pZFFX
EAwUT71RqyjcN22nr8h7FSJEyqY38F4+Rf7lATd7noGG2swKyJWiHorHnNdxu72dlDsnK9KMaKe4
sssU/G/2/HmQnSJcni3EfzSQq/yxgywvGt8cm302pmQba+J9kiosSB9ksuiOHvY4j/rdeCJyrE30
kTh85SMdW/2mS53UZJkn8rtg7R4ie8/UXKCmiXy39fLaUbkspi1fh8sZP9r67tYLV31ZQezXpc6o
a91CblEKgk0o5VZ7ywS8sPLpcG5mfXrL6ixViG83ffHiGSNEow2hLADnWhoffr5l2hwMNSwP9SBa
dsnwOYslcM6ij7b4ulW3GhM45YJ0WgAx8iL8uZeB7slXe3epIj1c6YzIpkvsDjJT8iAkH7wxRbj3
Sp3iOaIsjsD2XrCLMJ7ycvzeWT/Tey8t7+7Zg4T/9yLaRhCAPAUT1zt4/KocTkg+qKzHA7uGLUmV
iNu9+Yxqj2xIluABtCZIIMNc81Dfes0ZQ4EHamhnXHc5NiiFy3/pnm6nBVOhogMLJjmtBkuoOMgC
7m9mxDqRUMNIr2qUdKGJkPxa/zy9qkuHFnMWAjPKZDdZWrYqNDTGgkC7ymc6lSQv7RTpCMMng7Ox
0W+NF3hlZT1xt06kHC9SUQtFB5Aa92JXeb09sb6VyFf+wRxP885KApf+VPOrwa6rgRrmCRFL6+KM
1DB68QEBxY2kk+dQ3UJLACsYZQRdqiQSFpyZez3yw5HTKGhYOBDpjBxckfFyFSepO4hnmvYIhsVH
ih6kN11yfljXLcDjQvfqoim37yNx0i7bYyNHjyuVS0JoJzR23pblbL5VNsSrg6RXXZb5Zls8iIV6
5E6huYhGLxRhWxLJCXMB+z4TCO9ihgaMXFZx5vcFGRCfpPmZRgxBWhusm9niODvycvvaHx9AqD/K
nb2BuSWj6pLSp6yehauTXoVpZ/7cY+wpqAXNJubULQT9mEMaYdkt+JjxI1wDBpfsd3KPlVawNUyx
WVNKdrhLdEojiTdT0QEWyoulVtO0qV0f1e26zTE9Bj1/2c80xxK82pQpe+kMtovek6F98SfC+YFT
QzcHC6KFqklmoGcek9X3xNnxuLE9MsVftFMUwj9KmhNzYRLDbdk8iRZGEaWqk8ctTH4kcdcsutas
ec/S686Z++j3/X6IbYpqOzqIzghUtyqAfWrEFgSWnlGeM91h81AH3tbjSpE33ckJXmkxYXrd32YS
X919LBMR1I5DS0XS3z9HXAlrKqGuCHmpikn7e3Og+h/8CbQQ4I+Itdg3ZBT0u3OK8TdyDXy+iGue
NMDkvK7e/J0NB8Mmw7lhHhdTHAhOS46I8fAt/StF7woHoH0fElxKGZbvbpt5sAhbfILV5zNgCezm
HucffQk6DlHPHED51JgLtyKDUPcWlzuujJVCPY6BIJZq9+Tr/D2WwEOGFJUs3KbCpMKDseAWnZnN
uP6LJBaAttBlYeWmoiQUQL3xKRj5TA4Vz3avuliz+f072o0xqhf6fB7ZvH/x/mukF68wE9H1abKp
bcKHeGeyO+8qzh3+N+l+r+M/TyYtEvXz6tBpZf1r5MLbvRIRhhmXCIlgu0uvcbf6YWvcP6ppyWVK
4R9r1X3BOY1CCcbLzjwxP1o6ODJeGZO5BqHgMc/7F0xs/9dXtKFMePBMDhS51JuvGQ5i5lFHKEje
dNJM1HuITjpj2KXGt2jyU1JWDiu0n72irfSSVaa5IMeuDPhwpMF20olbl3fqfpyLI+t9KAjT3hJI
33aSMhbwCgRC7mkwm7prxw8vFK+pMy/uFbwdcVDSgWA/7ovOKFb4nU/FHoC9RspyVGhc7TVSNBjy
BKTSnkQhk1t2jdjAXekZU5YbXEGkD7opUl1IJSj33ql86kB0QxMzu+4HhX0wOpNLr3r6t1CtkXCI
YyZWOF20CQ9MpPfE9yleRyLU+VhtCTkSQVDMvsVhZnseyTzrFRWqlJSM8W6OXTKCnbcVS1rVt6hs
O/vyHHSJ1wzG8Fr+3qjo2KYnxyNql8sDczMd0W6UP4UMAcKgdUQtBOYhNT9F0mb1dcMM0cPGxTvu
V7ZbOqHrYznswPHhD/Os9OKWT+ZQx+N0rwQ0GmpJO+izIpi9oS2z+Qk9XoqxqC4I8ts+Z0dyotsX
nevKAIEccAypE+7aw/BgWJz0nScpXNhsU3ZnjMQrqh3Rb5IMweUXAEUi3njt7E7Cb3kZYKZm13ID
4IK0wwbdvgcMajyUVkCx3BmnNW6PMraZNcSSOXdzEYW5Ba/aPaQcsusoSHv1eExZHeoyDFbspIuH
dWykfI6bVAw/8lyXbubgfkTp2ZrhU3r56w68RjvHjzhBesoWYQN7JB9vMwyyluD/NBVs8Fe0fiDD
a9K5JHw2Nk0fgRCr4B54JuhPsrqxAhBX6DunRPgQRYtUlnbBUXxeNFRMF4u6yuq9dCSGTa931J98
gn2YWBdmYetq+3zWCeB2xfB+2SFyDOveumORPxi2ElINul8wqQp/DEDk1uzz5IKsOKAgtBDdA710
z45teyNijYiwk/+F0TK6thZXec8UV22gmz4amlawafxes/cakbXbct9q1DBKun9dpMfE0jGGQ3I6
clZYq26J/QKz93LtzUI6WGusk3EKKqX6aJn5tpfZE0W3yi4Gx0BDYqBIu7svZ0KPwFNMH7KVqITO
OtaumyrtPxqKizuUT4II62D7MltcOKm2wCyZb7gSKSWggwsEILUyt3t/m+obZzQYK1RdyjpX1n6n
3zf6yVPHGuf1Huhjl3n2oJ5B1dmLD2lQOtkI4YVZGdgktNUjHPBSygEwhSmqhybU4+L2cW5wXHYQ
9TJB/ofDTimpDZi774KliXyvZFaQYI8HXidETgpFDSZKeuPEmvkjD2t0RnQhuMMptnIadX3EHlp1
lGsjk9xh6mgWL2GUesDcSDvFtqOF2lR02SqCkGSUs64CWjuLIyjSgWECgDfa2bpW1omWebmEtk+t
xTg77d0j6BBidM2reTRbdQarEMUGJ549f+hzmPq8toVRffUq9gd0Rq+7w+BMK0XuprKph2jNC4Gd
8/0gcTryfe5gxJJGLi2qjnOFJZjRIcsA1qpGlMnkBlS5wzqMXpfzYxyC6teOsGKIDn4M0Bbwnipe
B5v43oZFsgvbM6dziJ22eWXsJhKjs+4HUTO6K+GY49JLvtp6yTn9GXCTDtnu5lH50wfvVy9JfYI7
dMC9Cqwm5U3Z8L/zJWdGIXEebkMfzd+k+f6uyhvI0LddHgpIFVqs8vn27bfxl5hgi57I9uGuwTb4
sf7eBAueGCEakX6Cj6y/FgAV/x83sZwUfwFV0ui064RQdRyNUvzl/ma1owZjrxFA+nTmwc0xUQnI
x0UzS5Pi4KNjnMvqojJMCTXKmwiDx4PNT4DdEwgfaWGOtr8nsVjqpUr6meNo/3Z98i5TEk2qn5IU
0z1+ycPwlCWUjIGCt/c1zfRzsIoiHC4+kNnQF3gDVt+DS3D9WiaONA6vhV6TIOb0Pjt+LdC1YtEk
X+lrUHovKpYPlPWouGwX/8M3ALV9sAsUxwlDFlwI9PSqp6DESKd7y3pE1iyV+AbGBwDgHZPZ8X2E
xS/0DjUxb8ZNg2VnnE/nnjltrW8r9gTBSQYuJw3sMIk4ZNhxu6ROisOjt54uFWvpAceP4TiGdcOw
SUu8VZZGoKVH95QhBbryRD7KPzXnNzQNxcbjU9kNcCdVsFAPb3TvVlTYcxlhU6AfA7mUF9NIvqRu
XXUzwXZBKc5Blammp7gT3texPTd6+zz4H2WWsqi62hCTyB9KLZoQzxhwV7bJfoCaGEkvYxkBdkmo
W/mHJ4U5b3vFqletOBVtD0M/JHpawcY9PlzlAT1vcQ/fUFb1fCv5Wxvqys9+u2HtCgu1xnihEMQB
13oPbNGwQqKZG7G2/sDn9fLpDwPj7Rz8G7+FcUo6GaBk0BKin8YwVwrSOrhwFr4LerA3cjDClz0z
cfRmEl6PeYSH2Nz08JKOnnWatJXdK10GaCBGFZWOvwO2cOQaZwiRQG79sxM8JwDd6WQatXFnfNon
C11cyUv9SRH1DTsK5pHAsN9qczeDGFq496bgYG2T3Qpntk0mxU7bsRCk2yUVxVZVhIj0J5eJBVz1
3MiQhJdIHalkvkiiEmTx+t757E/wP3c8eeCHQJCAt0SEzdoGaniPND9ZKhMdW8gF8AYrv03glkgS
QFKOcB2Gy4XFTHcRxd9vedeFAz0xPNPjdHIvS5tNdNgv1OkaM6JqA0YtLySwHx0bMuFB7Io8a6a1
41ME4ssrPx0mHDCWJosZQxOxbB4BJDMGlQJAqSKNKBmThwykqclQHh74MjbSkRYqq1MSBdDWdBtq
siRbGvjVXrg1WITo1KKUdiueH1gDrCwoxlYxX/2JauS1/b6TqRJ+R/cyuFT1X1UWEItSdiiIGQ1x
vHtY1S5BwuKff0YINNatHQYlNqe/lvIlUDTbP5LePA037y8ZFi1EYldm1qTN0lfazsiOzffSW6Gp
IINAzCerUM9IgQA4mhOCLfyU+H34u8KKKobOeF/8K2l9CAH/99rrre5lVZj/BD+P3J2q8wptJObu
XSWlPKx3ox/Fu2Zhl9xOap1KY00j4anTgXkpU2NRucvpF+tiUjNPLgg/46U6zL6Zsc6VbdCGSbOu
4QgU4Hdt0Exj38GUMh9MPIALZcW/j+HyCqV360/iiYMfl5U+I9O7L3KYF0AJmpw6rd9AGjqqTK1y
j/CFQMa9NaEvgqnwOKiqDIFJG1eEXGOwI43sK65vIc/pGiSFGnfs5FQ+9y5cOXR3toXuGdetu8Xw
wVftmBl2jB3DkKWuFuV1i/Hy9Vk6JLvjdpuROHnJ6uOHMCk01RSF+aansTrX54wmqmItSHRQTsCO
GnOSWiWq2mCjO+oCx3gw56Zuu0UZv90Ca6WnzOoI2AE09dGo4hEMQHZi+NS9ohUOtMS3iHLNEyh0
hqG/RJKqL3N9LKWCufuMP9PHbNrZ8wZ3HWv4QcWPTw27BZ/v9ie2iTRbC0PVQBjNdgBYAUPZgS4i
ZNm2RgwaQWIBQJvxUWK0FlS+YLbDa6dVuZ02wvfcV5oAXHuAOYsMfyExNdC9K+7WsQnUPbBCmuj0
5kfmozGhoIc7OUJI1E3eor6RRNCdqoNMTaw8jLWq6S+6d8tfSZcaVxUSWCmG3o7bFWy87ZnEGemP
ZL48J1r+PXEXmuYM4vkbd2ERkcuczww2jrp5nT/9xZE6qKJS2aYChUvajN7arneSY2j62N6gRfib
n9v8xJU3xJo7j8gPeRaz92V0RxhKD87SnmDlq25PCoSLaBDIzHXJtrb5esIoTPduyxudZW20frro
lx9rknMs71+vRbv+tEsW5x+Nbk64zMrnmQ6PgAg9O9zEBjro8oZ953P8YtCjHIaPb5Xm4s3arD2Q
E3CtNZ96u107NivmHKh9Kx2s/BvgUsKxhRz/jThAxZBJRHgOypZANGCSasCnHdkGVz07RLEX4rlN
Jh4ioe3Z+5mzaDoLWyHlMD2E7VUdNaG4ezljy0kCUV2KHX7x418Smq2vHwoxzk7BxfYW7DL1azpu
75Z5gd/IdK4d6gxB0gKTeBxeRQVfkbd5EV+9GpxHfSELfafXcXzKt7hP0awbKBu20qpui06fslux
9XtxX1UJbpp00OfONh5BZ8WDo3Cu9UkXHZyQ3iJaHXYcORTJ2fSRwSRXIpQaX1qNHYTC6TD8s6Zr
8uk7ZADzhmmiXzt1H5a2tnc1I2RxDAU8KulNLxYJUqEGd/HQhyk771oFeAVmufnLJhaddj8iAf0S
zvLe5qvUUITVCSKi4S7j5wBN0EZXVjLJfBZpLQev9jwY7agk07n6fmp9SjkKZ6RO/Sf49iXGNlwM
i1R1Gzlpd3bRLnXdVrGbJyvgTuKHuAHm6hPAdUWDCtlYREOAstgsncq/yNFQI/slOnCLIUx16OV6
f/rQPMlulg1XcmcoQx56Y+azu86odh0KIuStMCn6CWFd/Daa2Kl7LpCkLYFRigSbeYYllqG56fr4
5lGafE+vobcfe75DygXQyQGVhHmlK6ISUNBm4owKNi9KVkiwTCCoTbnNFrXidGnf+72+UZGeHCeI
ltHpNfnVTK15B8GXsle+k6sz9wxCyfpAExan5VENSJxgRrxEgC2UM8jWWfYIaNg8WyHLLzFmdDIG
zOj9qx65v8lxJv5tj5maEzTV4mQnNJ5XMjaAzIbJ57zuCSSk54wK3ibUE3l/itulzS5iv0k8Ga8n
ucE+2ygTo0sAkNjbPjqVjsqw8MITQy3QY1oWfHWIxh3f/nkxQbI71IbVcH7pkZtWqrUxNXZrI9ak
2DK5vibSZJOCIasS8C8RwhR8ohIA8Zb0oYgegzfnSGnGMy07n09HuNpMlyaHSyOBD2Lj81Ta3EHY
8PPtS3LxIcKNlzmoJdD5RRY0vbJ4lOKRc7BrrXvaDUX9kcePyG1UTw4r7tbqx6zFHnLym5TYNvZy
0QGBZ0wk5cE0e8LoOcXr7sioNDrpkBI2wiotmz1Yke2aN0pXRSggOkKweEyw6XD7aNy/cUYOogXX
MdwpyxtueLVImuuy1MH/zNanSAdWWqXQzi9RdEWdqvHB22LC//KPxAniuRNHVwZTh7YaJOFOy8z+
64+Qciek435USH2bIol2f4nzNMgwOY9qg8dwm7YwNGe0SI1APq67nR+Xmu6c8UXnOY588YUxJ2nY
NKTDSQ1ZoR8qTEtmHZjDjOL0+MaVtVNbJfMRrdzV+TCmY72KGqaIkVs8yj2T+GiPShtaHWYhfk9r
xiAXLj3pkCXYXoDBwTI65VVuVuw8c2lHZBe9EWqFf2+lVPSzyn5imcHfB//7qAAXcnCvb/cSrL7N
lAc4fo6ucp+jGBIiZp9YkQhjpCwgjrl5PbumICwL42xVZo2Fk5wxmU4DKW2Cui2RJYkgFHLzbNKv
PdGCWpozOq4LqFoRugAFJ9Sie8DyuRTQpiRPY6GZaeZYvnacwhSD/AH8C4m4jH6kJg9lZmHUI/bl
ZWFN/YiFRkkOdDuYvI52puBJIoXSDQzBVMEmY9wM2QBY6qkB+IrUGgchF1ZZwwlsKijLUHUA50Pk
x9IJCZ9KHLytEKX6vKxc0SnRAwNkw56Ih7bJD9RKG9Grygde1Ptz+Xk2L+zCHsG8J7IqIiCdjJsN
RBESMKoVBSRSutsXcCuI7eb8welTrpisNJtI5I4RiCDIK96YRL533ulpeJkgtWcBrjDjlySI3/aP
JgGEFGfct1XOQt526Id0TV51NVlrHKDcAmQMwaeYefQGbh8EFVFplKUhoFz62Bd/geyBkFaJazbK
ijZ0UpqfIm7d8+5Pfw4nx4k4GnZDuk9IpjPw1TYaPiJXYySj+mvWh8r/0RxF9GetY0iwDPAItFfh
2dyJpcYE05HTqtRS1qUVsyiA5UKOAQhD+haMJZqiFyeA9mpncHSzlrV7j0Ea31rFTVY+bILripDp
G9QPFW/kHj/5x+RGmY7sg2qkDimowe2EEhbMkeXYcZEJj3b6MNJlyoFfpHmmmn6iwOFB6IhGtpMR
ziX+iJ1GthMW5MhcigWRrm00YTPM0KVFparbSattNE8yfGrK3/H+qy+zGRgoBZSXyFHAaVwl7Blh
XhiVRgoye3mTCHaun3H3cFeWHb+msYvCI9NonvEbwmUX8K8oIbtl3uDEP8v2XF4Y+UQfTYw/BACZ
0g8iDTkFL3eEDjDMrLlEh84mVVGtpSg1Ju+K0onucXXmnDZXpC0tfKrIJbOVdWQpuJq6FEGB3Pqs
GQheGQR6/ruh6QkN11xCPtOB5m3glUf5d02S4d4vYCfNFM2NDtUrrt5Hm59IYSwnsCj+6On5baEt
pAfNnbZXGSHLQDWGxWnM5SdcyTJOFp9N0F8hpazCQIRjb41QGdDdjGAtqd5kYqPSP+c9JYZBVXLu
NT5tjvBhvC3vWY7aBjTTJaUJdDxMQCZ1aoPO1ywZ3Th6vkB6zO7GijRUZTF6DvfR07KAlw8xxmIB
VgpsdwWcaxT4Yj08CKafUltNAJtfpbbJgO2xyNmiExArAebWXjilLCXd8ExG92y1uJksbwbfrXiD
iSg3XmcsDN2AmcYGAFMqGk7N3MhX9LlRiWhxMpMuguualee6bQR80i/D8TKU3W69qI2dl3bm4w1D
daGKYhz6bRLcRvq0Pb56TL1J08HrBSqceyEEelmKXjI2CYkyehqY+pXW0rSBOMug0syICDroyaUk
ym3LOhSPoPCwwlniQZbgiYEs7dwIjLh/vXHAFRWIhaaNY1Y/V9RTT1qP+Y/B6+j7/huqN80yeH6g
R8sE7WcnOE3PwaLfwnC1t20k2AuzDjz6qDOMrTXRhBj5GcRRKRg+6EVM6aIvJl0N/ZZ4B8vH8w04
GVAINU3vNFT19QerW9ZhNhGT0Vr8fPw4HZTJqVwUepcUGknYhpzurKK3NHAKPEmF01vB1pAUIPqh
8v+54wqJjVjBuo++DQW3nqwCRn/4XccGi2gXU9XBfI6OAUD+IGkleGY9vW6ia/m4Mq3hSUpFpig5
bI6V2e3M6szZCG4pQ5YypUV+bwTvPr3yMPRIwnE2ZTZHdtDCnwVu2vl9KyHcZE0JPmvHNYsZx8cz
TkYMpfzWPI1aAV44vhsf+XqgMghoFXzXempNxIDX/NojeBT9bJhnRCCQAFTJq3r/Hx5wZQS+/BRq
3LFaYbsUkSkBq1ZQnOJUIBEbN9VxDhTC2QK8uEFJWHi0AprlKwC/oS6S81j4imEMJPgrol4xy3/S
FG1kh0VTJnyeiLvmVfM5q79w2JJ4vDdfhSXbaWewDgB2LO/BTkoURSf6yjOkLvw3FXmoh6GOclAS
WLYHePuCJqLx0O7x2EUFziq4qZAmN42VrlXuKPsL+UUlf2XFAqI0qaNXpgDAhdM5q+nYzJqrSJzE
HXaEh5m9O8Gxm1KSKmMhYmyuIdSsDQBiv4rKcI8LSi+Z8kaLUlCXWfgC1imckzzriI5HVa1FATeC
wWbnSC6JVnprl5uJ3RHB7HXRIiLnPfrzymUN4jZnUNOWQO0Wzl7HS3LKA9a7e4gaxLLvEomWYp8L
ziwcy36p8DP3bC1qvtxkCEHgA4m1y+Mn/IiLeqaz3/v9TURjVZ+bmFtgzGLO93CtegZnxY4lFaGo
ahFeljOj3y8/9hF0CrIqYsJOBOzH8uwP5I41UeRwRTcQc6tV+kvC1lIzRaThIvL13bHPXLUWwsgN
NigwBQeLxaHSkJeo/TEugfczbzKuuyb5wxulgetxGeK9EQuUmYieU8tQD2aZp3CKHpV/votNp3Tw
wqOMIgfm+yBHcl6IpwTdtU9ltQJe0DKjDX0Q9cRLSh3n4qEMTzDNpMJjW5Vjn6o9EkHAw92EbKXd
F8hKi+qRcuLI/fhhMuQeDXLx3Le2ntZty1pyacCTndyVRMR8YW+Pgx1m042akZIIcrxodRY67Kfb
RzARnZO2SwuCD3+BdrFxOFOfmE5HKdnapHnfkju0IlRQbQVNaRb9vOF2yl/HlHdZ6PbQ0as+07yv
u4Auy4GRTf2JwCcLO43eBcK/iNmm4mfoHzUwYkhaVL0XIvOMDzUg/i2AMFHWKrkkZ+hwrOBW2Gbp
UG2bIG8/UAChIf79GaaQz/nvfy0l4IgqaigjV6o6yVYrAX7kS8YfB8YCLF29RHa24NLKMuMltUx/
FHvhtWq7Ta5OwozoRpuxsAnPebRJBNuwIW0QuzvSG2BLsAiwXsn7IA+raVdbZ4+8RTjHwRDmxa1v
DjwNNXspUfesGmJEdqDlrS6b5lLzHp8SrTkzs82G78OxZOuWTcROhqEYHMFWhJd2yELndhU2MWuU
qelqGQ+S3tTlIepW3x7009okt8iCeGsHkrIGJ1+zCj2j74A65vdQfVMHwuFRgAzqCewQDavFsk6Q
m7v+nmJTYkEsQTlz+oY77KdlDYKzlSSagwIozW/tNqXgaQEIzOzS5/qV251H1R9VAm6PKeZaQXR8
kKMOwdLUyjVdKwxk+Jt/yVigFnOjLTLV+KJQ+pUwnY5HCGTOADH8zRRS7lzVZIz7AFIUkjVVdIBc
RDi3rOYQdpRKwvaVk3q53xYvuYS0IxLRqfhdDPj4jLuFHtPtZaf7HMA0w0Tti699QcPypuVH/o9Q
zA3UXy6+n4L7T7dcl+vmMNuDLKvEHY29CH6BgBzggSF3+8eb5OKt0BEfDJhSSNKpBcfRBNr1bktt
Df5OhdmqysCY+q3HZToLK5MSVECoKXYQ1cd7VGT+Bb5wtFDbqIAxNH69nCzPb+rXzsaEZXCUeES3
yY0VQnF+zlT2oEGEkstkRHblMbjT/xq2dht62cpY3EZ5rh9Wt/x2Cct6QY9TMTGMHwrViuhPYf8t
mwpu6XhojcVwWOlFempKX1tv412ZnBOJzLApEmEcaAzoXBNUSjyt/saS8TsZRV5uHJVNtvMmCesc
n37NeuDiVQITs7s1tCioJMvsoItdmtyBVLmtjJ8revwyZMd9uhSNjcvtqxtEaNXjZEeboM9BLyJk
pScIKvmk+rAvix1vYEb9ayAjJcj1AvhiKuCSL0k1ZjYQLBJ0tTrY73ULDqaE7v1m6ySleEldAlce
eaXsg8EvrAZVt3k9Jr/0a5jhoPIyzgfBbT8cgCC/unrxqHLHSfU89N2n4rFLBebyNw7mkK48Bq5P
CFtNJlRhKjwj9KYWISevMJl1XBwS4vfGliUM8Zh4Ujljq6VyhPjVC/VDAGacHFqDPYxdBtTbkeDS
ww2dwzKJqruJHi8Gks7hZQ8ZJJnTdAvlQ4XKsKJS8prNS4u40ReFBgnINyqH3jmdrxAsS2Wjbl8F
60RwCwkcGwjj7I9GM0DUM0xc6GNA1LH+TlJrjK+0xLO++fT7LBMbfxJ64GG3ruB1lnvPOSOS5QjX
MlsgC6X3FZOsFGyBk24nay2Vadn1yefR159sVcyHJPXL7FMHdcdzp5/2xtlnIFITjWY6yRne5cy/
RDsrkFQQfDzHSoKqWpINi9hkP9qGYlsfzE+KLJunamWdHcH+Jk4YVmvApe6pBadMduL9v6/0GdRS
0CIf6P9VQzxcl79C9aCTYhJ3gY67Vigub3QA0iwkAUU5EowQELjyEIRBelfh6KxIqhL6huwZMxmL
cSVZ8TnyId50TYla5iGDfSWAGT+duGS34N5htK2HlZABD3QKl8+8iN2m1c3c7Tj98wS3jSOBX2nm
qfxtCR+6bpZBMGskIsOkU/ZrYof39TqIWhF6kAywBdyFTsWTpgaq2vI6NryNazcqHd0x20tiaYXy
4IXil86Y+fVGVksSaCyiheXSoMDmdiS/xDT7NMp2nFbrmKjyHqX70IQkVSrhYvPCUL29aPcv6jg/
nZMpCJZVMBYylW6xHYWxb7ALwkz04d5ZLiOjcAhzDIDlFKM5DuVi2UQu+elwQvX8+jru+xWSAywb
/XKQ5WFGuBd38+8Kb8KvZL1N4EIg4xwuQPelJJQXZ6WryiP8cZKRLhbHO1MSOAWSNxoE/ojyJpF9
XsZr5OKllL3GRxuc8UT07vvP1EYbK93gJksxuybKH/mCO4evfdR5YIdkpyK88y+unEraNaKFpt0u
rsXfYbMppF96qHo0O+/seYimOvFTxCbx5DlECn+G8d4pNAmebO8xmwHN7TVDCXiZUba8aR4KjysJ
riZ35uEen+TtG598H27H4aURsz6mghQA3PEr1sTPDbgeoAha7o9R9q91O5IVFbeEL5qvfiQe0SXv
Bc5A+fncLPMOikqfClh9D2qgmAHCfD1fwihhe6glwnKc2mHmcjlb35AplV7FTSvsG1gQ8jiT8f0l
4PoSTU/FfDAN7McEoiEW5wDqgjIf+Cq4gnpm9aoHWa4g3ku5jP6dEg+pKDC+Q9CwDXNNLzS5+0hq
AAKLqDioloGLfwj9zS+Ana9DttvwwLFeY9Bf4uV223IAikb5bIZIc2KL8IC7ISzGau4E9AG/MMEA
fUIaMJKpIYINDvlcagYAEU2J9lTET3PX3gB8kiv669398Oe5m221yRK4HBJNnxKVwFHrT++mg0Oz
CFj3+cix0KOPAIdi+NUZamyA3A53+hPzBUbp4h9c/EsBNwFFif7ELZseUABcoxgCKbhMpEEzyTZH
pow7F6szTY4LA8/zsVp9v/koSZr79WTFfVM1DEcQDu9RVeB9l82e1AsBQGMQ3m8X2B1DmVzDATjV
ERnl/kQhcG7BWtsLUKgdjz8RCYPZju4B499j6b9UjUaDJ/L5CTXq74eDhw2pYdSv/Iu7Xe+t1gQ3
P7DGWUlUhdsZXby96rNTlvVpQmkbkzui2bopAQaxkxzIt2uwckp1du2+Zy/65b2t7Vdsym9BA5jN
dsSvKYBlV9CYjXoYrJkfpT3EhtBaw/P9gGkJquQD3nBk3jFVn4Y54WCJKFOtocTY+RVXqEMkiUN+
5HdOkcbhxRVtofHJm/sKbgvl9pvz2eu2ujhfGdIATbBfukVFT7WpY73T+OKH5+GVyEoICDt7q4aG
zqASAk6BRHFW8QBIoUdOPZee0zcFmBy7dyyXhKxSOigU3VrrWjjLm9seEboeByQtIorJ+xEKFrUg
voSmzVlftOJwIPR7EGMJhEXdfD6lxkQQaY2OkivtnR008olU4TYfw3bNCuP2zRNb5D3J3Tlge1Xt
TAy77wLV10g69LgI8+7cvTKlnXlE37jhx0aw99OYYryCi5ZZNSMBJRMg+XE9ulo4VzVo5Yfes1je
J7MX+QWEykDgPC3tPcCMfmTg7X1i3sw31filB4As8mThRjTFDhBxZsNmfx5JDAdbfBKDCwp80i5t
1+Jdwn5VpjE6+G+TbuDHvj2HPuym6fAxTk4tNjCGFSRy1XV1JrCEMolqQ7qF9RQwI/3b7NEg9JHf
K0bwL99w+DNOdmGBUOJJIBXwj2zsfcHd9FIKOdjdHEpkzv1KTQzAAhpqvkt3KOBol+VUlwnGb6lY
iUdKxW9zl0J12GHNmtLPml8QGNzpvtrWu0GgXVgpO0yQN4WK2f3oygYsXR0G3fep0/0hR9riLFZh
mpG4dk2zEKlYDE7cl4ZMnAxDLjQgTPR9gZhczIvByTP67X+q3mVn+h829VcWZkc0IFeGovvpbRw0
j/uL2eG8XGGP0nCKkTDKOsZSfz/EksBewc+YcwfoGSeElrLLSrSDQa7SIhjH4kySeHw1fzoSEpca
TAMQRotSqIoFVJadCZ7KhNyQR06DCskYxq4wTcCgM1cgK9zv+UJ7/Ib4wUjDwysQKzusewUtWdcV
N/WvdBSHEFszToDuhzWAv28B+Mr7hIQodnfMF4zKJN++PR6CSCNwyTm0//ScICCmlspsqJVGx3Ki
5l2ZrGwe2W5F7IboIWKHkdkZxNfF181UBZ0F1WP31GlCubUyCZ7xv0J+ei1QuJjGILXO12X/GRW+
50JSyLGzTgwDIBMNww/gw3iXNFT/A2a/Ua3jGBb5zy5lKJrCYXOPvj0hjNXZS/lzGLIbxriVj1O0
SiujgbGiezRMqDAnfYroBwGDlViD5rU1d6/P8An2x7UPP0elw1SAx1yflfm4ccSBBBsdPafd93fD
9DUIUZRmB5uBTOLKKokniUqpqXcsCSMDSe9GzrzEWFVPAZhllGFJg2d+F6Gr4pqY1ZnW0dMJh6Hs
knBfU8UTcasZY0EfTQXKGOxWaUT7RyLxnbeA5bCzsRG7R945kFTmCErJOhHujmOjrVDyyVGngbQ5
986L6bmcHvJPjCb05bV/Ny+d3iE14/6bc2BkmQq3v/9UClbEdU5CkVEEZzmWzxrT977JbzdVW+p8
4i52uGpm+/sTfD2CyJ8rFwyFagXrSi4WnxNXiPBSb2Rhzm2D9A4qoarFG06GZKYkGLkcr7muj/Dy
fyEn3XII0UT5U2J8vG35U9QE1xwBfWiyPfh+klWSP/DEs9uIIHqeOe6cg1IEHYnPZTFSbYfkvxJh
oT3jSB411XEmD93fZkLJ472waLyOLFvaKDwA+C6CyNmGwURNPbKYwJPp2u5QVSqcl/LgCWbq4u3r
N7Q++6bHB6FJNfG4VVE8kGTENPzYZRqW1lbv8sXD6t67Cc1hze2oIGNOYYyL/Q4NCemfcqXMsREE
KEfJuZtilTdErXatZ3k80PosD4K7+XpEEevsgJc9FEYQmltgfMJP4s3x8+OOjMhPWFUIMGOBynk2
Ynz043kFCa8frnBogbFr+g0jLrriMd2exZj2UbERQkWmQlcrM3HN24FCAA03V1tAGTAEMR/MusP7
vzIwSqagu6F/IXNv4dWvYBy897V9GVxIK/z1HkPh8bpZoEKoNgNQ1rbUlvmze9/xrrz3VxngepcU
T7O7HRAaGkyPQXyEgTyS43RV+5HI8mhAwfzMaGt3E+8AC5UKJDRWucZ5fSzniolProhBCkOMj18a
5+4AA+tgDZJsethlnXv1/vxb6IdmbJ/Rch5mGjR1m7K6oC2pxkpwmqXq7pB7fjGUeOimqyNmU9w0
pwcrgIYMMjEdgxGLQV9lwXhcnRUnoWNtKvBXFb2dc/3dw8BZ+6HUUmQqEOZzCLdnWVafYPeH48k8
tk9S2dHQ4mn/QAJ7Fyk8Jc+p/Nlvxlpd8Ffk+QNqQPFP3gIebau/c5B+sSsqtLE8I6w7BN/BVer/
nlcWZTS+5BV/6LgxaS/F716ahm7EbxXWTDzOdqZa1BwcXThLgBlP5X8MRhav2vlg64QBqSk7WQe/
zabRctSSYbkVjIQGQ8sK9treoiYYsF5Ourl8lEZOmf0Mpju8P74BUtioDqkhV7XmqKF7rkd1gAqA
IaCsJQcmr2HwQgWRafT4NBUQJVF/86xlhmAyRLxOTgoyqIE9AnaXWO0ZjHrnXIYMXhUM9VX7gMXV
Jxe3ur6CwZ4fWFlo8tpBiWrSNOoTUXq3x911OsNMmI2sNfVMDVXeJ/OPPgntSK/jUTaJnttmo9+7
CG6Oda1FaAbdGUOu142E0d9UAL8kV6BlStL6p+rId4uqecwha6H7/smSeWQ9k6f1prjr+1A+xtBn
ap77f9+xKzhG8aSAEGpLE7GaVHavbLDcvC36bUleb4PO4DEVcArSWRAdOv86A1FJ0/vp8v48JKaD
5yuI7au/uEn07IDA1tEUdZvlZKBZmCpehh4Xmxry5KmUZoQaMrQmSQoQ/9JEXPSho9qv/49X8uKK
DvLrDGK/6M1Rb/BuR3Nrg/ZIml+ZrZxAXnPSG6xbJJ5rpVPx7pd75E5o1VeacUU8kkAZ1xvxqUQl
dOvYofX8GVfLYZDgC4waL3TZuSzGoU+g5dZEI+EFdNs9EkoWff2uOwSPzKpGp2zJ95HSuUF3UIZz
gfJQD75cmV2bIosNArfOZerhbysz1kiwIyL6cm3ekVJvPmJIBIfq2vvVhSBUXoLo+LtHfz3H1ApK
arPOvptG4M9ul3JJSZoVALqenMcqvx/+DS778lZzCI/HB8oKNvj7Rre5uzqQh45AQS4iNJvF7ojT
vIr1JS2NJsY46bjFfKX4wnNNQMR2ggFdsRuTXTcKeDBFTYc4RSQp1igVKRqVWTD6osIQjcZPg7L8
rLK1G+PTk2Wju90GVzenpNneDtNEdrbIrIMmuUSz/++wboX7XNMdU+uigKgxeXBA7xjzLFumephH
U1Y6Lhg8enmduQLSUkNAE/g4s4X9mOPASvFe9XVdM/vACt+hgf9XZ/y/aTUq40m7nFe49rq3RyG2
x+igexYjkOmIWb8KzefVcy1/a1ZvueOG5eURWbOiTV0Ecsnci+uMu7zGCfGuIaA1mTMmGdiLTIk4
I/XYocfNSRSDiHdjKbHHaIOwRY2qbzY443uW9vT447Dcp6U3Gsslc4Lo5enhh6oDmM/tZp/rtcdR
ww2BQeFsZp3cEiAsg5RQu4Ad45NLdwiY3X52EmJc6plk6vEPR+auC93/0e2e5JUDtClHwC6o5zAM
F9Ua2u3/4Gj+8t+SlOUmhYM/wUv/vQ2eZXaUb2JFUAS4J5iCIQjWTXPkba/oNir/duIM+jzliq6K
ffAfRhMhZjJAOOJP1uSViX9h9RP9DzJsxSiKY+o/i0+4ORyJ3z6BpFmdRvxneQ/lcahe2rlgjjdY
eeBTXSY7VjVjAauHJ23O16eteNYd+A5J21iYLAM3D3x/wmNvD5c2LSYeGr/KgokH7Bn6SVXrIXx4
6+x/c4tcDE7wur/fDYz2RAt7xgfxi4EnctZaMImIX8V3Q7ZoqcRi0mu2hGeeL+xEucqsAM5vh49x
Sz5vrjkIadoggoNd01Yt4ygfF+aS32/P7R8bRf6UB7rSjtwJAVIatY7S/EfWhjhMxrbYUJnZidYG
GxRPGMdeS6bslCJXHDmPxZPxSPkEUjqh7+rMi3fVsOmuOLOMAu4x8H2QhDVAcUo3Foa2kmbSEX80
y1qid+nj5Iy+PGuaBHmvYjXC8+Z3vhikNzHcKxKcm90joExSNOdL7rmgw9eJniYbL60v5V+D/ykX
nzvKUOfTrz0ku1RfnHOYJ0/HZJJ9Yn0RzVkSV3O6d7zZmxb8id4tE2bnpOIRhRrw3nEVFrWsff9w
6n7X8Uz/qx6aRfGI2cQSNToApQeYmVFDzRtGl780oHnXkZfNHOeWj+EXgDO7yOPeJ/nDYUpLWzUl
47P7dBTUwDw1oCKn6rIK2K6AlyB/TNIVBptFbgiQ5sd6BmK39lTF2BnAWFZkY6nKkC+wCdsaTwvS
6DEYRPi80RD8wQv/R11eFqOLvXX79xQU54La4Ids0GLOh2GpmYg/yUPxDHe7EU+nPdURMiwyClMO
p8DL/rDpTATCrXPYxmzKyqwM7qaOxK5MHFd6rstWDJyvHHmjOMgjGDm8uP1uyyARF1g/qM1zp2Pv
PuCbrmeBHW0D2UOggBNVuQaeENOdd9WN6VaLqLcYdJZkK2TG2LDSg5ZrNa9oJZMh0hezEowiWz7W
xwnKMA5fpymok62yyftXHFTRS4LmIT1KTmk64cv4wNYyjj1vO+Xo+35cSFyt2viWJ4eLyPRPnMBb
AdcWN5NdlH2q2p85QEhj12je1Gn6/6jhns53kllUqUv/f3BGFoEJt9JidWkyIfTMnFYnTNXLFoPQ
nIIWihsuiJaAFox1g/OwsBKR917ihOMxSKHSUrGFv/D/x5M2tbjghgc/S0ODG1q6IJwuxCfBR9aE
uOGii1t9fi/8DlUTImyV4rKPo6o1/uhJs5s7iOM8CbGRw0Qh6duz9oS4TYRGodhvRYbvB9SG8LuA
fbKQTUnfX9T9JQk8DhCnZ1f+hHMrxf/wxiXAWuSOOsO8rLW2vcEWak49+y1aAI3J1hSU+bWBe25R
z3CT+9FVduAak2kKyXPcWGEQVzFsHGog9mvS5fmnndkDUCLV1PrmwD1cq6txheaqGHzbwf5DJA7c
xugcOxllQc5jF9OwgT/KVmdX+5nOjjpY2BgSUSSZlTSySGPXocHj/0e1/jOJbfmE191BxVLlYsk6
QevilBKjx0ntmQp0R3rH1Ic5m46gGlgG0ed4qM0EnM4zNwzpeBVSIhvK0/xdP+u0eXn3qvazyB4I
/FRFDoka04MuSvpzpaEQkQarnFSSVh/y32A3Icmfai2GKW/kb/Fn2oJFz7SqaxgP00lND3sjNzNy
MPRxVGTraN+mfX/dZqoc71+nEXRm4eSBXc4baEoS6ghOztAC5adm3h5IWtUwz6mfwyyS/j72QDGh
d3vdZePcDdDFjdVtLg6q3uLFYtzQfgh/2sKQ3dzoCpzq9d3TznVG2gC4WueXlfIcwAeUl2l82FVx
Bpm4cKrTQqqUbSRgHYwVsbinEMcEPWFVlgsnDrGtob06Q+SYHvHS2+utCURZJddthB0vHTCgKy0Z
D97EKpZvLiXqMnWzH+HZ8e2fBIvJ+LUEH0hC0AXHOXPSF17KBIs/ZFXcuUm4vtGcfhVi0tYXHbJE
PnVVW3SvKOcPCjaoep19Hkon+XxzLoeg0JgA8Yy/RMX2A+DCBKsG7OdiRJazLvpDYHFZdP6u6xhz
xGZ4wejBtpOkn3Ob564DKLAghqDhtZT0W48W4z46SO/ByqdGCpNl9Bb0t2rtC421ZL9V+0yBDwJt
fTcQs2t6sB/kfCzK3ayATsWkrWZQONYWZsB4QMQOJJWumF7/eb5If/ZZIWM3M9p/QLdlpEwXaMK8
pjU/dQdd0WuQv9To2BgYubElRciV71nYpET5K1NhyaB2pKSsBbB1zS1xUmRiM0MyrARpsrOmAbk9
2bIrnrS/u0fShDgyfGQxNtDTMvjpQJQPN4GIU9Ce5QM57Fd6XrC9xBRaPOaxLSBmIRDjhduKt+zA
wzb9sUSL0GPm3VZEX7ugvqfQ8/9vtJRrXLev61yJutmFKLGoQfzlWFFeu49TdVubxpS0LqmzeJJt
o0+fYqHgjoBGbxUY2+De4xL847LiQ1Lf7T5638M50it04s43C9k4lWMitOkueKj3RAfezSDgWZ0J
WySXOCBtkjFVSIdBfWaxWMOqmzmoxhPDzNDcdzm8HlKseXykjgHBYcNi5AMRpgb3g2ZFjJJD9S1e
nlDWW9zg8HyZm/LtOWTfyLH2EiC4MTfRIuT8h+Y1mCX3Awqzw+LozyeoKRSUC4hUFFUo5fP2xdHS
IXi3dGAOK8Eh2xas7t84C9buPQ0GerCQe6jgWsASnXhv5so8TkJWToj6USlUU6R02tRjfDjDe5pJ
xlLO4Qwn5tKxdiEgbuAgEM4zSp9TcL2f0dR1QdWkXpRL5lMgPaMElO2I0iv2z6g6humOPqjsV0lu
u7Tu9O6uKz0sdBtOBBNczZmCd9uaxdblEfdAM6cwAdrk4IoE/W3nU1PN+4FICbNeABpt6uuNt3uv
t4N7glSqlKH9Pv5kAi0mR8g5I+76rxBYhsUvXvkNeQ95e71TyfkhiefCbFm6DFJ12cLfQRXvlmb1
krj8q/03ksYdrYJxQ0DGB0lPE31twXXMtOM/ObBgdMYY8Y8yYTio4JPCCfi1yvtLAzgy0tfuVvsx
PEgWMrnQYzKMTEJWrmuyHDQVpS91wKroemcsItpIgRWxD/THUWkerr0fxc2ni1ZF7/wXKGhLRufQ
VfHkT+s78zDFHh8+zshQOah1Vq5U9n+/o1Z5iNrPYcUIlv+9zsydJUEzCaT5goC4ljWJyebeU0aA
7huWBy6TW0eTZdEFclYB5bjQdwDZPvm/Yp1blY1ZflZXk3fUg2dRD+a1iirl8BVvKKzzwOTkaEvT
nWuQGKKFWuc49GEq4Uv2LL4swhCbpETaJnBCC5ruq/lf5/OGnw6c4TrCrv2rBxNeJtVmm1vbKf9J
voD5BwJjf5X5N0pIcsdzV8G6gl8xKAzKCHRbkgKD/NRV1yLrT9enIxByoea97mnwW4qZti8jR9Ro
C+5PEF4imTbAIEXt3D7H5gzVN5u843EI7G4fu1hXo/pY0CF3pqQkyrUCPf4KZ/HcQZQoVC/DruJ7
4FhPOGeWaHeKWbLmJVO7WglA1E8oYzTqQpAs9yo2n4Nlpf2Sz2aAVcH8LLc08rvtKE/TpL57rq30
SQvbrdCxAJ9J7BHUXomifJa9vOgqUlBAWiCGNGTBjawKFoINoBCGybodf07wswlPTRmrE6YrM/hk
8k5YtaUupbGfjFs/cMtQorbriglXNEy+5NSUKrDDfc2PONeqLBWEt/LcfKydqVwu5OL9gB+Ubi18
bcv0l9vmX2EfkUz9iV+jc45w6bxIEj/3dPMOsq9+6caSYjWgLZkDuPUwJF5IJPnG6tooZGVf2jZ7
tt1SS/ry1yDWT+nus1NXXJjpKKp7tzDrRB8ySAF/GiYsijEX9gbhfMMi1Rj/oc28Qyo4UoFqdXPg
IEiuuj8NHJEbxBwLvJbq3GLsG/UiLP49GzEzH2CQpdW9Nsac/BLUdbeMMt4zhSaWxhFichSZ6ead
CtOnCtUb5of3cYzpYzLEffLAGK+kya9MKBCWUQk/FADZElQq4IzjZvtB1CyFCLY/2ClzHIMM1xsn
lSpQUeUfBA3wlQc1JTP5Yr81lzVnPgSWu/QQEd/WnLNhg99cwdFVXukWTCcQQHxxXWT5jalG9Ynr
exNpMv7V5TbOUb7iKsn6AWGDftKHUB4HnITeGxo+kuAIv2y3mFi2KAe/mh8Ppustq5JTVL75Ydz8
8wcCCtkqYCEjRm6URWE8WkTuqmb/phFD6nVb8z1gZ1DyE3qOmdhU59oW+ZOvxnWZMSj+IDQpNDmu
EAfpIIhY3ohvzyf+fvbSRYuxNehQ2QmEhUJz5WpsgIHdHcEa21tkJpbRvA+B0sB/kKD15jNpI250
Uf3f3m71TA96XvJEYcAOeq2QB94PX4mNB6DAgl1Oqt6NuEe3NtFfqGxo8uvsYVV33sOdumEqneRF
XcmZidE6rNzvpwHiZm9yQcgEuuUByZN4FDrLyx0X1xUUISkEKexXhJnGMhzST0QWsfsjditEGkKW
TwH3eVF/ryYFOw2jtZ/RrvpEP4TGyEOLLCqMwVrgtE62FH8L4jBSH/KrpZKKFejtCVpMyJQbNC3L
6zyhStl47CHv3UwGDzY81LJGFGR/Sw0Asjz2Km2GVOocnlrCNmkQwvKlj6AVVHDnHmEro2lhVg4t
6v3NcCBig0BZsxE97z1yDlRUCxm5biUa3Wu0PBOHFkUKRTyhWn7I+jD4zBEtMlw1OHJAnfycp1nD
O1e8CQ8Pl/VwT1udnZ8OtIDgZ8wT/38ofzphIWjFf1XBMT1BGD0FMvCb2wFE/ihfRyrQs8H+JTic
CEQysi3AXuv2SqFNG0FTKDJoa8fmihPvgx7dR0uEToZTroQBjCWjB2KG+D98fCoPoQmpmErkzP4w
niGFwzqLFs/TNfvcvW3SfQlc/e0UQw7UCrAA7iDXbKvu6uBfLMM8JJl0gmDg0WN+3jU3LYeUNFDf
q4GMfu/gk26r9rtwueX+jDKzyku3NX+7PG4knDgfQ28kDczPSILhPl9bwl/j+soFdpyXOteflU55
LWu2PhCrOPGvRWx7O/WaV2fAWO4DzpeBw0CVWmJX3uvwgpokUTY89L1WZslntVBghmSzdTXXh6gH
vt0WrdrVxKVPJqNECOdRFYSWwnS1zFEuH6Hnl0xlZp83P1keDYRMH1Q0b9+w4zpgWQYKlkTHl3NF
nyuwpeCDIAMN/vsJB1ubjZ99dZVKz5wY2IExi8oVICdcBZzcVmOQPta9IX4hLdVepHH8Gvh/4mfF
PwLfT2gBsk3rapvjrllFeAK8pzmIZ6QMPOav7h2wQg2HHBd5GVVeNIHWtImORLyxLOgJdnp/Cd/J
7QOgkZMrD7gNKJ3iGk3Kk/LqRJpX/1ky4Z43jyGhOSUXvTJNFguT8MUmkZdYPScb6/ggTDrnxzhJ
wNe5QmTnJR0xHCb86EzRAsTlARM09U4huQvU+aTI4XuIyR42QL0xYIk6lUVN5REFvE3gqV7eARVt
W/M/lNlM4RXOfh92stMWgJt9hfmc6vSMKuADIfQ8etNuZIbfMApjuWv2vj9+NkyoXPe4wsY1ulj1
7vlYJWcDVsJWpV5GtGgFtgL2r7JsOfo6Ek3lIoZjirwyszS4KC86FtMALSef5igJUNPBQQmx3G09
ww4Fy5jThGXnnKWQxBpv0eL8gFwlaUEDUlkMh1t0G7b1HOuxi8wp4/GQyZOCPEKmqC7VJsgUmmzi
0TS7X/g5b3UcVOymGdo5YcIAyJ3+r+NsfMqhWfiJab0qstAi8UaH6oud7vcqaN/rEY/VBZBrJzCx
O0fPXffDoTwsBBgoyGpEC0nzhzK0W/5/Wfcp1SBheRAIjjP5TQtLBUsCZnVAor9hoe2GBc45O+Fs
NA7VKfShkY69OdKphCJvixCMNQJROUOtIDj6ouMd1wE8XPYzfwkAzRIqrqdKkXExURuHXlag9xvf
1TnAgHbLYqLdxZTrAWRv+RRJ0hyPi0j2ftll4JceVXOjywIrGcs+gxy/9AfD03Ez9Av/TgRWPikm
VPDHPOAP13XVqqbhuw/sLCPw7WlXQ45YRk3Z95wDAl3JxglvWsibXQ+iJYIuuPeSvhnIO0fg6wKB
MA7HUCqFckpsMo6utg/Tys4SXtmXj7g/SKllknGyMfkzHXjBG5NH5k3L27dU+8utLepm87WYYsJa
LZfngNW5+pV4ltcZCr8jC4u1qSo2CtX0aMU0Rj6A7NZPL8Bp8YS2yhgSKNngmneERVl2VFPavyEp
r+N4HRhP4Sndx2L8tshaJkQtZsW7eRXemQ1tBU0kTl1QaUvZp7sF+Pqe6qUNlI4IdSQB7/1tcd6r
Fw1dBFOO+SdTxFpR6ipJ219uTtX8GI21qnaBc/ZsFXhAGxz6AvPseXocjk5+twA1ybum8ojQyvwE
G6wu0jeMRQweQDOKfRbwfuGPsFTSpNCs348HemgEIQjbO7izs4IbFvVNZpckHMwhFaDU0qoyzBtw
xZnXya/G38SGQ5qCOjG8qHXrvqATVg1nk6OpgsMZl5FpxFDVACTMJ89XEOTteG7KexLSF6lau+Ev
gExgLvwYYqgKCvgmf5Ha4nwy4wQnn92IKLG9EvhKFu+mUlfTHz01eNnnzfJLcp/MdJMMQ8C6NWmf
b+xw7GmnAb66+DjBAyHTiKQl/t8+ojoUgUtuiWfuzfcWMu0fGbj7fW9d/RfaNnbM+QW2t7kuuXyu
llCSxGu+IGoZtK0C7BziOLVVmuP4LfDEaApq86sQHivCVLVw8g4pU8G0rs9KT0b21Fb/70aEe98Q
/JMT2egV5t5pMmLjNhVJ2a+JeZiXm6m++BLxpkVgZKvaXH8CvmsLwlEqutAO8Bqz/p6ZHkdylv4A
KeHZaCe02NZzHscNa43c3QGgkO6Udt6dcon2Ib85fgrex5Xn7IWQHlcUay51G/F2QA7W9Ywx3cl6
eiajtEjeu/ZjahQfjC+JMmJmibX3J8XMO3BKSiczfyPxJ7M+YAfzPcf2IYLT1zkbUgD3zvs9e0mk
qcxIN8qchi45UXKxxuO7Z7ksP5rzCjsx5uxqR9tvZPyumX1VF/xkkRgYo7V4VFjaU+r3HZEnLWgD
JF7QH2QTgepkCtye3oKwEufnbTXZOA6a8QtlABkC9Z1mssQzJm9KvuqRDanjzm1Ftt4Adk9gpaoH
v9OceZao1VzNH+gccr7LwN/cI+B1D7Ly0knSW6Lx45mPBqLqBrx5PIdDvjTKj05dTfZYjfrjL248
S8D9rUbuYlsqaKbydYm//WolIPm2+kRQIcZO+R1dy7DUXKo1K+nzrQu7CcVQIBSi5XELrIzSXeik
w//MvO5+ORoHturoGH9PzRMuuJY3bZKbMTsCGIW3HM7CnTgfkYx/qSyyKYBDrzjPRjz+835j9eiI
Pf0unZED09TYs8AgBg+Zc98ac2yHmllXhy18hSoq3yxfyYAcKDoqfA+CwhVwY0Vy3Aa+v7HDlqja
ApK9kqEq/j2i3Fh7sF76K1/c9mUmltvExmpFAoYer+jP3pPAkjg90Fjd8cxvw+bJ4uTdgjANh1yx
Y2+ptXYA7opN5kHZIZOgldiHVJMs8gTMy4BWARgIlNrofsE8Kfn60BerjR8t/cWGWIpv6dBaNRuF
u9SfwqYU/l1xCnYAemc5boA2iuruZmDmMogU1IkIYWFGTNYggqBAYK3UQKyXNza7st2DyvpIcqRv
y+i1aA9RFjciRVnj4wbdaijsfL8KaT30ydV/9JXymh699S/GED7pvMpFK08V6dV/TdiZQYcpyyn2
pfU+61NguDa+opaXGvFmO1XzP1+1fxv6Gajj7rf+L+N0xiArqO5N6GRHl0x17T8azKGsOsRZaqWx
MkXJxRg8xkRcYjkwQIhqWNzNppn5JVWe8+bDR065oeRfQmVmQzWIMvwRoYrA7C1J42tyuZ4MsuHb
GuvkCDeZ6BxFwbwx3FlwpWLblH4wwN0UuO4SRbYzoHI33Ra/ZeUJ8WW+V7z+GTiYJHatRu1o6wdS
nDjAUbuaaixGfG7F02//Hxkq3nzrEZbAdc5kbTyEzdmLthgX4GaBaUMjjDiSiyrqbH5Aku+GhxQk
3ahvVMdyqXLIwhtLG6G+WXOMzz/2U45lKzWgo++5H3zkxAXBEX860SH4B6nFzCEdILi5r2frCqCX
1FBAuVf8/YX7wu26xXm3yJ+mMHHY7JlcwRKVR2yKeE2v2wiFZ9jxzLoa2kuTalLTNUufTrShWxxC
2XyLhiJtkGO66OPxWp4i5rZjHj7Gq4x3ZKLlW6XKAv2+qyL4iBMNpAYn1MXt3m2mw5rax43Gvne0
0CXhd+0LWgk1trZv/pqqjqwJXhvFEKyqYDxwTNGkC6c262Msg6HWy3nF1cUZIj8yluPwbhPknCX0
QkDr6gmuMSKOMRKb6VZKmr6NpWtrybefdbauCHTwSiNT2O0sdEKpvkIkKIDGd/Y0gG3fJKoW3oPu
g4TJZ96459ExNB9T6TPJZ+7aHHQf6z1kwnPDFV/lK0nen8Fnbu942RaoxkfftcF6+MGQ5wjgtl7E
KsP86vKKFUAPQ0I0R12Aelj02PSehCfzljzm07aHyPO0hc+bZKExVN5ul9hAzaJLSRJixkQ7vJea
tfXsdzjsBEREvEPaws74AePArsoK5uaA5C+ApWxXl9E4fKP8mYNbZsRYDLSzsp/uOlQR6Pulnmwx
5qoHLH2C+NezxJq1ThaU3Swvk7Wt9Ltfi8gvKqWqAXKZhU0hfZQs35vn+C7Hqy7TH3vuNumVsUE/
yFaHKY5Y6CYuodD157c2L0OX744g1QVT1NiwV0TRGS/Yq84EQZR6mLbWJhyY1SERuBIH6/BHUZAU
DQVjgxrFtOFb+64cdKNP26tAfEl1OKUp46SHQkdSp+TCSsKYYiqpp8UPIQpNk/7igX0S0+VWs2Im
cmgaosNfhwXDdbL5dluRrNKacgi/wjPDpNhS/wvYYTp8VUmok2DjnmkekMXjLrTAtoTa/Y7z4S5f
wvnnS5vXnZ1mkF0HWNnmMOmtDYb02wOE1Kfwb+SjA/ny0J6OAbdfwJJRlAR7F/D4stodWLOgydex
qwxRAMGF0Y4baTvzulKpKY+AJ47eIYJ+cdhcHitk4NtjF4LbHpqJgeQJ+QOYPYCo61SLTAXeZNzt
k1xzFYFPiSeV2TlsOuAUtCezxwBeGuogLvkc14A/fP6sVfqHRSnN5vlFjZPvxFJlfIxVwU4BN9BZ
wkGwAfMKEiwRNdsI9FPOb73xKqhmx/+MnxKAI71/gnXySH1iR1IOrambFqKgglj8zOx9sqLNuqGQ
ftZulDnJy2J7iQphpQhloqNCo1oS62emZPpnlZUxhxYlesxbjtsXXz70bwGoALJRO781AvHCJB2D
/8TDKz+RTm1SNguXZB+E3buH7gkSSsyOrKF2H2cqCbkZ40LwXjCK4GAJq4D1kF+pP0uTTcrfxlA9
90oovI6jrmjupYTatcQBOd3dYnaslRQHb7w5bI0asH1G0Twg+yIQW2hEMzdl3XzqdK1steIbwZVz
69Uoi6jQAzKivFCADFHU2JnPNidM516W/Zn7Sq+XWtlUDwQsJWG22A2RIA9TF9XO5ZhHGpd7RdzS
HP1XomzxMZY0VO8wsTRM+ft2yYN/XJUIEWzvy03y4roGOksv/LDvvG1CUVsf3b12OBxS61W8KBM7
t2e4duWl+f8uycbLJcmFfFFduX1LuJhYc13lWg4lrb47ID5nl06jz5Bvh93CK2izTwE3rVQ+0VA1
eWDzt61A8rBqykax3tVfB+NU8o/6TJh4P0igJ8OF1ZYGMfg4uZU/hpuqzEW8YkZY5JIt0bFPXosq
CXwk2H55YORLf2iKiHXj2su4qdyytlLhNo/FlzzH6qGgvvmrJTxRbeoseeVXE2YTU70kLieqg6sk
e0GMPHW1U/GKN9Z15Fu6HnlcqB7lYdhaLrjZOSccsj05vzwsW4vjtUhY6EcVC6lpnPr6Zidcqo/v
qeE7cXb+lVbDzq4lryAeAq46VpZYKRjey6tYik1CycmJmSGQVIqLZvhDpauLnNmj9kt5uCoJQX5B
lO6jIeNxaeaoZef7VRunJM9hB3ifubpQfOb8NqKFS0RVeo5nbkmrN1+qvZlgBOeE1MyqSE1IREUf
zkZ8LYjGzliqZH50rLmxEwBG50eOym2+yg5eR+TTj7Tj8VvOhR0OBsHtXq8mCeX7GSEzrgTqtr2R
xXD3e0D8HOXKDmywWuk4Dc6czA7suG7pgCMPh6gHIglNozXM4gfsauieL8ulaH8kCi7qNjqPIZVp
KEieFC+Xbvnc7MUFyjwHX6UfW/EFipAOkFrUCD7qEE9yiQ5hzYvXhuOuKowVeNIS7PtBTDgfuKDw
5y3YldPLCCJoV3IPU8YH1x2s8R+i9SfI8Py/lmpAPwSx45I7XmzbNom40hZAoVD4iKXvR118mA3B
jo/7dGToyRfzv21pGU1vjwbUQxOV13XMr2uE8ihq0NH190hLUn/vPYCFk0mIDa4fLW9RSECmnOeD
YjIkzpHG3Ln98V3t3nx5CxttNbMQQJxt4977b9JxWpqY1t6x5me1sLPJ49cjdBdcOGpasMAoJZae
60GZIuWo0rjr+ucvw36ec8GhhPfFy970jIWmxneBkhkSFzLLEajDbfmgIPPw2n+SYK9zaDgCusGL
b+vIJzK+4dJuepuo86HOS1kTgHHnanFUlLoyWaJdxXTc7FjF+BT1mN6qtJNzC0xH0c9MIef4HOCB
5r4nfDlZ6amiaee35IeQxCsU+U4Qjhmw7AQWp2HEMdumL8p/YbC7jRtIdPhkFWatTjq0mnkWgMpk
2yJbW3iFnDPYXb3zQkXWNO+H+2/XQjv5qYFUeuIJuZ5cHMntA6M/Ez6+/d06kD3qbYozs8VxOhtl
YURnqxBhALRJ2EGGQyoW6L/2PscpvfSuyTIZG7xBHSnK4TpkLMcyXommZD/icp6aefAHPCtVAsSk
6AE5BmtTELtyBzXwM6qvKX6A9+VFi+gDqLTrc8+orZEP4z08qHVy7RReMz74HT9sXt4YwfMAum4B
AZZ9+wTn1N5IzFaMN7Hf+imbKGLWSrB1jj6WzNFf+SwerQCfwHpk50iLnmc5QcdgyQGvd0XshFb+
wv2+chJEftV5CqgtHyVsewh8+GdRr8MXXffRy8+ocCN8irJtYqWz7VMzm6Gt27F7JDRo3Mgjvtxa
fSZBkQrwp+I+FTw8X6WvxxuHgMf9fBrtX6GPMjiMbBuCUhPe7i5qFC6E5PAptN38oz41EOfUdOPW
FpMTC0R4ex8q6Pydg3681KaulHd9KKs1gomVnq0tmI9Zog6zA6kH6U4zUFA7LIVqsTL2qDRWCVnZ
fcsZ1/wf0uEcpxSOMUw3fEM7KyBMXw5h9C0nV3/+dA538qQ6kdiQ/s6SvmcXGAX90Hk93fxhLr++
8V5fD6CcWJgNdraZNDAL7omCKptrkYUnkq0Oma40q/65ssh3LpZadhoXDH4IbWNGZShjp8ETd6PI
6hJb6N33hmyVQgNnfLNkZGryVWcSK/QkQkvLvpe2QhS8cRhFwQM+f21OMDfMiIW7RCHoRDUFL+mD
bbaiEjGArQVc3kR3FaK58qS0nPLlRjLfR2WXi6RKsp1A04w0XqDbloahBUTxneVNz55pih11cc8Z
PkWeo+G5yltyKQCmEsYTUdwcqp6aXFbG/tpN8F2ybyKr2bomOZwtVfho5DYRNyN1sQ2N9dy1RQQC
2V5Umqf7Zn3Vn2bD/JBMwj4/5ulIFmoiUxJ6wf1q2H/7x42unwDwDxhOglSSWIzXLoJJR18Gw7Hs
iahOohjISdxCEjFMjSVOH4QoXsS3xkFhkFbXgeT7QZL2B/vIcw+HtCwLLtQTWPsEM+CLKix0IuXo
oJ9wKMTHOoXUF8DO6R+rcQOqBpXzITLCjPPjeyJUunltNmJ2qk3+S75uqIQikwDdNwJd74uBAwHB
MeTUBe+rXjZIfpLW7E0miXdi5EDMVfeHZedYMT21j7cFZsGnmufX9b5VGsQyS3pwSdpsTi3yQzjj
Tq8xhAgcxauvf+Zmu5trTSUDrhUL4Bt3geXg0PG1ulDQ+8+3unOiypjd+Pbu8aLaLNlNvqIz119y
VIT65LJghOsIWDw4tXwDII71DKH2UanweWQzL0Td/bgP+la3SDX9fOYzcCpULme4tbtlKw9Hn1Tw
hEOMrUFO9pAAAi+YIDftHBn36z6KLBSOe3KU8GMiN4W6yR/h0b1mhegvTH+1mvdwIMNbAE2GBS8/
DJbMI0TULlFzbZpjeaMeJQM2AsMJKkMtp7Jxso+DQux4sfOSk5XHGw6+yoy/xse2cOgV7gvm564g
G/i8r69vfi+BPt8V7cSnAsfk1lwJFMlYNhAf/CLdaa5gi/0+8y4AsXVTc5QSJpoaBcSC8sHEoHSh
ixB1E90bomO0XXop1BYqfe2IyheNGe+tOwferWfydeC7TFBzrgpOife7jxDAWHMT1DmP8T6x6kSi
mW1UbkzIRp03/vrpyUhSTd9Ad/cTPIw8LiZH8ojPV9np972kg4tRfoKy0NYzHb8h3Qgn4AcSrEJP
W45KhNGTh65W4XSA/qiT145hkGBK9K6vdFXmbxXWIBUzVCcgIrdkc13nCWBmFFUvnvAEFn/NXo1y
V2f8SPf+ivmNLfQGpQjRlPRreOS8TVSPjcAsI+sToPZiHF/ZlneInF5+WPKnKX6nC0xwWwCtjSpx
Hj09orZteZvsMsHco0yQvEKmmd6gGAgo1dF9TSgT9N/ijkSsGf8wccoXJMmnGDoowwqxFgCMHD+y
WTTWelV+pAauoPN4fIFuBpeXrLD+IwAYwWqFocp0y2cY+KrmliGRB+NERZxlPbe2LhAmkiekteHf
Y80S8OczOj8FsnezeYsT7CDmuensj9e+AVtBcbbTvs9D9ArNoRs1diDuHJRHD7fcXZ2/eFBazLZl
7sv3zcjmuRp6MpXm0VKs6QbEcHMbqVQmRGcDgb1DdpPGb9ft4nubrlKAd8hnTZZxVNHOUp6PP88a
xNBd30OnJ0sO1aUMjglR1X5KfpnF7ClySIqfWl+asguW/gQZINdxureNQb7wnxq8j89zmzhKFaJO
aEXrwnR4ktHX0b2md64x+5p/yXzDYmge4wR8Dj6GEjGVI3iFUJL/yH8i5PLqwnJovjZlG0T5fT9+
F4tI6aRuv6q7vU2yRl6YlEh2HgJoFuo1Bt6tB7+/qz9PMoi/j7SCATwWgIpnkKhYkQUtKrrKhzZT
WpKSt9GDtZAZ/A6IjOeK+xbiWtp/n4mYm/4JJuyAaBir1KNiV0G9xRgz2RgyXtbebFBeMU0IjTjk
v5N7THJulvnopJgq5h6GnS/HB3YywDI5GdktBUQeRDFNbnNlwyC8DQYdGLEbAepMHw77+0uCtpL7
LNBuFqNfTATSr1oxIi5laUyXr0umhEOxU5ZjG7LTUo+DlvLLKI66nUX0kFe9soWoXyzPiGwTfHXu
xnlhj8jROoBbFyrlHBQ4CEc1BcfqdpfBjRoHNZ4ZBGlK5iJvBZes9F/Pf4uB+93KHsir69UijB1P
sdBRKcAjeYZ7jVe7gyx8xHjxerYd/EXdDaWYqdm/FJa9hrhlTYVfZY9vV5LrFVlAkfT4S9nAQSna
YKR4kXPqzxfBX9yB0wYmBTDBpNSd8VbFl6L9JoseuE5MLoQJSJDJGudv8cB7zcTG6LK6uZ9Pzci5
YOQpbqBSNS8O5SdeT286cm5Wp2ajiqLKZe/N7FDHoj6CmEfUJ1IX2eogbmmvUsjfRJZ0qpFXBPf1
J7Kbd3NkD/dtp2lj1SCXKLTjDnsx02g1V82/lhNLV1o/4+zjUsGBZbgTwagufTPTz+4PwvsGBLEN
/v2OUIFLZnENai9RrLxc5BkrgIslrzm0I9Ahua40RI1HUytk1b8B/9z9VMjfSrGFYp7u0BldfdHm
f/7x3PAZOzdVDo5vsm2sGyjU11L3GS6s+qYxrDcgGSDb29q7IS03K06f+Wv0yzJR0tjPCdLrBDdy
qKv0IhopWodRQeBc8S2q/9Gh5pYxoNajcE1OZFKV5JYQC5HyHRlnMAqnVijCwNUM0hCA4bwREoz8
pDQIyRjQhIYL/7754qtdk2WWLoAsg8JIADqyPDj5sZxly17wJJv6si3n4EkBOdYo/6OxkWvUV7fg
Bk2vILkq2J3FIq2Wv88r0b76sJYQESquW9qZfjc3/US+hBs0xBsnD7+xso6O2XF0sUI75cKA7Raw
C8K3nJYT8NJfanvY+L+wNU2X4TjRqXRtHyshdK9wtZxPmie5xPnblOerqEqwIYXDQfAZEpXfOjs8
nDh5sAAYZIqUWhtdHCD4NO61EYg5JsF8TQ6Ne1RBf7Yqv5WtzPdcOFdhxOgJI/w2ottFg/qS5shQ
1xic74JIUu5yNqL9mcp4HvDv9d2oXeq7LFloshFOehUFji/LI2fein90oOcSJ3/1/hkoyeG5K5+/
v4fv1AIB4wXGVpLBZsJAI2hTXqnTsE2iM4Fgat29zB5YVV5VpNcKwVNnwCcS0h/XevgNaiz52hqI
P2x+hpR8s7t4KNKS2F02fJCG6oWoLRH85o1KKG53GUbYyzHIpTi9zDkg46dRX39DP5oYOtQv4Ccy
7xltkf484a0HP1ncVoWnGZ50PSTH35d9/v8V/e0v6fhTmZilK6HPxBvTu02vwHVHhBf1AM+7jcdc
NgiFECpqcvIiUDzTGAdPHPLObW5eEq4BzCXqpLZ3zlbo6rlid/I/RggEZrEv5aWdZIOZv/Jcge8b
WaS5Sm9j9RVQll9G242jTuiNnpCwKwAZQrotbm8N9Rmun8SaZ8jyBwwkqtDwxdB8dcMChC2CJmGG
F27aGNn4SjCFM+AYoS2Q3LRrL5LF89CeuGDJlC+TkygUWabcwClUuI8dv8iTL7L8OhX8tennPWTJ
PNFpN34N4Wex277qTW6AUHI22G3FE5ZcHP3jSvz0bygyv7maz07QbGRovC9BdzFcRMNN1vwYsC7R
XxgqHdit/DB4r0phd8KsvjChzA4JynW038cN6oz7VFU6HDhJlDnG8nlBOSdCewkZyn4W624Bnh6k
qxgU5slU3V8/vRhlNlyjqKwlXJJCGlmxMXdT4iYri5ye/Vz26aPMw3ymgDAgFn5L1pdGHvdmTIEs
CDIxr8c888qGLw+py5xF7sr7uMKe7dxqJYz5mJ76D2QzxRmn1u8FWBmF9mS8E5c+eOSUgMaxA3kC
wtmOuWyVN+yem+xOHqIULkh35r4e1+N+efDABPkGLPgarEcRVbsyd7OZKfO47c778A0v4vsM88pg
0q8zVwkCV1RU/xntid8WMbZUEDh2Xx4L/Pb7Oe8vFAQEW9ehANulMFQ8rzsw91qdluo2OyFj4kWB
EGBgBnC5tssuSD9TNcsrK13kcr5ueCmLCOXeL/ScmtMS2njsnPreu/qDTFFllhYCE8qE4LpNA+eu
O3ayIOtp/69hAyopuXtqCXafEOZGSPEjEzSLuna1IBpQeN88j+LrAuQ7bgu4JuTtctUMdNI3qjsV
GHLRdWyvkKtpm/F5mhkdNrSBc7BkkiZEHN5tVUhNZuoByU6l7y4hWJLhBy4Sf2oJTQNdr9lY1qsn
HEUvPSR4nj7wGp2jkWxOvoZTwR9BKqf3b5oSqDbVcF/ip03eMp/f7bUlb7Xdchdn+06k3gm1pD8/
VwMsr4YI52NMkSmjC3J7a58ZMcQXAHJcqHeEacXP4+eOcgATJY3z7BewBdIH2thelLTPeGHGgKUI
taJWXbRHpyz2sJJvwXgEp1gHzx9CgGA2A7NIJVnjSYaHNeNOX2XdtDQtFXZLN0VTZpqkH0Okg5nf
/hywrcq9wJ+trCQ/+fN5e1rZrhimzAKyioSyhthpAfDDZJJrPA/v383YlFNiIU7QF7mcQGKw/JW+
k7xU/Lb322TNLL0enYNDljvn3+q5oP2NAFcnyeqT60qqvHsOOTYaLU0aHhg1s4IfTOJXxZInBiss
hwZpCTzQY3/7crtnjB1OgmE78sczlPFfr0WifQZfgyUORxPitvQFv7yuFOBbQEfC8eZnN8LpZEse
DJf3J62A2CZWmb8SBGf5S6B6Dktw0ZdjZMAJ1dEEqaYCZn76JYySUt/LYjWukxx8i0hyUINPkT0E
HUnqhypBNZ/8m/O1czIDasH6dlGlk7w+rlYwU9adjr8xPawCyVUhbVkN4yrMAI5aedAnB9DIoCc5
AlW8w67pFrgiGKpbaPtRlmG38yUy4WJAWHTLm2v43BMmjVDfezbaOfJLlhazCyzLASKR6TeH2O5W
phVXb+0K2Et/C3iB2qNLBdMA0do1QJOez22ZxUwny9WFrZo0J8NqwG9KXEFNHZGaLaG00iJt1AVi
ub9CUyGS4WVKFD/Tjd5jp67ZPEDhlflxkLieGHb/370jYo4bfVO3L7RWR0+BDFWkSr6lfphkRpO3
1S+6sohTa6i1dlYhUShUAzCM8U2GWHVtXA3P+YcvJSHAiFbj0NmkbVCUceEMa+hfV6fjB0M4aNPj
IkDe2Kb/EzU7CFqzqFJcVo9KlCbwyXLwzbHJhsWwtlDqKRMqKrGleX0PW2EZnuwqCsCOTAo7bUGB
59yrvz4OYAMSGBrImvVGuOFcH4PMA7qSZwkuqdqba45MMmoXx5Mq1ai/HPWExQGzyqSI0r+VoqXo
zH19sn5GWSlojwFMweWWeNkyUBPd61av1EChff5gvc+Vz5Is0abVfok4d0SaiXYKBVkeh8ShITnd
cJZpZEUfaGQ4gq5BmN8UpcqWQnYgVfGkY01JXJ6bleF9l+URMmcDzcAr3jEywG/VgUmJRQ4Hj2tT
RgupO/B7zG6KcR/LGhCniyOY1uljQRi8oruXZWG66UWsK0NYu0Gm+UbOoMD2wNPkZKk361F8u/NB
GEgxaMou8naophz6qq6xU6qXwF/b+XbjYNJvynlE9OtSSoNykBIk1YUpLKS502RNoc2wYJ8ybgtJ
0xaRZE9p8AaCpSjAQDccXvrhYaGSOgCoIvQ4RhPo6Ocn2mm1pDl4b/i4wWHJ86a83XnyD87x+MWM
UUrYExPFVWYSXstpR1VnVfwdru7fcXuioyzh2KF7VgoApKVs9KUBb+wr5qGK8fycTqd4pPxTuv7X
M1/B3RWXjpyJMX5gyazsWiW1i/bgLTJsnxu9bxeXjEH5D9X4MF8eYISGzrlVaZlVyKhwDom+D3+X
eOssMgCIczHRFswYrZbWulzBkciET3mMge0B8g27bmAilnM/3huehMwRSvBq0k2FEXkBJ04jBq27
LM3RMrpezbk2KW7HXhiLtMuzHxSIkJxR3qSQb7zhat8alKUzyJs0cADxxTa14ukno6NkQY0aotIv
bN+txlODp9mUjP4/o91I2KobIqJhjSO+Xnm39FO/Q9Hy5+H2dHlWfXGu/2q+mCwyLy94hBWEnnIj
eQdzfMOQnMQRLNeK80dSigedP/r4yodlajgxoujqwgjtnhMyQwK1F7npQzOyBHmU8oTQbPqqjpl6
udUE5rpyeqJe6idrTPajIcTWO8c6QflIKcpu16VXu0JlP0uzaU/wWuyNlVshNYa3pgdd6SHDJPsM
nZBBIbVRDj3ITPw0vBjjIxgoqTHhUhMzVomW0K0DRufBCCbvVBhi/NGIgcOAx0bkL86n50itN/Of
J0BCMWoZ38SXyYAFMN8VHWEBgaFufCD7QuRej37LLLfx6HPguPh9U++TkS3EK2Thcblx4/ZHbdiN
Ej5ZCM9hiWBdsSzkp9n3v+b5HpzcPA9ar1iCu1LMtH7UC/0MjWgPou05lThiszseEAQS6rGIqTG/
vak2qXuvr2b3Ujss0nQXt7RGXCgw9jjSC4M9R9d/qyBb9UVPxYarIcymkA0tYSyvtcEXEKKUj8dV
koZjZStDeIjfJ6MR1v8FSE5lU0Jr1pPiVfgDpSBHsPJ541XYAF0sSvqzLHtJIPEUc0L36e7zBdFD
0Qv3MlDmIsHcy2yoa3wjX96JYW9BnVWRMwsyu4s+lohFhtN06zsFy1pLLYoAO10Q9V7ltRSIhNTY
FDN2use17Nq4tpV+02fX7ssm1hokGmVF2VUh1Ie8VqUFnUbvEfh1beAO8FbASYdLwnDlDCjeP8zt
udIVXx+IzCc2E7wNG+r6mAi/vtfZp95mFIYvVmdhEhyTPwZ1UsYfuHvFK0OGylMSFY79HLuGiVoy
QBZUW/tuTsjOm9VUkSSPh8X5QLC4/S5Cl6pW+P1US1u3Tpdf5o0bYvDa8rQmcpQzsDJdgl7yPoBN
2xbv6LQUh2AGJ+qpQahv+0RDb0UQi2fz9TQVOA/8WQcFiEMp22NkGUQ2M0Nnx7eHpTpzkyFeyEkM
8RTUEJQQBLBkiyFIXiakx2RK1xvMxV+AAQgyoeNrri97isGR7Eg8+SY4InpnPw6EYnXK0Xu9KNfq
cUifu30EC6vFWfKobolh+Sc6S+IUwPxSZxhzIxTZw5NYFkUHHFI+vJz72eRvrCsY9yqeUfXjBkYg
qWbetDHw9JiGLKN0/QQVtqyCMCbVcUpJsDKaCxWqUz1+dgGiz92q0WkBuQZelANJF2C8jhAxZeab
s1SrUTIER3GRDWd9hLxzy7wTS3V7g/CZ+Pdw0DQeecCYvHC/AR7ecLW4tI4nnBzAnxFkfjAkQ8KI
s81nwV3FQH9vJazVgmqA56t+FsrrR+kia5Tqo1SAZstaoM04mgPPfq5oA0jYU3rSRjPTooktsHcD
htunwCIDMU5m8cAvA7omd5AoWbjrS53mxLqzSDVOoFKl4X/l+Co72WcRDz4lKD+QBOO6Z0dILVP+
qQb/JLUknLMXdz0HzXrfWyoZGBd8lMX7hoiOJv+AaJlxSUgbiyFtvy9uLURzsO+leuSsdNGQf0Q3
XkusGNKzyH1EZkXGg1J+MpXKPcww1s1oj7FcXA6tKUgbRFiVxWpXiQHGKi7cP8lJ+AoFql0rg4B4
8xbAsHxrwGGgkw2GHJy+Go2lTllz6XtloIqfKKQSGqcmlD49VmW8LD3WOztsRm8ZhbTCy/oU2Tgm
+C/uM7RxHGjGCSrl6/jFiRd5+BQRI6TvyVv2wDYzZo2bqVwlaDENBAWjmP+Wh17yEKCRmVbMom/N
tXazy/Sl9BkHhvdGAVqglNAO5i/bCJ463rmFsvBaD1g7v3eVv9HlD/93tIwvxdYOKAd2T9NSor3s
PHlEK4FnedOthHKhKdH0ugBIEAQ/ZC1fEAcM7Qa04AeWYj1jkAlQEsu1tmTwOGN9b+S/crx95A+j
s6HD/3DeZll+tF28J7v73KyyECE5QrD2BAhr85C8BPttgboxhAfa9RyLn7vGAgDmXi19VzZ9nGkp
Ag93ptcbnHt66197layE6tIJWgRcMdf6T26PARVMMXAOQDLEI8gpSxoyF6tvQFPlAEchWrAVkv5B
5nLSLGjSDm6pZdN7XckWu4rKa3ny6wsDmneIJ9bQdRiI4MoT6AUSHNe5PU637q5IochyB0drU/pa
IVlH4W//7cHDEA8iqeNKbC1uWfQqyZaM3s5HR4mh+QpBEA1P/9wbhWJJ9RlondlIIM3NJ+am0uAy
U7yOrLwhlrOLHvGW0EH3CAdy4UOrMhckDlDdahiJP1vpqzPydi4n6MtZUcbhjIK8c9F49vfHoy5i
cAUXIpOYau3DEzE0I53WLZ44pmX5MNKGDid/sPaCb2w93dsTcnuT0PdqPzryqZjuA43+3V+rxLpQ
Jz6Ihk5E3SHlovcLeixgauV+4ihX8kzfDm19dyA5YY+W+REIrVW1N3Ivq4aGwjnJNcGkyAIeO23g
YMG8LC7RiW7HYTvVcbnClDXNkVqrhuCF71Q1tlKG++h2QIPgIh59GlQPhNo7Av+AVPIU2kq3oODI
JG6PGOe75Sqr7GJ0S89+coTBAvB/BGmeZHDIcQCpNqDV6W3xazVZzMZEi4qeoMN1nA4clz3t1qU9
VKggXgndtOBm9IQsGRkttretqWdfrbkn+HiXh7lTx7yDUGGF3msaISYS5wfQUBqab2G1XnMLkpoN
aOS4xUgjgif/57e0kAqEWbB1fC8Aa/QGyyoJwJN18m6X5mlCmV2v84ZaO2ug1irxPPWirhbSMzjJ
gjOBt9PZWTY7zyurEWpkaLdaP5yU5GaOICxQ3cPLxsTP2WP2gzzQjj1CLcCJHeWcsgt753gEEJZS
XJXP00GsLO+E4xcg0Kn2AwCwP0/Phtq6EczRJ8fLIAhaxf3lWiMrLsNk4GeUMWo9ZlJeHnPpp6y+
KJ4eam2kPGIcak+CQz7QeyjbR6I7dgWrvQ+km9jSkHl7y2swyqzgW7L8itTR/KtLLg96co+t5AwW
V0J/jy8peLya9vYmHkGoSeWXtQlOmjdzg59zYMqGECH+1OOz9zfO396lwR8C/08O1yAX1Rk/tiLC
yENuInpGAXlle7IYT7Q/3TgOrDy+reo+DW8JXLzS1Y1srAUNIfOpEO09CJwf33LMzEtPaXVzcDLL
BTIPYh3IBligv2lNlMsXdS+HkwolyFt4Nz4D6i0je/wev7B+sLyM2OfbciUBglXxBvNKv2ePodDH
6Rrh9lsKu59UGE4KklEJeKDeHymscOxCBWLT5cqFixuqzrwNnqC57JI8628KTYjTI76ucSpSMY8S
ClGRmzfig9UjDvgFN+6/gkDdliu+KycxZ9x8Xa7d+6yjxgG+jKxiv23sdnJpLKNHe1/hfShLp5au
oKOvy5IR2OKiZrrMOgCyK/WOokVOS1qgW1UO6bp8z7/RGvQqCG5jqgRd/vDl3OL6IgpCm0y13cM7
VtAw319eec7kQ6PWxw4WDoB+jmOZuBfZWA/gApaJ27ojVemL5n0XaZag2S5x9zP8EEFAEP5uG1PI
ne8OeD2k3L5xCH/ua4/TNDW6pHZ7PXq0YHc42RVju5x+KuXqFPadIfb/LZ2/87BO+428yocxNBPj
EXZsvukoKckDsjph0weJDJRQrc+r/+3NEROu5RxiZZzpW+iBKtr6Pp7Fzbst8Cmaz38mmwRZS7tc
3N+uuqgyp9czk+44vmvxkKuF3xZuKk5uxnYgCEhEgyL74RZSiwQx8sJJChxNvvWngs+o510TOwQK
q8yDwsEvazZXEHGX9WTzipmQQhYefgPCJx6vPzdfPnjVkJPiuptSCuuy6oqmr1ehzJk/cZEyc4Nt
VxV4kg45KSpyBC0sivBbAmCTlquw0PBSEH4tzcICQTU0Eu7PdECuQeZlBSSB0n0PcyNQGpwMkA9s
3DMMG6ZlvIy+pAYjeR7CFFvGOqKzZSuwXiQSuMGhWF/+isx7ZcTcNn1geTQHYLOLbFbXM7phEg5E
Ql6sVdEsrh6XKtS7OvfZ9IE+skLSZ7+4TCDd2p9xhUOrH327OTvedXpTS9yP7nMce7WFwv5BwC42
1vLIrHlao9Mosdx2DJosqr5x2hi3/tBC7MiXAxiWo9P7quiSpZebbo2yeweL0xvGkyjGil0CyBOh
UusV61w6hxXnRL6rV/ns1E8XL/bH8wSGVvlpvt54TY5lswjbAOf/TVk513fMVjPBu22p64DJGU86
YeQthiX3MRMvR889jyFedIUektSOhUzctIYb+tJ3J9hFb/GZ94JyHdFH5Io7raenhDdOijsfCXpW
HdHpBgMCkh4C7kXBJyxr4/0tReXEpKNk7jSFlxxFfNCQV/MU7Sz9rrqdtEsUza4NmH8FqeG2EtvA
37HSWW4kDA/2YESWeBO4CfgzVJUgHY35flz9zSrIn+IaPv5NrEekHhaRCs2PTikwr1UYNtNFKnw5
tn/cNee5LdBvYtSdE/iMZwKMyh2GWHN2gVwbK3xUaqqa9mnW0qat3FgQEz+l+LBd2AiIMtZ0cHwW
mf4uEn36ZpynDd6W4S8vtLSGRE/uWkZVT8Nk9vB+0IeWvJVTvZt6DdsUDxNlYiUUHppHvagPCpPA
ImcCYHhZ7Ic81lTwCUv9eJAn6AFgNNA5mv7vpu2YaYndrKbMN5Nr2ie0v0L18/UFtfsBxaxMNq2M
TsPdOc4KLv24boQM1j0i6OfWSJGh5DonzFj/88GMF3L7HwvygzSA8lyqOgNmHirVX5VhlWHGlj4A
q5/kWD9z/6kCtw+CFG9ADYtLZXQ8Y5ecgvkB6MxUQcgyZ4P/Bp5q+ofH695S5I0mfLxL4t6I+Oce
gYFCayNJcJiu+RKGMGVsa8v1XF52gAIllHSS+tUMOOheSQBlqb49V6qKZI9P2vP5uQWY+cJY522x
/uqpcc5Ba8ZoHi1NVAurmA9n+UaEWJH+xd5JwUdzcp6e7zygGJ6Fr5VAjW88bMgV+qz6MyzasOR0
2SLhNLSca0bnkwa5+VnYPU69cZuPWUCrCVuu4XwyFTnyEXi6JymrLYmJrnym2AMcHp0bTIlKtmfI
wEt0XrgqcQ/zEEPIm2BQ9LsuArLiR2VycwPHGHOu3ZlFOTCi/APpDUp93mgVuoyF6bLSUY2+eyOt
zerLg2qao6ABq9gTUFHyqLs04uQjMwoQzr994GUhmiNAAXv42b7yp71/VbUC5jNnPcoq20/eJSNw
I0uzx1wjMy6lxjZkivf3rm7fEEXJBLpvvbrKwYY5d42mCKaqDUX1nYwUEzn+xUzByScn0XZULivJ
iToKDURqNMdzYgqWGYPnWHMg8ncRd1HkDcTUsUlDZ5fyK+mOglzoD5+M4oa5N7RorNE3tW839SXe
noU2jjmOp7X3D8Vn5Xp3ezHtmWHZOIZNWFycZLsvM7YAKocJaHb+SB4Cf4z4dqtChYubOpPEVT3f
ISjjpJE6dJe8rApjHx+5ZD0MpvHS4Z0cf31aqi6uJctEEl30ImcPiH7vdVUOdqbHUi0juSkQ9lwh
bmV0WrdN9a6LIj862JIsE7gYKpod4lAH6coEa+OZsuquxYsQE7NXgCe3guGiaIdtwgXt+8gKXagp
h8+wq6C8XWLdyTWNo9m5EIHVCD6LOI52HGKF5HDvtcKe9JlLqa/abpqJaEZW2lIswhjSEajP5GuN
Pzm6kgDBIDa/ckY0DNXS6AK4JttT8+Uu3h0lgjHBCMR29UC3cHHdnbOsPLZ7JGLkZKPkMoZJsHNd
ddgIKV60ZhRQfWGs1pmbbbEauT70KI/yhWXQNhtFO5H7nDA3GxrpwKzQAW9pfwqOmJPlJ1z2Bq3Z
cfko+Gm2bahf8RKOLDahZu+eAr1dff/rdtxic/BfRkXH9Mu0jdcop2sZ6yyRSnt50fjK296XocKn
s7Gq/ohSm+KVM24PPrVbpT2xpRvMq181AYGHNz4R3/gRyhPkINK+316DIiRihaVA27Xd1OPOcWen
CZcOw33op4FbqJF8eSLrF1NuTJbCJyLDsgghFr6AUkDDysjhDpoJTN0ni57mkHlKC73ShE8zkpmB
XY0XRKWj8GtX7BmubimDN/SbrNbPq7v+SKkE9EWgEB2tlinQnQlLoaHTVDSBZNJaAJvr5zV8XEyF
gAYbY18k5ezV38s3UtZ0JlrTHa2F3xyOIz6QNljl05/ZyI0amhDUufvhs6ZlWVcQfiGiBHvaDoNF
uSm8dFjKNcd2BvHT4VbvbQdLeiWr9C1U1w1bRCsxpac9oEXKfi3w5VlNfw5uMJ6nXSQK1/jWpKek
lwqz+K6Mp58w0C7aEzkMLsmab/2mT0YNSDLtIe90RGheAn6XQU8QeBg9jagQCKNDcVFJUmBisJNO
qiawLsWofI/1AJZSOPfuTmvNJRnNximwpHTP7IG6g7hDJIGIEKuQ1YRE8xx7s2UHiUICu1HOLyzE
DMIJJMmEStIA9xlbDh/SfgLcqdmlFj6jMF4sCGYc4S82HvERLijfkec3m3sNFWCKpIVLhTeClXsQ
IzCjKt7j6tlLgNGrFSTsJEbAuuTmxxO6k5m4Jz2Oojlw19ZGgfjKecvGxDkHhBZKeBIhSTnRt+d3
rCBLV+Q4zx/bFGAkdrN+LTOr329ZkxKZIkEIbRMIR1eDfToqVnHsQwhlGuR+TFH156pY07to37UL
n0QL5ETjFxLGAAzIrrCaqJPxhfnPMuB80Mx1w3OZ7w1Dr5jTWuP5VOUFP710RGqEt/xRzin0egJU
3iMIyQsrEtWLIe1xmkEgioCtauCrpk1aTczeAxrOYXc6xPQGgJfMhMi8x/Fa7pxui0Y/4WV003RI
Ywja7YZNXyMIchaCBDw4NqJu9uiwHdbByau5KTYBKc3a+fGh7bt5tPE0KyZjocWu6s9kGP3+oZoH
zfcETQoOIffbzbhmVThDk36MzoKMIj308iTa2L/50NzVf0GA6E+GT0UOf6tjByK/33fR1bA0sQZA
6uZLmlOBE9jCq6ZZjuCV5tfRnuOmmEt0mQyozRGpbzzkRNZ4yv3g3LzOjf5776VjYJQrHT3sDdNe
rWfiLwwBX5yyavNKY9C8fGMnmQ1IFE7aQgWCMl/H47O+B+hIgeokJFpbDE1DL8xA2OwL3Jw74KLX
Neu8JH+GpdfpBf+DjrccnSTxCEHkpwOu+YGr9Ta3ZV3+xtvcAALIjL3g7qleyhKYNonzQ3N64PUm
ZNAUyoLBe8TJzsAPJ87XpP/NPTlxATOvauYxvtnvSZ2+wybRY55Knv5hmDBFybyz+g5BQ+xozxnb
jutW0W7HKTpl2m+WMPrTvF6W56WIz29XpmN0Q8LrO8yMpGvJygh6VJKUSclSq2ber/q1AGK+kwxX
x2toZMpZhKK3VC4a56A1e9Q8ebuiaJsaS1CPn6d1N9jH3hK5Y4vdIwU4ut+EK6mWtV9bM/+eLHpp
WKHHvB/2hBs7Ygjq+ZUqkfno+mn4uX6ozhaEVy74fv3lpJzmnRwPiUbKIwbwGD3e3T13tG0SBbmb
nVNWLEQ+duhGMFZZ9Y+WN51r+w54hwMIKIbPonuLLb3BhM/bWzy5daBvqdb9bNk90uMtVExoJRZF
jKon/nF58MRctHzxsvUTuvqMhOsdtjXJ4+u9+Zbux/H1mMEH7kNhJtHAzZxhHNFgZbEkmogp8xVx
0TJPYOPaAHgDEWNeHBZfD68u3vDKmMEJqG0D7oh91J99ugLkWQ8iXklBNFBen9vHArb89w7OUITC
k41M2f6QmFYZbcFwIsDRepCj/rnTX3oy48E4XMnyiVztvPPBNu1wUXfoZJD7k1IDA/+Hr0CbzacU
sm3CDlssM4hqv/vSp+AJ7Vm/VSd3uE+d+7Lt1uCmYZ2tatc+HfEdDtaG7iPFVuTq1ZWxTPSqm9bc
KDFN5OVT2df4vCPvgfwOs4CLSS/un3BX+3Rg6hKpTMNgD5SyIxl5a2vgtsy213Ifq7q8ZarQWt+4
T2uPoZZxaBIdBrK+dRhTiHq1DLGSvyR7GzD6/B9z0x4mT+z0feSPtjAriqVBtoufRfzTnA+6SBHH
eSHTiu926KkefvtdHilwMlrcr78lERYSr7jyVNwqa4wBB23Ig+J7nErScqN0XvFuySRG2nY+Kmtl
cq7Wcbwz9vUtgg+eu/Yv9I0yCNVcGZlSpyQt4ci3nYYjDiesnYtApJn9vjtZQZhk0nTyBqPXJcAC
xK/FiV0UTyDGBqEVKPnukpEBy5WpM1Hzn96Zrsz0e6Uv2Jz+EAjcjzqkHqFu/oBzufi8QPo5WMAg
IuiSFM3Wz0xDyWQCS7vnCoPK07NVMtiV8TxK3QcUH0rSRnLiEzYg+8B7gSd1AMSrdIqGgbRc/7Mb
0JFfq0LNtvY2oCinqXo+ibp/3kj/mH/NvQP6qzk8ZLpuRjNEnbEgGUQ3E8Q7vQ9Xh691LadNGYCa
qKadDtrYzQAP4/yPwL/cIbjCOLiVa9AAaKmXvOuxXXXB9OfhsjPXfWrtxnnMMVunFh4yo0rPzcXg
6CNsZ8veT0VQMuD7+Ns98l8DbZ307l6Qyt9Z+fPBj5N6nySo4x73FsgDQZo5OLEZyX3NrYKJOXtf
FE8GwA1oKdgEStkUGxhVR7lPNCGvCzOhdGZGC+lxCihabdSoWc/ax8p361fv03wa2VWe1WCydlne
ggQTEZq4UifNZCNMCcDdcxQDfuVIRgDSC5oR9sadtjvBtrS0vNlH41MlK/dm0nkst4P3c2gstC/T
bgGmMb5dKkzZnfdG8hAipm1sjy8x8moajF9RBbN0flg8Szi4jt3OgzTNyyccKcdaIaYidOF8ukNj
aum7KpSG5xZiVqnvv23UVybVT0oVPzfMCSepnnBwiNAaeVGsUHsJlueTYGyU6q5DTg+p8NhiRSH7
ZXeT+uN7hhuGIH0LRdjMz6Dqzs4tT8EyGrOWaoh61RUgN3A0sFDpzh59GUqFfaUyHr7hoQjcUmxT
BbhAml9oiJi07d5yaaMeT/cLQJKpLjRgLuSAK92XIrraRsSFgLX2hT/SKJgpcOvoPFl8gby9g0LK
e5Vo6JoKbHeqkMaybOBo7cLi+kcDokoGn3TDltrXcBEj7paOO6NoN0kUIjctiErdppIg3W4VeSry
YYleMVF+89+67AiIGnkKodHOWQ3Tms+QTiit27EeHSRmufVqNZbKlykj/NuTmzZyF+9qVXtiglGd
ig97huk0b+lfBpnQ8fA1PqRuaJBEIFYkbxmQuz55zKG5TkZI/DRlXqYdH/1n218Vn9ojhXvX/rEL
h3oOjy1T/9k+2X+3J+Oc+qHtOc9KfnDseThAXst2fjlxmxqn16LlnNOS2/q69w/dvc1Gxal9wZio
cB5amfta9QVtucJ7FpAgmMWA6nrdTz5qOXY0qluptEJ+ZtbxCKCQl4ZqfGnlKD+RKFu7igx8AQKQ
KDMLONvlW2EBATfXvgAfe7ohtcAykBsgjam+2c+BOI99/+EBxhW+tv0CAvLvIOi9qrEN0zb0ZRE+
85u1czvr3plV+oM4UjanIHASFpMB8gjjpgbAUDbefE4+ehakJblliA7IV7J/wuYY5vXESBB798SS
Sz6lYMqPRvtfDNUBrp64foqYW2cQf37GJM9KMwXyRTrqzPJQ6Jq0t1RX99r8WsaVlupZOTjbmwbU
1VmjrfjcE+9ryHCnRbZdpfJW3nzifhZP2cY7KRKBLvUfSPz1IvKJpbFAhGqDl7Y9coi+5pbQ2R2m
DZl0r5ma9GuuC+VVIjzMe5j7DTsye7Q5f8+riHti2namsb4uAcHIy72IEEQQWV1z4X0plW00Mmve
X4FcjZCO20nppIIX1rk6Eurx6NY0zYUTuzQUxknc6n/P9dRWJmSPyjlL+H2UuyQWll7/doQCYwpi
UoPcJkfj6Kd7k6SgyCNl/XEC7Bn26VbyUwLq3FNmXHEdvcJHEPoETenkrCuE19+R2QEyrzeZGJk2
TrHFnltse1lgXCta0gqPdwnruBOn9uyDWVgSo3cqq+PfXpVwH9WHzmLNa+jFbE8lT0aS8UjWNDAP
VHpA8r9/ICiEYNLPORDfV2q9gl8VxoOUPW2PU9qhzB+skkdLbRudcPSrnDroDBMCe7LBI75G3D+k
DQQLkDKf9l4h+W1AmpSo1qE+xzXNr8r4gxGSnrZnrZO13UBKI3+8uBOaQoNamv8EmrAla75gjWh3
lQ+63VEs6hCZcu8jq5NxfeC+tcr0Gpl21H5LTWrRMqQVqhEnLc0uF0vABHCZWf4T8wSY8iN3YXSb
sHXDKJB6vUiX7vRHhW3Q30C3vWE23rney1YKmAZr2QbgkbDRnfYSQCT5xJKh41WG1qma9gHKOxh9
mSlaFxxn42zejRuRar7IfU6JlhDuXJj9+j6KWA349Ka/lxFDjESjhbW2TRw5A2lsQLr4huhVlItx
+pa4jyYw9yhXQXSVOMqvnLfoMrzlp10lSKw/HSDjtXl35wWdWZAynpRMneBqJR3NAe385TfPV7HM
4GW0+dAWGkdXHxMoFwuP4nt6fTrIriJO0ugRAVzFOukJisTS0amXPk2X5L4JYuFdPaAIIWIf+9ET
jL1NPkdE0D1cf2H7Vm4AEkzO48ww9TrmTUjXmg2x+KpGPr3DqbELmWC5Rda3KYejbpYKfAwmAHgN
RaAlkno5mzGEj/Xku4PNY3/RCDCLr75fgM0HIVnhAbPHuMxKr/eFgY3NnIBKwPzkN2FEh+HtfbLf
jV+5lgA7/SnZ6BLxyaz9U+/j+3pR4gHCtp1RBF/xY3mn/Uz3WIogAZg5W0lDtoEQRm9YFeqHG0k3
jRvOSFBKmiekeuzAiybRTwAPkoWxIWwN5czQN0I5TNHocZkX7jZj7nOgFKU59KEvpOjwpHPdebW3
vynRkx0jW6r3HGru4aIXKV4V3rwB1cxk8m6DPsVrsA68pPITLpz+pxlUANKnWbhU7KJtB3QLr6Y1
CCdc+khxgqG4Yr1s+9vpBpiNyGCbgjzlaSXngOozTxfMDL7wlqc4rfGZ1Co1dDGxgGWvO2XehHE7
IyWx6NjTvWnkdKK4AyAIZa/cNssatg5CBIWzUuLMQ0FCL9x8WCvq8KbJS5fHsJW+yWgukDdVGR8m
mcBDnYQCGOhhJUUvdnEfFQVyeQ6bIezGG+kivbUdQDem39Np0j85k97C2tDV/6vrKPdcFxb+cq2p
Q70j913UPFPi6N1BaVG2sNLaNLwiONs5ayCk7BFLGJvHVJqBqHd3vX5USOtbMEENlirkngCIS2M6
f43tUoQZQSmph+RRvS3dyCYC7qHzPfCKzHJ4meQYvVRWQeySxHCs3WJHc2YD147ftNDqUNQgh6fq
SZaAtFWfAr1cNGns69AKVzob3bCI9Uku/TaJzWxwUuipvY4T7vGMB318sSFlh4u/swi/NlUtN4Q8
kNzM055+0Ewd2DZOGASUwRVRws9U+1VyPfFrYSkSHshfCK/V4V7iyzzX6SmWGX2egNgyxwNZw5qe
OYnPKu0NV+jlhJ6pwdSbuSs2+z1VgD5kf/SjNVWCV+Vdrpc0+WoACi9wrIz1R7gGKUmrffPpUhaS
bB8+eerFv7IMmVS02hil6Bnx3d/DHpplEgCZ8c8ul7iUiy8Hyp+gla3uDPHfNGiRktqiWcE8aQax
zP+/lzfZWzQRRvG3hm1me8QM/uo8adSwlZ4cfOLekFiCaP09lRyVaUnANeoa/L28jAvUyHZquTG+
TUOfpAm8ak/JbJ1Hl81anNgSln7I5bMvgSOOW/XqXiyt5lgYOsKpsIN+UqQACU1ojJHPUQ+mI2rk
3FIj/JT64xaSiv2kgbTgCHZ7dnUIa8uMgoiiaju3j0Qrh5riDUjmb+aCzo43EPSHBfFZ3rNAICaf
YldfobkWI/tKQODnn/3VAFDhCzgBhJY9fafK9wkCYy7VelqJvarEFBqJ2qA3tSes4JGRHfGM9Avu
EV+lQHcq+uzImYR+cCfTlD2SiOJZS0vT5TVsOi0l5t+ja5BfgTtxrqT0DUOIViiXT3l7b9MdRj+I
iE5ZgonHwMlhg9d5r/yt5tJfhSEsDfb8U+6169fGQYEChiGnG5GlmhHZJ7F61yzXTYmCpfCBEPkM
l6QyTAyQNCu/JoNjItC6OA7rBT7KgK6frS2iGB8TY2Jf/bHuzL7WwP328qBgfaOp5+oHfdaV5wOz
x7LLzGgEhh3JjuA3iKl/HtSXdcn+X96Rzlw6grDR2jXpPLv+LT5kuVYAU8GysjXt7Vhm+IAaODaP
dS0IWMarEEAChrRajEn+flGaXnmhZi/T0URT3V3koPYMvRqhzZITYXbU1GA7vxxmZ6OM7n+U/53h
4l6Lde99DfVU7H/UhCKanpEtdsAqfD/E0sOdACwSu8UMP9k6KWTUniVKdqm9mCRMqb8KBmK3UX9x
JnTJmK/RUVdBQ3wi206iWuA+BjCkx8YY14255KxxhvcpD21u4qLA53VZhDw+IclrhafFDqZ/lWBI
/utr2EUcgKGWtm0uSFab3TxhBfDT7CRWoQeRGlQ6Y78gNK1mtr4Wq3uVUD2mfhBifYjU94DgnNFZ
WUgwV7ttghSIGQ2JJAj/fSn0zxT32P3B8Qy65FTzXqjRWGC/QoPqXbpEqZ5wcc/W4V8xcv47UPNt
5wbnZT33Bwwsz5h+OXaXWKextD7/lBtR3yhVOeHjdEa5J3BHeR/HGUJD4aiulF/b5Ca2Y/bEcvuM
LSi5ZCXcvWeRIB1rPg2aDumO4fLKClbn0eTQb/c5azJ/79SpdXyUeFeXEm0NuFnDnXZx+SX3C5pi
fxRc/VafK7H/GtfnObYecb0BjudBAbDIclrPN7LhIwwP29pcXevlAKXd4ij70cw93fM9Qb41FTYa
JdF/HF65bq4Hc06ACDTUd52BQ4uM0qq0ZpNsTUY+Zy2xdPfva1o8WB3exTg8vxQXgaTKtOtjjCVB
CEJkQRfG12CFxceGbdpBoR9VDk9mjPoBiv7dfjCOFOC8Z9EzalFwlLojditDfdbc/1vYE1Pb9Bwc
5BQJYl/kuiG3iCrZNh9vccWxXUK8wacm5yq9chCxas0TKSZgJ3Au1lavlBAWgyPBvEcfUgjJ307W
gtilfAU24ijFP+Yb235y/Id1dRPcTQ5iBEePE5nV5vF1sURPPLkpCeN0mtPGIUnluVweF67SliSl
/wVmpxG96Goe1SlBRyoTl9+Hv78H+MzN51nOJAXMLtjHw+Nxd4SC13Gp8iXdPxRSyvg6k143WOFx
kc8TiIY5CuYC9bldCoewyzTenNTBiVBjOjDk0Gtr+lJ5VtWmgtF+bfIcQfxVknJHSIDh6yVVeGfi
6UshvCIaYrbY8P7M5A+w3azfqi8cDffE1tIuGXOGfhR8b71ZbqBwEDUvYLPtLO1C7NTrvvL0RRIO
aypgYcE/Z/dcBgYEwLUf8rugbfoVT7MHdQNQtDtTiqFBALzO4JhJxTUhH8Kh8aRUrK6cIQ8MAPDW
5qHEi8PDzTSr1DKskDsE/w==
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�t��yгwH���S~��t�U�͇Z����F.{�P�C�a��f�,8�yM&�	h�WGO���s�(4(Ⱦl���^���������A�F�!.��gT鋝}E0:�ڡp��zshh$;?�BY(U�,���z�̆�qΏn�M����jI���R~���W4�I{h�Y�#n��H�:.g�c�b�P�2�C�۞6t�_��/�;�=v6�f4u`�t1�����|��k��
y2-J�G�R_���i	�\�a�;��)�e�w>V��(Mb���6���"�=��PW��[�b�~��;?��o5%�QQ=f�AjC껌�i	���k�u�T�kYeq�P@�� �K�+�e7=��YFS|��(뗰`�Ê���F�B~�>!SB�,`�-�G[�
�a�{�TY��뫲��;�����/?4لҍ
��	bo��&�a�a�h�Y�=�]8�w���G�^��%#ڙ�?Njяn.ǲ�t�[.��9�-�u&Ky�	0�2G��!�-�;l�� �H�T�����.cl�������� q¶G�S������y�C mm�Kz9��m�XL� ���Y�G� �e�Ѩ�w�'R2є�ohXg^:�?���$��?�	�A��![�ϧ:0]�H�ZƇ��������Su��ܑA���&�\�hr͋�R�Ǜk��K�ˏ��B���Zp/,=�.)�6|�v�񩅨	�F�$���7���WrT��aE�,�+�:��a������}���.�e�Hgl��qWB�����l�#XJ����Rt����r2t0��T(�$��,�m��y�d*�R�p
�M3؊$K���ā~gu���
����M^`>(�4�f���X��(�=���3U�ɜ�F1A�ܲp�&��*��B|:�HP��ڏ9E�#ВD�rH�nr~f8�u�V��鄂xi��\��s�1�t�怠�zM���\��k&$Nf��y`*�o�y�����{�_~;���+��.,�8�����Mt?;� �;gp6K��ޯ�q/���Q��N��(�Uw(�� �'Fj:�/:�T�.�{ Hc$�x��V<F`ePe-��"u���Хxվ�D�̨��mc#��\~����yc#�y`���/z[IĲ<1�Ȁ��W��"��Y�u*L�$NOC}�8�E�qQj�v��e�,�����ś��%��Z���W��|E����9�� ;�?`��%1d+A�Ɨ|�6��t�X4e���H�X�n�Vy���*V��Y[�����-��\�xq*���AY-i田V��G��I���Y�5��eI�BRzv���	��K�_\=6ԩ�1�y�R���_�6r�+�T[�PŨ���Vk�~,�E(�ƈ��o��T����#���	���/��Vs�K�]!O�����#�W�Y���Q����4�~5L�%�L:Վ���+����4C ����t�ˠjr� i��|LQW0.�ځ�d4E�T�Q�vlm��$�3�N`,/%ﴞ�c���XNM��F쭦��&�n�+��$�; �lK�P%pϩ�<Z(��n'��
�;7l��j��S&�4Gۜ(��Ɔ�FC��Gt,��{\QU�9}·M�Q�~��4��Z�#m�вԢ�!�/�`��޹h��v�V�W*\��nk�7�������yZ�>� KM��wZ�6^bMy��*�gT�-��P���&ӆ9nѮ����:��>����c���g;p��2_����$��o�F%i�װ�x�Y���t��)���R��M
���#��ѿ�hľLd�	��r�I���L��4U��������=o�f��Zw��3Q�E�;��27�)r�"�S;l)�!�
��`�Ù�8x׹�v �]~rn?.���X��L@��y��:Yt����.�w��!�(�VODy>�Fe���3�����D1jm,*$�1p�l�Oj(e�H�HJ�][�KgE�����$�f�=�]L~�uZ�ӹ�Z�����Vn�]�v���S<lp���,i�\ٔ<����Y{v�Yc�m�U��Z�pU��9H�/� �H��� R����<��f�b�-湩��A!��Uq���}�g18&�R��'�G�� �|D�0��d =��z,����Xc��ю��x(X3���w&Owv��Ш����̗l�·�KǇ4%���樓8��R�*�ʁ�⣼I���M
{�4_Aor��
�_ͫY7D.���(C�bm,h��׍�˷�x)h椞#(�z�ʯ��,.��d �������(H�g3�D��*���m�#˹��{�X���էl�$���3Y��Rp�MK���q��h5�Oȸ7�_��8�>OU?�7�|����M��b����Ov��R,��4��zu`��a�|��V���`�|�aҧ��]����9�Uc�}���I��އ�x���ێ��e A������{<o����q�E�����
?"��w�w���tT�d;E�#@U��u��~�'�,j<�Ed�N0���B�k�{��OF%�Ks�{��r�ф�I�)��UF�R��(���$�tBG7�_�c�)ݏJ��	��.�Y�qP����{��g�=��"��� ��ڮ;���k��T���7�"�(��Q��C���jB��#�`�^4EIc��,�e��!/$��������5/f���N!De����Ăhy�o���x7T6��a0�y�w�Hۃ��]%*1���m�e�kf�'��͚��#��;W���R漟{E+st:���?W.�-��!����k�Lz����������Ϡh���%	��e<�Z%g^�rLM����*�>�5�A��D3��
h �~�6i\w7�!��NR��B\�.oǏ�T5B����/w��P����vO�h۴B��9(�o_oqy����Ϻ;�d�nX��ƣ�	�=��=*��J�Hg��b��7���4l���>/.r�������xv����Sk�lб�C���Z>0��=�p�cmC��D�\�.��O�(>w�T�v@9Dװ�#�b�	"|OU�K�+��ȍ�s����Z'Ƭ��E�۱Z���x�18��u�'���f�8K4�?�	I�Jr�a�(����Y3&�����	�'�ڨ��Y�K�m�P"��3&��W��.ԝ��c����l�K�>�HO���]��-�Z6�K ����e܍�z O;��q6�K��w���Pkݲ8 H�6�ئ�8�IC�����B�,�X�^����f0UP�n)ճ�ġZ�|�/.>l�Fyu~����)u���B�5�읭�S���~4eTE�R�_gv�,���\��#[%��xOCH߸�%��YJ�|;(�ٮ��YL(���D��p�a����<�=�7�g��n䁋4���2���,՚7֏��IY�e�e��	h6WIo��_fk��e�-�b@;���^<���zͿ=��2�������(?I˪�FEÊ�����?I���_lDbx���|?]OMHZ�Σ@2^i���/'�Ef���8�N�t�f%e��=~�
�JsɅ��b�Ռ; Ih��X�j�;���%54UT��Tz����Z�L����������047��ƕ���Yc�9p�v�,ZX��̖�͹�
�뒙�X��r�|�73m�m�ЪH�J��M�3u�\���*���b��^����;���^gǝ*|������!cd��I�pْ�Xl^5R4�6K��rY?�l=_�+��Ǣr�SJ�r�92oU�z�#�&��U��⼙���aW��gNx;-x��*oT3�K<2���2k�,�h�;r���Xb�h:D^�6�����3n���q�n��vG��+��Nq<j�X��[�jI��$�I0 ��T0�`�ihO�z�Q<9J�i���~9�C��Y�-�@=�v��'�w��z+� G�k�u���As�g���a��Iu�����|�ځ�_���ɼª`OQ�|���}���J*�>�d� ��7�+�H�p�NP*��F�"KjE4!���(�a���e@�ZL!���՝	���W�+Nz��7���q�Zm�`E J]��vd�7J��P���ק�W�cl�hׯdS�`���k�{����Κ�JA&��ݡ� 2����,u�I5���4G'�x�u:h���P2Q����4E��%C��޶�(OB,�0��}�0+�N�ᝮ��3�;��uEi`��@�E�7S���^5��ԳE|\r�# ��� q��j���o�ˈ�B�
ȼ�ـuر�NzLg�\	E�`��[!3�Sj�y�����-o�`���F����o�Z� ����r`��è������*���@?
�D����`ԉ��n�z����[ew��Z��ҍ�m�e�$��i�sJ=̥�������L��U�V�>�}0���LP��0PxG��%g��mxȋ���ֳ�_�<��H���#^��$�_S��N�%����@��X�{�zE��~�g<�cxِ�FJ��Z��܋C�Ȧ��_�6��7��m$Ȧ
'c���|�u\fS�h�Y�
��Y�s����y�/e�ld*�6�á���+����
�aX��3�󡊮��n9�#3�C��!�IB�шx�"��J6���Z��$��^MY�Q����/\@�(m;Gl]|~���
�#�O��jq�
e'U1y�-(�N��r�q��"I >��_i��� "��R�dN�;�5g�2
 ��	}Q�]Ǥt����{��4��C8��@̃�=��)\�e�ѵ���YIaf;��J�ۮ\�R���>l冑l ��J*�{�$p��	'�{�i;ƞ\�����sū�����T X��|A.X������3Vl �7�	�U1D�~I7F����>Q�#��ԃCs0���V�Cj6���{T���q�����7�ɝZn O��۴p��O�	p 
���N����?B�u�xr���!�ְ��j�=�����zY���U"	*:�����@h��NKg�_i
qR���%u�)j����1r��/���ATF�d0U-R�Y��H$��f�"��\�0we������%�%M/�Bw���/QG8O�/R���M����Y�sj�[k<$d��ڽ���Y���[�G�G�r���"���k���;z��2��4�ܩY��	�լ>�j���p��I2�����J�a$}����U�)sEl�59�ʤ�W���k ���
K�7%�,rv�}���ǆ�Tm��%��lsм�����	d�����Gt����x��"y�FO�įTU�;�'��X�\���9[m��g��NY
�W~;>��v3�uW������+�8������A8�{���t"��Ȗ�O{�碌3�������]��Z,�v��}
�(�������%�������L�y���IWꈕ&>l��S�X��-��#�t	c�^,���WT@�r<�x��j@�t�D����aaF�1��寚�.<Q�-Q��Sղ�ûb*&���&�mN�����g�R�4�6"��UNWN7�`�c�Y;ީ�vҀڋ�����+��d�*�R��*��LΒY�<4���2��֢`&K�D��U�)���*Me]�;/	��`(��.����tд����� �f��v��ډG(Y�[�PUOA"�ڎ����˪a�p��ܡ!�����:��t���>"ԣ{�7-�
����j��Q= �S��.���8�:��iPkH{ksr���h��0뻠��˼IX_��1�^����h{�,5dbV4sH'ϧ?_�X�rH������7�1CYY ��	k�Rj%o�r)�4�c���^-�1�sc�aX�7�O�$�CbE�*�Ub�(!i�#xă'��js1ک,COY1S��F��~)�o�1A� j3\��L��������r��')RD�IK�x�� F�ۖy�	�Ǜ�{o4hq�̶��b�μf��b�I��2�\#���K��'�hpA�01�`��=X뺅J���0v�Z?)p�be�'y���I����.vb� �:���m��Od7�4�$h���k�A�]>���2�9G9����iÚ9�^o�%G�x^�|���_ "K ��:��C|Ym�:8�L �o��b��|:�ߟ_�N���"��,Z�����_���Z���5mBy�[�D���mU�4ǑM&��8x$Sb`F%:��[�:�S۳�<�#�%Է(��`�3f�b�|M��eT
o��KRn�_���.��o=!o����X���8�G�#��@9���RB�S�0��8Go%��,L��#6���+�ҧ�0R�?�P<2�I��r��Σ`���Ӌ����a�.,I�\"���Vf�	P:݇V��xB���>��)���x-5ϙޖx��%�s4�k��6:֨��8��IO��<�՛g/}.�^k�ir�☕t:^���׎�!�zn�Zc3� �H1��ί��DZ'�:�}ɴ��*���<v��i��_}\�z�X��~%��t0̻���� �*��{�m�ٮ`i��.U@�~������&��&�=�%i�T��;O���#�}T*���4��@�����E\����
g��t�����*�@������tFn��R.�|uh�S���K����	�X�'�T�1�+�����'��t!�9^�Ij���0A�������AtpƇ%�)�f�jb]'6 oC�M�B?@AC���d.����%N���%���爴�2Ĥ�Y�y�]B��-N����xBɖ��RrR�G����-����f�U����&�-�e������ )E�
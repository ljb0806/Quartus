��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�W266�T'�ۈ4/$�M�����h���R#��$-5;�tC���eV�y7SQ!��B�?S�Sj��Qv����N���s�>4>��d�R�&�K
���ڿ�23p�`M�3��And���CO��K���A�Z@���:{�����+�me	�L�cJ������v�#�}�H'o ��4N m�7� pg�v9Ύ��c��O�B��o�ɩ)��2��t�H��3���R6��'�ѣT�(G
|6��+�ʠ��@,� K�7$bF��v~-!b�yr+%V�té/u��@zN���a���?+`W;a��2�3�gӫ��AÕ����:��/	$D��v�ߘ������/����K��f�m֛Y�i�1�]ME�/O�1;�QJ3�B}����C��Ғ�2�P����Lq3
���ͅ|�!�2�&��(�]��Qc�����y��b$�VE��i���1,_�w?v}��5D��}/�i�#��m��=���Ա���o/�>�
�̓z>��ͯ��SPb�����y��?�9�~؁u�q��k�"�<Y�%|���KF1�q�4����r��75o)٤X&զK �V���T�tьV�| ��xW7U�Tں�"����b�i��%\s3�F��w<d�����>r�Eˤ��#L��NkX�t��d���6�I�ױ��*\���z���R���Vhw�F�_D=��9<��96���k�V&���E@ĸ�q R��;�xF[���9I6"]5���ɺd���:�N��@��ź������NFH�%֙*��Z�P�������l��(8�v���E�@��ſΕ�c��pT�"��#W�T0��%<HĶ�DAx���+��M۾�p�����ݑI�4���o5��I K���:�|chH\��eUz�/�̑M@`�D@��~�ͩԤƷ]-�J㕙�O~.��>/�2����Ց��o����7����Ux��QivL��Z�!�=|��yKm֦&����Rj�6�����V��쿠a5l�? E�Cߚ�>�*Ի��)u�%�_�gV+�Ɠ�_�^ٷ[�Z�P5�P�̨�����(
PϨΗY
21�J��k��TĽ�{s�I�1�o�ӧ(��db���I��Nmu�������Бr��'lGޛT�ŝz+��&:�5﯑�&6�m �v��3���%��ަ�^cY��	���|s��l�۠@�>۱���Q����̲F�-"1����Fٿ~��w.���J�cL������r�����T=�pavB��ļX�;H�v����QӢ��h|I���mbIQ�����.������Ѽ�Ư����i�����K��X��K
��f�H���� nR|�j,3���L�|�W��nt0�d����I{AГ#T�#j�O�GvN8:�3t��m!5vv�~�c=�C��c����SvqS���,� I3��HqU�h�D�.s;��<D�U*vۧd�V�l�K��-���]/��f(o,��^�ˌF�%�����OK �J|ɐ��*��e�ǘ��}[��tu6N_'u�G��O�u>VTl��r����D�̚� V���3`��;�dg��JD���|L�ìb�X������A��'����k����L�~���F>�
��r��ʬ����ܪ��5L$*p�\�R䰠��Cx��7l�m�.�Ƙ����]�H�Z۹f�#@���#骽�ER\�3�l��%th���PNE`_s:�����^��7Bᆱ��̪��V�E2��$�YO�@<�l�2�iђ�o���ԟ��7��8��w/~�"G.ꐤRH�Y<������D��lo�~���'�bs"��=�%�7ݘg��Р#\���E[���!P�4&���ݣ�Ηx/�S�iB��� U�P�3���گ!�Y���ͼ:��&	�%�F@���s�p�<��T=m�Kb�Bmc��%���ޡc�q�Ι~j�:8�%�i��4�֢�q���t�k��yE�PI�%$C�t�k9��F�1�q�)��/:C�z��,a<#�H��<lD�FNx�'���`���q�n�t��51�u
,[`+�'_��������W����o��wT#��S��z�ֆ� �A�Q�19Bf��F�c�	#��S� +�Q��gW�7;���"_�8��H8Cx�եO��?��*1���2�B9����C7��=����B�H:*���HiE�d$X'��eG�\@����^&CC�.�7�
�������}�\��iɂΝh@n;��н�!f(�t��s��ϵڽ#ܧ,�6�MkJlc���z�5V,��B���^����ؽ�*��,F�t6�]��rӗ��{��:a/#�r>s� �2��:������:\��UIP�g1�LwϿ����� 	��EY:j[�GH��FԽt�V��'�!��u�g*&l�\
	K����_��Kk�U���h�k��6�'w���p,<��v7 E��h���JH��Jo'�N��[���VʥLm3���b7�7�Ӎ[1��7
�N����÷p!ӕ$���A�N������ 2.�=A�ɋdB��q�4�����hp���k�T9A�H� Qx�B�lIP�pa�����Emݏ@v"@*�?��1����;�a�L�f�*�q�;�B|��oګ�zrJ��ID�Y����OJ�y���W����y��.���"~]��ݖ�ǡ�8^�SM���J�Emĕ7�@�7=�b�?L�]������S��f���V��֥��cz��CG��+6��2Й�&vǄ�Ϡ��:�f�h]1��H}������1��P�n���8Qh�!G��ūׯʂ("|����Еp۳X��6�YA�ѻ�4Z:�r�!O�����5���2��n���2�� ��Ǩ�N�(�fb{ ����݋�Kö�}�<� �K����Jq����EY֭d@=��D}���?�����j�B@yY�F����4��
h7$�������1��zdh��]E��.�v=�Z����#w>��X��������.��\�`��O�6D�I5�-㕝�3�L����m�<1$u�i3F�EX_��	��m���_���CaA.�eWjEJI�(��+�Q3ʻ��Cz:���r6�P�u�m�%�G�P֯�w|ڑ��;�C�{xu�������0�D�V�����6� �r�GtHɠ���B���O8��/��N���9�$��2�z,S�WW����b�j�@�U�5��$aw���
��$�:tVd%釱6�`�L�e7�EW%�d�Y�ɍ~�B��jt�SF���R�!�?�l�s��Wc9Q,�Ce�?wG�|�"����J^+U�"˭X�s�n,I»��j��Y>���濈�0PqKr��c�C��zj#�����j����1]�=�i"Fǧ�Vd�qFG��7��w�D��Kx \��PS�m2�?G��s���t'��C0 ��ыDS(��0Z�S��ĕf���(�c��!��ˋ��q48ֈ��R/
� ����s����ѓ��r�;��d�~�����:��؜�D6/8h�.�_�Ս9�Y�L�Q�{'�������6<8_!6�x��~����w<�BJ&Q����"��0�t����Z��Qࡆ�eEI�l�1���P�^n�Ĵ)�])��0)�9;�@>RV!�:��\�[*o�9����5!��cO�(ձ#�"������Jk'������NOk���k�F��V�P>�fj�&��0:���Rޏ�G�y�\)��rrJ���C�
����pW4 ���-Ԓ~�q'
6�
	�fw?���Ʀ�v���?qy-`�I&W�P;1������;t �L�[ Z����SoYu]t��]jӮ��+�ʢ�Gj>�uϚ����K:�ү��ݖ�(���>��.�ԗI�y�ɟ��?5>j�ߡ%�2(�6!8�z��h��:�������\�"W돨y�q��m)Hpl��p/����:֡��L�D�@G;]UF�[�G���U���s�m��/*C�������o�oȿz�̍��f	Fm��φ�ق���i�<�l�rGh3��Bɟ�k��|���N�_�獓F.�:���=��Yj�/���R�� 8dC�zUJ��/����VUa��l�<��X���H�Cz{G�T�Kc��;��u�b�n�JԵ�X�M�h4ڪ~��9r�zߞ���T�EȺ�uY��y���8+�L��J&xc���`A|��)����6ů�M��	����U�8� �W�V�!�����*�,~b���U��ʃ
�w�І���K]���%b8h'�8:�/�T{���q1�u�T���SHiT8�N'4'͢�x&�Ӭ�>�L*�n��Q�;�_Z�KM��n|���Y,��ewxY�}��d���ׂ�#��w=$����֊�=�˳z�/?��5k^�(c_�A��� x�-��v[�-)<Bƈ#h4�:��{�Hg���/ގ��w�Iq�(���
:�{s�z��
A&�*g
��I�)~P��ZQ�H,����)���ogB�F?ʌ-����,��T�"&����8�,�y%ڎ��󣸪��˭���`�O���'��:-�ڙ5I�g�@>���ʂ�����ͧPFl���c��q�
�c>��S��ё�t����YM���o5@����C��u$���rȸג�,D�̜���L�6�U�x�2b�e�؀�S.0�DI�[��j͍�{u���mM��F��V���O)�@X������ �������2�� r�_%�տ�^�X�n	vMi����#P�[�K��%+R(��֫hϓ�����hb2y����.�b�ܚf��s-��X^�9��9����bEղ
����x�}¡�$�	7g���g��B��_in�aﳧ`�A,s�����@��{�>�:����v�`��D��TK�W_����Iŀ&�p��A�>�n3��'ڄ�<7�vj��P�-k������{���{T�
!=�}�L����s�!	^�!�A�;�_�F�5�� +���#�tZg(�Z������&���-�f�P�А ����h��救�yu�;��ko�Y��E�*�)����CZ]����4/��8dy����'��ei��i�F�H���!6�#���񎑍���V�M8e�q�D"����A��V�˓�<?y���g3�<�4������f8��ϳX_�9�V��X�P?r.a�~؏juJGB%�UZ��35~��Xi#�2R�ݘ��q��Q�pd^�R;�E|J<Z�!�̱���hk�+FX�U�M�H$�9�����<�tX�8ُ@is���8�I�P��,0z�b��Tl&]��A�i~��B��5E�̯���
��h�n��;[-@�œ��H� ]�kl�EgG�ę��r$+$�\�v�mS���Շ�bdy�v�3����݂�S�)An����.�m�{�z��9������Y��j@jU�،�|�..�
b�{��i��M]Bi����
rū*.��y	/�*f)��0C�� ��1\ۇK6��\m%��Mr_��X�HЮ�Ԙ��K��.3!�؂���B��C�Ye��� ��J4����X="c
�Z�/�nC�ђ�@�=��&�8<3��M"�:�R,:S��C"�+�9ʇO.�e���)���_i����}|
�Œ�����w;�v��������#�7o�2=�KE�9W�YH�;��FG��)Gq �j�b�}�V>ӫ۞��iʝ���>':ѥy5޽"�{G����������v����{=�5�M�	���`�j�K+Sb��-re�YS���	($� fk�[��p����Tm��Mh��A��=��l"������,~`�dHi����m\b*�_�'>8_���i����n���:���ƿ�O�ƖGLu�*b�w-}8�"G�E��+��k��X��:B�bRn!p�:�^�C9������{#R����ZN�B�}
{�}(��ix6�)�N+k�xa)�gk�i���2�[��d�ܭ!x"ܡ�g��х�]����8��~>�1X8����*�;{���1�u�@؇a�|��ZF�ʜ�@�!`˹|�ז#��W�Àu�c�r��=ER�q�܊Ŀ�ĈV�}@����xq��o�"Ϊ�OO�.����zx5cv���
��K���q���g��-�����E��q[�?[8�h�>��gG�ڶhB� ��@Ob��q�$���U�-@j��J�M�UR�Q�C���h�/[��J��^�I^I������ɓՕ��2�����U��ｴ����7)/<N�����>̦	�ù>9���o�<�Aw����9�$�S@GIF���+�[�Lr�Z������9�˗�{�9��p�է x+��2�����q�����)���y<4V_
i	噖Q_������6?���u������BNu�劋�\�}��H�)�_S��2���7u|T ��q� {<G�c�ޠ�#��Mɶ(�b�hFv�\��ө�Wǹ̖��iZ���XM��	�A��@��$+�� �L�������,���&g��G�R��q-r������F`m7��,9��)m{�Ѥ|�gUk:�3���~]i��+1�J<�u
�P�x�RE����mq���.�'a��H�r<덢;f�7Y�c����h�b� %���=QS�&���	y���0
��8F6F�ڬ�`-��תn�}�)y�;��lQqO�:��'����L�q²!���'=OT�7=�j�B��3���?{fg���/O��>4rǂ�k2&���	�p��O�/t@����1},��i�S"e6���6#҈�RP����U�-R�±���|�].V� �~6��
���ZZ��kY����?_p�[��������P����/�5+o�Q��ř᝜�(A.��e���3��q�]�[�U�<�첲g����X����=#l�MVbL���K����à�����$�����%�d5�z��*�Fo�G�MY��e<�d�����j8�l�.-�k1��&"���4��N���W���Ht!�>�`2�6�?�Aq��D�jk���������Lڴ���V��d�a|LbZs��\lC���7��f��Ք�UB=�΀.vL��p�h�z��yZ���֕*ϭ$wo��ِm�lڈ���i��ԙZ��3ISv�%�I'	nr���ZA@���W� �|�U$����S�{��)��{;����ڟ+�j����)�D(PKI�kPY�g�+-Zs�14�\I.>E��-R^���ɗ��u�
�ܷ.N�N,Y�P�&4�:n�axr���F�{=۽�S�� �X��T�UX���#��=D�#���Zy�0�L�$9��w��m������� �bq�5�[ƴ��X*��4�����*W^���k����g�1�çY�l���)kM^�׺������J�����~�_��\:g��b>F��,�g���w��������OI�!u#`�IQ�FH���c�d�%���G�#a�s��u��D^J�0��D�SC�.p����������Ks�;
BMMM������8����E<���q��P�5�KM�����v�r y��~nf�|LBm#��K��b�ӕ�~앋�����ȢY��Y����4�E�yY}�]�n �},�^\�rT$c���*\I��q�Ɛ��ι�?k �gPA��C��x?i��SL�L��x�v��Ԥ�D����I�M��'�� ��7Z��\_�Hxo)�̌*#{[-���)=�bv0�t@�@�qƙ�0w�������9������麊{J�a)�'I0��2\�}��1�-HkO{�!���h!t���p�A��E���	g���Wޓ���ERf������.3��u��o�֡�\�͜�a���J��͘J�6��SioO+�I;�V����<����h��G]%�>۫j��1�
��[�9�Z ����&�]��ڲ��Y�:ށB�V0�B�E���np�ׅ$��:��<�|Į4 �y�
��ށ����e�BRdR6 �`���c33*�hv��N���|[��Y��Xß��9� �N|�2��������)'h�6�a� .�ҍ�����0���E�]Hw�mY|�?R�tk[�|��*��y�%�(�g�	�n��jH���v
�@;��R�<� �=�a���q�͋>^:O�THZ�SE^���Ep�?;o�������Ѷ_��� &T��{�2�w+�IG ���"h��C��]i����?��UUU��Xz�c�I����p�>\B�\����k�_}!�'��2-�'���5�IΆN���I5��hm%�\�kQ�}{PS�{��ń��\�hZWQ~Z�Kl��O�-��u��
�:��6 ��ʢ�����;���N�˙�<*3%���w6y!�7w3-�'��<>-BNj���jx���᫸i�LN ���K���'Eƪ��ּ�F�&� "8ţKN���aZ��j����qWR�j/$a�^9���q��><�?vM��f��~�/
��e�&]�i����J6����Lc�ß��%c	=�G�Iσ"��a��|�����Y���lDh���������4�	�g����.�������������	*���N;�pD�;xFICί�����-5���43�f�rJ���2�~F������cg� �&�xa~"��B�{�߱.�Ed4��aNĝ�ә�ltl���M �d���ӣ����I���H޻�_�⛮QE�ϘV�f�q$
�B;	�eX��*�/�Y����R�c^�h�";N>��Խ�r;�mZ\j�oU���QY"���F�� �5�=�Z����?�Kb.;���"��m��NΨ� E�!��4�a3� (��h+9?���FH�;��Wu��_���0i�s��:��:���0��%�$���f�S~�t|{+!O�DUǶ-hP�:`����n%Ssȵ?P$�D���ۧm���i�^Y�!��לǧ�S��I�����DP�b3b;�l�5������c�/P�}^�x�<Öu'�ln!;x��3���w[�K����\�f�8��U�;��t�#4���6�h��_u�Y@��aϐ��E�r���ƃ��	��$Kt�FF����$	�b�[�|���oˏ���VQn��fI�<��F�W��.���,m��˥��7"��M���>G	���x�f���dUK�Lu�P���@?�D��dB�M��$(�2c�+��#��&}��Vxo��% ��8��������N��|�d<�B~S(�`������Q�ݯ��re]+W�J.� ��h���q�%zr�療&�nc?�}C<$���hGf�K�@z]B|��8��	\�n�K����NZ4���݅Ej�C�2�Z����,��Hbz��w�l��q���Q�9R���OAhn-��+5P0C��l�!?Ծ��F�h޾�1݇����D�r�U��BI�EO+�a�L�
��I0�z�LA�WE'1�U��rl����Uv�{NIĴc�K�x��o�e�/��Di:�h��a��m��g��� zd��Z���l��L7j�-棾0�:p���w�ʚ� 9f>Vt`����p��&��\����qdΰU�2:i��Ξ=m��@�g_j�:X�ҙe� �5�{h��:��J伽��|{~4���H8o��_2�Ԥ���Ӿ��']b!=�y�y�� ��`��=:ѮlS���V��)�y%�9хn�;���"��-�o���l����e�[{��/%#��0"L}v	MXu,ᘍ�D�_�Ŧ�`U,doK�f�-,��㯝rU���i1��!���ؑ2�I˰U���>�4��Ji`�ϐ�'��!�����K'����!��O�[���2���B�������\Ƕ�B�%�Ex�;���!���e\=|)sDߡ�pv�����°��������dK%K[�8K�i�DSZ{�zO�p�U�;I�8kB��y��t��	�.�b��$&�L�!����E�r��l�B�=�ξTɚ1s� ��RW�F技姰@³pl.`��:%�����m�YZ��;�Iew�5▼�ː��:X�BR���B�`����)g��u��^W�4:�X�aC���Ax(��=ĩ�T���**�$�$����	9���o�M�v٘������'Y2$~�%0����a��DΏv�8��=���CB9�������9!?�����
9�R�%�m�8�A� �;�~xօ:~<T�!�{�|���f�M��[��Y�4(D�?O�����@D�6th>���,�]�����#�M�z�m�Z��&3���<'��S˛+M˜A�Q���Q��8t� ������R4��H̘T�{���1$��Ҵ�l�w&B|lԤ�<��g�u�-0;-|<�pn\Gn������o��ʙuyR�bʨg���#Dv~�s0��.�sL=�� �?����/�T�e"j0nM b�����2��-C����q�e�2������a:u����w\����Լ?=�{'����|Aʻ�6���~�e�!��U럫�䒲���&B�Joy�ڃ�^P�JN3�fYO+�W��|m]�W��@��Ҕ�D!���!Yv*�pG"���$����?1�2*�g�;�:\�hF"����hF��������vzˌ�\��s�VNڼ�0���}bT��5�U#`*����J�/�l�F^�~�f+�YU�>���ET�&w�����(ZΞ�	A�@�*��
�a�g�+�A�g⛸W4$Dc�7=��f�g_Ej���6�*Ϧjڞ��V������Q��A{%ͱB�Tۻ��KY�C:�C�n1'秄E2����+	�f�O�̲e\f]Z)��O��O�k7*�NK	e��Xp�l���-�Zy�i�%{����'��g�hc'���}�j�mZ�8�R��x�"!as��ë4q��OWfS��	]`��m�,��2z;�� [���<�ε�<�5uD�l3f�Z�����nŏ=�<@ Ly-��9��Yn�X��]
Q���T�:��n�=��diD��{˼q��#d��iS��G�~f�̪1�B:3	�2ŭ�nw�e<�T7�<���ZF�Gy�U�zâ�2���w�4)	= �-�c��P�eP���$B}��*�ѻpmq6��-�θ���C;df�{��(s��� _hM�i��5-z��O�\ "J2�b�R�<������v�����C�V&� B�9��/����R%9�q�����Q����㿥��ތnO�m޹ �WF�<��~L�g�N��zE�B"�q�ҥ��`����L@;����(!b��^ڣ�0Ɩ��z��N��v�_Zr�v:�vL�z(�y2̘���m��}��l�eG�Q�5��7�2�\d��*�B-��,Gy֯諵�*y�H@;�]�dG]����#'!V"�gK�l�c![�ί"Ҁr��ݷ��e_�[RA�)�<���]Z����v$�2H�WN<p������n��j�-���ۢE�N� W~����'���e����q�u�-���QJK2l޵T�����4��|G�����§`rǱ������y@r� ��c��������<G�
�O�׼g�(OmK�m�,���S���LQ�����u'�B��-����p`%k9�sY��w�e� �v;A�^��W����ѻ5�Q���� u]%�ܣ܌��ԭ���)�_�;�:�DÚ�tT�.ԔV>xh^�8�s������%�xZ�m���y��1������^�����K���ܢOv�[���=P��+��#F�ç�p�uj�hϱ>v���*��r��O��gO1��[;
3��0x
a#:c4;�&�:�C��N��:�	��c8���e�'ҙ$�ٚ̮K;m��#�R�����A��N�?p>,xj��9b��k)��Z��I����~�=6��e�-^;[�ܛW[n�%f����Wʾ��[�ۘ�$����:����S* :K�$DeL�WXpL���ә��R�o��w����'�������KIEF��}�S��Z����|�f�KGG���A��{�&��f�� ���;�@UDo/eem���Dҡ���U�t5��{=��cu��6��O9iBG���B�Ao��̟�I�d�r�;g�O������h�LN\\�g��d��	 ���;�5D�����]���]FeTY9�m+�j		NX�9�i���V���
S޹�5�w2�y��Z]���;�0	�c���}dHm�Q�̘G�%r��p������N���Bo@�T�i�Y7����/�^P��KY���J�ן!:c�4�|���l9���|1��5�#�8뚂��z���I�������6�E0��Nd����)�S�.�}Q��+��E��_dJ���k��Y ��v�!wO�/���9"����
>����$����d$>#����mr�=��k��'M��W�	R��
���b�N�2�=��w[.�h~���+��O&�1G�_���x�Ň�H/Ov��9.k�6�L�U�X������J"���ǭ����x�8��We�ʕP�dw�sN�Zȥ:�6�1$q����<d�z�'|�ϳ�Q�^�ǀ{ax��8W$ݍ���ϻqS|_%�q]��MD���
�c3��=pmO\�	`�	�s ��ʼϮ��l��J{s�u�M��v>�kǨ�Y�v-rMj��ѥ���:6,�����'�!bW
,!É�V{^�`K<�	�B��e"�2A;���]���	
B�#H�������ń�~�^�ɚ( A�����;}1������͹��x��]�*+Բ�,`*	Y�RB:��>��6Y�<%Eɏk�K��W�؋����n=��>|�,��p��I����C���#ֹ�#v*�H�=�[U�Ȇ"SIc�٪�������(���a�}�fY�l��Z*�z2Xi§6������q��K��z����ժ0l/e�Fp�º���񅨎�j���X�@U��w1��i�myx�Ah>Kۡ.�|@�ť�74:H���noo�������	��\��=M��a���tx�Z�(�Ѿl�o)�X�������Jk�O2��;[�lS���)�jy2���l���,Қ.��Li�62����؛�|_�⬯+S�&�Xz5�Ź-�;��}~�S&�F�ӮF�|0���3j��:�S����C�^7�8�a_�fhCl���� ��%.r��X��m7=�`ZI�֬f�C4���t���mƪ���%y����^_���V�i S���9k%2��)/6-��'[7�Ϻ{"���ɶ�o`�X�\���6T3&!u��+O��>9��%7H��XBF���a�jd[���U5F|�  ��.�
�:G��':�@`k����^q!�Ҿ��_ş��X�y������z��xs �
kg(�����ݴ�c����l1!Cs���v|��^�`e�� ,\wţ�����8fT��ߝ������#g��/�p�����;f2�P9�Æ�tSDC�9�d.��?#��Ȩ*j�O[˖��^Y�b�-R�8pv���)�"�s�� �-�
9h��)0�"�n�7�.�RL�0Ş���6���BP�?7�/E��	y��k��+��dmF�Y�U^������2�R�� B'��j�>�U�e�VR��O�Eg�FM��5�'gwums��9*�q0�|���<"К�G��-3l%�`8�>�Gg���"���3V|<ɐb�H��_�~��r� �j�͋v̩�6��Ԍ�f8)�c�p�x�;#څ�����Y_���m�e�:��ݭ���ر����X�K��M��Yax�N#�ć�i��	�VuB�n��h�������"�X������#��F�^=���M
�5L|hE<`��y$�#�,@����#���c#~�2Pn&gx B��բA�OM�3�Y�Zbv>?#H!�,Ԣ+�2��Cc0&�Ĥ��vkˀ���{[�(u���q�E�.���	^�꯴�D�H!�����ڠ�V�=ϵq&7 �,o����E�6����Hŝ��,b��o<r~O��#��.u�@���.��n��G)V��\��������4�,xcd�45c �[S�KM�?Ǖd�o�K�H6��S4��Q �:Vqp�����N5�;��WPS&!��]D�����M���e#�����\ى���=� �7��Q(G�nV�[}���Ma�4�#7ᝥ�>�4.a=�s�:K��~t(��7͉����܍+�c��"�"�!n��M�)	�GQ��w���:j3���7�!�wY\u��ɦ~��&� ���8�h ���&jL�k��3,�=TȐJw8�����-)����)����� w�B
ř� ��	W��kFQ˺���r�DIp�������p�&�w٪�ʅ>AȚ�'&�e\��������ͯq�����B��x�FH	S�<�L�y̘]�L����,Ȧk�Ԟ0�����K������+�-a���D�E��zA��iE��|6�� �{��F�Ą>8�~%>��~��(Kn.-��}�k7�������ap��讕�N��d���[�����;��/�+��c��k�i��S�5d�l�_�6	���4Q}Q>Q[1� ��=��w���Yl���y¥�c\��8�p�!�Ó��{i>C��OFɔ��Q�ǟ������MW�>�s��!��y��Zk�P$��JO�\!�[�q���[�g%��R�MT��K\NlⓟΒ��[����G���-�W�s��1l����}�KTI�h�N���nᶙh���f���o:�࿐[8e;��P ���$iYH�fE������r���T�~o���/��-�X�m������6�1��9�|GH���Ҡo�p���Q�ٱC�u
G>}�>���Un�箈���j��a�����6�Ν���� �r�yȰ�y��.��c��ϽS�=Z{w�Q�?���@+�^Z�;l��)_D�.M�W "&yy��ݨ/��1�ˤ�Vm$�+ �ݚ(�(�bʪ��h7���:�mP�;#��Fs�b=�Kk�"'��$(���<�_�L�W)r��b�%���@a����씮m�!~X���R���4b٫	}i�*{ņ̛��C�a}HbC��l_dh�e�D>O{��"6/
1Z�0R~[�n�q9YL�ڨ,d�K=	{ZV��M�s.�-5+�b"�����[u����N֕����;v��B��_(U �!Dӵ�A��\�~Oa��G𷰳XGWϚ��K���17�B_k�`��������ж/�u_�1S�-Z�{��Cg��-��Rh��xn�j��;�}�f�t<�8Da���7��,Ql��#i�[�h�Qn��K�|�� ͹�ǵ>�-�#-Xw�@� �d`�P�uۺ�n��r�L:Ե��h�~���z��d�Ő���pjhm���G�A˯��,���Ǆ}��Qr��T����rUM��J��jF
桃�G���y�������rjH�����G��A�~���1�B�.���qwt�h����͆�5~�$LQ��-�.�^���&�{[P�zJa��)�����옕_�O�0Hh{j���F|i1U3�ou�{�b���r����7L�]�$�R(�(I���&�-O#�T�f�e��k�#�����$|8�h+�M�;���Ht�����+��+h��0e��I�I�Y�q����K̓N���B�^ض奼�;�@T�gӈ�Е(�$ ֱ���#S�ˡ�ew���.|�����z�N�"�d�p��������H�����4;fo�U��߱SF��Ƿ��b�;ߤ��)E%5��jtV���y�?�,/Q�R��8#D/�h�7��(���NY�|�ord�u��Qk��`@�F�Ӧ��8\�;��O�t��Mm�@�f��v���x�ŕ�z�'����9�3Q�M7� �3���@�W>K����?���n�o����di�jP��Yxc�����$U��U{UUn��ha�I���{�m���? z얠�t�r: �昧3w��݌�f�o��l���Y�ltDq8#���cpT�/%h���B`����\�&��f?�=�*��뜴W�tB�N��F��^��_�\ô=kԫA^M_�ňԵ(�l��n�����a����&t*II���;G��6%�;$�[�����jAW<���,��ĉ�ZI�$���?Q5x���#�� �?*I������ͨ$-NˡR�|s�h��(�B���8��s	ճ��,�\%��|RN���:ٳ���O��!f�e���JhE(@?�>�Sw_�-�0���?�aQ��\�wY܃4�b��j�Rx��Х�F���o>�EDc҇u%lЋCp(����zW�I����O��(Y�� �V���&D��:���y�GĻ�i�Y�Y���s�+B���
��C>�tz�a�{p�����#r,~X����3�̉�ڨY��`� pP�a[�J���Q˛�mvݭ��b4���*L�N�sr��U�n({kk�%lK��6և���_�{�L�a�h�s���R��i=j��lrQ��臏�r���H�X��?�Ю��m*� c�˳7-o�\�5����2�0X�����n�2kǷ���LC�#�D8nu�o�=1x?�pP�G)z�~��2�\Ge�/'a��R����A"��(^ukޯ@r}�ɻ���r�s]�3��8�`��_c� aC��P݁�̵�##2��ge��x�p����F�â�w��.ONd5�RW��V:H[sa@*���W�yw�t(>n.�.��O$k�3�Z}����	jCR��1-`Ae�6וǫ�1�>�r�t�Z��O�<���g���+�<]|�p��5h-�-��}x�.!�������O���,W�cp�[Ō�/�O��)��gp���ۋ��i�g�>6k��e�Kh�LҴ��O�aSA2��#�˯n{���3��9z�oT�m?��l��H�X=5��֊X��7�ܻ�ض�t#��/�4�|*��o7� ��%�!��j�OZ8c#�%Yi�^-��&�'����l�&<�4d6ً�05	6��?���)����uF����`��������T<w�*�����B me�T�K�֦������Ti���:��f��ׁ�Lۓ����.���=&��E�xv&��[�I�p\6�©mu3�5����/"U��w��a4*I�<��ǟ��˱4��}N���6����fBV�o�%���[,ϋ=�h$Ds�\F�Q�%���#��Ӯ�����}���ѾmGBi�����e���j�����`�J���_��RJ�Ǵ� A�'�[���� �m�(��r��ܜ��C!�ƍ�U�eXs~jp����L4	2��V����H�g�Ga^��E���~����Lc�]�v:�C�����N��.�٣D�'/x�����ٓ^�IǢԕ�E� ��	���b/Y?3q�Nf<'y�g��k'������d���sϼ�^w0�ӛ<+sBX�So��u|*��h������jI�R��QC�� �Yw��]PWox����BLo�y{D�;g�:��1�6���% J۴Ь�����1ԬHA�;�o~��V������[��6'�����I�ѧ�n��<��p�Œ%�2;2H�$�4�KG	s�$:����"&�ve���Z����00b�B���2Z�Ƣ7���K+M���˹(J5V�`6��ͷ���d8�y�OL�>�YT����\����[@I9��?����d�x[�:.��[v��\���GR?���h#c1*���~� yd�ɕ��C�0��K��ڂ����_('F�h	����n��c�?��LMs��*���ƃ��~H���{M�n��|�Ԟ�)����l�TK�҆����u��d ��F�����-�XZz��Q݀x;-�4�֋ڊ�	�Q*j�M*�aN��c5����D�А�@��M_�Zb4B>F��:�����@{���)1�5| ���Y��$ �`�d���J� N�7PE|��9��g7}�F)7��x7�7��w�?*g��F��X[w�7R��Ä�����JB7���@��Z��lj2��(� 1��y";U ��������/bB̿�T�r��M!5��J�K�����������p7�N��l:������ӱ[ǘ�gY߂��	8�a�s��Q�A�D3�`���cک�WiY&��@*�^���<�(m[�I�� <q�`�J@/��u���� ��.����f��.Om/RU�&��Qvf���R���tR+�Uݾ���i�BT���
�)uQK�ӰPSK�[��y��q���c�)�(Y��p�iP��-P�"�v��U~B���n���fq>h9x�[�"�{���a��]�xV8x353���}�A���;����W�1"
�5��DP& �	�	
Q�H�cU%{(�+M�nw��3���A7���ܶ?��|pX�=#�s��&x6 _43�RPd��ZVs!��Eģ��g��|��%	yl��A����,Q��ehe�6���Ѫ�w��sZ6m��(
æ#oc���čL�%?t��J�ˇZ>en�iN7�����N7X)������=O@@,��"%3��9�T@&a��I�Z�������y"`i��+Ӗ7m�Y�<qh�zz�Z辇����F��[M8h�:�r�E���aZy��s���l^�7�m����Ŭ�����@��^��ڶ \�l����B.�oN�MPMc��k�#�����oi�.�y���O59r�(u��|�C�;n��`����X�B8k.c����؜��p{�T0Hc��eƱ���yE�³�Z0e�M��Աv>>�`<�<���]����q�jO�,��"_�V�����n��������)�1�������b�)��c7�Gml�7���f�,p�I�w��~��A�Ƨ3�h޲��m�Z����w�!�>�-r��2X|�(<����g���6S��dlb\��
�p^�I��K'*[�ϝ+��O�|�I��;m37��S��)X��o�W;�̸�s�/k)SJ�T_��}k��H�mk�;��D�=�ӕ��l>z�x�~{Ecpن*}���, ��;�z��&���,��/�����HbJ8ź#'�!�Y����͗�}���;Le�1R��UO*0iq��:g�A1�����:_�"�bi��jwF��a�y���yt���v��}:�<�c�jIJ����%
�{��xVgV�*��d�ks,�(����KSk�h�"J��s>1�x�)�ױ)�inK����Q�wR.�$���\DXQ+���^*fQ0�\Oq�q/H�g�H�6���8|?�o�i���J�7�|�9Q�F(������f�Mc(Bx����"��G3�I�5�5t��8r�lB�q���KQ�p|�
�\�:�3�HfF��Vi�&���צy�t����M4� �����.Q&�ʧ��4��)}��XX����s��B�r��*�]z��-�f���(�j� ��b�b�-nB��_�d�����8(�7�혆]����i�f:��ۢ@%���Q�l��X2��/i2�D^�#��
�||�s�|`]�冹�h��痁��^G����@5��רU\~-��G,�rsմ�S���,�yH<ۧ�5���$|�-�QWu i@6S$�9�3ѻ�!��3�b�(Gd�O�M���0¿�Cý�r����w���t�&�ޖ����/��Ŧ�2�؁~&9V�,���F<�I��/.�R��WD���+R���g�Ig�,��QϤ��Y�H�K��7�35z�M�Ϟ'���u5�Mb�E�P����i�5�7�	�64�޲�������Rr7ϩF�,�|Ֆ��8,K�!#i�w+��!t��A����YT���B�q�a�&b��N���:ؚ�541�s�D�I�µ�+��	\
���!�r�Z�AX�R�#��H�r����]��*Y��z�L��'`4ȴ�e�DYQ݉�T9��KJ�?�/>���z\K��=C���<;f��Ʌ{c���)��u7�j�հpئ�Y�Of���Ee�e
俫�&mA��
�����s���%[�x��$�ԝ�v����'%2���v�>I\�h�i&�g#h�C؃F�HM�ԁ}�5�hrܖ�j�ސ�2o���|<Qn�hn��TZ��c���p�w�$)�p#����x��1-�teN^�ߍ��&�\9Ӄ��痲72:��*9��-�.�eL���#z_�4I=�>��@Op��tpA�YV�$m���v��b��ߌ�1w�������疋؋E0+R�^���
"���g��Ҷ�\��|��t��^EHQ֡��V�־�V�����Ā
"!Ko	�͑����Y�5Y�ʹg"�������.�!�Zȗ�ϣ�6�p���tM9�{p�+K�2����W���"_rK%�&]�ƣ���{	�7��Ӏғ��)Uےd����GA����xȼ��1�.�P�g5H���N$8� >kx�bIqts�fv��ܯ"N#���-D�ý)W��(���#{�P�G�|�!�v%���g0p�o��*e+�Ztu��g����f��Y���!����j`��ϥJT�h�[ː��r!��*�[z\M�sl 1,Ó�p�U'A���o�u��S�u������F/Ei/%W�d���2w��K~�V�Q[>����/�ήµ:��z,Gȥ�{����S�+Qeɥ�tL�w�
��b+��8UnqV�&��s�э)1|:N9N9T���ɛ�~��JU����H����t���8kPdu�*d"�`���*+oW~N�k��<�.'k�q��*)�3������P�N�G�Ԋ66���0�,?B��^d��_�s˞�S���n����w#c�#��7w�G��X�/�v�$����ծuXU�D��ǚz����#A%�h�B�l����Ξ�yۅl�*J��M��"��$C�S�s�rB̤�o,��7y���N	��"�7l�"%�<(!��`�H�g�*�;�IR�*N�R��� ,C��w�iG	l��'vJ ��h!��5`���x,S�3�z�s�zO%��	/��r����N���#����k�W|�+�vD%��ި��b'%���~����^uo�����^�<w0�L�FW��uqX�����a�I(5ם��;ڼ���ky���GN�����6.����$�<���kݢk��
�[N!��+����$���x�΢�D ���"Gϛ���+���w��yӯD"91e?ƘK7�>g�d_�m����c���.
m�U'�����ZJ�T�&�Mű�8��J0�9T���;�Hȓ��H�4L�>s~���k�y`ь'	WM}Z˪��ht鈳��0}�t�4�HE�ģ�]<�$����T�Sv���4�q�%�@�������\~>��T��J�W(����Y�z1Z-�W��g�^�C�E��AEy��WIF+�Q�TE,p��TMgm�,F�._֑��:������d`@�\��_1��C�G��1Q��?�L(mK�G^
!N�}��b���񩍱e��!`h_���F}��m9���ǯ[�'7��w~'nқ���ɴ1M��L��p�Ki	G��&��?b���bZ�<��čҶ��q�IcH����P	��5�U�=Agosi/�����u�������,t7(��Z�2K�&��	/}ݠ���N�AL�Q��1��;qїҸ;�-Ղ�.��M�EQ��[LJ䷖L	́�ES�Btާ�S2�Iш�	.ye�Sz�Sh]6����(�e��Hۍ>J�$�]0[3���b�Ҋ��}�q�fѱ��K&��+��B(a����!����\P�(��-��}�T��_Y�1#���3�b9N�ԏ�HsU�.�T�@1��KV{v�����w���&�����*2�k�Ͼɖ:zN��-8XY�#?1�"!� ����h�K��b�u����_��fЩ�8��J��U�/��T~��=|J{��9;�������Q�b���&�-o
��i�6�f�)�����O�*�u!Դ��s%��oxG����q��з ��c�������}�3x�S���C����j����~�W����W���x���<%��H���M�P�C�/ص\�G݇~,A��Yzf��HV=�5�����x�F��U�Z����#b;ݧ���)��bd��;�/�Ģ&��Y_A��:l{�y`HA�z��Q@�@��ֈ�q8.�~�o�0�~�u��_���?V�O.8�C=��׼a۴N �����㈄� FD�jRuht�3�b?P�����d�DG(�j8�-�ɶ�NYyg���7������>�}�D41~ [�W\�"#���V���hF�L�pb 0�Ȉc^&���KWh���z(��.�)zq$m�Do�q��sX`���l���ù�V��W�hA���*)KС��nė�9�kP��bΚ�J�1Xޢ�Y���D1T��k�/�u?�iU���n��)^J��s�����y�x~���0!Or���"�ڄ�d:g�	��s�7Y���=���+4�|"��w/�U�
j	�A|]���n���8Xv��޿�=)�u�O����>�^�[8GS:'a���e��^Mɦ�g:�2�I��$h�:�H0�`N�0y�ȣ �����c�Z�IQ
����[!s�ȁ��t��x L�����=��ܹx
b�-�x�U3�^:��}y�*Y�� �Y�Od�C��'мsv�'�i���Ғm��x�p>d�6q뒋���ʕ`2R���8�:�Wt���z=��N�����"�fo��F_��$nbv��߉XURY�N��-�K�K��	������$L�7�6:YD^�5�.ϖ��K߳�f�y�E��P[�)�[Q9)$�L���C��P���-�϶�s{�T��0��1$�W0w��>�븺���\JK�<��4����Y��,�Ǝ�зr�i|}Ϻ�7p��ѵ�|	[cֶ��S���
<d>S�#4i2??��;R��r�6��?��mO\������y���|���`\!����C��Q�w�J����Y(���B�QOj��;�n����ن�pQe��Ac%صm�>�2-�󊛐��D�@[�h.��O�O�-@W֪m��B+T_ʠ�I	g8�he���7i�R�WU |�ǻ��d����).	Ȋ��:�X�0���ɉKZ�<ʗ�YKE�e�Nbv�P�d4=��f[Q���>7�"}���j8���%)9�����fʕp(�\6]r�J�s���o�*!u�ƍ[�Jj����n�A���Cf��)��+��a1��9�˻=g͂F�Qr���1��a��	 y��Ρ�!jvݵ|.�����3�}�>>��:�T]޼=��ØN`����}�SN3��4�"��t½8dʃ~�8kPߣ�kp]�8M�̄��x�_X�Y��M��܉�"��̎M/�֛=:^���JS^,Ӹ,j��_9h[iС��w���X��@�N+�(�	À�9-��͖TY	�@V+^�W\7�9��FL"oC�H�����W�\9�wm7m��cx�-H:6���h���sJr�SY[����'Sq�E��=�c"1"��Y���nA���9<w�9�8�&9�|ߢ�z1�2c��Ꞝ���9�w�х������2:i��+�G8Yq\�&�b��
�Y7���e����7'�s�֠����z�����`r��Ѥ���D������	�^e�fh���5���w)-���V�V�BlHsles���,V_]e���L5�Y�/��R��� 6��W��ʤqzB���)��s�F�ߐ͋�g�`4� �cSp����ܿD���hI�n"�7��ƻVe��o�C��rз�*>Q��e�� ���} �=?�s}�N�֬��|I��b������6���5�q�! �.����v#j��XC%�WPv���a���^���9�	5םݛr��u�"��cӪ��[Oe�/���\��a
�T>�l�ɬ(���_������1��Q <�*wsy�%x�j�й/ο���
��];� �1@���Yl�Eh%<l`�^Q' ߉Y+�(ǀP��f�U�{�������ua�O��CF6�/�����b�S|��� �s�ƞ�a�]yA�g�*?n��;-�ܑ�10K���Q�t;��n��[�i5�����7�{&fuȴ�2?,�l�&8�U5����I�I��N�]V�O�\25Cvg��00���yg�� F�-����⭷�[l9�Ql�=��_��N8��Mߊ�m��:�ԆfVh���
�]���ƣJ\
F�O�!�|����8	�2���=���Y0�����m��7ey�=r��D�#$?��d�i���>�_����b��,��C00r~�#����{�?KH��$����G	+���Ϙ�W��譧-��~7��ۢR���	����/�~E^���s&�W��R��F&��EBi�� ?}�𣟯��n�?���m�.�A�*I�YSi;]������j.Yo'[��$���5�#������4���z�
���(3��Aw�?���J��c�>:z�&`��he�)�n�?��3��3�����Npo~�����"��E��B�!�Y�aF�AQ�T��$�Ҧ�k�Os@�쐉X@\_ek���l*IVD���I�jWE7�畳\w}���T�񉄽I(o��"��l_�%���Kײ�?'u�=����KF�Md6�U�����!:���-ӗ83;���N�	A�Mw_�kd�N�0��ÿ�b';&��i��@�o�{8|�-G����*�q뇤:�!,à)�Do����bDt����M��ⅴZ�WH	'
�lN��?HꕜD� ٪�I=�ZR�-�[V���ĥO�Y�q��A���u���!)�A���@(Wr�F�}���櫬[��B��~�%5��j-���ב.)7wz��v�o�q�A���.���,F0�+=���,D!�Խ���N�5`v$����@�/�K�k�����:�����|��Q ?�j2��Hx&$ד�_2��c._��Wy0kH�F��� \˖T�/&`�2Bj:Bݭ��1�0�^X}a���!l7����rԲ+ʤ�7v�GI�B��=�� �$�
t�%*���=�<���:�\�d�*�uΘ� ���ŧ���-�Z<��դTH�9 k��Գ<I�k���.���Ԡ4C'�.]���d�z��N�X����ހ���>�(z'۶�hi��ZMۺ�^ʍmUX&�(LFB6���-*�F9?���ۙV����X�@5����x��:M��{A}���½k[��)a�"~����)�ß �/A�L���s(��;�˓v����|]_�6X�@��$I,.- ��r�+9.NCx�I5��ϱ"]���8��)��S�ɟ��a�����98E/D�6�ج��]�e�u,�(�xQ,>@��ᬺD��䠬�m,�ew���U����v��Α}z[g
�7�F���~
�7�=$9A̕Z�L�^Y0�@!����PN�`
D������EN��!p�%&J��öU���u��ܑ�[D}P��� ��G����:��_�}#h�ՠ�?"B��F�M�d�@e!�J�ރ=�A��=\�����b%Ubɏ%�		���_8�oq�+���x$�;O���:�a���Y8��� 9��//��Z� �Nb����z}A�q����9�x|y�⿦��t6��4XÞ+�:�w�$Ǹ�v��X�B.�G�|c�0��p[�[�7%~|���i�k�v��K�eV�Q�͜�̍��(h�!��&\|^-�v��X}f��9�J�����(uF&�@4��x��)#�H~���۝����k��3�A�Z�f�ޓ�b�zї����@�X>���/���<ai��lN�<����R���>��N�<�����R���5C�'���Ը�t�.���k�{�<E�Ɍ1lW�7�;<�d
��K�RO�,�Q=�7O)P������L/%澊6[��s�|�_O�����2X:�v�nvsX�ɚş�h.���|��Ȫ(����^}ۄ�
�ގ,!hT�jɴ�����M� 6}�Se{�&���w:Hfm�Zp�/�g��Pa+1=`_�����J��h-��Oqe@|�.�����#]�)k2y�Fl_�6m
��*���(E�M:2�xt�tvL��6D`�2^�����g��e����8<kh� @r_v�L{
���\�#���2R�|f����?D�M2��H��"Lሌ���������u�j�묭Ԋq�e�0�0�9�N��Kw#���?/�X*�*U�#ׅ�1�f��ƃ㷲f�R=8��*�:T<̷Ly����Ңpzl��5���c��OOiN�L����nx��W��WZ�Uu�8e�ʮ�lk�5�8E��b��p㢯,�SR��Y�I{|Y��B݈�"�����w�f5�׿����=�q8�[wpN�V-k���/�/��}#B��As�ؔ����D~�ۃV�t)�MB�УL�B=�ON��f��j�7����q^r�	!v�Z�Uк��[��e
����>_S���������p"Bծ�!aX�� ��G�n!���kU���+�/[UVU52�#��fH�v�F��'����tP� �Fkk��$A8֯�yd`c�׿�Y ������8�0D
ӌ��7d�s���s�(��+4�&ba��9Mz��'q�IS�^�Q��3����~�۸�d��8�N%q�l,�MJ��S0Ҝ�h��<���}��ȭm<nR�����i-gn!���D\*N�<�݁�eKj�?.a}qfsɳ ��읆l�7� Z�(�s���K�?����5�r�Ҵ�|<�H5V>Ũ�(�8��|W `�[G��Z��)Z���2C�A��Q����xF�z�7�ڝG}��6��)f:,����n�@�,��Oo �d\����	oЧ ��uY����T[*h�cM*�`�OG'}����B꽎�صf{����+�})�h^��`�i�שבٲQ���g&F��?�$[�ׅ���FJ�/eY�;�jd�=ɡ���]UBT0��X�;7�]V4c�MK�#2��. 6B_E�����n�Fr�(�L c�����`)̈́�}�{|�|�<Sj�����c:8����9���m^��#�
��*mH��F=���L�ь���f����O�a1�qP#�ͰA����#����S!fhS������u�����ﴳbb6Ļ�AOX�U!�Q,aH<E�损]ͼ-m�SW��Q�H?gTH��W�\��1������%VԻ��h��m�`��a����rn]��S�u(97E.G �:��RP)	;��v�`0�bHY���(�s0�z�4]N6��6s	ɩ��o��6��hS���<�����Ék����."�r7��d���EFb�n�Q�lIn��{�Q,��a ��B�%[�0F��驌����I�U���XZw�����lbl�C�3J���=�g^A����_`B�u�;�D���z�pHvzR���>�~�s:����｛�8��:��m��s�����Ɉ-,���r��~��Z������i9LA��?���K^�h��GT.��m���RI��7��	��p{6)40�S����1�>�Y��vQ���e�� U
ŋ�1%�2!���ue���y���:I��t��G�X
7)M��a�3�@�~�5� �qV���:���f�#>�)�=��A�&���-L��:[���!v�^��-P��(>:�֢Qq(�-1�=�[g?�,���1�@��t���m�|�4����Đuv��z4��^T�~Rt_O����Ц��?�ᩒ���T�c������<έ��>6�6�)��?�#�Ӓb��2�p�#�֌�L��aO����m���d�(w�0?��(�5��c&��= �5�p)dI�h,۰��9Tн�Ȑ]+:e�=�:/A�6����v�8OJ�A�4�maj�����ˆ�I�g8��2��a���H��w	��?$^�v��*lb�?)e�n�>��F
D��i�+IE*pq���,|��6 kB<z�rE�م�ض�Z��h�h�1�k�
����ɁtF�أ�̂C-���p�g�K!k��}.�< �{Z�"�h#ny�n:��6��h8�HInt$bʚg:��r;�.�*���a`��l�'�0��lO�Y6��pn�\�M�zd�8G̽zI�<~��	�Dk� #��֒�H$�'�����G�0=��`���G�f"3�x��uy��R�j� ������۠)�t�������d'����\�� ���e�|a4�.�� �pˎq�� ߶��RϢ$|jR�ТG��?@��Q��MB���^!b"�d�S#BG0�9<�֞c��x�*���H����O �Z�k��*��c�mt��MS����PS�4*�H��a8G�;�=<�����^��V�,-l[�����,AJ�j� }fP��
��f`�j"
KF�D�l��I�7���{��}|�ʝ�3�K�O�b+j��g�M����P����F)�y�e:���	�;?�~����0��o\?o��Qt/6���ܞUا�yJ��+J����ܹL�Vs���wF���I%�Qf|�-��`<�9ʴYR"{�6N��	� �Ո��}E7����3M!����-;�<��I��KU��i�rֺ���6�j�J�!�<jO��H�<sZ}�zv�/��F3$#%�������"l�
�S�wx�n"�P�S����h!,� �Ҷ֏�z�S7B�,�q�od������^�5}�l�cZۋ���J_�.ކ���p�^b�%�%D��%��.�Cc	���Fcx�P9.��ulO��{7�V����|��>7�Y�_���kDH�k�U�l�˓�~W@�τWܭ�{^Ձ�3�˘��&
^����<���Aa<.9���ˈ�q���$���%)z�i�L�6� Bˆa��g��&T@�톿�]��霜��6�5��W�q6�,�i�\ğx�<C��ߝo�(8�k��oNJ�ik�?0���2T�>��dĿ����:�=�X�#����M�g��`U�W(.{���O(�5zy�Ǻ3e�*x��I����_��d:S� ł.���f�w~����WL�w+>Jg͑ž��X?�C��҂u<�a�S�P�����KT����XZ�C,u�`1��r?t�&Jᴅ��C+�K��7�Ct���蟄��V@l\�1]��j\\o?�	�@��4�|��ȧBJ^s��k�<�R��ҷGfr��(�dMD�d�e�bA^��~��$�Ĥ����||A���首ܜ��^���h�Z�=���!��W���"� ^{T�<�J!�I�Jg0Ԑ�����r+���C��]�o���������P����;��7p\��S�QUA�ً��.�B=��朢b��+��T���Q��K�ﲝV�LX�m��-�9fy~+��1J�˺6q���
��.���#E	t���~t�.:�E5^�8�wQ��BV��r������Ek���*{�bfB֑��bD�B�4��nO���Q|*��?�&��J_�X����ri2�1�Q�t��?CVDϽ4Ã�!k����&7�( ���6F�ܡ��?����QV{_<s����A2�Dt�nv*,u51��*:@���s `:��O�c	�
�3��Y�8�}DB�eUF���UG���k�ܷږ�g�6�nP�ǹÝ����^]d��B�e�p�Q�EM���;��]kI�h�Ə�3g���歷�����8^������9��Yd#�59�)GUΆq_�@��%]��[s���f2��{���LFQy.�
.�|��r�����܆�k�=�rs�kSB�����S#g�c��H[���O�c.noj�ANS�����@�Y�-�?�1�p5�|�t�\~�e��I��\�`fڶ�-�Ù����D��P��o"���x��A|� �o2HS74�Ȁ��4]� V,���;W�������tɔY�XT~�;�7�D[�S-���6!�0N�GzH�z�"i�{j?�~�SH��`�:�w˳ծI����ۜCps��j�â��KJ[(ڔp��oX���{�^������\�ꎆ�H�b`�F���6��I�4�b������;��ys�z�'(ѵ6��t�LU́�a�Ye�dY��+�$-�r*ޯ���-��d#�$�v��V�~�^�l،�җN��>3)F��>~5TH%���%AQ'��\\+���BDϱB�tz��c'�G�yY�Vd�:���c�X+Ic[j�q��H�x�F���>��oQ�uє�r�rafGp��٨@H�C��Vo���y��R�y����\�0ĭRSy�;�[�g<���KF��6�-qk�> ����
��tʗ2��G���_u�W�����@�	y�e���l������,�'5���
F']c�#|��Y+�Y E��<�=������d�]��ꕚ:��I�|�:��j�?+�m�UD��A��W�]	�!�07��azŘw<������汢D`D���v�L-�.���3�8!�	�{��k���sZ����7&�w��5���k� �&b'ѯ'�3e��C(���h�Z6YIX�lׂ�_W�4nuքB���!��pQ��:��0[nIyƱ]�>�]��?�3��*@S���"p����m�h���g��I�݄�H�J�׋4�[_�l򕦏8���LYy��ѳ�v�����vA�YV��X�n�,	1bS]6U
�i�m�J4A������@fJ+Z�"�bm��3�*(A�+q����%
� ��}����=Is�6�9���r��k rt����E�].��˚�w�n[T r�g��Zn��#z�uS[ӊ�y�vj��Ч`�#A/o�k��ʐ'��?�s�"*#[
��nY:�����4p4`�[%_�W����O��� ��t	>(�<���"��)k�����YLʂ|V_�=�����>~��/ڷ^�A��-���9;�����pGߩ�kS�5����c�]OeT$�i���c�b�rR��"J`˶o�c+c���.���1c�C���7�?�0��U������>�0? ;�w����N��s�K�s$���B�T��#{��B�0� ����,�ﬥ��c��2��i[���"�� ��A{�-�����Ҡ�U>�J�۽����ve=6!W �O����ȐB9�m�	����+/C�;�Vi`ɇ���n�RF�y�lYR'9p`+A�h�Bg�	�������z�C>�˙���R`��H�s�V��[$��Z����W�E8 <�� )J�:�`�`w�i|B�j<��{�6����7o�Mi���[#���<�P��m6H㌽� ��)#d�e�Z�i�����}ǯ��H��Ӻ���5��=(����n�#~�=�����!q��|�)��짂;T��+$, we!���٬�Q���A������~���)20��6P�#��N�[*�,b�N,�ة���R)|�[�~fl�;(Ă�`�XuI�(��9��d=��
�b]�YbP�������s�-$��N����TY���Є��4�(�� �f�u��Q��䩸1� �o��Ԝ��N�,$@��h�C�{���@�u58�j*�VF60pCK�"߅����	��ς���˜Y��:,!���(%T#p������R��]Fc���	��ؘ �c\����kH^�΁�
D±��
Rb��'^���/-������W��+׭������&�`��y���}+�7�����&������^O�kfd��9Ne�4i )�|���q���w.ar%�Qr)mt�գ�
��q���"�������y{/��,CX��Ys&�� #Ԥ]3gSv�R8�Q����d�^���OD��I��2��c�m����}�f�M�C��V��ia��]j�� �'���*�"�9n�C
J2���_Z����R^#:�	Қ�����o@ǿ�\�Z�wM�ˌn��ey��=oe`����Ob�8�~����W�Xp�����@�#i ����ߵ��^ڌd���>.
C��n�I��2+���fQ�bի~g8�ND �`ܗ�vlݫ��r?�=������Ѭ^��V�u�^A{���e��g�#��{���z� ���E�5���� r^�߶�d�(����љ%�YX��Q)=�aK��^�v�5¨>�(��qL�#pY3�&j����?̽J���#N� J���Y0^��>y.�+��='�ͫcs{�&)#��J��_����W#�S���X�"ߜBs�'�2��U��s�_�RQ�����R)ϝ�Մ��޿���S����m�RDNK8W�~*d���hd�V��F/�
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
byuLOm1S73HwUQhSZQ9A9+z/8fFlpdRpAIIrK+0xyzQTTwryO4mWCRXviDzKidFHJ5SOeCHW+d7a
RCIlvjIFfDTB0nUKK5QFLTBv++mLIkbW+FxUdk+MA1kbPAuABWY+ViHNNc1v38cEeizTajNAXksZ
GyORw8k11JA2LzY5yoGDzl4Z0rW4g/YEKm6+jAn+s3BEoMOUvkSRGBAhlqUVqCNpVfbQePqGZ2Xs
TJAY5PjDEK+WrN9KSOsUqj5x4dJo3ZCAqUMdodosy6Yaum1lTNMq1w6KYlPF8/oQcDWo55WWlXtX
uOWTOWSD/8J1oV7VzHbAqB8elkpWq2t3eMcbYQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9424)
`protect data_block
hsvqWUiwy51EKMvihElCRtOXW4ImccsVQkP61JxrzWmWj6GY4L+mvKI1qNKShaScohN0felXYxLR
mkNyUCwYWIYaqB2jitehNjE6zJ50eFVB9jPgXDP5qY1tZ3KJ1g4MjtAJPNwOnXonoeTR50dqH7Zo
XRC6sUf1Jzfmj9cwntQ5V5vgqEliAYV9DRFpstYGm2icFC1Ixtg9j+tb2RKGO5xDTKv45WJKXXuG
nJFUUYHOCRh4RvgoF53LwCasA3tIy+o48tjZQGASAfiz4mn8Xzjflm3PiAPWMLGN8gsPehvdtGtH
JwqRTiOgRKSgtb2BvbWIhsFC90SKJcWCgHusMZVI80hiRBbDwl1tZJ5gzFPa0ZaegdrfGUy8IIhv
JdFgBlJtGXApR3l1uiNOjc8rIx2GpBBanuF/bYsQnWRQEvOcq5mJXsQGp5JsAS6spzNLhCC1dffW
00qgoVVC98scT7eGlNAHxwFVob979UE4AVXHRbuIr0ID9fa1KzuR4yfb9qXLmUwnzhqMR9iiJ8It
4cowMzL2OqmeXWpclCkPA5lt1yakPlzQND2gQWOIwlzQ9hqdhwRgl51d5wyoGcKPwL1Ei5hXI0Rr
wnUKwsufg9njw3ch0DxZmWu3mNpA/dtZfigPlaMcsaSo88tmkfMp1DCptTm67zpGdFEULDxWgEKn
xw7/6LtFdE7zr7ofMNk6h7BX+EVoN/ZbHtFqsCynETE4IHNuqMyqfbCu+3fPGQVnXC46sI4ku10Y
nkn6uZadN5c98BTUY/JMclr3hPKJ9H6LF7AfiHLTsxYXHC9C7f+qTzpfZx+/q7gr70LjfTZ7GgQE
ZjBzPl+4rwsxxG7BTNBmUhHfRE9HAHijXBA3Wr/bEtLFKTIAnZvbaw6yB/xdInDi03utJMlNJ+XA
IB2ST5NZebnuhqxhSoWehGakcA0VrzXS8Mz4AE8cyVFhrpp44EvbSpW4aoQOtBSWYHjfYAHuBB1z
nOfpygLVQgx+tjtSDiFu/vI/4cuxLVCPB3Nchgqay+1wdAwuVTPipZKdMyIEaOmMjIGKyWOkHHjt
4e2BzX0TzHltdMTm4TngQD4N8ep78yaGBs/jDKpn+Oyp9L1QWBK6vsHhU1eMVTmJdpkevtBoT/8z
geuRw8vEth8smAZSGlfyMqGv0LavUPcgOuSmIF0V4WUeyHVJSkyXk0xVoM83lIJhesvXqCrqdo5q
/sM3nCv47znfA0DhYFElXVRTIIxjb8vP5YPL5FXry1lcYKYooh70IURb0tEYBXBDgEBG1YAWEgUj
ujG3/9F3n6qA+PZ7F55t8PvJJYAQwLJ9jDISGRLopVKt6WXc4lekM+kwQRHJg8hK9m8TkeRYpUHH
yfEAWNUUaDqwITGj6Ndvys7xtHkcYzbXIpeZnGcmzCI59PPkxC5SHsiK8AwtXXL2ctl9iPHorxMt
fDnFcaIPdzqp2RrWSDEkFRBQ+xZidi6Rv5elS+qgqW5FSs5bQxx04zWVATq3UFIzChWMu6N8/Svt
4i027J9dz8IDoV0wYxM+RCbMilwpS+6irun1lPKDbiD0kYJ8rrwc4FjD8kbhKQ5Zja0flOyV+3cj
lSFixfsbtDQWLT0K2/QHnRscYiNbTiBu/6u0n/Yedn4wvnJBo7HnuCFGSe+vL5jwBqqOVxnCp5aK
BAFqwoo2A+2zvnyjWR2ltA3EV5TPW3RkgqpTGqCrAhY1yBsHrOJc1mDKOtdGw7zLfmtx8ZCMViOx
7kovptzjqus3nSj0k/MO7CaJAwZcXrj7mhxSQb5YAvDDafR6LE1jgan5odioUDnvNFJsOv5R2n1l
Pua7zsfpjYapWn9k3dnfBsDvK4meSrlCrH8vvOs3fDwfBkF4m5wTXHzzhrA1dXCweUWjbUGVFC1u
zglIM8ck2oDKDw32uxLAIZcCvx7PV2umGxEEJGmaWADOwPKUunQFkmmJyMHraqo+5ZKHQtKYrdq7
HOmSMFSNUvNG+qSuMIaGEdVgx1KKvIkIi/HATjEtY4R3EL2llGmRVaUxUcuPllHc9TuPCeX0gx6e
YBfRN6BEAjpFBhhhRX3PLm4OPpzwkZYLizVuNdF/QPNRTZmMuAVUa3kSqj560Zf67PmJ3cME/WJ2
lek/CCsF+m5FnlRQNflMdM+d/r0o8FI4tnqEhhKbIP+Y1D30fU3t89kvPS3X3u1RSBpB1/xrcItm
qOToxEAkMaeuDekv7sBihWpAspoPNjg+hjkpo3oxgQi9gzxdacUWig0X27P7tSfuKnSzLfZbZNTa
eRRkwSf/XPdIdI22Hhf3LmvWeTRQHWYgWJ4eXMyWAsi1QGQuPVtGgI+iJal+09eRaoQO6JmMIMmY
+/VB9v94QcEh0AI7v2K+gIwV1cR9Hl7XzxsZ/X3QKpmP42We9Sb0iW8qEK7a0nTcO72f/XhibMip
RDjGaFsvxBc15EAPMmPv+ZpsO+SeU+TNrH4hA5acjclv5zhRiO7RYf6upXHMbiGwavcewJD8bwqt
ynvoLuhUo2mIG9pXTGVv1qzglvXxjEaPwFel/VpBWoheKpX3XoL8e5Ja2uGPszu+avDyTSdhPvKN
mVsCjRspDrQjh2JyrTCTU4ddyaeSlJR8F9sxhtBcPa8FtfdawE/VC40jeUmYTwrYJowea4PTfXfZ
Ueg7X1rQg+8JMyBOXa2kP256OiqeAz/Q3g7HflAfXLLq5FB0zQaNIoOwQ690UTubOc3QHx5xarMi
O2HBjoLTgUmByU9pm6ZwmexhZvR/E7v6W1uyILaD3JCMkJnBGzKQmF76ANrUVGFig1IwozIA/EH5
apR2pCsvisuHdpsct3igou4JSSUmTn+assOd7IfU3UTOt/o4tK46ZcCu8HkTbzlF3FQsu4+0PBzF
E/KpZJFGEgMZ5NBuVw8uPtwNPnEwGfejg3ypBkDSijXpC4lWx8/lWIIujz7zjzC06nl3ScAIO69R
3490X82rRC9ukFybOSJItniupRMV7KAJKG7eiWKzn4nvLbtCERQVGFa35u9eHI7f0bSTorHlFZT8
5YepLDt//rvGtqaU2AZ2OZBNGhKKAlxtZC4Bg4QPpxCwvpx1wQMWgFb3O1XQ7P/Rkd112ypARTNG
XX+jyI/m4lUQfQ0k3W4ObDKynOi3JSxz1ymz2HiZv9LFrXBOnFC+ZEJl+BpyjzIBq2y/qw+Z6kRF
Ags4L4oENO86Cfc2N7tU3piHmECyElY6FUFIhrl9znZKJLU/ev2UJ+3QtDIa4FdPL5rpPXRfsOHO
n9tfHKZxrRlemlCY2tI+pIi3grAWpkTPm1PRQ8RYh9MBPYdCyP+tqkKkmdQgQuVPDrHt4J6tcvK1
eb/cgSasBg+ZHf+Ml4MZ3b1TtQ4z13DLGXY+7cdgNVaOIo9WJjF8L930IDz+0wZJ8n3tbpvElAGS
5zbQLSU3w4/V/21OgSMNohP8D1NgRst3bEUBOQ1twyrF12EW0N5ocSmSQSL172q8PvAcid3ALCF/
Fga/XUQlZSvaSuajoCA5kwdjM48mhTZ44uBUGrJebNk0F6C0q3hUbkzb5eIqnDVpH+RWSgsPU1el
l0uG4Yj1rJnTVBCC624C3IqyP29+BzSbOOGmW/FOupR7rBOhYHgZODOz6MxISfso0RbVa2fomBWM
ZG0FoBSHMue7V1AIh0+NH5sM1NkPGepfooEnqjIZp8yqsxdVrX+VvWYgCdmMQM7rAqCoRT0j7BFM
c9fi9WL/P+fhnC2znjyie+eJMRnox6Rp1Qnf58Ec+jLQKgerefBCR1eibSMcr5MZ/imOa9tHEM0x
DsTli1GkOJFRQzu91FBcypkn7Jc4My9hz5JnE4EUCb8MbdFgxPPDXs0PXyzCV7LMfQHnKP443Fjw
hD5Ih9VAGI2RaPlVZKrm38u8JvFu3RygER2nMf5x2MyIR78cyCl1NAK5P0DYkX5kAL2PLnnkTumB
faUy1xrrgp8t47d/pbczHbfajk5GzGRz7T6/T4GV+K2G2zQ7CvYV+gvH9wep7WmoUpl48f/OJ/+g
rBvMClZRrIZxqM7S9wMYfPwN0bT9xszo66O3e4J8i9tyZsioNdjfz1hDAK3ZAZnNiiTuS637sEaX
nPwltB48kmtMNsyrTgZXBxh6VVKaqAKTw+CYpaGZALNwgxiaQ3XfiSiq/VHq1K55zezTArAe3CyT
h6kchTW7B05ntQ2uUkYrmJamGWXegiZjwegkjSMePyRdFfUI9EbQcAD4s3GXHN0+FBVeUd5n312z
+P3lVV8P/W8jBbRaFrnBiM79b1+Z1QB4geCuWINmSwSTtcUAZVDrbdv+MylSfRLfLZ/YoF+Fu4qD
BHISTUSiJK/njk2fSOb3NejCqU5QXVBbbzPfFPRi75P1dym8GNPf66ihKCPTp9KYkjw8f8h5MccK
1KOS9mkufJ0apc4g+92mr+sZCltVi92LuX0aBMREoIky86D8jc5BxAHYZiCww7Nvdg2Kd0eOe4Gp
HbIih8IBwOsuTFSS8WfqClgaqzJGZAAISnS56+qmG+QphZNGEcbMK69lgORHmEpdeX3TtFIJVwGJ
4LY80KCnv3dVAf33IYDSAK6nsYFd7L0SalFSmIy7AbSF/pog0iegvQv7TvbhKZGo4KSGtyt10iP9
CqmRl+LJHghkJqXg2pwwZCzGh2IyfIHiIrnotU47bxrM8jRCU2N55OhVjnxz6uDJ9I8xQfSEn4Co
wM/hCUsE3ebGPgesvkYpy8rHwHDJeg7WZiygrhLWc+o6O08GPX6TO+HMe0Y/R9FdhST7az2IHVR5
ALBaMHSI72qn6nlph8cAzby9gC6IEYK/lGyUVeuiRKbO1S/3kYnYQGf3RH2kYA6p7JAjEyHg7yYZ
dOsZ1/yFV3C0+2TpKWXWXccKp5JVdZxt8RJhnq91g3sGG6Q3y1nK7aXImAU++N99UCZV1xCNhJLZ
+952gsjh+seWF6q8logev+oAkNSmi06lX5l04bcMAP03ObGeR8r1guiLvfUOCkRDuyBrlu/M+xSD
sM3mXhNYeZElrmsGgZlx2rSXjKsR2obKQuZk+/X52U0xveVmjedfkry9REu1SBZIByK8z1oIMtd0
VkO36x+H5Us6fr6MlHja5WenTMDGiCNo7aDuF0CXUioyJnkukWouVYT4vXW+QlC2SCqMw8EpPScW
gNvg4F3JnOo99wbGFZw7Pn4RvjHIw7Ua9b/JkzKsGVL6v7hkCCCHmTVVMh6VISWq7BAgdDNz1buR
Frh0tMExtcmwrMHDRqWSXwApWvHv3be/lKd/P0sFz8ovUSB8ZWMG6PoMMab91EQkxVWpAzC+pJGJ
YFHcsVYkseQZrcnG+vWc1HR5GgKwzgV/OTtCkbjwxlkT3QiBQDPRa2DZdi9KISOFWq0owBqpVCTH
Fi9/otfz+Jm/DqqPIHFQbZZ3T4prVAIWvTjwQh6dU4foOeCN37Wl6ASHOwchA1Gy+z+WP4wbWxgt
UlNDdhXUg1cTFVyNmeCBPy1+G6RS/kzBRILJ48KAE2eQFDaClc8iDY12DLSJGvS+uBjeIcXL02+g
X/EZ6H25MeGBB7ZDCq95l/7+l/Y0tIlXmRvLLYBASsickp1xewinvlpjODh1wVJ8ItrPxDr65Y7I
yCPuzNDexINMDWL1HH57/1CdHAvA81mPTGYssjIE3fCw/diJ4pyzjcfsiQaGgFYHJ8+BjdxddZIb
mdejq8PJErAz1fPtmYE3rrb70EEUFEGD8K/VrXsTux4lQqvjQjhv0GL/8cH6k8OTAXjmIeUxbgdi
SdiP1MZVVHMYKTjBOFlKR+j1kG+msp/prulDiYWBu7ncpqYgnqjQfO4tyHd5EVhtBETsxLHCGViA
vP9mTz6WvhPM4Fg1ct55bj0TVQsqbtkY/tLJbFScQFW3NX+lsICIMSaU+YUzbeuauC5cV+0nF/Fg
F6W+TB1zAqgjUPKatuCNM5cWKUxztw7URBS7Si2rmJf6/RecXdzKGyzzQgVu9UJYM3efQtJcPLtu
EQwLWdTj9Gkwd+KLeW9BjL5LTQ3cC1gV3xNt6RzQj4Mpoo/gQcERweRxFhoEx54r57EVDxGLqCx2
/FocLUGyMyVcHRofCrisUAVIIRzmtK9uJ9Yj5z5pKIwYvEpsovE/Z9v/StY6pMrGe3RY1IBLGn+z
SkU/sN9wxJ5hLW/U6iExSgiTz6gNpnN/bpS6YFbjYm5OWKYXJuwf3KtEvFzrNJ3YVVsehSNL2+oe
PR2QI0xJi/xm17jIxZUjFIT7+Sc1GpE/oQ83nXeVApuYnNPE5YySLi7unzayKnQQVskIVKt7/N2n
4LC9jwhoJW0JgVpgmZFz0OTMbZiCAISnOPLwIq9iFsmCSRjqhj1OGK5o9TeROWa72heyi1C8CHgW
864HwlAFKhGXZgmo8jvO70geH2Qe06u72fkyr/JT9LPeixkKOWpsKjVhJA8K5wGO7WWU/bV4sp82
2ZV+844sxWz/FO04d9uWFUH6bDjyYv5uMaYHTwpeWgfirAVusq8RPd1hbuGSK123YoaPPefapcuQ
sgQEB49OZZIWb0ynvECOrDXjaXSuEnDL5RlxqJm/08sOm1i9n6+lA0isdGOf5M3MU9tIF4CWbUPS
f4MCOCC5VCqtxsXKoZN6HnG5kXwHOaS0TX2iGcAoq8eV8aFcdTLF8kjbWR8iyC4URas2jqZxxRNU
4N+e9oaL13EBmVglQsz6hM5b2E9V5OA23aOOfv1nZTP1bO1DRDVS5wT+k6IVEVO/gJqNrnbNCQKo
J4w38YTzpmgjhWR5/02uryxM6rbiOmfZU4QLPKQ7X8NlmqNw9JCuGLe/6rvL7Poc9F6C96gP0w46
nC2mKK2WzxhREkybyDmCiPIUOpbXcI6DQIHBdqC7/1A4VeIRDJY3om58rXSe+iv1fxikbmU7Y0xn
ZcPtVL41aE82mkZQ5ix5PVK8sRbbHZSYCRGY+GT3bzKA6ls+nbvutZmo1WtIjcyLspwK7v3gmndo
9uShbs8vR1FkHQxTJBcV+btFSYd1PDwqhARrjYJwlIkhUgipqBTn9YkhwLl21Bixa27VeCDbU9MH
r5UAEntwk8ODC3YOLsbkYwARR7dQ5VEByk79wmJ1ROHGynvc8dhxAzqNxNG0hbMv+zD/9/Vgq7Gk
vdSDyZVSv1rxskfgMIJi4Bsr2XeNfYS8S22vPBBu7/DlqhcM9tLR/N20F9yd7Dj73czez68lG9EN
4zs5GjIDZAmmlZ3/vpzd8ScqMRbKAwSibwWgtrm1ieQzT+8ay7ZZ2V8zulFjmlcM0HuLddSygb2r
sB6SFItM4hxf8WE3awh5wsN21jrkf17U4pg1oEBB9dEQ9ND7vc6N42d3/AdjjOF4CTQ/fbyCtENX
QCk0PyOe8w0+NrCUmV7/x0p5TG0DS9evEDrjp2CMvLV6b2Io1EQMp4i6TUakNLBEPlvmxdKF6LaJ
+onQb2mrKmKfc9oPFX7Kd9jBkStmg8w70naMdY+JPwb77lDJo5W2XJMKg7QnVGFndrxYTCjNt/00
toqXrsUOUSvOnMYHtng7rPeMk8tVNNumwgtd2a1QRh+NZwhbPhOGooDOLN6DlOdScoe02RRGSFyl
a9zdSxoLdIShFjvYV5QLMAnOjM7Z/Z4QxyTjIN93T8ErI5zRDnfSf/YOc4pB/7aQyds3/NBnOh++
xxs8kN5BttQ2zAZ0YYWucJtIJPpvIgsZOGmTKHQPdW2ev40jF+kxQxtq+BUwynAYUrhrhEpNaNyI
XFhwBg3pCSf9Q3dL2E2TYVRQ5xkw3Y7O6HfC7rWXtrtoPVVcNzIPzjVF8Ny150Z/CAP2vHmaRo2c
u5+UtmLbhOunVzvFNXL1+/8k/aLOiCrMo/x6g0aQi4jqL3M+Ex9z/Czdc3BuCNi05NlGW17D0V68
LH/sKSx5xKV1jd9IYnK+gnGheN8fnaGMxki+TH6qxjdIyQJHqYF5lj6unTL56MWl/q514T3xEfaD
Qx/GBw4hzpVIcQnZQkoQpl231PdB1PnZEpufEyJfnqyEuecT6+Xv2SJJ8BmRGQYTSB2uqG0kfHgn
ovGlpQZYP3dAUWhnW4S1OwvPfoZAHwQtwvXA59ybgVgepdo13iE+Ij3kTRTB8Udm7dVlDo9zbTfa
egdkSFzCoUoU/3KxDTOgqtIgt1aglvzzL+l0QexcK6HNi9FdSQ93flch/50g3szLJLg5I15Kv1pw
Y1IplAEEUqGAiLNyC1WP6tlX2LQcAEvaTl25gMPekg0xco3QuLRwp14MlqumGSJFolOwLOo/+uFd
wCBWSM9BK4lX22dlCPOeiq1OVjH7Drl4HI8OeMEOK9yGxFHIU3hcvtR9sk7hqIOwAebi4xEfRiVj
o/8xbZad9v/7YbGEvEbXMRrk30IV3xv8cBzrfCwj9Qbholpi857AWwnxkr19UsN8DWpT71SeEk2S
j9g83tg/5gQvaTDpiEE7JsvKI0tzgyo5C40NlK7amHQEKuG616sKJtx/5L9b7uAUOQAVusGRTRWg
fwTHiicAORjx2XSu/AwmE5JikHl6Fyr6evzFqK2DaM7V9xUK/Hut3QLs0KCCJ0110qW60mD5lSo+
03OTLGdohLVUM59X5BThmNe6UH2IDAR9L1d5dhmZ8Uk9iGYUSRyNmy3Xh9GtH8B8CnWcVohfjhE8
JBV6t0qYl8q7D19fGgbE/Cjnke685DTR/hwG+tR3bC0AbVhB7iKP8GO1oQdkcBAg/n7Ear4csIpB
eqQFRlSA2O7yGXkT4DRABJ8OHFAICGFezc/KuyfcB5T0H4vJ0opS9272KOgeIRarDfLzRp0Pky6u
gQPrYa1ZhouDxEKAiObosWCp+AYrt3lIALJrwHi4d4byDX+aN/lbT+JpOSem7qChXJYGeWmrRt26
tP3+xgjzQMEWsP1/CNJ9ZUEmWH/6H5kBIXZ249/VKADYAeKJiRpEODYBHcrxgCPcVHXIrs0fSecj
VHUY3OW2o6djvl8gI63EjNTzCgYXTfZnoc4OTvD6SQFsQjyzqpkph9wZoP3cL1AeRkBfJzt/wnpP
Vh3Et0lfXFhfEL0hgkjrkEN2tX+40DVpfRavBakrSY95DIsRztn/fUwU4sPYp4NduUdAZkb3MRcV
yJnQDk4tshYiJcZqp255LlJkGKdjchw0XEy2VF4bMAUbfdGxxtyQUWcQFsQHQV0itps31WE9BZpd
mN4YEMBMfZMwOLIftNDvdLFLHlqwGByrxNU/LumMhbMskyEDbRzCGhTD/UcZ30GHQRlrTswwbKHD
D7jTi7H5KaxcWYFPk8JaVC4MTcDb2cRS+e4G/mzESaRvbp0iyK//Ck/FftSBkeX5GfQRq8ViL44P
WFJX6DtRCHzte33kBRmf/kXt+D2Sli5+LlOzMRnppdSot38TQ478fJ2SslUAONh90BX9sSM0qjIR
BeblWRFjU/e8Ea5LLOD8XR0vjpxwnspOMjy5m9k1r4W/PdrX1AZUbpT8G9pF2UU5imoWo3goRzB0
0d5pRBuKR6Q3lryWS3PzkZ6JC5h7g2iSUe0R4T0y5bLlqQ6e1+ORjmZI6kNSwGedMbeyVWaWrata
0fR9DHlUMPXErodxda7XkpOMqqTCT7lNeIlWAfkmfVJJ0aSBd787kSl3mtpg3YUKcQ2zVn+kqRac
TCXrhSH9YE69hHqcHNFwMHkZmcdfs8BxvGVVKzU/ISyTxJ0cwKOfdpdkW76Sf1IJ5egrTbcHYFGG
f708TUCaYdOz4qMjsyqvohgNVUtW/8YqTCqCQ0yGP8gxb5wOq6HKpmmIOZP7cFX8ik5QA27KFKtW
LK12gpplJk9yiy12+0cq4epljWDFz1Cosy9MXSHCq8PG34aAhP7o+YS55yn/hxv3Q12sM9l5C69r
w4scA0TjUnfNlotkrfFjRIsJ/ygi+aQ4XNgO3a0cL8fY2u+akfs1swlDGxVgzjjXHdDvGLOomehx
XpI18aSQGDu/cIrC9zlcMxKdusD5AjcI3pDnkhHPr5A7t0vbAV+f7sfTuaerkrO8Vk1HNeoWVSvS
+12KpohKwLb8HbFEKc/SgOrNn4CeiI8OS6T9cxgM/WzbPsPk2aU7mDAkGw0SSKx/g3SUAIBdXxF8
YzPqNkn15YLG6DxV/2e7WUDPEQxgiCLCP+suFL4uHUlY5ZJLb18Dhrs0MOabWOCGVEs5135ajaOL
TV1Gywt+NlXl2keb8nx4X0eFTdjdnIRlu9m50eWGyX4SqTL1QXw3LHyqzfgcQWbSNh6vLxT+RcGd
aOXOMk8NJAbgYgKZ+blwa77b5acuO+WILQnM9aQMVvLMX9TyzHctT3vuyqpxUsia+9ZwD5aCDd9T
l7qI6UvT2ch5MTafSHFgyYbxst8FifX+3gpuAE5B1KxLPqME63WgTTrkN/o5Q4bWe34ayEl6DiTB
dHeAhf3Wu8aTz+Xak1AF2EoavoPb+lyPYZx1YYxDEZWuomSh30xIq2zNZu9bGjAzrRwwO7TzJDAF
bdrHu8Bnv4mf8NsQjVvCRkZ6sKSBX0kGsbrzPnviY4oD41fo/x9jk+OecMRJcGkAB4P+GhmyQJOT
50bCo5j74F1BJ/vRj94nCq82Rn52eRZoz1PNjeVyz2NdMeA4UDZ5BTNF81Zk2KpSO1OJHfZX/Xhn
qfHo5g26RpFTKro2bjBGDNHUeYKCm7DFmWATXCLkttCimoAyDHq9t+yHa2zzFOmPcapKXjA9ORPJ
zbSHOvjDOVkCmJXfd1Cjv9PcCZzPJtZpHAQQdC3MIdj75jfCdQGf62no46IgmREcRUnzTHPZ4Tv1
h8Y72O++hboMiAAPad3HFRz2HOvOA+rLxFi+6t1cSdI0XymPguv4nv4SXpozXp2gdRqLnGuNBunG
8YWMZZ4x+HfZXknqpxorIs8N5ngEwDYXU8NWe/EtbVykwZHa9mu+dkli2YmDLKRtxzUULLBnu9dU
d+eT4e6dheK2X+/uXW3DnN6bfcQKPconaLLyczWzsIKhbfTGYSk3zyDiLnSEbuYJQ5UL5iYENLvE
qsNBO3FJax/eo998ibTpMeD+d/GyHz5qTGgcsPg7bTsP8wFoZ+h4NVALAWfKeH/8AY0A0mLNwrW2
jeh7xqX8jdbOBgJ81xhZz8W4o6su4A5Whs7hh6HvgTwTmZAbC2fOM47CNSXQKVzv9iwJ7sW1eiNd
f/3ZQNjNwmuaMiACAL2MAT52cEpSh5etiyoAHZSHZPs/LPyrpDwyLMv1St0WW0XfbGiLPVLvtGFt
EthADOoJtqI1LUZ3MZ9u1n2sKs+ZSYAaEwk38KLOtwxOaCB1FVCsf8UdrY6cT/IWHqPdOo3L4jeD
x58ih/vOqNcYKraAYKFnHokGUh9eHM5TZ0fZ0F0iozNdaQBF5ija/fk110b7r+iSI7awQBadaiy6
PUrG7eQFz+aOFmexII3aJWtXa3jk9fDqDONwa/FoWDAVWCFYj6h4lwLRS/J+EKC168IvOhzD3pVT
1rGSfNwvG1JZV2bOOLDPH4TN+e/DSH8V5aeQPTcjFDignOL55eFObS5xAkMI4n3Ic6YZ62/zGsgw
6c3DxlKJHPB0XHDbhGezoe9WBWQw+tlhhqeMIW3JyzlICXrb3YfNFsLCuAELyyl8VAbaODEZMywk
4XFVL1p+6wGtFR4FK7rLJjA+i+GqApJjZNXIYecRW/r9nsvl9IYT3O5BISomqG0wmGSl3mbSLgHr
O4e8BlvmfozB77rn6pkAEsE9tRBG3RAy8+GSyAuktJx5vMYKjEjIz2dCEuccBfmrKUozWY94YrEP
KjVuOxfAJkg89xXN2OuLB4liSE23iV2X+iYMzWO+fCGGcyUCEupBEt1fS5enBlOiD1kK7xMUS1G6
n8VrPiH43zoC9VOkNzZL61zxHcakqzeUCalSOOStBaWvrv2RObYtEora2lmLJy6tnNq6cw/RvhtX
YMJecILCDbl2LCYQYhKDJkblNEaGEM/Gn0QMB3T0jgYGTzLkEO89s/DgSpiy6u32DoCfNVdnc8zJ
AvU2bux86t8n7XKz1udNNo1BF9TDNy598ezNB5Xab3yVNnMD637u7qKr6xXaVDkifk5Jk2V5NglM
AajDUVcXjtOsjL2vZTJOqgU2mZ/c/fg0rsraILiEDF835sxfI2eudVaCcwpe5dYT98loSz6WKlCB
u6mJWuxdcuCcaNei8JItB+TYvO0pjX5b2lbhm4FEWhDZFitD6+YL+g2NHCBIKbQ4YlCBhLQ0t8Lc
K/GCY09G8C18Hpvew2WBNDJau4vmLSFB+J8WOhFybV+Azca5XjAsBLeD8zNY4yjd1CpnzCy2KHjs
E3Fi6RpQQIjQhFOM3LZ+WQOMEtwmxMXL4jOm+H4wZN6XcOPS1ObVoLSaplJ8gxwg5fyhdeF08S0+
GW637v5cciRqyq+MkVy5Zk2O2W4KrjXBw6d7Hmx5d49LqiTn6a+ndxZfpnK2LMayA+yJBy85ISjJ
U8oBoJE9tHh9JQI2KXGdWpUwVty4bauuGO72WsV8PK2k7J5XXxTdrzGUcdgv2Zbh5ZjlZZiaCbej
YSFAE0Yny+Pe9m/QNWIhQhR4Gw==
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��F��g��^�k�<s�9�8j]��y��7@|�G�tO�;�L5zAM_J���+#y#؜_9Ɔ���D��҆]�I���������-��XL�G�rħ�b;?)�t�
�~G��y�W/2�g�y��)�ٟm&=%�kS!�*c�=���u;�755�T���/^Cs���U�6M�����c��3�3�03��4|��˰�QQtżW�>\�d{8�5o}�ZVu��������)Y�i�c)am{Z�=���~�ǁ�j���x�w�]����\t�w�i�o�c��`��I׺ң��[�&���9A���;�r�U���6����*���>�6=�w��q����=���V���_����b�:�r���Z������i#������EE���A���x�t�\�s�. �����#�.��0R�@�칽�����=��vQ�|������Y&=_��9$~�*� A|�D�*����Ϳ�%0�ɯ�H��e|�#��إ�wUMyXR�Z��EM�'4�\	�k�|��<՚�P�P$�u,y-�������� e�ʧ��'4�v,陉�dc�r����x&��^���@�+�E��T,dz����B=�t��G��?6����:�B^������+��dh=�����?����w΍#�Ϲa��Jz�ϒ/�/�l�`zYb��fa��mR1�� ��xݓ��\����<�͵b�Q�k8A��F��	�S����)�LRB3��_�N�f�+�v��s���٢KX/W[LX6��8�v�!��"�%�_�9 +.�MA��j�П1/����uE�3#D�M,�D�p��k�1�q]T)x`�������P�(2v-����e�Ш|�7�����@. �.}�(�8�<����~�=�$Zr�D�)�c��:9�!����q�y,J�;Y�&�w*Z��<C� �hG$Rs3��K��tC�ο@DX?����Ξ�ZL�	��w��J�^���Q	F��w�֢D���I����EBXV9)��öᠧ��Q&y@�r�)��Bw���dr	��+ʦ/��Uzj@���#>y��C�#X���|t �{����/'�Jˤ#�H����1}��E�Z�K٪wj� ��l��U������E8k���p���0-�W�oOe=�������_����_���upK�zsN���	�f)@�}J�����DVĮ��,���`r����K�w�"�G�8�a��1�?��a<�g� {)b��p�`]Ǎ��&� n QJy�K�;��j�J�4����7���b����$���0N��ؙBY�=.�:w�����w���!0*x]f H<�`�<<-�ٚ�A� ����6[�la�؁��xc��njB��?�ѝ�����_"�@g?�rb;�@@��G��6q�#�f@���>�+����{/�r��G�U$�z�&�4��%��%l9;����&V��M�ϛ�ª��p䨛3!j�8��~̻��;����ΰs5�Sݱ��v�����I0�??<�)БxemcwPt3���4�-���G(#�a�����6������דQ��6��.s���]?5��<�F�",ɿ)�mq<uQ��ȍ �Cg ��B�"O�o
��/�-*ɬ�c1����K�K������]�j�'f�7j���f��n�fv��(�[jNn�������[�a"�'^�~/V+S�����)e�Rjx�]����aQA�h*ɀ�TH���z9��WU�Ky���"(*��9���c0�Q�LrEc}kQv��~�������9u�u�/}�����t������f�t�s���j� ��� z�/7�D.K�u���">��Y |b�-�__oS����炨�`?*f���ea�+�qA�Hp�B�V��(v�O����?@��ې�v���Q�4�uY��״-Jz���o�ـg�]S�����Sa����!�͓���;6]�G&�gvÃ]$�"ɳ��d�t�  ȠU1��>8��/�Ѹ����vp�Ί���bL�}5{�s7妙��
�c�F�/���՞�a�lO���u�$�`d��l��S}��f/Ɖf�,���P�!��u�6�A�nY�.�:5a;a,�g=�yo��5�?W��O"��6�*:E7䬬�s[8�
���jO�S:	W��Z�|�e�,l�2L]W�~0�"e>!�3+-\Al�`���B�B�PB���� s75^�$N�,��h����;���E��X�{%�E"-��_��ag��#s��<D�2C�WE�3���[z[S�&��2�UCpSYX���*/Qi^�������ck+(k�|�"Zg��e��{��Y
B�De7�.I�c���K�z���kԷLnRA}�"�DrB�clFG�ЀV, �ƌB�Z���Ѯ�r+Oa���4��Fs/E8
ͺs�|�/P��>�'����6E�FаR��7�x5z.5�Dғ�*��z+y��b���eyuH���x]��#�9��϶p3GN�iru�!g-��	�H��߳��-(�����+��,>ǫ,���E!���J��@�|�M�\�R�& W[���F�XmP!�׆�B�&����c�:�kq�x-�ZF���[�C0���3�_�F������5!��9��@�RHgI�*icO��� � �n^�\�9�{�=$�0p�Yؓ��eg���f��CD������x�T�����ۉ�UV\�w���md̻k�)ُS��OG�%���З��g왁��J�*�Ep��E��Q2��x�U�~*��4!*Hܥ��p��b޳�f���<yoI��`��>�̮��+Ep!��|���rA & ��Z�2C(4���r���t���*�*�JC/m�DJ�l��	"�������i����MV]$�Q��Yd��Lh��y��#�"f�'dݢ���=Y�� b���@V	��N�aMFVO<��F�9��{;(�V�t݋�B��B���u��Y�4YL?�9cC£�f��H�x|s�̋N+M��>�S�](�-���n��"b9��%�������=^^���㝗������q|FG�b�_��KK�y�d9���Ȧ�$�l��n�oD���+��?��K�s G�;Gc���,��ظ�պ�]�R�p�*�g���Wq.#���G����r�_�k��T\�a���:��.�Ӧp ��I�M)�����qS`�,MŦ_*�f'Wʽ����yn��1K����y��u��җTd.�#S
&ݝy��\��>7������P�N]�A6��aA����v^W��A�Ω�N���2� A@�Ds��H�]� ���tm��C�/��B:�kr��ǶM%8���&�K�*���ʇk2��W��Ȉ��_�����#_7缣�����\��0�]PF-���C�X�χ�FU)����ң�mΩk|O�[�����85$�V�ʱy�e:W^D#�#�,`�Qz~`�-ȹ(C��둗t��Wh�h�����LW+���ET8^zY=D.O�G��u���d�� ��Y�c	��	o
�Mv�-��I�n�Ș����R!�b���~e0�����%�Eo���K*kP>7�j�b<�QuvN�ds�/�����H�w��u���b3o�_06M�/W��'��׶�f�-}�ݶ��
9����	8��|�V!�'m�l��u�~�Q��&���*�F����T�9�� �V�n�l����\�4��9i���(��Rh?�(1�;̋�����8���[��R������"��$�JC����d�vo�ՀiMf��-���
t���qgtsx1�Q�9�2j_2�)NJք7�g���/\Ȗf�*�`���$~�V�H��*Q��*��0���4K��u�����H���{w����p��h���#��7�TZ3��$:�N磨&ug_o��Դ��
Jab�3/ࣟKhՌY;���)�O�Gq�r����fѥ�WT�U}~�Ta�N����k�p�T�fC�b�F&�|w��\Is����t�	x�V�ç0�׿JJ��od�'@]�������I�̀��^�^I>!p��hG?�#	��u�7. p�� 1�\Va>��&T��Nv��:���z^�
؏���*i+U������_���2 �N�TCz���R[Ƙ�w.�b����#ˢWl�3͞�C=b�i����]Z�	[�V#�P�{�O�D�V��O�p�����L/��lp���b�.�n2���T��a�"���#�".\f�t6��hcE��ۘò�f5b���w$��,�����-C)������3i���d[Q�j���7��SM���h�*Ӌ�5'�Z
����9�QN���cT�K�0�h�����+1�,J�B�Ĳ��J��+p���] t��"�IMk
�����s���J�Y������'�_4A�9�9�v`ፃ�La�}<�Y���班Q��s{��It�i����G���E�(0��2_��H��l���	��q������T4A�"�m۞-~8����J6[�&������<�/��2b|V�����a�;��cЅ����{��Od��厕.�X��ѓHm���wkt[��e?���p�#�����߇���s�<�<��L��-�w�[a)D���Td�]a&��L��0ѰN.X��k	i� �篼�EI��۸N��Gd)��8wc�Ž_LDp"�(�_tCI��~۵��i�FiE'����1dx3�z�wR��f��/zY	&s��z�Y,�E�L7��<!��ڣY��D\�xs��Dҗ=b��!�j[=6��ƷC�S9Z�6�1�
Ӎ����\B�f��3��nW���_J���B`��w��� ���tT�"��g0�{��� Nn����uI�<�g#m�Ĉ�f�(��l`G�.S�}�������zŤ�^��j�)C����>>���]�ӊ�[�^�o,~���F`�jj��@v&[��>�	l
�T8�6X�S7��ֲM\�,�3>�O$w�=�Jvw�:�}ך>���GRgQ����K���<A�z��\���;hE���/۰�N��σ&��k
�u];��[-1���:�}3l��e��v�9�pz�:�Rڶ���O�y�9<� ���T �j�ݨCؕ`oK��2+N�n9߀����`��jd��J�T���洡�F�B��b�.��}��̀�����+�6B˫�b���AF���<��DC[��ΏL@
�(�VmH����M1,�Z�!y���oS��SrFj!�T�>>�(��+�ph	�:N}iB�z(����v�ԙd���w��c�bsA>��
Ķ���ā��"���4�E�C��q����k����m�K 	1���F��8ȉ�9�֔8�. ߉йx�:��D��iͫr�l
��&���?�i���Cg����K���|6�~3�IG�	h�T����CK*{s^��:�W��^��Mv\(/�6�$�"�7�x��%��0�΂�<�j�FџG�n��O��Ysֻ��K�9�ʛK������ +����@����Yڤ�����7�,7��&*[>h�<&�Y�~���L��kQ��N��s� �M�2v��R'�vr�Q���5F��,�@,�2=8՗:F�� sO �1fc�����v؋�7�Q��Ǚm�Й-����,3�rn��r�t��_�JxK��O�����N7���$C�`��"�wP�@��6/K�Bf�����#�P{�$8�7�U��&N< 2_
�@��PϷ�UxJŧx���I]�V����+�(�h?m|���K�[��������`p�'u�^��AC9�>p|�2a�x�%����
���a�:���?ф�
��N#p@	n�g���N��r���y1j)g��C!/qB��VW��D7��0��D|yI�P'��Yr�?�>oj^�`�2��9�˴j��;,�2ڄ@Y�\��oC�&��"��{
�������94#�5��?���\=Q��3p�\��u��{�y�_�t�|�́ܙ��`]XB��#SD=����r�i����rp��
$�a���Q*��B�՟���B�b�MUZ
�#њ�x���̀��?*m�M�(B�f�>ԡA�.⅞ʬR�������PɎ4����!��V|������j�L1�N�1E�&&�EM��p�:�?��7�)S�n!�6�o��f�g����yVjY2i1�v$3�Gsz�&�'��`�O�p� �c��K����f�@,K(�	�),���
���م���޾���2�~��B3�+�qҺ��[��F-��.���/E���*��.,��٭rl
�r�s}h�7o����0];�p�c�H��g��yU�#��џ��$k��]�\��qf"�Z��vɭj���w)�;M��i3�;��S)�e��6C
׵��~�	�x��|P�{�G��� mHz�2#_V�6̿}"���Kpz�K:?�/mo�fS��-s�d��M%y�\�r�D���;��ƪ��ڨ��C��j@����n��z��x�
R�$@�a��6�	�r�ԑ��ƻh)�h�q�u`�.���ds������R�� �]$��~�Qc=�zm�juNa3r`����^��r%�-[�����:���h6F^�񳛢�s�hAPMd@F�G�#cD�V�Z�z*���nI��J[�lm'h�$,�� ~T�YƗ^��Y˂����k�'�7�4��Ǐ�o�f�a�
+�A%�m��-�Gy������k�倏���o5Y�-$w!)��[Ok�
�f�Ü`	�=HGݔ�|x�Gٷ����������5H�~����x�8�4�Bz�}K|8*]��
Mw���{��Q����=����ba�T"������ӄ�0�($��d�mA�ɳ��@��G4uֈ���h��kHq�E#q�����	�
�������W`������F8�L�oo���y�گ��� �Z�����2���V�)t����a�O{��	���)Ԋ�a�uYP���IH��6�(و�*�މR�B��Je�S���e0+LR:(�ӝF��g����qd��e���rηI�w˺�bl��o��`�1�D�H<ּA8}2���@��b��y�_o@o7Wh��+���2�|���;���	IP��l�/�Ot��|�s�X	1a����;Q�Wx��������X����+��5�5\乡=�4=�U8'�,�@��Кr�{5�u4�i�N�D�������G�z�w����M�M��G$C4�0��Q�FrOp���-�n!�㸔V�F O)�z���^�b0��jj�U���!����u�E�͡g	�/���U�g����1��#;�m����uOˌb8s�\�_E��'c�L�A鉓U�1��{�ќ�;2��g����}%8�j���Vꑀ+�G&������T -:,)8zP�I�!��~#��o���v�����)y�e]@��������:-������c
�z��8�*��h��RJ%��B6m���4[i
:v�ʑ%�b�}k����Y�h��#�6�w?�T�g<ϟ�+��z���uw��p^�\{/V	fg���O�a'�W�Rk@=?�Db���g�����¨�a�&�_CD͊Up��Y�_�o�C b0Z��>Y=
<�G�[U�*�EHNg��7,a���M2�	 ג��`��|	���5�K5.<���a!�o$z�X�F�xY�Lw���8D!�\^�/�#z]U�\��I`l��*`wtGpe$$�Ty1<����'��Hh��)�]�aO/1"a����L�`A�/���i��k�@q?����MHe�Α�U?F.�2#�te���s})�����!�HQ�6�.U�E�K�]���!�vS6J��"ؗx�j��!9�O0c��ݻS��7 W�栭f���6�b�=b@�Ļ_`�VE}����t�FK�j�f����� ^��>{�=���jx��5�*�m�oB8,���U>x&����|�m׆[cz�WG�`!}8����\�aڛ���t� ��sa%��(P��RRP� #�k!�����!�@8�v�pM:�Ƞ_V����|���zP���9:��Ѩ伔�s����Ӣ��Y1L�N#O��j��L���'�3�Z݉M4ц';��8�"Jm3��b�/����&�ɬ�fm�4<oa�@�!�[�b�Z�U�G�����:����Z9��[]v�x�	�pCl��o���G��U�<�^+��0	��5��s���a�p3:<���w�~�N�̥���M��6�ď9�}�}p��h` yS\|N�M���6��r?���;��wmE��N�0$�1�ˮ`�`H��QC���8`�[�܂��)˯a��KoN(��0Ǌ:�'�QO��F*o�U�+���i��f`(�~׽͇�'��Ϩ�"[�����%>f!Y��=�Tu�Ց�J����boԅ��:�=���.#W0�T?�㼿�uE� #� �����:���'�,|���W��u��#ߍCc)[���T��eY�ԟ����U@//'!�.�=!ݔ�C�=o�.�I�{[�v�W<��SSRUI��A8���r?��$�ߓ�ErK�4���t�&&8��1�h�IԢP��Z�C��ש��+m&{�@!��vg�Y`��J=q2t)ɷ�:$���K��0�o���{����S����q_�;�����Q,t��F�-��\4��������o�ZA,��[�^@͌����{�� >��&K�_�p�9�܍!�*����P��f;�vM)�Pܺ��7g6�^���/{ݦg��K|Ǟ�v�y��H7�)"��r&���m�ri@��te��\���
)0T����bC~�"��8i�'
�To���lN�B�k�CC��G��)$E�$@�d�NG��M'z�����h׶9��7,v&p�E����2kK;���N7�M^��mv3���P�5�}o�\��S�����H�;�+V_q��;�?tļ�\���G��t�B����G����4ޯoXn˶�9�l�Gʾ�t
Y��:���ƃ��"��>�q�>��=��kb����{h6��L�sỤi����w���Z�&CGCr�L�K���y�~�_��^y��e|�8,��8D�n]�D��4_��D�����=���i'e�C���!~�Y����ʨ�<�`����zP N&ш+US��q��a����U���		�q_!Қ������b���q�]q�A�bG)�� yho7��ؽ-�R_�3���:h�C3T	�8h��!�Y=���s��R��MQs��j��1�Ȩ����:/���>z\��SrM�D��ǽ��JMY�r#�0��V�z�U�#��K���m��EƴZ}�D˼;%���H�i�U(�v)$�<���
͠�\�ɠaH�K����T0_�V�N���p���oy�M?]H�e�lh��GnͶ��S�(��/�����k+$5j2y�����Z�D�xa[�cX�f]�7`�;F��zw�a����Yw�Π�-X�׵�����N7`��j���m�B���t[�DIw�L���l���Ig��8��.2�t��8��Jl�'�Of��@�N(�_�ӀSd���x�-}�y���oH�?��[8�m��@+�0�/�����1Zt&<'WT�D�V��Kw�h�3 h(1?]��ɨ��2i�!!=�_.� � g�fl��lQ�yx���H��GA��Fq�"�+f��I]ta���W�?��[��W�*-�"��Q�vY}k����/ʔ���������+Z|�}��4,%]@�z�V��F�bq�J�O ���H��r�,��|�h?����f��*v"	�ܠ'I���ڐ�h��0�(k>� ��kS-?���i�}�p.\9��t��FT�j }$��JʽB1Etܷ���V�HK%<� A�3c��7���x�h�.�=��o�C	ݟ�5���v���F�fT���&����>��A�Ǎ�Ԙј�[>!��M'?���qS#����k��s�U
�)�WQ��Ғס(>0V�+����#�IK�O���Uv�t��ue�L�$/p���P%�Mi���@h^�\��~�+������kp�wK�m6b�P�}DF���׶���Q�{0EH��"+Xm)��;�\�]��M��o��\)3�|4�ϕ(*�bAF��kj�:4'���=Zb�B��+E��Q����児L�� ��<�PP�
 ��<`��_����|�C�:!ř;Y�B���'�vI ���8���G�E`�2�h��Κ�L��Z�ۮd��%"�^�����in�l����_�~�^w_X��#��Z������5��ҍY��3�w���[��s�E���3������X�) �"�K�H�>�R����}שm�$rY�ӌ����X�Mf&{��H�#�\ƂY��=����AP⠘Y}g��]҉��#�!^�Ϡ�6xE�M�Y��)�$��R��c���H�2��R���Z�/)�4sЉn�O6M�A�+�6���I`S�C��eZ�whp�Uw!���))��K:�p���p�?)�\y3>�����}���񮴔��x�7В�O�똂7�^���GA�z�t���B?��������Y�d)�]ư*����w�$àE��
HkPъ���9��/=?;v1�ZS��6�C��&�ԏ(T%.y�}�aJ�^/��n\R�F}���頶��b�D־��%)�Ӗ�]5BW�G��}�&�R�ص����;�`���{�z��}�#����� �!�����<l�He[`��{ARc"|)VIw	�I���M�֨��e�cN���1�l^X� ,b�H1���3���K(*qU��Z�DI�=���bF�vLC;m������o���g$iw��kL�,@��{R[!5�֕c y)5�L	�9BE~��I��p�(����:�-��<�@\���.��g����/ܼ�(�$�s��k���CZ�-��<+��[@c�[�k8����:A
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`�����T;�x��Zg���)U�b����\C�]ȧ�n�ig���uWg����Gb��i>������o"V�SdsR����r�x�����5�%[x�
�e`J��:������D��%�֯qd�����D}`��н6a�_�	�ͯ�m�B�jpG�zy��b:�1v�cn��H���G�#T���n��-:��L�L�;Ha͆{���{~F���pJNG���&�P�>ҿ7�Hefv��po�ڐ1��R����J�䬝|�-�|���/���'O���l/��Tp�i��7Z��Zx-~�P\`J�{*c]��RȾ����%�T��I����$:y_����_>k��R|�!KXEɁ+��J %��:v���5I��k��뱌qe����jA|4�T�>�R��@��$�qj�i^�e�^��P��坞 ��3���9%:��EV��'?O��O�����c�]�k�)���ٟ��I��R���C��p�0ȳ�<��?P�r�{��o����g�JBLH�*`�M�c�0�l��X�B��4���bJ���a�^�����Ƕ)�)�F)=���$���JE*K��'���N >�>Y�L:����6lp���F�V�I�1�{�v<#'�@�x	X�;-�j$�-�=�	���V��g��ŅQ*Z��>q���׹ss�E��]3�<m{?,����d��G#a�0;����%/����N�e4���-䣲���$U�)ӂ��Mo�d~���E͖�<�t�}���=�{�pA�G�B��z�;�Jj?,�F�7�������gu�Yr������)�ᮀ�wI؞D`�%S���]�]�O�m�ޚ�O��f�O��<����k��}
���>��j.I��L��zǖĺ^2=h_�`�i�Lkq<�������-��O �#�b�}Ff-��G̉Yl�\���GEyY����Q��-J��lA���9���̑��y���`c��-GHM?T�t��C`%�]N(��qҷY����3嶄z埼#��oT��~��\�f���r1M]��?��+�O�R�{���A��:4X�(�����g}��m�,_�0^
L��E��ujO��I.,��s��<F����\�G;MZ�{����%E9"���dS��M�"�1j/Eb��µG��]��P��^��	;��U�a�Έ_EMR2lJ���Ɛsρa;�KqE�o�b�u��)��ie̅6RX}H&��^>��S�������!n�SD|�u�1o�~`���Uyi��CqA<�<3�������*����Ex��Fَ:�ؖ ʩK4��%�`��� :C{.X9�&1�@����\u��|�6����F���� ���D�{�����R�v~oPnf�{��ulX���S�ؠ� �v�6>R�9�	t<���4�j	�l�����VWз�:�^4c���v*i@G��e����Aq��W��}�~��5���_揃e�6-c�{Y�-�t|~�B��
X����{�1�/�#+�$:��I̘��>1�OC�p8u2���^�2�(N���w�q��~��{,��P��Ұ�L��0Q��LE��������kd<�=C�����ή=v����.r�����
��Y�mҏp�-8���_~�J����v�
��$�د��X�S�VE�`#-�/�T�E��n��f�1�3I��bm�#?;��怢e��]�L��LA����1�|�y���wH��.�cZ�+0���$���T�qk�f�Y��y�'0��7�~��T�O����m!6�����eOz:vm�f��huW��	��̾�{ז���� ������M������d	��vS�2���Z��й�GQCΚؓ��H�_B	��j�%�,ݍ[O�%��t5�eα�b�|2����W~8.�N�������9E(F`���A��y�i���JwUȑ�JIG+j�x����Bi�9����8n�cָˏ�D�tJ�
m�E�Ay$\��!�c��M����{Վ��ߢ��&�|��)�N7%�ўJ��\U��o݅��l1��{⦩P8� ���6���2m�<�]�=�1�1�8o_t�B�w�m/|IyN��DIS �Q����t�;kc
#0�n,��Iv���ʾc���g��އ9���]#[��*������?��b��~��`9�G���zF�:�����S��,��(�2ɇ��.������a-L�*�,�eSM��M�'iO!�u�9��ݓ������X���\���̌�rb�x�*�KIm�³~�F
v&�%'�u�g��D�Gc�^�ޏ�ۉf>q{�tWT���I�A69�T���n#�OGG7&^��(	���cIS���n��Yjf1��aL�n�b���,�bࠆ<n ��XJ��P�`����=�wZ���I
�.y��Fk�X���)?��?U 3Y����y�y���mJJ���@YƤ�f��hܸD-k4�:�kbxv�2�\f�iQ +��;�#z�h�/8ݾq�p��Er�?��[�xZ��f��IH	�����51s���;StD��!o��6��@%����Te%1A�r�A�:��*�;�1g�X.T+.%+
~=$q笮�2c+^5]���C�������d�-�9x�c�9+�����<v�C-�ʎ'���j���d���k6J�?���#�aY�I��GA�w_����bb���L+"K	o݄0���� 6k������;���Q�2m�Xw/��d���ZN�J�'9��S�[�Z��5/�5� �������+�h��L";���.8�p�����L�;X�]��B^�������z��,�DzW�:��Ʊj�wG��vΰ&�Z����� �ݹ��w<ֈ�e �}�;ztg���g��01Ԁ@7������y��sD�(W��	�g�W'Q���쪴�v��i����<R�d�_q���tc���r�/�$�̒���R��0��2��GW�\�ߴ��v͹�ܣ#�\��ᯱ#�0��Н��]ԫ�λ��p�M��aF规W�d��7::^1���JÌ�S�3b�ST�<�m�l}�~��!�4o�.a�Rbo�*)�w�i`�&�U�|A]�`�0���ߋF���P������U�{��j�9Knk��<["f�{��P9Z�nv�.*�d�ҍ�<�?H�2U3x���m��J�0�tF��a@���>陌MsZ�[&����8p����M����M���I��꺯g.�V�ߠ8���ҿ�QH��9�_T5<��K��Pw2�|�>Kt� �*��Xg)p�3} iA�Q��s�.JH�Ao)}�����9���av	C�==S�vJ=t�*�܏���V�u�K�G��,9�b5ރ�?�ƉG��-�����_JM��!̅�[��$��1�����k�t�|%�A�8{��rx�o�ю���<���k�3�P>��/R�W��u�a�W�'�0t��P�.2@�bi��L�Q��hr�*]��֣�f�=ǥ��l����a��w�'pU������,�ǌ]����̺%¼x�����N������;i��ej��{ɋ����X�c"ޫ��8p2�uQ<���������Z^�iu��M��i �?�����@��4���7҇Id�	����M+f�U:�fB�.b�:K���@��LH��b �Ĭ�8@�M����dE��S&��vbh�7e�V��=h
�����#����a�h'��OyỴ�$��)@DW2xd��_�����+xws5�N�>��Kw!�B�z���:�)���	��� 4�V��^��	Vd�T�ld�-�7*cL��R��?�ވbծiT�^�$�q6�z��Uk�4�%��+�$��	ş4�ȃ+LH��	����ܧ$�>B�������N�E9�X�����a��kA�A���5�^₨�-�,��7@4*GH�i�nwh��
�zT�lQ$b�+k(�Uy�����o�πB���P��x��<8�C:�~�Ml� q[�C��C۩�/�Y���nLͰ`ئ�� ړ�$Ue6&��b8��j�9�DJ��4�i¼%�b�ȭ�ʃ���x^��Z32Ǿ��o-�c��CO��8�rUba�/%Ǹ�AC�+�!�+\�����#��=�N�L��#F�O�8��l/A�tD ��T�r�NY�")�P"��\�����%<Z�-�Ɏ�X��8:ش����s�`m\:�����g���:�V�ޣB��48�����N�A�?餲:���	d�O����!	_ L:��#����}]X����g݆�]d(:��Ni�>��
b�tβ�*�_K�3�0%R�iY��7�`t`�8Y~	!<����:�S[��iLʔ�Ӏ�b��unF�*Z��l�8hsK��;OU�vi��2aϲJħ|��=,/�0�r�}F���ԕ�%`�V��:�ih�����i%�۫���wX�ʗn��s�iM�{졏���6���i�"��Io�b�[�3u�>g4�i��P\��&���eB,"mH����`y~d��4�1���0U<Ui�+��z���}�?�ȣ	�6ؾ�oܬe��BzR؃�3ƛm$�,<Uk9�0���z�d4)���UND�?R=���*�X��a)B`yhɍ��A� ���|&drsB��)�w+ L��ZI~Fǅ:������R�����S�jx�ط���)�6��ve��Xq]4����(π�v1���ʓ?=���߂n�4!������jI��G\~}�Cs�Z%��WJ8��A���zU�w�UH�!f�B��O%Y�5|� o���D=����U.m��qT�ˣS�tes.L��9�8��=��?�_OT��&��;Hx��ڰ�~�"���<8]� ys��4)j
dr��>����A��5171�D��j>���[��t���!� H�\�1��K��ON��5��DR=��[�����  �3r�����.:�/�
<�'�����܋��*��"��aG�.�%C��3�@���cJ@��YW����|�%S�ͳ��~$'��`�$-�X�����,E�XJ9��4�f�NR��;k'�`o
�t�i[mVvd?����(����2<LήbP���a����e��E�=�r踊����p��ѽ��"'wB��"�M�CdYj��hQ���Nʶz ��m�_��O������_=bPi�LG�=6Ƙi���yKsC4�4~�k���5u��ޕ�1#�oU�]�����1;�=���d�7�) ,����i�J�x ��u�r��Jya��O�zl'57]�^��5��~�dk>��.]waq��C���7�*���Q�׋=�^�F4Qmk����r��=���Iq9w�c"�Eo����9xI7�a�"��&|]$�Ĺ��
�3������s���6K�u��QǹG�P��W�G��\�|�T�/q�%L�1x�k��q�V��=Nq����7��շT�md����$����/괽#��/���IE�۵x�5�>�a�?W��`C-���,=L �AԒ��?�1db�`��	�e�'�0�7⹣��@�Ƶ���qIu�:�Q
�C�qb�3�b��$�lSMΥ�֛�y�ׅT��|A�ۧoǍ�M�Z�x�2���#;��@{�DB�(��V�����3�8�C5!Jun�����K�~8����R;�rʧN~�nԒoZa+�6���D�tQ!S��YBAH^|ǃ�i�/Lzȓ��;$ے�׫�1��tתft�r��a�&,]p��N$�M:J�n���K�I�L�<��<;��7Ț���u��<�eR��+�nF�N?O�T���:�~oۇ����,���(�%���̢c�Ͼ��16�>/���&(}�S�K��1u%�{JW��9E�c*�9,	�([x*�?���p4���L���p�ɜw.\m*ؓW=�ȃ��bND�u ������T?0���g�>��/� �\X:��
E\rF�;�Ao���y��7�4#�Pc笒8f�GžOQ)�>���W�u4��m�7�|7����0��^���Y���dJ�X�?O��T�^������wҨ�^���vM/ɥGv�Eo�����&��܇�7!�x�}�o�H��*�Zs�6�GhCp�4�Ņ@Wa����?R�'I��G�_M�W�P��/
�چ}Vڲ�p���e�*T����Ǌඈm�m,�������g�ol�*c����r`G"do_i�߅�/y�j��u����6��r�J�bHt�]sn����o�F��D��Enr�dZ����9��z��W�[ A�o�����Q�%e詯MN��+;,*}�I2����g+v�.u1��`2x��T*a�w)����R0�O���O��6u�v��n�<���E���"����)#�?Q�p��A�[gT�Ty�%*�[��3���t ���
3�l���PI�x��Y#�w�>��PJ�(��晐gL4��R{����0`��1#"�7����� ����5��vb�Q_����E������^Q���m[��-����|�A�×��|T�O1S�h~,�1����v!���/B�B�FFdP�3�ܔ8���*<S�H�8��P#�`R��Mos�sU�
<�9��F��k[��ן����-[6\P��$�p�<����Z4\9���G��[� �[&>6W=o��#���b�Jk�~�� %E;��w�3�mjo-����u��0��u�̈�����EN�taM����n!Ȣ7����먋l��[��N)]���O�),id�W�'9o�uAQ��q�;�	�36���C���U�NXeA(n�V)��V��WKEC��S��8�����r+�Ć��H�	�� �K#(��kC�UQ�����7r�`�<�Db�#@���^!��0�-Ԗ�KDq��a��ޙ�yĸ��+�_Κ*�Y�UҲ�DA�����)/o���	�8���\J�n�-�~۵����|�K�,���in�Z`ݢ����oz�">�Wm\^hC�:i���rj��J���ɯ�a�V.��,����Z���ʊ����d�%�������*�A[s)K��h*Wl��[�\��4}g��)�I������1��+�����Ȯ� r��<d���TN�e�`��Փv6♥��X>��S�߷M���������m�F%���6�H����}�?V�!���F�HSN�_�Ow���$����6|�f
�C���\x���3��DS5=������O��Vמ:�K�u�Mh7F�Ԩ�"�3���A~`�M�����qapyiU
�H�T&��G�~�k��Z<A���6A=���+L3����gur ��;Bj�B�hxf����$�K��!���/��"2-�
��&��s7�W��Zj!4��}d��=���[���������ns��Պp�4*�s
������m����7֭{���t�HL����nڨ�������΃b5��2's}�c�;����ÿ>%b����7��BQixP�Ԍ`�{���9��
N��S2�0�}�D����]Y ،(D�[2Mu?k@BQ4�=����)���O�n
���'8�'���{�7bA�� �&��o'N��<��u���uM� dANZ�SR�Y�`�4�Bs}Bp��[Q�r
�B��Ҁg�`a~ t��b������L�Q�%�������(,�t$�ǐLg����� ��Hm�%]�����dK҉IR"O"��w$�A�f�PI��D�p�	�M�4K�j���ʵ�`�Cۖf���^�B�Y�?�7�VU�h����g�Ŷ[� %� 	�1�����j�.޸s�L�~�$VU퇠Bu��- z�m��~���d�-��Ɏ��P��A����IW�&��:�������%pL9���#��ˊ;>lS��Nˆ�����XX���0�j 0�E�#b�>�-�z�vU-��_>C�3���=����j4N��Դ��U��ƿF�9d0!��G����PcV�>^��i.\v���&l-ضX��2�h�,�/y�����C���t�~I��j�f�K*@��W^zu�VZڗ�{f}u
�a;GX�y�CQ�V/ J����	��fܚ&���\{.���kc!���"���<("�O���|�F�$��	N��4�N����H�:��{��6�9�A���XO)3036��ޝ�,�,��"#
���琞��@�yK`n�4�e�L!�nm�7��	��/R��q#�E6��v��s�L�f�g��7�_O�C^/��(�"?ȯY�N�c�K�z-Vm��>)�C%�;nM]XJ��+�ѐ�
}uz1��k6K���)\��>7�Hk�=�~O3O_*^_�,�����{�,�[����_U��+`�?�����0��^20�1�U8��]�CO\��M�/&a�I�GXψ�Ѷ$�E��<��x��{�}}�-��+=׆U�����ٿ|)>�4a��,+�m8w��[�y䗼��#`nʐ�Z����'�R���[�t�|�e����`�b��V
������ �cR46#	~Ǔq���"S�)s��N� k���J?����O�1�]La��f$�b3���⏷���v �R�f�/��Lv��)D�p��>�&�L� ��?S�-�$��ѧ�mRJ��pٮ�;f��Q$�L��n�:ߵ��R���q�Ua�2�3z�����k��}��'�f�R>-#_�[�vxs��K�uK*ax�Q ��P������ʕUݯ_�<���$!�
��%�p��0Y��'p�	������o�����c���sZ��~"8ޫ̄��|'V����Ю57d���:�"c��0��_�`�"8J�6��v��H��`�XMs�;��a~��j^Ь§� ���!:�t]��W�y��a���DcOk6#��H�$f5���SkYsC��I+�8��NK��w:���H���,���2��{����ёuY^@�ϟR���>^�g&����Z$]n���Z2�΂ء��Ni³�5_:à�@�66�8f�̍�R��M�����f�^��>O�X�Nw�5�L�7T�����%��}�<�\P�('�US�׌�L�xA���hE�h�!J���[5G�.�_�E��Ħ0�����˂�K�o�\��O!����A�6��!�hѽ�ZW/��l�,�+3O��e�hO�-9@��E��b���[;��qP�(E�9\3�9v�����2!�x&o_�Vhj��̀������C&D1�C��8I}O����ㄜB=�1�.�#/[-��>�󬅋*�-e��/=���>�U0͞�4^�kw�Q�V�u�s�Uv�Y�!Y �>~�{�w���{��6Z&Yl������N(����:��j����z�k��'���"T�zK,R�$P���.q��iYq$Mi2%<�Y���B[-dn�oX��d�~,�h��ͲZs�%%H��䴻~5T���<֊��*�V�n/��!4�Jw0k0Xsѥ;�쥋���3�hߛ�@��ĦN�`S��G�W�͠5��|�ld��W�9���Dc��&X�z���DD��  O*��vN��F�雝sh�FL���Y痔��/҆�+�ςR%�	~��p��_o�������Un	;��������o*.��ڕ�
�5�0���R4_�/�d?]�n���Y�Lu׼i�!m�$��2�Mw�ك��
��=R屸�����[4[.��-���}�.��5�N�0��|��� �.��6(7 �s���'L��?xu��"�?�@��f��$��OăY�8������j�	�>����7�i0��{׃�m�tr�&��:df`Nx�v�5�@�G��O��%Չj����;����e}�Ǜ�פ���Q���z��ĕ����,}>"�N�W��&e���}h���*U����cL5�U1�B@�}�?��{�n���2M�e�D��,F�/s�h��Q��G q��G�Dш&i��-��aKp3$c� ��H ����צ9a��a��ss4��"5��{���sM���h)k�H����%�JoZk�Bƞ�,��8P�1��4��/�T��դjy�̑����X[R�>�<Y�x���j �VV�"Ŵ�C��34����z�������ѲTs��;8�-���E�����Y!w�ȟ��Ez?�S�C}4�o̞t;-�;`�^��tn��d\�*iTwM0���R������i��K�q oFLv� R�!�?sS��2�.�5�,���J���͚?���=�,�=Ks�z�3 ����ܕon���� 6ॼ�I�4�p<oE�ĕ��^r�UA��Z�F̀�^b�q���G$+K~�h��^
�߁������X��xD���l��I�=�:����E�!�� V5�夒��	+����9�И�Ý�Lk�۫��)��'�+�=����oՙj�S'�Ŗ���g�A�idC6�I�b�(qac�
��+��im>���<� ��2\g�? �W�炛P�jwS����������eǻH���?�ŷ��P{PM7��� �O����]�0���@9f��A�ٷ%!Q	E1�Q;D/^u'��>�{bDd�h�wƩ�2�M�n)D�  ��=���	GE��ߪ��n��L�5��z�#�շzS�0Fx���ڧ��c��+��M��=�wczt���G#�aFbl-��֡r���2 ���a�k��Ç�=�<�"�vJ3B�QW�=�ڶ,"~���@���յּ�{��ec-×���-=�e���N'�
����0���N;P=��'�b��Uz��:�`j���ʕG:�Ҡh΁j��w��%��T��%��V�X,��.�ә�������C���qΫ�B��R�+t��/��N�iw����p�^�@�K������?-��`"����Tha1Kũ�����C��x��iW������k9�!�r:^.����[Vx���&W�������k	ѹ��d�4��Y�|��Y�CNaQ05����� ��Zb7jݿ�Zu2j���M�i`W�PD�����$w !�,S�nf:[�&� �G�ˣ�Z	/n)���.l ���O�Y�!`m�^�rrꇶ�]N�8�Q���qt�np��D�gN�]+�~s��{���w�{SJwD�m�F�YI�q�������T�!ӷe�b
�'���';�H��ls�pa�>.�a�U�Ldjs�
�q�Zc��.W���ⅳ�,^�6�G�RRlm�.�s�}T��ɸGU�#�u`�"�'%�e̥���ٕ�j��������Z���3�owKu�y��� ��[
3��	p�u����g�,N-��2n%�(�
��:'��<���i���� 
����u-�<�7��@�X)�M�Pq�l˰�= �������x�p8i�)� 6:�$�z�R󄥬e!���l��&VR;�xʤm3�=�֤�E�����nI�O��T\\�s_T�j�I2�n��4N�#�У��ڥd�݉��.#S��,�F�Ԣ��q9�yA��89�ˤi���0\k@��	]�}U�;�,��z (���#�:�Hc��s��c�]�1��I# ۉHL���*H$(^�N�������"�<�V�@�i{�7eu�����$Ʒ?߬NVh�ꙕ�>p���A�M���רO�+RW�)3��0��ޤ�E,S�-�
$��;u���]~�/㹵�%�.�S >�,g�#Z$`|�]@���Mm��q3��+�l�����K>kd7��<U]�{��f����J���^{?��ޝ���[� �V�]5�9��(KZ�ݨ!�v�
�m�.�����."�|��nc5�����?��=��;f+Ta��<t�T�c��a�ŉǐkxd��h��Wߎ��M���:;� ���~#4�8���U����M�!�pǓ�x�*=z3Iz�Pn��J<`�e���OE��	}�_�A���5)�r��U�I�u�~�PO ��U�q��bm�I[�E�6��|���\��v*U��S�d���i�uԱ�hY3u�W�;C_n��G��W�ֈ�[�2c z���˚{D����p�(�W|6z�6�w��;��F��l�fFn����.p(tɯ��K8��n�JI�6RK$�)i~�z�"��'�f�ǳɪɌ9�FG˓��^E�bۭ��O��%/�0�g_�$�)e�"��㢌���b:3���Z�MfQU��E����9\{5�f������?���6��l;d1��cQ	�mY� �}���P@�Th9/�ߓCB��9w�Ek�ޡ��U��x1���@�����EO�~�z��������X����W,5�r���3?�l�K�u�(a^��9����~|�����I�~�DF���f�4��{���S�+�Ԟ�
��Mi��3g6
0ռ�-����!������pu?�z��_#�yv����k�5��d�E����w���L�!f&�%���R��P*s�����i*r�����%Y@�&�U�L�ǂ
2)��l��f�c�n]�R2x�E�j�~j>D�\�L��j���Y揥�N���}����q����R�!���H��[�b� �25X9�z(��`�rC��r 6��0���$湁��h`���Ԫ�2��/s}���x
�M���v�%���������P�A��Y��F�� �xc�g����w���r�Q���� _c�w����g7V�^��B1�FX͒�,<#�E�j�8Y�45W"x���x+��7��� ��N��1J���+��$[�W�24���kN���c���V�N�ޯo���{$�kO./�Ӑ����I@��(R���-j�y�A�'Kw�r���m�j��gG���H���/�/?�P	HY�w9�^�獏��'��@-�u�/�=�ϧr �J���̑�4��h=�;#H�b��Do�����L>��`�P����[)�����C� ������'h:w��c�9�b&	�C��s"��Ԧx�; ��m���Sqgms��%X!s{}%��f�g_�є�n^sz��]3��	�)����Ғ��(�����Jn9g����@i�d�Y��%�>��>�8�Q�<�����fϱ\��;>�=�9�H�p�$໋,��K����٧l
�aק	������,�ҵ��(G�E�G�����7kP���6M�+� �6�/T�����X!.@���Xh�4*u��м���&�3�}}�%�	Rw�PUO�J�C�7�V�����Ȋ3���f�M2Z�-t��i�]/wOvFf�-I�{z�5�� �zl��W�Ed+�`�j�Ҁ�@'f1��)���6Y�l�6�=�B��$54C15�"����[�a-����28k���Ǽ���ԯI�Kpg�������w9������7�_}q	��k�"O�JC��-)�#������.S�{��C�מ��%��G�?G8���d�+'��������Yס�R��C�.�U��0�i(��z.H����ۅ���ԵZ����[���tC0䴶�=���8���h�Jz1C������W)y��^%�duhD%�o�4� !b���v�yO���͟�`1�zr�|n��QY`�W|����ޯ���!>��H�)��A�F�#�-3�����#4�W�l�|݄�f9u�����-�<��44�TZ���+�d*8�;���t$��z���d��s:���wl< ��b��sM��X+l9�=#@�"��u�����|)�%���w�C�)��?�gi��c�U�f��C�~����M�`�14�S���z���+vC��g�b�� >Av�ccL��ƶ�[Z$��.���f ��7^���m�4�"H��1�QD����2�'���JK��[��u5ݹFi�K)m���Χa�Y@w��([DaB^�H��YB��}���}�cCT����cp�_�Qru�@ر�{5�2n�,<��mƘ��>�<��:F� �V%!f��ۦ������H��t����;
�` 1�"9��k��K�?��$��jFm�����ck,���w�Tj�H+����f>�F���,QT�Í��-!e���Pf�n��?�?�*�1Eߪ�=GTڛ"%��N �x)��'4f?�?���}�Mfl#�D�&G}�V1����i��K�ߏ@��b�|A����ө:T�=uP-�Յ������wI�&x��u��z�E��u�È��K��_S:)k�X!���&��pD_���v4%����(������v`���7�*�\�;gv1���z�Z7�\�
؁�vB�_%����& ܓ7�2R�n�[��)����\.~� kBSA0Gt�yuZ� ᩏ����r��?x�@���<�й߱�����V?J�3�w��1?�I��>�G5}��z���2�
=�%�&:�̧"Šk���ح�Bە�ZF�5i�2
�`�ˠ=��I%�E����*n��`8�-hZy/��+�Ot����Ϳ����ȷ����B:-:
�=�E���֦3��G��W�b����mmS�2�r:~x3�0�WÂx<�[,��u�?�L���Jۃ�f!��Y^�g�!�N�R��뷯6��o�]�&��׎Db.��yy&��,�K�&��-^�dL�ZF�$	�B M	���"�O��%^�"s�>`B��#�V)���n=R�}��h������_���j�o�i�V6/��H��DAۙ�F�;M��Ś=Z��6�=�P����Ԣ�s�*4��cG����6�i���`R\
�nʖW��!>����aY(����4s>�����p�Ry�mv�J%u�u�0�7;D��JK4��n����G᧸� ���Ƨ����@zf,��d�<2���A���HZ�
������qw�v�t�Dc'�ҷ2�� ۯu�8y��$�
a��v!���so0F�_c-S=�@b�2�!$PWᾅ*�yV8����3~WP�mYu>�U�d8�'��9�Q��ȹ�B��y���բ���b<0�;���Rţ�C�ʬ0�gG�B��\yY�7�c���M��e��U$Ɏ(Q!4��em�ݚ�9 �Q��U#@���ST ��1o� $d�8oد)(��,�'p�I��{OF)@�1k��{�R
;�=2b+��[��-����]Z��䜁��n�3�T�W>��Xs�5����ك����6�:�z*U�c!&�=�Zm$�����A<b����5�u�1�<��q��ڑ�՛�"��M�N��4]�Q�Q%�۔n#�W�H��-jFqdT qd�藼���Ɖ����J��U����'8�2�
I�Z?��#�����mVW_�S7WN�#�7$(�`���kZ���j	s^���"ˡ�A3Tn.���d���������l߽OLUd�2[ڳ�<�������dѾ)���f�CC���{Q���:����^�Iu�P�@&��pt���H����D�#�;~BT���D��t�?��+�'�^G�g��U@��E���+�7����ev?�@��$��q��K�T��l��!yʣ����%�~,E����b�=*B�-�S���n����w�c��$^~���4D�k��2|��⣛Ih�3{��l�9�_6;�,[ҝ��l^��$s� �dz�/rޠ];���C�w�?s����o�O�#�I��@��\�T6Y�|�c��e���at˻]ƞ�P���IRE�f��`?�����J��)(}vnK3���pHL�Мhw��:Y���Vz��b�D��-W��։H�W�Z�2�/�}���7j_�K������q��-Z�kZ�/U��[wc���8;�����,����Zu�����J3���>E�5��:K1�kt[��|�G(�8�
�A�A���Z�����36w��n�R����(��F~I�1�F�{~D� ����Np�
�y����d�Cd�M�Zp���|�̠ghNJ���j��A��}��@�R�N��qik�`�F�T�F3��9�^��6�|�MQ�A��**F�_�š�
 duhQ*�Ú��lb��Ͱ����*��z��C�b�����2��R���U�Mz�5cN&��}ٹ�����S�l9'�@˟��;=�e!t�k}d2�¥ŋc'�E3��5�ʦ�z,�Wγ�楌�ԝ;�쯝���V����'M
�g��n��?h�İ��lJ��Hp�M !����2,e��ɯf)�i9����ӝ� �Ҥ�W^<����p1�m�>������ϙ���^�Eܓ2˝�i����'Z$2o���XS/�A"s˫	�x�0��B&�,�%�G�.?��>Z�7{����ߴe.9;-����#�����u��Ƃs�����u:���$��c���`�:���Ӫ�x#����u��>~������-�ur�aN���v���C��ª��_�<�=z�K����4\L�2}�_p� �����Z;6vZ�t�P��u�L|XW�C�U��4�tf� }OS��8�<|��tPwO�C|�D@���U�L{��v�?�V�����eYB�Z�;�|�� ���� ��A
�{׽�����sg�CI��;�\��~l�D=W�R.f���y��7r�yZ=,aP������&f�0?����hLƍ�`B[�~�����y�]S����Y�4���a�t�q�l�I�|k�����=�z*T�1���O���9���ћ��P�	!��y��H�I|jg��;D2N�W%�	��"n6��j~_l.`����4�'jo��H���[�X�M�! Np���3'r��)N���I�-kO�%Y�F��~_絁�=��
��c�5t'F+�^�8��l��	r�JM9�mJ9P��I�n��@���~UB����2D�V�<q��J����k�iL|x���M�Q��9k:��[���[U�}p�C�O�����q6�ryi�z�A���9�j��1?1�T ��Tڱ+p��V���:�E�x6.�0�kIt)��V�?�r�����x�Q�ݦ���F��&s��ټ���
"�hC>ۻU0����	4fKN1}�`����Վ���0��B����vy�[����~u��"i2���B��s`��
�(<6�z�P�ыo��h�:�!e��u��,Ju�~���2aK�
̕��{(73��Z�CJ�
����)"�x0�nFȳ�}��ߠ����[b�%��$�P�g�������������g���bTV=�Q=�9�p�kl�p����Ǿ�جe�������Sx�=/'kD�H4{�IT�!���/����.86��sz� �f0������?
j���0q�{�a�X�;uon�Տ�MB:���#z�T�x�>
���US%L�Pg��&��'����h���i5DoIAԉ�3�f���p�l��V�A`|m�}ű�
���k>B'wuB+�+�:��<!RG�ζ{�~�_U�ѳ�)	�9�D��o����VeֶRU�@x�b7��RM ��Mq٭���d�&I�΀n�+$ٶ��b��(���ɂC��Įf�>):s�)��J��~�0t��Q��hFƴX෇��a�>����6�����$ �$T�@��$`�΢���uz��W�$ß��� �z�|/�����\Z��ģ���ډԻ�\Q�NZ �l~z��� {�݆�1��w�_�kT�#N��FiH����95�.�i3���|�-�^A���ֱ��>L2���%?��TKO���?����Y�S{a�HE��<�W�tt7HpA�(|�h��	���)���З�/���1p؏�������\�K!���S���_�<{��Cu�e����or~��t.�}��X>��f͐oT�Z]~�u'����q>�R��
���'�_^�3����
y�231d\Saa�A�K�8���8J�/�w�M��CX�R��n�D���&8�W��pHh�+b��sU�}���IM�mq�m~�Jp貑�М�m�B�X�>�i�P�6���A�K��#<S�̓��A����'�Y�i�)"H��Rs��.���R�ͬ78�!(a�L"Mы�[�\�7:�0�	�q��-iw+�������B�YH�HN�Ef�'�P�LX��>A��!�J���>��|ݒl��Ͱ+_�'#` ��@��hn�����cq}}I�q��� '�3��xK]C��������k�����<	7
?p�JV`��x?�)����ۑ�K�\C��H�������� ��ߎAB~ƺ�{~qj�r{�d��%����?(%�s~� �~���D;���6{3H~㯟S/�1�4����_WX���f��T��`b��Gޜ�8z�k�gv�m�R���#�ȹ(�m�ΦL�z`Gw���3"؛������0 �C��
����:D��@}��� ��;��և^l����'�6*��X��r{#V i�=3��S'P����8bw]�^y��D�K�Aa
�Tܹ�����
��,�DQ�]�HeP�5Q���O��\Q�w)�z��ga���l�C�X��e���1���,�F���R����6PӤ�����=[�Pw�����p�F�x^�������u�>�����Ί��R�Z��6��O��`�ձ��1ۏ�oE
&&eS}�]��q&�XB���	�4&s�`x��W������=���Ƃ.! ���-%��+ْEf2�Ug��;��LʆjX����xJ���c_��q:��˓F�A\z��qə}at!7�6�\V�d߸�2	�у�y�vӤ�*i�g�R7שL%�����#��er�a�JUW����D�'��'���d�zv�b)ũ���s`w$��^�һH뤩Ɵ�	�I�=(g��٧�yFAI�������.V�0�T�w�-��%����:Y5ڛ�/�d���6�ιp�W���L^��=2��j�(A���V��x���"xwS�[��3��㋦l�=+Og��h�P�a�o����*��Og��`HѼ�����ʤ��U=�1�e��(t���u��O�v�J~�	eJsԳbhe;�����@�qu8/��UvLG`w�NnDC�7w��qH��t��~��V��c
�6%J��}l���Vsъh졨�9=s4+�StՓ��#pd����|w���ޒ�$����q�{+��ĚF�
�Oz�5c���tQ����
tor�t<ܤ��T�1u�Et�IG�i}[���.��	��ۤ�7z�S�z����Co�<�4�<��P&|B�kYhcO1��45aBdE��%��Gc\���{�NK#�4��p��	G��H���s��4�|���q1�\�b�<~ȓ3��)!t1��/<�}�d��/�/������gp�]�'NP�x:�RBi�N���@z�V�/.&3�Sq��J �˛��7eh�,��XƖ.�}x�c���*]h�:��OĪ#���c\�'�_E�àld�ޘe�ȹs$aG���N�#%zf���~����������ZS�#ǻ�;y�J񇯔�6Α(`�b�� ���ZS�Z�{�bսX��*�l��5)h���sI�X���V���=5�x�٠��Z8+�˗���NEZ���J�*��K'/��i�B%7�II&Ju�V�-=��È�����^ʈ�fB^R�I�ϊ����?�~�=#����@�Ö^Fl�ͳ'XP�O!=3/�(�ߣLw�L��|���@����FGUM��v�JF��:��8<L���Sݐz���M׊�q�?,����hL�68̊��&�wA�ֆ����xXф�J^����,De���u�e�)pZ���p'K���Q4�?E,�n����t�xKj�`m���%��%6�mfbc�\ZyCH�V�#.m����5B0{S�K�B�����h���Sw�
��$�f��]��Xʅ���h�'��;�#	H�L6���H�H~�������z��[���'A�!`A�a.��t%j'��Kk�p�@z�L�7���rM�F�:a��]4lEh���_H�__&��#�޸�ϪLߦ B啙N^�@şV4��^"�d9�Yg0�`Hq��e���q'��gG.�립�8��Q(Ā����	�x-bĕ���(�;>g���[�o>)�����Z�`󴔹nFO^�`����*���vH_�n���%���Mn��W��8|0��Yb� ߆��n�^��+�$�Z��0�2�f��=`:2���2�RYb��6lƏB�b��}`�Uŧ�Bv�]�Z	�rŹ�G�(�
����L༱|g�A Dב�CF����1n��Ә�'T(���S%J6��E�%�h,^{i*��!��ܹ�8��X��3�Orևd�� �݂?uV��ءΞ�T����F/!��;Q��.�w��#�O��M�Edh�d��Q x��h�����S���u}Z�Q�Ujp�JS��Q�iy49|15���t���Z�M;����7�ӏ��I��Bٴ�[]O�����[��S1&�F&zM}����t�z�Vf�7T����U���PGX�F�ƕ��z]I9���  O�)hr&�<���7����6�'g#��"�z埁������P���停ޯo'�obDĔ���Oϓu�FOkl�hT+W;PT@��� m��/�_J�o�Ƣ���k�9�ӓ�eO� OS��rmA�S��ˬ"�dѦ��ls��w����$��������g<5�d/�?���$���a����IHE�Ah�	\G.�n爹tp���}�6\H}Q�#�ǀˏ�_Q9Vs�)rx{���j��L����6�%E��eqiğ����.tn'A�0����c�g
����gF��<R�����hb�Ξռ��Ez��aS4��BEj�FG��^�IU�I?#�L�/kE%����c>'��S��j�C��`ݙ�Ԗ��hC�{�Һ��^d��KsH�%eYH�JH�茽/��D^}���f�k�`�Չ��|��oŹ�OzD����*���ugvo�7ΙE2��z+k�l/��C�tj߮�Iܶ���v�m�0/5��yf���ϰ�:��@=��E�2]`1�^��<��]�>���j�3����S��v���C�o�rkas�Zx��:P�wD�֢����7BKg���&N� �u�M����e��	�]q�|���@߭+��Z����TҳBX"�	��w;�Hf���@M��� �h$!g����e_e9���lD��/��k4�����a�p�00����h�^�"̪ Oմ�Wj�*{�1�cT�P^�o��/����"���|�"�T��-�d��:�@�]�X�8ڇ��Y/�.ۿ�~4aK\Z�רּs(�� -�'D�>�w(���(�dk���у����Uo����@.,�S��݅�!�&�Z�B���qĒ�_�ױ]�m�!���nMJs#ϥͺ.X9p������[�����+���DU:��Eu�tN��T,O�����.���ߌ�p���T)�dH��z53���}SO�4l@Z�K�'6�wC!IƉ���%N��.u�	�����e�����b�+��7�Zf>����
 ���꡷��s�����K�¢��Ͼ�k���~,� [%[ed7���h{`V#Ԙ[����s�<���c�Je߬����+!�5���jQ�\o��l:d�{z�f���z%�Sm�?�y�R��4d�Z}wR7��:c�>�:�� ��L���/ĉB���B٠>����Ce��!�:���+�ll [5AQ�|/��`���Bg�Qa�=���Rm%�<]�(��,��H�yI��k*N��as-��=��r��j�C�ոA*��1�t"2?�Wh��
��+Y]�]O�s>� �����CC[~��{إ��6�Nr�^�="J~���n���]��@�(,��{}�C��w�4�o����?���L�/3lO��sx�T1��p!�7� -O̓N0��dn�_�t"�be��,`�c���f�_����f�˱�Ƃ�W� ��~9Lə��(#`�EM�"J�����O6��1ï≷\�\�܂
×{�ER�8�� �֓���K��sH-�fk �������nr�J��Dd `�!X�=��{�>�m���Ŧ��뱠 V!w����b��;����DVpSX�BٛQ��2�uc֏��`�2e!{�D�C~�9����X-|n@
��Wf̥p�o����q9%=i�p����_���`P�������PMa���i�Z�[aw�Jx�Ѿ�y��o���ĩ^sz\���n걥�c�O_h��$o&�-���s�@�sm�q
u���Q<8��/|ih�/�[�{aM	CJ��kHi�GY�j�d��v�_�{"�,@���E��7�X�_�fĊ;�O��M�C���c儃{4�� \$���]V*ҲV�୲Jn�HBƂS��uQ�(�x�i��>���m�D�»77*m;T��xrpn�������
�!"ɺmxc Ƽ=��Pás$�������zu<���{=�%��,v��J*���>(j�"	hNF�[����πLl�@�~�Γ^�
��&$��6V�E�<a��	��J21��zk9��َm�QҚ������Ϥq2�Q>9F�p+�F��+��3�E�k-|����y(���ڑH/�%�W�H-�\�v<����X�uѡ��;+9����v��W��X�FqӘ��ڀ�f���Vm�c�}�h�.���(�P�~�4.c�xS'����4�-��w�}��=�,g�{�y#��f�Ō�a��`v�{K��uᣅMD&�A���'��%�;��&gGpS�SD���Ǹ��g�ò��&*\�!̃�!i1�t�Í�4��kT�so��%A?��=i ?3M������A�D?�0ވ��*[�1�+!����8 � J�Ě���+���b�h�B�+�? 9�* �>gj���56��E�F.&�P`]\{6��kf��i�<��������f�>��X� E��� uY�K�c��d�lC�}ϛc��π���,s�A�tI?\��;� �ܩ$�vj�)�ncK���;���ޟx��;��)�ؖ�������nJ�
�:��m�Si��J�K�9��-�B%�(v{���ZM�����&��r��$�b�o�`y@���P8�?ꋗ� V�wl�]�o��b�ksc����(3��|���M��<Bv&��p����̙�/��PS���9��T_���(�h|9*2�P���Oħ
��A�1����{�|�a��P7z������۫t�(�>�J}��F�w��L�}z~�|L�L0#�98	�>wJ��܂��ϿQ��"����<�C�wPj����y�)_�>*y�8T2�<tk����e����Zs�k}���ǀ�:�QS�ftM� �̓�p�x�������(�a=�������&�S����q�����(��EĎ��Ē	L��CuЊe�o��$��n�9�i�b������#��}OA�a��<9>��)���o�Ԑ{m�co�M?�0�5zˈ<��F���g8G�|����4<CO�]XbԖ0��t0U�FgΒ���$=�W��	�onPH
@D\(/C#�����Yt��@\���
�SV����I�����A9e�+�,��w� �U�u�s��X���X�zb�I��]��G� �Q$VFW/���
��y_5^~����ՏE�w|w�JU`6F(�f����Fz�	��2c'��1���ր�7�!����e�(�Z�g����/n�79j�͉hu�v���-y�P�+���#�;�6yԼ�#��_2�L��p���_H�Q��)��+\����ets�O�0��P�	�DW�AGf�'�b��<zv�tv?����ےL������1�Է��ZL�M�DR.o�-�y$�- !��v�̉�τK������Jv���U�Z�з�Q�j�(	��`�0BF�0��֙�s"N���m�����wu�i������IN.��<��4�n�p[�L�nx�V��t�t���9yƊlxwz�F%�In�1�	��"����ARDҦ[+`J�\�Rk>n��V??`>��JŤ������xg�Y$�XN��	��[�̹D�	␠����W�L�q������cW_�m|���[(�L������&��n�@�s1�h�u��a���O�$g�N`��/�i�B0�������=�	�,x�6����G�G�5�ISC�<�Ӯ�Q�}��9^��4��ʄqR��5��UW�3I��l��_.�]T��/F�@����!�����>wG{v���*@x����	�����3�?��N�uE֥���QoN��y��%�z�S���:����!U����5o�W���V
sem���@�p$�r؅���Yi��+�vH�|���	�$�qrW�����_9�^�u�N2���uGZ�^�K^R��|�z�a_}�t��J��
���"��Wѐ� 	�e�����&����r�?�z�e�P+E8�����PăG8%�5 �Ċ@{6�}�;	���B��E<X]Q���*!Yc�Ea(�/��s/�cr5����ć�ۼAF��vN.Y��.�\���xFŘ#����]Z��i�@z�{�����*�F���F�,�T�C�yBY�'�������Pk�wo���]j��}�˩'ԪP�C-�[��f�������.�M��d綡�:�j1d�L�l����>Y������2�TEy�T��9�kwl��K�~�\ML��Br�!1�ߗQ�ɭ��ˊp�!~�>\
ƴw��M.�OY֏��H�z�2��)�+�Mh�gc���I�x�(G�>Ӓ�"ew�B�,����[3�eֆ�-��?�p㦮iŎh.�:|@�Y�%��|Bo�
�LCĞg`\(�xeX
[~6��̨㣇`j>P��ӢX*�nמ�.f��*�HW����m�:��������Йƚ��� -�e��+c�-<�^����h1N����<�~-#o�������N}>U՝]Oz���n����Q��Rb������U�e�����^�j�@��}6*%�U��u��z��A���Z�V	��*~�K�w�j�VQ)N����7���v)ջjQ��zP�I��,���Ј&	S�����4?�{�1�����x�	�:#q=\���K��L�ی�Y�?���-��F�ၠ\g��W��`2&?��b�`������Ҍ
�˹�{��m����/!��b��|q�y�!��l֎JA5:�8�u�_P�U�s�]K�$�z!�]���y�l�>Hcʇ���h�}����ڃ��r���J��x@gD���@���8�5C�����SL$�b���wyj���Pdq��^c9_�V�"����#\bD
�'P)�2A��k)u�:�3�|�G�۳�=J��0�m�NB�j�0�?Ð��$tdi%t�S:e����=xlQ�~!|���7�'����2���&@�g�yEYݖ�>o�8��\�\Ѯ|�R`>�iK�2��*Cr9U��KYd�Ias���i�3-��y	N	yP�ѽɆ��DB�!+�̪3y�H�O��H�RyoӪ���P (2��:$R�zŀ���v��ɚRf�+��\��=@���O�f=��Be��	��Zj#�����*}E��7�LDdN�j��7�Va�?
 ��r�L˛fNJ[�_�+O������6��M0�n-��.��"@�����CLc��K�����VP8��֑�) �	�v�O�|z{��;o�� ��4XR�'Y���KF�H�5�#6Z���g �)b��?b���A�{g{���B�n�@����jJ�z#'�9����x�q�����T>H`�e�;>½٤�"[A�	p�lR�{���M������Z�t�*uc���Äh��8L�s�s2X"�54&�<���XWl=� �
|)B��l��T<w\Zl�޵��*	�6�aǇ��DS^�\�f��m���.F��h�q,�{�iD�x���Bg1�oȹ���v��	J��~��hɎN%����y#���m1-n�.�Q��a~���vE��ꮄTU��}*=�p��T�%q^t��yL�
J���ԙ��?���8�������̋4[���r�_f	TL�؍\Z!����@�w��/���T96���@�]�AӪ�H,j{ƥ}j�l��H���,��Z�����V�PL�JO�I�������V^`�?�Ȃ2��h��ʷ3=WdE$-'�2b�Э�8ҸI���(��|�1?�N�$�?���!����=�>�mM�2{��QiJ�ۛM�6���G7?���K����>�~׿��O_vy�ῶ���wfo#9&^�vz�O�l#P�Pm�"�潥ph�%��-�������7��p� .v#��ԝ)��&�d��1��Tΐ��B��@����0���}]MhKe�m�}�O��f^aƀ�I��`YHl˕Jġ��������l�z�{�}��;�S��	�\!0��jr�����}f��\�z�Z�&�����/)v�X%��lU�WL8Ag��������~�񽗑�����ҦHHj��]K��qq��hi� xt� 7M���`�!��=C�,O�j�t��[)r�՞dY��/~D��3tH�X�a�А�&�o�Y3����2S�^?�<��:p��U��R�2(��K����x��g԰�WP�`����rOi�n*����t$">հ�q��M3c��M�L������|�gd�߽�xT��
�V��B��;����o�U�H|K_{�"���){2[O��б:{t��#1c� %,�.\+sӇ�Q
�o�["�z��s�&U�$Gmt��/>?����� �;E�՛=���g����D����$����!�s�?[���	��j����cխ�5|g���v��"3��4v�^ﾵ��QJ�����E#��h�G$*V�nf��˯���X����s]�׌mKF?F�o"���6����͖�o����X�a�9vx(b5�;ƍ�fV��'�q�L��T���?�dd�����D�1�s���ȇ�W_HB[	��Я���J�w
�ք�ڏ��^��N����p��F����
Q�z�p6f��l��V���㽄8�^�}\��p%	��W���y�<�Y].���_qX?)�ul�/���+�=di���添>����ՅQ�E�h#$
����W�wAb ����N#���.�J�G&T�S��,�nί%ʌ��4�*�>��S���VjnL���z�%���gVM"إ�r�ddo���և�5���̋F�� �b��/r٭�@~�0�mZ/�6e�������8F\@��a��<�}�O'
�ޯ�3��yp�3$X1���Ү&-W'�aK;�h���1��2�@\��C��P�=)����a��N�zW�+l���S���B�z,]i%U3��v�ʽ9�I6D�0��$c���7��ЏW��v5,@%��fo�z%-GV�fG���y��S�� (�ے֩!P%Rh>��nk�}0�M����@�KK}�tɯ��h�����!t-~�iՑY�شzƢ�Yƃ;�&�G�!�5	��sNA]�\_��e��+V���4�$�mq�"O6��iG1;�2�􃻒�U��z)I�3�����D�x�2x���vq��)(� � y96��ӭ���<�]hx��caQ��}h������a�]�Bu^lC\$B����X�])��@5���AR��N����?�]���˓ɦ����P+���f�F�^�Sy�⩁���qj,��a�\̓S5� ���b!���"��Y��=SN�]��g��x٩J;���o��Ԟx�E�/H�)h3D�ѳ	@b�@�I���YQ\*&O�E���>܋n k�ݡ8p8��Mt��-B]������}q�R
��,Q�|u����*�s>w��3�M��M��!�2g�Q��W=;�����H]�ș`�Q�@a�t��ڤI���4�rd�gg8�h/���\��J6d�+��2?���k�
w+�gSR)����[e�k��<PxQA�,r<;���c50�%j�Ŗ�a�L,�I�=�M�(,�Zv�*:3.9\o �O%���M�a4n��~
#�!G�6s�-p%(ڛ��#\�l�MhRB�����zG�pzj1+�ڟ-���b�#�&ӹFO��\������zvH�(wY�`8���h�Õ>$9��;���mk߇c��DVPO2�[����g���+ps�~���y����r��(]Q�d��o��M�6P�A�hq!���F���̊�w�Z
P��4g(������!13Q���死�s-�����4���"I����v{h9~Ma:�@;7'cт,s�,bU�%҈�T�������a�2$>����MQx��&2%	��Jf�l�W_���G�ܢHŃm�4E�%�����%3���Kܤ��X�����_���a�rZA�O���)�b������<l�����/�� R��f{��b�ʘ�O���}�p$F��fC���պ��/'V*8=A�z�x �r����g7s]�RՍ;�o�A��e���8�$
$� M�'Sn�D�p}�'eY]�~�
K���$�ȫ
�*��f����:��:t�[��3y"U�<���A9�����.q)�^̅�q�l8�=�J���؎���;�}Ϋ�I����nK��/�]a�[� �,׊ٷP>��[��lt4G:��-��������+J'l����C���ҍ
�N����/��E9�L]V\�`�SYj����q]�d1�?m6��ĥo����d�.�~�Q�^���8�qւT���=�bK�7Vn��%t���r�]����j�2�_k[Y�?ٓ	.�h8�,Ϥ�`���l���<�,�$�jx3?F�P�0����{"ճ��f>s����h�uv���*�9+Ew%ս����|k�bj��Tиkƪ��+X��/��,m�g!�i��ӹ"e����Ƙ�ϲ�\�
��x�Y�{�
�E�KZEI7S&����m�\o��P=��9���A�=�Y����)$H���,�g|pu��4n��4 ���5��h��H����i�N?~�7�%�U%�5�.C.Қ�� x�p̵��b&��97��߳V� 20­/���H��V�1�0:֢�u���)X,Rӓ�mOS^H�+�`NB��� ��?���\�tɞ���O,#,=�[��7��In�
�����m��*���N�A�Uz��hu�?�U{6n՞ :tt;���c�"�����H��P紖3�忾��V{C=bx++�N�;ǁ�����j��� W��N�,OV=1��-tw��p��YX���N5�?�%��&��vPf�*uy�H>m����Y%��~!�$�,�^�e�W�5�ƣ���86jl\*��	�bώ��ɢv@&i����5���2)�G�_��C�Lr�I��Χ�-c�R{t0f���=.�H1R+�?L?;P��4� �D~X�%���vX��"Uh�
�:o���a�`�tTA�0�BC�4o�^ˮŧg�)ώbJV�Qv8����gz(��Z^ǫ~SU�iK��l��B �A%E��[`O;�ޝ���;8v�@B%�x�d�̀��{ ����}�j2]/�A�* */�7�B�D갌ؓY��LAذ}��-/,��,�՜2�y��~;G�����/b���rRŦ$f��%%R>n���e��� ��[�bC�&{��D5ǐat8I�|"N�PD����+�4�z�s|��S�4H�~���Ѱ��د��	n ]���?�9�_7m9W�ʊT�I����.{3�(�5�S�5�_��X`�ر{��I��w��2z�|8�q���M��@��~R���t�����T�M�LL�B�DQ�:<<��fP�ha��%e1�orKh
X`�,&�!�Gf��^n�q�ƱKֲ��^р����p��s`�9�R�L.�����֣7�˾�������Y��
��x�}Dk[gK�S��S�_�B�4��{��4�t].:8����A�M���_f�GO��V�`���.�BO������UBO��fd�����w.��κz�������Ⅻ����N܏-�dӎl��(�(�2F/G##�Δ�x�*�A��V�y��~X1�#x�������râ:@�bZJ��7*aÂ�Œn�#� X�7Ƈ~.�h�=K�dپ�t��&ض�\H��Po.�>��"i���{��!	|�:���٦��?�5ۋ~���7��vK<H��� ��������|vU;�g�[�ؚ&��a�lL«��LX��������,�K�i��"���w��v��h_ ���mu1�|2�?������Y�]�E�F\�Lk����QHC./�c;��;O���Q��?�q�K��Օ�V҃����[��oF�m	q�����\��r�-�b���}^'�V������'���0��ey6�ve�7L��n�e�����N
V�n�#fk�2��.+�l�Rz͆�������y����sU/���E���ͳ-W<��f�*=\��1N�O۾G��%���������'�;��R�NA�R����C����2O�ͪ%��C8���F�B���Ǻw���ځ:jJ86� �>��E����C$����&��"���A%f�=2��,Y��g2iR/�� 	��03C�c�e�4�=�r/����u�TEc׻��h����oe�zE�r������K��_�mq�󛇟(�Q&Y�'�DY05�ӸaX7e+"I�a���	�P���d��}&��-ZGXN�Cӿ��\�l�\��Ți6T��I
I7�{�P؝�y`�])8���Ɂ�-V�YWr�4WFz߶��\S�S��I]���Q�b�K\ Sr�&�[�S��t\��*�I�/j4]P�Ǡ�����#�B��}�!�@R��3K|���I����FN�t��
'��R�l�D�+$B��'s��LQ��^�I�HLh�"ӆ85B 1@�F����l���N��ʫ��b��v=�ň�4.�l�*WM�D�6���g��"	�)�p�VR��ݛ.+ �����7؃K��8oC��n�eT�|֕��4N���go�p�Y�Χu��o�3�������F��K��][��$�+.�]�@�!_
�A����?�ޠ� $9Yew��%E��)j�H>��u�:�E�ǃ���0��i53]�5��+��rCf4����^FB��p��y�HՆ��I��x]S�S�R�	��̺�e6����_��Ƕ��G���y�Ӯ�[D��I���D�k�-z�c��i���>��
^nt�T�u���
��dSUg�0}���T�!7�9)u�x���|�\���eI8�Ll���y'{f��j���o�1��~��7+ �S�羪���;u�)}�7,Bd/������q�����9���tj��`��P&njL�)���ۖwe@��%�\�z>���>��-#*d$K�5���S?e�6u ���W��ˏ���H��*i9	�M�ʰ���ij�'�N��pȒ-��ݼ\)������qSOG)�������A��N�ߔ�6���-�����9J����B��NV�WH��[9XN�g���a�ά�iC�|j��1�zXM �o�&"L6��]53�elr��^�%��0��gz{�����Icy��%���������=�y��T�7"l��^�D �9T�]
^��J(F�A�����2���¼	�e9O )�9��V[���k!��En��oTD6	�ڞ�������6D��	Nv��E;Q_�<��|[ �#@x��됙��nU[��L�����֌�ևb�L�􂑲y�yc.Vk��g2��lQ��
��6�[Ȳb����xϴg�ͳ̫�
%�:s	}QU����y�����`b)��͚��8���9�Aou]Ҹkn �g^�J���I[ُ�y�p_�u*u��J��ę&��4"��I�w(�*��
y��$tv��{ ����^�w��hF%���ri�W�c�׬~'�GJ?J���"S�ǅ3"C����j���/��r�����)6��w��puR-ⶀ
k��`E�4O�;��y�_whd'>���P��>R(�$�Ѥ�EB��Pw�
&p�X����E?�U4�Q����f�� ����|G�Έ�m����^�#���F�>Ҝ8؝���
 c�;�]�^��0��_I�11�ʵQ�T�����{<���q��@b���BU�45�
�P��p��e���DI��FR�SA�m7���V�/�o��~�%M:3��-��-+<��+�N��bs�I��?�~�#'�C�5�sH6&���8��GH1�ѩ
�a�M!��Q
�`z�_^�����2:�WI�F� �X4:X�����\mfz��or�g�!5�G�BT�QW�>���ۖ��F���o�ʌ$Ъl���*[�^d�h��)OJ(�Q/^�Ue���ܣ
�f���~7bPP��W�
cZ���=��M�1��5�2N�C�'*����j�	�TmХ˪�BȻ�|��hz��$���f�"��Iv�}�29o���֑#��B\ʁ ��N�d�Z���eL���#ĕ�m_Qh���P�+�:HY����Y3`i��[tKl����v|l͠�̰nng �l��K�������X��D��(ħBL𨬧p�=? ^0�6�9C/�F�@�_��Dd�w���x�
Z�-�r������7��\��o��>�n �HS0�m��ʊ��B2ax�-��P{��SMǎ���#���ѭE��A��?��Q�W��x�0�Pl3k��F^V���	5G���Fz����lű�dhJWc�����
S�#�G �i��/܄3]ʴ5�XE�:������>��W���r#���G@�c�����+�ƅÓ\�Pp/.�U�R�z-V
X4�Rd�"����V$������3�$��$l��	?Ba6W�PU�OYs���9�r�s/��[����~*
�9�Ž�Ǒ�_�0�D|�^ō�QH�HsI����C&@տ��ħ��Q���;uѬ�M�y���ޥ�ʍ�s��2�Q��H�d]��Ӆ�.]p?�]p[�j�QH�\ya�xb�}p�k��C��y���ym�;-����%�����,�>�`�R��xg��������lW5I�T���q�&a,�T���6�K���G���3��C�����OB^����o�6E����(���I�N���u�!��y�yiien�0'�Y@r#�܆y\Rf9�f��nM]����;��j6� ����x��%��|9=����NW����/�pJ��U��d��yCs>�F�b�pu�Hh
U�T�����7ΠG��	�Ȳ_o^2��%t����w�� 8l|]�	�?��ǪO1�A+�ܐK�"�i���q��#�}y,�A�Ճ)0����sʳY]�HB�o��1�� �.q�bU�V|ڽ�.D��1�@ˀ� � �3g��zF@Z�X�/0�p�uYZ�T � �	���&��b<���E����H���3�ǳ(��p1��#��f��/�9�xUCAM��s�{�	z�*�������[݀�ĉ��+5ۇmki���m��{8���F���KQ���3N��(r��d-�`�p�8�7��]NHqًR�+Tq
���	�rθ�P9�й#z y�:��`�/�T�N��? :���<>^�7��U@�X)u�r�2~Y�Xc�R�W�bx|%M��h�Y��xPF@&)�E8b*���Bt��:bz��%:�u�X���2�F��+�|�kB���Ȕ3�d^�\6��'x����W	�%�J �?��'(�ua���g d��<R�����3ߟ�2,F��k���Xm��%�g��//��2��2��	��fT��n��}E�1��jd��Q_-������+��/�=�Q��[�HM����e�P���Ԩ;S��U�(܏���&	m=���#}[6Pk�6�B��!A��+�LuKJ���\س�OC(�BN��d'���S�<� ϰ��T.a?X�?�BN �Tcr6���p"zc���Ⱥ͸Y���xB��W&s߱[ȵtxYV��)�{�҉)P��#����N9P��W�!ŘN�H����o;�4;�Df��S��t���:��Z���� -t��%}nM����9�Hr���Z ,��m+ʖ/0>&��V����'h�D1��+O5�Ufb�����J�~� !Ġ($��f��U�o���s�#�}�8�cN(~�j��T�� �\���Ѻ���SͿ��v?��1�r��Y@��\˖%��@���7�P!��5a#��@��:��7O��F�i��G��Xg�_)��|���&M$ǝ�{ j��������J�2r�Z�0t�}Dn�5)DrbG�X:��
���HZ�_���kS�/�H؉Ʊ^����Y��U��n��U�!C3���6)}�dˈf%�&�N��$��O����2��]�$����{3��8��v�2|T8��SD�ڛܣ�=��ye�Z�zJ��mۍ�"�L_!Z�|��F�iy*p��C��iG)7T�ٖ�ۼ�ܩ�Ņ�����R�ѱV�ef�)�zb*���_p(&L5[��O��� ,��>�{�o��;�H��{�����D��/�Q��*iu㡶�m�	n�F���0RD}-y[�k��IQ��Dz���P��R�d�±�%8����H��}��Z�a��禁Eh�4��O�����iuD���ī ���5k����+�ϓ��}��-W?��X�k��D��n>f�t�*o�;���F�d�M8]�%�� �!+vf��ʳ�WЊ縉я7�3"�'�8
�T���1��A�m�kT"0hHi6�������}�ʅ,�������f�'_4W;���	�A� /5e$FX��C�Jv�P��kP/�$���F(�pz_�0���{�=6��Yѝi6�zY�f\^�L��n��C�>�Z�_���jTCgM�!���46�t�|��g��M��IM��Pf���8M7$���d�i�w�"%/���Z}zv��P��S��Pq�X���M���}��Wue�tL�g�Iu���̤�V�8A��Z�?���ZF��ݓ��&B�ze�-�G��W"`	���;�����X����Fǖ)�:�$Ov��{������)�c1�h���u����_���VPVi$}�{��ړ���/��&Q�t��|׃ί):�j�Yێeȡ��QX0�W�l������R���umxb�Pa���|�
�WSXʳo��b2ë���^{w�{�Q�K@i�<�p�[	se�
ώU����塓"g���q�"�4�P�OF$�.��)n]�R��&&��SQ6�G��
��(%{b �҉�7ε�v3uĹN��i��$j
��Į
��&��-hc&�+1�wT�H��Eקv0�܄��O\�w��4�F�����!XZ	B\�����	�]J�J��-����Y�� ��{���{l�h�iM�D��b��H~�I�(5���KC7t>lЮ��
B�`�B6y��٢�g���V��ִ�@j���Q����&d��aW�*���Lt6%�gg'����3b�=X�2�(���ώKi��7[$�y������nTXq\�Z�}ߐ�]��,�����q�$����#Ԁt��|�J) }�9nSl�fF�.��eq3�7�z��1c&���Q�$?ñ�S�����>@�hT��{C(�K��i83>˨�G�,m��m��f�V�t֨t�4�]lEɪ���641!��u��"� �ή:J��˘���Z3���M���q���c���a�_BTm6U0��F�x�����4�[��ׁ��w�x��(�,����\��bi>S����HI���1��Z�
�ݢd�ؼ�ՃOΈ�Ў�*R���'Y�A�����d�{��u�Ҷ/謁
��j�QYC.�ж	%��\>��˕a�x���;E��� �E����Ą�a#�.u���Xx���@D$+@��oؼ�����ĕ�0s�h�bx�E�?2p6<w[@�4]��z���	���!X��>�=̃�az��m(��ȡ��� �g$�o�IG28��s�R�Q�F/q
��i2�^�D	"�6�o�B����o�b^b�ʓ��җ��\Y�������]^1�}ʸ�z�J�����y؛�F�d�)	HJ�6�� ���H|y�_c
�l��a��Eޘ���1]��E����b�F�Ps�7iC�)��� ��V	�Aj���5Ŭ�+����h�{Q�^�Xd��a�����fs�o�¯?]=��)��S���&�UD���OhI��ϸ�+����nY�8UG�!�~��A\NU4E!S��)����#���㳓CA���3�a����5����$@{'��~Ƚ<il��;ɇݻ-���Ѷ�G�.���#�,fIζ+>]��AR����\�,�WG�[f]��I뺕]�ݤe��v�0�'_b���.E�DV���G�D�f�<������TlU�<j���!j���|.N�_yu�&�k���w�$c�����I��:�����0������
vڈ��E���9�����Pd#��տtSF�27�����g��e�;��,����V��.�9œ-�/$�<}�����QR�[��;(�^U�:�0�`���E/ߡd��pn;".t�ێ+:t�R�rrV�v>uÏ[��r��i�T>�����;k?���5@�ȑ9L��)R�!�n�V��s�E��l����ȫ߂y�0���3y41��s7*̊���7W��p�|z`0�I�y
��7��B�eȐ��./d;�� o�M[v5c9��)���3J��[tvY �AJﲵ5�\7�J�4�lO���M�'���B:���6�2B]�����M�ю�@~���z1^uE��B�w���������9s�Q���J��<�璉��@v��L#���7�~;��/�F����9���Q�L��T��^�!z�e��~;�wh�(C��N�G+lNLN%�ċ��)�NȬt� ~�	&�Q���C��`ͩ!Aj����w�+��c��&�U�4{���
�q.���W�D�ED8��qft�ɲn�ʺ�\�x#փ����m�	oS�ABQЉ}��zؚ��¨s0{C�ݥ#�"8Ĉ!�>?�񠨌�j��/�Ե	?��[�w3��� u��{��1KĦS/�,5^ܪ��U��� �L6�V���i��е�8���� T+w�i�r�]����d����l�ʠ�~����ϵM�ބ�V��?W,�I[i���K��&ʶPl��9��9�s�u�^x�������
����쯈�q&���5�뤤Z�czw%��:�P�>6X��!Y��>���v6�]80 ����&-�Զm�A��݂n�Y%<PU�;k��ێp����<Ԇ�J�"<��c�PYK	[W�6��U� ��O#|��@Z���9i
�g�b.e�Y��|e�����PgN���~Q�XF�
BVr�_-�Ǽ���ژ�������V\��e`<ÉO�V��{���7���`�br1�D) h.�����mR�,z�o�N�j��l� �������l�}u�����ٱ	)}E��X�8f��w�n$��U	Y6m�3���wq�@�Neu{#��I}Z�;E�u��`Yy�<Bj�����D8�W��N2y\@.L�d�3��xu]�.y�R��J���ֽYᇶ��F��ԵdJ%�}�Qk(GbĘ�-K��S�ߥ^#� ܑ鳿���Mf��u��T/�/o�o������IO�������|��f$m�O��Q��H���ͷ�1���}��'U�5\B�Ǉ,ӏ��b23(�T���U��G����~7�|�����N�ҁ"� )��?�-�=s\9�MOGex6���,�9e�0�g�
*��aދ�FF��o��~�}�<���}����TH���}w�s��B�+F����y����Z����B�"Xc�����*<�~�h��=�G��*�E���/��Ԫ'�,E�B2���с�Jk� ���8]�?��3Q��V��W9�������rJ4��=�W��'�ID}V�?�:z0�C=���@�1��O��eoY���0Ƴ̐�t:ab��	�a�����Ǚ��9=5E�a�w�SJ'�����eSܽw�䃆n59�=��EW��� q�z���d�?����J��ڞ��Ae�?(���}{ƑꓫD��ĕx��W%z�h��%� ��5��� �X]"B�:[]ST{�N�IcNVs�=�x¬�3х�U���T�V�g@LQ?<�ho���K�C*Z���#�@�ɘ�wd-����4�I�?�'�hp�8l9L׏!ۄ��za��)� ������dY�^z��I��*�e��2mIv(���1���ߦ�^Iz��;@r�?�J�E�!jD�`�Ӛ���.�h}:XX�`_HK�@ ���;?'$��X��a������J{���|�T%+��q��*��2��ա��Z��ػ��R�[Y���q�?V�N% X}3c�O�ٜ[�*�ےb���\'�!x��jy�:��@l�`_��D��]����mt�'��J*#�k�1F=N�O���G|�+���n��[��W�~C+����!�U3�S�,�ʖ�T�|��f�6-zC'��f.`���p��+��L�i��\(|R���U�EE�d=RRh.�l�J�y�Ge�Lշ��7`q+��
2�	�j�$������߄�a���M���F0_
�F>�T8�7f��ȡތ$B�p���iԚqd�rY;fBjhej�DzL��$͕����m[8�ťYO�紛6�2��-	,������i�18S  �M�K�/L���a�gJ�ʎ��Cܐ3�W�
�/U�>�ϰ����Ayr�A����^�C��Y�0����z�X'�����'z���Ɋ�\�G�pZ�&%n�O閩��'J���}�.,k�MG(��d�Y��yΘ
#֧� N�܍]I� �zz;�ڶhT�Ӑ��>�y`F��Ǩ�!�
�x)�[q��b8c,E��T�ͽy<.̽B���ox�t,��_ҷqC�n>2b>%���T�{A�R�eu������ ����5-Y9R�|��t��%zk%��`�S<��m��%0�qf��G�9x�o����[��X���[-����/=ؕE�j��>̀�G!)�3�%\*�-8,���E�Q��N3���#�(�Ku.���m��4�]�c�%�棼 \ƌ�4g����O���2��N�T��ca.S��R�]GIs�t�.XO,�a�U��X��Һ��c�a;�=@b$�kʍl�)/����V뻦��6�)x�ʾ�#��0��Vz�	*w(�x�����*�9�l��J�� @��*̜Gʄ�9��X�B�c�
L~���VT;Sć���M�Ȅ��rL|֋�ʞidÈ{mV	�70��E�[e|64y��T��?b����P���/�����ב�2�z���6��
�3�_��7m��4���ٿ�{�����xM2����V�=�R�u�<���ZL�8)�"W�y�Y��dB"����K����>���A�F�^���x���=��Qz%�"Y�(�A���Dj�(a�o�5?�_�m�����%��R;:��������\|��S���#����ԋK� ����V�+X��ac�u��ݓ��!a��2D��g�(q7�N{����}\Lpe���ihqkO����G����ӎ��r�X�zY�?��$6�pg� ��揺f���
�� I�L<��#2�(~����.����6?cO~�/��8M�),ƥ4���.4u`Ҩx��
�3��o���{��@�#��j)gV��074�^"Β�&�x�b�6��E� ��pl��`V$=�|^��2U��ѸPI�8�{	�R�:,}L���e �� ��F����gQDG��r8GdZ�h������oH<���/�[�d%M?��X�nD�g���u�|zk���[�Gc&�r��UH�w�[����j���ٯ�^��ֈ�����J�eV|�4տ��'փ�ɸ]���	IpȉMt��U��
O�.+���t��h�Ʈ��Ǚ)����ԑ�7?Q�8O�<����-���\������a4Jx��V� jm�����b>�K�d��@�A���Y���n@#S9?�)*�l3Hb����|�H��G�uEy�:� ��:�؝w�v��
���}*����b�,AP�-!ᥓ���r� ϱ`���[�q!��+�8�_Hy���0E�!2�D�9�N諔?rW�n�)�ӭ^�d|ˎ��`0�+9~��u��1�V��k=� r2�#���r34S��\>4�[����_zYk��A��!��h�9/�����qA�b�O�p���!�a���^ez���W���a#��N�����{��!y���:5������lO�T[�	�O[��{�X�gmD^1�D�ڹ��k��Y;�k׃�zb���!�C ˦N�z;_�xt�t����"�,m�c�]Ƣ���>��bݽYs9��6x�ݤ�q�!�y-���z	�A��m>2\cg\���X.��%���<��2�@ձs���[�9���I�J�w��}flbr~?����<��x�bQ[Ha��|� u%�0@�*9Iqz�BaH��F�>�)���.�i ��C��AQ��]��r�^�˱KF궥t=��� �n��Ո�L&5� ����/ El_i,{!0a����Vʾ{ȉqH#i�%���$`D��D}��`��4� ��x�B�9ߟ��o����i���F�y'����}aJ	>&ϵS�٠N�~��}3�û$F��"c��H��Y���dÉs;��'�pq��`�RO�la��c�Aq~����>^���!�W�?(���_��O��;N�섟1+��rد��_��� k�AF]�޶�����'��`���D�a;��Mz=|����x8�R-�.�e��Y��`�
+��"�;/$��Ag˫�[�үN�d���1�25Tl�o��S�D��w���&	��CP�	�$Q,\�v4��۰�a��w�5�w�	��]�r����l�_�}��5*�T����_�A�l0Od�
��K���:?���YX��H��.��/��J
��	����=ʈ�9��Uճ�
�?�!,j�j��ʐB�"�^��D�ꝷ�P�F����I�<�fB�Rԟ��G j���9c#�mH��6��z:�}M�[��ȕ}���T?�[�D�*p�Aʾ0} D��Ρ� �'k�V�}�j\�ë #��0c���x9st��b�T��,��TЋ
hT�&t'r�j��E<�י�nW�80Ou���-Q����m�7�5�;ߵ��z�◡���y,`/�))RR�9(x�iC����  heU{
 ��#Z���P.���~f��B��"�&8��`�1w����|�dد��;�����.��t�@X���~���*>ka��p��?t�XJ���J���C2C��,HG�1:����"V�r�6��GF\<c�`O]�Z�wD�繉�����+B��b�z�Wtn(r�(_t��j��*���Se/�[�4��"��E8 B�g��u�	�����o~w���r3{{ȧ<�G�~�3�vX �4��k��_^w�@�6~c�z���&w\劔,~�p�Db���_�"My�:$F���}�w$�1�lH4�8u?p6�\�0���i;5M��@v���Z�UV�q�x��I	��!_	���OI%�q {�-��-w������� ��^-�3
��`��Z��9�;6x�����,�1�x�;{�[�T���$���#&�=��֪�m�SW߬o�G���貟+\0�0۟�!W74c�� �������¡Mw��7�yYn�,�u��+V����&E�S�g��嗕y�K����*Q���QߩҘ��O���%EV�W���^?�������e���a>A���0؉��鯵6?�ƚ��d�mC����"����*I�#�!��&��ײ����4�i9�d��S���
�da�ƫ �2��h�����>9z\s]���5��"D�~ӹ8�	��5�-i:dA��V8],��~�iH�����s���5�:¼�����U�[,z����[P��Pm���U��{^>��L!�P��0h�QȞO�yjʕG�Շ�y�w �ۧ�|mQ�&�h�3+�����K��m��r@g��W�`����E���>�cǸ���Ӱ�%��D��1�)�<�8�F�M֭?���D��,����%�ͣ��U`��3	�t�a�l�bՆ�d ��^�5[щ���J���ӛ��|,�� 9\+D�.�b�]��)-bCV��bj��w�Ze����cǚ��PY�)$�{�����]�?��B�WqR�QUkS�kaFP�Q�'F�l���'�y����������!�L�s �J@`U��f�8�槮��*���
+� ����`��B�4rZ� �ZC�4V�e�-�F�Ǉ|�T��9�p������hF��첩�M���r��b$o�}%���?!������띿\
إ�?�>��U�Sۺ%��f�i}\�}惦��tcP\��	�Y�pQ7B��v�}Ъ�g���ĪJ7^��RZ��ŤY+�-E�P\���9}���A}���<u;��O��滑N�dKG�������8�װ����xi ��h�Z���'��H��na�>K�`���w�%	�CRy���?~T�������Q�q��o,��nog+L���J-�FsԈD�C�S)��pyǄ/�[ʢ�ی O��_'\[[b�fH͘�����CZK����-UA�ȖHgQS���<e7��0q�i&Cܟ�$��a3Gl��$�>9J�0����U��ǜNRE�_V��_�?��g�?�&F�>��Û�~5ՙ� )��]�\��厙a�d{�M��L���+Ȝq��K�^z����sFb�zW>���v��Qn���\8�ݼ��_7���"�H6�s�M������Ҽ�l�q7	z6�G��Ś�c\W8���=�N�� �C��~'�`�P�V�ƘO��+?.I�&G��Y9�08l	�ԣ�=D��`��|��tr����e��o�M�z�Ĭ@��lD���I��@;%��P��㵌�i Ԛ7��0/�.����=��J����<�d1D�� �9w�l>�!�CI���>wۿ���9,��Q�	J����k	��UF�G�eu�-A�t(�I;9ˮ�"��{�x�gý:A ��3��6���#W������܋>����"�6�˖K!R�|��A&&O����a�YY�'Xh���2�\��~�)��)�ʲF�~���< ܄�N���Af��w^�)u'��P�;*�!P����O7��f���=��ja��=�~~e@� mW�����GE���:wH��0�����l�戧svT�tTY��N{��������lݨR}����a�?z��ˮv|o��*<]�]of .8�7�ݚΞ��?�J������.]�v1��� ���������%�N)2��
ǓM�������!V��;�e�ոWt�=�F�F����?�Ϸ�)Ya|��th拉��jS�sJ!�PY�:����y�"�+@� ܹʢ-�	r�(�^�hȢl��M5^J��u�Ļ}�凍���s;7�N
d���#G�9�"��m~~��D�gy�w�trYE�xJ-�� ?\����Yߍ�������%�����p�y=�Ǧ���Lɝ��A�[!í(���Ԡ���c�~%��媴1�F~�T:�����B�g�T���V$·wRQ����`�q&�C��f�;�y{��s%�}�g����aL�a��ũgZ%�t���d���};-o��hH�����M��*���0�ՄvL��h8��[����e��D�'�������|#���&w�+8�\��rU�7� ;{�ɩ���[3`os��4���v&���_y��Y��PD9��L���:�	]����ՙ�	/^=ۑ��|����s@�mye���k�5N���'Q��.���_�R�>fV;fA!�x }W���	��A)���\C�+͠n�pE�|��<@k�0'Od�@f9�\�J1�J�|<�+��
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��YNqeb�����-���	�^aE��u\s�=��4�4�5cR�jQ��I���Aѿc��tͯ�8GdPT8ȵ~��Gue4аB��O��k�!>Ny/�0�7��~ef���-ǌ�h�j�g.��[�v�7�C�����.�E>�/���g��`0��O���=���]X���eWVS��������C���C����H�ѐ];�[z��2^��~������T3���!)���@}��8]�����z�'Cݒ���
�ZmX���H�����	3��S�] �0;�7𼼦4;�	��&J|�k+��KK���M���̚A��Ӹxx��E��D�`z��>�\��	��<P��w�o�!�Y�S�E�۱^u3DU6 u���mc�����<��rp�t4� �}{�ʐ�^�vL�I:j[�adю���n7f�_b"��|�5���SB�n�萲z��1޴���qNWB����a�^��dE�m.��M�����[��S�/W'��(�Xu���q4����0�ڑ�Opd/KZ��X<M���Al���7	 &xqP>��.\����6�
�����b�p�ʥ�a��tTameW����<�v\�*����c��_&����ݼ"\�z_hʏ�LZ`���.��	���a���[��}��`ii��謡�RA��.�\S?���.�"d�����E ��_��f7]89r����`ɻ�~�)�t��+��<����1C�TzIaeD�����A�$3V�9�Y��bH������̍�r��y��y"~;z�)����ſB�.�f�.U�j��c{�
��s�rS�52l��B��
B���
T"@��:���}��v�0����;��Y�e�RC��Cy_�B��n���KQ/��`��?;��ʀD���v�3 ��_,���˹�����(1d��;�4~����n����<L?�T;�{�� ��f���1����F�K�d�{QK���Y��O��`���� d�-��5<�V�91�M��)|��R�Y��LW��E�cxC.�Q9�����nn�T���Ok輲�X���H J��[�7��h4{ c�-�s^�K�1|�&���EV8�,$��[OABv������d[՟��+v�0^ᒒ�U�p/�r6�s[\��\+�yM7D�B����Z�H�:6p��d�LF�\���հ9q�H�đ�$�Y\2w;�������c˽�bb��J�ǈ �U:���B�E����9k���SI����]�����V$,����b�=�p&��F%�"�	��<'���A�s�قJt�Q�����z�Y��H�Eb�u���J���}X��1SI��L��?/���I��j@�4������[\f���!�^}���~������BVzՊ��
�P�q����"�)�pޭ�$��ͧ�mѣNx���,��<si�s�,�9x�aW$:����kn}
��rS�jmʾ��m�e�,d@ZV S�Y���6��m��/Ct�?go�I�������Lh�T���.�\���t�5�@�f�9���|�@��w�u�@�5�)i�z�Dj����u�	m~|�;P�%�4�we���.]��:;���|�+���z�cLQB7.H���BC�N�f�a�������Q�7�xU�h7�11�d�!���:��� ��H��0�O�bt��A1$@{�╸U��q���֌��uY�}�7��5�u锝v�A�h��+٩��r͎
�s�Mii��֚Zl
ؗ��~A�N�:���6Ehi�)�K�u5v	�Vq�m��[��_�O��\�Z��
�߭�k��{y����_I�+�J�k�JK�s�$���J��@W�lBB��	ߏ�z��������1NM{j��ܿ&��ܙu$��#�Ǻb��z����[JÍ?����|�����u�,,Hq�� �2�߳���)�*��܋�Bl�D� �3�FyB�l�Mv~��~-��t���
���YA��lY?7G��^�( �}�t%��!��ڨi SxQ���?{�3�����uΡ�1����~��(VQ��,�;KT'�e�K
 n��tE�G�O���/��L���+ �m�\����,�g��~8OY���}XD>48t.�n�ٕ�
P�֚5����*��r������^kM\z̡���'�\岎'^�����w�|�?��i���[������{��*Z��RS����
���D��<27m���0�ġR�z���M}6�P�����X�|Y3Z]�~
صµ�b�QN����N�f8C�F��{ �7��l�\���<�o�u�]i�A�� q�`KF��B�۸yܙ�a��
fLY�����,�5>���G�\�y�*,z$��%����p�$����x�!�2��� f���|���y�j�͘a��0�B*��a�SZxG2��"L���1�Uw4����&��@����U���)M��q�n>�R�P��� /����t*UU@�'�-��'DvL�Ǯ{�� �[U�e����쎼�_s��6-���kHO��[G���t�ߖb�S��s1!�b���I& �O8�/<>.���0�c�
E���m�ROj�9�����i,R���<_�����<'��y7�=�`Jfd����)ĝ�X�/|o�×e�t��[�`X�{z���7��\�Fϡ<t;�Um5t˄�E�vfN����,9�	���ao�T|�q"bF�!���P&�JԟQ���6���wG]>�[ �3��=ɓ黑Y{�k3$��ri���ud�T��+YO�����B����Wڦ)�T����w�I��xVzyT��`�r���@�O��=�;�LT<SM"4�����T	l�e�^��a'V�E�0�2.�z����;e�E�{���!�a8��[S߂H��y�d�EZ�'��S������d�T�R����0�1C�T�	�#�f|����< �����IvE
v[41oj{�
�u@$Dя��E��S.Y쁜<P-�ܧm�W~�S�6���� �m�^��z�$s္Ӫq�	�� ��vl�����}N�R>��i�7$(�A��
�'�KdIf���Q^�Xg&.�\xQ?���W�kv�]��N�h�����Ry77��m��G�����k.�3d�%E�R�O�A�o����� U�o�2�$?�,��̤;�rE�o��|�ͦ1�#7ǆ����6T��d��;�v6m�&Un$���6�y.�`��t��������T���� O+8���`	�'ēױ��D6h�E	�� �E�g̨֦ �u��'���d����k�[���Հ�E����\���=�"�L��� m6��7-=3(��S/��j����i� ����������ċa��_�M|׫YF�下���`��'�˃���aiq�vVG�#�˲�^�Ф-�#W!�mE���0�Ni��^M5��s9����s|=q�I��	OZV�ط���K�r��� 1�a�kc$Z�.�KƮF�[��GקBy�߷4�(>���N1�O�M<U�X�ΎÃ���FR��cV�9�#�_��+<q�N�r�,��&�*�נ��A� ܷ�7�
�f��iM���'w�f�a|W����8x�c�P>�9FȔS���aY#s/U&�������r�,��$ŹnI���$wht��(�F6f�Ӡ4��v���~S_޾�mL�۝�w�#{G�Z�h�5h4m����E\���"��.�ts�I�+�so����J�Q�m� ���`�朿��u}	S�q����HK1H���:�ɻ�6f"y�$C6x;�ɹR�$�%�B	��M���]�oB��Wk�2cή��K�E�����bC�9�c*���E6��WVq������v�ON<�!�Hh�p�s������<̳��0=�2G�:h����*�  Qyo�"ҵ���o#��H/���T��0B�3�0�#�6���EE�JV��O5�����g����xQ�2����gc�n��t�x�w������u�y�*gw9�A� c��F�����e�����ҹ�u@S^ .��-�O�oAp���#tk�{p�cÚ�p^X{����*�,Y.���Td<��f�-�>y�#�1���_`H{C��;"�����i��
ʆR-H<�ED��]�A�|^ab�����Q��Dc�*��2��2�Mƍ�=�Y4�s´z߿��0d���ՙ#A�{*�)�fvY�-Bu���g�6�n˼�+c/C"�H1�lE�wI�%� c�~p{�!A��3�mX��A�Jd�VNi�P���������o�^(=a ��SBX*��X��%x̅�k���S�����a5��c^+��Gò��/�]Q�6���3�7\�;��⯼J�FmjiNv�p�lh#���6�"���ÎfXt�C�f������2@������q&M�NSfg{�E@I�A'3p�a�Ю����lQm�r������aRX�+~��%F�:6�YojwTh�v*��_���&�EC�	�Q�a���b��B�w���|],	r��?��!�� g�F�b^���UcG`�۟��b�����K Xʫ}n�w~�����\��kd��b���?t��i)k<�\�	�A��-ё�u!n���	�yλPq�.k���0G ��u*����n?�Lo�9/����i~OV���Fcc-O W�!j[����Z�
&["�o|�/oEA5����q���:����|��f����:F�PT7���ƈ'��v����P���l	���`xx;{��<Q�c1\��:]��
�<���" 5���d�B�늂ެ��''�Y0+������=�?�{)9��F/m�k?b'㏭Ö���h�r�]��IѥL�M^䙪3���B1m|�wR3&t� ���Xnr������V#��#a�����^&P�sNG�̤��3�> ��(�/l� _:��<����۠�A��r�[�>L�.e��/���������z҂W�2��N�̠��������l˅�N8_p~{|ߞ����}V���*�=q�;ו�MGF����#N�ך�3�&6^�S?�3�	���f߲�k.Xsd���I�Kǐ����+��ň-:�oTޱ���۽����0��sx9cu<����+CC�	*A��uT�qbg�c��� GP�+p:V���������z���R��8V���!�j�RP�@VN����]<ޱ��z�-�H/��F҈�hs]:���a�
y�NQor�sZ�/���v����J���(wT��/<f3C\^-~�ڝ��K۝q���z
L'i���ߏG����.BcO*�@���9��f�Z��u����ߐ/|���]9/�f��L�a�o�&�!)�M1��i�m�6��l�v�3$�'p�V㾑�Hyn�~�e�:)��vVrzFĕ[Cg3P�'�Imir>�I�w���:����K⼠֘̈.Q�I��gC'�������U�:�@�Kb�:Jj����庿(���0�?5��G�nH%v�Gr�F��O���d�W�0s�]�j�}k�I�xu�#�:U�|$j���@h�!�qǠ�vN��%�̺>��Nr�x9n���5'�$2$%٪[������a� S�~Q��*��.�ΜOz?	�����Ӿ�;4� c�R��v���H�j6�5����'l���>���~����b�Lx�\��
h�r@*�I&4H��c+NT�,�K��ϵ�t6p�5$�r��Z*��j�|{����l��*m���Am�RYRd�;Ts������m�}Nt;-�v6^��KL�3�sp�B��ж%�"ʫ��p^`b�|q���22�V�G77��c����~�Yp+��]���BAS�2�/�#?��zɬfB|�%NêpM���L񗺈[j�y�F���-Qtq��yǧ>�k뚾{ꤪ=q�&�E9�G��R��f�e~��������g�1�8��M��\�gɅ�i�$9s�R���pj&5�P�����k3ڣ�)$�K"�g/8���
�u*h�~!����I4U]�{��a�}�����|��/�t�6����Q�n �z	�o��i�=�	30i����fKe]�7��3P��
���U
[/��jz7�K��_�}�	6�����b�u��a��cJ�Ƥͻ����\M����ǒ����Uu�n(?�/���wl�6��5�E�v�s�!�^�Х�Uq6�*�_���"Zc~PG�y��MQ�,�[�-]lF��>ˁ�R�e|��[��#�����,A�u�"�5 /P�w���Q&,��q�c�������q���ѿR :$iY!��$\W�moMV�F	�KS�9:R/��Y*ݚ��4ڒ9з`����F�9�7����I��X���W�9k��1�y���]]*C���dëLT�L��lpn'4 (D��=���o���j,Bp���]H�Mpm渣h8/�p��U���;����Ǹy	������0(�1��r�U-��r�<P��}_�,�7Nj�~wp�b:z-"z�9��~��z�$��ա�@�ȋ+�wJ��E�ւ!\�X�7�k҈����U�a�k%|
�0�}�-"ũ�t΀���N�ݨP�6r�Ew�p���a�p;W��!ʦ�>�{,L��/	Dtt��<�D~�����X�`����S���,�X�К�3E�(�h�e�� >f��'G=P���:�v��	 h�E�;(���0�v��\#��|m�0�L��0���W�.��ld�2�5����y|2 '�ɲ�4xE9��j���g��biT��Q^�h�	���U����pR_���]���R/���?����^�u׎qo�#�����`䙆Hw9+|�P��d?->�N(\7���[7��wn��v'q� �Y��=Qñ�0��7�*���h�D��<TaV�r�єN$)���eJ;�g�~�~2nsJ��A	V�mŮ�Cl�IP��L'P<r������-��*��GW�?i�w���D9�|��ƌ�l�r��qT�s;Ą���w�p�Y�W8�iD�������(p�c��w���}�ʗ����6&"�g���`��h��0�:��C̀v.���ZS��K(=�gշ�F;3A�L���;W�m����t�/��%e�Y�@�Q�NCq�v���q7��&�)DLB0����0)زʄ�cb" b jDR�R���a{ՑV��-��KY���ʞ2�<HC����a�UWKea�y�g� ��$%������>�Hx�-���S�Q�'�˜�p�яGi;!#��ʉ�2l4D�o�����R�3�eJ���g�]�3�=ݮ���wL1>��K��[���sGRޤH�P/�֔k[���pUC��	�؟��V�W{:�]M�6�z���w{�bb\�+�d�B9����\a���Z���=q�}���1K8�0�R&_
���Ʌ�tM�DJ# Jћ��K�%�V3����pw�*���i��M[с�5��н��"��ֳe6Έ[�fPp�����Ґ�E/����,#��,��k�hv��.����L�z�0ݺ;�ܵF�f��D)��c�a���(FPP�Xn����z9�����% \���#02�e8�ͅ��	��:Q�l����T��a<����t�^����̍3`/Qd�z���mͼ���x�?LQ�U�'�L�\��5-���Ȉ�ݻjL*E(�~���J�
b�
2[Q8�p2E9w�͸Ǟ8kJ�<������o��cC��n��F<a��	<Τ6K�%�#pT��������E9b�#��{"4���9I���^4��z_����s�}�2��C�b(����h������5��l�Jbk:��O�7��v��k "�#^��@`T�ej�䜟7�i�/5��Vw�(DCɠ2��ԏZ
@d{6,�@ls�n�Zhz&w��w��.�N��`��:���/Gi�~ɓ��O������b���]%{> �h��9I�TCg^b�c����Ԫ	N�ا���<��0�-�\���5FtZ/w�[���Ϧ��ǘw�e� aD���S?��ݗ	����Y�Ba�&��]W/��J-<����>H����7�p���_Ƴe��/�z�-�� )8=��R�^�9��Z���L��7P�ES��`HC�%��..NH���<��S��֗��M��%H{y%��,֕=�7�G�-	�hkْ�qLV�c������=�q��_�z'h�#�t�>@�b�X��?��var�wt\�(��җ=4��ͳq��
8��o�?��֕��������!�����>����$ҢJ�TC��ұ~*����9�<�Qe���S���#��)���ī	���5[��V_5�&ZS�޾b��ĺR��=�*��ƅ:��1�x4�����mb���x�l n�5�g��Z�=v�X�j!�o����tZ����2.����H�$���,^YҀ:U�
�+M�3�J�&��G���4-��� 8a��j�Z����Q�Ѩ_ؠ��:��NF�:D�:����-�B)~�u��?���TE;�O.��ì����7Ojص�b�=��|��v� vE��dQ�8-�����8��[�
�=�n5�v�Z5�@)˜s+'S��EWy�a�!{�ۄrH�s�]�i��#�W��(������p?�;����!�n�pt��@l���]RXy�E#X"rư3|u�-�&�@�1m��3`I��KBtm�]y�����7r� ����߃��dAf_~-~�Fg�ݲ��_�Y�]��d͠,�;�EM����;�%~�� װ�g;\���퍽�MK(�8$.��������@�fH����]z�c̢��O�#��w����y����:����E܉ARHn�fK��bh���R{_�N	��b�2~���s�ng1�U�c����.P���3��O@�{�}"&+3�(`̋�Xui���w3U<���C]�+�-�!v�ġ5�-�����,��jY���n���bZ��p]���+ <<o�M����=3�W��vJGoG5��Q��w1v�YᝢW����g��\�]F�����%���p�igSA
bX*'E�-��=��W�m4��L-���zK�}}n�`÷D� �^��j�x�^�v M	�b�۷��q��Z�J5��y1%/�e+�K�=�^�#=��/��s����4s|�����e[h���w��?��G��9ߔG�"���4*A�#�`�v
c��t�!��ً���Y��IAZ������^��p��q�
w=N���9�@��<���#��@ �/��N�'��&�"Z���u`lMt��!�g��i~:�o8�%�Ɋ�q7�K&w�_���Gs@���H�M�@T�h/4��PY�֔�yyC�8??6�ZJx���Ub���>s@'5�Ո'g�2-���r���:�#B��IB��L܎�*���ƚ�O�� �1�B�AϮ
'ح3��)s�un���T��3��R�>�,�B��y^�K���Ϭ����/�yp��1>���	��{?|�k����&��;�uWˎ-�%%6�h�u<���3�[�;�� 00��[8�έ� i1&'�0�	I��7��$rc�kX���]�Pٞ��z��e[�̌�ԫ{	p/�P����z�*�_%N%"��c-�� ������\Hmd��cȾ;P�g�#j�qA�,YC 9Y��@;I�F���1f� ����s���)o��Īek<��-7`:I�u%c�MY-����+�o{jW��F80��ƽ�<`s`���!�0�
r��QΓ��Cr9Х��^ʄ��(I���N�)�W�~>h1�)�)r�^�Ðq�fHl�$,]��Z*�ـwGJ�7Z�B�)r�T��]���I�}�����5it?�S��Ճ�����dy�y�4d\^Y1�/��P��1�ۘ�?��*��d@j'�g$���h�WmՊQ<��!0���~���ۅ~T�AO�fh�l0�V��̟�rՃu61����
*�ȿ��r��fr�����0�+�;R�P�����5h�J����h�2�jsz�"86c4�l�ٗ������D�(|��1�܂銌r���08�8?]h;HE�1R:j`-pϨ`�z!����D"�Y�
࿦��|�\:��_��̬>fu'�j4Rb朏�������.�Y��wm<�30m��C�K�o�s\�&:�IG�=`�m��[����E�S�6������[��
�U��ݱ�i��G�s#�-e:52� @����~蹢@.�_�IR�)�B��׀�9�|�joqM�ynV�$؟GL�/�j%�����s8�J�!
������`����Xi�p��{`y�b ߪ������t��_!���Wz�k��O/�hHQ�ə���F�$�-�6Y��P" iL�ʒ)Jš�6�M�}Yx)x� +�U��{�>�=m�Tf�2b�&��+�<Z�
��@nشa>���į����o��{s��"�����E"Lp{ۤ
[n���Ĳٽ��m������}���Re��GhV�-�����WB�vw�m��\?�2�9�X��Q�FC;՞`�TY���7�Ȇ*J��w4��6�g�c1:�������T�w��ړ�g�C/X��91�& �ے�>��@(��b5�ʂ̔C��N�G^TR�#�R>o]HA��Ŭ��ؼſ~~z�c5�Q��(�8ph������f�m���L���r�xb���w{a�hٮ�a��h�/ܶc�������ƙ�(���8c_��[�~�Yѽ���{�`V�e��Q#�J��-(�H1�`���]����~rV�S�.k�婨|r8tԴ9/�U@+�7Rk$��QM�(���g�9���t0ɚ�'����M�F����q�/��<,���n��Hf��Cg�XK�0q��H������O��Qm�K�Յ{����p�jL/G#�5t[�6��H�v=���Y$�]��$���`�n�){*K����Z/�-�r-p��j1z��H�9�G�����J�� ?l���J�1�~�n� "��0�	K���ޤ���m:zS��J�Z0�����}�8j��ON� �b6
��ul��``�ש]�y^8q�g�0��OD��	�_��\�ij8�/���"KAI+�N�a�_BN�}D�s�+>�]�={�`9Z�fl؎M6Ņ8o��K��(��6W��v��#ށ���k���ہy"��J��]�J���r���_���!��	����i�{�_ޙ�y��F
&�$�n�✥����R8���A�-��p��*��?�3��#�#ղ&�%��Gt�D��}l�+L4z	�V(�l�2�nZ�c������z��$�F��c8������/�K��}`T�DjZ��/����Ư��;k�����]wX��3�9q&�5�Ȝ(<��e��?4>�ڹP���^Y
�H�zQT��V�v��jPD��o����n˻(s2�y�v@�q�AeR�^�ӆH<���Rz�}X!7��.r\��y�"j��˱�����uS���`�����Y��%Ǫ���ӅZ�Ś ��`�l�*kY�&(��A9I�y�+ ����Z�Wa�(=��4��y��x��7���uB�yߚdH4���<�(�����T����-ܹv��2���{���w��`x��� ="-�(�fE���7�
�Y��� ��,q�"6M�$�:
EhK���f�[i�^Y���o�3E�@�g�o�5��oz��b�Y��tǁXB��.ڷhV���W}�9hC�e��+��2�-�� ��LPy��¼U+ \\9�����wgn��������e�\��1��Kg�,���P�v:�a�w�/��QR�@��k�����
�op�u�Z��#.a��5�F���d'�����ox���!g*T��L��#���؀wm	Bi�V����ux���bm+���4�KD׫�L.�u`�<�+d%1hw^�D'����|�0^�"������~�������y��,�Lc8�I�H���π��UA�PaK�����\խ�k4��t�����
�b�M{r�ez�#9���T���"pX)���A?��a���b�e>��u���ڜ�v�����a�kN{+o�y��>u�˸�5�ӵ=���Nˮ��(]:���P����Q vT�����Z���(��Q�� 󬙗�Y%[��:S���ÿݗ5���!�?XR��G��>�����?Cu˫j����u�ْ��3�Qe��k,|��v�* ��L�e�F�Q �����]��� |"�'ʳy��JY�蝓"��2t��ÑN�|�I/pCA���)�~��t��������W�/���Y��51D2���m�MIWv`n�2�y�E���U�iB���r��j�)-"�H޻b1!Gx�WuEG/��6c�%<u���[��j�Ν�u����]�̵�7Ɉ���h���}�N�y{Vȗ��!Kc42 �O�����fb��#��1�/ۮ-�<]��hn����Gqo8�@����C�1�\Y�u���vW�VB�=��psA�퀳XH��&�(gq�%G�gvP�M��^��W��T���c��n*��������?�#������(�4j��b����>t+��dK?R]>o�Cwt�1����L<��cI #�A�r��Fj�LU�yۡ{�����㣽7L�i?�Dհ2%B6������/BBS���br\~Ē���sdP|�ߐ��ﱦ#^BU�#�����cj�,eD?�V�s�]�B��~:�N`�-n�_������%=���'�Ĉ�=,�tgK��@c�L.`y���HR�ĸwDzӏ��"J'�oR��˓�B{�C������෨Ԥ8������"�2��Vk�W�:�A�g6ikE���ڋ��<چ�+ٴ��S��+\N�0%M��{�a��	Z1-���$���q	�?��<��1��u;p�Y��FA�ka��+�Y�Fi�ؤ���QxYH=U�!�dH<"i����E6����^�R{��h�؅�!�T\���ߛ����,�Ȗ��O��T����Ք�댮�1�*���R.�V9*�!Om�}M��ٮj�CG^�A �^���6�U%�y�,߇#�p��'ow�=���nW.���7SdPP�ք����e��s���ec��X���w�*��(:xc��쥷'�Z��m�8r�+)w8���8�IUUugu��qK�m�o�N�1���z5�)'R�����ڝ��B|���o<ؚ3/)�X-]G;��'��b��ƭO�|�����靔l㎺2bg�{�0�(�5�� 	�d+	������f�s�:��͟�A9�/�c��IL�<x��E���oO��t8�H��'l/i�v��>�\S����!�G�k�0�H|r	�|�k8T 1�z�,��>�g*p�e$`_�#��G�#q�v�h��V�(����L�Mm
Nu|��-�qQ䱒��_���͆�Px�����_���JX�&�)o,K������z�Iފ�x��
�
��%D�&��Xif�L�i��!��%5A����J�Re�|kx�2�T�c��~B��k�#:�����ۏ�7�V�@G�����л��O84i�",��l7�R�J���(���T��ì�593{��vo)�7��B�Y���s2-�le����0&ˑVK���AK 06���ڔ�'\0e�[K����g�A�t�&�A��!�9ù-˳�Ss�
[�X��]��M$��c�b�]����'���Jq�b�����^/����A��R�w���<ǉ��O�w�\��>�������� ���`X~I5s�K_�wӡ3Ar��}�*�jT+�B��$_�b`�r����D沉ݙæ�t236П�%ɫFlۨ9�	�����S<���ҽ��QY����%��T?L�]R"�~�Ѩ�>֮���(:����[� $]�&[PB��%����f,Mp�NN�a� �Դ��&��e!��'�Gk�6(��,��:���4沕}�����0}݃���`�ίC��B��Ƴw�Ŝ��L�cE����o�R7@n1iy��N�m�R�`9@Q�yK�gT��?���r�|fq���=zģ̑��^J�-�o0�V+�S�{�r>��?RS�����Xڣ��)�`"盛��F/jD�`�筨nA��/���Q��=r�ȭn����\��u$�E�McPJ/��R��L��Q�iU�%h�;�TLtfpl|*��
t��1_�2��h���.�Q*D�3���֨�qף����f��:��~{�cK܀M��=K-��L5�s������ �,{i�ԃV�vk����D���N���PP�9p�ZeI�g,A�h���g�vı^)a���	Y�q�cZ	���q������,Ә=�͵
�����D�{K\�C�Ǉ�ŝu�ƦloV��1�]o��
�:E�_[{&��R�4�J>�gK]L�2� ��;��d4s䎳��H�E>pu�¡��K�� ���7^&a���*���e�(To-ԭ5�z���=?nE�e^��/3\-��N��t�%v���➓&P�f8�V��,j()f���;öu���p4j�2�˼�QkԞ���OJ����l�Y�z�FM�@���i�'���Ek&S�s�6��7����7 sN��N{��\��9w�J�˼Hu��.x]��@C`�ٔU~�kV}�o�9h��r;����]J�D݄~���\������rh��#2��Y���:b�5;�����G������r�g'~�*�Qܞߩ�[4 JܼQr�y�B�m�P�LA;�=�=���d~��%�ϩ��6�A�;�#�4c��Wl��X�͏�. �%)�R �{��wG��l.���>�[�+=8��<�����&7���F�C-]�FST�f�%�lO�k���U���ڦM4Ўc�	�h���wl�( �����zg�޺?�OQ���3�����l�0�bD3�%��I���Ǚ��^�Ȇ�Z�c�hF=(c��\�D��JNu6��9�`5��/fo��2C��@V�GwA��$�,d~�/
p՘�Բ��Wum�&L��`N�q?�)���b�޳������X�L���d����SR��خa0U��3Ĥ��*a\�?f��D��k�n��v��������
CiIv�mx���2��$�G�õCl��Z*�Sϑ�sxH�S2�Bt<k˳��U�>��{(�E��c�t�e䮅�y��I�����9��/�-7�+t>}�|�jn�N���rA�����5�O�8���$����݉:������+��L�V���Ηބ�H�ui���j�8b������l����[ZCH�^�(��-�d�2I����Z9���� n/2��V���N K�%_�\���<s�3�kQ�g�V�_��:Bh?h%7�h���2�F;%����Y��x�u�t/s|�R�"��}?�2�X���BB����j�|z,��HD���h�����͒�T�3�	�#=���XN�ɧ8Lr�9J+"��5"�4{�ۻ�Fw<���ڂ�;���#}B�����G<1E���X�co^���<9�2�!���?���P�b.ƽaTs�	� �c�3	�|j��!����e+&x�
�}���`:eV��BL3p����?_ �������@|
��D��������~Y!�S�?n;�{j��q*J����LQ�N������fl���!� 0<���!���<b����Zţu^�R��Jw�tҘg\JDLݜ�7s��oю�~p�?��V^��"pUҌ�_ۓ�T��X��� �(�57z��)�o���xkk���5| ��Ǿ��jm��|S��8�JtA?W6�Qv���RL���-��v4����&pn�47�Q5�|kvJ�a�J��M��Y�����ٍ㤮]J���4�����)�ގ�&�:X3��v#p3���z�K���:���;�>"��I�y{gצ3 @=���~;�\<�t����<���� �~���x��φ3R�tvQ��m��k4�l�	*��p�
(�q~ݢ8{�2�~w�M
L��48Q��A˂?���z%m~�L6���[Im��F������2�����f�[�7��k01��s���#��xʚ{�uJ�0��hƐ��n�Z��NL�~�Z�7H�$����Ԁϥ�+=��M�y8(�"�8�1��8K�g|���9T�Ε4�0o��`}���-Tݮ��F�H8s�"r�2��'!8�w$�����w��&>�& �If��xkz��i�@�.g�:&�26����`0�X/���uم���ةK���`M�r�O*,�,�qhm�H	:<�R{�#4Ň݁:���DT���K�D}��)M1E�&��-�A�*�{����Ϲ���!a���j���'ܡ��n}���]�#�1�G�!vS�yA#�f���
����~>�R6���J��ig���.�Mut��q��������u��B�v��X��߸T������8�O�iO�r{��$Cżbp��v�ެ8���^7����Mz8��K��5��/��0s�$�|B�YW1�	*
��4��%X����
 �������{Y� �[�<�8!m�U�k3I.��`�C�l�Hn�v���]��v�c�������6�!�g�O1m~,�������t�6�G�T�sd�F8�={�*A���E{^/U��]\�Y�.�׺O����[�m1�!�v�W/2ɝ�vYr�(D�a��}��:nL��B`n	���1�}{�ls�	Δ_�ԁZ����h�:��닠�3%F���S� 8b�тD��`�eZ����.?�jH����%e<E�=��R��+���EĠ��w+�7�V_�Ə�ǜ��l����\���I�wr<	�Y��u`3j7@İ�ǑSL�w����N����ה���gPv��Th���	���=Q���	w�����nC8Z����5L��K�~3B�ߙ,�6��Oh ��lcK��m��6[�a���� #���C�,����3����K�JZ*x���O;%��?B����ɠs�(�f�ì	/xt��l��e�z�^�	sw��ę�ƀ�pn��r��CSLqFT��&�z�d� 2���)�$;怺�'���$؇����ԣƇ┪�t��)J�xM����N�I"6٦�A����H�"6C����Lm��9��F�D�:_4O�bx�Vq��XДbH� 8���f���X���	2�~RF:ǳ`�^x���r���d��	�adM���u�&��I��eg�}�[Њ!�A�B�]��V�7��1J���`ȯ��HD茮���>�sߞ���*��a�%�zu�T�m�����u���ΟCD��tJ�M�
2��,c�GB6O�y���	v���i��E��/��ۙ��oEsξ�@�VG�P��l579{��r�٦,�yM:XR��sA[?I�Ӎ���H���)�p�M��I� ��y[���`�u�蕛���-�a��6�+t�V����<xf?�cC+�!/�:v0�(��6�I��O^&%^��*��Q�Lǯ��i������VX�g-�}RK<SF��}M�_�Ӌ��c8�i��q���`�R��Rt�UU~b�q�h�5��r�{���l`���,H�tӼޚ~��#���"(>@�����"#ĉ��k�LG6O�e�b}�;I)DH��T��U�姇�R�����!��}��!�J���Pgؓ�"���1����1#�r�-I���1M�Pd@�p"]S��1�D �Ͱ*���z�������{��2�|�^���ZA�Z�������i�צu���o>P����{�B�Q�����0�va�����٦R���O�#U"��y��Q�O۟�Bj���"�_�E	��I�A�#�����c&��N��lc��W�d��×��
ψ�
):�pz^o;�o"kL�,W>kĊm��MFi�#>�M�*B:�`�<�6��5ɀ0���jp��5{Y�-���̓R�n���c�O�D�W�cf6��?�p7A
0T彰��r7&�6+�d�B&Q��=�NF�2P~ڽ7�@[��V��g��d2���[2�6'j�@[=!����׸���1'Ҕ3���W�Ax���
��;�#�]�d�ք3&�	��o0E9��D {#(��\�CA�;��w��M�����,ʑ
{Ux����p���S�5��J��"E&�� Z5�5AKWW�5<*��n3۞,&��,\k5f$�o�Bus�{\�~�bXJ�jѢ���;<�p�%�8��{U\G��R�vjq%>n���Ҥ��/ۢgG�ŋ��7�������S���L����-�Q���wv���}���W�8���9�E�^�O��3ַM�X{I"c���;��ǌ��y� �L��������nS4��5=�	�Tb@8C�����Ʉ{��fnoNҢx,e7�KQ�&Ep�h��y�둎k�N�ս�R����܂K�C/��K�yKEפq��m,��͢�#�8�b"��<��O}�@��u Z��S�nF�iW�	� w��@\���؃Q}�l��gй����r1����)�?!��i^=����^�[! p��x��F$��*��p ǠҼt�!v�bjlv;�H�+��<H�vy��h�������!;o(L��I���#+2�y%|,������*�B9T��ܹ��d m��57
h��@A�ԍ�5�ؤ�gGq!u�� =�r���1od׉��,�wˇ�}���%�i��vw^��x+��DFC<Cܢl`y�EU�B(v�������b����WfM����=k�Lc.��71�{$��؀5ʩ�bxkjL�d�z��қ�7�o>Uv��V>��!�g��ZiI��yu�^.�Xq�<6�}���!��AS���O�Qd8�t��s�v�0c�3���y�2~aXP���r�f�D1���W.�bj[�����J�W�:�����_!Oj������ �
���^��>e�4@s�f��H]�>��S�߬��3���������9N��ky�)��� � Z�P���AFP�Ӕ(k�	��8oC����0��۲E<����,ȻKR�v��ނ�z1�w)g̟���j�A�H.������t�8p I7Q���J+j�����<�:T��턦;�Du�@�K���!�P����o���|K����2�3���5x�>+��=�C��P��N�K?�%�
#�Bv��R����ɺ'y���5f�6�0����q�Q��]�Q�h� �*���H��T��"Q��X�2�p�3��/x܏�P��	RlI�ȴ�YI�3d}��P>[��g��*���T!.�A	jC�1�L�[�����ˊ�q:Е��J��_��~���i�;�W�5������P�㈳^JbYg
�8{�$�O���w=K��F.�;���t6�������*U���3R%� e��ʚ]m���=�<��F�<�&ȇ�M|�4�\I4p��E��9���92Y���~��uP�Ua�)h�>Se��w�!�yb.C��`7������
D��/f�t�k�ѝ�z%[�]�؝w�A
���Q�d$Ќ-�{���` ;8BQi�	-dg������ABʂ�z�V���w�"L|��-q�l�S��)4�x]�U����ư�%�)KRDG�[�b��!�%�&���S!�;��vư�E���E~�/m�� �Rd_�6.�U�X�Ɩ��>��cS�2ǧ�eas����ʄ�_��ze���W�5!� ^�bZ�G�ui3��~�M�����.��A&�(a�ܶ�'}���+9w���.�&���噺?K뺌�d��_�F�_�G�|����ro�v6�8�}����cx��À���������Ԧ�x|�4��0�7�$��"��S�ϾP�%�J�^�������3'r`k�>�(L���_�}�/��} H}��eD����w�+� �*�2��Ԝ��<���kgӶ,�k���r�%���W�ߪ�����R���Ե����GK�h��aP)ۍ��T���_iXU�Se�D���2�����\�g�ɀ�7��-�Z������7�sV��5�n}�Gp��������3B���%�if��Rs�.�i���k�)�j2�:�W�_z��@jʤ��m>&��V2Ͽ�h�w�Y�ҙ�"���nd�z����_o���'���{��S��(�ۛ8H��2�XM�����xQ��0.\��OV��|e������`�e��g��B�go?_q):�@=߈��9�6���N_��>�;�wc>��xD�������yd����U|I8;��ќ��gm�:����_R�ɲcw0ݪ\SD�P������@e��C�]3Ŭ�T?�ǎ�+�|}yg;m
M�r3�&`�_�t�m�W�ֆ��i1�KQ��(�mDTL�0��Z�@�x��8oE1�XcS/��q
_8���SCl-��i���9΀��(��k�����c�{��ژ,p��m��s*�pxEv�vI�^<R����v�Y+��w����(#�����[KAC�B�H�J��H�X�1u�*#1�� ,Z�\��М�r�1�N ��x�oU{tgu� ������#��oW�%R��\�ou�c���Yn_R�	��$�׋M����vݑp�$��O���T��s1=$�|ǰ�@Ǡ�u}��T9�ܖ>a�r!�lO�B:�\���no/^�x��]�>�[������ҫ�t�wơ�|��K�B����נ�	���쭂�$�ͷ2�Q�Cw�z�6K:�0z�5$��9�;�،���J��˘�� %[%d�Ez^�NWo������w� PK�|{'��K"�4�<�0�Xs�k��u�H��
;��V	'��~�k_�V�;0��[!��#a��ؚ��2cjL��ᡃcBqĈ3���'�%"�G�[x������ܠ�N% >�\���[��1�&��](\���e��#	�tSxC3Y�f�e�
�b
�`J{P������x�0�w|l�L��Ul���6�_҇�R��aܧ	����n̸��C����2�+�Oh�ĳ�m[.�����S=���R1.�Z�ryW�Ǒϫ@���B���v�So~Yz����꒣���TB���;�h]�'2�e���p�iW�糔+1�læK����Tv�<���,��VN|�����c[��U���;���E�:�8�F0�Aࢨl˯SD��0�	S�6��s��J����g��:ޕ�ޔ_�*^U.���8�+%�ØU(��k�Y�� �1w��c����\L�X�ϐ����V7-�uȟ�)�Ҹ�x��J��=Vf���,�`����� Wd޶����I[AXF+����gi��ɖy����ؔ��FNB�_G����(>B,2jT�����≍}�r�_��~a_HYҭ���GHc���9�wӻ�gS�-�ls�ȸ�Z�o����T����h���]�-��.J0��b��/��?���?A-uܰôe��%'9IW
K?N����L��q����n�+�O��1_A7�"�QՌ��J��
�\����B��-������ߟۉ�������|cp�kv�	<ي*��)����!s����*��f�i[�j��j_�*fRp�Wo��	���7ys�m�)��v�` Zɔ�]k:�{<jbB�Yp�|���&-A1`f�� Du�%;�����>f��Ɇh�KR�țR^�REDy��i߃[��~^-�o�җ��@^�:H�@W>_--�q�Qb�r+ȅ�6�~��ob�yJ��M&�7B�~5���D��3Z,�p�Z8�@5���&^h���e�.��	}5EI�]7Ή;A�f*�� ��D��\��=m޽ƴM����d̟���J�<����M�v@�2�-��"�e���tׇ����w��y���Y�΃���*t �ذց���<R�����i�,�����w����ԍ�)񮹩3�
zH^H�mF[�v��2R��!�E=�� \��]38�|�;�N}M)�Ί��5�W&M�9��V���]X�ef�ӭ����帓hEHա�z�:<ฅT���(R�W��x�'�~
P�B�
t�6P��N����
rF��d�x�-^�)�<�-ᆸ�L��ǶM�u��{���!uF�D��q\��	�S*WqQ@��4���������T�6A�?�pB�Sp5[%HT�v���6(�#�@�l��_���v���+��-���3�$��XE�[G}��#��qIl�
�N�Ɂ!�K�|a,%H�M��tyϞ��=���^>`7f���+�q�I�uGn�=��A�,2ܭ$��Rd�[���x���T�%��Ug�/rH�?�H㟄|r~(�a���֫��NpC�"7�����s�L:ڻd�4iG$3
���< 
��6Kw���Q�璊�'�~8�����������E�vN�'���?�Yt�wMG~��(�V�H��2�-%�h]Ϫ�=Au�P��O���.��ඹo##���U��D�R/*�n�8������,��"|D���n|S���ubP(���rX�|^�^I:��8w�^~S��� �V y�� $��n�w��G�������&l�/3��۝�j:|g�г��l��ӔGK��yα�V���'�'�yV0pt�8v��׻���rJ,Ŕls��ڍn@��a�����Ӟ�Uh����	�2:i�=��c&�Zi��,Ѫ��/��#G�G���a%��H5���e�"�� '�7k��R�Li09���C�3gdbRmpy�E�c����h9m���^j{�B���ßm(���)�lT�����r?�VeOR6E)q��*�À3�A�0�}{��xO*uϹ��D�f�6�EH9r�U�G��g5�n�Y���9��}�L��I��B��bẒ�,_i�Ճ�D� j��z�ō!2i6��ʇzc�E��2b/�LM�7��TǾ�����)�k��F�.����9�u�[:剼���}��):K���ISٻ�ӫH_��&;n;�64X��wڋ6٫Jp�R�t�E5�i5�%���A�X0b�4KG���$9!d�t]+ק��l�z舂����� �i�k��Ep<67ε�hQ�\dk
3�L��[�^5�l�ӷ�b��wQq���i׼�ŭ���#����)ذo���r���E�/�����S\��G�k�|xe:�i�n�I�2d>黎��I�l�{��ü������������h>r��"�#�PYb;/	�?t��+��{󍡋��3t2�i��!�qWp�JW���T�E4�E�e�[�]�L~�����V�o�N��P�m(��.�fi�@ç��U�R����|�d��+{d��	�bq�{>ΦQ�v�S����%�� q����ϝ<�*$���K�#1&��
'Yg[v�Ò���\W�Cg��D��餱��$��	n�!�X�P ���������Dٹ^�7i)���6,Ht�Mc�u'<�A�|Ft�� �k�_�Mr�;��d����A+�YЛ��$�HM}���P�`���X��{ %nI�&�e���4�$bE誕�C"F�5Q��υ?7�2����������E8�N�k@aQ���ysZco��q�kU}��/�8���;�۴ظ���b��:&�@f���w��8�.���m���A�sD%�-[ UsE%lg���Z�}C�ϓ�#mFǘ�;{Ƞ�v�I�2��3�䇲�Z�R�������t�n�~�4�o8����.VW�=`�ߏ�y�M�A�N슂��Ϛ#э��3O�M6��O�]�/f�t�u���"{ω}ҧ���iL/�.�t���K�3���/���h;|���sG�&D��O�B�,=��ۚ�cJ�5f�(�,�k�f�X=g�3w�H|�H)?�M�9��f���� 4�wmv�e�i�:IK-R�i@ƴ��0Rn��v�ǘ-DK����T"e!�K����n���<H��+	a#�<W��F`_`���7�Ok���p:��v�VO5"�|��VP�6{�'L��!��S��K}��	�NmY�G���2�ux$T�,Z��
k �om
��ݢ������܅���U��M���O8����E��u�^_Y�hoNcL)�7�E��ڹ�s�Xh%2���g�n��L0Ԭk��K4YJvf��= ��At]�\Ǜχ���)*�� �K�D�3%ŧ?Ұ;����=@�>�6&b����́S�9\�f��~B�͵{-�v��Ը���s^q<!%9��|��\7���"������VC����ΟƲL臓AK�֕��_e�1���_/�]9���M�B�Z��������I�rl���X�����|#w�_�8�H,�r8v�����ߺ�C����Ne�yK��(�z�E���l쏃�;�(pW��*�y=~ܭ�������i�PU�}h���YN��~�DI�Y��!����8��`�\Εڹ�@�r	�iծ-˽���0�5���6^�������s?��L�Ofd��� M�E��/��.�i�r���@(j��
�6����<�`�/�|7�ưX��-��v�-��)hV��������~�K"0�	��7�1����iO4��&Ra6k�3l��VeO�\ay�/(νLl��MԻۚl�Zjp�YK��[��r&��C���4 �їQ�IFXs�C;��ˢ�U�����<��'���J�*h_�}�V����\��MK��E�S�Y�̜�^�{��7y����B��K9�®��t����=aR�x�l�˖�ׅ2�?k�����>���6�B�$S�|Ӝ�S��~*ha2oTq���ܟpd~��H���;ґ�W;�V���0 �����9&�=�yk��/>���H��0Sz�vH)8Y�z���#ȫ㩓�ӽ3�ƥ�$�����@��+�b� ��ro�v,�.��8X�+��!ig<�K�M��cR�=2q���|?{���1d���\{�L��'�p4L�I�5R��XՓDO���Ŵ�?$��uF+�'�k��YS�/� sJʆ��f���eM���IE��|���EHqj�� 
�Ĩ�i�Ҫ��顠ڤ�17����H4�f%�d�V�z_2/�p���INe��=)jtx���F~1Y[S=��� `��	.o�D��+�׿��×2�?�\$�is��A��ucC��v"�\~�y�P�����kЍ=aӞ�*���ùz�<�Ԭ!n�l�t���1���P�O�,[��8���8���!b蚮�XIH���i�.��36�e�q6�q.色)�,F���s�I��,�%FP�_�t!݅�w|k-E�`*\�y�Z�3=�r�M��e��>���$����|nl�V9���{6!5���澼��$Ҷz4�M���ha���d�var�����wۀ��]_(�}���l�#�~�*�U�R���)Ye��:v��]@�s8i����W�cj�X�HH� �A@���KC�κ��Z����l���T|7G�s�����("�F�����
7]T"�kU���бW���:}���p���8���;>:cص��E���7�xH�FJ��b�W���!�Gc^���W�F*z	�_������_OY����a���6R�VM�3���ȂMT(�b�R�$�����zb�#����KFAӮ���{���0sc��q�y�"F��zK�,�zN�ĊM|l:����+�x��������Ϲ�\"��#-J6;f]������cz|����#쁓6z]a$� �����db���$�Ly��*%܂�,ˣ�!%̮I*VB�%B9��-�~DM�Y�`�9ߐ$�:�����E�XFl5�爀k�d�@�r܊|�~��Aiucy�,u��·�픦���qw UXg{���q.�)�6dd�6��h�ũ�u]�~�	����*j}y�qQ���� �G#�����+� ��M_2��v�N�PVD_��:�X�o����ԠQ���y������?��V�f�7��ѝZ����	��n���<b1�ݹ&)��7OW�q�ñ�W.z6o$p�^��rX�Ha�U3������v��L�
w��L�l��A�ȻE3��"��㛯���}IUψ��J�7���g���U]��0o@#(��A�+�'�!�`&�7���y$��;�����5����-���i�)-�g���z�Q���/ϓ!��/lf�Ӽ�v���-k�?~{8���*ٓ�$ɏw�\YnO�8Ƅ�0��E���;Mɼ6��4�z������k�EJ"�c�|�O�#+^��V'�"_Q4�ؤ�ҝ��S�@��lr7�:�@��K����,Ĕi��f�]i_7��4L�%[����3s��8���(Wʣ��僮�h�����T��f���S�g��I��}�q��4� ۩D�!/=��-�+����׈q��rC
�f<�*:-G1&�=<8�� ���pE��(��9�V��[vTg`�:0����k�MNH^è�T�7�#/2\o\F�R(�[�}�U��[ұ?��
�{8��tˌ���/��헓s��yay��`����L��������.`+n�En��1V��5�M�����m�Tҙ��M ���۲�[�Xʵ���(�v��ﵖ\�I����p*��,j��1dB��t�5�(�����+4޹��P<b�I)lV�����>N��0�����$�Z��~8��[�y)�Heɘ��9��S�֞��<�S��S��Yd�Z��;H��m�݋��'w�x�֗ч3h
%Xɡ68Ǹ�<W�@�a_�ܵ�����#�a��qJ=�Z~o�H�R
�q-�a��/�u�m}z&nz�Oq�]v�=�W8K��s,B���_��v^	\����p��lҢ���>�MR���@E*�������Ք�h��1�AL]�[�1&y�]�:ifV�\0��\��_D�Ԝg��Z��#^�ݯe[���F4��n��mep_�o<�~|�Ϛ��!��(���[�"�}�Fz�T"_-��t�i£�ϡB�U��¿!�6�{�J!��' A��������HHc�
���9�R3��ZQD��oؒ��%�%�nmA��|�h;re�ſ�bl3B<I��e�)V�\k�}�������/y����t$�ŕ�a��W�M���/�����v�L�W�Rk;��%�v����-�|/��IcD�H�e$�����a�|Ä��1��9�9���{�r\g�2�[Nt�T��[��	SLAGt~�~�IGR�����UJ���A7@�P��P�}:rJJeY.���A�9=ޱ��mF��f��&��'/�6�Ω��l�i��\b�K�g���͢�]�Q	b��i�R4�@�������8����>�V�M���\�n=����.�~��۱��!�;�\���\��œ�̞��h��'�V�p� m~2,ʄcZ�]GX�`k+���������ۨ鑯4�A�~�.Z���E�KhW��P���b\��l�I/��E�C�K���Tq�j�!;/x�o�a�+\��L�]0����}��݁���Nƻ��{!W�	v�a���n�d;bsD����EFa��֊c뢻�Ф�Po)���Q�?��8D@���hI�T�$5��H�T}���x8$�U�+@�w&W%���:��i�&.���yEn��}j[N���FHyU�F��ы��^�������q�?���U�e��ک�*FR�@���1��4a��-k9ƱQ�݅��
 $�V���"I
F��u>j��{l�`�@��~���Ib�'q��@��`F1��H��<�H=��߽W$�S��_l��Dy���\`�䘛&a��N�U�ޑ�����Ɛ��3�r�$�BY�GțV�q7"b²Z,_�=��h�Љ��!U�8��t��)>��}��2ͨ���;��W��W�5�i^�����2ʎ4�>�v�8��g���9�Fq�n�l�i�2#��S�A_p
��|������?��v�4���`�	{�<��¡;����]@ݤhx ���͒b��Y)1�j����!�Y�$pk��D�?Lj��^5R�����	��Q`c����jr�%�q�vEa���Ƽy�r=�y�D����&�-Z�2?�b[�|�U?4䢮Z�9I���Ne�}� K�u>���iHB��%�e�ha��w5�����n�w0*=�0>R.܀郱�ȹ�8ȣi.������gb"-�^�I%���F�O���/���─߯��Gr��3@���YH6݇��'Ԯ;n������Q���.K����!�����m;��D�ԈᩕN��G�
�h�6��@��D�������\�E�u����_F�A�_
��EZ1�	͆I��߃)���փe}��0vk����
�\Ĵ$�7�0��]���Oy���ڸ��(�"W�!�3jgS&,m�2�����h��/rj(�wR���Bqp��������	H��dK/Y���=�/�?��.ٯ�
���^6�aO6o<, \��:��`<�<�(�خ}6��\s��Qr�X��� ��D�>M�p�F^�yM)�n��n�l}�@�A_�2��,j��1������,in�Č*�1)I �c��d����Ǿ��;>n��|�M�i��Ӫ�i�����޴D��ݲ�!�qp�)��Ey17�+u�c)d0H
i��T��������6�����~6>����'jV���BOi���J��c��9+[EKa���! V�o:/:EÃE��*Z���Pmx!S���N��I%�i��S�i(��9��D��zǩ�7/�e���6�������%��6��1�e�A�|��hDr� \�������\�=0'��jI�w�t�<woca��A`+5�C��/�Z�J<�1!X(݁�"�����T6:w�V�	P�H�
��(��S0Ҋ���L���sf/q��m{�nmP���Gj�=y|�*�x}m aB��uF��� Å���RrW~H�گ|�B_l4w����`$��E�����7Mb�3q�p#TB�D�����pڵ�
��kD�=��)�&�1i|N� �|��X1��ז�­�%\$�TN�q��������|:�_V�����a��]����F�Q��;�c2B�;�'$��R´�Y>趡 V���bV���x�tY'T��d#��7X�U�J��lM-���}6o:l�T	??�.��8�a�uү��N'�/�	/�c�Bb�p�w�t���M
�Y<KO$)�h�H�V�L*�����Q穳~�(�Lź��7>����iǘ��Kο��������!,f���	��cV�x����m0-'�B�L�
�h���F=~�>e6}���������/ĝ	�p�-�
�F��U
M(W���E=D�����2����6�]ZZi�b���M����\���ū�MiI�{-�����Q��[�3�s��@���|��3�Ɖ�ɴ��xe,�]��BI_�!}H�����ú�ҼC�pm��Uy>��?q�d���JI�ޭ�KU-���n�p�-dt0n���F��&�3����"B��Pv��q&�W��$�]~%a��T���Ɂ����q�63��h��(�°��0$�Y�PޢDKq�L>ۂ~�5r��||VR�W�����a����c��\)���ͱ���u����u̒,�0�\+<@���sq;�x/���Xw�?�Zͪ���=>ʎy�#�(��x��|��Z�����83���6A�����m��;������M�f�n�(�]��>��$��џLV�T��m�?NA�T���#ȏ�5rqu@����YB�wN�GسL<�,��D 9�t�Ī��C(�
��f8H��֥:d��)3�S��0�A#�H��w����9��@T��0�c�{M�����S�b6�����a��'���3��Wm���g���C(�n��z"՟Ī�}w[L�Ac�0�@�:��,�(ӟJa|��K��\���Ei�SC�Չ|@)���OBdcdVx�f�Kf���X��.,meˣh0UUv��1�^Ǥ�
���jK�+'�&�/���\��vl���O��q��
����N�+u�F:�����yh�o�<w>���~t�V�
POG�N$x�sg����ԣ���qI���Z�|�ء�:�@�Ϗ�l+Rz�s�NK��!8~0�<e�&��pG����WQ�0�!��`Q����u_ ö��$�9E��f��-'ԋލ��Z� �htB4����i�X�c����p,��(p��^
g��U�U����f�d��|N������)g��-��
`;�&e��}�`�!�-���nf�LGN�<�xYi�L%\!�%�Ą�Ax��M�z*~ґ� �5sr�N����d��� ��?3�A���0	r4��|�P=���"�N�֓k4/��0U.s_�Dm�� =�C�����͕���.�\F8�QB����@����Qt��Z�պ5�{�T�U���?�8�7䑊��QL��g�u%c)D.�j��!�oJ5.꤀]�t\O,�W/K�DNO:i�~��jz����P��[�R-���I��'��	&(�0�X !?a#H����g.k` V���%q)`#�g�
uo����ǇL��h8:��I�]���� 2�F:E9�m�tI 4��H� �˚␋�hK2��3�u�Y�Q/�}����1|�|ns+}O���{����U���|�t�huS6��/ALJg�燉����m%��4�A+�#�/�o쇨[Hq�X�_y�J����q-�L��"(�|�ѩ'�G��7��ȑ3,ɢܑ������$\m��gT%�p%�{�f�����:�<o�lq��ۗ_�a E�l�R��(�5��M�'����ķ_M��rOg��-7&n��!b�n1�9.3�%�[����Z
�9�.�F���T�ar�bt�b.>`J�ɵ]�_�zbJ�Ũl�;��=�MJf��=${��9��mUR?s�5�-�����Ψ>m����U9��B��H�L.y��l�p�?K���q�I����M���|��P�H�e���H�����:�����o���x�z���M��̸�Y|�X�q7Q��e@,	�V{�P�8=;&����opT���
,vu&���'�N+<�\�����~Jk�)��]-�
s��Qxu,з54�G*�p>Hy�,:�4�oGȐ��S�2P}�`௡�6�v�q&>}`�3�D�Fi\~NA�+�]�\�����べ�,~+xt1����q�'�w?�3N�λ%�)�m�:�`Rtd�>��1;�I�:k�/�:��˼�3�p�5��%�t A<�	��fFt�Ml�['m�}x~c?�WEWs(�w}<�ܲ!Wm�T�1t0���!Y�4|��
z��*xM�z6����N�V�Q���UdhP�. u�C<�Up����|�\U�vZ}Ɯz��A��b��gI��Eu���X�nP�ӆ�R��G`�䭦H iҠr	ͣK$<m����6F~6�?�"1��E(������dE�!�n/�eH;�=R��%E�@4�K@ш1wp��&��P<I�A��P<�G`V��4܎���a���5�FWT8=�Fi'M��X�Py��]�	���/��~���լ���B�����h$�a^DU��UΞ�m�8-ݿ���B6k\�|�~!Q�]����P.dC���9���������l&}�l������ߢ���t���j�C�������:���� ��]b��ЖoS;�ŷ���P��z/7�����~�7K� D���@>!SKe��U&�_�#܊�p$J�A�ׁL��.�@P�PK�3�.�;��I�s͎����o[�!K)��ŝ�h��ӵ�s���_ � ���x�\*1y/�K`Ο|�7���	�%趼����>c\-�N��N�:n0/��ԟ2R�+�wʐ#�K��DP==QhT����=���G�(f�D����<ç�mh�zHqU��<��wpsh�)���ߺ_ƥ0qׇTg~�h��v��m
	Δ^?�L��s�m8�J mD�����y�3pJ�~�����fO1����#M�s��%��xާA+U�.��\|v��Z�� ��j��ج��Or?�ɖY�$�!X��?�4'��w��1�&dk�S�k�����rJ��)����9s%��+�j�B�����Qq�Κ�V(�N����P�����ꅝ�����GL(��%3w�w&�x ϴ��Rm P�p%�;F�\*;��
�qW%��%�`9�;���zq�و�ɝ�akZ�����O�)�Xh&�i�g��!��3�$��hW�"ThI#(��&J�P�t_f#��?����&�0߯� �`�d�#����w�[#�Y,U�<a��>��mD=�AP��K�e�����4��W�V�g��jB"���4����ЁӠ�=����jG�����D�&� �&U�_}���t3�H��ʯ4��&�i���b��U2s�u<���-|��d2`R�g"�S)��87m����Ry�;��ԟW� ��L��i6�B����+�Uld;身����&hJ�Hʩ
��=Jd�j���b:|�<����_9���¿�a�렐,H<&cN������A��;�L8���2-R	 �y��̿1�>���N�C�eg��>��@FfѠ�J!�&�F��3�@�B�M����׉��W�Q�/T6|�[��7g��Mz ���GЩ�]З^5�.ZJU�Y�͐�AN6���]��U[@��\!�n�yQ����]#;\��i�����2��Q�/��d���
[��-P*G�ٷ(�lv����N4�*���Q���m�{�+�n5��b�)�(qv�V8�0v��l������( �̯����+�.+p�{O��3�MK@�ݑm����D.w)�^?V+���;�i)z�I޳�9�:E��2lW`+Q�/	»h�:H��=�ADܶq�y=4��_U'#��%(��$H��܇�"��|Q��gɋ�Sn���-W���%F�ٷfhiH�}J��p�Гi�u��{\��]�窣�/C����7��S��Xc;m���Bԣ�/F¦�O1��!�񋶒<�����.ܫ�^u��rf�~�?���K�Z��H�|�����rĸ$�ʦ���lf��%	��D�v���s���g0p�m����E:P.1��;+D����2B�"�P�.��!yktZ~��9�w)Ct���1^��a����(���r�a@�6ns��~��/<��Q��O�n�"��;Mf�@GRW��NyШfBE�0ǫgYy20!�Io�s�d�1,�������"��V�J�7r��]J�8�pJ��/���J]�:��cu/�nek��J�x^��}�� ��"P1��ȴ�/VWU�B*�ޥ����h ��� ���p����캽F@S��-��oJ3&� �<z�\�+�C.��,o��K�Ż��=�,�H�K*�٤���[v�e�޷�ەUe\��~��\���'a�;��kq���>��+0C��j�����gW	YELT7ozZЂǎ;BS�M@4fC%�B�+X�Az��9bYI�x$.�F�Ȳ�.l�˼�0�+ER2�u Oֺ��z���� �)5�<���</�0U/������Ez��<���P��#�� �:\Ns����S�j����kIa
�ߧ:�%����j����rL�4�H�~y�e=���M�;�Σ{�˙���߇h-����y���g���AcQ)M3�:���	Lq&y�����5�P`�4��t�Z��_�}`��ur)4+a�9 �]r�!���u��b�;	�$Ux`��I�����C�b�36���C̮1�)?�P|Ͻ�=�ܳ���,� [f=E�"��c��J��'J�/��E�Eqn��|�믨x
�m�]Dˠ^�Z�X� e� �a�I��l�ƻ�+�
o�>q��Yx�|���k(�y/ha�@�|�mg^mɜꒃ]�Q"�Y{�<
�6ŋ���r�YO���{�����R0��f�m"�&��X��5Ǖd��7Xza���􅟠H���<5�I1c(C@g0��� $��Y�9^,5���H����a��0�.bAO�'	�L���aB(}d�RMJ}al��gM��Kf�mФ�|�����}<Y+��P>�C:?�nb�w���\��Mi;�0*�D^	�E9m<����'5]ucJD!b�9����I���Q�����&��K�;�h�ye�`�[��&�gn��d,�W���<ߙC�9	t�k͙@;d�Z����2�3�˝�2~�~��a�V����`k�|yWq�F�8Q�j#x��R�V�5����v��r���^�S��CX!r�c�\>��8v����z)��@t�K$Fg�m�$� X��i��2�P��3o��2<�7��[O�V��+)�t�˸��TNOΧ|�@�x+Ғ�c	݋@p"��a=m�ߏ�C�u���!�鞲F#��#�,t24�AP�9���l`1�l-�#7����h:����f���ߢύ]���IN+�v�=��rMs䍃T�ޗっ�i�GZ��nk�s���j$��a��v�9���3�S/b���2��$���2/��0b51����#w�l�gό���ygsj�åH��~]�VW�x/���vi��h�Y��1���;RU$��a<����x��L�@�H�YQ�=H��9L��ry},ؓQ��9�h���1���Y��P�����'�M��L�}���,x�*XD���a���W��?�G��5hю׹R��1<�=���%^�s;�����da~k�ԙ�5�)!䬭%1)�x��"��XB|���A��t�J𩌺Zx=������$��j�;�q�|�/�e=�����#? (�)Ŵ���̺l)JOo?�6�q:NCQ2%�$��B'��ֲ�[��m�.�Ԯn���p�Ps�4j%����N�Z�Fw:��[��d�-x�¹{�0L�[�}�9���ўn�@�������7��!`PiP}T6S�J�b:�^=�"Ƴ,�����ϕc�&(��з5�H7�ȴ����)K���<�a�0���{aA1��^�
�<rej�������v�3�;�13:��'�w"��t^�W>��vjb�ynM׳wW���k��A,��	�����{�H�o�3�ؤ�����������a|����^��1F:�H�r�!��IF]��0`2T������eL�$|�s�$�~�i̥�d��&�|�B�x�0G�-e^�]�ډc�j�E���(Ī�RB��`�T�
�kRA�p�E�#|iR@�X'ertjQV+p��4f�vf��=Z�Y��a�x�!m�����k>���ڌo�z�X�4a��"Y��u�t��Ǖ�E� o�鱕ۉo^��~"%?u_���7(��Nb��;]��x� ��� ���QΌ^uO��m��0wl�)�hXj�í 钃j�q,"9�i[�r?�EݮqԳ�����i� |�}��tSr*�Y�O����C��"�,��sԒl%�A8���
��(9N�^b)�~����^bi�%m;�9G�B�α=�������N	��1�C����e>������:�Ч�yz�����>����� @���]C�/�p�x�3�Í�Z�ᦿ���#�T+�J̒A�Y���}��Z���e�0���,����7�������ݯ����ڝ*���!�t+�ۍ�Qҥn@��J�mQL����r2ItC����yq���9 7G��?��=Д��X)��{�1��hF�H�m�v��FX�3����t|Q 2#"zQz�-(yF��ű+�ipٛ84܅7��_�j��1��w�c�� e�����ukx^ײ�=W?�����Tc09�^����8�O��Y�>B�8���*�n_{8Yw��G_�O�5|�Q�IN��̯/{��)�!���N��Kԯ<g����D5dO=��庿K�9����(�|�I�T��>�س��>�pw�����cCs�d�x��;��V�VU�Z'�3.�</F���Ҿ�������|�>L�B�f%�*��Ly����"]Gh�U�_��>(�	�3M�)I}8x5Ŋ�S5�k�H��+ީ���h/�c�hν�]x�.�W�7�#��`��J����2�A��A:c5n-�H�i�=Tv\��8��өZ���RE��ūD?��	�[�6�����_A!H�rf|�?s���xˡ|"n�i�OJcs䬂�}�:Y�񁨎1�͘k�/*�>�:��S���x6��Zk��撡�HU >wGw�$q=Z�jG�����"\��u�%�Ѥ`�qv)lj�W�%w$��-��#"jȩ^qnh�}3���~}%�g7��c6p]��ķ����_�1��	�L��_D����]>%�$���>�8(11hrі��_⺁���)4���Á�ɯ�Z�rȧ� �?�a~Sa���x�D�{�~>�)�&���H+�zUiX�nШ9$#��5q��e0�_�ሼ�%�x2]A��m� M���/�s\ �����}���E+��9B�� ���+@��2�f��pW�́{��v���9Я��Ҋ|��@Pq�o�xhߤf��~ۑ� �s��A����������dT�m��E�Y��k	��Z���ͧ�)|��U�R�� �R��Z쇦r�NLr4�7"(K0W`��<_����E�=�DI��jX�0�T�P>H��]$]S�`���q�.jG��@>!� ���ѭ)!��)�kD��#ص	�N�X���/$ �e��s�����3�����F |�Ѭ���%)k=����d���DU!�.���2Kޗu���B��ĉ�޼zޛ�]�^8e�*̜d���lCw��s�g�b����|���(�͓O��3�Y|J���=~���f^e9�'f맱D��{qcA��m�
�ŵ�����w��]�V�L'��^��G�mГ�<:>�����xi��p1H[�U� �d,5�Y�����p�!+ХD_���닒Xp�R��U*I�:�3C���aU�'���2ge�-����I���HFY�}44ԄY���Ү����,��o3��@r�t�ڟ���s��A9>L��Z�'�V~�+x�L
x�T����#���-�ƦKy��ܿ�ԋ��~ޥ��R��M�m���k qp�DA�d�����z�}��[2lU��z��)E
��$P]l��~�K�_}�HT����+���?���lz�b� �d�4�!���+�������kF��Ψ^X���N��?��t��B7>A�5˂|=�(��mA�W�v"�\��-�v�sAD�y��L1�E9X,�&�O�cs��*���	�힀�(L�`ff����Ma�F����O�d>�6�j]��� Rď��k�Ɇ���t���[�i�1依���=�[���b�����Da��W �����׻b� ]��BwXP��I���	�1`��=b�d�(��Y ����;�a��l@��b��=��T�l�����g��)E�1=���H�#�oP!�xh�+޳41v��:��X�T�ֿ����Nn=�0�kG�HJ��n�i=𗹥�}j^3qPֹ�\뽿���Z�o/YĹzi��9�t�}�4Σ����b*ЉL�1��K��}�J�!X#����6/��7��u���T�
���1# ӆ�QƏ��Y��Q%.R���݉<�]���H��)ǉe�'_�a͜{BC�"���e�� ���?��m��:b(�e�9���Xfے���)@@ǻ�N�ddf�(�4Ih�����k���� O�~sE}O�gq4����&k����n�K	��	�,��t(�!�V��d��Sm���N�Q?�~r����U ��?jslS�V9am�������#
�Wd�%�"�%�k��44ǎ�6����Np`I7����213�U�����L��־f�bGp:�����*���6���G�Z�/�����Y*Y�룽�"���@�@J�3x����Ja��ҭ�.:�E�����Va�w>geS��� p�$�ex�^ՙ[R�M����	2�oY|��(>�j�bs�~,Sp�_08Nl�ޒO��j$k� i-��P45w\1)0�����x*�&tF��G|s��s�ݻ�]Ϋ�x��G�_�����N\0{���+b���Sn�4/G�e�Q>;�����j�:���J�!ʹ��kE���Z\60{bk ��Q�b��VO,��o�R�Y��6�� �#���k�tg	��'�KF4�O�M<5�@��⥏ �Yh��x^�	�2i�<O9�Z(A��d���0�tn��g�GU_Fpf��_���u��N�=�~����'�1���H{s����@�vg:4s����O9���EE}�0O�JU��L����}j�3	�S����ڭ�y����f��&�(+l�@��N)覃��^oAU�!�P��Kn���h7�6p����F��v��޳�p��@��W�q��}T��0�4�F���HH��&�s:8=KGw��N�O#\��b���Г��%l�.�^��>Z5�s��ߦ� ����Â����g𷻣�pب��\��R�:�5�L,���E��Y�*Ry{��⿫)���r�.\ WGԳ\Q����~
/0�w�u��`�����צ�m^��Ϧc�́=w�'�rl��$G�f�`���/����t���M�Ŗ����ɾ����ѣ��˚W�����k����\J���RK;��/��?���;�X�a˼�%$yj�L����C;/�gIԉv�u{��I��r�����]]���+�����-s�L�����jw�Hd��'��B��	�'(���z�g�.�4��>�y�v���(����˯�Nb�T�՚��~AA(ARp�G0�s���v���,�No�Y�"�k���GU�l�k���7T��F�)1�sO�f�o˳�����W��*9����V=��g�;#�Q~��~�l��9�C�r��+BU������ 2߸JĂ��QyG��@zn��@W7�z�"?i-����y�8E��sX9��m�����?P�)72������H�d�B�C�w�����m,��M��Q0hKd-��Q�c�>��b�1�MUU3���K2�v^��Sl>�lT��!�������\�'��mz�Mxo����$W�>r���Gm�߷������R��$.���;R1j2��A�I�#�����>M�V�c<�����Wǒ�%�/�U#Ä�s�.]�H��W��ǿ���t8A�좟���0��zA�"��6 �[��>�q����G<����%q��	���s�W���,gIr3D��%��C#X���!��K�,��X�d�r��^�G�oF�J&|����n�6F��R�S�+�k�܋�����^�:�f+����A\��$3��Ĉq�. }'��;�*|��S�Q�q�+�:�'\(|+9p��𸤨q�A�1��Vy�r���	,��q֧
���^�c@��D�c=�GF׉��>�_���8�
��c�4b	��'�����1Qٝ�W.?q��Kռ�U���	MR�_��U7.��d�:�-(�&x�|?��%�S�������ý��x^H�$_�3$~��'�$��]�	�i� ��(�Ĺq�o�!�Ѳ�t�jRv[��ܦ������]p��3S���^ڙ���t��@�s��={��BN��qUK{�"�o����{�ėx�,}�2�?�:ʢ>K\>�o�4~Y/��x�:}DZ����p��LP���S�G\4nn���#������,o�4l�x
�ծ���a^�����s�7R�-��!T�1�b=���F�`VE��^ܤ�V1��)����F)�=n��;�t����n�%�
%�80ľ ?�ս
h�	+r?�xx��Y�*x��X�?�q�s�g�*�n�0�Nɣ�j&K��߮Q-�ןQ2�T�9)����&��V�-��aꤠ����:���,|�j!����7�]�t�9�QNq�T^"/'J+讴�!�[�������'vSMW6�

-�9 ���p'�T�h���;�T#� ���6�-�z{)�Jg+{�p2#�xU1�L7�de�|�`���n֐��xS!��s;{�~E94�lu�ax�sn�ɽ!��F	8�\Rk�j@�gv�1qikX+$m������
]�*�ğZb>�?�_��;���&��u[W!�өH��O,l���e)���,.|]��0�m?��dp�s_�Z�ߗYT�Z��^"�6�*O�L��=D��a�WG��_X����2�Bj���r��W�}N�g���2�@�#�F�@6o�Gh2~�[@-�;��Il!�V@~/� ��A_ܼ�Ʀ^@�R�4�Jpd�5�D4��YĪ�����,d#5W_̹铲��f;�aw傆B���+뽏Q��f[p*O͡S��C��D7�6�;�2���N+��i⃆0,�Zw9�L��&�=�K���n~EZ?.[Z��u`<�:+6�ϟC_<�ZԈϴ�HKT�$����p��<��j��+k
\�z��kT�A�|��r�)��Lu��_����&eK}���<��z�F�j��v��[[(zm[����O>���5w;�]����*X�ߚ�#=xx'��SzY2=���K*����wf�qX)vs[���=���lz)'��s�t(ނ������#f(���	��M��yޝ?o���	ɞ��H����0��&�[�0Je����iF)'AJ����.�qBaeA~APQ��;�-ͼ�-t2��9H`�O�
.�R��MY�'!)=F�ȃ���2�Yė<ʩ޾s�x��J~�a掽og9)k�|k,�iE0K�If��_T�W�0�L3��'��o%'�ꃐ�,�7�޺$��bm~��]綅��,����wi��1;�4 L�X﨩�i�Πx	q@�m�0d�\� �IH;ޣ�r5����OGȶt�<R-^�p׬�ʰG���M��-�0\�?�C"�F��f]&rm�l~��u��"�p��|Yq"ވNɨ*;�!9pp�=������+�y"'��\*�o��GSx�	H�(+`9Ճ6��<4iRl�d�Y��΀LV�)"��!�E�����k+Ko`���w��<R���
���>�����;�}��L�$��x���Y�9�b��ʃ�p���NʵY���^�baD�f!��횪)��nN�x���!ܲ%ڛ�)�����+�􆎎_�s4>z����0��"��FnȘW�`ڢG�~�j� k�Y�A������Vʑd�jl�vcj��1#&w7�e 8�����@*���䇤��+ŵ�����SYϳ�����~��j��Ĉ;$�.��m��/�gJoƿ�&t���"�h��xqy>��y9-�U��#"��d|��ỲPη}�����:�0�y�|�,A�%�܍�<�0��p?��q� �?#�d,d0��\*�/�^�^YĎ>~w�)���gΰ�����jW��l��DJ^���2-j���Y#�H�i�#�*��EĊ��9]�
؎�ݦ�FY��x^R�l���d4MF�²I[��.@��WjA��D4.8��	�xs���Nu����֣+
�SĈ|�S�,&8�W�W����h�g!\�-��w�&b��;�j�Nb�3�@?�J��>	�B �����}�Pk㏲��y��	)<#HVZ���+?>��񿩿J����DZ6<��R\J�C�����6�:"�����Ȟ�q7P�x�Σ������ە3�M��>��`W�T��nn����p!������tS�2筏LH�1��|��Cbu�"bu6��K�F��
���i�6c�zf��'�/��_CHJh����S��6b��F�"F�c��pZ�}߅�э��2�dc��i�c���(~�C�C>�:��#M�ȋI���5�8оՈ�}ޜSPr]ߵ\!�T�(���[Ԅ>&o��9�tYߐX��@c�0`���T�/�?��������f�DB�8�;KKW:�S�A��_�Qs�c�`V7y�$8�r�:$���I<�݇�De��[Y�L�bT�$m[{�/c�~~jNK"��h)�D�E��\���M�����@�[�� ����&X7�虓���M��EeOҡ�)֒ڒ�A=m8�G,�3ugP��ր��bz�_��w��o�|P|�_Kd�+S�W �ᵛ��2�DT�R����y8���Ȧ�2�N������WY�.�ǬP܇�l�љeـ۱���G�0sė�rE��
]J���,������
�sK혶,���θ#�w~[���o��g��]�_���	rz��|j�;'���"*Ǵ�X��FYsd�W�� ҃�o������oB{J�`3�L��y���_��P7���&f(%uڌ`�Y�ó�?~���3J�/U.�����S���M*R�$i�^[�g�#؍=pU�Q[�e��Ba��}~��0��#������H��>�퇚r}�c�+�����En���*��`,)^�D��=a�jR���C��y/REM�w��*�	=�$��w�2�k�ݼ�J�!�4}E�g��{�08�Aֳ͈�L�Tf�$��[J�����`�ʉO�Ѓ6SܞA_���/�0$E�
����V�櫾��f�EH�! kh��#Р����*�z�g:�� ����kG$���W�n����##��u~�`��:Z�4���c�%��[4�!�����k��0�Z�����v�7F_>[ǻ@�Λ��O:|��q��8�P-�ݏ�l3>�j���$W��42B0�B��Tp�:i_;���S�L�qE<z�&Msc�8~t�QʊZ��~�Y���X'(e��5��Pi��(�˿�o�e��i{$�G�l��'p��~��m%Ir+��G�`���Zc�+��}�]ȁ��8���|��ϝ��>��Ƈ��
o5=6:v�Y�[�����W��Gp3�۾8�n1$Cu��y�}���~��.����۵ic��d2�V�VP.&�U�ȼ��œ�d��s3�5<����Q;H#�b����2rI��*܃�m�Ʉ�X��0��F�PaD��g�N�G�R��R���V*7ϱ������0/2+��z�T��RIػv}:܏;�B�weᥨ�o�Gj$l�M��o��5�.$��w���7��p;�iX˙m=�b�XUNBo�J�n���aa��:D3pɒu/�Ĩ"q+�A�6iKĞ�?��nq�%6�<���qPZ�S�fw������Op��o\��/�,Q�yt����$���M�%�A٘/�~��3_}�3@q�9��`C���0��X�!���XD
z��~�._�FFR���ا]n��L�8�f����Cˍ����Ѝ
^�f��E��L[:_���ډC'Xzm/g�Lq6�á_c1}�H�N����x#��ד	�,nC��[��M�@
���?�zJ^��Cȯ���2b
[Hkzҭ�}�7���o굕sx���k��4*�zl	���
>df�)/l�U��e��v��F2]p'S���v~�G�������Rܖ"Z_V��H�q�)k����� +�7����:rY�;c�X��3o���K�z:6�cb����J�ᇄ���w��p�уaۙ��k�f��А��3�m�따-�J�L����L��O���v\����,�L�	>I�tlB�%�O��䆤�'���㕥�P��W��"��/�AS�E얭"�ཋ� ��vH������B�����ú���G����+¾�
B�����aɺy��.j(6\�����<��1)�{�*oh���63]U$ч<5܋`� �����Ћ�.��2+ͺ������@�C1e�Bo�V�6�o�6$�}j�����<�k�UPl.�J�#L��T}v5�jҦ>j�:pMZG*�t~�9�g;�syoEҘ�SĴ�$��� ʌ��y7A���1 �
���(�AKD%�8�����{b�dE���j�𲅆G��('o���wZ��d&]� T�slg�b�$BX���'x�A��iӶ�0!�$X�n�OK����f4�W�v�J���Z��l7>������\�6FKRV��2�$S�(+�����"��'d�U�૳X��)���������fV���;g��'�|3M��ϵ�:�UN���h�/<33�<���'^ƨ�� �ש����5]m���1_6�~�C��:�͑վ�f��9&����v)���Q7� ��яYg��/�EI�	�����l)f8m���)��,ODja(Cc���iF��:(��5�O�3��mQ���h�ށ)%��$`=]�ۍ{�����w�q��J]�1��fR��
��~�#0�\��si�W�O")�%��}s:/�����ۿ���|	�y��>��eH6>0�u3��pUQLࣘ��H.������.#�g��
oO��4�����CDD�ſ�Uj~ѭ�� @GW]V��uߵX�zB����#�s.��|�$��|דM�X��^�!�c��P�Й�=]��	�q��j�v��|]���=|&\Q�0���Ƨ�U��f�ycJ)��t�Ft�*$��q"�$����PDɚ��!3��)i0�����*A��Q]3턎uTO$P�X�J�	�bϕB�xnx��^�CC�=M��$	�������1S�?��j��W��/׎52�y{��1'�0P���6{�Kz[�<D�d�&h�!�,|kdܥ�b+p�x�E�K��Z
�s	m���D�P��'T ,rru�'L��s��w�%]cۦ����]u\2�[�^5O�ϟ.gL���4/��ƥw�S�����8���^#�G���rƆ·W��Z�,ɽ	��Դ����n��:'uH-�g�i/	��R�1T�ˢM(��"�ǩ�X����`V@8����j�gj�����W�2�#t"�3�eoE���x�Gw��/0
�rT7&�8�]Wfl�UZ��e�S��'�����R�S�DpO,�b�N�|��j$���&Gݡ�_k8����f��m�5d�fM��h($�'��FqP�|��z<$C�.���H����2ܝ�H��ѪIzF,������҆�����%��Lu5�؄��?�+��s(��۠=���ҷ�IJ?uq�p�-� ���Ol��>~�U�jV*�Ի�Α��FV�.k�cl�,�o]���P��CjN1�w���冖� S̍:C����
�ه��$-�x
���t+ဌ%Gf^�����3E(�%�>2_Q4��E��
�)ʱb�����H>�I��о�!GBG�/Y�k���([X�!�Mg#��W���r�!�=�a�*6Ep5�|��Ϸ(�ӬD��&��v�*�q�/�r��͊�3f,	Mj>L�+CͿ;o�j�'t��^�{�9N��s0�{�)%A��P�M����m��[$�;�������h�
�'H�q�w׮�y��]o���D}�@:&C�n
������Gc�w)|�Q�����>�=��N�G�P��{�9��f��' 1	��ĕZb~(-e�"Vj�皋����X{�҄- Ek�\Ub��(����P��n	zj)�����6sɏ����Yh���+2�S�9�Ad�!���p
����p���ׄ�/_IS.�G<e�֖���>�7|�R6<��%�?<�>nu�3WJ�B�;*��س �5�$��7�萄��L;#���Ԏ����X0��t��\�i3�����X-���HH���%ʬ%A�g��i�N�Jf����y5���S�P�I�N��wu|6}�Ñ��B�.�CBb�9�g�����s�p�q��?r瓣�1U	�ƴ��h	�8���5�=H�罧�!���L�����}/�"���W�2\�Ž*��K��gl״�׎���l�kӪE�ѐ�i�%R!���\��'6��গ��B�U1�,$N^�x��(���#{����_�U3��X�b1ԝ*pM��&��b��l��6>���a̽o�&�����*z��QȔ%[�ݩ'|[(��k.0��n��B"-lo����;Xinr٢s�B�@X�`�]�o�v�Q\�$�M���o��^	�V���P� N�(R�:��5�|N߯��A�:�Cxܲ�T@ƭ���C̸?ud�[3s�?Z��/\�d���v3�\@&�!�e<)�6̥>TN��|nX��'�:y:O:�����uU����3s�̙T�{L�#�]���~����2��cC�B�'������D�;���-�2��K9sʤ��QIp=U
`SN�=ٻ�s��f����A�]\C}�10֩v�Lk��Nzɘ7����;~��TӲ)������E���7��3�N��ڴ��8Լ�Ģ�Õ��A���$��iվl�	��#|=m:���
Kf��f��,���q����Z�;n$�����3�9 ��M�KU^�2�I�������hTZǷ:���X�zF_-h*��N�LÉh�ǯ���X�����`�&{���/7��.g��X9/�%u���
��lb�B��{G2��|Q���������7aDG���F��xUatz"	[_��MƥA�]�j��_F��=�}�S�PqCV�S$Xb�Y$�s�k+ssv�3_�5�v� �z�K،�ͥk��k>'��MTMIUh&�S�~B��=���	dr�&���j��'�M.�2�ӱt���U4���
/������Y�+` f��޳���i�Oz\6z� Z�7��V[^
��WOJA��@��I��	�Ļ�4��#tއ��+��{
7�뙔b �sP��t���xT�k�B���)&J����G��p���
 D=�c9�l"�N�zW���߭� �[�g�hܓ�K�����kfo���ո_6���RT�S�?�v�ֆ{[�aAf6��r�U����jhT�5�٣�U��8_,z��-� jq���v}($�W�f%p�*��U���m�=WB�lv�(S^$<�"�;Ք[��5}�W@v��[�����o�,ׅ�*7'����#D,��%O�7�sL���}?\�[&����}2���Zc��#
c�C#fյ�N�r��g��4t�}�ִ-u�q�w"�y?��l��Q"!/��T�0��A�p4�qZ�9��Sv6E���|e'��&q�j�EfMq���))�T���8��1�3�j�3D����(GN̐���D��!��@�;s�<�]��#[�4b���	b��D�~�H>oHb�I����haQ�|7�꒸@p��h�X;��1��ǵ	X�]cq�C�&��1�Lxds�x\�
����"���$��.�Du0��7�W���Q�%L�N���M��>�ۖ��YMy`s��5��v�h����Z��>B��r�AoLN���|�������s"��K5ϐ�?F	�.�ffI:����Ҷ��0<wM�UBl)Ҙ	��7�_����	L�N4����&g,F{�@l:��Y�����d�5���Y�돮o������$q��e��������1�b��r9���
���T-۠�5�v�<2΅���ߛ��AƏ�<���Pс�{V�신���Ō��b򗩜�yr`2t	�Kk*��%)g�Na��,��"��}E�lK���h�r��R���OK���I耔�qiШ�g���Dl�|�g�ت�5'�%�w�����dvL:Y5�W�������_}v��\u�K�@qGe�D�o�*"�F�/����hv��`ϷtE0)�[�lg�?��CƂ�����y�HQ8���>}ׯ)%:�H��V&��+�1*/&o-'K5�0��,���:�*����]���|����3e�ׅO[ ��%/���xCE����Z�R�$�+�ˡYp(���T��������s�&sI��+����D
�܋�l���K�8�/�$^#BM-�@9=b��@Ϳ�ީ�M�|P[���O
Sr&�b��!7�������O*T����6J�e�+��̇n�̓ۢ�4���a�&�}(�F6�G&����on�s' �[ʸ���E�f)��q.�p ��%"��m�C��������k_����K&ZH)��>Q�� J�y�:�������q�MF<�.�5h��p�w�v�J`�י�b�&�7���ZaWv9�{�a���4z�Ձ|S�\[=IB�'���E��r�OY�9�8�\�>Q��|��ԙ�b�n���N�AG��9 g8�#�-a�<4�r-Y�
�Тc>bт� �{8pL����s|�w��}��k�m��je�����.#gϓL�M�x��t%o\��̩�%�c��K��a�$y� �>9X�u��u�a ~��(����o����dW�!��B����{��ݸ���5B2��*Yu
R�1#��TЮn�Sd}6.��ȟ�|$�p\�FF���}։��K���ҸVI�[����W/�.�.Dv��/ȯ�<uW�$ u�K�=Sm�s�ؤY]r�09�+4��f�#lh�@�w��V�(���]=��;[�.��Lo��m��%x��p$C�p�j�kh}Y�K5�Tg���u\�++~�(� U�r���c0Al�W�{fX�����V4o�W5ŵ#�r�4?���b͔|iG`���4��9�ر�Z��
D'�<2�8�D`�'�O�x�NrDH� ��M��LAB��n�/aO!Ȕ��YCX8&O��;C�>��\�hT�?'\���Xh�)/;3x�
�Gqu�$yE�}�,O�	Yfڅ���,��s�t/�"���� �����O��٨_yLP`���Z�0�3�F-�('z�t��C�/�h��!��ë́kU�e����7�`{>6�����p�Sa0�?���k�K�o�^[���P�����3��9��v�(cz��R9~&���(�^*X�v�P�qg�<j���)a��{��TL
���wF�[�4Q���R1������j�zjɾ�<��S��݌�
V8W��i.��kYZ(x퓨t96���+E�W��	I��c�%��h֚j�2���l��'_?u� �2�7�hMuw-�x���	��U��#��
�k���Ȅ�f��~�{����u�oZ_�X�i��r�jO���3T�>g���I.Ia��G�^�3�*
�LȉCl��k�!��Ogb �/�c��4*iWU�&A���$���.�R��s�v��W Y�r���Ѹ�&�+i��q���Z��+/��jC��B�is!�N�~{����HX_���T
 ��K`o8Z��C:��p��QZZ��6�>s�u1�ݛS��f�������S�r�0��G��B_OmmW�t���>|MZf��ree���Qi��^(�D�}��Q������ovu�=E�6Fc5�y'1#���5���W[�1.��&ևw ��gP�,~_�ʩf'�/��Wֲ��|�GG��ѮqM��4�4���u}�E���{�D��h�� m�/|L���T�jr����zM���M��0��ץq���t��M�lU��ϓ�I�w��bS�M�!i�u�4gg�a�="zZV%�iKGw0�+�N|{�����XD� �Žz�e��������݃�m�64�|��\��D��DZ�zX���d��.S[E��'(�J�h��#| l<UFd���g�̻�y}\��.W�ㇵ�>�|kj����j���O��S-�C�@��ƒ0��0���uA@(;1�8mɷ(�$��M����\@0)�-i�2Ӱ�Z���@Y�flթ,|?e�G��@7�ͪ����v����	G�n���1��8��W}N�Hȓ�/R��i�f ��f��2d� l9��J��Y9]#�����0HO����9hu&���?:koI0Q9t��E��4�3�Xe��;��x��/w����ۥA��!V9�*���x�]��C��;XObY��R�,�r:D�1��������d���R�ς���|��0kc�ޤ_p���TBab^��b(j�R�����K��� i���`�+�kMЦ&�d�1G�(5��B�2C�4k��9+4����v؛<d@�s2ݢ4yj��Ŏ����VX�>^��ᚦ� ̍�b��ר�<Q]�>v|dIq�f~�fꚥѮ����T���z;B{U��IG�`��}&�b(�ƒe环�Pb$�U?S���9,W�8���FU�"1ռ�M!��z�Q���	^��. ��κ��=-s�����9�� �T�b@�wl3�������i��[�=�J�N!�e����6�!��s�9�"M��.�D����a���Y���v7��]?s�g�@\�P�?/b��͘>�s^���P�����b�b5p��z{1@�z����&�y���E��f9Y$	G�ZMt���m�-3-Q�o���]��>�
p�A�2 `@5a��ا7|��$s8q��;�̯c�\K�/��)V&�
�$���lV�g\����,���1��3Ȇ�Ř8I�%��q�^��社���*��['���p�(�g>)mP�`�W�	����j��J��/ZerV��h�!�#��	��<K�zx�I�G���\a��/�pi1v�P��}B��}#G�!���	f�i�~�_-����废c�C쬽n;����.�Ge	��~^?�>��Ә٬12�tW�֙���M�|2��y��B\�l��T
c��Vp��\J�&��-N�*���y*�/�{���\��w�p�ʷ�W�`jlf"MJL�ʹ���ڍ�f��ۣ�u�u�~[#벡E��i�h("3��t=\��kxz�Ɂ��ݒ15��dJ��w��b�ߠ�
�-w���e�"?���FHP�Ԏ��3ǥyr8��^'��H����ޱ��w6�残��!�DX�aEl�\�HL���>�Zw�=%��=Sa�2��@�OY���X��Y�C��ז_4���~�,~�+y�#
����O�t�hX���)�M��k[�O���갣h{h٨� g�{Mp]D����lZ�R�U�Y�`�*���5�H������w�6@[Z>��z����^)H����_�v��WfK 8=XN�r�}_�l�"ȥ/��4�����dy1T
5FE)[��&�����q��nұ�d���I�_~�`O�`r�6^�ϸ�خ�!�/v&����,���~�:�`�f��m�-`*�Ԁ��!��.�D�t�"IК�d����v�p��?�]��A�"��>��	ںR���?�ċ�MՈ`�� ����ܞ�\���  -�%����H�❵�{ܲ��T1��1�A�O�U�y��M�V�n̞�J��^�f�rsr����q��;NGcݍ��~&ԃ��=�'�26��cu���L�t
�hS�PѷlH8�[�E�Şl=�(�{a����V�<�K�@��Gt�-�D�7�Z��<S���4<-Oa[n��Fm[�<���<��=����_i2v�1�����w!i�<��� :/���_<��L��[��8^�� �w!���>#!,��/;�^0��
��3���[&�Ǧ��r�Q_�!���u>Us>3~~����48��������w4n�:g�_�c���)\N��	c��۾�)�\Ɓs�eFO4��8k�,�u�\� ��F1�%eꀞ����d��Q��R�̒�tm���(ڛ���Vؙa3�2o�(؛Dl���E�����'T�&H/%(^��,�������%��%o��|δ�� ����+����!4O��%.�NJ-u�];��z>����#z���J�5�v6�r�}:��HQ�6�E�W�]��H�_��HB~C���ڃ�~qߜ*
�5�d�ǐB�-�|k�3G�6Ϝ]�ETi%D��2z_�?����7���}�6;;KCEJ��;��q����K���eV;��IpU\�_i�	3g�Z0��r3|_+qs7�����m��P��Vu0�P�r۷��1�v锭r�hr
E���M�����2�h�p����="z���2/��g�C4o%!�8�Q�S���<����sT��j���u)뼙��[�Y�&"���u5p��-� T�a�z��a��!�7�$��E`�4AGԖ��V)r�,��3�;o:'��/�ۼ����BX�v�p�e��M�u!i�=	���*1ÈmO���^�G��S呅��(����0C���Ɋ��i�
B?�|r�*pɤ�����w�$t�{�z��˾ �.���0zҌ�/h��;�%�8[�.15���2>�a�:��C-B�Oܕ]�� ����$PE��_���浂�z�\�1w[(3�0�j�$�N܋E�1<J����Om�s�,����'�|Z(O��$F�������d*K9��, ;q������R�sL��<?��@L��%��_bҰ��?��
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y7'�cq΢�s�+۱���lRK�s�]=R��!�����,��%@�������˔����DD#L�M:��ý�᷒Be���0�� "z���A(I�^�0^^��ѐ�!��D��]�Ak�6���]�4ʳ�03��ּ`74AjLX�3��N-7�CY�����UNhK���#4�	n���J�]Gϡ��l�_��'.�%,�Z����2x��]�]:��
+>�K��C�����7?����\|��(=�>q/����"?D�R��C梶�ƙ1�����_a�rW�K���������v�\|��D�T&M�om�Y�n�`��	Jk�ՏE�j
�1֋|hP�	� s�$�
2f)�;�5"�Y;���\�z|,��~N�S[8\�����^r"+�ڌ��f�>Av�s��D���<���^��j�OEf�ײ��I��>��W�Θ��Z'��/!���ܙ���+�0o)[�����C�i�a��,�/JQ�5�
<�
��t��[ʸe�Ò�p'�P��?���l׈���=������չ�eg�μjw�]�)���M �����_0R��Rο�!���]wp4:�����q?��p�@�j����=����#�B�N]y����G���M:���T�V�zyw�O+��^�0m�l�]/�@_���_�b[���.��6��N^�����P��yu��lP+�F<�Qr1{+��7L� ����߲���D���=�����{ϟ���`���7.��*I3RG�7d�-�{�4^(/�8��c��ld{n�e%��k�*D�&(́TG�kB;�~�� ���1��2�M���؎�y�1�c�'���H�x93K�ї_x�kFb>Wn��n�U&
�;F�0�Y����nq}�Vtp�F3ǝs���R���9\s�Z�t*.�4�$C���;{V6����U=�/�Qsi^�"q���~�aPV���2���9uKA�0���Y I�>~&�����N���v��7J�+�'����1��ɇ�Pwx���o+\�� ��!��z��e&�C�MP9�);Ciz�<F�Q~��)��E.��0p�ꉔ�i�r�sQ�̌����x�.ȡyc!!�w>g@�ɩ���ȓid��rv ��!/fL�2~@�sl�t���¢#���<�������F9�1��
׳F��=���qk��s���^���}���F���l��r�����m���\��K�� W�Tyn����ourIH��q����F�� �tJ����*C�C^Ce�{PIE]q&V�,5��g�>&�Lf��y�v�K���A?E3/ԥD溝�pc��g�9䀄f�>)�5+�ݲ���WՓw5WC��ks���a�2jfuٕ�ob�����&TD�GU�A�DYg��k�h����]Ԑ�X��DLטee�'��@#k�K]C�-��=��U�+W�0��b5�w�JJI���������iм[F+q�N��n���?E_�%Ӗ=���Ɵ�$�qg�9��CV��i� '_�V����a��U���3	�f�Yxů�;�swj�2����oe�}/��u4삩B?��\�P0T�P�h���!��(tf�C{�f��.ǳ�}7&�`.6O��fj�K�W����i�=�5����HE��w�JS�i���"�/�N���
}Wo�"}�(t-�œ��(�t	�t�Q��������]k��#�G�.?'RZx�-k��]�nCT}4�A_y��Z��Rn����uHi%��:�X�O��an��k���<m䙡��������i�&7ǻ~7�P�c��I+��v�
E��r.4HcC=�/��ue炨籵}�8���g�*ac�
fS_�!n�(��r�����+��C@bXBiPz���`��f�a݁q�8�R1���O��&�3���H��ȝ>�j�m�>-e8΁����8V�K���;�f��!�u�<��^��4q|�a���`&/��0�Z�s<	�I �qz������� ��e��}�h�b�������`+�}3��'�N�x@����cI*���Q��v\��6��Q(A2X���%E#�?���r�+:IP��!H.�0�ob�s�m�֖�O\8sը�����X�����Kz�L��ݞ!}�n�@8��z�<8ej��R����UG���*� D�Ա�H��0gE���/CX~'���zt֬�ֆ�g5<����i�*�[ ��R]�o��XK"��,#�D�V
Q;$��#�>�5]���U�׹ۿ��кRׯB\X��p�aތ������1�;��$E�}m�����{"c���a�i>.�Qi�|98���OO����F��OR)�������7MI���������w�l�
1���o|��S&��|P�� ���৳W
���=ٗQ쁮4PL(=(w��_���g~�m��b
?��GO�6�3�qT�o5%<@�&uߡ(�;}��_�������G�����f��Sv�8"�c�jM��+S��@����ۯ��c�89��N��f7!�;�ޣ��n�'l���O~�����g�fR~��̯��n�pX<68/]J|����Z 2bM�i8�S���oK�+A��S�=6� a�0�6Q�����	zG�ә��'"K�t�Q��49���g
�#���ފ�,5i��7^c@t��#�_c�$��V�/�B��J��.5�(�������Я�E�B4���J1a6�����pK��LI� �B'��NUE�1�)�Ek0���U���3�������I[O���n������ZX�n�Y�!ig�V��[k�&Y�ˑ��1rŀ`��G-i(;�iz=>���x��<�Qw�U�U6��:���󯔜4��l�(��F2
Pr���smPI��gnN4Џhk�Zn5Cf�:-��B���@�	<{y4����#/���o[���i됵3�U4���H�:Z| �E�V���;/����d�0<{��}�p��5�H
l��82ޙ}:廣B�+�� y����${��	^+�^;��?��?SE�E��k�-�]�/Jm�x��y���6�t�~Y��ث�Q�B��T�G��#�O��Yh��Aϒ����SU}d�� P8�,{�R�\�o=�?YFf�L�[�n�\�N\��X��n$��al@�\Aң���|6�W`����M
�"��a�^aS	K�U��`@6:7rš�uY�R���O-�Y�����D�n��� �%��4���4��ث:�6-Юr?���
����Q3٢�M��0F���'964�?��M��%K�X:bv;a�4�hzO�t`��m��j�$[uo�jAh"�|7�7M+��:1�}�~A��4*M�ʌғ�x�DS�s8R0y��{g S�>���֏Aç�2b��>��G�[㜀���E�ad^�����,��E�@��,D'x��5����׿H��v��ܾjq�������Px\���������
>�V�C����������h�
��O�A��3��Ǖ�kz�X��
GĀ��ZEُӱ�(�"�1l9�z�&�j ��F�f�wXq9�� ��K;����`
��\Q�m�1ʹ���?�K�r�w�-��O	�wS�ݽda�!�M&Y�XMŒ�x�*��r˕	���q�bv�c�pqqZR� ɖT�{�@��A+{�ͮW��~��r¡�U���{V�r��/S�|�Ʉ�[��r�g�2�d�D��s�����R�5���gf�z�#���@����f��w��'_6 J�,���^@���x�"5p݀�������>��t���S��L�v���,D^���R���֜���9�m������4��۽X�~�I�T�xT�~xT�� ��~L��tO�5���Q`,�!qU�
�#U�0f{��遉p|g�k�}�ћZ�]#`��1�z�k�D��%��;��PT�c��i$ݹ����N:|\�L^�L<1�o)U6��4��$PMD?Z�冻q;���N[�N!O��R��f�=�V?>�rAv��w��9�9N`$����%f�'/�lR1��� ��0}Gvd��c4�l��N'ā�n�Ϫ����w)���ª|���V�� �ͣ�^o�4�zR2���n��(�ј�J ����=ޣ��auR� E�sp�:ܿ��€r-Q����
t���
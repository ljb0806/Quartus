��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB��1��F1\HR��`����+�)��#�2_iW�{�pOB���3(+������lc�)g� 7>Ox��������L��*6�du��O�?(�	�5M_͍HQ�A��x�e��!39�}���[0g��<�>Ѫ��*��_*=]������&Z��*���㳵~�p7�u�ߴ���5�`�k\��J��j*��c��;B*6��[!�X1a��
�5H�hȿ��ų�7DC.�bM�۳c[�^B���5�B25d1��{�ث����N@n˴��W��FVi��"=Z�~�
$0E>��Rs`
��"��4�C_y\{
J�96��^�r������d�T-�B<�� �C�`�� �6>�li.��"��2���N�J����w�iRM�!ǎ$����$n���?�Q|��w^�*-�F�i��fG�TD���Ó〺�o�l�KXγ�멅<��[p']hJ@����Ǿ�`�G)챣�tIdF늒�l.�+�7�ߠw��T��Q����9n���ͥ�1t˃�Y6M�mX[���G��G��,Y7��r�d�lL:�R���K��j�,�Tsq�"4OV,?������\�W�J3`���5�0����4n�	��HQ"U#�����,�����{�	�o"ӺW�E�50�mn.�E���T�@=@����mF�3�1VM�XV��G�BA�� _��NfV$k�c{��@�2�)j�=��
�1`O69����p��+άo�9�� )8�%Ck�Q��i���2�w��Y3�8����
f@��ػ�z��`�n��,�E�MU4�us	�媧���J�!<"[�M"�c�*���o^0_	��_v��= Yc��mċ�(��<�)z<\ϧ�c���!��A�J����f`X��&���4k��C,����N��ߤ���IzC_��n�ex<�p ��X8*oݱGk�q%�ga�"޼~�3�Pg"_!�]����0����V��K"��K y-	�ϕ��`l��,�"nb��U� �nx�KNGL1M�bD�FHK����`��Q�H�=��bMH�q�O�4�ɷ���K�������7!0�����n��UN�I�a�]WR&;��(�Q{TӸ�s	F=�����!iwKa�gva7����(o����T�O<��}��_�dsD�� v����a�%��J�R��+­��Ǳ����7�!�i�>$Q�y�t�5ɡ�}g�3)�o�T~@������:^$͞��ط�E����@���(�W��h^r����Z:$_���R@�lmGqӗ��z/k:�觜Z��[��s�an���bR�e,��$:W�d��v'=�+Q4�\��B���;W��{�[7���1|��[Sv�
�[���!�5?���¾�b�X��X�L���:ꌤq�H�k��o��P�+ ��>-Rt.�?.�����<:���!�@��43�Mv�n�ſ��?���?�`�M����`Yg�~8B_<�#I�߲:#��xCG�5Q��S\;ڪ?2�<���NY�K�������i]C��3���'��^���`Q?!΍Cu�+��+�`��^��8�FT��F�<���d�m&���UK��4��_o��}"��	�=]�:������+�*S�wY�ܽq{Zx�� ��Ф��'Wm"����~�a 7S�����6]ѝ�7��3J�ޛ��&Q�w�o�=f�i����}�i
��ж=�� 	�w���B����x*h��_H֪���Tz6�4���<�!P����AT@����.����E�rc!��Z�� �TuΎW����XOZ5�:�@�fl�*�2���Jՙ�� 	�4�X��,͕��i ��/�X6��o�neӁ��a�j���x�fŨ�I�mw!j�{�h��q{ad��0j~�R�G��K;5E'��ĢU,,��z5n"8YDo���h�v3���U�*�οU��!�����Cxf���4{<�G�8SL����L�v�>W
Fw��E��]�.>�%�c�A��Y��L��y!=�W��
�Q;����b)��i�{G�L���\ٌ�d����Kr$}-�K�}N���Ƴtұ������wA�R&x6��VHf��w1`~�<B8���]�u�,�D-�Ƕ�PW(��uuNI��V�y
7���{%F2�j��P(&n����I�
�����	����j���;����
�Hb���>�	�
-#ߘ��U]g3��� �YD5���z'g!�/����	�$/܀R��wN��*�mA��9%�Ә�<w(;:��}Ə`&Ht��Ōc�^����.�}1���M�IÔ豔��5C��/9��\ 
����v&�ώ�HR�I �n��a%���E�E�+T�����!wsg!9��%z�T_��t�y���{]!5a#�?D���A�)��0���6 ʃ7?��L����K��E�/����T�d/��U�@��P@!0��~�	�8�C���e~��\%(u��[��m*�����Cr������F�V�����[�P[՘<VEΦ�8hL���~#�J?Gy�ž_�7Ly�W�DL�����D�h�v&x��2�9�����Q�!0pT���oc�CC�ְ�m4��5����Ui(?������b�-�P���I���CN$|�KĶ���d� eןA�4�e]�ݛ&og��?�����;e ҵ$�`]�&�q��
���=���3h����(?���[�P�s��%�H��� ���q�rL�ek=�E���-= 3��ʨ�⵨��6����=1����>��7½3�3����@��������n�u���`�h}�Tt#�^��y+W�g�3κ��"��Ɂ.�Px%�y�#_-��П	�He�8�#����1�p枃�x��|��K���<{�}�p*��p�Љe�O��m� ��+��Q�4��B7C܎n��ϔ5[��ʻ>����w�������f
]	9��IO�;z�*
���; ��I�1׵i��/��$ �d�.���E���ՃN�᡿�{��r�Ze��+09M�ިe��D^X]�Y��<��۟QQ4��Z��E�����nC�n����+}��N���)R����Jk����-+ۧCccN$�屔�8���_8XG*�T����A�;��ʂ�rB�uN��Y��v��c}���n�Z���M$�ާvh;���p�ʤ>�Q���h�c~~�N�!�
g,��
İ2�9$(��
����!q6��y\A�CV�9�+Hz�E� �x)��pR�\66T��rKA����W^�)�.1p�-��pX��e#�h��L�� �y�j����Q��]X�H�Pޭ1�d�Ķ�m>���m����ud����0Vy%�\������2�M�$����	2�x;�K��uy���9?�
Q��*�M?џv0�m�l��A����]�Mt���0�5�����L>>�G�_�ɓ��Y��抲;_G���L�\��x�K3��.wA�����B�&>��Y�X��X2���^U����^��_f��g5�kJb�TЅZ�e�����MW>g���������U8V=�����S�M��,N�m˟Q��9�oq?�������gT�� ��5O�4>BOĕ)�:��/2�"�8�J�|b��Ey9�f6�X�.\0 )�IVXB��;� ���6�M�^����	�c�Ү��%�~�� �!U3]ȸ�4z������S�
�l`�|�m�" ���ˡez��.��r�����gS��~�ώtZ�W"�SrN��\^?�@�s�q2�\�2 ��MU���(4�p��"/bU��1��
*n8&�Y���u?��̂�q�ڄ� ��v�>�%�y�ҵ��$yY� �P��-��aÂ��X�cF���)���J���|�GA�N<x���3R[Ys��W������ܡT�un޸���Z�sv��$�k�T�+�>z^�<��^�S�9a-@k��E��b�u9/��jq����u��Ph�k-5/������� � �DU��kЛ�vB��_�)ȑ��V�Q����yI����,>۽���C���uW%����k��n�O���bQ�����d�lt��͹e�10-�œFZw;��-Jx�Dԑ͈@�p?�fMs�;���a�p �k�Y��|�)P�C�v:����r�3ȓ_Ű�I�<,6�����3�̀�7����(rSi��v��f����x�x,����~9��~�:1��X�9;L3&�+�x,hF���HO�o��Ri���HQ@�?���B�P������@aߦ�`A��NFH@���4��L�y'ʸ /pM;p|. 4,��ʯen^��p�'\���x�>ڱ�"HF22��HV���!c-�]�((�6TD_gS�H����dr~��~��(���-���M��ȿ�?7Y�{Wj5R�s��!�Ц�7_[��cIr�86����[
�$H��7����,��_�0�ş�i�tF[lm��F3��O��Jw��L/)�a֍'�V��&H�N��&l�Ě�*9N��h�p�x�����R�c؃Hub
J�ʵ�9��Ek�LE��������K�VB�[�kC��W�L}¦�c���K��M��ެ��)Ox�+��U�T�����!��j�@h�z��[�&6���=`�%�I��e�n�d/����HD�j�����,К���eI 0��.j�:�2@\�0+Q������^v�������E����.LY�y��D�OV_�*�SO,��k�g��o唡������mL�k}��'CF|�!T�o��g> B�P 8�Ĭ���|�׭��)����H]�	����U�r(��h�I�<�!���̬M
q��	�v���{�����~it"�����>�B[c��W�Ґ˨��3�K�1x�5�R�_����W�9��d/
:��&�Y�x��
����PFs��8$m�{nngj̨�F�*��b[��۪��!μ�2�u� ��C�x��ĨʊE��K��H�
�8U7��g��v3O꙽B�=����0�[40����**��5a6G93/-��2U��üq�9%p��MtC@�RJ�v��	�^�F1ؿ���Ki7:��'����fټ9yժ�^�I��X��
Ǽ�g���婒F��z�ą��*����T�G���멄ƨ:\����E�/V����;Y���D�8r�T�o�"8.�A=S.�s�B$;���(�?N�x��@y"�s����bQ�W����c\�xyg~�y��	�6����M�/��w�X���ƨ��|J ss������v�Y84+�����"����fr,��7�H���a���4�
�l0���E�
bn����h1�;�󒢃�_�u�Ǌ�,J�
B�y��Ae�<N��"��Y�����݀���V@4���Nq9j�х�餍�/cp?��#�@G�ݹ�ʜ�\���M��#*�����6��\�"D{��PyP��5'��J��\d!o�mn�.t�j�;��a�ԍ/M�5IX�%ڎD����4��xF|��߿VpKZ�vyb�u���IH]!W�D)���aB5���R�"�k�H�"�_�9 �������"5�]�w�Ud�3\�b�e��������:g���b�.+���Q���gr<5�X!���&�8�/9˼mİ��r}���ձހN&Фs$h��b�}6>�&�܎�w\Em�'ߙ�"�,�B��⑫��e�uߣw k���E���i���(�%|_~���^�E��w�=g �;����v[�eqD��J n$��{�a¾�p��=��(��rorAj��[[��+���Հփ)T�V[p��);NN�5grA���R��e�jʶK �^\NQz�a�j��|d>�8�����\6N��C*���r_6<�;}�p��5;2�5Y}���DNo-��,Z�a�!��,�ݽ紧���5�rʪ-y�kD��2��.�����.c����,��Cq�M�������c�*��e����i��PC+~2�cS�E7ւ��8=Ͷ��{¦-�{�%Or�
�>�b[w���>gT�I�o��cbœ(�]����m-a����7˕A�������/�}T�au�e��0����_2:%TAc��xA_�S�v��L2!�Z �A�̂N��K�O��.B%ۂ�(��s���sgüJ�H�����8�>CC���p��>�1�(���@�	ښ�8/u2��uL@����D�p5��1Kt�NP,��o�T�������pY����ǃ�Ko��d��0R�*|e�#��Ǳ���!Pؓ`��0[��^��)8�4��c�����o����w�zDI���J�/����q�c1�~�X\����ĤMM���UKa��X|`b,w!�~�u5�}�K�|Z���ۑ�f��A_sa���sL2W		ӡgQa�Jt�Ж|C��3ҏ�b��sS�6bo�o�$�.�jt}�\H�9G2�OB����Hn���ՙ�9���5�ٲ��a�J1�yb��L���F�x�=�Ahv����K�7����	H��uų�۴J�<���dM���Ȅ�!(%�m�1���n�����-ԑ��QZ��t6��6=L{�¢�C+#�L)^��썂���n���_u�J�xn��&o-�~"n_�G`Ϧ�C�iT�.��Z�ؤ���N�,��cs8���D8٣{�m����h�(����wj[�Q����d	$F��L���ξ��8���u�B�&c��Eq%_>��o����)&7�"�on,�|Znl�J�?���������0��k ޤ8֗�I�����R���~��b��,>MV�(e��F��ض��I��I����䏮٫3B���p"jI3	J-;.j�e�D��(�p��:S�6Xx�i1�����c�����AJ*,�Y�Q�O995�՛�bP{� �V��l�`�yIF�DX�o�{�J������3�^�|��{�P�v���(�k��_K;K�U?���o�>�C*r�즄��$}kO�����4�Mx~�X0���ůH�9)�hs@�ZH
ɨT*~XxB�ؚ��P,זma�kC�C�hD�5��}=b��	Г�Oz�y'?��Ż�,q��Q�e�4��>!��!��rÐ~t��M���9x��fR�T�he�Z@�͑VC5
eE���	z��G��E������E�t(��/�`�v1A�A;�Ҹgx�'6p�2�lz�4��U�7�1�8L\`xw��86�G=����ON��
�Qm�T���8����l-�/|3I`�
q�r�bi���aQ���:���A.����+��H�Ճ�3��a"��o�CM�ͼ,v{�ҖX��*���6�}؅(�(OkzW��Ʈ?����?Zp@�g����d���_�n&h*-��׬��+�N��Ď��D�qv�r�*���(��R;�]i��0�x�`��g�A��*'����_;�i{|K�}O�yDo8�J?�_Ƿg1�歹�-��@�<d�.��լÔqx��?4&|�������;�[QD�ۜ83ܧ52�x���]K��k^��M����W�_�-�m�5��D_�;̉���<]KOA���j�ڀ� \	�.�O��\�����l� ��B��ޣ�8�\@�vТb��I2�ـ�o�#o�T�?���u_�a`����$��-�����O.~E]SE��	Vq�~�|AZ���ѿ��0>	ef�j��"��/�0?������A����Q�v�^��^h��!%i�BW3������3N������M^���EF��#���و�ROǤ��;N!���*G�\�ع����l��{���eFXoO����~(I�
y���7����_Ķ��&��� ���!-����tʂ��]1S�U�"s������^���|�W4����:���'E��te��)�.V�]y�-L5��j�E)tC{�_k�5���wa)�%�š
K(f��-��
;Td+����G��̏Q�}>�Sq�Ro�Ỗ�Q�h
lΏ�E!^ �6e��U��䔅js�s�#�c.��-L�Gr/$)��k���D��b�D�!"p9S�+	�[V��$�%$��n)|���U���*�!�h"`��eQ��4w��1��Tk���:���,�Oc	
P���Ȅ�}��� ���[�b�7�<{�;r�B$z2�K.;k��eA����VX�6�-��g$��7�?"��7_f� ��f����2Sj�ۭ����l�̨�͸�z�B���B�i��z;7�;H�mo�e���%9{=�nX������_F�IN��6b*��֏�	:iX\���4�'�D����r�����L�
��YX�䟥'�Y��n_ݥe_!-�F۩�{�Cl�EKYM`?���@�cC�ԢHt|u�R�Yr��ء=��Ct'�L :l���<۰)(D��6�"M�1��P21��f䜲}�6�kjrN5���
�{h|�e�D��A�Q�
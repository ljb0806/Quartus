-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ESKa+Lkl7jyHBypqpBRIIkoF/tGUd54yziFYnpfQVqwEiETjxN87nRxfoB733xTTbYPsRyalSC6D
+nWp88quzCmBZJU6MIO0By/4VP4VH7RlscWYF9eTrOWG3rn9UzC8Q7sBu0vHK0O0kuCms6m3JiBD
pDp9FBPpiOtoO/KuRyUnzs0tkgvtfeM07TDJeKzZWyzNxiHOHBKsUjJHIzZh+rE1puWPo04oa05J
AW+gLg+Xsct9egIOwRf/Ey7//oeuvpInH+P2qRTvc/ZZYGjSIpNa2Tpbbt0Ys3+ER9bfIeuBRBZ1
DFI0bI5tT7Ap+1WnTjoKuDOaYELMXpI/O8BNTw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35184)
`protect data_block
fy+zq+Am2lzwD+IMISCPUdLgsraSc5SHiy7lhhu00GJQpAoQBmYE/GVbuBji41qWHPFaCh0aG+fx
MRdoPado5D7s9DMyxMQ9SRPElVLrqKm2e0+YShiV7LGfmeU/3szJeTkf9WNlYe94jOpIrzzXguec
NbMP1HJjHCkHhX4goXhRYRe21y9ols+MNy5MgR5HcIIDPNB+Bb0hrXGFlC2Tu3e1itbm9YwCgyjx
ah536K/N6xBmDH1kSWwxg1eymWuOWTEd7b4ZRcMJnzZ1P6kknT33aKc4CE3GfYr86xByloX+okeh
1Z2H3BiYhjq4HK49jbfNFYJ6Q81EB/lUBWT7XWVrEzAsITH2VZljnaz6dd0RzXX+rwdJ0ALdCXSn
ZGKrWc/oQEaniQP6gydW3k9icDzvIl+N4fRfh7MhZSYZZ5ybxkHfzpztLwfGoYDINwx4jDrYuflD
IGFGtnyyG5CQdDyDOG4nUEZpC3YX59ZPzA5EYqPH0FPOR6vM+wVQQ7VQ/HcSe9jGXJGZ2i1D6m+l
ozhxg6yH4/GFPrWWrt17PDIUR7a7GTlRcWaEPs4mGu22VHYJyKTSeeB5wolU+1e6CjX2f8uK1gD9
XhGvRvSIFuZC/qCmtLmzpcxv9ePML3jxxMTPQJWzR4PeCplkEGQYUV9dO0Y8cZT9xYFzm6WH3ZcJ
RnfqrVza52gkiWLVPYuTPoPJh1DYDIeLr859alJBWE9JtK9KPb6XmxFmxuxSzJAXB8USqSuVHQrA
C0qHYSbaDNgiDcEUkyZUSQUr/JEppGQ2RqcJxj0C8AItYl+ZbgU08ZZyCzHx4PINk2DFMhfQ+Ck/
zmv4xdu9i2htueVIg7VtNRYSeiDd8ibwELUvFp4AnuuFPC9h26vuzQ0za1eQox26emmhUgsX+qvD
0zGxV2e3cB7SWz/T0QVJ8DNZdXLFdDdfLUG2oxAZj7cQchfnyqRrweJyLR9k0zcOmApTFZgT/Ra1
0gsA3qrzcH0iWU8IHOU8N//LvhIL8MVtd+OwGkjqwmLXh95ZhUr0eR8npHz0JRbkfeagycWZhHud
xjCDtEIL3TCq1r9SJzUWvyT63VMIaSvCLA0ZkwPReJ3X5n7T7kWEUcwzhbtpjT0kKx0tSvw7wyqT
qPnE1IcYUwwjHPJK5FmTYU4zrbjx688bR4UHFkvSXrVnuMvsbR6wQCTN5xvWt/xFcAhwHB/zxukR
P6JCPc6uvQacY1JG+R6BqPEyx0MplpJwrt/Ke3avolUuE/fYIoKBiINnfCIafN7+tCnBdJQ1Oa7O
pS1CMMdMju7A3XkGXbqELKMdD5azKkvdV5sL+v3XgyLAUut7Pq6jVHgXu+SWrQ6qe9DRYLYp0ErR
AxTdtX4OK3IWb7OZdFxL9KCe6ZxBQLyDdaxBdHAN0BQQcfi0UcUpJNR4YLeg9rrQK2zzwIK0KoWZ
wj8S9OID2tI1gUqKiHdmI0uV+qg1zgcgEEDkWHRVREYZu3PC8dfoYypw3RCNGdHWmvI8ao1Kbyjy
nLGGNpmQ7Sd6/APQ0fPTD/5E2NLr1OWhSuO2O5pIWXASdw+4Aa47Q5sGEK1u/bBEcoN8ih4XV48M
HGzXpeTt7Lqnq9TbE2vIOQidL0YBmXRfytu+3OR/avg/fvimE3Nq684w7+hRfxN90NsaCbfavdKx
POO7jqiC9bBzKK2xnPSof28NjTuJaFLibTGTkv7IoSynPPXx6RO51R/1F9xHHIaiEjcWSHWx/2X0
p11keumrfsAXJgSggnWTMRraBoNwvDgiD42jjQ5e6FOCAhvMJidBVbsKnqDzf2noqPlqkVgLxy/m
ezy0Z0cOhZ0hbFg4okhWjxau7wIPtn9mgMDogPikT41kSM4JsB9QzRQlAcA3hOpZilBHzCAZSIve
dIi9wPAuVEFVAsHtYcpzg/0cbqwytROyjjKoG6JeZZJnnwWqWX1lel0carifbn+0zQiP1qgP8suK
WbrZErSXz5S/xbfp2Roak+vG3B+/1G6ckHTMWlWB+K5Ohmwz8S6gkj/Ady0ACe6Rc2e3KewDYLLX
rbzmCiVkeFOxYFWd9rY8u2yTs9cZvfclQWfrNj0ccgmjr/lp2rQBWyBJfIgi+oRGO8JWmGvicAiQ
AOjN/CewA3wRN4KobwmbLG4Ly4RmlLVZwiVqjWzXER7KSfjfH6s69tXTrW/LEvHB4krQwJPZuayk
lacH5i+ImyQo5ZO/g7+uMrj5lkKl0udbL7BBYJ3SvNHmowyNHMq/Np+8AdHI+9IsHJBFwSiA4Pzk
fnLKJZU5wuQ+zeIxhec+dpCcq1or5W6FZw7yUgzYKaKiXKp2VKttHBngYrCmUoS5ZCCL0G9YrseV
muc6SkyDQk2lUWdjXLo3PRSdK4GwNsyWs8YqfnqrQ+VdmUnEtZyRh02Fz5f16Q5p53oeSeOTP6kt
HmwSygClreJKNULotUg+H7WyYN1MqbyZQoT0a7UALTSpPXl8GEyyPY7ZqROF5e2gYvGQvhbuLGr1
BnQNr9F70RsbbcCLAUl4WgBb9qqyBojXSRNIpjwEX6IflMw+Ufgx+B4VMdRP596re1Xral2UE3v6
4c0RbGpuIDKShIj7kxJe80WxWTx+iwJDH+WL7jf9Wlkc5bP6xHIBD87TGEsHUXa80mcihjYCgoKW
2Rp+F40+oYeyPQJ+4vKNkdFPPfZvBwEikrC+MiHODmkw1fnpnw3JG5JWpD5eN2276Wx7cTzlvzzb
BT5nAvWLGhHMkbOPJzD95R5VGspFrE6VVsc9G5xjifl0X4vpp5FAQuSmhxdbHgvd1TW+9PHft/+5
sUMZh581KB1kEGf1XFgqK0ub2blq7wbz2GSqhu5bus3iRLVTjF3IlL5LIceCYYaz94dV89cEpegu
huCT8KGLOp5FGjzVC/QAn4BLCdqvlyCeQlXL1bPUNss3kSLMWISNJmRVvj/tKR163YBQmxvXd432
z+qaeDwa0VmpsUWmGt8dk9YPZZyUNsTHuHVdzswdS/4kuqHMSzpjepWfaiVNrn2OqO5YZ4NgpWiM
qVZKf3G3OiX2Q7mKrZB7FKw3WrxRpIlhQl/uBL0WLHXQCW36WpDNRRTWtMxhNzGC4en/QZewMEcZ
8UgGkL4t+dRy2sjeBRklOIypp+HQNh5AbqR5JPA/8SEiOF9vX7fI49fI+1u6ZbFadgxJNKpByzjR
TG41+riY24WSLBlERi4HSYTfqTF8jITSbUqAk0VFEuNaoJKc4Fj3Qx8KcJPlZ8eSggZlqVqUagbB
8qL2dFdUMMHNP7AGzvO4WR+dY+qFQP/mPag4BPSHU8i4SFvAzkqHAS0T96BCP8+AhoVdu95v10vT
8GmS/t2FGr9Z8scO6S6Y2bXfHR29+7st+W+eyT1mAD2GGgGoSCxL1X+5lDTikBmB+NUdb2ukzwF7
01KfsHWZNkE0wo2sXd4GZpGitSZpE0afreI0CNWd0xzW0D9LbCicef206FfJp3l8FdWzQOSBTUTY
Flz8aFvX8uVvqIab9TlxCtS6hzEzclAUDeT/UBGP0sipUAF1BeGZnYgoXa1nJOTdiZJAvPlaRN5f
EA9aC2snHgqVgG2NIUZiJEoTj0qorFzvO5ngGi6ytjiml0N4ncQ8BAxnxG+hB0+Xvzu7roeo60pl
IDjKxdWIK3ydLGt9qiRea6+sqwyAtHRm+UODW57iuxA+8fDWFQn4PZyKVoCo430hWkyzEbbn1fiI
lXYhrAi9PqzzIch20n5GIs3BpM+6+hbruWdRfxZvJJa5svMXAppPmdbHw67WNkPn/pintI6vbtC6
KxAELbBgsL5eqxu4CZvxI4q4hQFFWWsSCEwXhizyeD78rPrI39/ODEzUvAvfPEqhFmxI3qQPJQmX
9fxZ5uzpfjb5ifNqXX5zDEETQd+Q7ifPXEIY4OdZzwp+yxQeRFa10LA2kTI5se+AvOyE8+Y0VNut
UB2saBv7S3LGbyS1IvcV4n3mHryZN4nDWuYdumpHkD+Rz4En4EO67NifMSa5jBj4zSauChd/kMrx
z7bLreV7xBN7V1IHE1IyIu8kubC5F6c4+7ckOpQjDB3IDpjXF7Cqq/wFQy4YZRcP4pTGuJBVQLEk
Low8p3lPx+TCPJT2YKubWueZuqmQvm6Bm89nRCej5Oi5ulMgbJ2IqGs76gIgDRImY6Ko+T/UNIzr
xNfLwwPziCPGVxnsjs6QMp1yN84e5MmbubPcL7gi+elP0lNhcNq2+O0pwhHQbRi0ybzvB35uKEm+
QOxvflMDc8x81qDs7kbvkyjwNlE7xCEuJCTwM8TDZ6ohx/igFdaWkweP66E34V1GBcKBtPKKkSa5
yE9e3U2bH32AcCm1Yn8ZVJaXItTOs3ie5la5l0oBlcTqwRpcRI+RWslBdAe/YwD43UU3Zva9OUIc
8+zgnVsUnWTmAd/y4T8eVTJj0nS/PtW2SfhD/NcG8+ysu6Hkm8aYOeWpRXvQUXlbKdG3ZAJJY8ok
ilRrFFuwnpIYv5ZxEBtNrnD1DfPRHrHZdAusMUiKFtYs3aMN0Kz9waxpPlVy9hDwpgOGLdvRnyW4
ZJUk0PXbHGAQPgJAtu/hk780Ica2qMLIYmJ4vIScXVcfsoDKMdvOG/MA9yqcVfjzOjspjGBpHbow
lq3sil8kWy9Lt+kqfuq4FVEfL3Dm7rKC37LVPoaAA7XNS1qxIocmyC+9qfK2wV/FKbYBAhE75afn
QocJv8qSBG4PP4tmENc05SH+k4wbQGAFtgDQ3/sc6XOpzu40KmrcnT5jKprETp7NsH6ZK4aETxOS
gtcu5wJoB2jslL5C83EZLFgbfXH5BSQMBWEu8xyYe1/ztD1SWKgXFcZJ2PnWrmX0WMpSQJxldrhO
OIkkh72BjoetbsKuS/FPUvRzwiyOHWgp/L8HoNGklxATxz3L8tb/TZkmPQJTuD7n/bAV34wFMv2y
4eA+/1860rXchkvSVkrnk0sZMdDnmzRam+VYPwNvbUGR45bxEE7DHDmk1InfPlLwFZ3jKrFn4xCF
/CZgU2XimEJzSv1Oa/YmLZBZS5xGnsQSyhDQTr3jdSScT3zQ2D69p3OBdCh39iJ7LCuMT/I148QF
cl7iwHVqs2kMJdvKv5NtZUaRCqtTGI3Rnwv3pny8AZWXw48zve481hvnQ6x4U+9ZVWYCB98lITL9
LDLUAqongsNmFr32xn4me1xA7zcCD2jL7WKgxCQYvI0+gb0yCzn0Ik+yMisCeTSC1soXPX1QRJrU
f2lcbv4GVB4NXM0aNGuKnr51cl3idciHv4cBrwy+v8QsF9XAeemmOlTWIaOlU1EfhhwoDew7LK8+
E1uup7Zkl1KEEpJJ0LeB9msIXYb4wRkqgmny1Utw6PYIoz8PD99QZXWsh1ee6t+AgUSsfjvD5Zqf
cVR+XUhHUl4fYvyWW6m0mVO9dJSwoJ4/ZwgmLZwG4GqSIrZ7JGJM9wjwQoEpnWReDmU9BTy4pXnb
7x4vMBUxab2uCHPlHWE0Nybtpaxy9YZT19gCN0/hgESxgBMutwgnXTIs7y1Nys2deFQga49klJrq
bvy1tUqSk/WJdCzTYCvS54XqWz/ZpxUagPLN6WUSW0OgitPJrBFqoUtAZyx72fHYCertoD+dJ70d
azu477a0wluddudpmIa4H3YA3S0Xw5O77VObWykKXG95qb+sLL0AqEDtVJs9BJwIA4SsoIvzKavA
vydv5wDvWoS5fMCZHb81PZmR/crcLud0jeDyInwXEMhVfqZcVoe9EZf721KGvYd8l07krnZgb40P
gCrcF0amGrO7fESeBcGfY2sdr6VxtmNvzw3GQjec9EfeQCTKQGWS/0lb21j6QUvENaw74pHPxg9e
/9qMbhPQLSQusHSwMS5aNVSd+QX4bIzRzgAksbgEZNZJz4S4I2he9yU03d7DXSbpK0qRTLXbQvkP
IpyQgzR2kxDjnKGAO1mftjny8R9Di1WT3CR8KhFhNOCw9suLH0l1LuGXGKlXAYNQ1P1hFyKUUCM7
pFhCJIllG5RZsOwgK2/LP6oYOpfDFN6+UxHSnUCun3W4NNZKxOYYXys6wlZ/gZHdVlCVERZZq6bF
bs1NykSiXZPZJ27ZrP6aJQA7OjixPeIsxLl1gsCS+o8YdZ1el6bZrGPrvRAX8uOJBPVbH1nBnfKA
CEh7hEYxRELpUE4SY6xAn5Y+Dw5eXU36WsIMXbkxkBPK188cKN7rgfVuDr4vVYJ4aqrsioXdbJof
i/sSns5O2oEA2J56NktbLAljwP2s+5+OXJBF4fQF+Qw2bQ8bLTb/bVHDa3dlU6P8giEq9uUBZCgf
4C7jzzQCiU1eWhxOqTikPyxNuf5ibIU1IXmuHx0fOsMLebsBpMg1ll5nDFqotB2MLXNs5pbxxGci
srssZ0lfJJRwjlh0BtjMjak2Zb8EIVX5O13Wjk0pao4s9uR25VE5O3xEe1Z/YFdXiYL12/PJJpMR
azrM1+gRtJfDU+TPTB2Trkz96mW5yoOZP1I2ClvVUB0sXz/isu2NjLBVMKDFpUxwfVASdFpNCbOw
J/5ayY+luGh9w9BCfW4IKNKMfRzS+QXdoOMvtJbpPBfYjr2Pa0VYUzDtVYHvTsT8IQSTp3qGmqyU
1nW1ILo3SHO2f1xWIfVoBBHwN3QAmAhyjrArP6Emml8OXEz4cy/SIKhvuCZj3BYh6gO/5oUjIiWF
y1+NP0K5F//Lx3E1JzAbJLy9asNBxluX3NbjExnyJcO80s0b4UZV+vgWuRqsQd6J2avxbygiDgqH
a9v248b65XjeOCOJoGp09ipwGWpe+uNNvN3jw2DLnycLmOqNDvFvZiDQsJlQJ3jDHChw8ZrxcZqL
8sm9sIODIJBfuF31F+jwLvzitvPD8ssW7q662wayUiBYF8kFeKAktOAb00Kxvr7rFKkOZ8fz7+oR
CmFJjIlAQOjL/hg9ixOD3L50urWkFiQAx+O1rnELsk+3CgK9zahAwCF0oTreA20vAjWWIOJXBawt
5YpjdTIufmYT9NJJtIG+Oh/nwGOl0qCywQiOYQX4MiCtHT042quRGpQlXpgK6DaXOduWxmfqC+SJ
LpR9JCU1fAOVRQLN+SqjHs21n9+W5DoziBFVrmeiY+fz4oJ9uCc2iSWOWpGN8JAsePUWXEaca5DM
xAatNYz+Zpxg4uCnc3YsqDWZfwF/Vya0A3ptQ1Uv88gRvMnx8bHUqZe8bCJ1mGp9EG7AHZhnXnkk
XvBfvqbPWTuMFxq2kahFEm5fLIsWPOxV6nj/z7sL/nnoJTSU/XA2DxJyN8Al87qrGTcdRDShRhDW
ViYgKC0hYAu9YEZbPRJ2WUd7O+ytdusFmC+nKG+dJezd/vWFi0g7YGp7sig5YhtP8Ga4Z0+L8F8Q
vGNqJX2Prdx/2aVEwFvsE/jDAwGobwZlKaRHnLnjOS0pFQC1o0F3M35ultYNhtSz5AAMHuABnAWa
NeS/ERjldB3Q6AkRJnsevA6O17Bu6dVPVopEbCCvc+CfqwA08/pAtyo0TBHsNAEHNPmbJ24Ndaqk
lbS2wx/5eU3UyJPNd4f+yC8CjhX8GmbSsKstYSnepS6uM8Or8yT1aAk9TkDG9tsvcSh3plOa1oxJ
rjZdxVvPdxm90HmwWTkXbCUbnJUdAW14UTC1pm0+9EUOvkmVXxsS3DIb06AGRtX3aZmmrAxUYr0+
MAwadPmL8chozR45eZUeQRhVTREAN668FhGgopoNoy7PiCJY0vhf2jThPXPgd1zz4IRZTqUdRvoi
1FwpnJDfCP1sRkr0YOa3SQ964RH9gety+INeazNsaQcjVWBZARcHMQDlYAxILBiH8gniDUBbLUno
MnAyTrMhwUT009C5lFlaG3O5LILGx5Ip2zM4W2oagpbAf9NGuw1vxl5pK7hkCdHLAoubdezfHpUz
9i/RFsjxEnHFgfBmE79TjjN61kURxpFE3oJH5RWIL+s5zv6P3TGusYGGSXPEM0lbLP2RDjKRCEXU
HeLp9Zslsa8f2iD/2aT6N5ReeEXRlfJkypfrm4px6AmSDBUYTkaouSKDCP0Fy125BB1o1ayA/n7q
DKzaoER8rlzT9H0ONwLsIWpxOtzfYT1SOnC08L2MIufE+HFI7HiP7YwUFqnWKe/ViDg8/qhaxlon
9ZEZefALHCHpHKYnCL+oT9oGL7Z5t0kFT8ZuThfhmTKAPqBl2mGxueq+cAj5UfwHfSRSTqvYXHzp
uZ2Y06M1ImsDq8uLYr1dj0lIQU7eE9dJzF0dHwqJGTmrmFnJz1spFsZHPZD5ck+JjF1ccGoc9gs/
Vdo8Ku4bH5HZsm69Bmc+J3Ow9cP7DDpXU/mUzIgZCSBmw1PZ/O9rnno4hCh9/WlQ59V3PkNSCJ1v
guWKJcmibWwKTIT4/RGeEXtIgStpWtjEsE0unKC8lyG7Wh+mcAQ//tIVZy1dfzfw4lratuHNF30k
4sC+Yc/hnUO4CyjjUtlvVRXdGl8CXNnZogmD0t7uae2CaZ9DbSekLkvcbpzQpLp7uMzpfHSOWgEu
GVtR3zPqkCJtTcHlqCoC0azYbOJQDpUpwKvD2a5A6uyT+jRmyRhNZxLe12OFflEMrHlKBLVENlvE
eAbbtp+vzJBGH77hJ1uwHWYlTk8CBKKuc4SwohYYbQg2nvWG66IvTohD4WzGo94zFii38cpNbIek
v3PBL5xYQh9BZzSwCwIt6SSz1nUvjqDZwVJDgkLN3xwoH8GBdcXBS1cLi3WtY6DpmWeD0V0b8Wa+
AJakAeqjH2dyf+gKiKPiY8wRQ0m6DGTLbTZd4holXN1mQ8T3hzdHuDBmNQ6mFhixyAGFHMPKSOxP
xgCrglsvhUDTlyXDl0rBWASvC2ndbvor6pT2TMIuYLOngqSeNFFrD8zGeGIrXslj6MHmwgDq7Wki
GJ8rAs0af9XOQn0w8HfihmAVG33lXQYGzh4SOqzWGmOklHGPMw/Q7IO579Y7Vb8c135LhpCTQywp
I1DLgPqF39v++zMLArUC8Xu6vzAJgFy7/7qhj/IxshkRbRHWc4tVbZh6Cs1aOwjDzM4EuVdjdUxN
dVAuvBr8WlEe+Hvcc3p1TAjlHsZPxz6lmCyeKB1wWMUVzLDxPEqnNLqfdvVFiJxBfJoFhNfsHvKT
9JX4KLhACHHMyULLQj6fACVc512l7RyuAW4kKAEYikLQwKDw8Pr5TwWVlLPJ4nDyo8vyVqb2sXcR
l3KLvfHvSwbMB5CHLOD08FCcqtyTKwSFPeIAh69FJDTUG5aEqQiujkOJcWSsNkrT9HHgf9faEeUe
McvTUPcZ/T1wzBMSFi+27T/PouNaO74nVvPCIfYYLQrm9a+yIUrHzBSBLvSuxzIZML2xRx4oVCLw
zUoba5QMozXP1vwyA69MaoUsWDxKjP8mPiwreq03T6H8VaU59S7BFeFhhBd37jReqYkxCT/IftG6
kellaA1UBmgJ+Ij3tgVdXeKVxnDp7JQ8BnIFW4LQ5Zm6j9ejyoNDAePtxXG0670rryx48hja47Lb
8rHappzOzsBd+qig/xn/5QcYWxBxQEFA0eZc7gqcbhsgzmnRLMFyyW//DPiD1u2iH2MSRGdF0gYV
3cQ69np5n/DmbeBxJwz68cAM5WFCg5xfFOBvynBvizURwsYW0k+PIBZmbUJCmXP6UHejiusoQjMz
ZhtvVKdJdyGYNh0yB728OegRluIM0jwGPu0thXBRtle2EZ9Kf16CfkuTX0koCEJMjQ3bX5gu8nHM
H+vEEE0Un94Ky/i0YdJoduvoO8LM8N4j5ProVTRAMLOleCckDh1BmCZ6HCwGUoJ+8L97/6Zw9BmH
T2hIP32y6NPHB6g4Mwech3qGZQvAVjX5vu7NIAqJuzFjRJ/3UCVIEwtQbMo+O/izY2vk+rXju0uJ
FBtijxSHfJz8NXGF25YA5Um8yS/kF27pcGJCERr/af9OFbhsK1Uii+RMhG+vhNIUG3kjFHdAqsqC
jRSu18sBJs1dN96OoaJzFeCUVVjwk3YFTMqG5yeZQl12fFCcq15ZQVbXE41FXxj/e8f47TKF5kJH
Hf4O90lL4WphX6mSQIFHWinXZ6fHXTzB0aqkiFxAjlK5xl/aea+VWHrdzz4Qi28qRYgE4nhr8dBJ
XqThTsOQi0yHj3EHbdm+EvoCysbglGy+jxxILPA8NcR+wjnR/+2DBRaZpJM3GM46hrHG5OPEh1Hj
YRAl/m8CvZfO7FMW2kmspABazQ3ycLUwIfs/h08ajhvTLr5a8vzNRbu0lVv6VIh7SLCrjy6ZERsi
D1DfnttAykq5forhK3lahPYO6EVT5Cf6a8RJNvAor0nslSUmifq6t9WXCeUu5AL4Go9x8l/WCF5f
QgWtr5QZmilFWpuZc8Q+Di+eatQf24RhKuOh0ZRZ6zjpF6YmRZ9oftVI92eg8mIFcYHX6Y8Fwor/
cX6/y5BlbZJCKghrzjAn2fIrrhgxibHX3o3KYl/PjB0vo4LKUIlLYY7MQK6yZO4vyFwnumMA658V
ihhjnz01Diy2mkG+LcxoSknoNRI8uWQoN9KKmtzJDRvI4nFht4tczJA4Z/fiSmK2Z9NmQrNO8ux9
m+zAI204Iyql8oVcCLN/HPviCnvygFaTeK3PBhu86I/9DMEe4bi1oKH4BkZEanW410OAP3oiH2p7
pu3pxFNeJiUylV6g8A3w7Zq5lzZM7XeAe06hppmVVZ84lDy3aQqVfKJ0Gu0ap1E5nvwIssoTukzZ
GIHcgedhTVxqj/gaip/SnX0VrO2BcAI0rinHyxQEMy4ENFccUUJ5Q4NJt3Mjn3JRDHNNSHZOfe3I
PXlPWq6hVkTznOqP0n9aEnz2Z67fTwreFzM69rQnWr2l1fP76oaeZcA4By1OsM3Kfqef8+NDGRg+
11M2yp0tn8f6HMb9ICGS51SM9lzN2L18NQWs6d5VD9LQRl/vve97p++ZYKp4VojciYlJKrA7tK48
TGJaEUekaJ8Q/NMbrKHTualwBvpcwz627zCKx/3LiPzYoUHekpc4A3okYNV1ULh7Z2Vz5O7CWgf8
5pt1DnXXLyjuAFbvK63tIYR7HNhIsczRBC8XCVnPLh92Gw1QbSeGRyHg3a1nsLoI9Ydu6y30yviP
bX95HEaiFkkwQY8nWPpu6w4VWRbxvBZegXHwbKBqeXBkmCLISszQY3Yk8xrC4XXEkZ27JdaPV6+X
GNRkwEN6gTcaKInMzM4At8rl2y1w0PdGgXvwFl1ez+UZyfK8E2OJ+J/WAZwVnR/UkaRSKK+19HvI
tbtek3UrC0ZwgH/ldjR++Q8YhiVIKsj7VBbruChBT+gPq96y/kVc00dG6wKxYyURl81snGCEZQut
sEIqKFxL4oX5/644LTKOTh6/nSFSs49aFpjvdZoeVgqahptBLwkUqEIZe+5fxGUNLyGEUMhfGDFP
CffjpD9r+8W1RCj9JahUOj/SbA1fCtJK8NMpnJfj5/AXQTmF/cnFP74gWRvJm/5hI5TDEGrgLL+W
PMyQ7S0k9DBH/hJiZguNb0BJhJOsuYkpr7isNxwmtE82ueBG3GxXPBA6t2DLh04RvpHX59xzEc03
kFSdfnKDsF5YqV304rm8FaHjDZSBFUyz5H77jHWZxM+a/ZRmdAE5oQRTqusBRdDkizyuG/mw/Vux
eeLIzeAri3iQNn9uprurUGri61og0ipL23xW6Q9QvAuHaAmpxxGC1SSa4E+cJJSyIbpm4bzuWxp+
GmsnD6g91R6rFUztUXqd4wT/hflNtZw2aCKlQv9BQAYvQjbOISneeBKzmLYqkbUpHW3p5ey/XD2o
yThQSqcL+GRE8+p7CyWdGqsHyGVfwh359g56fwVpiZ+j4wrfJFQPfvekWNFCsPW4oWrklxEZG/og
/ks0LrWSwPgVCSsFe+5nCQ4ODfG/dT1TkkYeowTXXrHWjz2HNmH43HFMfkfTuT4bEIyal7tWrQIf
Ss353VOzJVDOUwcdUrxAQxQFQZDUsWd4xgbNsZ2sKuP9ega+tVpOsz8vWx3dt9ejjtM2QYgUGnaJ
/Es+FIBdpt2mdfHT0DFz4n5b/HduxvuzEhu5+B8yHvQZnQzHZJq+i5B3em956dSBik9TwGuktVN3
GA5ZkevdT79typ6U5ppuu0NPzmhXTXcxgeQ8JVxEeEm4x8EjEi4VXHnnhFe4MgrfvPLaMXhHLrrI
KsXlWDdknAIe27uTLlj9IfLP6TS+0U7HpDOPlmovu2fvwQfRXBsXf4EDTyGbuZGV2btx3/LUojKG
DM4ZF8DSXrl7g6vFID1IcW8ekVDFMCWSXgcvwPNSFOSTdXyA5q0/XfHlJNI0HdJhm5jWsQjLVwbg
yb+Xn1OUROyz52yyw4PIJUqjKlszyhfXDmut3P9s1vj/CDLprxq9fJ/GmGigo0hEB1QRN/TgplJG
EnE2r98m2DoGBFM/l5lSYMCuA4Psbr9ZbEYF93tL4Uu5kltNMEkj+bQFSybrgMy+AYX55I11ss3j
9U35IUszrR5gRTk7q1wfluOxYLHh2jg5Yr4pISdh7mDhRn5iWcMxdv+dusfzfKuQt2zQa74TUnjd
vM9zym0B7uYJ1YCGqml2Gd+Ek2hX8wyYshIcDFDkN5+NUUmdFWqr9d2+gCBNpcOydRuWH5diEhWx
TM0DUYdsz93dHdcz/w0KEgTKoDen2EN96AhqislT4uWwDHCg/dBudsObMVeIOemfP537dWaq+WID
LNKLCYp1w4WLd19m2atJqq28iihvTyz2iP9svu5YdGaKImiWxX3ArV6/wcATkSo7SYcmgW0w4s33
44VjUu0dNaiD9/+SxMOIawtAImr8rSpDqfF0uxPQILcAXO3LfrPiM2QkkJtiL1WXzWMq5NmcxG1n
bEzYg2h6toNZ8zO8dJqSENE6KlX8Pwzd5N61BJ8bmEM5JWU9IMoeNrDNfDFrIq/rkz0mE1K7Fp6y
+u9ILIWLV8ZlmTtT0NuwrQxy6XvaqHxWV0dgmcvaX11r7aDHl1pul28yFwoAMebTYq83DGaeaVIB
sRgh+gzAtEFJsjXtO1uSKQJWCS1o1mxudnMfWWoVstuJNaJ7KcsY3ZO93KZFVogBmDE9UB//Dpu/
cZ63xyk0F3iChAwyNvEQRDz0lh8GjQuFbWE7COdBk89ZZYzGCssnrHl1uvqqx/EQH+Ut52Tu6WXQ
3YVKkaM+61uPbhMHEYW2/d4ZM7gJfxpj70tMh3BnVUerX0MO3TBO2n4OWnf6SwS6MmbePNJ9ELqj
WyV9EaRyYZlKM+Djo3tbLzm+uy9/VjZlGgWG2eIj/bB4g49AZiAvcca7H4r5zxFLiAZz/UqumGdy
PMqkI8CbVO1bhB9NppzbcPzeGrvwI04McyK3dohymiMwsJamqIscUFpUGesZIO33eI8N2SSjfkio
G6ph/B505mX1lORxiUHYmIaPEtAvqdbmzhnKn8Kao3Hct9ysVgjAIxefgX3p1KsKt2cJpC9l65n6
pdg7MMju1nljdqr/uWDR4BRlDNnXuCug4yT8YmNynVJqV/aRZ5IkiFpMfpemWdSLX9zZTUziCCsR
8hGN/Dgi6dBhO1qvDfKSh3W0Imc7YtdOhEU4McbOn58zKvAEGdVmUm1wGqrfHW8cXWG4u0palGHa
PSb+WnWcOIG7VeuIhgc3kR37Qh8mAAn2WIbDebYmpFD3eWgW7OzPzrLiKfN30BseWDUuP85N34T2
1sX6y9HDxSYoIbGHk20SaH6+kzWp2WYJa+OiF1OO+JfppssC6fo1izc7CpwEjKWQigClCLVCrewA
SHwWHTBZ6Gdxxtj8ry5kwM/M3NvpI337ACqrQsbT7MwiGBRfdQ484nfBydFG61Of8OWW3/hJlqnU
x4fEgFji8HYEuTxXZmRsluK13Ho6zGWqf+tCJE4SEkaH234P6C4NHD7SHhj/fvYs0xkJSAyXXK/F
+uUnZKI37GR+/aw/d1JA19RnViyUytW67Y3xu44Uklol7QjELROgLtqz9xHx5/wEzWeO9Nx4zYpR
bhIvC2GjgsYPoIWCp5JwFTqMV1tTn9rJWFYeHuP7gLuKIuOFJopicrR11hIA9e5UsX2Fq8+mzXvg
zXYnCgxiGxm54vtcneFt32nZPtfZj6tc6Xf+vmE3YcUpqq6kTwOk88AH47v5S2Q+SsttktnTrIFM
eRmJaVTt45Y8P/nbq+qKQh6f4voif+Vi4ACTlAYLUtg977ignHufNRuzGkXtKo3Yd06Z5j9bqnNQ
MTY4SEaqRxbjYlzRpCc9TLLCHyvu24WJIS+N5wGr2/Ep2zcgVsMLog5E4J0+LJyCabOKNNknla+P
FSc7IXT0OG8JFB6+Y0eWKgYvdU62bbCTVL0/t6wUl3XAXMtqIuUqMgsahnKWBWKxtpOQmO6IWYpY
JA7h26fX4he6GrFo+vuDbehYyf7etj29sT1LA860VkbU2mljJ9qtK36vT+i3IjcfRBuqiQWhYvLZ
VgMP9X9gNIIsOi24ADQebbKSZXtDMRHNAGYkGEi/rx+2zAkA3KK3Fx0U3vlWV6IsvXrunhPqCSyL
/5SkkB95r4GTqYDjtfhupPdDAdvwzxY8UI7iYkP8DYNYld6BHP9ETIxyKQhUM7UQAq1jaq57mOdo
djR2q25KsM61g3kK2hIC1WtBWzEYFzFZ2ysjTuEVmTki8itIxqvhGzOZ50lQ5LiujWlwDuTJyI1r
w1Z6nmWvhrhFkPSvVmelfQrx5n13mzZt4Od9kfsUEkpFkvly3rp0BeXZzhkFhW5UUjiuiljp6TYN
SSmgpw7CEU+swY+eH51QRWkLhimy4mDOy4UYKbgCY4ciAxwvsSurAKIQhr3KnVZ+mazZT7AWinma
jaiHaWPa94NxW5Lpj6r5DF4qST3ICCEs8+1y80K4XRTKnq9tTDk/ZMqNg7f/JvEy/0UsuHvWdS90
M8dVGtm53D0avIg1xGjSBd/8lEOo9fCSR6IQruS6/H5pCJ9MqZgKy0dpscTY4QUONePzjoC2XhIL
sQKgWmJlgJS/kLixd6XkVraUNHltO3vG1ru0U225YW88n38tlhrACm+4aCd43w8pFEYG9Dbqe0BQ
S3j7qsvnybr5LyxIszTI2t8prqjLO3Ofpe6JLY8AjKO+o7Li3RWBy3UvDo7FqT+ohEsOmNpqdRYV
RuzsnSDvmh+kRQM4oo8++raIj2bgeKKQ+rUFp3emKRrF2wEGKzH8YyPVg2YbCCyPdfTZPeMd8PJL
Na4SXiKtIko/4BvNrWfDNYtHN9PSrn4Z4emLSEFV56g8IBBlYfrQu9iXXFyjwOdzgUq0s1S987Bg
GSbSmcDMIdWixGe9Fpkun5BjmLGtcx0H7ky1LhmSIJgYDbAbeOI3bfHzU/Rj/kU6ZqskFQhHmJk6
pXsTNeVOKB/AkjXqyZJ/Kz0Aay/rbTCqEBMEtTaekvuBrYHBompbNigDjcJ7ePiJ4nHJD6WqMn2k
8ghSg+B91M8coVwjOFJ+YYoE9nk5iAVE/SZORhjYXUmddXFYuhIzo9PY99JbgvWHbQ0ff4S3ZQ/g
LwtLEWzuTlj25vSeMXjzKwrAJNHn8lIUhc7Yss8nXuCJQJqSTZtmBrzDi27JGj1me7Y3x2u8CzV/
k3LSvEW1I++D1jfEMgATxtdPrJ9ffhbVKnSjcxb2wqpeOZZApn4s3ePun8VMcA6E6XzPc6irwM3w
vi0Hm3oQri9HEzxYKDJNwu1MSqkmRFzuGY1I92LvONwe4BhSRsJ6bRZxSXX4DCYzk2qNvB6+GRZ9
48HTNKMUjLb48OizmNwZDoh76cHRwG8jZhNCvWIViate8wfETqkPv30IDeRjrv2frvwB258QlXMO
6q2Z6xBQ7uYaQQY5IBg877tcmTk2cMfco8qFtlT0l2gk0h/nca9IetlvA8lrVSIX9PV1/dZCETc0
hW1QafCoDEFSYF12Bbo0JnMgGwrOmGvAFgMrr6yeDP9zgd3NYBFoZHconzedutveDJfEFfcfUu++
EzOVr92GSjEoVd4YHJtRXhd9G3ERjpcxc3ql4AQANqIYEtvPSOLcQV3zctIt1xzW9ClVk6DRcp1R
+Mo8FOopZ+hV4fJvV0LgAkwNZZzjHT7NvzJRISAMXL5Kp/clSdju/6HKOfoBbyVEmSJ3Q2DroMF2
m3V928L3I0z830CsM6l8EfRnAISzqfadSoGLT4IN9ZgJr6bLTA/glIvW05BsjBWI8v1UPsYf2X93
Qg1T0geXRK75MlHgqqLa7aa28XGK0OW3MIOtYw8ebhRfB+8gNPAkbNyTvehmafWfimaTvha7r37+
U7p+5qbUbAU8U+zJG5jB+7ryj3W3Owx55NQ3MXXS5V7TTZA6Z75U7W9JsXIAeIggTdBd5wdMccQ+
SFHSHRfCka0IfTKxzWqCc2vUzTpTFF40rOEx2kyxI+hUTsLtdDj+V9o2wS/kFB4tLxLOO52LKOH8
istAoKGv8MTI9Et5le3NxqSQpQLldKTdEbztfwe+0usUniRqk6tSB0Gx6qvmHv70Vuy6ZnEGBk9y
vBj2anJjCNoyh4UBcNyF7/EGFfQXX6X3K1YkasSlSCWkdw5+SzeZpPzLJbX2N58b5w7Cg1lA34Bi
os8dFQEs2HKU3L7JxvL46Q+MS2TIssYkLiAMp2i167kt2as2Hi60T/swqRurikM+QhqnL/nzc2CS
KgcSqdXXeClBRmUkk7eB4NgfvAm2upmqHsthIEbzjI4vxvVF2KQRifYi9zvnOEHhGy30ByWhgmo4
h++3yZ6CW5F7CvXzpJve6cj1/TYXi9g6BCQFKAlm0E8HV/tf/sn8Stx4HRZXXgZjiHfUFERlNB/E
FLj8WBrToZJbEccdlvYlV31FvsqYbf6YolKJqDHwu7BtRfU9JXZ2aIs9svr/6BUS3bdNubbPR9ef
4anZs/Su+tt8JUp8Xhklr8jaggWdlo6hd/NOCEAZBDNVtvXu4Ht7EqVCWB6KLDQUEfWEAx8l8fmN
GaPyZtUXp4/7Y1a7d04ccpASf1g/6LCy0+IceDRFERXjDd5bRx4dUmgv4nlw5Ze4xCOETEwSUdHI
1yEosY00PFmM0cbCN/8KUH0opCpu5E+ggIO9GNdnjmQtx3M8Rf+FdteejCeomDlZT1CNzQSmNJ0I
wMRSho6/tY/P52gcpgY0i0a0nMOo9q93RV/cVNHSicyvlRYz87Qc016d2CVIPhkVMUg0zWqp954G
0mWtRloy+AGF7DYw28dZ+VAOn6MZK6ipW4UJndZjDpgKLyzaVSwS7EQEcOyK5yVlqihWiN5AvN4l
YqlgjyoeAqshuS3v4tBKEfjnc0m0ewNL1Fv/dE11zB1VB2IYZ99f4K8JWKeOvECm4FvvFnPfo4YE
DGOLGNqPiT+NaXaR16zh47xRaDEDSg7rCaFy1jA9bZbbreD2WrMgAQUSvGpvgcxmwM2IJWozXWQQ
n/sUQL13/4k78f3eGm5fOJUKIYeoD++d1e7IKAcxYIREfW9yzfcmIYZhfW8HYDTDf0EXQFraAACo
Pn+5ns0ybKsFPBCO4AE4DT0giuKcl2lO6R+ivgy1DcVy6KN/vZbekngYNWSMPZMWY25iPZaw8Cy4
6rLd2Cte3qFbNFQs+1KuTTAOTQyuKtjgGabpE+DnyfO7j9g/NODIWZU/8ZjStfAx8V7du6CHDzpc
+vFSNybsMXhd2cYcth/wPyL+GqthOR/r82AnVa1DraEpYePtpCOGtd6bvgII9HM7lJaglXh4axpA
R2FibjoOnMqDR8LxdZjjdpYRlHscoXcbYB52ILVfTyCZWlD/bwJ6GaYUagsT/opQUTNlhnAEHqba
68EKjs8IiDIQvcKp0iXXFDi0slhK0VbVaNSIcWhtYLZrzCgvXZkfmddI6OitqP/qCRUkvvbrSgNU
q/aj4fRWAKEP9xaa6OnYFe+CUHBLff3WseZviBbZ27YFVfBbu5USsHPpmEPG7xyKsvFEj2e65nRR
WjBXZxBi6gUA5ZLtDUKRQT3ywOvqSoNbuHXyG64B8sf0iQLabTKk9Spd5DpQyUMBBAvDV6JOQHjB
4FbTjvEeByv2mmaooP4twYA8HUaLHrW7d25pIlsUNXpe3AlRz+6aGoLMlperau77y8dx9QH9hJKK
hRQj8MdL4gUB7xUaepnZUuYZpFwdyOzRSEz8qqnWjznOSlrP2S11twV/P9eCMqsPEHZXYVQ08YwT
GQKXPchKQaF3bCH8RW/JLqdI08E2hEFyef8DWbn3jr8InQRElXculq87ZspdC5BIO6LFPLhZutyS
Y2J0cfEmg8nrLkuVE+9FMRxFPRAWrGpVMpT585Cyok2d46C8GrJy8uZpnrN4FXZWW9sJoUL3lo6h
lHvrwn8Qz2Vgab94NGNiCz4xomynwE9WXrM+ygTu/zbXldCYF2Yo9lSQzbQfNaclmtbD3H+nZYqS
ZDOJgQbdhY9NRqHfqx61F7BjO7o5vKAUj/Gv6wWd4DRFqi2bENOp+iz9vWaR3dJ4ii56xMm8nHAF
zvfOTQO8EQGUNsjQn6kJ73YmiRcBXcciif4CP/JGzZ5SjkIJIIffaRKWdlocqCmyiPih8vlklihj
eGg2pFCMNMJ14DC+fny8AsXbB7GD8IeD0E51kZ2rpH63lNIAOMfF/kY0Zgt+4bNRhow4IFnBjGpk
Q3u0PMaO+F3J9JM8CcLk3wsk8tDQl/ddcemSB2bK05RD0tuUKaZhSWyx8GDgP1OlJsyvc1ezJA9P
/HPesnbZgpjdNSSYRZgqTT12DhxWfyTTY0OtYVLt2KcPCuSth2yHAzA3Hkw6uWJBQ+5w3iOt8d7A
MJgpoVA09v1Inv4emLHuPC1IKjX4xGOErL+ZEoo7nIAiS97uy8i390id25IXaKq/mpPg72w/zU6x
qGZbG/KHa46N4gQMwxnhFIc4N2kxvin8qXNl212A/f35ZBkRapue7TGnYyh3ssExhbU47HSnZ4sR
mdFu6E6SN2tWCP6CgKCmaqyhFr6Cdp9RCby11HPpZMVnaTd8ZRL48qDZlIGaTaXji3ihM9Ks+UTs
lmtYXv77cp97+9sZ7Un2Lu7+nT/l+ORL4/dd5wlIfcY6Ahj6BB0tS9TG+fQxabxXVAp1/DhGpTg3
q3ppGBFcG1xuvXByLDIiCSMx8eyCfgf2aGyvCeVfPioCI1Mp6xh/CqfmbpgXZOfG2PL4D9FlmuTH
Orl449mEDQRj2/mBQNohEI4LugUMlxTH0bHy8vln6qggCk60+O6sbxVKnGf+uZ2PlhZLXvzQ33Rw
1SSuyUHaVYqRx5p85hynzAoFrulWO7GflkH9326YOsw8sqfuyOAVseebKqoiGPdkOVORqW8lo/0Z
i6+cTnZxpCNeYr/3KLdBTLbDg9EzJMlqRlFdRu+O/lpElNNA1GkQCl0FI/QvHASgQyblqNyDOvyF
BKjGa+SzwwZaRW8cZy5QBZH9KaCokPRgwlr01mKfxgil7ySprTJinAV9csIgTCFy0MgY3zwdVakI
aPttKB9GhJNBvP1Pwl3jduOCqKQuJHk3vGv3fY6w2+OQ4kFI7+fhvBdot9MgzZjwdvSwCeVNwXAr
KTGnalUYCZ8llJYQzfXkbOzxbupA+fPme5S6EJgLM+po+szZNC4Md+WURkVAB45KGP2HYHEBuTSa
M+u5mp6U2aIiEa6sfCTQDMEh1kZ/f+pM/AHCVB0inWFYnod9ODHD45jTnwOrLdx4Z6ed4g+K+qHI
PjsIqkC86tElpCWoloNLFjbiZXUpyYzUBAcnSe6gyBSuKk5mPNTYdvcCZX+d5bvmzqY1NPPEmSyq
4RBymh9cO8IiwSOiSeyClPhs4M/jvkD+mq29ymSWwlpZ/VWwIPxMt700W6+c6miGmCZozP/0PgvQ
VljYBQtGOh2uJrPw+nG6KZxmLI1uPxw5aTDm1DN3yKy994bWhHwdNGQmfxPRggwWt6tUOSTy19H2
m+qEqrOy7bnvB4gwZgPGnYUD4Ce99wL8B0WAyPQ9S1kcm+dklM3a3HN6GXRiK9A+G4aYiZKnnD2I
SbbUpF7/siMqhDZ0oNwHw2DjNztmsk+CL9i/L6WoPXwCaWMIbtc1XZbxr/mqjRat811YJkaDjT9T
qQwGqM6tsmp72Mhi1Nt6QX0tt7e3/kq2cXmUEJGiUzn4OjBGpeiEDxTbo/XEqadq0FCH0MPUrl+j
nWzjyAbfNpskt9fjVCIVP1JYpNdFbx1SoqCx88tDTQxpEM71ViQmY5ElSeNA969n+ycuOOgcN11c
sNWw8QWjHIv1/zC4wKgBOfKBhet0DJaR97N1b8w24fiZ9qyWWRhUL2HC6wuz1632/YguXXnNzRRs
2pTbly0ipvsnRqqannD+XWpBny6bwDOCklVIi9KfvnsJriXdTH8wA+/BrfMi+ES/dCcjDA6H/VDs
Gc3PPLFehmMFC9PkKZV/nVBMOnppv64Ymdz9EvIBEv5b+nHXNFbv6EWVFjO0pVUGlg/m7G0bnT1A
s62uJVoGydlVdojcqFQsr49w/DWFiemF8kk5AKHmH8K0EQcWzraZrXELb4Cnkc2dqsv3yf1emx13
0I0U+j8w2I0TRw2QelQtoDOUy9k0aEvjSLqEOarj8d29s5OU9jOLqOYuS6whbWltz4RN22ikLn23
n2ZCb15nC/gTlA8r19c4KQguslaakzYPnnP20cmhlJZp3Z9asGwHGssvV2GoecS+YM3brKT/wY0b
6ON8N5xuR+Wxn6sjU7Ocda4LngYuTq4VAmOJ3XM+gL0OdDU8Hr2uGwWRyftMTCNsqhUDfuTfPfMJ
j2ZtCLBYRLpg+oGN/KZiEaACkR/ozH8ygGNvmaCORE+HcPIbmt5JbmGmyhKR70uS+nE7L8Xn7lqp
JLUxrs4d/9+6BPBX4A246LPZudZJ4+eTxOdGg9FltFEwmNIGFkROF0bd4/DAMaISkusvtqTYLqlE
gw85tOmquDMbI3TdRhlWWmzti9cIpVST9y98OaGhfnOnSDtmvT9CIjcHrzOBd4kLD5BYwILTOBsV
dTr6j2YYI/d1iCe9tfyO9H6wzET6JZfdukmc2U7pK29EL7RRQqzsv2q0e/Gaw4SuRoc9saoGPxle
vpmsvyiU4xPvj0t9duPXz4Rx4Yo/yew1nWRwgLZB1Rm9ImmEjCKONm7WcaJrLQOz1qmUeux+EgId
3EHLIohWxRZt19OKmN0kn+8lRtzsSgIsq4zTTmHJ2+sbOmdzD/61rprHhmENRUI03C3PooKarXoO
43fZ3Vpr2u5qpD8TUi+YYhz6wrx10GCvtLSsQEtAYxYrOldzwtv/uNERZ9nWblfe0V3BjQ5yfykO
36HoHZrrqVbxWOez+kFj0BtyTvRSEjXWwKLs5Ht7ZQIyOB4IJNr7EWi6f44vLW9BuHSS+Ki+lneD
6fQ3nJYkMlWyfTc0t6ZqHk0Rh+eoILTG1ohwBVUpn/tqV2dxcRMvyUAdTJ/RbmhONQjy2PQkjnoF
S7Gp8oKUifup89guy/fKTy2SCv9635zDalus+eJNz4gCtlWkgMFLc2Nlz21kTySUPvQ9xEgytTUz
BZQDusUXe893X+oorzQh0g/OfIoRLcOIrUjCTmShUB2Fyfp5zgAe2v6izXfBBGikvYNtjxibtKHp
GT+5llQ4o0AOwoESD+QXXwtOAkFJnxpbAqjEiaFnYad7E/LhzfvGvNXvn2k+EBzChmXQwkWUVKW5
zrxWzwroxGfUiFEps3Mw+69WCos50p1F/hs0ZCXE8lLM24+QbBdi0zl5VLYnb+gdhsFyT7YjkR30
xJCFckXo4EJhhi1zMblj9fuLU6ziK2ggmiTW627YbmvXkRL+jJYOfFuHf3rfQdrH6SBs3VxdEKJ0
QILMTR5uohNtBySLlQbXUN5or3upNeZ4ph33Y6Of47oSMMhQ2XKU8UanE0NiTJcwald9KMt28SPW
pgAJnHjzUbZ77u9/fwLS45YHzPM9+/w+L5p4W8ojhit7xtWCtoLWqDx9tW1Ewv9SrrEoZnfQ63zP
IVz5Tot06yVrNVbeb32+fspDDfH65fC2rO4g07gVbScMI+JCEAlwkLdpAz04HyCEcr3LzsiN0RSa
PRO/BmMi5h4epGeZ/d7GiWK6SEIiDaEIZzwB/LSDBNENXc3L0KY1uuTwduwqTChUHo2rMn0Zm51m
HAPfBtyYZb+Ys8mjTJ1GkW16Ritr20YJYTEEEYAi8wVD8zqh2iunbP+txmvW/433pJOLEGJIgwgG
/K0tv6MVJpuU0Rm9bwhldnL49S0wEOCWC88r/YShYoJnq7dXTbSvq2mt9rIPyDA+eNfS4ja2Jxc6
WwtOkoLxNNK8WEbIosVAjubuMIiOnTMH22izIikIUNjT12V2ZrUQj8YAO51p00k+OybeeoYlpWfx
mlKR7g4gQIgpiaR8eW1SpxbP4fJBzuIAr8NWFNazfpu5ZmDcA4MbYjAjLskO20+wGk4+SC5EjT0W
zFpLbX/3MPRJScv5R4yRUW1KCBkvw2ms0oWB5WDHBAvAn/HiPp2VttJukv0kzkZgaMzJ8NLFZshy
1vUNAJ6qcToLoy/lVKHk1+UXNcnR8c0dlB3i53rKxgl0RNYgvlgXmk4Fr50+LNpsDhQDMsagOzjg
bvnaodlnX67gq3L0pvP3I3YTI3DfVLNNcM6OrQwNRWhiG8n6xbdyERaCMJ/cDERG3+1jNypwmJzM
V1wFFuoPdpIcYaRyvGXVqfxvcl9OZzPpxs+KaoEBrzoRy6a6siuQLYzSrdK4Z/BO5XrobzSdTHXx
tX5l4HUZS6somQBex/Mi9LuBYavi8HUKtFsTGHSsGwzdV4+0kaILpOIsTgW2EvH8EhDRd+L3ECoY
sPCzHHYrDKUe1VwlvEFa6NNJXahFIEC3mz9GoXJiN1Rf3u63CwbdztY2WnZgpduaUjlzWQuzxTjM
RdPGhFOr/XqIDLQVcFgv71GqMO6+GBRyQIY55dpckTeyGTTtVIruhxB3NIqU1GvdtKYXjOmCoihb
gztKdNF+P36Bcwk+3KQtDLWOacAnM7UysHrPrh02Wylpaw0ppNvrXWFOJD63fZv/FIqvlrkufPSF
kk/X7X1cRZOu5Y0PfRJIfCkZlPvGMYOPArgcx2pt35HbT0lUwR5FwfEVNOKy20o5MX7VKNKIj8Qy
jnABWhJ3VUej/MuVuFBHO46fGrx0bBfQlE8iZHsjPKScmTXCv/F8KV5rQWaSOGRUrQhG1SALi2LH
9n9GsZu1N8wVwd6wDuxA5wycMiiNd91V9hJL2TYhMfXXvWiMJV4jGAXxqrH7XQIVQ9ks6PTKNIKS
lL9GEbErqf2ZP4hVPoHkp4cH+YAO953Ff3UNmdXyy4hkYDvnOdohLngjmELkMUv3Ah1GPXoBmc4e
mGLRpdHZ2zf1tBZVwfTJkUVrODg0CIbwHJyEMNcG8v/+QK52hhFx8v6r1uPoaZjIrRHIgM5AJM6X
dNAeiiylZcWH8A5YeFDBd7e2E1CH/2hR9zLv5K//+sj3DRCYF260JsC4UwEHaYBEtmqZQjh3DHub
lK4gcTeBkTNV8HFlDL5Plbe/+P9iqcogDiIOEndCgpCx082Fqr7lalukhvJHtti1LvFJRI+N9soM
HkGigCpgr40/gKtB92ElNy+WVc0xLAvECVSM+Oe/xikAnUBJQ1JBwhC0jrrWqXWhZ9itfZRd8fzx
ExgNji446J1XPEdc2IBkYlGVsnRGBaaG4qPM2KxTyL5htfEKgvH6acrSUfAKmqXSVibycmZRz1tH
TOdv7xk3bz+Jy/dtqcZQkngo84Iz4znBn/B9NFAyh/MvoYLb4H3i5ntzLJLqSHFfjhT6ixNaaMA2
bgOiCVGtrxHptlCflOUbwV/N5bZIItL2Maxw6nDbBd00qDauTFsyxDlh1ME1x7N7T74gAD7LCS92
WxkOlJvW/m1hPo8S5H3q76oUv0vEuf/07UPywc9dBQtOmqNO9JSSzG22AoDSEQm/mC5zJWVVPve9
ByFGStr96uct+HPdOqO4HE+yJvyL43kOKCcBcQ21nHNaqxxH3asHMH0hIZsIUs1rpsRdfdjPR96k
Y0yrYSVRn6FJ386rVSV7vQ5hYnZeDt/27f9vMse/MhktDMmQ4AX+Z8wGJv48JqXMIh0qJey9KrLP
9zakLzhdZotBJXAQpsW8zGhhO7nD//0JPw4ggNhVFftk2U8UGpwoZZerhhZAECUeAqS3OG0m58TD
Ib0sq07VdXVCfenlJz3BOFU/D4AXt8RroL8hPYS8EAeqpRfsjPExjZ1Mk+4FK1SfzFW5+lKII2Qa
2+4bRZhH8YNNaxN7KHGgHlFx1B/jO4xpMCfIF6ApOdglhEzJOiNzvDwuSN4uYpuc8KVlZl/EdMDV
lh/4a6biXDm2uJ5eHX0sfsNuXrrUkG6Z71Xnqxcdzd+kjRiebRkkfoug783dyZMJ64GsITlYOhYb
MKYRo0FDd6QASFnWAl/wyVCYYmf0NHF93MzjQ883rToA25xL3XkYBLi+9MpaaE3sbnvDdPS3/zTx
ciooLLfkTSq0hR4mhKK4NC66Adyl68j4w134RnwJLVRHysYo9aWYiOwMGkvqNB2ximdWn/VRsdLs
totiu+tiAe5Ld4F9NjxJ2DblsfWM55zMAKfc4t+ZnrIny64ygHmX+ujcnUQNEb+zXIQPwwHK2brO
bDqdyKrLBT0+WFKouJ6YmN9wUdfnudLt92TiYB8fA2WO1fuyY1i5p65TbqyNanYEiCFsMLKoxpVT
RPth+qtU1yHvjNVqz6pt9dY0ax5aTlShrfGtHW9qYk9L4i8+9PImYEWoMHTxFyyjG6NU1kVlQgNo
UlW5EA86IBEq29epVC9dhOHkeRuFSlCE3DaWbdnx/QRm+dkVsN8xOr3kk5N/9tD6QaOTEKJkKvnb
i7rT8YfoVVGpHNWJC00NUI1xwhxAatIj0XCDmh0KCnbs9mWZ9aqGt8BWeLcp59oerIv16fIC8xSz
kIK3MdoZ/fT2dyR90kLpx5KQ7J9+FyEpzLSG07yMUeFwwgqzHUY6niOmhF8t5/liR37etmgvIAD0
0utXlVa06uoHNbrklKzKXRTl2pNm9ZXWmYMZgAeX8S8xcqGdB2ZQ0zlWwiNvI6mrZUATbUYiiGgK
wHh+u68BX1SUj0iX6/YBWQxrfg0b8X9UsA5WArDTq4r8OzlPFc1QJScBqQ0izhX6dv6qyX0xyOyz
YBoSoUjYgA1/MNiXwPm8ZeYijf3awaO4tD05nF8n4I6Gfh92yFjkLWhyyktrpqNrU18+bvrF2fct
1PZjCj85VqC41u55DFHkUQ3PDFqmkPKfJAtbsNwogGsu+qUr7zfhc5sk7wAw+nFsNCitQW6wH014
bmGutMPRppyTQZZ0nl1ZocyN678J4ZVk+nttCT9BKkzXeDAi5hV6zX0KxS0klOpjO6io3NPA15ax
v19TaTnBbyOLzEabD6IeQ04iKRgu9Nwycrr1kJJHThfzHPXqKYUZFA8ChU8IRopMPF6/R3MqO7s5
H1q/KMuX0MhM+9DcBhYh7Nvws2WmH1ngW76FjJjVtlxT7shxnDyeIoKwDPVTE+ROWKffLUjqfSWi
rGjFd6nh7SR/nNltqVFj9cAU25/0q8HYySz3EFqRvU4DmCbWcc2VyDWZtQBHicyIl64xAmFZILuv
9OVazt220D5AJiRJwp9Y2zceVz8Rve38ofeeG8LZ0h7bbzBx+iwaAER1A8BCCqaDwFTtYePFFSq+
2vxHB4OdgfSB8X8iqOZCUREIK/jQhg2nhVZQcDfPOc10R2So2grLfQ7aPW9svaw4GC357x4VTIjJ
GfPn8aUnnSSejH7Lb3mZhkgTtveggpCurzBix71J5HO0E145UcJkixHlyZsQc6hJysqusZcvVlth
aDKYGjnpNfVNop83d2t4xRJWZFXzYkBmzFr1iLcdbUUgoX7VDAKbtxiZDNlESZ5h2y/SZGFSU1nR
RFrPQuHe/1MAT9mR/WwVoz/lGaHHrtE7lDPcOf3Dz9pKgpSTUjQUdS4vXe1gC9GBZhrtsoLK6aB0
F27ezFlLoUEMYIIqwc990MEwXnMtdkt6Q9leUB6LDec2UUWz40IWrPV1zSwiIgIsBIZ21dIY/pVo
+DNW9Folzl9bYd6SW/Px3Ex7nTkGgVXQqaQyhrl9406JgvgRCIc5E/RZdBS+RLcTCyEeoXkKeYfo
6HkIx/duUgywx1wxYLPa5ppOQYXiat85EfGKrrljEYx5t0hL1xyP+SlRUImGi3Wsk88coVixBN82
S+87CmCxUP/cQtqCZTPeLSr3eGA/c6OmlaXaaHEUlzvCVbIw4eVXGcq+cSNZ1RYMjhnljt7HDp0i
i1pN+a9LTi6K8LJuMUOgEvKeEEDMNZqnxRM06sr0eixFUoKhr9FQVk6sMiX5ajo/n1F02JwqyXGn
bRXwyFsHbEt9wJg/muWc4DWsYHjR5N6iwHfeW39D1Kt3KZ290JVK5McMVMois3cNn2FoCyb6jUGS
jM3N+vv3ZElJAaMS5NVZgMd83mQ+l/znswiEanIYQr88SWNK9eE7GejZx8HGW4or+Zn+0r4vmMOp
AGb7iYQc3Rv+oT9wH5MjQaWoGYWCXLF9TwtOjUA3+6A4IXR2BCPOjOa+QK4T3AlxEmjY4DRn9oM5
ayL3c+WwrV30HpV5ulUpVLj86FPMXucVNETvWZZUV2qcaPOmdZXsF0bfedvT8IkNXuLqZPUA0zDx
4/gk95GcSiAdlqz2osM3ifVRcH1e6oKcZbH0UQSzZCxNlhgWyAGV7VofzUJZacNtMSs5pUpjzl3C
cBwkRw5ddn9gSxaNjEqjjPJGq5UE+a2Whra+jf5gBuej4pEkBrfcKJbv2+dOVdG+XcmK4xLktk3T
s/ZUVbl7oNbcVPpIbPs4c/l3jDiPT+SUB0ULToTiy+N2HiqteQKNHxeI8GmwvEtU5TGY90qVlPce
8d5PVWe4P57n46+jY8jSD6Xr8qurjA9oyCZc7xKzjMsMmsBjVu/3i9hjH8RiJY883im+WRUNDAqM
OdAShrHOJchYzNCBEHo7kN5NIMfwJbpTk2hauN4j+PhUOz1oKWWYPkA+ReAPwwDb8F+bw0BqaqTe
sgquQLmzgey3Cl0cK7NCDTEcLCzRzrOl2aBZ27OtTYuFGTszpJx/PpOnppDj7ygY1LejaZrlLFow
SUbPCyDPBVroSIBaLUOBLpz7W9tXj8//n/b9JpbD0e8n1Ey/v7tpc21JCs90Fe7meNdGZUqJIsZG
dCpaUwXKIM4pWV0BUaQi66pvGpvgTKPdOvu9cqWx8mE8itz01nDTGsXO0oFG0Wirhb9DGkYCfGzZ
hGZnfUj1lJ+xjIOUW2QE6G53AFoDjAxCRFqACMDeetAuaQm6k5DEsQWJTTplRs1QfsYSSsMXlmAH
9srn6HRQt9V0cfjkWo5EutsV/l6p/XOhDvd1D+/WGTbR4atSLgKe0CJuSfk8KUpiHv4+omGd0m0s
AVsJE5MeyAIcIO3G/FnAMEy/kz0aVXOTd4pFsYFUBGkXAfzbnAMBiCuHpC3EXvspLBUn/IbO+/jQ
R8CyHVaspazg2sbXDYqqBRATkypThZBUeKAzBDZkKLGLU3PZuLWxNzqoHusTbu6U8sSrehI30KhX
3VCDXhHXPLuWj6PYPkppjHRnWJG5KW+14w2cgZJCpOARhY6x+21bvUgkjM5dPqH3q5hpgiuxE/0X
+oAW80chsRMklnX8baBDR1c4pEYZ10+Izf+nXNkpx8N3MlT1NFHYtohDXQo9WIwpNab60tP1g4LK
z7H9jccIwl/752EwKfFTolqCN4XLg1sHQmLPK21s2FV3geum3qia9fvLhS16oOGfSg8WexxiteMq
WmmwYpP8CMkeDyrGWMfK0Spni50NIPt6mpeEEdVKJehjlKDNOwr58E2ihPGsin5MJ4hog0BqzOn6
BKTFQsfk2cYCXrMAiFFEhBSSbld9flbR4KGr7mEmVvq8bHgxWs0T+mU+K+QOsj/xUvOPqZq+oGVE
AY2gGxCQfB7GYzU6pZ6A5ie74jmwzoVNtMhmTQ34HmsFghZeplfCScnv+oretZjcbuTe1R+SIhm5
DLnGUQrwREcyFi5bkaS9/QRVB70TrzEO7uOYqHeJBZiVvU9h+oQFxgr3oYPG8R9msxLBqiWdWkv7
bung1OoY5Iubr60Mq5EvtKga/DIM3s/4aATclQLiak1uBNsK7or/COD++WAxHkQ5LYW+XugapHlS
59bPHniIn5DLWadh8KCNim6xfFLWscxqaVqjXhokEoO7nTb/jfTyBmQQPXOUtLyOwtbvvIkIO1x2
Ub6YCWYLoqVmI0eIY0hd4+LMeFAcyEx3rYTbbznH/bBBu8swoHHrSpppXrhm3axc9vXz9oAP8wOZ
YwAYKgBilArhWl5h6x3Rl8oi/bTWTpXzw5NSXjnm5Xb3t13GWzjFh2ESmCdjGGKkRw/vdQrIQFIB
wk6um/qKBd93LvdMU3Ge2Vv2p5y3+w7aJq3yOy/qP825IvTAOw1Vtd9nl0Xjxiq+Z2tznp0FD4bG
p0IWpXXYH2/zEc7LiJ3vMTBY8mnmihl2LyFS38GHhRKlQhvd0HfqyWEfOQUaqw9qsEJL6l82dDNs
w78DTd/u4lOYbrZDuAb46HT0pqzfZiL+QUdfq6vWPLIdZGT2JcbYKsNkp4y9I1ixZPOa11YphMAr
3QcYgGBh8tajHgYAg7r6mLFucSt8c9J5U78Izt6Q71k3AI5SkH+Qfacq1cLVDMW6+iBb0Tc7MHnq
RWeeV9rc5qy5N6MhkymAlkgzLReWwFaWNIDp/ByIbXd4ANy5T4jbBTu8e4TPp3W0sDvuHCR8YIhS
bWMCmWpUBXylem4iv5SpaGbvZq67ZPXvCkakiThd6AH9nKaFbWdaRdF2y0kMx+0GzZy005Q1C9nG
pARHer2sJZSloqT1DQ/X751Bi7Ceqg7SY5H2+kfZEyLZetxhB0xsD7XlDZ1rXNCwjLOXydndd8j6
uAzy2PtKUdPnamZdo8n+xmRDuxwPa5xHMCnu5C3qKgt7hBoILo24x73NsdEkN/TmfPbmVhxH/2ZW
pNDqAuWO4KHiu0xrpb6H15qpCKD3VCsoEGM3rzZHFmMOZV9aKu5TVv7SW29zlc6A90BchOzf4jEL
Ct2pzSnQ9Eck9OhP0MgoEI/ba/1W0DiD1n7SwtvjqxEu66eXz8QfmgTMgPGcvINHiSnHRNhMeW+v
KSm5v/ICJ8IBh0Nuc97j6vfUWzgi1K5gAGk+8LfMhFqACsfJUzoaYBHM4bxItkyMWLGSHv2gl1ZC
1zmlDvWcbeQ9jE3zORX+FeZSQnTEFPyZF/Chm+Zq1CNEVQ61yNXIF6/vD9wOdlqfKN3nGrL57K4t
HBCHpfkLo3VZVm7V09kRPPc2tFUkshxl2ok/gV7OzqCXDcpZFHfQs8D2mySTiUNcnYGy8ihWZ6Td
OFk719D3Ld1ThUeoqXEqlkvtxbVUo3+TOqyENL89lcfSYf9dvhOvyOGr9F7B4ZsGBheql1g0lybs
xLa9uKChOun8R8Iy1qp237DokuAyl/CdwbFHfud8UsiljZpczvTRDCYA9FifwI4tjRLAFWOMSJu1
DUjPz4WTAiAuZW4cBsaRhVn48zlbXMAs7CQOOGxORSLnJwI/oQDVH5PMlbfcuczhJ0Y38SAcJI1K
AL3DPUxFiwCTKbOPjySleu6vYZMSCfQ0CrCBI0cccDt+raQTuOy+w8KWBFlAsa3daWv/abEbEEGy
i6oeRzCG1dhQ1woq4KRTNf4iaM8llr718C41jzG5Z9jM7124O13+qx1PSGARBpzZcQqGxJa08XEf
LkaTU35jDpVopa7KM2CBbQ91X+e67aq38DwMgG/rfR9tJdbV/COnkpPeHZWc2WH6Hgcf4D7Mlpsu
Z5HWIUaTdyaHs94nKOKDFasuEykbiauE7wUiVRj4zbL19S47fR2KefmdUKESmjQ4eNztJUoCsQS9
b35fcV4AQdMqY/4dU6rmtygtnbxtewxKiy5nUxY1L3PQh6RAB4VSfklUQXGrddyyo5FjawjcKm4r
CjuK/M5b0rhcCpfHwgIIWX4o7/7Vf7UKfwegjFjviN5YF4c0nXU9gDVnOSwvZRq0Jyenvog8srwS
/0j5P3diJCytMuxS59+b73PP+A7LhZUqxxRWtm4cwjK1YK2xSoQcNvT5YzLd6gojvXwAhdAjSWeq
D6v/G+g9oCp3kXhMgIP4oo2uv86NMXNCM2m4MPP1CL9CtuwXuUg3D+dlAJ7Ar1gDTRI0Ex7oYRtM
764FzPHgGDVk4IWz+9Rm3tUSqV6cWlbRut+MilW43vSdMRtiSSjRXUcn9nTl7ZXbwIOa9JkUDY2F
0VaLc4Nf/1xvXZO3P3kNzUcPjWDHvaZECHZ2ZBp5G69G0/qtvFmaXD2ctAP+ipQA9k82qp9cFgw3
FD90aFTuYj163guV3tO6/qEwu2rREahqPUn0aVjNVfA3vOQYnhnslsSazAMh6aJCDjl6pAvaev5a
JjxjxjW2o2+DEO9Yo2gvxYnufFKZE2DPxPU3rejSGh3LmG1Lb0L+DMx3qA2uEjBMCr9/kG0Xs8oa
xBU8vBxenswcJp7r2TtaG4U5i3ol1AqAX0LjtKPd0iDF32sqkUim9NzpNWwQTyX/V/rWeOIx3icF
by4x7u1oDdRS4hDLjQM9eWqIJ4GWWybE7VobzE5uYMGeaRzP1mM8xmWhTo1s27DGlQbNn3rvUwwy
ORgMKz5VEm8Cn9XRmfu7CNdD7sqzZWah67bl6QFeWM99ViDIK60hy7/epVBOK9EkSLCGG2noDJAe
gVdnWdGleYk594oIjemuFywn7TI/lrsZCcQQTIrX34Ufjqct27NgDLh8bd7IZdsUqEVlr3ebyN/L
orHrgJ1CcXUaThlV3M0SJLLVWx50omhMRQK/6M3sISXZ0nN8O4h9OcMeok+d4fC0lLbZq73DYW95
CYcZonCuNbX9NiUcs/zy6+jYKaZB05NRkVuiYtj3afjUkW8fgiTrK+p30866ehJSrE4AWAEeHULZ
0hOz7BUdg93uNZWLWVGWC2K8Yed24FQPP0kWWIpK/U7VCYVNQa15M8Cwj20l7mZ+2zzcsnj0mDBw
4VnBA4DOszoFo1G2lhHpe6bF9/pwkp9LqdnJrUK7BgpUYsEniV39sBbI9MkGDNdj3i9y7Dvm4V+Z
bQOZQXkSxMjcYMb74gygqlhmRy5R0kcB30hUHoKaXAyID75f8OYW5EM7JlwnZKAeerpcrs5KA7/9
mrgxU4bwVsW4JCQ2J+46joua5bQTsGBcI/KXdFUOIEce5oJ/TReslvWzELetF1cMgF9ViutvJH7C
sAgyaIYB9bIQyIrw2ROR2R3a0old5zhAD8ZGoE1EJcCMMHo7cc/C2L1hQRJmUj7Ljq0ofT6J/9W+
nCnF3Wt9f66bfEabp2Rk9gVzutKlcWYi3f35zolgWhzhMiEGpB2Dpu5D4GlyfO1m/V0pXgRcDAx6
J+TYF1Z4l6KwCgeaY3n7r50mLy6VUQhQEO4Hqc5yENzFyldNwRTZlGrux2J7MEMOmdpkxv4dyxwR
jZETJ9ZL7kGsyV7tPqnWofw5KiL8iJfSjJdz4h2xk2wmBIJOaDihe0cYW0L6F9TgbCGvEAhRm6/v
9gwaJPzVl/8K3gc6hInP8kBxC0jts6YMFv+zApsMwHJCKZ8AYbSEMDF5y/R+fR4aHES0WuPIUUHK
iNzX8fVqrZ/b3NNZaFICt7T1MvhS1v5mxynBjRDGhm85QozBQvjTyFNvcSbI1zXjqZcK2HyPjDQ0
UkdNGKEqcYaP0mBk6bmW7c1/+OpZplFctzEehwfnglZ45V3fc+RSVbK4th4bmhx1wsGrN1ZgbxjQ
BPKgDvMPVaTG6YFLa+oTrAKsJ91O61mUotLySR7xRZphjjZQfryrCNFBOSxwr6xCIVKn0Am4EmTJ
yd4Mtz9duP2vH3bV0CHnpzoliVXMgfZ3KoLFLQTFHxmcxDdp3WXeR+e8AOYHoP3gAsAbwyYwVRSK
w8hxU6sJEqZmVsiZ/79fKTUbam6/2jTovE3yXlLS4KkrF9G3AhXkcmRr0KVYuzaP6CJ3e3r+gxsr
zxxctMVTaT2TrVOpzZbs+SzUfhXNJ0/snOAYzM5NJ0ZDS1oSMqzMRH7MjlkAIuHWFyWM0kd6KXQ3
1jKBVabSm9U0WmZ+H4ZxyHwqmxrRWQ2g0NJd6XXEED3GBTBSRIAtKjF+iEOKcOFJpl/FMs1GZl9y
42KGZihRaVgyL65sKDufyPPjIZU7I3ekE+ecM3fTfUFhpzdMD0fLabaASTakh/v5re45JvTv1IeC
nI3XTOCtKtDtQD58m5eNFxWniC+TXKNzM3BeOiKU8Q78AsuPKlHTQADRRNiV9ysBDsLLwGLetHyZ
kr512/TDkfE8DHfqSUn/ppJtDlnLnPqURuf3iFAXEffhxfoTEJpp3Uu26C0H/nSj0Gu5DUdFxlb5
0qKkm1B3TaEcJHVzJBj8fs9GoUEDPFb6FqHk+JfDI5djipoJwEvmw8CF609gxD+5DEB+JqeOAQRn
JQVo6CNNzKJSTOda/P0aUQmWyKL2WyMb7OF1XaV9I3igTzY4X1C6JYCMyDVb6la1py/0lCQfvmPV
pFD9/CwqaTIHx42hs3L6TpyigfJokaXCPA8oQyOsPHpuBSaxMMyYqXv+o7qHmRZRoG7E1LgZsrH4
83V/haJkKVpXBHIWsaxCNwbVm27nDRBA62iD9JSM6kABdN9T7PunXzTJDyaamWZS76AjUT9DRIsD
api3HGbaqOBuOPpOoSeABJi8Ez43GynP4isTWuLvFGO/U4/3O3R2GQR5mWvqOmThf1esOQ6Erb7z
3W+TndxGzbFouZRhilWrtaWNh0Xg1PuWDi7Zg70PgIOlgxZAIFG7OnZZb+6nnONnnpznoKrfuBgl
sFQExMGT+/4oAgaEGFdqmJmaSYFQDAfwGy4ALZb95R65o36HnQcVBYaoLhg0Q5A4L6OfpoBj6FeJ
wBKzs+FTbytho0UCIHt5BC1dhgHYZfVF7u7Hrretnbjck1263DAaN9G2/tA2YGEc/sWDm2ZTvXiL
f6waGoIgD9qfiQlgS50YuiLFbqEp7DJt3zCM76p9uIlHXEuQIUTviHzFFJBaQCcUSUh+Z2+FeBsH
CtPknCsgQKIAEqOlKmoOYrCPWVhtuI104PHeHmegzu4EjrkArxBjJc5uH9uqjf2+SP8aUHS7AqYd
q4e4YUk7XQzhUcOCV9SE8pZ/q68iJRN16aldugoBR3E4qm6TsotO9EgQQWZeUpMHBd5c6fZfjyGq
VQoD7nPh5XCGhmohXnTjvTBAxGgST/nnk4AKFeAroTXbU7udIlDnmue51OHLmc2xVFcqndL7sSEN
GSWxgn30hHav9jsmkUVIuVLJH1lHUB4dX8evSchn9D4rPg4V/qS1ywcCVovIxgalue8T37yjfGfu
Zj08DsMatv0cutwgkpPYUy/XyUUhOykRgBAgUFx4YkGVHkhQnfLrOPWHdKmyTMucD+7cSLMIOY2j
WkA3W/nQNqzvDA5bLbr9MSYiP0+jt8KQ8/LX+mdrDYoqlMiYqs1PXOfCASsP3R2/hRIPC3sd6d81
gU+MoT41i/yLfPftbpFEuuCy9Xr5EQ4k17SE1Dd1f3VeqMU77qPJPX4teO9qZRL+MqPeUPvsQdF1
7DLNTtnS8Fp1EMVhqPvyeexynFOIAPpfxCJO0XVIzG+wNhcF0kdLpFTMZM8JeHgBDqMd74RK/o0F
xgg+kvI/2NNcE6vQQkx9tCCMo+KAHSXi0yPV8vcCs3Qs+avnDfK8QOHlkiQUS0JZrknQ1ZbuZqto
72MyVa0uVoaMs7Cstg3peKVkn/LjpwAta5x2o+d8jfE75dB6iS/JOjULNhB1hulBLFBUM2TZq6hg
jzKsvUwMIW5E1pe4JKCFdSEu6h2zm3t1FfUX9HVS9choXWLRIxvC0hP6tDPQVcEWEZcTgIuWzngj
7hQjmtqGx1FEED/l9FQXVGKXCu7UTwCT7fxbacGWtsADcaSJ3QQD6Rz4783oo9CkDOyaCGJIJVIs
31m8MRPJkZ26Ar2T/tvBmEYouoVXwyu9ETGPt8nF3A9ghEmpZIRMfMvLNr/37SxO1LnfvQbEkCQS
ONbeWKUs3pkZq92RvG6UpPH0BJDCLcSYcikuJKfmvnzcKu8g/FTrf+PTjvXcmFJJ3HqIqN+0Z5St
xUtLg+pLp28/4LXvdPbPpaySJZd5fCYf8aez2HjRAg0if8zC1si+ugzFL2AJiD0qKw4Hu7doXvhU
XzlO//vBe5iwVgUZ4SngiSzaVloUVKhR4dmvr3vzn4lxX6MqhlHoZ+8o1NBBG8ai4mQhijC5hoq+
ghkkcdtblBURvJmJCOtCGdvZB67oo6TQxr+mBPE0sMKEC+DJAYK4ouOEE7gsxAnh59YjZQMfZLZ0
4p80RfYcCOXUilE4pvLYvWA8BAh3wQd7zJHTp1mh7nqrABrGPt9QG6hkoaS5kpIzYRNXmvcrSiOA
830gbdr4w3DQAVacFYZB0DhWVQtOLYrLfSn2uui9SRVyI/xmQk/hNGTXI6l9O+g4a5OfFhNcJBJz
7V+B84Y7G/hga85UY2WqIVasBSRInXhA/2NcWglZ9S+XhAhKKI+gwbeAL5EnUODzltCAJpQDjcTA
MeLscX3PPFb7FfHLWEAKqbLW7v63H2Bi1vuM9ooU7gOkvpwA+o/d8eYp6+7/4r31z6ry73u+UPX7
+4rSSWflC9TTTbU/73044iDM7G0u2i04MJh/S6c4QU+bmQnP/fXNuwy676W1EaSnSOE2cMTdVKJ8
ztpZ5XOkPrxEu6IjxcxXAGzxOU5RTrVrPC+BiUeFZFEnm50gOU/L00I598JXSvyZoH6IZU7V4pgn
BUeeboWNcbTnrDsA1DSZFi4sxtCRvG91rhlIRs7JAOtc/jDHZEhOjgabhdYEFfNXYJGXaUigwVUN
BRLAXw1sC79+Y9CywEoU+9JRFboVfBY+bfIsoe+6Bupu9ANGDdMAvQmeDqnL0y7d4XhMUJ64sn2j
VccNorseBHrPtaELP0PzuWb5gUExi3iZD2/WTiUxI8z2jnbukRyg4tf2ewBcKPXXfErJFsoEZcwa
PFs3v25WqWzq1aUOGsdtMD/rKxgdQE0eFheykUzXNaE+GdL/MkW2JqZrbcIZB6he+kwojkvU2S6A
rIpTRJzkaGOs5+Z6Qt0kURIoAcks3NssUFectAo0/P/xwm7qrg/RK7VfsxIN/9MLZSDJOeBBkbo3
u3LAXkZoZHeWwdGl7v6OTvHyvWmtI8YGRrXLM/koRvm0kPqkSIwV904tYsHihwVLW7ES4Odpdzlj
sPplcYXj5I3emVc9vfHVonwM/u4LV9UuFVOJ0YyBsRYOe883sTdCR1lLuCoNVqsVsUinhtsTfUuf
XtzXoVMg3hEf/+M0XooZMJxf3e8hXNLnCK7wy56WU9POzbfZsCzHB86wV70mU6JPVOaJ6HArIp7v
sWSeOMpYTvvA5KVKKtH6pxIhEB9DySS9ooF7e2BZQbTtU+eFZ/uNXcOr5xeTxaaVfrzejX6ZXOBE
BpnB5bBzlFIIFOQ0XZEtU1DuobW/UtZ9QSbQdcJcqLzO1MfmXiK3t0/BZovfE7Lf2XKV9pRyg77d
6pjaIZa7S/0NkTHMGinBBLX0g2ZRUobVXNUuKWuzN/FC65Jq4m5yjuerl6a68D61qzPSVe5M5pYh
ds/aC+EBPrbzf2hXNs60x+dzACYLdWNySrcDUjeFATxucWTrztvDseb3TQ1zkaC7jWEDPoe87qW/
8AolZK8R/J5dhx6t4XKMiBnclsgdMfQ5ndJV5nVCdWYIqefC4N5RuXmsvJ2RIeiRR/60OR8Ds34+
05MLlNfz0CgVO2mg+HCCaJSurCt30+LpgCjjvM+l+Qws3maz1Vp6+zdSeAcBqTG+w9ZgZ8KqEPht
UxYOiRap11ZxD1o+oKdltBhONVi/hdiEQJnkG9GwEDxXZGZ/duSbLW14oYxZvkM25QJObxgUGhPA
vDYQS56Pm1/8DSPnOxXkL4CkP7Ok4wfoTEcmyoaUQlrUk8mtHmz1nSxvaRI81h9a8t2KohMh+aYn
+MbCkuMUyKzQhOWmKK57PNxw416KUCmwf00+l9bbCq3xEiOMbpDKmSIUx+jXZAtQER00EHXvIvzQ
8n8GvrwuXYA942zTkdsSLh+t0BPBvAy9FMFk6VKquoLppksyblzoYbYt1cLhE3i6eyUiBflfD1DF
KXXaSSsqs/UFheghDd8oROHIUtB04KMcnmY2Gg2BqE4NH01SMcjJiia/IzAPbA4oBntUL3XXjAOw
QpegSt8H8tSIXxCbneeGYWyNaoH5uQWV1dPHdTsdNWjQFMNEHjFDlwg0KZEpT/z2WOD3E3EtYNLI
jj52PKyapRcUPsIJ78qb4c7JnO0dmvEyA5mXJcz1vifUqIwNW00ZnQ6l886IOMHI1/EEHtEWrgEH
DCEFeIBYBgLkv6StIkB8HhpZVN84FQo0tfl7KkFK3KZgKpJVyxYmSB899T1tNk9uPHAA3ibJIAse
78bBntMqeGYChv7J+St0eBQnW3qjfHPzLiYSSEJ04+SVxf1xtH9r8v9Wbs+awFGPJ76iCcoCGwmt
wvCWy9mRKg+AYE11YddzLXqyo2D0GkVhGCpH7bGfp8fKVeu1P1kHq99DOopssCeCj+ttF8EEmTsD
w+w3s54BnT2scng7M+Y9FzmVV9tnx48wHDQE8IOgiFF88NNykU5gnTke0Sg2HzYDX5ckYwvDnvvu
RBPizPNVxQJFh1SpFgp5xVuw1GSJO29RSCoHQj+gUja1ORLw7e6ncFW3UolzuznBFmjksImqAMcZ
l7IHIQdnRiZ+4XORgAclN5Y0+X9aoV2GCaIEYk1sfuLcsToMTMfVMsOFsf4oDW/D3lazyX9Rt0yN
SzE9yRN9P7WHguM4SPLxTR1a2qDitiOVDPvzBAwIsx6Lk93cB6jAQ5hEyVZNUOHnVTnrswXUO7sO
CbX0nQeQlyFFWE2e8Puov5R+MAHITZsjeIjAIiz+imAft1cuk7k7Bqr1wXX23Af7CrYBWjaVuToh
WK7XIaRYh2LlibY821vdXFmk2EIeq9eXDHQvCt7wpcwhLMcY7rw+4uWRPT31fJk8eAD/4LvFG7/7
EqkIKfzfeb57AmcC6H1camRXDv+fCaObSYCYCaNZ1Z7NzyElaE2udgVWoxYVVSwzg4N+i0IQrJse
q/qm+T4Nm0Rv3J4R1W7UIbajlHVPqnkEL5+0nOHzF4Me+RAoHAC4YD6G8qtldd4PPvvjubgvJIX2
B7KGClV2Yi/WeaEvBpORP/Jts5aAfnaDhlyxGG83UQWRU6Xy8AsdIbHv+Fi6/BumpXsLK+spq33O
e0zJzT0HsYAjrGug6H4tXxZUpL8HsUB1hI0Wxoq4COSNZaecEyhNcZIdLVglsx4M73oAKF7SRY2g
GFrcq6t48n+veM1ijSMDSjptTRU2lY3LiQe9+fjk/pLT0Kj28YSeTpFoM5HWOs3fXO8jWc6gOEau
HFz0OCFUkEkDGyiLz/Oirne+2XGNakdpSO26XUC141JRVjGO42Hkj+nqG4MMMH/HDT4rJJVnQONg
AnV3lyGMD035PQWWvXpl+r7mtRx0lSouBgsCn3J1aXhXiZZO2OX6z9RAT8tM4H0OjYWf9NqP5+Lh
1edPmA+vtMO/nUDJwcAACemhsUjd9fWA3A6YqO2YU4mDH5wJBIM2ZUEDeDAYunyBR6W/QsKc3iJd
hYXmTFiuB7gDvrPeVXlXJokZGB4H79sw4Q/yGv7zj6ncxqkx3bP6Dm9mSaj981lYyUtHAPoC0+EC
fEhe/waBauQq92v0I2DH6uy2Gc5K92zJACt4DcTSdhIf6x+NB/lA24CUCxX5CyJGK3ESTbqIFv9k
KlFCfA8VQjQ/QbHbkbPugISf/8mSPOM9BK03fDng9RsvQv/avZjr3M1MA1iqdbZ2geEnWBc0Ip8a
Rs+e8mS+ntZMJ5hdz/fxI7VOW0DIxAGzclsQZ8kZKumTcFVNf23qpk+Eu0tjEEZHhAKo32VuWOZk
CUBvteM/fYzssxN46AZaqGxIoI6FX4GdM5N6WRzRXXR77SLH5CIFZx1r/foY5uyb2pcGffkW2uiw
fd8nz3nir6tBHX3sIgayPnqvWCoZSEbf6pFW+iY94QRVhIz2EQJnQF5gKRDDstZ5GSjtc18BZTKR
JOqNU8WVwBSYzK2qtlP9FFYw0U6ellxddJctfS/BOCwGoP9GCLoKIiUOcKOwE4Ew93olp+hhxlhb
Dz38A/RdAXKr9D5WRUu1J8Q5sXoSxt3gHgneZA2ydL+EjD76ZqbcUBVzI9M+lDYVT1l8p0r/hSOI
vas+JvVR++J3Cs2tXx0hNdKcqgn6DRjnUF4/OK4/ujmWsgoxp8esFGEU0TJhWOgUGleytAkRzHWI
UjW4vgPePjENk/UXZQg6VTNKTBSJlVdevFnBo/95sNbgXrEFBE5mfywxMhy7Z+YqsjGGg183Wu6q
OLxrlBxwocFo2PXRM/2PMN9gQcug68SPREhx7MBx+wQ5A/CjFiX3LbhB99YFAE0JW17vqK4G9smU
3kKdMxkIzAidGpBLXBOdR9DIQg4Y9e+oZZ83ETbN8Spko+tvuDv3UosAxsismfyu9sUpuOvSrt6I
3lJQkA1vf40zK4nm8WvGiCiCjuSEt9UnYRgH5+BNaty3I/Tw/NR2kwafO1z+rFJ/o8CFMH6TmeDM
0IR6XjPw8Zoj/63kPGS/21bW8GjbTsW8J/dI9HTzsasYYikWGlt5rE/imvnXSIqz/cM6g2n7RGbW
2vflj74VdHqJr/PC8UIi5hHsk3tYjGMMztr84IyYN+eXBZFNdyF3o0JTz/fGuiyE7icvsDAigVf9
psmbafUcFHEpIM0Cnu5q3AzaAMPI+GqqxeOY8NSdTdP3P5lfRfvZl3VnFQ3opvOPerKji+kL28T6
XZMCaaS1kD6UycH4GEx2fu4UDsN2oC3zXREP4qowAAtAdcX/VXScelYf2NFR/rvYIuAAErnmvbHe
ZekCl8PXMUkOeLqre7GuIc8slyMWYbp+65X3cYeuPvToezt42SzmYBE7KNWyEuumKuEqmvSCGO6D
WKve5RlJF4B4gONWCib1RkDz9Xb2ic0c8mqPsgKZyzYd4Iu/EGKDaDoei2QK++AbCnP34J5Thfn8
ESrwPObefvPz3nTNQ/35TfVSQ/OP7NPu+vY8WgUv71qxDDNtsUoax2dLXIH8zSa9jH71tNWtQYNx
xyhUnSB/DFSD80itRGCbtkG1zSPIBHWbj8I3UBOZxFs4jFsLslcrNUA9oAImEDKLxQz4sBlyaNDa
AG+Q0igHbjVVZfZrXjaO7rmoAr0x1tqScRM87/HHa10/5okEPNqRYt9b6FxxAgcXnDgfO3LEq6ur
cnLVDuSXgdJYLqYZ+NR167yCyz/zJl4BIc2xiLH05jD+ya9+zYtWftRcurjnCpamqL7sYoNOl1RI
+QZ4qSNiy14JHcuZq+tOpyBClQCKL7gJlIgYfQrmAe5zOyT6fRchsItwm04+ZC96HHARYVsPAaQW
t6lxHmobuE3VdCNo2XFwQPRokOVFBbSI7ZKZJRFM3PBXz96hHcudy0+p3hajpyvJbl9EJQJ4HwyW
5Tm5T1vJTtPnVEnWT1suVDxnZ4tRg4LdBaCiKYleICRqUu2cfU+b3nDGr++lr/ndwhf52Nhdcqfa
tc3dwM9sh/FWpj9WtxN7JOqSmJLPCVTYrjJfNw7BK+dcotPCBPZzIB7RCa04MSekKBJbr2FfkRpl
HVyCVPj56rwG1Wb5wEMKwHNvZrHTk/j15SmOVHEQDx26ClsOvQq2Ul92lH7a4GZ1MLchTeHnop6f
e2tvAWCBPcBfDKf/C4XYM/aa7wkXErdHTLS30Fg3qTamBb/xA9AnHmWQ54ByqsF5uFog5Svkz2Sd
9M/rTyaKs/uwicYAjlsT1+6MDCUcaYN4+NuK5CpoHcbtmVMEaScNf9C0oUwtE5ZaC0aM+9tN3obR
LdMrMxro8RHVKidjTyTLE2M14Pr+g5aBzSHZTarECgFL5GYTbK/XFXQBTUSt0CeoFcpvXs+3IrDV
K0aFK4oljxafTLT9taKGD6hN0sYNIIZJsmBICb5mx7Nccw3v1vbD41FB3adDe9zZPpKPZjveUS+W
aSEpspAqyg7joBM3VdWlb4hAlnGxv2GK6uTUR7WHbZiW6aG34MtaVUskR0mraKj4bjXrAbc7ba9h
FhgL9I5D1Pbd5tljAdnH1AbGdUxVtq2Kam+Y5f2J4WH7nzAiQFjD5iwmRYkTvXBMlIF07uJPt+I6
htuUT1UVAYaX0omgCSE7P9/iAgNo7p4DS4MtaP9+zHxfzvzfmfbC6xZ+hrMqhpwyqytnTOcVOdTj
P7KPcNLaAzqy52aGn41+dReJ7nU1UybHDBdkfoHmPHDtC9F/7ItMqqsvtJt6bPhpJwuZ1ZrSGb5N
8cMkjjmPZoCursvk+vrcuNiCX6jrpRJIJyb/xJeXT8XUSsSFDCb2WFdyDGyS1SQZh7itJjTVpswN
+eVKgbTf5M3uYa+z98XRCB8aw4CRA9tCXF05wsMa7LfP4uW71Ik5IT90RSeHVH01xV7z5X7mhXkO
ti/AYmQqfQbER1RIqgNTvQXTR06g9QXYJoJk1siJU3zDYMzZT4ObtAXuqrqLpgtfq9Pe5DkDNhCI
HzuEZaYF6lbHXgcuDdZvIfXFTXFP/vnIuV87orRqVAAX2mEDc/kpBJY0paEna2FbX9DxA4hIN6Hr
boNc/PhDo4rWevDuCdUinRUMIhxx6sAJRVbGt5GcVuJ/+bmSLBZ7NHY47jfk6dftlT8yBemhXwsu
QApum1gvQe3C+JcHQvxg1r67JRy9mlpcVfl8XvFE2r2eX8p6tF3seJPHUwi8i4rDrGUPh6JrpE8a
FTKO0dSpH0ljkV2veea6HgR7XNohqG0QGlUUG6JBLwrWLVhm+e6raE7xekjhjU5yHYxXMgyrg9WE
WlZcywUAYs0iXIk09nMvZiaKpjeuz8iTaQVVUR8GxLx3CUh4kZ/Eo1q2OIIVqEJxkMtIs2AEc2Q6
OsrxJ+mu8Y6kjCR1kPda/07YWnKjvAIFPBkwHoFuoyrhKaNx7knsV2kgqjRIF++q/9Zmv1vPkaDE
3zt5/8On2sGQMpkZ48wrLalHUMoswfFjLbCZhsaiOqbt72bkrJh8HC4osj2YLnEyENf9zvUM8Asy
aoV+ExfJCHXAtcYXMMnjOKhRow9uRdrmLizsL4qjoKUOxo5u0jYXS6v7vLVj0C6OKvro5Kk81fRW
Njn4nFu7NMTJR2Fb7nMi15XKXAEpZqJcFd8sQum9O1bzTZ1URS0UcV3TGuuTf233viVaMiyiZXMW
uDntWtAor5EQUZibmZpvBObOZpa3cgWzI+rO8In/VRXaJOhov7ZoAAzYj0GgcUTBke0r059zXhoW
xB9lVGhqDvh0rYWIFiOS+YNnnzlvJk8bg0e1+ve5ZSHgAmvwSmCqiu4AUh1m4kvFERkvOB8GwI7N
+fH4xA72brqtkgcFi/wmvdaIE0eQfwebXoqF+jiAv5gb34YUTEBqbbVWGPGGPGFfwa/2msuhxA4t
8tu/j6eR/s3tCEckyg7aRLowvXkmXprUmN1S8pk/65ktGvsEW7RGXcZzkhfjCxmIHs9pwmacukSQ
Y//nNQgKaxjVSQJ89eze8r25+vTWdiP90Mh3bG7LEGpDoKk7GmOUQPSRTaOm8jS4HNVMH8on4n8b
XgPmUzhexlUNVdQ4eTgUiBwBveJQFLIO/aCDCeyh4dllVHumrN1K7V9c4flACtVRcx8YpcNvh0QC
T406qgtrMblqtCse3hPSrkvBLJyAbvZJpoBAYdm+ngs1GDjSBaUVBxjodud27BBVx/l3vK9xthPb
9P4/D1UL+sWStBaHaKUqdXKRn0niJdtnmkSuVqwTDJfrNG2+lBIpvIFM9DFf1DIHIabSbhvmWEPe
1BYqv+mREAxXzJqF/EXdM2jV5aBco6MiRZR6tA6z5qWkhNDthkvUtN0LLkZgruKjCWEszJa5KKNT
qsLpc91/k/YPRP7WbFWEWkZEDy9qp7ZyXVQ4LuU5xuHdCGPTpXA7xeu9PIFp9pdQNl63FqyPL6ie
TB1hKdkQk2i6/17AnNHfVdu0uNYvetDA4Q++iYDtgVQEFbEM1zWFy5cwkH71rGjUAiJzl9EdsjPY
RXlSI3WsdUd60EaNo1lvJKYEfhrLmcfDqSOuHbjuHMoSzTpD6JQwElZKPGLf5qivomvHrv4eM9c+
daWKrq4fo2S2MavuzIKQUI7th/OaW3FcJxlRoyJjOuU6JKN5dXX2P56vpM7NXunRpGETcflCSbKE
4VhyW02XMRdaRXBiJzqtuHz6jGHgtZmciMb73eAi91hki6ohYwyYsyhztU8AB/ug8eaWNZumtzGy
pXKNi02Vybj0E0wblBymfQ6qBnalGc+AyQ/O5aIw0JKAkkbfUL5/hieEayggcg9zg6/AjonYMODl
6JuYD6NNhk6VZbHAnzwj6GPPl+k7G+h4j4JOghG+fk78C8eQiO/HMVw5EHjxzRyJAb3oEk32SrXQ
aESdqvQ0yT1rEJPONx8L8rEH3TSz7wFdOfZ6aiQM0DljN3nYbHHvTykjFXFapeDPxwZjK9fNUbUE
TMoiCcJ3R5LnD/uS0LH6u1ZKq85CM3oPpmWSV7QHK/YcvuvAszp9fHQMdWD/+ryI3cD+dCPnIEgm
TQhHBPhs1sngnCeA8lS58rS2TbkDqLugLDrs2KJZUIGAHTj4QDW37tfFDM5GVgc4uXFGWgVzb/Lp
+/IAe/DI7OinSQd/aa/U+pXNQmhMVsICpsY92ECY/Wm30v0AThq8TXTYnwvMaDsddw9EK+wHUjVU
SjLHP8ZVCXntAtqCHk8VtBKMer3+UBeiC1dZ0jcZvhfNC8FYVS/8YU1E5qccakv/yhNSU3nVIj20
m7+yEgATwCtptCSMIdSX1caOdvh5woRpJQIQLDtSltxh6K+nr+yvflqtNrng8TAVk9rhM3VKF57C
8E0g7mOMGQdyHoe0r6MelUNcwl/AVxrn8sEe4hjqTsljetNWRlDl/4FJLZ+bcdFejct0WtLzrOKg
C5FhrvPJTTBc4yeGGs9bJNPD1hLOeaktiOeBtCeoPpupPubD6Sm22/NOF7jkylHedS1HkQXfkCZT
x4EwadZco2guWfOcKcPvS5nH1IQLBQe15g1Fs5KZYBlmspCzmZZ4QMNaOAdNUGOP8XDz4wZwmRCp
csrL9az/6gxhEVtWbph776iNPQ/9GEWYVydG7mW+Ki2ZSKuEIXzPsWaqQtmYYqVwku0FT+aV9nM0
Y9FoKVXjqc2iiO444gjdENH9BWSKfloapso+sBpojOet8xybv+hzXooyoe7Y9Snb+lKJ2Jn4B8SR
Jkh64Hl+Mf3L2RMW0L5hngGMNkvkno6+P+OEmvIG5exawmIJz3iOBwyTgipkekyRPeHUOwhaJzCO
CBehpwJubcyaZn0FJ23ya1XtPPvL94ONCrSKwSl3kJNFN7aGnAAUfWg9ktUZMqw8dXuE/J5scMPJ
jAGtpMbkweeHEI51/8WstOr+CHgqn5Jm/AKbbNABdS68GN8eWAcpn6N9J98PBg+0/pfQ1Sc7ZMmB
AETbMOnlGqccdkvXwlUkvdWbcPvV9PWQx3ONn7TIA7njPVJLXLEtkZJF+U5gXiDUNSVDQOXgQ6G6
sQMamY70ekOy/laKQnj1WyYUWfNyvcG8Z2rVYUADjA+C59PvFUSqQpy99dw12Er2Blot5fqJwlLl
Sn7F6a4Qt8PFjgrR44U7xEImh/ZIgDcXDhTHH/L/Rq3/cmwjocwU6nviYXDpbNnz+T08KGewYhPx
7Do+u5J0Fs0yMbHEW30DRAIEat6YbqQfcACl4gd+et4jO6+pj/5tJCEmWocTE86gB0JOr7CLN4J/
IQaJNdlLKRs3LMBAMhLuAPdRuxGltEVw8DlEcoEBJvCjTo4cSsmn9/IcXVhovyElLIkmEAf5ht3k
/XbTUBj925Dm+TIYczdsMGJxpm06NSWIXDOW7Iibe1rRlbw2z1Wy5HfM2Ksm7576blgDxStGPG2E
hDwEwI7giDdcR673iHC5eTIuslUeMrBJuwa+xj2rQDk+yYy73MGSyA4z692kCiiMqhNFLwahUfwQ
Uq7A3mv0CCS9YmzVrxKc9fk9Nt13uyz3XrtBWG2SGQMMZMu5em0J8ZEdGxZ2+eLVD2Ht5cpcQpBC
CYspidfDizsdmfftSJCc2XdQtH9ssHxeIqL3j3EpkrhXmcAXA2rcdaRLZcsfLKIKGBbsLgZ/678P
Au/c3Par0t6NCBj8H7LUDcE11ovFruquWq6gYuB+fefMKglQ8qjusIHnMjimxdvz7DLQo7YRBLd8
+8L+cXYc9dIv9fGtq5yI9ccCsDsDYU35iWwgRD7/5F1510bEYbVXcrf/jG2mwsQXXQuBZgZNX6rJ
0G/VSPei7AxY5Xw7Rz+mWtrLPnFqjo+9HmRsUGIljeNVpdElq/KoMSnZFgjNW5zZGLqd2B8X4CsN
heHZhAkcy0LLIKybZMVGzg+FbY4S1WnCCzmULy84FJDh5jNPWmKNxpfuEJdi8E850RL52Mdw22km
s/o9iVel+hBzWe+qqpeKAMRGiphRGPZ/jBBoxYSNhD5vuGU7WfNKQ0gzdXJdACr7TTfhLv4n2RbP
8cp31ya0Ab2c5H4QpRFm/k0pZBYMwEgawJFMKzFwY7IoOBuXTbY8glTqEe9je0B74sLytxD86b/X
3yNLkp0NkyMVnVKyzEOoMPxxiwI3OUvhFuF2yEUYLHM5L6QVoQN+pL0h5y0xRFkvsFo0W4e5lTm/
LDnKitzyS8P+xqNcTnJFSoIibeOyh0eKCboKVwGmeWjwpse8mT0+5Qlw9fN/dNbFMGNgNMa99V09
Kp20R1MZrePo963cUvTY3LXYOZBbwQY5bK+rWpBdw/6KUjcifM8U6yW9l8qbEnbPorerXNs7JCZk
gqCE6VKqIhVPzyC7fQWY2lczk9yLg1RCESb79bgMFFQyvs3lLtKgdgK7zApvdVMwHcbzNMg5Mtib
yuJK2uf8N4UUjOVCu5crogvLwnI5z8pDvkVDrepkB6AbUh0moUWQ0wlNsD7u9cfuII7gtAUDSIGb
c5986CSAtgoqW/DXaI1uINkjgkBgvDHEiNUwxXXt54ujldsM+emh/Rndhxis/KaGm8Zcf9nKo/Q0
AfC3wMxcqhEBwEt0o9a/zLUie8Iu73kFJhHEK1TgHJnN7gVOORGT7TlbLy1BSGA4JxszNaAzqFDY
8+lrNKlPd88KTezT0ao4qpxi3htXw03AwNAiN9iLtclgz8RO1np23vfkI7x6XQkHOiPDwBwwFsFv
IzP6xfxzS1bwnfF1DEiHCiP5sAXBpkzMTWGKRXB9QqnRWQ2YkB2HcXbXU2QxfdYHvKvxZ7cClWYi
4VxwtiX6wI677I8CavjoWwK8ERPy42id8e/1qpvnDxL7mRGeqQ7JozOci+6LqBLWwjCwS1SMVj/u
YFY/VlSo/LGtvzFirWX7J0BgvptaH2eoFR0CjNGbg3+5V6EEDmM4RcnZkDrS5F8o2QPvJRvcr+NH
oXZDmpeXUf3gN1JSj7Ns+xRgzU5CRVrXlopd8yu0NgryfICf0nZKr1IHPELTBET5IT4DNKnqjakr
FIx3vuNpeaXQHoHktS2ZHyKLtlsoCNJo/hIOHvQT8EsWR7Wd6dw45II+k/2qUZoScpX/uQD8HVw0
YiAJX1YALZWVnbU7WU8JY2/ta6gsGpR97KlZc8FOVuZhuN3yuTBvM/LYa43sbGVxLrzwH/P2raSO
eObvTp7MJT7e3mpTjrEkDpITT2cXLcjCuTRC611/KJ8orPqnqOT0g95XSH/SBp4qmOKBQbr4sbkD
IzF4YzorNo3gE4f09W+vNMclbQGYbRmh07+dbJr8AXkKOXArpCqFAufFZcY0nZ/fWieejsWXGZr2
6XzrZzmqHCxNfdLM9hJpcaO0uAgcz9RrJIR4folgM4VQRGjiy+8y98IBcVU7JG0ANhJ2vuLZoPU9
TrNCK7K7+o9eOjO2rdKT7oXTM/+ZeNGi+4iWPl1uSXW2jlCIycoNnVC2QkDZrS2eO4iZpDPCCJiV
/M3ILl9NovVvv7DM1b1pRkXzaWJHKdVao0720CdG7ZzZmwHH2ZaSNPY6oP5nX+un0F7eeMfKiPdh
lBpGkqGuSMCz0trV7uy9D/7TvEqydMb8PtX29s4epnRIcs3o1UJjQal1ypEnONmfXuu50R/brSQv
f9IKS75TUauyXMLk+vTaTM3i6vcJ/v2abJu1ulGKu5Nqz8so0vbqVl+ytb8LDVkxgNA3i/m2nAsf
gYYD0aoRTz+OZzxNYKJIVPC/PGKgkIJPZbQl9HS8ml0Bdx9SFFG/d+X1ctxGFJMaFQIUlzls0ZN0
TEUo00AeYgFnSuvJ83DVdHQBs4+lc6BaRDKoKl38ttWkefAnXadZrL3x/iWzyAyIFabqJBv0yVCK
8VbrRRzoNdvkGwCWZ/jnYSWv4SALbWV6lrGty5cjWyntMYFHUrhd3L/YiKwajr/RuIwK+zdFaDwN
vw5wTDgf5jpbXSCh2X8idgponYovxNLi1aYRpwu3siBmAb8I4o/6JH1rdN7yGrS9R63WJ+gndvV8
+B2GUUuh4LdXaoHQM9Z5cDUXCBE0htQILgajmC6LJLkWEvZR6c3F6BQPmC+CP9lttZObKBvsj7V7
k1ofEag/0gx8wR+t+s2IsZStwKdiUzz9Cx4OH8mfIodprmqgiQPMZDs2gIbwErcw0Oa1J6r/om5j
hk/YTwo6TLGpKPfvwaeH
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�*��A]�~��	�y�g��s�{�y���6e�<b��;�%���f/�r�X= ����'?��T��92��9��;E����T_�V�t~���f�g�ۦܹ�6j�����O�fꉞ�LaUϼ�!���{G}2�I�3���u[��F|1���Y�'u����~��L��D���25H�Ђ	/wi�'��Ғu,+��w�z�zF��PW���×��R�xͤ��"��Q��{����ʺWB��3t�#_�YT��ܛ�Z�q��KV���m��2�PT+ұ0=t��+\�U��ϱ�F�G!��=T�e�w��3�̝9�=
VX�_j4F<>���Ư���4�V����4�������%�C���}��Œ��pSSVi5f�E��Mu�A)'��`,u�Ӎ�u�d+f��i��
a*�0�����D��j�'� ��Ja�:��ᡝY�i)�蕁+�`z�n�~���$@���Ʃ	�E�K�K^�x�TPe^H��&C����Uq�h�h��O:s��M��.��,�>��Z��r���n!ֽ���#��@���������I߆K�6��D�zf�K�1me1?��S0\��Ȯ9k���~�`xS�k�>��[<��z�y�J<�dv�3�z��=)���A��kfHx?�Qzup%�%��/���`��b1��ƕ�@��k&�2�/��8�~�7�!9��p�-��\��Hg��T����N�w/H��X8/�:�-������8�[��u���v�-$ׯ�)�WB�������G1�Q7���f0.h����Z��9N��^�v��r^u�7��w�p�#��p�KNK=AN��k�m�L��k)mx�g��?�bG-���������(W4��xM�UCg�FHS����#��]��*�9%�B!���7�~�V&�-""��<1�Gh�厇�Awӧ]!��iI���ë�">��!A�32
��[���?�mJE�{����b�ҽ�Y��C��K6�^M���4sQ��"��E	�6ؾ˥L�z�1��S��Y�!V6�Z%�R�x��j�~�SCك��X��<��b~�=]b���
1�� ��/�
�>��w..����ʹ\d	J�� �e?�ho8��_�C)�����v�h��@
c�ઽ����]�߰q��=9���\-![����K�\��ePMV�4���-����+��e1���hy��S�l����͂�ԥж!͹(����.ߠ��Fc�,�\�m{�0w�9����3O)��d2C{\�ւ�M�����(�ƻg|Y�K|<C7�L�ص ��A�7�$A�&��;���KT��g��5�����q���m��q�
��dh2ܠ����R�T�\�vY�RΦ�ʡV�>��25u̙��ï��ޏ  6�q��<<�#<�)%���Ҧ�^X�9��X�2|���#��H;<�-�&J��X��<*��|�� �:�w��"����f٩�I��,!��[�̿p֓��^TON��"����`<������N���+!��!�m$%ga���1W-H�ˍ�?Jfwڢ��G��%�(Lj#(�� 'f��S��u�h��哋��tA��Q8 {��(@�c�<�>>��/c�{�bV�!��az]�Vݨ�V&P���I�� ���M3��o�u_����Cv�v�����0��u{U�3�b��-<�L�S��K43��L?�C�W)h��z����@�I4�`���Q�j���~`�
`�4;2h�N���߻�:����a��r�����P��
7��C�%��gc'$!r"!{�nOa�;z���vU��6*!�s��Xg}(zX ���v��C��[��2��L�ш�˃��5<zW�[pb���i^�)'L�$8�b�������@֝�Q�$���g4�O�V��*��4�ݟ[}�8pBW3M�v��F8Pϰ/�C�$��7��V�`CX����8�t[7����NVn��9�ڀ�q��޸k�����j�+��6	�"-���|���.�T{�_������Zh~����<`�3 @	�G0҆5��t��A.W{��/�7U)�'��S��]�l�c�)�n�P�n�x����"�nΓ���'Tɜb�[��C���{�xe{71t�D8�B{�>ݭ�a�J4L*v���%`j�V���X��z�Ã۞mL�F�.�a��	q��ހ�țNI���3�3���?��7���s�s�	b4I|D��w�t��Q�jx	�pG��,%[�C��^��C�������(J�D�jIe�p�
I�H9W�xW����v��I��h ���*Hϻa�*�YB�g�X�v}��	L�=kĘ6�Ŵ|��YE�H���6�~U6ߓ�~Cb2c�&��aͨ�l��AuY$��zY����5#�y�����<�����1�+�x��9�)��`�<ׇ������r�ZT����}v�Z��gŊ�3g&-��򋣹<�$���a5G�����B�!F�UO��g�̚��?������3��]�g��P0���%��'����=d��#/�
�h�I�)|���V�-�N~E���6"*W9�lv��!BH'�B������ck�Χ���^������� ]���9�ս��g�����ס�  � 5iP�a)ב�,%(V�ꁐ[3��n�����EM.�2��T_�>�A7F��0+��4O�	��RM��H+ʚ�)t.E��Θ���y+���y�5Xe�4ҙ�b�ӽ�wl'�J*���i�o�~�d%�����Aa�۾�ú��jm�q\�ğ����֨)�}�!ω>W���
�I�4��]�� c4iMi��o��:��ef���h6��n�dB Ԥ���F���."��R+I <M%��p OC/�h `��ȷ�*�|2B]#e�]ܔp����_ڬuZey^`R�=�8�,�pՍ*� �\-]�Q����a�uXz��2�2`��g��7��,����?0���b`��y��������s�&<.�{���i:�������*��E��96�ouE�.2+zc	�~lH��2�Є�q��9N��}/oE��JJ����b�b�V�ǬA�J���p-n���P�<&���e�]U����
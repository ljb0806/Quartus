-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
keHULkZNBc0taF8cENDDqqUP/H+NKZqmauuwnJT4T7oKeBvy1iaPqlU3Nyid21qFPvRqvcy3l956
Wp1cV+/ynVTRAAFRTyBQpKzFJlthTaOo6DLMVR75Sv9pIJKi59i3Gl6LzSoMKe6InMw20Mlf5kqN
qw++Sz2sFS5wieksIt+7htnwFm4ZFubYthTeAk0l+q5XZNu19Jbqu0Cqf/tsFwJVMhmSWcoLlNw8
mnD5m0zds+SyoGBbQrtgrguPGgxujrcBkZDM1mxP0rpNKoG0P3PN7B4SoiHdx1ecQ+jp5bFpnmnC
5X1ooIQ4ImYO42sWHAUO0cxfhvQkdaRAEebXyw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91552)
`protect data_block
bZh3k7CpRvRYmcL+zcZEjbhSm7g+zjjM3cHow19kSEtjsRctRlIbb5j2JBpRo1ttKI7tte1HVAP9
hob+bT8re0JoSZhi/RY6BdlXu38SEOv20YaS9LMxffa8tEWaQVCd4UCrfoNCr57Pv4kBd7SHfeSF
Revv/cD4ec1VH92HRkkMjbLtl0v0AHjXudS79zr1BnBiv0kbNO4QlCqwDwYCDlEqsS5gyfVnB3ZM
ZtHa59RdzfwTSKLnbd3+Q7duAr7CfKqU0spYjbAejc+KI497j4iML+8sh2hS0YyZA4mX8l64iWqA
lABn7RbfjNfNLZ1w/d2DQfNKP6Cp/deyNNi/vD9e82hwtOBU/A5e+X3ed5xghQ15yR+PxbBnJqDT
Oy4zuQnyG30ISIcue4fXXqlpMPSxkP8vAV1dmZEcgGJYe3XPIaT7ECFIt6VGpO0JdtIT+QGxQYcV
qCUSzsMCrhzquchW8dSVWfSYIqA67ZTJHE4KGfcFSoRyiS6K2F91ypeCUjsvqxomSarqKEC0yYuM
Ba6xoIZU+X5NaBfwa6AydjyAVqDzRjLf1sLe00ul3YQv7O7sLtjSMjt5/yKxk+DWtH8mpMYq4xl/
1ARaE6lozMSy6322uDNN3xPeQgk+8pVJKMMNjL5j1vq6yO9UkWYsvjFRiGu5ZB5sEeU6Z4sBwOM8
/P1mO0K7ky9Vtj45hozE1b6rtz1s59CPUrRMjaTEBkE0jZBw8TEe21ib2mAq7bTVyCSgvu2AsmCE
sJmwNbKEFfpEI96PI4qmH2s0yvEQvcZ67d9Bw6eZrdrd60oZf1+GRlPxRMtFwA6xlVnE8j+gjibu
ygUCRHlcQTwQQ//WdDJdnE/gumGryHNkNbCGvUZ+VhrvELyYZz3V1I7KyhrGe3AgyrNghrN/01oF
w/Pd3g3sdlZIFQaAVaujz+7wuB+oGHXB4tLI09AdsXYyypJoJILe0TWODWHHyjToVT0DHRONlNem
ex5N/0edv9vso84XOCTaZxZ8RLTQDOOR501qOajSMUQLGKJXYeizPF/cTb9T5LpWUpEcP7Ry7ej2
GWa+lCr2TACdDlL+htCxde7o8ymow437zDJXqbF0J8ZEvrUdBAdHTZr+kDCZAa752WnjTMv6bkue
QxermV5nQoIM7U6HwRKhnXsTau8B+JhJw01VsJ85Kqkw5uL5tmPJZYXwyBbcNI3j2xtcho90tBJ8
BTQ2Ucsf1qwrWN+M8zQ3WoidgJUuM/2D51/Puf8uZ8Dts61YsnoFJRVLMnugnkqjL732GxZqH7Ux
vx5oniatnHydL79uNgcItsa/jvE0hbBg3GfEf93B/L2d8WKG41k3qw4Iwx7dyvHtHkoHThJm/swK
iQ/iG8aJ8caxpqwG9JW7GvI10CgCaO4C+Nf3I/tfc8Pjn0BhojCOXlfFNNaQo6/WDhHe3TkxHs9f
BpDqc40LGFQTfrG1hyokueHQWzBa64A1cZ+wsAmdUzAV/2TQElaCgr0bpi2qurCjOpvwOy+eehRq
F4K4pzmpUMIrY6L8qbjzSLDTi5JYi9ec12Hxa171WRH6mHkb6ZrvjrDEn44SfSYenBMSixEcfHG6
dXiBl1vMLeVRDQAudcMPUjkYk6xk4Fyu14vOIPioHfVERKyZpkzuHi0kVgTkWINX0yvZY+Zx4Xdl
M9EJ5PkzJONYa27gjMWcxeP1bdNURTxzPYaY7bHUnIEfhucJ8JMnXxgQzOScyNvrQRWUf+AL370x
nrBz1dAZdiW0fUIYJyP/JL/YdC5NEgXqFuXfdgikE76/xiwFLZp3ZJc33pt0DSbVGJAsk3mWWKv5
GBIz0xZIgQtx/3QpjRHkcb5nDFCloP00sZLIDrTSjeuIBEcqYSsbzOwJDMd83YuHpn+ZhyMcGmG6
H5xqiYnE9hessDXo8POElxdXNnlpPFVB90F1q+ODDUEqmMDM2WHn9QWu/QAxUyqliK93ynJoUxQa
TdqLAbgkougEGIsMYZalKJxpbHMeVyDwqfgyeh8UDZ6R9zycweDR7IA7TTcVuvloGdh34FMl6FCj
GYtNKY/2tnD8OAM9vY3hPNbBDpzrZKv+9tLvZTIx6aHc8YNxTf+I4TjQoL15Z4tZWBanvmcHZqtz
QDMKx4xW3RFWDPvzi2rx3z86zWqhJGiDyYmQPVMSrFrP49HiUKC7vCH4neeKR7meA4DDpygLTVPP
CcNcDnrfClF8oHqPR/nLaGXPwt0UUt702wHWji/zpyzdaBNh6f3+3UfnyIbtpviHd+LQ7D0QrscX
5yWVBjlN9FynB0Pf7kB/e994j0NgTUpMY1Gr7Pi4O20ZYpgQqti16TK266Qt0nnUpsvAQJFaApJ7
T338EuAIPtVT3vqEZJ7Q91WavdhvJ1n0V1+4A5zW8+kL0NmZV7ZEaUkELriuc2eUVOBc+RYwLZoQ
nYuYp3SdZ1Z8B63lt8osrUKT/6+RUOXwdFWuDCbWdunsmjTTvOuOz9+zZUuZWyl3p6c0lqpUv2XL
eQiJQ/utmF0oMRKfu5zMFkEzAFk9btGup8M73PItj7VP899BPEnddER65H9uYY0ptVWezonnZED/
/k7HjElra81GvFeRUNgq61/Eq1fEUxfXcIfSbztnTRPF0kU3D0Ks96h+XTKILB7Jr88fsB/ou5ZR
DoyzTlIn+j/t3PYym6pPjP62l8g25Tncc02WYKE55tW1wJHFb9R5fETWiBcVVYMZBtyx7zw9MmcX
ko1BnDL3+LFufUwSB96CTvP8ltvVKu3NjAx7R48sUrYWmItlbX+tbgeRu45nHwIL7UNXVTrt1KLP
hXmrV9rH2UA/w/kncv5MCBjUKW9xt3GrolB4M5+oJNIsOYh7iMgNgenBUAZS8ORHNOyyueHZ+WLk
XMW6RTjFVykFvfVN0aqUSkJxZBdLSNJmGjO84MBgdxV1MMZonzFPlrgPLSV9Mn4rWJmEbLIcswHV
cOsSuc0NVte9Ue3Ojz2ou+ZUaJSjYkaivTEeVCiMGalubPdWY/3Z1prd4FKu3RZO5xsn6EzCJhms
sInVRSUyBHTNhmvkyn3Pej7WrCBjolUTqwUD95Tr9cgKEAU8DUxGaLTeVOwahZajwekEsWAO+Q1E
TsEhJcGw/sXf1n5Un7VfinPgLi8bF6Xez96bOyycVS+0Ol8TLL8UgK3CBe9+00WybQ4/QDGr/IvX
fYWDf2de3T48pZ1MCxNv/5Nya+HiVgVD7FBEfXhDWzOOz8wzneA4IobxquySK5I1vYcZHzYNcXhe
w5gXswfJ/ruUuzy3NLzyX/idCd4HdePQfmmCe3CmU2zhyIIzUfBZdWzpwcfWRayCnExRRAqjuqoG
6tuHEJLj0BAe3JhzMnn59LMLXR/a2rkzxfSkvOoEwqznKzn2McFsWFXc5YCDTTPP/b5nq62jy5yd
2GH+x3LnR1DkmxM1gDwvdNnoi9ahYh/8fCU3OyLGoz1jH8oUq4yvJPVI20iCv97VBQo2fABAAGH5
lirX7wfRX2rNRR4aGp+i0cZ+090xf6azh9NpideCtMIL0ibYfooI+WaR5m5bwfOblRwwDucIHoQj
f5Bnxez8i3JUZjRLCYA+m3IkSo+Z0NKBnhXP3zF4d0Xlci+E0JWrS4fsRd/DnO3tpRf3sdTu0LvY
4QFJTPDAAc4L3mFfJGjbKW51pImjkwxYs2UkFZsg3jQ6WMFhw4S3NYdYdo/4AUCSVm06sjSxRbaI
Scy3z/X3LA8bfio+ZZK9GwTRe06yutL9ZLf8F7yVnUUhkD5sm/6qXx6cCAvVAJ192ARKyXGg9mUh
2+hvbuJLWWBj3Sqqr2tiKSinKgR0nA3K2Fv5pMM2knLaRZ+S78eumkdYHnN1qW0YRtbUvTlsJSUI
4EiQXvwOT27hkiGtof5aWDv8Sy2qaroMi6QytHBDsEvs5dJMb8sgi7zNChwdpCSnCH958g9u9WFF
7tQnWgn9bUCFJg1IjObWBGc1VM5xHrYp52K0Suk0WWAgXqlPB0Ly/RGfNvfVP072In9jfFRFDqqK
EXFjyjZ7qvE0lGML9ySSrYlr+WBl3tjw8uFro8luQ5zLVUesSwU8YTGIXpFwLHRMwzabLQEoF3vl
utAJcgsIYtlyu+LlG8SdKH2uF3pAYvi8CxcLkGYBlVh5DGK9n+WfXorR/B5iK3Gpl9SDt935kkGb
kd/7rvicCdAX1Otm0NawNoNRYEOz88kBZdlRyzZSl04P1sgoaCiMIFwp9jMnoicIavVB6pZ+LD1z
1FMKMuvTty0F3DqFEB27P11byn5R2yxn08gveDoHD498sZ6JnODw3aZ2TBV0GNWd5rLc+qF76A/y
+Q4WYDYAEW+e0G9BQjzS5pTnBjd8TFF9eyEWjNnHEIHFkjZf3rUcS/xfvC6MbcHXJPdqo4QVZre9
SH5vKdDCXRMfu6t3qjY7ZMjgyv6xIaO0xYdrCgxQ+XrEAJCRNkKP6gzHFpCH/KJnp+7sKJetJadZ
M75V5lR2BF+iU7jLiQp7PXhqMjCzvPhUpzjo9Ivz9+D5dxwzWdHmi6eyKo9Pxiy6TJ1Pti5ezwp6
uvDCgKKJyzT8D8Ji5yQgxcERhuC46BiiWQizg83Am1JNhUvBVJevZ7aZfH8SvVfTcxrrC4NL95va
ecebFUKcnXz0PRhCRa+LhrMWvI6nt3FJH60ftzGIKiU2B4DOF5HE9B8GbNRVJ7OjtmD9JonOKnq6
Aekf3vx9zLz5TwjmshLMdT5mPO9kaEjZqIYpNmH1z3w+8dSvn2yxIb15P1+LMzkjr8a6osKzpPNx
5kh7TEAOb+xOBnj2x4kaRZ1FEHStkueICkBRsnrDNDEb9BQdFPHAsTqpoNQ28YEVXvG0y8feko6e
Y0KEExkEAVQCdwSijjjw/0qHm/FNM/5yzkN9kDxL8hg/DL7ue/Gh2wN53fJ8XdzKeMnMCCTWvJBa
eyXWfpIS5aPsWWN15YRDOelHVhlKm82YWPnng6IVJkPGWKjubP2RTpu4lMk4jd6uCqOSPWCvqa1S
K62i4vRu0jMn2nLj1p58OsY1bM55W6M9gHXjfoFQQTlEf6Vvwqv07nC7e396ItV/ELowun24lDHy
36V5TK9qIE/ftUn8gMf13BX7U4JDmoKYvss7sLqpDRZ+afcE9qhffgF+JzOtYrTDtCwa7ixjab8X
HoHeOblIKIPK8kOpaliN+Rvet7hLXgPEK42GfRBEoU5bb89yy6aYc3CFtW11a6tscEuK892Af15E
jJYfOUCbGEZC5f2XfkIUiyZCdpu34bP1hqPEOm1fJxdYwfpH/2bTGHTNFwT5TidEPSl6x9xpXGHx
5kuMn+z4Q7N/AtlF0lE5zzPIsaKs0BVHAAi6pAkzO+BunetyUspEj4znaKmdFLApzuxWDopQjipr
F0NMeyt6n8L8aGkVC/+t3D6HjyW9++Z8Rexyf+S7AQkKqnASNv/8RBwpht+xU3mOaYHxzfmahLoV
Np1hK09yvWY98rG9/xQGLjWYRTXgQLXOgbWenjRJbvoxzSD4yi8IIHfOJHmZy+afv5YBPGQp5+au
CgPyXY8qM0f2m4QBgROsp8409K7uDL0KFFpni2VI+wxl9BL8BviX8V2GXAUdnsnQZwsquErCQZAI
U6K5/XCaPG5NAnmg/It5Ze+S/614HtaAB6VGPOHelIU6M/K52h86tvTtJJIPRl92F0WhK1IWn0+s
/xwzqMybg0AEuf8/OKVBFd3em3yNmhPD25dWlbobmcC70wyh2cLtQE0UCfziABlmuyVDK+CE2CHI
kUNvXlWnqqFm80+4qSWM1xTKX3ppctTOmM6Uc+cGsQ+wEtRUhV/RUN5BhERbHyN3P69avIKfxIyy
SGx9bOEZjrHFlRg+btX5xBlNG1JgXtDpyEpoH4l/xnUhHmb15+kvEmkYwmRg2qBAre33RT0RIZ0A
BLsZ2xf3gXgiXOLFMK7jGlWF09M2dVM4ofdQa1SlcwFFd3rOzHFEToHXhKQWdWyhpM5kCVwBtKkn
yVcAaqb78FZRBsdxv9SMh/lhbWa3YBSA9cqxE2podDyqFmqMJT8s6+X/015PUjWXFGSelX95PlrN
tCTQ3qZ8rh9Ohalawv3ECiNOv9SUo6LFBrhZlLC9sanleLdLDaGBA/613pTYrOeJr12701x4QuNd
cnOZfvi8X1TG+os7yQAQ6Rzoxo5v/UxKNT3cUzoVyYkz0AQeRsYuE8aI+JuiZZwu6Xx8/LsL1wSI
X7V/Ka8jEAfCBZiIlWRW3i8BWpEkfEQkLihjDApG+EQSi4+WHDa2cQ+HQZj0fOdqXa9CTcwlcmUI
clajyRUjBiggxkIeqmCowv7YATtQ1EMjlX2XOPFv+FVj7xvpaxE+7HY91IA2nvc/v8SgS5HWca2G
brkbmFGoSf054v8tqLzFPWShbP8yBMz2A4pbnMybFn7yX2P+uo8BbF5CQJAcX/SEjxR9Q1AQbMEK
SYtlqd41/CMdRvfcVdrt2jIuJjrItQ9Qy9nwL26O0m9b5FLIP+LARIDIEJS2r9nzEgR4mk2J5yoT
InnHCckWCrrCSDROV90nF/w7IGg6Uh0/K1M2fT2HsfeLan6VJw+YwJo2rayYxXrvTRSNAFVnIjoO
EOxvmKA5D3K63sO39n181eWoauEfbMZuZ3vBYPDQCUdyI/cANaj8JYi/0UAdvX6HzGxggU0tHCS3
Nw9stxDsqaLU0k9/EPcpaB/q1qN85w8wCFEXyp5BIfPuEAJYkvaBnH5PNo69IM49G7UdfIzM39+0
5qZJv6W2+rdHmx1YnaQq2ahaiiPyLRZsMv6FioMWelx7LczZB9K+7xh2jKYC66X2fSBZAiijUojT
FN0cpNnVqojpEmRlqmZzLIHCap07IecX4Vp5HEWyo8VG7Mtxxei4oxeAGmDSw1ZOnBSqwbvKGz0U
PwPl3ZwgnmmW4iVfwPCFxInjncNDatwUgRTRzY5xSAzEzk0UD7V2EvJFYx4mfffH6r6NnaOAkmQo
7E+jc0IDXEn/EfGyJ4u33eS40qIcOdvIZt3yxcxWsOYJwPROdLMMcOiULheE6QmxbNVdVzbvujPA
cQc55nHG/q3m2I7Ia7SZaD6OOSPsC1O+NEuorpUuxZWLF2JYD8/9rbcuM3wmakJ5QvbO40wWFLz3
bd81ndkJsfMyKLazcLCgdHoL11pNnmgFS4uW20IjeEHGu3iDhjdpvQfRC46S6lNoomExX6OTHchk
Psd5aI1Hr06xObYaNIfgaarOfcZ7ry31UarBavD6sWB7Q4Ha5Di5k4kCSA/78CZRX1OZQY6N6tIs
Q2MPDrLv1EIzl1jn8asaaAlO2OALv7xQrCpyxNf4mZR0+05w8n61NEem5KBpR1axh5GmIgOHTp28
L/V3Kihoiu9vUuwOyrZhmLlcWsypwM0yixonkg0H1oLEZKMXScCGcsitMIkhiUY/PjQ5N2SBLqwO
SXn/fo55rKBHcHmeFzAN914m3sJokDSgOQvm30DdkOEc8PhnzSP8hqKnmA6MBZd90Ofui4klcs0V
m7Axwso+gZaqGt+8y6E9e0whMWQt6VzbgV5YFv0ogovh1nKcWE64be1KrUB7mlzhHNELYVtbl5S+
/qI1vq/vqyiTHDGaZXI9LNZAdtobclDtPYYrhcZYpShItcPF/rA6iD7qDhZMV97oFXRCLYlpDWbV
NHmuiwmFTKTanwqzDyn/87wLIrQr4ek63HczTF8EgZHKVCLafI4wbmXmBh6+UIlH0c1ZcpTg+LO2
s5N5h4xI51djMchCXO1apEoXjh4sYmOH/rZXMMNWsx6uVofuPAz1IpsSs8p7Kv9OTqjxlXQfFBK/
P+Wlat+eGpgQTfVntv2bCPwcB4kl75BrX/z8ovYJxn6lCvLNU9nl7jO1tWw7hXi/TJgHC5Dt7s4+
/tEMXs+lpzf2tQh13an6f7FuH7w5Y/otfqVSwlp9c/oPKO9JUva6pWQc7bV1gCVTFQVb9YL6oQXP
Vp9l7uVvLVS2rrfFbWTHdNnKNmeOgYhOgK7WPLSO7OAUsh0vgihHMbJ/crl1o661E9E+ka7fuqtY
fx7WToH1Kc0jHKIsf4Ge0QyqN/L3gUdKdT9S/DqGxzvw4mTM39FSGqX/zNMk05L+SnFoEPoK0eXu
6o+FfkEtI5REnoJ0gc4oNDQEsQvTp+bPvdvRCmDmgbsgm1RuoPu7HBrgiKYGWTGYpc3hBxutXzdT
rtNzb3zBw4j9BjKWtgNuRYqsRKza0JFMYryzeVgb9ruxSZXIRHC1H/M4/sSeYFQHTp4tfiG8uKZe
Yn5HCCGaKs2cwWRT+7VwVcVDL/yKYe3RcMTEwp4fbgcyprm7labQo3sp29F9rLesvrHNjbii4hGt
agqXgIp35GuCV6s4eMKD2+uLrDWoPH3kJ7zjuArF2xcU5u+D4fJHmbWHn2n+l8m3QE2Om6zNS3B+
Ot8SwFcnW7G7/GMR7lc07cFcrGfUXqE214rBezgcfVXcnX9sHDWa16VErmeskZdUmqi+JruZkPmc
pha7Z5SiXvhSE4HWTyLP/LpnOuIVLZj10woSxwaghSVz9sD4Vdtn6PxjxSDyxiQm+rVoz7vi/jn9
7j3rEj0Rmy2k3B02hXBFhBV40gBAxKIO4jbRI481w9hV5vB3iG/8X2+zEFxOkJOoqUzqLYpBhBNl
e4NT1Pt+5x8cKWve35jb24w+7mPL9N7fl/CAU6PHwRhIgYGOzSfakUrkffzR+8JnHSKGeTp8uWTz
GhwZApx+u9RRlda0rm5WvtiKlWq9QV+PyywTcrx4CJPSg2Jp2RCO0xqStbLA+pUp5zMPZYGO1yYo
lyPl0XymagNmExJ0pZ6mP4c6rN/UsmXVqUzCMgfkD22csOX3fTlPYtuOhVT7GMhyzHi4k7FMF1H4
pe9ox6yB9N6KOkGVw9BaKXVOpve/PiHwCkt2VafpHqhkNNQtpOkbDjTGxGvqQE4vcxUE/2G3P/hz
agEUXhkt3ox4CclEH42Zf/Ofg6WFZekJdQNOtx24wGDLrf1HkuStJieAexJfLU0wEi1TXDglC//Y
wX6deLUo6hTjPSUuMm4smGdXtMxhKP5A9aBMMWK2ZFFm8wZ0c3TUtoA3CbtgXefwae/onIFvlq/3
ydAJptIX8hROCY4Pqm8teHm35nzRr5lHF/UZD5OnTW2FUcSuaLVTKdpPFI9wm2/tTbUHZ4Mv4w9P
+eKvZEnFOl8TEGg5vEAV41HQleF6M//YgqVkZWVe2yKGgdqOS+MWg08hcdbaPxvAKaQYXW34Zw6Z
JukXiy68MJqSkbuxvjVQbLcy2mMLhNRijXbixeeEUvX3eAC+C7J6QloVDOZFfDQ94W0KN+/MYR62
cpaEi3REWmMQM32Mh2zzX6Otsx/aPXUOgmOmvYgFLUrM2/QrtR7e1ZxooRSfKsHztJPnW6cM19pV
BRq2xy9m/6kwood8vk9QExHl6vQKWOWxm16Wy0+Mn7tlLMukmUl8OaR98CbzfRTREV8GXcKtr8jV
I7VNILNacPNdvlnzkVgoddfymFFo0oGWzSguHuO9vJC/SowON0hfoTikry3Dk1q4Dou1+vSTcEG0
UYU5YP+FHdlVHQepxPKVd+jvQ2Hh70TLW6JKBKlO1rGsIa9KSaGppZ/3ZgDDEvWAz+J3r/LXhGIX
dvtAMCXsbJM2OTc9mpFX9GO7zXoGVMYIW7eUREEb/lnDrGqtSus/kTdVs+SdeeQSTGx4eOl4sPPa
nvfrQv59Oga9/N4FKAkpGEg/RnGbfnlQ3ja2vI8QEBNODdqT0jdTEp4dDoTnhe+fFKRetUEG4oO/
sl6z649AlfWIZCCW09XChot0vrIscl9LtNo7zeZAlMOeG58DKf4psg7hJ9wAnBiqSspSA5STcZDg
7K8+naObk0nj/FU2z7p36hD2Raa9ZQinS+/GbAHS9ajsiROWuWIdGupqMOXbgJ5DzUzbrLaBJaD4
5o/QXepcb59pXlLkzPTBnJRghSdNHrczq/i4k+JxDd7Pm6QcocrUffdVO/fnlN3ERQHEr9n49k+D
YW0o+oTaCfZiv3jqPOf5SGMXxt7zVdrBUNeGGuXv/Kdr9SXtdji44xwJRg+o5e0jPN9/JY3jbJd4
z+M8kAHSx3saS5za+Nzn2pxTcXs83Lv/NhCEmXN+T9rIA4rQs3n8vh6EJtY7PGAf+ngfrK52QJpi
OO4AzgxM2ndqZ0/IVODNSBNbBtPiVHhRbLOssKXeJp8avp15XIFIUx7gDY3Bqv6z9TrubiarGqN0
0pHkhSkO+y+Vngb9fZiP0BlIy8aihlecW2jHSkXU452X00/qkhHBs0AiUSMWGm4H09x5ELIBADFW
2JsCao5OwAC6paMaHEGK/RiqTsdESrAuw5abcGr+M27CkZMRkpepRhVhma5pSvo6QMlQCQZy887B
+yD8cTW+3nB7Uwsbhvs0zrQGXBeG8l1wGnlgEmKrUGHq8/rqZP4mxdVRd4uoBrbHSxT8dnkoxI8e
Pn/BFV15TPLXWMHVWuVXKVSWsoKN3X3jQnYa3gtt2yqpQCynEEIJyOwIyyoWdUzIlk/sxeKUZ6sm
WM4qgIsmia3WgmrtFCaSsQvsEg+SsmwPEiLJXUkyMJTj5mCpg9hN2P/psF/yhTbrl0hzZXNnnDXi
TUQDnLHmN1qRsRPPMjrxjSTCtPhYVmeDttNOVNcIpoNPAA40IVJKFYBf+teMSZZ8kiqAy2yEFdVt
Tz12+BnsebFlY3paq8Lm6d4EHjc5wesSChUy+TdcU/5XvjFBEWQ6DHUlwtjtu9FgCemAfOjAlfDD
XmW4JWPQhsUMArNmyirMD6QoSfn8fGKSx7d1YPRn6ke5whnCRS+/0cwvOLBtEv6asI8nV0yI0zTt
yvGlMpNp2ZH3SSKwpnywKRHzov4IDm+KTmJ86wjxK+d0F80BpV/aw4F7X72H27KSawPzRPMK5GSJ
ZQYN8KE+8KozP6fL6d/4edjmeDBAIMZlyfh00WdPDle9AwUjx9/LAm1gYcRWuTfTWnu9vnEjgZgV
ojW365cCSI3UclT3JJabz3iOMpbNJnuygd3f/Qyn3fprP43DlgDjaucA6t3S+VYXrj7K8BH62kQG
Mx1w4SOI5hXyu2duWR57vFv1TvpHzwGorCf/OvoROSnr3LEFsyFK021SzCI5efpLd22YHTea7PFQ
95tdhztANhJbYVEQlNMg9YJwGqqwXUSz1LVAQ+vHuD0CV1SlhFwB3B3nmMrTyo5NFyScGGTN51he
HD7C/exM6+RcC2sZucPlVfk7NEzLVhC1mYH2MErIR9LfuTxqRR23K4+lzJis91EuIl54CtdfO+L9
oZHV9HlxxQDjq0S7+X4yuM3/3LUb3s2j2Wt66GW+/8XxbSMBUunvwjbflw3J2eZm9Vw/V2mMaWGk
2Y8k0YwebacGrsw9LoAx8u269hsnPcexviiaPiGbIrCSx8qNJHS6bAOeiWx9w544rg79ViOvOWxP
nApKKyQhgFYx7BaOkVSui4ou6GVejowuZZBkb8VdZKdmfYROX8w4f53VlYZtZHP76if3Zvffur95
NrQHBURKtP6l9H3nt4/4Wg/MIsCVkIUpfszOQ1A+JpYQbxzhlmxXzxfpM9cGp9mArBowQZVzQhzA
J/TROMyzanrrPy8muZNq2eyjr09spxkBzeOuESETHfeI+hEzLKLBrP81f8bPw1KSji718NRoP/1l
K9jKUIKqY0sqP1R8gg5nu4C8Kpl53leddkNgVEt6Sxt4ZHreAOdWYsW7mBPbPFSkUfQSsBSKa42O
EJ4V9POzYHsi8pypbDZqlkNZpZVME63BJQOHAyQ4QdSltMv3uPrro0g6ob3lg1RjNxKVg/41iqw9
6J0qHYQJ703wkNA18H4GVaXaU50t2L8tj1GaIvAaugCGh9ksBy9I7UU+3NizzNkoQJU9daq2oJBM
FiAIvMynpkEdZldJNOv3Z084HsoooEYmnjEx5qOmrV8ch75zF8bLl01Fu9b3Yude77Sro84TEHSv
5nIopiatpKQRP8s8wdjgMk2Vz8DfWwwzFfi73dsQtJpAf92KTsEnMEYfTQg0sOeomgoFJrckaI5l
XponQqYkPwFHhp9zWFRThr7W+uVLPkWhOLDKhICwY9T69qgPtQwZFZhMsGRmuwM2dhPPtRWS09eR
0DSS6GwFvK1pfZfcyltMRuTDHJGsQR54DIZSMqfyxRNDNdm59Nh2N2odXQmFECZGnuFqWNEME5GF
g0RvtNKOrwp2oDo4oIecVOo/Pv/j/u/UHlEOmPeKxH60nqxLiGgFYUlBjJA+0qyiR8o6fB1gnPiR
JjgRj1fycOOTCEEkZ3su+N+FxnZU8mj21Wb67wEu/Mzh5g94dPBo0oJ/GXR3kVBa2G3r3rYyJlvp
wijlgHd4QxLDHP4Q2A0f18cnoz+i2zH9a3WZ7lspvPiMu0QBwYRDcOKthjKZIaNSCdruQ30jJVPZ
/eseXjJ6ParQasRFCkEIEj014sw1i5BOnw+pwCLPtl9b5Hpv4AL1VpC7B16JuweuQkJG9slEFyFq
DVhRmsNu3j4SbIHYkTCP/Bt7+frE8zsLkt6dy9TQ9ZBVTaNQtbOhVeQREoc81pq3ZTn0Vpr1kRJR
NXTQu2yc7vWRRv0gA/Rg/cyOhu63ztbuhd5Bwl+TC0en8Gzajz2EjduVYmcEvxuaQ0g6sogiD2nO
HZbd3GLsEghI/Bsoqf2aYZ+NuEAepONSLg+U2ez8HJt8/04hkB510B2AQKnxUuOCabpbinj8qP08
gydzZaLsqrLd59kRrmh9bzNRK5N5bIIaTttxVnEBjW28qSBCZ0l8gLnlqDAF5WXR/R+Sd5Ed6ZUB
s+qV+Xs5om+YirJCIdA33Z6PXiZRdLravytT2HQTGLaN75wWe4E7jTypIhmoOidEROd+IL+Jn1SH
t8ZDdhllrd+MHE4JUlILrru95itZAr/lk5kH6hxCFAE1SdeiBnUUhFY45sIZoTm56DmE85SX5Hx1
31jS3bj1e5otBOTUrHlDna1WZ+/bOn616qnCHIew1/YuVBtkYHLJAT00532lnktVm8e1ohdWYA3q
zgCz0h2XelC0YRgY2SU80BAR/6n4uplaC4lMvxvSrZ8w4+OpyLR3ZldG5QIAEPR5kgLicEJ9wHDm
5Kl43/llkhTOrOCfUg8NbAL2XBY8o8NyVUCC51LyDagh3yUewE+lVr/1O4OeOrSvTlv70VIpN5Z7
vUWuA1E9vo3OZaXMgStjlxwWgKEt9/L5cOtF6Q35bTCw7++poXlDY5dP2Ob+mkgzo/fXNIn6renb
SK75VoDU9HLbSV5EshUuk0qSncLxBTRPeFUSN+6yS0tPyC/jX0jAo7+6gHbWHU92BwVCGWJhFpzF
oYSvzNBmn9RepKv/MWMoMXhKPceLDU/i3x+xxhvSN/pmB30tQgzfmMRnHZfpJAu4TaozCkGUjG8G
VhCymJl3EeSMlSceBDylcOYD8UTK/mCLfLpgzPNcVOwLfCwBIxMsA1NZ7AopSppI1rhuWZfst2ay
PRGPgNhEvhGqIny5GCLC3GzTWi0keWDFizmO2zqYqXHte3zlD+52CRn7UYPqz62Mu7bB4FTvKvAr
YoVxHA8j9kx+aMa7eJjy4oA0pokwnhNUBtNt6h8kgvcy6DcWqlfCfKRdHfYSUEOT/AsapvbCpNoV
4uvquX7shfgKaLvpI8IIeJ3oRFwXC//Hnla498AFLYsC/ZtPVjAKv8Fj+YH9LD+IZybKQa0qEQ5+
EoCOul0cuPBtjNOyGwhf+qd11eZfdQefYd/M061bRA07R5Y0FsfE52A+BXpjVqMnzb6thSEZkZSm
jdA4Sm3A4HRicUB/89uLpcxRyrn733L8zStSWsR+YcpF1ihTbaZ67sLxu9CgbXavWaQTDK+ySvQ/
Dz1CgceFair+5Rb7fMpJbwm8cjS+Ozp/XfdPYwYqfvCbF6Maa4z3BwTCVZUc5kVA0syPfhSCopKe
kW8IxsgVMH1N2Ho2Z1nWKHJZeVx3keuQ3j7g/ya+MCkRRB6ze2DESf4Q1KowcHvnraIu8kSEbHKj
LhYa/kfXlvqWaJn4tkooJcUngkYufoeRCv2HxgLDCWd6Wo3fD8GcQN5LpAFyinx7JQasc2DEU/w1
xp35y886aa/j8PFB7zVRs4NNzY55DVEYLI5dMV5WxpOypGdusC+gaNB3bInokKVWsVv5CQPBRwPf
cEz3eZPOBwDPtB+V7PPrKfhO+w/OzC8qG0I3eekjuTvuFYwWMxy5AOEOzufSWyJehNJhh0Cj+nTs
Ay+KSSNvP13EGaznAweVv/laTLddTOHwa1wcP9u63Hb6GXp4pTt/eKpf4nqv9uhM8zEkCm1DTz6e
wa4pv07/5rTe750WghB9c9zPk5gkjVSp7nBWj5UYMhj8D46pnsBODc5z8RKiCAt9XQjEBShOdRpP
wrhZmwNsLO18EHm3z26DnRtF9kh32HAfyC981E5wJz6WVqU588r6qi97ymThwxl6XKFl6E4fq2YS
JKSrVqXn1tA05bzPD7ZiEBDSOxa4Afl0PxtYI6oVj8v2+aylpTTgyifVL8R3z5JKYDtRMPBJvhkx
oAyHwqdb9shNsxOhbPGAV5IiKgA/hrRHNmPbACl0DxfCTC65Zuc55yMlvQn3jeUfhgobTZpaypIo
T1G8qY/Lb0Jdab+gnxM+ZnAEpoMi7j8KLjFBSu/TzjJj1i6Gb5dvjmOX/MoKork9K31sVjGIiS/6
BY3xPS7byzTdvKrzfACWpMj/gqntcetpCfUU8PgDAnl4FX+fQuWb/aLU06eaMJx4ARWtFtl2vn0I
EP9w2qJ+3o4bqabUQwRhWB6wkX8vuhFJozPlrw2YXiAzSJhsv34Ck922JonNmjkkOzOrHwg1B6IE
YXyYNhj/a85uSFETzxZl2D6CneW0Qj28dN0C17y96bucmKhIYaCg4lptLnvSpgI8dYr4SZs/Y1rK
hUzQ3EBaFMKl2qltq0BAH/9sWL9Jp+wAdQbyf0pMdZ6wviAEkxdqMBAOKyM4owPASSh6TzzF+174
nR3YyLv+7hb0vjTmy1SeKO4FUpSNyOrMILXbfNsd+5BY8GfroLdmmnsk/cQt7Exck4hAd10gz6Tu
fgEByUyv+sd4OjKt5Sq0v1/QleCafi4XIuHpxqYXOtgoyLiRv8egFtVEIKOiX2ntJy7NS1IRLn7n
+6Cwq2DLwVBfoGld6/lf2sxWORF0d+OOz68IQMguxBhGNYVIJ1MmGSrL8wMft7PTDvr/URN5yDPf
Xou2egohHDSMfa207WtL7BKnLF+oQeg2YUXFBZhQBcWZQ+eowwbV47z/30CvFXY5iH8mVlhKFAxo
2nhjh47gxEHIkAS45LKeJAzdkqBlz+3WuZTJAcbWo9PoOflFoZo1uINe6fkC08scfyI/xhTERjBa
lse5idUrhQ2mKmuw3Rl5QXAMxx7tBaS6y0V+k5K4FCf5ap0LZ9EKQ04NBWsev40kcuOfnJ9mBSD1
3ktTb44Eo2XkwvhPuhJuiSqNaWd0niDnkKj9ISr4yQP9Rd0gRiswoxpDR5spqmQFaJj4CnaLLdLv
d4BIxd42TG3YkbBQeYNc/QaYj5gCRgb9ubKTIDewyztlazv153/n600rCHv37m6vLEXVpJVSC3fx
KC4jMJri79zUIGFl8EsI0xszPIaDY+Vd2VZT/NZqjOUKFkkMOR/U5UAZe8X5TRAij/UfxEdAlcPE
xDj8mFbT7r6TMZYhocmHCzhzIZPZ/a+VKiFCtu0cQQ53fYxlA9r4z9hNTSUORpvSbJyt/id28hax
RBtRgtFLP/4M7bWSNr6T3AdTUyzaqkIAMPReyh66FPv+BbZLXq8AcZ/vzTm+zkGZli2hL6sRLbm8
Mldmiwpqgs8IKfUOoqqGVfj2Kq+Gqs5KQ17UF4o5tC2XXZJi7M1NbkCrP005dsDQ6lcEObJ/cY9Y
3ET0yrvxj/iK3GakyoddL+NhXOHoOXMinkalmPqR3MBNZ/kAsAEE57XQwq+GTJb8m+K7XhVg02JM
PqFw3aOV+fneurZYK0wQ1NPKSmzlPbbNIpjmQ7zznB4ez266loF1JsgHMGliadva4JnRKs0umqkO
TVZHjympvpZqcMAVAl28/4FafcyZKVr1dr2fztjUrQc/Mbmvcnj73zPzH+4u6vJLtXLjZasjskr4
xWCYP1AtJG6IPSK25HMZMxkUUnJ7To5JFNSQ/YGsW+2/15CR3YF735/VuSGKKdUA7+3UZqhw4qoC
rwDWOfQuZ3e49pFUqHOpBYb/tKO0nc1hMajslBtf/RbmWkb4vKalxs/YZ8qB6Smp+RQzxs2vq4sP
Ih7R6l5XR73baeMrPhj/3XvHHQlSXNxP8wIkL7B8btv8xt+Nby7BrNlRhmske/C/QV/xAz/eiH1S
vorqZxP4Ak2X8u8yhF43VWnh+frg/ku5TMVEMxNZxkA3MpwoYMzbgyxdrMPNAkHxkYoGGRTu3ccz
rnMKW3+BKz90iION4mz0ZeFKbTbY9+RO92uYc6bzurV5LxLzrYdL+htX0speXRkOh8DhAqek2lib
VSIXR5VWlzsT3DJ8RTXH7klTLQduXOioY2m2/ChJ5mzvBkpCaibRtkU8O40rvcq81blThANodDtW
SH8FA12YeAtZ+MvpWrLLGPoU0kqKwPMimYWkQpNcvbDSq2DISAK3WSf9YoCLWrxfVidBiOswDjJW
zvd/bUgmhRmkilZTeg//ebbg1sIHE9rfu4nVaTusjK14WQo7OmtnnS8SqXCJd9SYu3xB4DTsRU9j
tY0mXjqoklzcrIGsen860bSHkeniznAEKAWHdK0vvjgaqqp8RqGka2AVY24nNMuRNsNra7FLOc3y
rUm5Cg51HG2iTGvZr8Vu14HjNNccFiHDkL226e3Ckvcci9cAOsRFVXPsKGnEjQ3Jz8ZLO3p65/DI
GPAgIIAgZJ7tVezw70CzN9H//d3PsXhS8KY3UbbCZN6LFzwfPOk2CqsY1/7IbJcDwFSCOsysMdEF
9UDbunmhWnpRdvLMET9vWvJHX6jqceYhtOHAqJOTHeHG0TqbyylUmESLBWtr4705AcmrJRL8N+Ns
oOyZJZBQwwM8XGWo2PeDdVBCNM6DFBi9dqYtOGnMp+pc+6xYV19zFSx1rtyDJNY82wFY4rGFSLAb
UW+Ov1G+rYpl4BAcRNJj+Dc2r72bTv76giBump7uwKvN6GkBiQFUhasR1I8UlDuW/CGbtiUh9Shs
xbiKnz6yjMUxHT/vuNRJnoxHvBn8HIkpCw9cKxsPJ9qflzwpXkYYKDC+cIW3uBR3VQImqx1ucole
ElmCMRJOsoXzn+UFq1MvV3VtlxmyMsqww5f/KbK8Tp6UfT0mVhAq0zeinkHNI+NiSnv2zFo1QvPq
3gYf7cGs+Dtll6mW6RyZeL+UTDGUNdbEMd+Bw2pyFHGKrQP10wYEdj3MK5GabTGy+f1KZeVB1M/b
g3uZM0UJ2gpJW+uPZ+L88uPEWxXb9z7JxE2ON5VOv0VCvFXYcRxoPPqN0VyusuQHTMcpbuy5IQ1w
IWYFTPOrpWXxrf+WCVy1KeTdqKrrHdaeKFnai3+yjFFeT+KHNgO6y9D7yuwTYY7GqnhHEASD571q
b+qmkvg0s5slsMuQqoYkP2kXTvyuAQOKBEjhT8kQ4+J3KcqO/+gRsun48G89xpGTlSh3+TSkKzpa
PzH2S3JGt6vuKB7cMJLYomF14oe5eKdmvl8kr8oMqnAnU2gnEqrAGyNsm0hveF9bkFvWpWVwWs91
nVDA1+TtUJfIW/hcBHUpks9uCHZt/bru7L1coOceep/QAK/cDA+lbWpUlQ1gv2we0bGZDc7Hlf5S
B6ns7diy4Vp1Ig8x6BDzDI83bkSv5EoJ8/c2Ib5VAll6paJkl+4ImcdmbkvHJokcz/xkMtvu6sod
EsOIP3KFzLDaP5FXqhqXWKkykLNgClrNswsKTGgFnmeulc7+kG824HVcr6oY+137fkQ3sAQKALJT
0R/1xzG6ebPWWNBjB1X+ztT5r2bv1IQbsGX02hYBKNz+v1SOIohTACEAsJR5q/IC8qq2+Yk0hvc0
oDL5uMx8yBE77yV3baw/X672y6neuGnyYU2UZbezGC9eK0742r8J7y7URF8gMtgOfWeOGdsctHgy
UGphPX5xlP1FTdiGAzKYmo31VXd7i6p1Qc2cGDQ3Jnc3mx+iXpcslqXMOHttzYgiEwUDSwwkL5J7
2/Aq2M+a5e8qNIhdhUFH9XzQvSfBL2S7h2OKYotkNRq076a6yT9xB6NQ9eJp7U9C/JlSOLh48Ig1
+d3QoOrkgi1Fm8NLi8rAcF2R7dfQ2qbPum7BW10bzNUXNYrV7gGRDgG7dcQdoa6SW6E0Js7xRlde
RqudvNXKs06gaXpSMw4hCINeyK5yQqmXHTQcEuUdNsm72ewuIke0hWKRXzJqLQxw8hshBcW64dYN
RUJ3Bn3A+NAmmwjm9y2AnKF7gzkxd7wJ/U/BBpIuB0qiNomGj4K8qf7/mm1fCyq2lrKu5pB6JJvQ
Ad7yTQCAWyy/QVssZuzzeYWzzjiL3PVXt+0EUVzrAVIkTFpX6aNOVf6xlK1X8LD1TdIa9q8HFYLQ
7M6wLTCuWbZqCrFTpiS1bhQt1/Abp2snfcKuuPObnSZAoBl8kpzdEoGD9JKAmW7b98ri+X/XVFXH
XUlzm4TScKWfv0RHkMazSUMOpIVr3YZ5E4q4ilv2a96KPmID0pjlDp6ZWN7xDS1kLcyw7nNRV99C
P//x5jk25Mb6eaUJt6ZELBHB+XEYO1xTqn6DLu2cbHC4mhL75wSAJ98z1EcVqdIHSACUJXBtsWwh
GWbEpdurSmj833/aFUTmXvkiLARe5ojl/qyclcKWB/JRYC3l9QDKtfqzTpo+LONckQqecJx4qd+h
2Za0LghQmf1ZuudS3lr9xVZCHs+VdibU2LhEKjBg6SO9rQGjIjD5ccTj7AocJKJzEja/oeRJkKkd
oH2WnWfPA3Nd/SpJggcCMybcvLn5GcHlKX1DOXycKBgubgt4uPU3YXoIZ9kpyFw/gKKf72OF8kdM
4l58cYHaovlnwDuQxaWHfzCbQoc3uMZ0eOdi/zJhQp6Z4mxnvdw9/pisIcwK5EqHFLRHD/A2+xUC
ecFLoqW8gnwmyAlNJ6g0u+636taRNp0sObJ9rLzly0HmFRZqhRuhRkRKVZCIfid7JVuNFY8vWV8u
aU5yvMmkhqzKz4bm5m6td4GzDZh9x9Q44gLqOo15YrThyXNthACvLClMzV+h/N1vPuMuNxXtUS15
T6KiOqfdKNZ5z+j800ccy42noebrX2KRoUy8IMfx0o2ggfh097PtQsROe1Tc49g4ZRvm3fUGSYLx
RIYbueTbsESqj1RfQ2ODGrafL4ycW/DLtSy/eQCmyAHGYHNR26XABjfKRJ6cmzc/zzPvrgNHKL5g
lNub1Yc6WsvO69CHl5hYCpQQe5AHhQKoktt5xL12GfvsRnR9esAo1sOSRmiPpfeDGJofNT+s7HQo
GZ7sL1HSBZmkIriZYbU5ACuLQF87treDtu3jpuCddsTRbzeSiDaw+iZ78DDukOTNPu0lvW3mjq8Z
2nQg5JITcuU6p2U0AxVBbhyATCisZOrk7cJjGoMe7WwPToie66LvhiiHqjuJUavt/0D9evAXqljs
9x/0E/KyC/EAxMN0EemcPiOfsN3be18VJJOkvXHMyAgTWTZhFkn+F2DLDbkRMNtV/qpeXfEsTV7N
vX3pkaptyq/dcNp87mdrjBKV/atDdX3QgTZiKlwMpCJwTcuCDYFx+fOsSLt7LmhRSrDueJtQq9KC
Ioqqx3udjGILa1bvGmeINO97PoTx/WEbwGwcApx3bBJiWAyoiRtbyKJGLpPSnMmh0oVOsFAydNcq
bf31Xrb0BvxU/g0auK4LzXd2vggvNx1mZ0Y2//D2hE2HzZ3X2FLFWB7gaByqkzjv8oxfmyTm97/S
xR0bJNXjiEQ5893VRn4KZNjV9Vx7lMbLfrNTrOmgVhzIDHTaDt1bq2Z3Hj65CA8brMYOqp4QEF4P
XlYpR6ysp96yUoo8dg+Wb2gAWwnU+Q145GZACB3zX5WCEj9eqFkqQsIhNHgXkzNBxgaQXrzPeBSB
B6Ek4xWuaBoX8sZYXTIuFRiGKuolBmM4U1bC/td8Bw0b4Eupip0NS1eY5dIqlX3oc6UHI0EyoOks
T+voWu6qO9iEzwAHq1nGlF09/dOaKFqdXM15dPIFU4PhNiYTr/U74wYsyDH7nR9YgHxG0vEvL05I
czZwX7z24p+SEwLtj0N673LOfjWPqgq80OL4uPBgjXl+X9MdnlwYNb6feOHu5XnFRYxpC5s0LNV7
8yyx2WYgWUBTDaR2X5Giogq8K/OrTEgJfZbfRzOqeCKL9CFLs6An+gxrBmzcX9cWxXvO3r5JrwwO
Fy2mVmUYRIrCs8N/n6dWdpqQppBOn26nnoR4SkRe8bZossABrXmd93auXf+99O6AJzpoV6kRVjZj
PEs3zNpo4Up8H3PPy3PY6qs6q9zC7nyBNeRt5BTFYDnYjYhKOXL87h8n/p+5yNqFhJ4g+9DjqPDB
Gix35JVZjsaiOZBCQR4KukfpbgULVYa00GG8zJot/I6Jtq4jl9ErbeeSm3kIrRQE4wdDuUC7uWrY
l6Pqhat+HfkZSeOQGDv8LmHDHeXCbg0zy3dXDgD2kPCLXExkVjWzrTsEPa2Pj37WRVR5AwuSQSIy
xSPt/jNiRLfj4umdwbn1egLSdKZAPHKJuOyjojtfkEW6LXIFhCFIlSOViY4N33A45za4g+hO+E/R
2+aNWbwHrt0ekbXTZPCcyd5YwTfEK2sFYXyfhKF8w9ADVyDsEQbUGz4JrIsqqJ3v+Df/vShChIGc
dYcK2fpWhHF+Y2nqwK97knN4T0+qceS6uPkvS3VUUe33rtZ1YxwldcJv2PgDS0ePjzv6nheBc8kb
XZ+v+Zw/NUJHErB1pvR51W0q1cLOd0YzDpDlY4QclyKTGzeSWszd2QJLD+RpsnUZ9P30d/qS0W8e
YQgX/k0mHsvVpphDZl7mcB3pxLK8vdae9N6hknX1YZxBQasCDuiEcrSdlmrbqoaw9MQhYDhgFf62
yk5bBzutb9UAcErgvmuyVCW7nV8S0US/EP7CWuy2bEyQt4DY4BHuOUhXbIuIPJTtokUgua79AaBy
fVW99/+8sDSdESo64YaGqtico5Bs1wqAKHzUcmFJLbTt9+fcJmh3LGcTPZp5/5xN6nKyohnOA6nf
cTao/fQmTLQByUr4Jx08/KfC4BK0tjmg8yc7vetF9VeIcFu06ORtN0VlttGAGw98Nqk2nyumP9yQ
GsWji8FNeRoS9L5H5mbk1jvyrq543Ry4XaJIPIxa1P899cn8xRGtjMqNYvw698RxzYC/sV/YiobU
0jtHgGCnCzdWuJwIw6tm46s80q1dT5hxDpEjhs8MbfOq5PEHIMftuFL6XdHQAlQX5oyjjN6MHlei
h5pk193H4BCktriE3la9eFgTOq21ij2/Oww2gJoQWhSzjjZFVKH6If8FbWfJhdzAGvXynIPR/Fp2
g7IUffBt5uBv/hHUcIncKseyzt7y5BW99+oGOPs5AeB1wFCbH4gaSEMMwjjD85IsIFE9dPdPKIbV
ZPPCiHuq2glJETjdiBkVzX3IPv2XJpiVeNwdth5k3LHbTl2xFRAshmmXEr3jIU5fCY1UoaQVFawA
hdwh4ZbfQxwPyz+Saum74p0vZM20I9W+Ovhcaqzy0OK08nElPiXN5XwawDFLO0FTG+svsdsnG+5d
BLQA2QPqDH2ZofbVufAaOUafQdRlolWC5rn17FypiYZjnJTneNp9/vaF3giFWZm2dmeW2tg4d4rf
iFmylMfkpPFj4QAF3AcMSUDz6H6iA6gxkob3zM4AcQx7iWutKFrCJg4r+z35XsDl2+bc3IVPm1pw
Sg4qEewbL57K80bhbn5jDuFWLwI/9g1y7/7KUY7q58GeWpeKU0j5JL9UPzSR9Cuoyu2kDQ8hi6U1
cAci3iHBLP2XIIr3v2AyIbtMmUNrZ7ELZcy2rbHnJdVMFvUE9NSBAxEdDwpyKdIm2DwfdM1T04hw
uH41sGx3sEPqFZ7vDZoGVWJYkeoIZPgvLVcc53oM0uN9ASBSqMgkRF/UG3q80wyZlNKTB0jhq4NL
+G5whZLjbNWkJmPJNn0kENEg4pjYFe4/2A2UgnL18BwbjbjJ7QvqyFa7NpcXo5yICPnUzCKMN2pl
BPGY8lpYqq4A6RNGkvuqQPH6jfeRE+mKDzZ7serPNVC6fBHRT3/qBl+8mWRdgNJvtKmmqqYquQ+O
S2koET7OntUaI3IB04JsOvQZFIpVDLlIiUGIu5UUJzw3+6w7sRg2waj/sRRo//4NxUNYjnb/Vpvf
VYFgYCeXLzNmpMoG2YLuhEk9t7Q9vQeF/ODYgIYWoMLEEXcsQt0BJbEceLltwevQQhKwN1/ULVZu
Bf+EIoO9THr4XPvcP+fr/0fboEcUjxnn3hC0WhEYtd7g4wj8mwxSYNi165mwdLfHzzfpw84TzSsa
fQRLsF9jBBrYyBI+YH5LbRUGp6qiaPsDOrKw4/GU7Wv1xbwaHT7rVKqAUuJSHhBXTKr5RQ8LMn3Y
itzOGJDKYSPc8g2rO2Wdlmt+DtHN7k166AWW2AYheHN/wNTIhtHJk+1Xn1jYiK38Wh06Qv49r5mX
r2J0JDOrr6ChJVf2WTmeAdN11aFtOuGuM6/mOJyDDk8YvexGCpx2htgDsuxTEmdNh2p207mfq8UY
XuDfVpB7d/7CA22Zi1gSkvO7SqGHutKXRTK7NWSzS+CWZsCioSnVvcz1nmDBpZ3FWK7zXBF4UwOt
Xc8jH0X91OVi3IdY1n254wsAohc4H8asVg3pcKgID1QIPX2wvz87Q1eXQt+5qVGGxTAD/QV9GQvp
jlKC22+/v3Dve8EnEIfkxdZA2FiPeOnDklJEftKPSWRXucle2anPV3EYXTmM8RiONA0BSlEfQdtm
kVeBS1WlOaCY6jiseM6rfYwWdMCYtrZkz9Jj+7AC4A2e9FeKGuh/ElZZO28XRKT5GW1jlxu0hEB2
PXqu/oJvZoBukn9I1fgwY1IHR7qONs8jgetjRCQNRQ7Y1Amvj8v8LW1JVy6tlrLdRPI7wI+dGmak
oKP2CQ4OmZx2cxs+bHU7Hex9THE8Sf3EkI3z0g8Tp1m9LQB6mVYZIhKhejmkG2XW6MJDZ8FB5Ax/
QNYlt7X/8TAfWo+WrBirrk4TCpoYPvwnEhD6u9yU+7El42g7uPZoYet7rL7K24F8s6bmifW2/mi2
Eav3SWMWhPocNcF3bG4L8o5ddfiDZmLbq81ISeuE94j8ItC3uTqNYiMfSbHd/T6VkvVwB4xZH6bn
4GKdT/WQwH3eXd7WlmVANK65aLLgugDJv5Y+FNCklPJAxv2m4H3+sbgMhW8MFL+US95pQOMhpq2e
tuRE62WAsMQHLmA2SBIMmBkbhNbb6Z8W3q/K0WU4SDmGTNGOmMNigppcRe2acHMisGpxte8jBL2e
1MLUxNOu71Ef+09a+BmURFHLaIpqu9NcKbT8ZtJmQbfRdYUfTa8kEKhbuYc9/kqs55wKbayBNb9O
3OZ9g00DrYHB/8RwgPS/8ZvxHZa4A9UstbS+tBp5fls/sZeCq+wwSProGH+cyQAS2CQ0XUNrTpq5
CvOAqIaRGww8fnClvMKP8DrQ4I/cF415tPY94P0fLW6a7Ma03Yjmr0CdWBvqPfTKRs08aBcd7t46
bHuHI4yi2Ay2Gt3sM2aX9qQvcUhTvt7qYyk2ieAbDTWg5Uo3sXTf/sMaRNg9fVT1O7KH8GxgNNUo
lRo1Yy4tkGo5siZH8/z3FcSBGIYsDuQN7XF9crKM1S5SP3kuBQHsoYdSPsonrA5GkzJYOifRvXXv
u2K090UoHtl0mqdor76oVEhjiD9mpRc5FbWmYb1136DjcYyYe7ndWild4flRwcLWDQ3Bq9NpFjDk
lUaeocFg2x4tK3fvs6wjU8RsY7TBIWowhgTJKGeP024KBrG6aO+byQa2dd/fSOGH5O1uWN6tNJPu
03jNDeHo5//kHn6cxB2gZE0hiVFQBrTM0SE6M8p2va0PujJ/FZSD4NC5e6r1AZQqxalqhHG0ySPW
fkawMfUYTRR1/7oqJPdaY/y9XAf9qxvrA7Jh1d1HjHH0gxSHHCsREiwpTB1/3qSTFglMSZ5XXG04
Hbtx6WjTQ3+DUHrU5xoWl15Y+RDZfmEDISPAaOXSMWTyGBk9WicO0/DBibHc1dfN9px5BnuxqvRI
RSSD5Heit3g6IzHon90sYL8wPthl5oL+Cqv9wDUSJgnGq1hnvdaWioulOVgpClh6mNilMukZ5CRN
AFmOHneS8Vxq5UesZzEL03Pa8Ip24Jh0nMPBY1AnFHVCyuY8nk3itzoUvUwBduKSsY2PtvtTtKKl
7sHmP3M/EdverxmiAl4oPbbGSkFDapWrXmmDnQbGRSsULXBTHy7mPhNhOICVZcB7zHTTXlAqfHk8
CMpAkl7YvnPz3Dv4h4Ca2JpeoL8Y6Ggcqckx+b+ageiUVYxBEaMnim8YQx30YhK2ojD2Q/YAeTfz
xlQM8hXG24V1GVcZZXQ46CTu39AWXuSrGcY9Tj44GfarvGi+BVok3sdwYpN2lVZxeqeRa9QdUYvl
erkaP3H5kzJQci3BlbiaVHjwAuuXS3UBW6kDFMYtaSdqUXskfoGzStDrV7laaaWAeONA0gfCpZrR
OFaE9JUMXfDWoyp9hO141/A8nX4SNUeghx5iooqtJX/zSxpKcAauboq8AEj/EMD4zs2/7kx19qHU
S3DBHI8ewlwOVr9lUD6Aw6J6zrL4BtcX26C+9uD6B8QILM7ltco5ULHLYx7H8k3ANPXgycHGEXgY
SS1XH+SwuoYL3i7Obn+hiu3/sOBnHTLa0t6e638I73wqT/qod4WdVMbfp9g/vYH3S8AhenR8nDlK
pb+Lr55Oxfg97UqLCnbDCg9lSRaTjnFw9GusE2Wpa1FC047f4J9KlD5HPdO66FYwkaEoNuQs+bHg
KTnft42zO2bCuRp474vM7zPOQf4VUdIZPUbJ9SC/JxVrnm9IsnT27yFhcpr6PoJaBrtAR7D5tW46
JWSX7ZBOJySA8Wtq5BqJdFHXbzxt+rVXOERG9uvMXbB1lYGXhwsrwBqhcO9cWVWbnJxU2BLmfI+Y
Jexevwqy9X1EyJ6ot9HbBiJimyt3INsEcO5mgtteeLa2NX7mTZOW0VXZbQMi6giVhkbhWoe+uRD8
6a95MqV0izh5AQZV+n0FJrt0urcClpoa+xETXDXIedcmo1buiJ97yaJQz1SNNhFKvYCo8CgRYf8U
OgF8P0DJWBKI8MX7pweh3p4jBusfWFxps2KQLyuIxKUURiJuCAxXILc5XFrNJc/+Ni9+H+Ro03W8
MnsKxVhkKyJ4xn2eXFBtPOd7ZsE6Ppcx9S4aBMC3S9MozfT605jZtMyPGwBzZnLUZ9cM71qYG8u2
WaieIIWNVU6EeoRMJyBLrL9IeF1MuxAv7F1ngtJKf0l/UXMpSvzet45pK+XDX99iTDnmEUjzwnyr
n7xrBG6H0ob/QHk3jC0Ep87Abib5K7r5ALtNJT5QbAhRcv7KS06onr6s5NzbttUXtjKQTmmzupQ/
Ff1weaJQ0n8dRdGw/zQCcnOte9D7NV/GL6vO6keUooRmkOcgThwiEVTpLevYLhDFflYOgimcXAYN
sdGs9GDh7YlGV2tQ0H9ss2lAALNjwQmtdDam5zZP8C8eNDs259cLWcJqvIhYlMUde61coFMgMZ5N
HiP8sTs6OVc7Lkm3X9tAKakCfq10l9DbhSuEv8OgErSWOSAxsRmSx6uxlCZrMY/gxXBc1txw3tw8
Nnm1zanFtu2jXl7rz43hF2El4HETxKTuVT8bupxwvbUICYXXPSRcXt0D+qrarD4eB/3TLBGP14zR
YP5argPHcRATiHgcnFkjP2ExoMQUkJHTdE+CUNeQihdCRww8Op2Pt16is9YBRe/OpLALEI8l7b40
4aU/9rp+4HjZFEYJtdD/kqGyPytjl9OkFo2QGEYNZxaG4AFY7hG7/H1ZSLhAlF+psjL+htvmn9b3
N8qFLwiPkOUFL2WNpJxazOVx/NV+mRkHvEdkUm8++DYOJvPJT+Z2c2t0v3EKw4Pg05+/uC6dmMlh
b1deSVE8MATfTh8bT68/6X0MAf60uU+tfVH5W0UBabXNNsRnJir4TEGatRAZCu8IDH+Rizs1jk4l
qYNKbS3QhNZcpbDctQcyGOhbbzlTFjygfRjRvRh7H1nRRuoIMBlrEHGtq80XD1qdjt0zF63Ri4YG
39PX2XufkvxzDW4AyW8uRug2kTP1Y8gmRResCNJSSvi4DTx84SIou0bX6vDcsWsX8lsGip5rw1r7
RWJRjWZBYpCAyABp94kQR1oBh0DOJoGFNjcZa7KxA+0UnWC2GIvcrYj6LUCYzYt2Zhh18IyyMaxc
YuWpEjOtShNxa5OokgU785uRxe002tCi8ar0CDN31tcc4j9ENdhXu26t87EIVngdHCN6nbqpkUMj
2eE0u4uHEgM0SiC9T+mL8txWtlTIGV/LoBNdcCOTqTMl7eCU3BE8BaKOIPQ8NLmQ6oCiWBC3EyBB
JkBIRM2fZcXoyVPo5dg7f28N5uGcjn6kp8ZvDB2OJquznWcBxnLoE7OLfyimAw3AaVOoz46G9C5I
6fng1w7BMG3sieD8xofrP7uTjXN0itluW4XSr5T6GIMgARc+Kg33bOjWJu1j32EWiNWUVh9kCqdY
f/frDHPxUpQLRQ2Dz22iWA5xtkKjmtA7k7TwJ6b4V1Mh2+EFYMgKz26Q2HzzdXp0Va5i3X9dU2xI
x8e5NoGuehwJqPF6RykAixhrEdi+K010QOJUa3hgjxhNiII9wcje7/5ge9AY+B6I7iiqz5RZehhG
DBE9nTcY8ZXVcA2sTMef9EjU4I0Ugpm+bF4n2NtW+HXcElEtj6/RY1tdIN36dtBhqCEkyT9tYIB2
gLRuUlNXIz0EZNofeX8wKqW6JJfwTzeYShTdgrFhMz0PIOGEgeq/cCs54vLkPiydpKzXmWKZ2Ocm
yFWYQ0jsr2AvYt9H/1Un6u/mPMYBPr2YGiZaKb0p4uZKyk2LH9I6OI0NB1NdDjPF47M6R9Ty8cBc
E9E0p3IddtrtUILbKtlCbC6yj9KtkNuHdlHc/aQpvkL9Y7LkNMp14ceDNqcIASXje7l3MQpAxjJX
KS7oPgMYuw5E5ztl0ydVLkWwp3pJCBnfSlCdi/HvDz0u8seO5AdhLn+yETVLv591BTMhOTSH0Wjl
WtyF8UOz6hgHQxnnWxE4ahWH9sj/4MaC6Y/VY/uw3qnj7lMY0fePun1VY424BKqZJ/tGLXqYzkSb
6mwZ50WsVVGbMSE4eN8G7g1IRdAC8bKyg174hmL8vxK+iHQsSLy10i2KwK9y1I3p4dErtZLno4jF
8ivKHjAlVELkA7Y1RnK/RUtPqw/6oMSe7szOrNLRnYGS/EMmRacHo7hC2Y3voeB5q9431x9HgpkW
C526SUCdUZXt9v8Cn4Re/Dg9RnCKQD8zq9IJVW37y68Wu2Qhyjy4PfPkD/XEJB4jerUYfUu1HpoO
PA15B3rm6WwEfQeFV+Kcmrmdk+PBs78btwG2nxjCy7fW+gR+tUuuLw9XOZPEvlJETLcHI6whQpUH
AO76CV965joz9YUrVEOELxen7EoLEg7lRLSw0xw3kBssCMGjC2TPJgylqM1PIHuM+a2Fl2Bzc1V3
dGFyRSuiZAAtV0rwWQ5G0AQvSQY/PtFFWC5tUNGLTNnguEWHy7kIRdfxWz6TfUhPcxZw5CLMBFbi
JEKNVPxgYI+eJQT4rHXe76ngNVPEi2alIukndYcfWAS3CtOpls6PjDrsSWx0EmM+x2b2LbPC8/i+
6KLq/Bjy60nxbYsehvdYl0H1ODVQf2SCp9m1wcOh4reNz92uvbz2C+eMaTKTcv/SE8yn+VTnE8uA
PLEv3N2qWwGOzfrydcgieviWhXCFBptn95nhbyFgH0Z7uoe1tVaI9nmNP7/hq3rTQa7GIWmhG4Rd
LwB1UUk17qLBDQYv4tatTQdjVU5r5tiiADnpmYcqVfjDLV1uruJLeLXTXnxGcMmWmIdOPWFhDICF
vKH3+bqx/wBsUycj08UHkGkdS1O2QlMwoH0k4r6RS0gqnb0l3b6kX029n2obqAKbrYYspA37jzGq
EaOB/BAyTrWNcFeugHocdoaIPvOjrqVGfngqQ4iumf4vlXHZng+r2hJ2tdzmLeJ0V6+t6pSYBtSN
yJEPYoELhtgsHptONDAUQwcWUlw0hmM5M8prTJKav2naV6xfPgfOJqd/QNza8vXDMXz4nOYPzFaO
u0GztQHnJNeoKT7/3eOZD+7lbAXv79JGhT/cNKW0+cbMYbvQbcj7WihjcKmeFGW3bEsQlmUt50YC
qlNRNgooxUX24GSx6PLN8fjTokQu8dV4Ss6fiFwskOngbYuyw2QlRfZ/ceF4ocfhMawoXCCnOMnZ
9Mcl7TXpK/71zVdtVU4IMQJUP4BgkD+kZbgGKo56PYJLzfhhrdq2BVszWf5zJO29BL4na/dDuSxf
oTE8FNNN85fxyJuhM2n5f39VdYXoOWoDHog40GPafo4sp6YNSxM/ujk8h7XYMQgUevZAG93cpUVo
Su7ll9OeUXaoB3Yn1/W2zsh/RMFeeND39f2QxXD4wZ3W3hJWoMZioAR5qM2ugbeI7pauTANL8Cmq
tPoN0wXETMDE/tfn1qjpOn4mDiz1QIUPmLFbFrrqS6d/K8BuGb3YnGP+bCTgdBoOnxxfbzac1+TA
xEToHCi9obRvd7dRgpVXcvsaPh382q454EjvUoKp10fFNAibMCI3AV92N+ZRSfU45LAZmfdj8A/c
onuANa464XYMn7qCmkgDg6+xcB3/gmplSFaAe27YKaIAZJfV8RLxw9KXr1x3YHwaGX5CSYMQ+ojs
2vA01vlL2nWA61olvqhD5ah2sXiGs00PPyJGbKRRjlUE22eRgFamgJaAPNte4Cq3RYFbhBQTyxnE
DWLQAqbcmOizxh6PnJbcmC9vXw4yNOiRjtqLQ+ZYe173S3rso9cE6wQb8THKRympbFXcXI3VoLK3
iwp8BkLW5nezag73mrpYJCtTHcSn8kq3vEIIjMIdXfUds8u8E3we6Dmpxpu05NWMK79q8dK5/VRf
0W/HRutgtndy/AT3VOX1q51aZuIfRrZDkrvgqZhT5ub0a8TNfK72ECEscqO/vXQxoTBVj9+F2Ezn
e0LFvkGfHn1T+4RarYz18RGq06ubd5oQWxSpyeHqsafepDUdrCIZI94LUYhuTpw4Zw2oHr1fVkJj
Szfvvwo65mGyLRZslDDmDmzgk7XD0vW6vLa+GovWOcXKFqwcjICKfPYlHzl7cKaC8iMQvSi3k+uo
P+vaCfF1S4ad1vlCVPNWMV1v1q8xS19mKL4kY5IVxQG50eU9iq+pteo5QjmP/kcYpCKzXLxUnwsi
RtVxpIlGzdMgcgrmX82Nb61ewOdqWwaGgI4makmknqv5wfYxwjM2QZRq5NO1/+6bVhZrv39/7ydR
N2Kbnzn2eQ0AWZviBnC2K4vN456v56scPj0WGaSPDdm8Oc3G7pl9BR+S8j7ie9NjKSZHxM/O/EVB
WT2xVIEMNUgkaxVFA99KQrNvxYOeRxWapvFIvaAftHzrAfWvpijEFV8SY5kDoJr46S9ep8jEQhZC
BmJ9YIWKYeooibWlsfqTqZmuKnEeU1gyHgjU+d2ZaZDy7jc12EKxRJw8a1oEPGY7pYFEuSseqS/7
w1+t7/bdY8+xTGzDBsneqFYV2Lo2nr2OklcwYfKBebE1wV0F5nu2t9CGc2FLw+k+4/ml5v1zLkmZ
Sb7BMqZpqHNtlkRaN8lSb5mYkXGpjF/VHBTsO8uWR7ddw1G4z+EjzWpapx4GOaR4N0vJqOiRbx5J
WfowpPc5w3xto29sPce5FPvGapFpp5vk0xemtwWSkoJ9TrPycYTj762oC67RxQEASP/2RCzXOiqE
/tCT/+InUuFw4HtDJyc0My6EgbJ3LYiC/PzFeVUn7PHYYpUbsQ/BDYIZSFlMbar/KcNuIKfT9v4z
b7Rjh52njGLJ0z9rOXHAOioBYGC3v1dBnrOeyDno83eccwRS8BZSy995quMf6JHj5/kU3cH/OWLG
nLF3szRbryu8SUxpzJPt7w1SxABiiaZpj6dLKJMZm9u33s0E1RMb/grIQNny4Bko6j8uxfJJxxGE
iCyBr6BdOyF/+aosp9PimIrjvnieR2Gy0GtuFd0QJUuj6Lk8aIPEzwZ931Rv6iuo2f/8O0Vn+XDL
LMxQmnO693NCGrWDHSeOSerVVVM/DHBmjcI+L62MUIJa4DrwQ88LxngVPuMUUszDdAm/Elk5uTBU
KEJkNlp3Tv0UDTSFDKBz8+kzhcsLldCm05r47wpyrY7tkL8HCv8MJwr1DpmVdsvBNWa5sCvDuWAo
miUwYD4nU8tXO8ewRLn3lyiHpDIz/sycDMYNcu7jkn3lEmDlO9hEFAiE7OiHHm6Jrnp/MPMfT4US
wGQCwgBjdSswi1QCJR/8ij3NHWc9gWZj8XqLMh6rRboOALCxGGpEoMjwb2gIOsa3gMs/AY+RqjYU
iAWRGRHvhvjznUUEzSaNX4YxK5dGqWDnUGFBIJpfChQTSVohI+cUdm+1dpKBidFKxl8NZbIK1rnH
Oo+HYGNd9MNjiRA/XCw/sv9rapzNJjc6PFVa6GbGRCT2jmlOdhLx394c4UWEfMkAsqp/LlJ/IPhP
rsRUw5zL8qLOubn579OqRudEIY/MKo2X4k0i4xM4+7NCdYOVr3afI1oqXtc0B5u9kJPNnzxfmRKx
zAxJVQt7DmS69EDAlD7HsQPg6YC9hz/QHcVPwNzFXE8seQwk5DOp77TIjLEXO0pdeiWJdeRifBho
jDc9+3Rz8BZwYmdNNLauYS08v31LsyF7sIHp/mnZP3owi/Efm+O8+GRGIW+aplp3clVcM6htkbHz
awz8DUvNphseJ/5B4Mhv83wZvC473VvMGjI6629BsOZWdcedtSRiaSu9ehIX0jKlQ5YdmtBKnTBz
8JbDIYnNYtjWTJOKU8NMJIhaG2v8N4Roc1CfsGguXdnUrFnlC9XR5N6NWe2j0vtjXjWV4XHeBX1z
SS0PXo/rnAryVOWFmVoug2dB4k2QF2tjvzHE1NwdWi2pQ/ggMlKJanp/zudO48z2knPjp47hmHus
n2fXmKxHs7lxBOue8J1vZJMQgSVH/6CcfBmy3AOpRjx1psLV2Rd/R1PUBEhsf8G98Fwu622iSveX
e1lM5KSuWSwjoFK6627C09QrDUKs1ZYgv7FfhfkXEqgYpifPlyjVfmahBT60WXLV/Q9wH3gCxswR
KH1aTza82s2E81eSQd6qePlRdyMZXHsxIRbZOq/fyL1eICx0Ub+nFvx3ilT+kibSCtkNbhjTP+Zd
AI4FwNuxTHF7I+2gDnaOyfyZ7S3ZpAfufSj2r9pwRwMK0wBq+LtqE8muKYv5NrQVemrN5UdfvqYP
xXKQBnj+XLh0jeXjQ5vDDC56WlX7PvRoxd8v0PhygwrDwhbIOaPBzhkBxejPFFp9+CFFYHT8iQSO
X6oKtIpzIlWxo/XWKUBPXoIKSP0/779fkljW+BV6UuwQzX8LSdPZ6zsbk1jdvDGZ9wEzt433KYV4
o7CXxkjjC2NTwjsKp/Ek6QAPBCrE+Bwy2htiizS5dpK6hZLWcj5YHKPbeTRsEIbZfFIA7YHaVk++
vvHK3OVsOu2CT+DqgXW9eVLzHgPLAkb8fYQVQcEJcWh+B9A7XrS72kqI+Ts8zyecvxQtAW0GjC7o
MSUkG0ovgsD66xzEJYM54CriKUhNYdYGnyzK2JE7x5fvm9Br3BwOdYMgd9uOQ92kZj5QWMQ8af8G
iarytbJ2uSJXI9n+cgBoW0AnFck9iXvXDtiT7A7UAiIRV0GqWqSDcuW2vbpAX49J6c9RJAQcIfov
WyGh7HazAuKglmLFE/T2NSSgtNQO3DesedagkNDuky4igqr5zDBDzDjBYv/eBSkipxN8Mav6XHIR
+3QUHjnl6jnKv1Ac+xr3Rq4uThi+QHkEFX7g56NzxdFc5UKs/YrN20xLDb6297liVcgSps7jfKzs
I6Sgw/VNu+AII+IYkub+kskREEB2/n8S1N0tzVGMp6K+UWdT9HcF1a+/N89uq4P/V+Dpds0FgTXe
e1f2EPhh8SUza7Yvj5ocA2fhWinYClM/gu96sDs81l46JXSim2CZlGlclYGpTHdktZyC44qSdJHe
vwZg+dMKoWE/LJe3Xnhmuw8M0zIoBoCwtlEY3/0LbUTsGNGOnLzPH9xHmnTjQIX1kaDg5UBe6AwR
NpG0jUe1Xs+IER9K5XR1vNPATychigI8viVetj3bq1ZzPG6/VhjNOvG4AY7+HTmxyA+3Ft5GkgaI
gl5jXmHDiSQSnO2tnPIZKzdp5H/BcSfXg8GBMszwVdIbS0WdMP24RxwtKOK6pEYnicwajELYTeDr
33yQRxAv2iTZzUcWiPBfpFFKOSQLdxEqnHxm/i0HukkwQ0xfeKi/41BDBviPkbr/OU4ifpO9e6wp
JhE0wqTtWQ2gP+ReqUVMmeGO0XJeQA02DRvYmqidFyboeLyVIooChEIjWDel8m1VT4CzHZRVKjFV
U3VghtYzhQM+bjP2kfRpu+HlLpV1gDW4KSoP8LcuZgFEIlrRzE4am8kSc7/aDprMZ01LqHV6nxS9
Tz9/t2ezRhRSWxK5R+7vdgRO+jXPbjMWGjOWyBKdTEQ+fUCoew6bnM+JKxgO3GOcAl54H/fYV8wU
DGpVZRKRNowecWBJgPNnFgYmfmvS/G6nxZLI9DzZ2aB2qpJO+sj0avP2XNB/HbJAz1P8mH0U+L3O
t5QOA0RlSmhGp0OJQYsZR7sGPnrQKzk8Rm9/vZ5bGG7ComNHaYYUBIxdTfO/cH8KCm+0ua66NlbY
ct7pz/B53KL0vNHKnZ2ZM28/P7y6A9Ql4/Jet3EGDFuhiWp2LX2bW8jS3i+kmDLlsUm79BtisYTI
jwhMHjmK94uSleC+xOFCxDSBaYH8/ELk8VbGyuOwzP2vrRxkVpT4AbnvoxPIQBx8qqpZJX2daHVA
pQ7J5QOBGnO1wYGtA9mPDi6n+Hgc+Q1hv+C5os8n3++QesdYRlOJfx7KHMUnmFKFgJ5qGzXIUiq3
b/jnyg8dthTPNOf9Q6bR8zgZKI47aZr3TzCO5VUPetgIGAuU32CU6r69posVFRKtWfPjqAmaG0gY
ML1AcYexgRrQmw1j8Zi0WHjND1bmdfTOcawOwL0suWE69n8CH45DWkgr33+MBXTk+y7TqF5Xi70/
ESnwfLtqbS0gd3YEzNbHT0nmiBuUi5CmYMIk81nEzJ9+5PC5oBq9cKzOgpl9A38+l9sa4he3j9cs
vmGB5E3zQV4cFo76PYLj+WwdcwShJEtitS5PJyr5IA6BRLVXL8quYri+1K24BZBjmliCg/Wwybp8
uuuT546WgQdVY2BIVAJz3A+RbHMnwq/Ixv6CvWY1PCLqHlOlhGr77Qx4xo155UD0QUeRA9WP4ccs
FwNcRUdV43hYw1FUtsMkXK69MK36YHv0qAR+MRgDS8/EY89ywUzAjOcdMDI3m4d/2MPG5WoA+5Ek
8NS4W4VTba4aolAfydAfUm/Iadii/GvI/NQlNzXPGUKxLQlmR1N7ZPLS+zNACookfi70QJC61VsD
SgJSAi2xlc5CuYXDJ7Z3e0NTaZqBdsSKScAq/Obeae38sYVvvPn6nhubtSNCuEqTNb0nfSFV58+j
mBPWcofEu1ino0DJFhGs0aMTgVYbdcCPetCt6gZ18CJFlikd7WuXI32kRqscTfXd02hODkLcihod
bj7yMCgHtfCFIoUVcX55XzRTi3QzL8pPWTpW566a25hGdUiWHNELORdt3PQyGXbAR46CTLWIT1Be
wJZyiN+XOsf6z+WgkR+QBOBneFcB6KtuZeA/ExERZ2uHSL0kx+y12KBtU5v3dws8jm0C4JtkuRek
4CL92pW+7PDO+QO7lN5cJIbT/rCRWPw5HIJ6RfncsSQI+mvrB1c+kAsVEePCILMWOdbYoa5tkhlY
MfAAq+rcTeO6BdS8Okctbr9tcyB4x0X6s4nnkvtys1N2D76FGhmULwGalhpwbt2JAPt0LoVSooZB
AeN8q2RsLDDO0cAEojoRIZr7mI1+Ti3xnkLbFI/BxeXVL9dwetaURalXS82q2bwUklcO8vfkaNkT
pbmOAlJLiaMNo/LiAs3OFkkxNgiphrD6HNwM/Tewfu3iszdwFsbtb6SDKlEy/aft/7yIXSxAjzmu
GQZ0mUauS4+7wFL4t27W8d4+ZOHVv32S3YPTLifg4hqDR2PiJ9FFPs3bLdwA695/7nSGj96/+6Ux
GS9oIBdJTUDa0OIOfLU/ljA4MZqfuu+UuMGjEw55OoYhu50PT3sdGAtdtMMNeC17+Iq+m0HuTSCf
P4YVY3rtJDmlzoduHHD9HQlCYmBRwSFYPeIXj2c1S6Ca3KgTASUZQQK0owC5NJcx3OUAPnrvfJXY
XCwUjVFMqW4ZI86Xb+EvxVSTUT3YcBWG4DJMHcGSGfwEfQHteGff2CKWhygavPsctc0e/VYtPBLb
rPV5cxmUsOYkQAPpJ3nVOS9wrGgfmIcBvEbsiWR0Tu5HYCpdoK0EPKM+hqgfTk4EpcRlEI4F83dF
LoKzReU59lqROsUreuzdI62mOO9v/zh5BizopGRpDGzV9rPv51IDL5PXDxkj91xtkGC8mhiWh14b
I2eEPLYDF9/FgtTtk+UwHXwAycKuC/Q0PefAM0+s2zFBtyFcQYe8r0gCbgVkThY5y4eEcyA/090p
IQgvCtdzh6yMuvMQ1GnRexOC9NqWJRIGh6Yv1GZniL4AAl6wKz2Caae7H9HgoUWPJaXZbEIVF9cR
AvWTusHEQesQQa1ZYjaP0LvH1bXuliDruPuvjNZ4vfCp+a2IPFa0kjvM9WVWn6deDXIEjzZ051yB
45CXcpANgGFuggaIuy8RTPfYN0b9h3bGy4QbMmSAefNIbSSKqWZW+hTpM+ssoB9q0T7e+zC1R880
AtQP7JEfS/jDs4KSPf4EZsD2eLe1t3mjSW4mOSE+GSKTAiH/E3UcL6EXB8RW1At8GHIMjNc9aR5p
tZrO9aLDIPIGxCA1zhlNTPlsFwzCLJQKC1BP9hTRGggW8S5O6Pc05SQLdCa1VYOcDMxUCl1FeCsp
fJJvSsYNEq1MgJD1967Xso4lYTsXVXbUfy3XrbFm7cXTHrYrDVZ7/bgcxpGpk6o1bvpVvMyngzM+
Nd5Xp3UyXW5nS3zxkcnAUmPUVqC6/CwZ8NPFYaytjS2msbewpW6rZHIunkBKPf5EBKD8X6xd6DF9
pT4w+mEKfBvKgf5EgH6Nhj3v+ewMfUKSMccu4rooqWIXbvxKcY5QkZ6gcikS2VHZt0nHRQRFvmud
VcW3hWUqsHF94mELbNQdQUKnlso6yB3xWmIzbSME0RIsNmU1FddjD19P1ME75n6bRAqzLgOgIS8+
sX7/5ow+eI0KCWCZkokHSzX4v3Hmu3koy2pRPvnPsalPlviENvQk+0Ci6Gz4zldE30I7kOBQhrPq
XC3hGw8FrR5VaDxXvSkjcuWSNvgFVGIVBurzzUbCRFgahp5nVVnhzBxSnS6c/6eoqFKr1rPpigLp
ruKdYMDDRT71nrO5zPBB0HVEMdigPKCSlj0EUiVZsMh2ul9uAuKaWbsrsFtSeVuihVTBO5zI60lx
2hp8xVQgG/76eS5u0TiT8BA1Wvr4ev8aWiSIeiz363SEVm/F4GZAjFRD5g/LML8FLEurqyf0Wlcr
pU8+t0hyAlNVnX/zTtfN6G+7eJezDyiZkT5IpFvB2hWaGf7tGmdq+zc4WW56QFSKrNJmt2USUzwa
nFWTDrBw50dXZZ8MO5F9f6n6YvoyY8mcAg2YSqOdEyKqCYG32lPxvlqt8KfeuupWSHo+ATcG/+gH
2Y5T3qVIS/JLJRomeJq1b56Yuh/mahfDxvypXFCHbG7l2zWjkBpAk1ShdybBZBf5BXpg2Cr4bTk+
NpKxr64XfKx/y+mlxZG5WUbnv1k2FaGwPG9rGWhNaKhWE3u2gRIgUPQZbmuyiwyfzhEDaiURvKva
vi7TLzyOihj6gQ91SPssCKNg+5Iy+tLjvVKm6WJqXRzxE1hbVBFWjyqkOhKylRn3uBuRInW3AfmZ
yhNC79xwkSsslE3X+fXPQGe6xZ9T6dv44Ac97kz9RN2DTEuPMRBWvdbYq+L2gXe2FP6Aj2dWmdV2
nVp8I+su3SXmiREBEh2Cef8a2fflLV5WFNqgDxX24QRnMc8CFPQeJimCsCbfUwNoRrxEdzHSbRrY
OcbAlbnKe2jx05c7LFOkHDZfrzbbfw5LphGI6pJVcrmfWDVaqYwk9FzICraX/IqmpZ4yveSKtyLi
VV1vCrSpie978PJjziEchMXcnE8xJ8/Nw4QxrCb/V8HC+cZj1IHOaylhEY27Lkt9Bq1I+UegA31R
r0E5bEKdtj5xUq/kRqPLtB7jBqYrkvvp7f5P0cHBcKQ30fUW/Co+MeObqwL8IuaWiA59JgZrn4OZ
pr7aRySJjAxDsUAnhiGK2oC3AMPfq7MHVjF8tDdT6C8SpSSBV7ELLeA1TLWka/0Y7+V6G1uoAacS
YIkfcDCPxXHO05pdSeuq2vj7mpl36/Xxy4co5WSl+uixz8uhK1Ro6w4VjWEDPWuUTou9Jgk3OoeF
79TitOHapRvBpWwXzzB4eAoYwTpXU6WYgSLpMYyp4Bk7HzsJQqW1uJauwzCzXJ/tBk+WDGMMqssG
9Ch4P6NMYs7i30g2i/vJ0ths4LOYSEY+xc/4fBGfgHZP6Dj2g4YINJyF2+xSVBXKLmaRlQCPhIXV
qxmZzafeQIpi197RW+VrhxypnXuZ0uwTllHgoS1ctXRic6Y7xsxsuLuTIjJFw1vS/HUS1DL/+OGj
k/IuMVgvSx7SxWXgNmDw/kDPSA4rRr/zu3AG7YOVtWNKH9e2hMbn/A5zs6zCM/fetsnCnsorYy1l
OQnflm1F3qs6O+q7hkrLfKe3f+wgqSG/1G0pn5FXMow7Cd0JTDBhBJ5sZBLvA8bZeEyiX/qr/hbE
ZHm8tOvuxq+SQDOUPmyehMPhLnDPCmvq3UB1fRUp6+/7LKwLNJlnM/fHL/MnVPIKA2FvTnf8DExO
NmrkZlse4Be9CX7Mt8FoCC97DhG9e10rfQdcM6TpiAAyfDTAdMnfZpXE5vk464t0M12bRLOW3Hus
B2tjBuGqfbcs0y3cZjQy9TaRVxm85pJ1uXJM9WKPUwPpNPCMm1dMP6tu5ggGQ18svlCUXtvKGi53
iDnCCog+OaHAIJsnSxb5a8tLtt1uAKNwmXGi2xm3rMmojeYnvH9I2DwOUKxrUWWN++5A327HWbEM
+/MFKoqRubaFGS3ks9NTB+QhEiL9mUPnZxImcb9dIw10+jUDthDgQJiwYepAGa3nzq3Q8zQR8cej
vGLHwtufEdiMC2eRfoBvIh/tEAwoqGvo+beU5q4UbMCxygvZkFCKZkKaSPI/q9HD4HDsAvHtgY+H
gz4KjONW3vGWf5zt3R4Oui8eC8Ybk7myEUhQHys/h1JB56T40Sx+cds1dOOiscPTvmV8AfWcLgO5
F11SHQcaMOUZqHMa6ywnmP+4LYAroKfCDAbV/0YOaTNm5LwTXFq4f9hOc6ykbDgy1tVsuxfB0rsu
OUZsheStVlTyxfRMNzpRR4YhphBalgg91Uk1qQGE+m8LWvG+v8gArqrWInBWa63mQ/9GLapeG7Qf
DT85vEe0bwM8wIVbloBZgrwKmc/u7XCgXsnfXyBedWj6zEke7ixGfLM9S/GuPYfeDqhvECsBEMWb
/rALPFOHBLVbfYWnT94Gi+2qSmsmiJzxZPh/uuee9Q1N7a6TCfmRuI2OQyo4+6CLSM5wg9piqNH+
pz/VjQn0y17bjdiE17uFmU0B0l5/tXT/3VwntkfouOxnM++Pp1P4313Kd0T4S6HPlo4RPyjXrP9h
Q9nq6RNgK2UmUlVXLqD+WXYV9Du+Fzjhk/dUUcnqbHTQMGAaJVbhTAh2HoHfd6EEMbfSbYcF83Yq
WLHSeAvRO+YO2Sm2pXF+j86CWBgW3ze+TN/kBI9hBgHh2H8YGOlTm5slJRSrsEHxJfFZ5ioVeeLY
IzkBuBjj6AmeQKgLMJoQWu3X9cfeACEcMLVdi1s2q9kbobpE7u0VG/SmQNolUJPmjBL+GE0skv8B
l2uYBzRR8T9fqhfN30rQwiO3zuWzMuvICPp/1R8aT1ug8EkqDKsTwtUUktpl5tOBUuyXvmr5GQP5
P05dlD0Z0Ld3WK/GURNqVTCKLUn53gf/3T1owetO8jXg5Wi9BlzI4jDKfoM6R6g524w4HI2rIx8Z
PFK4dxc7e8HaBsbzS+6LvK3CoKYZE2Qo2xZvy1WqoChCF708EMZkm7xryRZwRtl6Q3LNmoNiEPCv
0J/lxFHHZ9mVBXK+o7AN3eziKxryRhxbeAlgY62neOboXkPAufsxfAPuX7Y4NcnhI49J6nw06dlo
dKqbZkvGkNiw3O+ZsqwMqFRBLW+pg9r3D60j1P1anPOIEMAnGwkUizg0uA56o33cZ/9M22NkowdP
1mxgRsJQcL5nCNKzdJe85ubqkUWzug/544hp2nqD9cb2wpo5Ba6Vp8cwJfC8lAjXQ9WyrefBSc62
/PY/gsY36UYgRKHju0JbNHjdM6/zBt/DhAMxvm9MuT8LK7ReFP33VYG0IXKOXJ8+D4v8J+3wIom2
aSaltcsrl94W3PAnf/7c/j4wYEbpr6Iuej1So3Qf8lPb6jpctvSFivEZImRx0LKvqlP7aMpn8IQ9
3H/F5kgRPJdi2h+19X2QZtuihhg0SQ2D+d35PAlLUOLTw1SyD5id/wTyvfcRfJrp6/RmbN7uKTSh
6Lctgj9hlJiD6GoZ6TOs7xqsLYzJdwj702/2PdPPPfTHCc5e1AVaMwrQeXh5R8Ex4tRrH3bBqsBc
yEj3b8o9JdPzX9LRMKwRKuLqmrPmHU5pnVGDk21pZzR32iwvIydRIc0/iobrg6JU0tVVir1rAWSl
74Szi9wkw4Q3CAOZfp5liWlBt9RX723F48Ck788alc2XJKWv2RNJh+YX7aHaAVKwUWtSk7LET+e/
n9viUKogRUF/FzUfCnXpKpoo9b0/CGUBNYmtXa4WC9e2fUDgaBapapDqwCVFWWKd5XS+Yj5Xv4Lr
znvQTrBdyxaWPTzqRHsJfkik6EQC3ntfwG9vgBpuL8YespBbEqnjBGj5IGTnNpWp2pLyAjW978KE
bf/CtaNFCjqulTKpikPOxDuVAttaOqv+VUNtCk9ZKCZcvgtxzl1TQlKyiePKoRJKSukHHuDIDnmI
RIyULLjj/8nqhKcvZ0r0raH3PPM8S+oYldC1PEtXwNj6G8lMe+bj6QEpqlnJeR1rIZdQW0qlg3V5
Wo8rihA0tmIssNz8QuUTprEMqIylbNph/Kx29upeMRAVd8zXFZe6Nn1zxUzIkUnq8iHjws6m0ZxY
pUjcXeA9UxtVeo1Kca6enpKu+Fvs4D+xEEd6KEIcuclV+XIsipbokPdSV2/OJsACvtsInmfXHX7a
2RuYgqD23fIo1RCZYbZ6G3EZFJ1LsJxcnhLJR8PwTeWmfGKr/kBcKttcS/kL6HHXqrRyWUMsiySk
tsIpODBAvhp4vhzvv2CK15sqTa0+Ydx4jLjsaJhUN0lx4cEgFK5lAUuDjL51d3VGF6DN8tFzt3O5
saAtqVUvG3UeKA3/MiXdlrh/Aoyzt6UV2bsmgEU6OMi48f/4R5lVoTJoVMKka+GTAz0VDvXJ4K8w
EFKwch1xQe4vEYweM+fmsLwCDdvuVjkb1kKTb8/Vjx1AZu141q3P+krtHiz2Fg0u+NU5lLgNfaVr
EzNBaAWsdQq8R8/2uLqe/GRnkwLJnNxav9JvlIr/EOmwomWqybtPpxCC122ofUse0ejmkSIYXIlb
z/xSzRg0KRNdAnODp+X/RVHe7KrUXZDhjwaGdWKED0XxHIYsoeZmhj1DuNpS3cyspRtDZAo+373E
W9rlG1Mpf6qDuYNW0TJ4N/q32RNP1NdL/jxBzCvvyAYf3rTCBQQJa3LZlpebuK++eVMx2RaXX/I+
UdBh5TUJUUxaixy5lxqusYKiQiyl4ukLz8HI6B0pqi6QDP1NDc60ZITdxMIjHjT70r36AvxEvZPX
kL0vLkma7RuzfUDHAGKBuGtlSHGRQaDiIE+4d0Qk4WTpp5lUnDdQf1mpxLntXbcPwH3zECuRSB//
8nN7JBUlvlQDpKWS0NdLvS433uxuOUGTgvwx40y9vIfbwcIuLJloGoH+z/V3wN9oSvMSMTAjY6mM
2i/5mOTqoNdR44EnBepZQydwzW91p+vGZEgW3MDhoFYuLA2Y+bYw9ss5wdPQA6j2gWBzAraTRaY2
Jyf7zbkJev6eSdo+dfrQIZtHVs/jPIGMpOBXFyqV2WcmMC351WiOofXVHcbNP97b2fE+W5Efbh02
6W0AYj0X1EKd+sp4SeBwndTQgMdpkvdtAT+Vi81ckeVSbIduBzuzKW6U5hLnwYZMpZW+SMGFoX7U
tqE5GySBf/kIvNNXJICD1LIbHuG61ASBHNFByO+P7SHRfIlvukGiRaVlqwx6JqCoJoWtWbjnELq6
Y5QRifRy2mZaIq0YzBYx+GnOy8btBVrrFqE1IEaoIQn+6Kl9wwFI4CXZOkK15uDNY4khr8brIuVz
a8tbt9KU+XtS9K02qGxK3DOcUG8dyQ4kzlE7E3K5yKf/C3hMqcIhLH+ZqM6hM3SHZq13UE8B4v6t
v2Ad+hy2kYpfz42YHVPAMQ1aq9+OxxsgjS2wJA/eSOUfpfQzkZPChXh4OApZ52l9SS/J8PjVhZjc
NL2uocqBrb3ZK00HugviYKqJccKOAwEEYvr6MSUgg1NHrPKOFiYAWQwXzD7wv5IPt2zbm/dY4fMP
xlvhMm1hFRtmjxcVtGi8enw1PD8O02VBEIg1Ly5k+1Ex9sbGLocy3IdRXJHBr6n9/4hvn9HGUayI
QsFMvkLSAV69hu03nRr8tqkS6RW6T4gqu/Qsu2wXOtIsApulwjioRzrMUj9TvgGN5yZpoRzPeTlo
l+AdYgLcFAfsv2OeAv6vR160eztk3tAM4dJvdbWJvVMVefPTrN/gR92HHaV1w0cyBlV3hjJ3qtJx
BxFQlfuFPfNPHUZirZL0VmnFB1dajmqUxC/MfuAlth9+BBC45ys9CnPyT0oAtQ7rITtRzb58AkXg
ZgPKDeKuReFR7cJgE/UIygnpNBecAzqP5PH/A52KaQ4W/2V6VSCCXxQvrjA6B4TcbwamNFsmmOHC
x4pQ+y59XFNSpmcDEjhS4C1nZCXUEarP8alFfNoYlcQ5mkaL3qY5L3F+gpCJD5nX5O9VB5VC3ilm
luCeGe8y2RMtqmS7LKNlof+WxrL1PrqgOCPBwXao6OgXLCxn0YfvbAAjTAfygZGCXXnhJfzhXZW1
od5LXpMY605QC3ml5b+Nl0RZR6QdCnp4o8df6HvipowG9mmhrVft6Uep89CkQakfXmPXyK7sb2Ap
9gRz6me+OqXQPRziapp3ICqXqtPyogfUMiXamX34BM7bJOC1odnkeshPHQu1yqow1deBPRpXZyAp
oXKg/EHBiWF/LhNogIoeuVCC59FVLkBnRoqjrwpLfD11ScVzx2QHgEk8E//1GmVMtdc9HmaOTgkG
tTsbodkh90CH+kOfo4jQjMyxBipD2oe6Yd8eSLo/oEv9F51QKogqCi9dWTsbkdrO3CpAWs2BxzXY
9DlJ1G2xIAmlahJnbg45VqTGDy8Uu/8UCsRLw9fx4b6iTat3rPjKWzwc+yxWiuR3k5Mj1buN2ojN
LEyjNG1iHmgjFeXwwC5BgBermy9zRwtMHNg5icHx9vjbZKglLxrBRgUADfpbR8Lbpb0LSn/WSbxX
R945//81n3UxyEX3C36D/TX0g9n9KYVAqAmBomCuAuifln6WrPmLUy3UZg7FL1jS+NobKJkatNUr
rVBpJ056sZW5tmWgNARw2LzNonVgJY8Zr7pFEfgNrR6pxKckre63Q+FEiT8C5KsOrl/cPWi79JMr
hmlvD+GLy6iR1POg+Pc8xr5wpajHCyvzK0GVEZic1VH8UCoWnwxjfRm3wwEujhwDJ3MpjjN8t/wn
InhoL9KCufSrVelYr4xjWTsm0hkP5KfktH+uPgp0NGCZKP9xtr2tBP/K1n0qSb0o9Cj7h4DYnvh3
M+xHFGQBxRG65kx56RUeWYguKQlSJa+6LHGsbYJsxTa3/wfSMlpqo/wceplq+y+fYneF5rZHBaNf
CW0oszsEsUUfZLClRCj5Ho44w+9nrv+OWglWdb3tZ5y+8lD7GbvsmQPWZ+LacC/FL5MOgj6fGZ1T
GPjQrCcUPAixFrSLUF09UlJYKFOrQyko2+i1b9RIeSaxZIL70Bs2lrmiMAduDv1rVZ5HnOD7JJu3
XAOxNhrxcia7wkUl6oVB3m6I/2ZMTXWZhjbRByELD7Yk5+Rg9vdOHUT4T2mkAMFFPWMawleFWD5r
Ih7W4Y4YqaiGfH05vU3Mix/RkemROfF+L2chq/Puv9T/4XiU//yQurPgzb3wrmcWwUXCrcT/6cCl
IcJgJxkjuXhAAUtT5PG1cAkucrR+860ZRc1FLoi32pGMI/MQjvAG1eKjqDURu94ZoY79ZAVrU+JA
XmFuzdkTcWyXcbJWRw8nsC9MPlbH3H5IwR8aPdobzrl4W6Z+5/D+QU5j9pfMdHSRawAiFnCdVGzw
Pm8JQI38pK4M2ILXSLwwmumjWBG110CDF2wlb+Llg/vQxRbh3LqkmuRGTOsTdjO3NFpFcAEQBy1f
o5UDi/BxEYINfMDMsG1iZz2JeFGIfxtxgH3n1CuCol5qcaZ+lH82EdoyrzXXZoJnYIhijtbK3Q8T
VHktTIsn0IGYMFJptL0LJUUgUB5useqc7tbcXZGKQ5fUNQmvGXFSpp+3V+zMJte6074s170CaQPv
nZHR4C6USDCa0HTLatjhRbp6I7Fp9vri2GuhZfaawpCtuELnAas78Z6Iq/NVtR/1l94CIoJisNe2
LkyQil9ZVjP8qvREB8DV3wXD/fKjV2T0NkKIEV9gZR7dM2wSImWhcFf2JmAIQ20++WfYFRnlula/
Rk7j5lXGfbVyOTlzd2aMMZ49kXRQmz83NAGnqwoqlRUfWEM3/1q3/mx2M+PJHNIk4OpIDGN4U2Ue
HPFaN83r9dLfgwpx8VqpxxnSb08PRj/UELYmtK7vA3zwVpSifR+wjx2g7jfNcYFBLs8+nYrFsi75
gbGlxDz29RjR2qKaH69fVGzSU/bTbd4FhCCc2Qpba8KwItWOKVnlB4U39pFridtWlYJ/vlx6Nr6C
w7sm2BbypXHbRAMW9KPnXR292QNab36LF7m2GSZLwOjnbrpTAqeLWYD7sUgzEQChjg1NV6BqBqwt
fZfx0siZuYLaf744KXBJAaqI7n7o/90PbQ5gktYpnBm45FR+77xtXnrjAHdNR+JxlYFO03UhSbH9
ppLFYM2MM4SXl6hbX38zP+OY2QVjA0vDR23hg0PmfupoRdLcz6P1pClhJofrq8M9biyTN3YigogQ
H5vld6jcZcOT2AQq2vF7OVnVei4k0gRAlKMV6DW/5DjdrPWl+usSJlgu/OSfDrcFnRcYXObphgWH
w5Q0pTIZQlowX4l1bx68bkledKCKgcgNpJVdsNdeZ1sXC3ON2uWnMA8okUMHYXG+i0TL/YOJ8v8T
WdKeAsVf/46eEhN/lilLRrtv149EALTTl4dVVY9rWQM1N+M1rJ2ftPMKoB8NEBSbbAJAiXiKBVkG
+VFey4uDgHvCSEbqegoi0J3Fe4PqhNQdpAsjQ7YJADaDHX8RqH2TowSUaRUzZutYMfAFR/VyxaQ1
6AGoTe+nrJfvxrasPsBRNQa2wdYPYbjAkCnvLkSUMzSMMc54AOUa5cunq6DZsUuDbPSSUkBsVO2y
jc+7YMGDUjXM2knjW01gdXT6+rzjeSSNZeOpEVCB1cM7QY5mqUUqIFnPJw8024V0XAgdYIs/hTFp
kE4GUP0koYm7Atg2BnWS89nIPwdlJHsStjAmXUyJr1VXPCmPFDsxGX2J/IMw7ldisJH2/VzgMENC
l9f1NfV9qUPQnzu9PhjtMXL0jORJS1TiRb1IWsSJrHSJHBAsaN+w06+EqlbmFuJliX9t0y5lpDmM
jB10K4tKZLATOm1AwDCJ8kQti7O3bTTivxJ09qryZ02obsD8X1pkWtH3agnck9XMUWi8QqZLFyBz
AzQVoDZNLJI02chQhlWV1qzAKaKqK5MAdZgmNKUYVtFLe0LLfBsPt3MTyUriB+xEiy744vE4oyc4
NqJBPCw40G5kzaO7vE+aRazHUcEDDs3hBFCmZ2sztxhctEoDDrFP4jFcl8z3zYWiVhUS3IrWJ5sj
W++8QxZskdb71E9+CAjLtxi1mQYRVZ9iCjxDsj8JXoUdCimNmdaASPig6h2LsFDTHcxSWmr/djH/
Pktu2UgcsLx4hxUFDfiwS6tO6kON92ksR+j2TPxe55NHWQfqFXmbZxZZcL1t5m0dhat0pKm2fhQT
y+Qvg7I6bFs1A7gZp6uHOrQuISfBHjH5tHc5PceCDIwM8zEFrxBtzn2AZ49Z+AAuWvRli3q8RcDw
TtzNPhP+I+4CDC1Oqz8LjMd8GjrI6RGoemoKbS6RkNHteDrZuf0yqWDW3Mg9pw6JY+sudEILmkd1
/qAVLb5r0pymZRsHujY7SFU1kU0p2y44fhA1kJ/sowrsiq9eG8ssg2wAJxx0QdxO8yUI+rkJyM/G
7EWmQr3fZcZL1n1WdxBXo5HQ6ubg5+/gW+/oxsfg61hrMPzWBfJovvgK2meLNnhX7BRrqie5gSvA
Aja+cmrmS/KqGOxfeXv31ZfWTwHWSDbkv+IjUYtSCqNaqzrd6iSY2uF6z0x6zMPqgx9eTbfcafFa
iVvqgxDl/bcj/dA9CJeFbUhV7U748cFdjvojrEggUF9EAxiq2fDaPp+sfDvcst/Z4iF+BGMQNh8x
FIWvOEFaCHnV9vPdwkQvrKukAaHcz1XGtH3+lvhG9vFNPQi4Z8LIuJ7bi46lCEINzbdYc+moMStQ
NtzhfHSU2aegCrPcdy3m0FGOFlQ8HdKv+L+axqRyjfmCHc4l/J2Q9rlbglZG2VzUbNst0DxPN+f6
gMhxJSS+rzyL7PlWt5BRxmhgLDsNIAsvMDROlEjwuBltVDj3jYra4OotZ3FMdS1iUaWVhBLVE60e
f3vsOWeQ8xiFWR2goUNBNTej9PAvHn5bRGK9XPVky0MweNVmXw5PFbRTzZ8Ypk2xSLCCMOooA0xj
umnyLoRQl015c1Hz03UPaglBQX/GAjShPleYccptsVzrngn97f8UjbAbAd/SDb15T37cm8Xecr44
Ih5sSbjNLm+oqp5ZWIXGH3Sh9Sy+7Zaznw4IKo4Bnp98MRu47rSudJUMd0ZR2r4lDf8dl14Hv5Lk
n3zmZBL1UKM6be/Hz4Lv8f5Zy3sr4Prv7W5zj7YzFLzqI1KdqQy+oKX9kcu3Ns+6hJ8bCuhTcZWu
uE4WTqMG+Kj5TKCdGbKsGhkFa1thfdP/akE3IcVGrFQmdukBaXPW398ugDd658pb/DetGFKJFlUj
rRDicflLIarxrO+Vfol138ndUrjDpbcLg3yVEct9S0QVCw39DZo7gv8/FflG+3IAMQrIU8lmn19I
r+qOIXa0eAXGdhnFMG3umOKMINzezwJMrrLqm3XBDuzr+pO7izErja4WRbh8vfnEdGhkmjlLgKX4
HcVUX5xQDXImj8oRtAtypYfVwC+hFXkPTwf7Yv4AdZXXsD/W5iAu6gbS3UGhtw0Tsrg4bTxUyAP5
demCPm2pNdkWoi30idPZlIeTcTchuOenedDhyuJFgIDurc7BJs4DnZvm/OxTQSPiGg8D+o5ierjo
FH1Ubpa1zAwjQ3xZscwohIgyKFa/OZCJNUiAtJoYoYTlTVYrgB1yV4ufeIDS5BufqjaoxHzP3J+Q
Eq1WXGMEzeNvWbiFLwchWPWXLt8Lp0YkT64GBoSGcryi5a9SYfesQ9QhIycqSDjrvnH0wGT1Mxsa
zQlzzFGafhqYgwY7+eITthg2xBCtrYtJLjS1wNCRjpr+h/O5T7M3JUNcjm3s3kjRlTDwY5Sh2bS+
qKvmzJvca/dMXLCG2wvDi7xTTHkOP33tMA/ojYbtsw2YIzgleKMSgI6EvU0PUEd0Jj0J7WSJtGMA
k1DAVLQzw3htUg0tHunRbhY2yLH4B8LUE+vWM/5Ez5MHuvw6oqCy8IY2Oo6Go/m+OjvJUeAUi60K
+SJaXO6nONX5eKuY+8oyrHNKQ52N4S4ciKNDngwzWcL9mKBn23xd9+DSGzCSqT5qvVRmWQfZho3V
LpZ9RM2u1jq4P5RNC3g8vaj0R1rPEn6QyouOut360rf5vgvBBAAY0Au4B6UNxpZ5wYhxRbpsqbGE
Ie6j5iHRsvg6twVdzufko/q1hhqws/R7yOZqUawWKYMmLPpFTxu8WhTnYccqHN/TBW6M5rhjjRJl
J0AD1c6Yi0uncyUTjL3cbySO6qPSmZNFjjsvDKSiTnfr8Ct9zGWxQC0SJ865/goBvpacAE7qKkHf
JP4GjPxJmnw+Q4KvltBkQyyVlZ7w/GZ62sf355ILTEw/12mdG7PINEMrQwtXNDHvTMK4bNSZtzXf
fPWKakmHgfCxQijGiEiN6KDPevFGr0p3xGzJJhMFAC53VV6iaPARj3IU8PnipdE5NUnGf5dWssbN
ND958w7wUhcARrKFf2A+K+OvGlhtLOqY8/LdGwtliiqM4Xg2sGnjzn3b3HmH5VjCd7evPpyach5T
3Tg3GR2A4gdiisZxaRuAkxGAOx6hyZnHzxZazYLbxoQ6iEFLclUT/Ds+/5vsYdgBJfTD+Pmj7XLe
CJOnLtUVb6pCvcElS/pRIouGwt/XvHZ49rVGsMNeivIXc3Ag/mqPKCh8RoN523g5C4dQ5WKTsdSi
gPE/8pTFI3lFi2WJOl7g0ZgUTXesOaKhLsaMlBZ/Y/nRlyjHCwq/NOteKWwhPSeRqwZT1DM9nHGT
IZ1tOxlhs/+lXH0nBolO9ShDLNTmGqqvhC4wfFVg+XLrEkx7ZT5uQzt/KhIOJ4hePvKcjK6o0vHy
3+TtpLsEeK7fMOQ1NYFDYgv+S2zZIs4koAlWgDpI3qP6IOPkGYcdA0pTLeV3c5g5Y5lKsIk6ZnkW
VnPRjSE7B4kHv1NcKtOOeWBU4pleepV8ZNSwnRQfmJZHnqh4JuwkBuBoudBZY2jrSlC01DFJrDBD
JfDCZAM6kl25CrczuuNNPpp7y6c3C4npHBez0ew2ykKQ3YvwTC2GmkoyVM5LDLKIlGwq4jnpFrWj
pP0qFEgkfgcsyI6EaJCSJ+zFp/jfAvwLWEMg7haDrwDgq6mc3ZxuV1XcFY4ysJuo0upUfsRVKHVI
wwbkEHrkEGI1xirrd/yRoRzEJBG/lHDikgAtR09rc7v3qNLGB6lsiZznXo1DCAMxh84O/ljGou1F
tzsY4TQqmJ6jCo5LUyGHflksdPLBM/46UAsFAjbiZcKrE88DtojM9krbUyRzKkkjdAwxZvHoKX/2
UBiQQKD3Fipi8X9pznHWwwgSLQPfY1MDIpMJCt0BI0Lu2KV+A6Oz8lnWzqO+2huwzwIuTQ1xEOYN
3WQEN9rtbb1bXpBI0ynL4f4/h2rPM/CJaMiIOqiVMQjSG2NpPGRPgHt2PRf/mFgm/o/kHVtNMeWY
pHSTiG6ZF60WKxffm5RdYzLmk/vAKwtLpXES+382PAtY0KQkbWnhs+UOhmSVcdL33dbxXEtXIAkO
QI3typCIQXFzIi5Ta1Iq37CyoP90AcSW2zT5JntmRaQQ8ucN5Zc75+nVUlTBlARViP/SattnPFMI
n9RoqCOyuwbLjrBVL+GsaG9x2YzKaASqFSCEAyr8PPBdU86sGJIJvGTNtzEUKhxmU46XKe8LdTg/
LwSAqhkngQKT31Ob0e4BGeMMzW8U3/UgOohyIVlzVfe+/gylaPa4oSquhdP+ncvw64AQGdgnEQju
C9HTOHacQOkqZeaZ7JJ229btkxW0MxwZnA+eBwOXm2velP/H18WawU4czhnOad/f6U5UIWPfBSUA
vzm8+4Hx5uGbVao2uD5q/b67IYn34LXzMboftSSqkQAzlkbHlAYSnXVGw8LRj53ldetppKjpWtau
d8I974oOoWGIUV/pSvbuoKPiVFxBkEn8w6nwVGazHCTCt2BsW92tq/IK/jUwylm4008IXVSXYqkZ
4T82qytxcZhtg5Y+ufOf5TtN6yFPUuVwmMVWeaOJp3SwrjN6nh6NxX4jUPZtcacJNb0TUf/ZrLYX
JmIxvx1RsEOQnVWFYwLT63za9f+i4YKlpB3VrdYGF3p/vpU1xFkauNQaSGY3Dg/ZRzgFGhy+5Fcx
OjvmiVuFIVF1hR334sykK3hCFJBcpbO/wsHz7i3OfDbrFtF0EBhAetCKVMyR2quG8cxa4w4idZUM
JKyhZwBYSQM5j5/RlcUZ4eCrZa1o4OQRZMeupuKlclknzNfdYZz/omzZEhEMarJQPflEeMrvG0e4
ZQiv1y1jdKyEbv2lMZDeSuIoqVj6lEsmM6b9YIT5RlH/Lzx1NKtmqPkJd4e0QqmMHtun55xbKg8X
m+UmHQU5oKFa2JS9PcNyW2tpx2C0zsRCjUpbIiE6Tfw0KX3Z1WXooaArexcTOEgL6Zx0YA77GkqQ
HkxukEn6sdjAhH6yArBFGhLYrgeVZ1lmunrDeACvG9q7cv+3w+jKXHzeH2RfF4CLKX6rrUPlNhzU
j67Wweywtf9XKe22BAPtIa/F1m7Zny1NPmynAgTWJnevwbzSixDU4Oi7i3qCzVMSOAYPa78u+HXu
huh5n5t2yFl7EWWUEau2H5IDDVxT41ajYmVVF1Syiuq6yQQdtCB3a+AaEvRirS/evTDGQNak6E4+
UywovvtyTvLW+FlXaLBs/5RUaznLP/llPczg2fF0oNQHVG35jUjcBpvYztApsuaJQGL1/YU+YY0o
X7Znel3pApAlBW0MLp2TEOxm94nY6qb05ahl7wtZOHd3tMsuz5Q3VoPhYPR7XA3LgjLkYTtP4KQf
+gBl3YBWGk8ct+u04phdofXuClCEwKh10V1BI25ry/OZ2JcBBr+LlFELppxwcPRWb9gFjWui9L3/
cRt0e20mgn66z1kRJ8DOunAuxGHW0S3ctQ5LW++EzQJjfIVgZWrYUR7V8MEOSw1bcrOyVrG8EFZm
OVvFGYx2LmvEWgZ0obkfb6vdsGUZqbXNXon1I/+ddPXhPn9ygdoL6/+LM5wfGwI65d+C84L+7zTr
REFDPjxkonc8yMpvMNsOQZ19pYCfzmU5A9QUGs7rSgBk1p4zj7NOsig1tt7B8IHzfiTccy1J0bwp
LAYrVCRXuIynxKDOnA3yY4rACAfD2+Do0ohup3PLe557rUgnz8lWXpVfVCf6fCiYFFNGjRKffL4u
GQAZHLl0Dj7FlUQIvx2xgpt0gvNKIq9mTCmPZOFQ1ni1GpeBwbuGchhxGYrbX8rY7vVQTSTKFAXs
eLzomJ3WEpggS9A0leNmVP71CUDZQkxsqea5gP2B24cmnwj++RWUAYCM36FArUBhetwcausNUOfm
gyaF0kOMcuNC1j1BK1Y5Eb/koU8kMfHzTIhQQBWWzKE4rHWCHG+AIQ/38N58K+kXI8dRsyfqejer
egkMyonNhmPnqSPpzuqbF5vbds4JRlh5o1np/fNafkX/sWMRjdoNlE8I1ZJuW4Hydul0GQfMgK/e
5IIY8Eu3Nlf+/6jOvHYTN2Kd9qvt4gwF0Q549d9KZhSGZ+/H5Zc7Sy/PvHgxxUXy7uR5AYhfpHQD
kS5o4oey3I/cDdzwMgh8+1AKng8pebVUGBxpN6IEBRoV0KQbyIcpdSkvz4TnERFegP2llCnVAU9n
/0bl5oTU1KqH2BiC6w9Yjwl+yejA92UWAqFxW1+8RV9BQc/J8vgzkwhjhHvsXfnjLmzu9HLF4l7U
nYa4xlUDoggd5eErNTqmA4o0GewTTWiDaCOAvAvHT14deDcJPf5xTu7Yi7vK4x21mvTmOHT00bAU
g3AnvNSf8mh0qSs3Dv5YAiFSyXUSSkSqxJG+x7mciDqJWTkpgwHINbXBdghMlZOdvEGVPGf0McEf
Cbyqchwsd0BsHyp1g2Gm0fQ26ejzLZSKj4wn1768AmpkUhb2EEeyRk97tDAyN3/8fWaYeb5giFcB
JRGfysqgdI/0W4wRuF+BNb3AsyeI4wn+bhtueF0G2zb5jTZCOvkYdytF2YbAI22+IR41xNvGPsRm
b/eMpJv9HoG/3VNiuaWa/7CesrD0akdy1bWpRJCcFxSW6J1kTfDQ9fqWRfyR4B8jQMiQAeY9Wfzh
LXxdVQyBNoq/GMLu3jJtugoE47O590adShUuwF5hoLqCpIul4IdYiWKqbkhn5NBvwVJNcyJlGF3O
1fHocIbb80vb+B79kyUW5acZc6faYoy6I1gJlcMvhFtOG2nV0kWmp0sa90zIuQnj7l38fBT2uzaY
DKeeK/fQafcbBAoygUSUV43M4jJ4V7SJkyUX9EtWK0TgNmVLMqamuDwABBTPob/MJ27FH/s7xcap
OFMBWz8q0QPiX39prdjazCrTAe0vEKc78efvm4InL8vMPo6mIXz/qIS0E9MKZsOCps18/tKWugc1
kvcD6PPS6HEwBRq9NaP2KPBbbb6u98TpCK15mStF3MSNu7iDzRvji6hY+NByM+Y/xzhw+Om8Frmk
eukkSypUqVKcCdG+rRC33BPSlsz1BnyJXLoe9sWhYuL+bakYAu2+HnOpn3U4perciX37PyCQDgs3
J/c3SHnQWia1TGyqBAPvET3vk2lldwTXlv1uw5+9g+S/v2H6RaHkAsbRO0fWyRbgmMbB5/gWaiLs
8ZXYIRnGGm9DbtXi1oZq6dhUBKgTCja+ZkzZTvbDe1Ppzg+qAH1ESNwLeQeOmEbY3rHMdBsZc/mj
vSxSUDALxf/LEjkjeaMIoSth/r9Rbdr2M12yZwxGuvZHucjRMbNsXu9KMnTunYnx8Wf068mLjNPM
rmLzJ9xGQd9iM/Se7MuWa1oWRA4yV5iDAPVBYgtSr5QJS/baYJcCsgb0MdQrUofF1I19/oqFPmAR
4xCm53VF5JF5G2grwTzw1YRu/H2yGnCDBEc+TNUYk2xIrPOtrTc/NrAbip70HN43N5Bo4Be0JZXV
JtSZJ6aou0jEpBiYtjTx0Hw8ynarSKNIfBMbYpJFm9u3ozfFELLpOyJJxKpyePdtVDfwMKvv1sCy
CrCauZXw3PPLlfU9uGUqbbHFc8bGcDq037tNXxfck79RscXE9QWZudYOcutni+MJw5FbUUpxdqUD
XKF2YCtH2K6xH14g158ot5lvp0jrHyZ1BLMrzHbG0ZXxoa0vbFTbHDaWy9xXP+5ttf4+7btKTD3S
WcsdHCp22SUTTX2CF6wu7aFN0ccccS6ewoVQcC0P4hJn4TK/z5oITPcU0PIn9SDqtS3+liyU4Hcu
jeGZo2GC37ZCe8klGaVxRkceTlFxm+Wp3+ckJNdFMGzZI33Uhqf/Ds+MFH8nJQMdrZPoejjcZO96
1g6eIHlMKYFLOPLht/SPIj3fwnTGAo3DzzBzdHuUvOrCRC5ibQPlIoTxaivthDTZUW4MgQT+/qOw
oQwFPOlF3YRU6N1e13LWzXROWcSmb9hmZh1gkV50swLvQltBOw8g0dF7QCJ8umVRzRUQmJ/qMl4n
IEpL3s59alkC7FY2Vd8ISBmniYgfyEO8HMmy68/h/uzRxvI9AZoyrcl87YIwADRHAZ6IAxbkreKi
TMJafFiubtV+bGqA8q3Ifb+orD3mrRgKe5S4ifnzP8fMs8pYrplMWI9opSWpvdd1tSUY9CA066oh
2W8ehqeg5Y3iXNwuscgHw3tTn4fKNGnzgKuM2r+RoLUmNXq46b4+voIN7rbMiuLQ85sfu3EeMPWq
zpHFSm9PRCxKUJcCxubTyaTl6RKx8ShHE2aUYbW+tEoIKHH0lTjpKY98+wtMngAiCD033GDTE4PU
t2L3Fc2xHZEU1MpWkd7L2kRlwJJvKoUQRR5jTR6VC87W6Cw0/Vh0JzVFnikSIZE3uMpRAoUJhs4b
4+cKmIp/8Ue0ERMkV5pcRnzHt68YkkFf1ilTU5Wr7u3N7IMq4jwgo8EnavnI5SXUaeyyEuvsnuy0
IOP8aBW4OBiLNBmIZL47sXdxwFgd3yuhmjne8qviwVm7/lJamQiPGkUxdjyMNBrnc0cmL+WvIV34
/9SPp1DwwiAnSa+x1Y9q5erpivda7ARPwcuGeNSeba4v12lGYZsymcw8lwB8zZA3uAIBM1FuTUe0
qFDLKKRwtmKuStm+TymmmqZFKiTGD05aF06wHDTBHQIFPOLa9nwYzCFMoQ1WCRrUJ/Qoi5wE98Ul
SckHJSBWb+8C9RSvbeL8N49hifkp0slaPmAGQaj0DCvYXx/jrxyjoG02ClhQNheTKhVViMbBDjrj
oERlTyR6IQabb5Fo1QPBaYLmwNHGnBqUoG2ZOlqMN95NvraNrliqxDL8G+m7tqnb42w7onQs7+qM
j1ZVYbKxM20T4eBTm5UxizhYReUU8bd0ZLy12ZUibzChqKfdtg5pDc+cruWmAV3PYEkshr5eXo6r
+v5jV+XBLANdh8nWc02AAJBgZ8Bz20ptTZJd/X58U5gj6XMR2OGMi5Sl+muswl3df7ikdB1PYkQh
uoIUij4fmmtjBC+KTj48Pz7s/0tyQ/xhvSKBBE0iXf+b0XYleGj9FhoBR9hStU1fZoSuh7O+PFIH
o9vkMQOvkIx2Y8JCc+Zr271A5TdbLyBH6Js3StN3EyyZ9WGjIuFPoY16Om90ZZ9evtk8mmEI+Jkq
iNTTre7z67DVgdexPskMIplKxctGwU3FdQM3CUzpjcxo1lYW2T3moDt+2swNGaXFkP2ZYu8qEKrt
a+R2O8Fw9WCITau/B6zpf7OdbE8nA+HGMBQ1YvntYctbfyZse1SbDPAoGQj6Px/5dbotcGZXp2vn
96uReJYmbcawMTV6fAND7gpF3uEeMq9srJdW7a+4JeKlS8mqs9HjJLFb/A1Hpm8AK8ogklpLs5ix
SbkJw+NSNk6JGY79Vqofp5e+7e37NKPT70A4f6EyBpH5Rqu5X/REUpij9DKhL5Y7pigQsHgP84ty
SfC7HxP3VrKYedX5e0mVz8q6BdpxlfebF1mtFNObO6h57vxnOZ2KWMYfsRVnFfMoZ8GHuU5wpBek
xR845hHWV9wShttXrJMemFpk8T641/l97IWp4a3C+aN9gOK7urT8xEgBn00stqEcs5SUb8KFsZLV
8O4aCEN2UVZtaxBImjsN4lYdge5YXFRY2eq0+9m7LktO+Hqk2a5J+aK21B7TpFMq9kBKCDNuFIUp
UcUM6sJ6iorLQnLMSo5zE4mfhZRDDeykia2VlymhL7/UmNSRlWAMzd3tYiOjj9UyjB/ljuKbdpry
X4xect2Gy5D0ovI6UHlCNIgOe9UHdkLUpH64oMxyd/qMTSn38YCatWcteTRrEaDOeruC8LDbjNrb
tFEDvlAYkmLGRrpyDBZE6bhyJFhwEEVbY1scH0JKxn+k8WfBiZk9YLolm9CjojnShp29YdfaRGlY
mKDsuMiW/HFuflUCvm/JSNrwyHBwDp/S9VURI92u/A0VUjtrjXsWs1lRsk4m4rzxGl2mwxirkyo8
MtSA53chqOuxZKKPbNqHyTAoUVCWw91O4jH9nmGe5/uV74JDM+iOaqvPRXCIacbYUIWbKmiOBULb
E+aWiS8eBuvTj8donTA3QTRZ9IgG9Bkucowf2/rz/oyhJyGe255KQd8ct9WLdk5ijdfqQerfjphw
UMjHtm3RorymvGKgiKkpGhYopQqtlSPVAEJCGH5/EIU9xClpQ2zZcUiXBU+SbugAMHY/p1bqVQp+
VIZgxPEm/+7qGp/FiVnEyy/sIDoxTP46V+++RXNqGkBXtDtGwNW8TrOjp3MqdYEOFBg6NUmjCTLk
6lq+tylXu97kIsnhKZSH4yUePvOm1nzNfkZlblc8XF0DkohrDOr1wdnwF/w3AC3u4M4T2XMAsQHj
CUlNibrDGIS4IF0nHTw0yM7o0sOX2ovRRVyft64dY1C77nDDjoSId/zjk9jILJwiSEctKFDIv0Y8
9xABuZyhedJP261FkzpJ7GZbgx0BhnxhQa+6lks7/hy+pUj4Eg/SmN1/tDEjOscE4WP/K0ryU/sH
dN7DctzUpbsq5zAeaMRKUKD7wjZwIy/30bDRi7n134EJfIvGvvKcHO79axPp4Oeb3S3E/6H/+2Qz
oS2DHuoH+Eg4v2FvEdX9dGeEzqt/ZzBKCnd/7jyblZkbrasRI7YTW1QV5OI8QXf2/JGSxshPGUoY
yBAfJvbS83BUmynXmlOJgPPq9C9CwhNHnaM3iJzkhyRu19bPsRqtxcYt/8w2tBhDaHBxTdabUBHM
nHBcZ0gOZanWHluSWZcO2Jm//bpfULZRh+Qtpx8FUfMrionddPx31foxN+69UfgJgJbiWcc6vMI7
wDVmV45jJixrn3adzehym54CTcbYNlETw16Hww+KilNbZ7UX90l+7nCR0f9lJ6khOLsX5Zz44UKn
Kg3lPpfoBDMuvBx7eZOnYQCkePFQ24hRh6TAcWLgsvgVlli36e8Xx34mL2hRhGLQ1UyrrbAq0zzB
ralvKykEUnfIX2Lw+CCFF46Vg0EilVETbg6RLZiXc4nq4X3hFKkmef0MjiR/Px2LkgES4N3QfXuf
GTR1zmb+RxT+YVSblphyh9pUIpoGgcwomMiDp5Z6AI9gIkPWwYib/eoigQ67AcVcEzae+p5oYR9p
qEbyLkwKDJP/eq8VuWinaE5P5MiyVG5n5sGnWooNqZuHHiYGi3/JNiFwt9MMY0wq9MFCSun9Oith
xcuohSoH2hNTrVqH4xOwaQbRJdTu745K01yj86iNnTHumEwnNtL9O9JP1t9XuTyPXca5ITPT8u7H
gh4pkau4Z52P9UxkHEIf9fQU3gQyIRuakEKXx+6S1ujGaNwnj9km5JIpr10Qb019j2o96bVDwseY
i3SxOzPMeq7ucD5BD2MyX+PjuB/2hoM/68wasqz1seAp1CBw90lirIv58dSOW8HO12NDCgkzMnO+
bWRqhrN0ePNcO/0epwR5H5VSFvoXkZialY8AxBg/Gd7iBuVYqtGE9EQUcy5VS2g/1nf1FM3ohdsA
1aENBjbP2GRSJiB7L9OFZdkP3cypyTn4qp/tsDjeDJmaRHtD4Gu+LjA3Fs8WEijdczHzkeemV06s
FjT4un01EEiQXcNbANt0+J4xmw33PTZr3mZUROW/QZrIVsifcoCcr5NTJ8ej12QprBCzLykZalTx
zLJn5PFFHsAoNZ2Fsz1VBKEiaumketo64LscE7JLFIMs9NAt9Zd7NKbZrxYZj197PaSVVskMnnKw
QkN13exORxsBsMkujP0ZOGcOB23zCnZhtwfEY5gbXELZki9c4J7+uvGV360Dc89W0zHmaEMY1dXX
YNoOSSSA3ST6m9Ul/cKu5ACRj6z3Qdfbmr61ksm1YlXrKel5TnJiwQvegn+7PnKfYeUUOUzLoxst
T0hiYuuavYBSlbQ4+NWL6o8IwNMR2w3AwgwcxZmmSgj89TafH4dx3cfXV85nJDfz8xtagVZQmwkI
DnqN3coPTulhYckg2i+bGaysgE39KcsPWBLzhowLG9Ua6Iy1qBDHgJx5wzQIzPlrfsQapFjOaTSA
fLnOWwHOH0ECwo31v3iRuvS6RCmK+BUbpyjhDBzA6lPokjnGYFrSPtmf6Ug7V7il3qQcrcSH3nWW
R46mvz2iloSKLK1Zu7mDzjX60lP30hRI1ea0wlyBioD/dxtcKzFJ/Q4U9U8G+/mLJJqVuSm0pA/f
rg2z05bo3trRaPjJtr8LViNuof5a+V6r+4A2An/N5tLilQ3rNtSJv57UQYiphtgDeeeLFBdGgPRn
rKgL5T9hjmgumSq6oSkWSGcvO+Fq48Z0mLS0q74YxMRPmEHT1fV0rgEyBLM1/CSaerMmg+5x+KxX
q3HfICP4sE3CaYs+/HfzXhnEm6wIF5L9wefE9CzQnnqga6WE75FDey0vv+vdwRbZzU9uv29L2wWB
aaxJDd5yWdTgxrtmsOBXshICm5DtrEI3/+Fc6FxRdQdPLVt/E5BguXxGwJxalnHSB94M4TyykhJP
eNRbumgfln34cxllG+SDKBa7tGMKyzcNuoG5vYAfsuGSKd+VlUethifn9P95a/syWDX792dgciU6
L1LI9v01+1IPe4EQmG+p411RlTY7TIDgX9qbYcQqlrL3G1df82ZFfc0PwL3P9Mam4mLR1O0TyXzj
zWHVX8rVDuAP/n5iwhAUpeMuvlmwz5q3u3Z+j9rDmWNYJWGhmGsIJsrrEnQoR/GGKmlL5CMqejrG
svEiYr6YYgx0wIRs67kZL8f02OLwgCG9u3uLaq4hulkTU8sdqVq55kKAGfJRKME7EsEPLOnufOnW
yI6o5EBKH8q0sMKagtoKQlBt0frtm2ERwxrlkrC4/3YxZG8WZ9pGlvJo1fqQBMUg++Y2vehOf+pr
HSRSZgifY/3ikW8rbKOtBSLds0saKqKbeIHvo9ZBC5ecGhkDta2VdRAvtXiMRdt350o1syYwqXKa
XJGBLxHPX/vwmuRkALAWhfufN+/G28/aTEPWVVL1PhEKDBIAswOeXFgXTCa8R5puAhU2+cr4fd4Z
CweD1LqMy+Yzoc0y0f1JUez279EmfK2+kiFh2FCpNF9mztXGm0zZmPvx45uANUWEwsYUblXUUDNo
OnyHuuoFp5A0HsQxsVad9+cfkeM+MKeXfvKYe2X6QBGuGA2YpZEZW+Xf1Km5tP3JCfy3uqSwjvhg
i0QwbJNq1CTt3OYFRgqMdt59R4F8waBH96p73IpjrYOgAqp3qauX72Leh3/0xjZ7inE/xFLqoW0M
3lhT3x1Qq7oIZXmzxDu9/QkF24ayGfRVn1yDPZANgHuOWLJGr8nE39jJj16FICvWBxHdrA1mM17J
/j88MDn4BdqEZFuHpI8P+WcGeVEjnpKjth/4md0vm3+K2sFZB4BrvhTSI+bkuhCCX8mW0LYqvgAb
h7rtavFXvh8STw+7bT/W6h4K3Nx9KLTCDk87HfBEcjAAlGKNvReRUlWdqXa8VaFvFvM1tc+wzAVc
YC4G1Sjqnk0eFBfgEMsFu64SVc0VVNi1yng1D4m94dMqZ8oSXwETmHGCOJ58Zkutxa4MFt2w4I2j
Ns7caHM2q0pYH2ic+k5SqA/llSlG9UOddebSpcsMvj2aMp5+EMNPj++Maf1APvTHKiXtCXUya1Nq
JtbbypMV723nuqHCuw3sMwE/FpIb2zX+zVbDTUxlZgLO+27Sq0VuUm7MbNUNJI7HvcC8AVo/EORT
NzCAnnmRCqoHUp2RbRsHetRjycp/lOejBBZe8KG7867F9kdnmP6CW8J31qKlb7PXMoeD3RQuH+OR
Iv24YwL1wdBs5M55rhRZAmuB2LRSwyPcLGzfs3l5ycEzFGmejnimwg+hze7ftUz9yyQRrdDwoYHu
ucuYcNtf0FUOF8O3m+BbM8xrP9Afwqx3Qc27kmI8LggJxEq5DT+6tMJ1N8TvKQHdLr+BHWIHTBuO
ZoUbKhtiFOKQ+yh/9P3KCv1vIdGhXf9cYk/8ek5qJTr6PAaerhHvQP0mnzaX6nvUvWeDfD9nlqAq
3p93+rwbUtE5KsTa8LCqtK0BhvYS60aUHHmdrszGNUQJFXHSZXpDsBt4jMN5YyQpGNRB88Znmjpu
v/Ija6oXxSzgtcQbtFeml0L21CzWB7fttLp5GCsesKUAq/HAZZBlOl93S5ImRLiNOlMerR1tUgv+
ZzmrGT2cp2Q5VcRzgNvgEwS0yBS/uRFvO4l6CvGUerNZ9gl+jOpmwtFk4N8UmvnnJC1JO9IKMUb/
YC1sL5rMOct3xqjOsXL/CJ01GhqTk5+8EHymcYIz0yGqLL1PVKo86/I8jGwxm08aPh7ZdyWxFjYT
7lIvNT08yEko3K33BIf7JiZpEKURlUuHVPW0rlUu26GWne/PFtXUFIZSar0Hfp8e19JHeVjcbM6L
fBgBnndi66a4ZPLZjjkkn1pBh3HfozyqhDsqiaNXzeVMl7q2xG/y3yMdadCUlV80u/DN2Eeu+Xpm
YN7Op+opsCA52CdSSR7kw2noCdRZRlSDMkexKjAdEH+Nl4URIOCcUK/n7WbWMg+e9EvRAz9pDivI
vay1TJKE4wbq3P8cfEs2I5C3GhvkC+sO521X2kxQ/SX4hADq8RDPGEy8t72bmlvXX18JPAs47ClL
jIWZR9CwpZLnZ9tGeP52se9lYSGsiFH0JqE26HsyFEmfiVb1G+1TnAiyMFjK+QsVlQUUE6aFg16V
KFMbdy+LK1tzKFi9IllWrxm5jRJjEf294uSzd/zCjaalvMCnTEQhLErYO2gaO1qjM/VNfGQcRE5Z
c2CtcMy//hr1WpKdWEjsrFGGsX9uyjovvV8HPD16ofEdN9rkITDOdG584tfylHhjNzMo0JJoFmgY
Z6jyym6ez6Yxc2z6rToCM2hMn5kUsgYBgA/ZEADIw8OfQnGsVnWvl2QIj+BvRjdRs8Xy6slC019x
TzUhjgtJaLH/uUgmts9kkuzg5wP5hHaPMXEGgZ1DE/n2aC7e0zFMNz38b1MoaSdrTsuEMUtgUqBW
JM8tgcc4xuXCylC18PSxBY1BuAiHMAgzR/L89luvT0o5Z/J85MVmAwKyAeU+y9W5YpBBA7rlHs4w
6DYswP4R/6t6PwwLB67Aqiu6yiGWYJJBUVVXo+riP0EFD2DC1dgm5MZUz+JN2Dcviot8/WBEjYC2
AeAWJpUwi7i/FicQf+l5PcJAt7mDXBD35bFMahhq1/LozEcv9fx6KmmraN/IqHMag2sPKGMjIT9H
X9XwH7s6BSHRNCqkTCnvo6KtEeqo3T1XW2yd6/pm1igy/+k4FR77bf4kRo2DqtSF2cbQWTWV2uU/
8EtyhXDflZc9M1twZBsxUs/JSv4C7Oa6TxPihLzedEH3sUZDxgvopg7o5sKAMITwJkrESmPaqeLm
lRrCouDgtrGcrISp0swhuw1rfQL2lFRntX7xaAsUaRh3EcaoXMUBJmepSYvJ8U8C2vW9Mi14qTfQ
+DzHQOZv7YiIECqfg3K2ryiU97VeLwqGdbWWIOxPJU0+6qYS2OmMU3bQiZoU0mOV3NyEoQC0YWc0
z92eFhbd8SpiPUrQJK8jYCEPkJgPJwj08uv68LILE9dE15d4SkMPPdF1i+2toldY30IMDuZpGdrY
+cTUkGP2ylivVz8CuCS/1d9w9o4bb48E+sLSj2jX9K5NkdDABFcFIJV5IlC6j5TOMAH3a+BhIde4
lXRqhdwvlixlJbN1NPE0VDXDSl3mThozNL3a1gqMGNY9ABuU74j28E/8XmbM+OwvbOqNe6dp7gRr
gNZlMQIEWQBEQ//vZN2DhSx6VqoZqwAB/AZ/p8tHkXnVUa81SZQ3UshAPz4lJjOVzqiFH8suIUYz
3UT1ArRP/9wok66pkvAWUrYde0WGzTo/sLuFUNEf0B3XuKRpkjzicBzRpfKFvdcT+QaL5Ht7bEJ9
GXiPC3CtwQb967b4RQY7TBeUQKnRJJvDbYBTd1ahCiwZD97+bimxxL5rbn70Jp88ueu1UvUJ2ieO
7u5OwW+U9zEAyhik2qtwuVJ2Qur64tvvgvwTHpkAb5c0psT6ea9h9jchJuSZS2CJ1St2eBjbFSKD
qhbRBDj4l1uxb6UZSh08p+y7vH8bFV0ddkZpqPPCBbUpFT63BGbTYw1k2Ey/BwZ5mmjhyIUbpV4h
X+wSUqSSBdL/Q42aXtZQhTdSdovb4bZEh0LJXvwxjVpegSAbEoZz/27G2LechZ9KWoqCckeaxF9o
3qDtqNwp7xdj2L5lB0o6b7YxNhAdv+dCvDrJVqM7szPlWQCJIQ4CLcmBPIpwQP5CdgICutskDIsX
HB8wmYAwxaVvoQIEgEMXMQPd2Exp5UZFLxhQG3XPHlehra0ToGWC60ixtsRRb/xzAGwa6HUbQ7ar
OYy5B7IGkVOMEhTrcdll2OPjI2Chqd4ehYaV2iqpWvCxOAQJ0lge2CfUzT8ghkvcWKtXDBbPpU6/
BwFXWRFm+l0z7Y9mYilQaHrXNFdnxkgR9CgzATEtmvls6hRiLoKDBiOTFnoAagXjLJ3b4e3B+krC
LPNxjohK15NgewyLl6lJbP6T3+BD5OOHTcEy2PA7ZHYXloua4isQ3XlInFO4oAIXGifKIidNf0z6
T5RlO/e0zqF1x144HUG/WemorRptHrgzkChXfNvy/zDpyTnXsz4GcCbNBYRHA9MwQPmP4e6WVRXd
vNpWqWD6TSTqyCQVaYDgFszzuaNk7qOYqN9Vk552Sq/EZyStl1EiD73RkpzwXIQNSyUl4PXKr1fa
ihagjqq4dYJLRYzeUl/7CcVTTrTugBYW5tjTAKS+VBVCKSq1VZddRH1yLUDrEst4T5v8XSExKhUO
H+T2tS/C2Q+v7YApz0ZUeGNWxsYX27dspzp/QiiSxWdJ5Ar3ArVjaIvCCmdHtkYDRUI1mSyy3XIh
BltFZUd9v+/mh8HynAWa6WvyTI7jp2h1WtstoWbUf7cirnH6+/AsQ4qqweT1NmmzVoIGwLbDKVcq
1svNh1rwLUxcV42qYQ1tjgOv3YKUFQnNZy+u3TVMnbXU7g7S9OVFIaEfP+ncSWsuxTraTXhmGQj2
Lgr9lBW+xtVIopSp6IdguV5E+7ccLv32TK9cmLpeLJeqtgTdZazCRIirRNbhb2a3f0GtkRQyL2cs
fMT903yzTp9hXo1XXW/zScV5NygkQk8QaG6Y1Vzpp4lraZBmPZ+oeTyF4xNtDdFmC0FOahBraaBB
Ls5NFYZbpHZ8fXhRX+VpkfCseKXd21jPEkoNxw0Xe8C0uzCAkPjtjjLxwVKxE2+mMyRAyPe/jL/z
SCvSgbC8LyJ2fOPGmG1RigHeDBnug8Q5KguQXefo5hiiHmSiTlRa3ewDEV1wfLuRHWvS8PRnRVw/
j8h//ocGGQa2UyGElUK72f6xr8zThhfYtWXi/+KnD0Yhp5BMSyto25xckcLXI1l2QtFwJx9bmJ/E
SaMu1+c5LP6WSPvBUZbF8PuHAh8qBsWFgeKsAgG9sN+/Dtzw8CgjwHd5ypElbfpjnDNee+4Ob4Va
ZR8Ip2SPYIXl/5N0IC2tcHYD23lhdCDbfAGM7ZkHFKJRpDvn4xv799bZm6b5kgXBq68PjLelUhB/
8naiul3vw8CkXJDdWS5EhjU2eXOOD5n1KO/qjlopNGQ4mJKf8BW8I7/InnZ12Y7lAbyb+Zo/dpl5
NciHOXy5OONaInOKfOJo/vuRxHUXheHlCnp7NaZrbgsnLKYNpYVHXQC+H4MEbmuc77VWTGzn/cAD
MUNKkZkVoBsymgHr8Prwe9QhJBrCIvXhRrJ1zhx0l4wujX86VEaXbCtkOEUAX+DRtcHSpt4gkbX9
YQvnIMk5rgQ2Vs7i543crPilfe8n4gqMc6ZJX5Yt7A4tsw1z8+2QV3FfZp201gFGXFWsaJR9+H6Y
iepARkhH2wRdhGy5Y0D9Mpp8XzUEv6usc59IVagmaOYgw+4DWe+8tT+ME6jqUlJ624Ljeu4dLUVW
/0NjoARr8YQckQQWvSAG4Yo0nAOGbqUHrSZaPZSXkUcMCGmT+V2mV6v4Disx6pYmFUnhfulWfASC
zgm4DUh8lwwaKii8Vf2E++xe6s2TK5kMUpg3PNLwdWxhF0SKc2ZzjupEmAzkNDk5Yj4poS2STYCM
fcZUpfKDhMH1TyEynBJ62TbDhIDvYjA5APZOq3Swi9j7NkYsz1lWaG7z6RtHUrjFgWl4YexskFjB
j9r1SwCEVZw2IeX/3LTY51wkSC1zU/AqrRnfZL64I8MykYa4S2/L+SPGfKdDFhqRQ1fKFCqKy+4O
31oro1m8845s0k6ma+VItflrnicQq4kBKylc3mXhTwIUAgXKBU4ewFQWPm6911qmArU3itbks+JP
ykUhV6viSqzo1KlnUdc+FUU83Vfa6lmsolg4UxWFcaHK06YOqwY0UUL2iLHl8vxtS+G7iQhYxBrV
QhniG9VQuMM1eeV05TEGktgzPL9E4Vm6Uo0OQGXLydfY+tzqHp2e5n4p75FddX16dVgcaAtPA6rk
ZuO4jMsDu4XcQFT/my4VVBxn2UdyRKoeiTIqazyk39sfWI3NBtnGOfiFkv5fIm8CLnFBxF2/BHVh
8FcgwRVC+DD0F5k4Gv529SrtLWJSOXXS+8mwSElfIzyDVWnAaUeYI9RD5sVyVdb+FBNc7ptXK8Af
xDS1yjfrbSki75sTS9X+vePm6th4FTxhr9Ay5T17MKnQZiYbNn7ahRf+n2LTGrliEMmMDiRBKAhH
pen3ak/iVhe/Hjka+8mgeoolcAEJ93vS6Chc6zch2u4L/0PS/Ut1pV3FhXgxSQLTR98qFClAgbUd
VNfxu8RO1KULKzuEg2ltqXNNvx3eOsjwNzilGYssV89IDuCXDSZ83rzrLGk2yyJCNHnES50V1xIJ
By/L88TwJmTZ8M2xJN84IWUPcq0stng55I4PX0Zf94fsTw4z2eYCQBwmM1lNKdA2IAshkluNHbSb
cvtc0zX+SLqk15tvIkiqfa8YhMR0sXNFbJKzacCDlU3feWPmogi0e8q8RcuYx5sDkzdVmY7afdAH
0xJS/vnXbfEnUKHF3uX+JfCDrgg+eY8yNQ+6CYTKskLkz1qFcWwfhUrBaX0mvttxX6OotBE9wWxw
rfVRfvba4s+9l2v0+xQC9nroWn7xvuf1DKj/tc48FoC9QYRBKFiVE19pyp+avrksRe9/p0xBqoqm
8pLeBAnhmoKLlJSJZKRL24G9n/vcwdITfPlZu+bUATUjPRpVlTq8fCtEtCIjO+VrA5+AF2a/8EPP
p6nCBYynClek4pIVAybfVdBvVKr+M0V14QvnUYveO8O7Bbu5zQfINrR82fpXxQPhS3ZOH2AT02cT
3iByhB7uYEerJP8kBElqOIffe5kOXkjwVtXk1dWfT1rYgZU/LqFOMCmTtPkdwdjxbw3XMpXbaJCE
KFiL3HrJT0Fvh2IjiDTAhU/EvIyu7ElyZbAbMMrDB3jM8evjIxGhBL6oy/EmtdUcUzmaWsoOUZpS
j8FjvtqbD7K9I1QIVKdQOTxNcvyuqRRZncEqcaVNuODMNKJD5EviBuZQOGO+ZM/MuTArVhe1ZSag
gKg4hgPgZkI1IPzyNbgnVeYiZlBiXnJHND97tZenNVJ/hKlaShidd7Dzj4qEGN/VWL/81L+2J2hj
H2lqL4WH3M/MA9usRbs+ppsjcArxvpC2BqzYlMSe+mMXoXFrft6ls0CGDL8jo4bCHyWqrgV91e5x
rE3XXOk4lZ57vGjF2Cotzw4sqluGThLYdSQhXc9rDMpCIHKsqAPw4iOvhyx/CxbXAoRxABb90nQs
5nFKulAPvUeqDVrezFiEgtJkkM38wvAcY3TSFfo/LJfscHg3Z9rPMKhOPBkcymELVBgYAuIuqSpR
cMcpaBu2VpJOAADKZW139szHGvb9d4pwxdlHF8VHPq6SsF9OO2khc2ZxpyrRJw7+unpNrLPRE/vk
TxUZAGpkQgEs5OwpIVjVjlo1662ik2d5ctCl9O+aYtH0Y1XrZlrO9OtJmtVbXPEiJ+d2bQxH3Hky
2KDBpCjDnUV9Dj36H0aguUKOSXOCcfc9QcV0l7JVNS5p41PH3c7PvT4mr6DYGiBkQEr9v6vIOPbc
exNjr8wIeDwko+GGgcTSGoKEbmScmkv94X84fq9IdtC+wz7sNukP1AoAADejHrby/OJc3u5jc1Gu
P4UdaOhHZufgk3J+pOAzQtfkg3WovXrQ0efclZIvbr6u/VpvYzkDW2Ojzbj+1Nrsl6nHh9BZsMiO
jsLTa6x2stPi8vDOBiqVBZvIt5DJeGpD/loUJeS5Cn5LQz4JnP7uhavKYH0VfeWNfGBowaQk5fBh
0HHzbdwKErqE2SqF9g6F2yqNML0SEMoNGJYEC1kHyShkE7lqSy3xHOzDlm8dAQfjp06oWOBysZGt
ly+HrelLvTHoVUq90jUS3HWVyLySiuHIUyFlhSzjn5CODD+X401h2Ea1Oom6O/qoy/3Kkwr9gEIg
vuXeeTY+5EH0B6otNCPeM+/Bt5wEvM71vbOwudrN7HkrD/LdJblhWJJXMEIzOJq4TDY8WbMQ+2dv
sOjsRKot4GBPJId+nLPa/kQujmdvpsYt2ulL4DrReH16PyZG1DgE8uCRfe6zyJiksONoNO4f6fFR
E+X3y77sv9vYQiDIBuFAQdlywLjJjOO+1aiKlnBmzf3sF2Rt/IxTb7U3AULhB26J3MnA2Tl0jauN
8IKznJUqgDmo17ltDxPz06pg/5fdEKRSU+oMud+eWvp91KcE4D2ZjOiIuVW10oz8kmLPLJXocEPx
uKJq+Y3SrmecBOfL328x3xB77Wxu4/PxTagCa129lcdhcyoSZXzAB3sldDqhYVP7/54fZfZfhxv/
ijncXEyCPPjkPfMruYliUJXe/1DyddU7SebCAihD5KW+Dz4FZccsjtzWK1fsOsZiQfgS6U9IPKCm
eFGgWYOfj5Lu3kCBNpkMTzX8icvwFuChHs+V8oEHEmXG1BmIe8kAIiCz/8AqocZ3zbKsKorBZRQn
9LS3FGimPBoWJYJl26oDotuDYMNBnDYtzwJntGv842OaHDETMtza/GuC5atY4qRynV1TV/ny5+Ly
DAfu9p4OSLkUM0gD4OVJ76QSvKIXP/ArUpc4E+6Z1Mh6BonvLqZY338YnAez/Avg2i+7KiJMIKwP
CjlkJZumF//bUerO4kOdMx0PIVKGoIQIIvDbLfCCN/MmuDrX04UtudPfeiFAQSJmJZmMD39DAtBA
EqITDVgky1EsNjpEdJTK/lI6pQ7rtHdfpTLGGpNBaeR07cqoSBTJC3WrpAhFGWZSxVIicxeQTRvP
whXdXaI+fShd3f/h/pA+AEKA/xaIyLbbnQki74oL6XqLDxlVMSKcjmEKZJ7naIKr6JHzPNSvoOEU
+Nv0KJonj7RQ48O6Fvc5whGsGCAP5sOUPDKgYp6P8lkUxiwwlWfwwkPL16JxSHbSvGo55wLXyBff
1Jg0weQVuQodpT2llGLqISUUktdrayp0d0ow9lcmelJKdAepOaNNNV9getbPZgVv/Re5VvzSyrWc
joGc5rGmg/U1lzg3MtE5ZH3Iphy4BtKDDwDOlNgb1Zwsg2QtSN+JlE+i/WsyjuDq11CforYBdtxw
EJ0Do7lwpSBoVoFQIF5Y50VtUmicxX2egqZByI1SSzLKL60YLkTgNriABbL7pvjKjO06cS/nP4aa
YTlpMLjfOXZJWRXpJjEFsSfKiyOWIfp1axE9sTkgwETUjCMIZzgVLBvW3P3Iqolg4SCWfZiHLjwq
dkC3H2pD8xlH+3C/BBOrwRK386cEqILmegJv1m/0aVE6/n66WLJy/xTh2Ul52yMc0ZPRcYij+uzH
oFObTDBHx8SBEP4APi6szgUZtcS/xV+sn0zfZkKpx2+t3okjBW4h5JDvlns6RRsOsGXf7lDrkZgB
jEzm+sVe/FWIaFkGPCzdX7HXWKne8oJV26+Ijzo57R7d2Z12uAsl0rxO4n4PyKz/2qBMYDmO/6lz
w9/TCc+4Z4DPFO/SWeXhvOXONDjspw+kKAZcE8nUkK3Gdfe9HH9SolzkljeVJPYiSCX5BqZSOYq5
nyf2ooqpwCP65SPwhCff8vc9lZyxiARSgRf7+4tg2337NMEKdqz8TXG5jkogrAfNUK4GV2Uv2iP+
CMRtvTTrGhyqryk/otZBAGf1jkXD9G9fHoCNGoR/P8hwVnTnURMnPXza0+Q7EZmPj/cS+FCS7jEF
WDM+FnuC7EsnyBC+EfuKdi9bj+lfxfqwaG4FvwAvlf30nHxFseLFPdDVAhoZrH03V6nreS5+e1xL
dobhaEKfKA9No/bX3S9NiiAZnbEyLc6jEwNaln+q10/+mnnjCwPFRfjYKlkqxFc3l0r1cjlxsJHt
mTzyKnypG56eKck9Y1ranxScpx8xWI+jDOsVwbrzSXD+Bqe2EskOL5sfYSatH0ap1bxCAvv6GtZc
HVR5K5rwvcybn5ArDWBqJaQULwcljfsPhCCTsUiLvyzBq2uAFohZK3wjE8+73PVMVtdL82l0CLi8
pTGVicQl3eN1ZZJHhThO/NjVWD+sPpYzlUpGlDdr+R3K/ojSLpXhqf2S/WtvUiwIfHjC/OvWCaaX
bkdSA4k2GLu6S+2sAtLCit3yIgnP3Gu8bQWbum9L/l1Gq7hTNp9dJOZyW7ns6SNYToXc2WD514Li
tH4syZiQZHsdvLhUiXBPXqBZUaNJW2W2Capbu6oMczUTYkArgn2NfEGaTFgjTbPYfcnVEL6qXPaR
TpEcuj9VW6sbKodpb8YdE8xFmBeCeR5PDpsl0c12Axtjln81BZHxVyPtVwTuBF7bLn17Ng6P3dFa
0ynfcsO5+rSM6N98+NxnjDipke2gSnw65dd5cLYZhycbF0fdW8VmLMY0IMkpinyUuEUrzjq5USuh
Mmbi8GJA1SgwC2wFY9e/PWYfPMhMVl3rTHpU9hV5baaglyr5MOY7Dkx7FeYsXgVwtfAHnMdaCpX9
Q+kKrN3pJzUvZ4nndf5xIkECKKHrPQy7B6yIDd7iCowVJjUU2A/lSi7QeiyJawVrOwWlWCNtxaKC
oHyPt8RRQwQxv7Aqipo2U6FQqItbJsx0L8nT+GRm6qbtkYsF+GINIeynLrgyMRsYVvwzHhMfpVKg
MpYspPnV9uwHWJsMwsjax4ZSOEInU0QRxcOqTokBJeKlqXE8JWa+gtQUfRlXn03qnwCAHZvoAum6
5z2QZagbQcCtac4k1j1aXsVQhylqCtwBRST1QgkenyVZHeydO7gk/xjdq5yO/3FlDVFR3sSRj2MV
r6ezmnplYJhzmpaaejUgS8layT9uOp9dqMArp62Vrg9kw8JEKfrxw5j/o+ch32D/4QsD6GozWc6z
glOEsx1kKlU/V8y0JgekJ4FVBVXCgIFuiBO8ogAQkV7eqzpShuPfT62ZtQCqigGGJ2zH+95QYGl2
/aoKpgvjy7fX9sr2IqyIZp4j1p5cU9BGFITA1i5jGaBhgnzoUnjM2Y+PdW2e2hRi80/GjuRRqHUO
rp86VIM24LZJvbcoEqztuu7ELf1kU44Wyuc1/u2h/uux+aXiyoTh63MxdjxcGR3EY6gGqa4xIyMV
5wk+UtRnDQ1HMRZpjY2iJe0ifQ5ChHS1ilBEN67dCtgZSCkv0QeRBx3iiNC501ucUptweQ9ZRXCr
nd2CTUPIOhcmy30tkLvT4Jk9KgPqcUdWDOiSPQTYZyPnQZ7lqRDYY8pPzJYPf/6foDJbV4wOqilk
qEtxYY7JvrJUyFSh4uEpM9fNDNBc3zLc/sej5j22i9V8tqBmIysI1CE+f9mmHazzeGDWzodWAz9s
uVsbMTptOKWR5wGpTQv/qOutqtEjtOy9USebxbLYATHXQQ4dQxgsowiDUP6p9e5Jldajo3VXGSIR
wDsPyrsvUDt/8Rt2bjSQX/JEzL7pVt/+sQ+KyhvxjSFF87A5dM+r4BsWXZQlKV3Y6EiPIJhmkdvK
sheNFvooQndaqkvlwY5jmq35GcafWEm6SaFsSmkvwwBy3UJ8sgmVAFslvqMGzDe4v3RBTtoWdyYw
iFU333SMtACqqYUCinvkCXgwKRLi3UHbpKrCzxgTuRo0ttRnB4brrVHqClptBRR6t4d7yGdMdJRW
2xPjmJxx+QZcWQSZ2jpMhaj5IptlRqVT7W7xuniNvcvb6zxQMj4qEQkL8E7Joz1xgvvu7eAAW8RS
LSpt69p63PsswwqOR3UxSwYl6QfpYi1fIqLDj6Bt2EPEwYGHMg+DauldnCc4cWaRRBjguf8YDVrl
8Jtw6EUHvNYVA9F0XtBHlPyC0IeU+L8HG/NYAwcCcRlQyWZ0IEZUNxbrCvzi2wrA5hI/LQpkILek
q+ADWDnpWhwK2ibZwVSd5R4Hhw2oz3Mw4Drpf6cSJvQXAtkobKvzJoVGUNq3e6F3U2GQYcpgv2p1
3dpOl4lLmvPiHkO+qt+kT9PW2UN3CukWYORcwt+vMwpE+fKxXXn7jal35jcyrfD2IBSm8Xz6pmmQ
Q5spq9z8Ij05barCOEvdSsEYiaoaYGtv0rBWW8RYYjdlGhV9VoKT5T6Nx5qLOFHNXYnmXJJJXMPV
G92RwrQ0vHo4IVhzwng8IO9raEgyDqASBGcAFhscC4xFMOvznHqwwXRSnBMFeYlu/ksA1UE2HPLi
+jzXJ41Bv1iftuzIL6O/oL8FBzAadUU1QHMJtoOUWX9gXGzfBj+RIeI2mW5WfyNn2whWeD6Lks4m
S+m3C/ZQuB9VOcLpGyE147UFOTIy4ZcvZCYtCF569UMivqI1gWV6Hdi0OhVYfzZK1j75K1l6UjQz
8LI39iskDCjQx+HjVxcsRwqdgws2a0Fpy+AKOFtVPTgvU68TgmCcqxzzqjy82t5b1PWzz3yiZKYB
8SOqvRXEBtMT1djfyNO1VV0arMh6618OQyvy2lxMbmBei5ygQEQErpBGbKVw6MBtw6AGJsgywKO5
N4HDBdTUauwpdTgx68OWTYD66+e/5T/JsvdxCgBNWUyoKmRkR1Fr27/YqCcr6Icza2tGfqgZp/58
9rO4o9yFtGcb/Vr01Zi577Fjyum0ipoKEsZ+CPhXTqS+xAyhhhUb4mC0szpMtoDYdTWdmZg+/dTF
Vm22bIo2JOhwvIu20jBOMLRdgeeyPAYdbOy+RzavE6R3vfnJB2IzRH1S9TZgDnw/I6vpiyOrp1Jb
PbP6CHa+z2UrLW0pQssDMCU+f2tGFtfcNK7y/XNsCyo2rnifr9jCHvLDKhCsYzjruBbTaEJxA8y1
+uP440RtBql/ENtNuvpjMRzY/NU1bhrQPbkXfq3k4m2vc9yAtvMZ9TxhzUVDohGwDV2rG2MvmoIh
ZVHRZRkaiymm+XbgoFhW+k/1wMqjK404ROVlDI5XJDvS0tAjbQbzjViwLrvT+jMKmk2BTUutWf8T
4MSmpwpY5O4r+JmsQU9gAu2PTVT0iJqxRfnIc1NceebQXB+wHPl5tbqHaVPHuI95TAJRR6G51taf
5G/XepKWMxuRpOE/FzU4frFfbhUupyWy4pvNEgiUlY9XqlFwysTdFkSVW70uJlGW5X5/cF181Cm7
GOCpLvqS0t+cmIEiuUdUSaeRjwtX2HsOYD/HOX4wgw3XCe5UVPvljWXa+74+kZ6nkqRNiVHZK6RQ
XMZ7WRCLiMKuygsWVB6qCaZ+rhva+65957JaIA+Ekt5Zb0Fc0+hzlaY1rHrTyzaxIQbNzXI55og5
yhDvYwrVEFv+D/GZes3NyLIsdLq7kr0GNZfQWlJhksathgGkjFE0OeAI15YbMOmOT+ey9q6GE61W
CxctnxJ9FvWZXr0Pvrm0uWVlCOEFYoToHhyoTcTv8A9/7/9SefL6hfdIe1BxMkNiica+mi9YJLUb
gA4mCU7aoLndw6+0K1LBqWtfBRo6C+G/LR1dN13CRR5zJ8eKhGTRRDeGZzSiCmFybDdASKBJ0IRo
faSFQVvsWxfIHS2OOg06KWOnOzowOsF5TnlTZzv49ACd1X1psF0fRq7+9Ll/QK7h3VQ+HLoCF/JF
WKlupu+oJJtzmDIeSm9YS/x1GTpSNM8Qas8f5p42/giK7J10Hvujecx+PU+eNWL23LGvZSCMDjrw
rAWCJof+IGXmDrei6dp5zAsMWE6bjNeWQPyPtvugHnBvNtFez163ZTsgh5TUjyGITPSRI/YeJPu0
jybtiCa4zpmtElKwOSEvzoaHVc2+OuT8O1nit21qK2Duurxc2/JbCNzPPuAv6OhRKCVWGj2lhKCX
/CTj8u5lXFWMy+AwBGyfMp4TVsIEU1oAln84r5OgSFY4Tb55U5TqzUaMm3Mvkmy1mxkkCQa6DNIM
Pg7BTRM7HR44pelU7jwG8IF0k6oRWuy0T+fwyUXSNODzPuX+gNupzrloCLVktoHxIuPa3AcnOgn3
FdTFiDV4zGilttsFVWNx9aCIULYvUotkRfNyeKEGjHZ+4DEdcAcwak1pP+L7fJ+qRtY8IBXKjWDk
KRUFGOzHdT9NAHYrZsQhYwiaqC2SIDHwll5PTEDlAZ7t4UTfQbQDIoIEZXNT11E1mEjDPa4xb7Kh
sgrO5nDH2OsWqLyi0LfSsuplZXcvZ7iG085ehvSi5V+cRKlD74nMMTVs2GxebmGYPQPgE2IbOMBn
jWND7uxL/LE8PawyttfAMybwCl9F8XmoWIhfVqIH0+xTA6PFhA15HRS8i4tPY9YEpl9ejTZtLIHe
rFyrr5yhePcxTI5shrq7FWtXfWqw24PtpLvW7jCT3zOVhbUWCHkqEqry57W0fkMK4Cjfg8gle7Kn
vY0vqegrQgEmTnPTphhh+Zh17Jl8MmabiOQ3iQJuYpyBkv6evnLoMw/28ot9/Q6MaUJF5p9mZE/l
4eFsVNfyQVMW4EBBHZg07ypqn9fzZILKjvsnuyOmbYKq70R5na0Ge/cjty4hj58pGCKvIcAOD5Wn
cZWvw5P3OF1oSpmiWLshyOLpy1eYrKm0NqEPfD9cRCi5997bwuuosn6K8rwhHnFcvU5CgQ55XOj+
Qydl3F6rTTmCIT6nSr5ZMI1yELzAg1QF2RU7/mE8WlIXiv0kw+Qw7RXTdN1WLStu+1joOJAf9jYe
3xc187u5V/wDX0VegRKpKIqwhnz4x4oIlKJ60s7034i9/jaeZljckYbJbBzlWSzt9zI0GqRyIBkQ
UC4/yEvY7HoaPVFpBeXnHlSqOki56KrhwzMuetuj7xc7LwCQXoqm9PrJJq/9sqEIy0Y/L52j29rD
CABW1bjhtPbbV3fDHfV/4eTYmZ4lIcCjLYJlJzz+BlyH12RHboOni/CvTXRl32ndZZDxzmKElCRi
Ugc9QEWQZXXDMn9/i5HvUfeZc816u5eseE3EJS8kpHFfx4/cL31Su6Ph0eyx47vS7II+cVXIYOI9
s9PEh5yLyVJezAqzl1LRRoj4srmanc8YkrW3wiSobf1rNe8H3IiUFE5l/8V9ecY1BrEHNNYf4xik
HssPAuqj6XIqgy3E8mQjDtcV93/HVlpD9XvAgVxPk+0k4trZPkjeHsvZ8wbQ8yDqbjqsQU82QrxE
UW8xfwuZXFsSWTsNRRBB5vKHq6TOIcoZ0b1XqL+arWXQAVEJYrHcAFo4PnAp5ji0wx7viuuKjt/Q
/HiJzQUhkk52aYmp4QKRYS4ua5krcHQ+FtPdchPGGDUOlnJqaJPqxOGwJB7pavgNQCngeyvkLgtF
u6QsQH5z4YWgP190Ziz5tl1GXp099EewVWZrJP6eGFf4cPUTdckW/DxNW1/cVy+GWqz1yMA7GhgI
y8NYQHcPLrGp3ceIuWy5O9pz2rUvt6CS9WLzEmEYrRjHlikER2uo1cuo+fzoswkORPFBBzc6FIWw
lTR8U0haV49fCpCaL5O1u0sl4AWVztNKXbZ+NpT/d9HAp46R3d3MamQ2e1R2sdf1XgWr6WAzDkVC
2XoLGCqx/utJSyo6XSE9iCh+s24kjaJlV5cZnVkpj4z2IONZ7+NSQyQl2RhRTkevm4JVrrhDLk6+
s3T8QdQLclgsexDBN088hyFly0+I4+OmrPLsyDG1UnINFBrVYU1+Mnwksew6I+GO+xWWn/rTl0po
2oE2Iu1av5yyec1DJCOm+9rO8LFpXPK8r+NCfUPeEpJoNdNwS08yzQodj7ySojP87oRZNMdRZe6c
YyAVbcWKykRIBRz/5t273LBdA+yq/aEE1vW//+7MSm3Mjijh7D/ZcN6pXcJfWhidoxVVUuv6PWDU
V4T2MDVvncUruLM9UR0msXeGmVtUB8gm3KNfF3euokD5VyYhVA+K9ay4OQ+VnoOir6TZKQb4Gs66
StT26b4+F4g2wSeK59pGqGvtYuDyYgb6zb3l2PNG0YNfU293XbeAzZRBvLu0mxxy3ZlwGoKlj1Os
m3eGFXI3c7dXZ5ZFURrEJ+QyeuRD/FQl12918NfN/+VOuD2wx3yEBXgv8dCUP10DN1HAMLdsBlK7
Y172Qo4a/sWyLbvMHlSODhPdgnLM5rxIatPW3DfntAxLDCcrsRD8btTZuMdioQf80QviadH5D219
AHanSJ5f2NwJxy3f20+BfooR022Tb4Y1KiLFHCOQe+dhu84wNm8OiXY5qyVSD+YBC9owd4QgWZOx
J7PUHhuV9pPLxxzqMAQm6dbGwZYaH04U3/VUAaBBPxpJCp7J+kHChta9gRno6WhhIAqLXuDkHmZ5
HzKwkKEoO9wkS9GPSIktNX/tHLFYQaLX4qOghKipCbnJJHLpoinFAkHcZs8U6Tg/c46v4kv0ZxLz
Kxpalxs0fR0Nyj17VBC2zwFfIDXpu0nlaiVfbn0u3q0PV6ulgpdr/OwlnFF/0TfGZQk+uKovtQyd
3/6bHmqjSNLl3V2sq+qGUEOFvNyW1BUGt0AYNX6Z5cfesQ7gRTzbnm/Ei52Zwh8HaBW1An4MUFs/
47GBfvPvoZmxW/2TjGF1xnsGxU/5w36ZV/IDah417qLOY1jsZD0Vu12Y9qEYfEtxct2DgCEy8KnH
P9cuTiEVs7qjoEI/FYtx5gD+lvbwpFE9AQgu8nj2pSyTmcoTD95q0keYCIWH1U/yBzY1ZFvYhvKK
1+JdnJDrFr0/UAKeHtb9N55LvlISOQa02awUwr+CDQlMvrqrSZri0j93qzz/aweziJIXhkx5a6UL
AqfnzdfrjWJYBSnSdBc7kcv2IgMUFjiJUzRjbkY7eUiyQX8G6/PNflSGn/WHD5ECCWfR2SCxTu9v
gzHACAGSEfWh2pyhOcXvKjaRj0WUGskhbSWDI6630GBkjrJ73QMpY2DRWc8nDedbZdVFhi6/n0Q+
hXx7vo5BplObUvXQmSRA+OqlJng2L8d70HPobJrl7UPyl4KlBJSwtPkd4Y+uiLwWMcll4wu1Dihz
G/a4KsVpN3e+Su3u9ed2Ns28S75AQWJyJdrgsFJcr+sk6Sp45Nz0nFZTUPj7z62xKG+tTIGG4Gpj
dHiTUA5DyIkWfUeJErc7umyXS66Zr7kfZisRxG7GEYXlTResw7xcXi/xxaWLh0MvTSeh58S39/tI
KMBH22iBIORi/9fWOTpxrb0W5X7vEKkJPzTNLmleQGph3RTSWMR7ELFi0H15uyXKB/YXvQFZxC3q
1WeS8CnuEVfjqvndDsUUeJe8g7/rZAKAt+VntZP7UHl2919m54siwk9Uug2ffkO66yRr01RPb5T1
YqJW871S0SKZgrM5AyWrdd5NhHmTy60eQIn1tWofP4fbghqYaJdOa5Gd9ppTd25YSU191KLkqze6
vGLrLAqHN0UM0yscdCj8QsCgAlB7DACHK8k7q8jrEgBNLGYMmWlpYEa17V/M3XNgGykA79rQNN08
iFUmekJ01Lh2pstrkwBvx17+xsXPRLslJ8mHHgha+MuHfZSpmEks5SkV4xCltd1Vw4ehTOCnNOx/
T9URx8SJxT+ORX1f1KiI/GUZNjC70OZEx+lw+uHleLNoyOZl9JaXld2fLBgsO5I0kh0skZBrO+5N
VlcDkJTL4/hrzN4iaQsXC2dSH+m785DRNLUKzNEZuRCS80JWM2QO/vnz4b1t+TmxWHyOFonIzrYp
tDVcV51LM/dKEA0ExuUVjTzulhm4vhqoW2qJuVr4G59yKf/yUQiU+GtVIROGxt/plH0cmZVwUWtw
rgFybvMF29rHBN0thJi6NimpKPPAqnowGqwFrO5C//Qk0acVmqXORzNyjB0fZw8ujScrVyDSVg02
TZCGBz/8kawLj24wLIjD9DMd4QgqZOEtYWdapBZlXBmCh6dbBGWZNVOe9X4C3mvbOop5b9bUcawE
YYQQoRONS0kzwjRDObVPL8GxOfCXTxHQqKkuldCXgRNUo0Uk+u1KIYOMv7tsCNJ+XlbJ3O2JAIP1
tkligObApp5g2s/uU9w/rbayWnmMCTQDWvu7zgi9qywxRxXbZ8bu0J2duZ0wFe4+1GjOzjX2QBx5
QitL/tSraMrHhE/SpL0LTwDokvZfJi8+OXIYYdSfbpNu03RXStgvaBuuq4dslbssI+bWdMyQ+9Ou
E1KR+yv8QN97YcGgZvU9Jiqu6fjR+d54wdAaJWaYAoS+508lryx93FU8iofwkZRPbvJpu5VM83uk
sbJ7QokIiZhual3+Tszzab8mZw64hhDz8zVGSPNlj1cFMIdPaw07ROuoYY+57jKCu+vcdm5mwYdZ
AqFkmCM7ZuGkl3gTWmSvA5yX3fBxy0AIu1s3pK3UQHFWcR3hC6fZ/jmB86VWILFDg0Gpid0nSDhq
X/p4tbRDkWqsRErCFDZzaklP55rN+4jkqY6Wauz7wzPJ88ncWTabDWw0D0ggdwPqsOKgZEOm265u
VWL7VcvtD3/RQBAG1GzkdeeW5knTIXA+1RL8Q/LNpb3WjH5n3sX+H31dDoUjx+3kwsan6HlcBfX3
QXQ42A5tj4Zh5BAaIeFbKUsBviIevMSlqdWLKdp3STtdjnNFx2/VEMl1mIGoFs0xRiH2hfgnvrmN
jI97u1mifsHQe4pnJ5mhKspZJK67S3gO6CPYMWo1WvE3GpQdJZCk4+VeafKb3H2SXdELAP/gWyrc
1icHn8d2x0Di59JYXSlQBhcRyZfY3lilSyrh0CBF9FyYunCuvyvHhmRtizE3X5+V5pS6qm8lAv++
N8cwH7WXm7A8M87VUY313nGGIvBa8CiSTkEVlVIfuDZ5xuaU9RtHzcwXvbXa1/FNUkgtD2SNks6z
YF/Px31mcVkqUBk1KxxiPOjcZd/aC3yLG9vzHCUD+6YJpUeRdtpyJSRObU7RFWp4t9nk3OkNf8sQ
D9sEDiDKbWm2+wHSG96vKmaUUup6sQ9W3U5lEo7Sy80tjKRSvkpKu+ZXMfgQoxnkBYafYhh8ktir
ZiOESRN3WIoW+VfwBSv8BHOW3pCegT6VxLdLT7RaMQMFYVcg83t4n8nT/zhLrfYCGVi2JU0JR5Zr
fBbC9SF9Y9KIqAAiBKhJku9toiwB2VcrwpD4xbKvL0PGHLKDNQPorfho027f+v/AOcnStFeLtVkH
SG0pN27nS/Qtf/8jiYm2fTb4LXMxbKHWDFzWoReCpnFl51TW/7huelb+WHq48wyuLLAJ3L6aekBj
ofj6baX+rmXRM7leI/x5VV4+TDhGkyeiEZE598VVrwx0imt0iAqFB3IPLHU7J8ZExPbl3MtpPNdZ
mkM5xvUei2rEhnyxLGCemvs6W/d90Zz3aI5BxdAerCdwzp3S73HO6lGi6YMAyGNshwSnw3dfJI6m
R+KJOJNPoHH2fV3gOCKVfJ/8P7PChUuyEBJiuoAg9x8nnrDlf8TzIL+mrK2ohsbNfyvGpycRO6ba
yu5cgmTwPvSiwjBPtz1l6hm4RbwEAgaLcEeF3ZbPZtzdUFyhjrg6fHtNEUYsRPmKNZ4d/gG5C/zT
G5VKS8iQzgWjWFruZPtnLj7GAj0qn/uM/yvd6L4ekVkcgqfRVOkTgA5VqngmvXdC12ByIOgK+Ln4
bd2hZNmeM6yjlE413MN4xqy5PvWtGHz/veCjMR126Eqs7RBHPImYdxW3eYYpyP8sSepx3gLEMr5Q
SH3qKssUx/IYQje8ufUcAxGoL2zpQVdNkC9Nzr27Oq1z4JuFDUZ0y54exgIoPnmXRp/+2/dlGjpb
4vebH68vsJLepuU5J7Bq43d2PEh1ennE0sHlsAo5lDwYMqv13kZwmMXKISiULStdA0Vw3gHy14lr
rzoZFuxsOR99wu6nJDHhV5eOdXjbYWtFyqLC921ins2ZKk2hv+baVetjEc84ZCukk84SQRG0bjSU
G+ljg5QLeoi15lAYgj1pp7cd8V08K/gDvuy4nVN8NxWawHPshP5Sh4LCwttV1PH4Iui56Y5dNnAl
tXBqc0VxW/F4BH7kn+5AmtgHdc6UmP1Sr/UsrfhakA9SHMUVGQ8qaGjRC8LNMBrVNMM33QfV4Rbs
N2Olb+YXVKJNwQ9nUTAuqZr1xLXx3IL4ogGBc2WPp9UCI3YOY12akBpkhLoj8qUkC7HehY9C8wOo
RBKS2gjJr4u31nUtXbjUhhgj0p06eJ8m0ZsocTkrok6/JbCaU0MR77i6Q6HUREcmpp6OZqe35ZCz
M0uB/jvaRy81s5V/kOzQMsj96FAPd86iNTUzhrVeHBGvexEWTagY9vU2ZlxqYtqcSB0djaJAaaEy
LZFgI/0+7pzvmZZ/OwJRih1LwxhX30vlPOH62eSHH6FHqRKpS8BsDw3oC2d2vXj2BVvb3cSKlL9F
e83k2Z1vTcIg7Kk6Avk+GdqqLH92zAFQZ2miaqK3GrefIs3El+aUkSxsXRkaCLSks4efV7xItRlR
L/bAwUfF/y4AiAD8by9QKLpyzAUi9xYQ9yftWHtWl9HEuPnRA5lMb0NomVQw6iz0lWh41ZAK/unF
ofrDNVh8qkwHazaKQnlt+nmqNa6uxtAKb2cXk0IZG4PsnhQqFZ+3T1PugURPwAOgt0S+HDnEmCvl
6V4EWQtFvD1FO78KL5hupEadUJQXcO9d3tlIm/LJCNGHKwUuBAJ/fr1mJ8gcMPvnQomlCOQd8JlQ
45t0ORy4Tc6CYA2z93TCqRipNFtJR1uSqJqZhl1fx2QNXjRG04jIx90u777yPriQhl5J343NT6+2
Xp0WrAm6+jC597SBcvhkZeUiDkRkSaYRcqMHKBPx33/q97EhxYfRT0RtxkydhHCYDZOba/nmVf1b
HL8w/kx0x6T4Xq5zmcdyE8abH0jiQtRRgBOn/9JHbFOsMlM5XNTRUTRA79QC0R6VBJBW0OxpBaY4
yTTptyiIsy3zDPRtfjafpj1fnAef9BvaB82/+gXz0xvcmRC7ZI0RhxysDMBNgAa5GpHNYtpcERGg
kF7/aV/a6bK179acmlLyLDqEplI1HlSfMJh3XPIoIbl85IqMIOG7MCdQEDdTuAjUDiiBMDt6grVX
ZuQAq1UtqqkeNZPXuJcq8CENDnmUkr7+Ku1JWN/YHlItdgkQDm4I0Ebj0XO9wNjkBBocBYzvwE/w
PqNZSjvunr2kEmmW/HsUQ1rEIxVgY4pDEJaBWT6mpADkzNumg+snjvID9zB/T0wmgIm981yh1cT9
HP3GOZCLDm5gYzncXy9qFPsGJzg1PUzTfzmq6SE3S+mv2rXlU9Wstirf0GYpRpWiQA+zobC2LDAH
hE6TE1v3EkS6JSgpzmwJ0nXvrjdJCsQK4luzFeffQK030ohc5yL7dhgjXA++K9Ry4IkPiuI6Ip2X
Lv7+PL1qUxrFWSD1pqJNkYWWyKUpljKh3ZjeezBcFZSKtY1eB/nHIY9kXpu41y8KU4/xok2dnRta
PMiWP9N87Jm/XokmzsMcP8Gwmwy/MEzCBjm6PWm3KmB7bG3UBGIoGwYvwv259hFGARwTJ3DzQ2iR
rS03FLEaFZz1vCx03o3O7UgtjWcRBTAcSfO7OYTJt0eTPM4OatWAvfF5pPqZcWLggmQxgmmzhwFN
KZyuFoXZFBa5KziFMsl/gWK+gYTa3Z82Tqt2BbFstWkDgJXkywxle2E5atx6EeWlLw2fy2HqtpeT
UuygdNPuNQuW8HOFtfQEEKU5+KoTa1nWe5vZCR/hbOqkhaVH+AL1LsF5oVlekv30FAtAdI7Vrg6+
PY/ZhnLvknxVuBiv0n60euTXA5LNRYZ6G1L5irIxlzo6jH+onlkPf9S8v5CaA/8J+9MdNQKPAibb
H6HhrLDpZ/v8pmhUGoG43voFf9Pf0kOWs+jrN3L5cA1Mrx/kKfV1rW1vXFV4ZgAN4ICZwqUkMw4U
pKRuHR0mpFSWrMr4VRSDROsbkaogVsHpYncAgYupIYjlmiHG8fSd5DI5A3U2Mwnvz8G2l2oVkIV7
WY8WYVKO7eSn/j5DbwhQwbEWRl5bLNQjqrRf9H+whbVL5ZPD3QtVLJ5ClmsBlINp6/cGFwZPu1AF
d8wj23EBpplXrR+FjYQqwnN1aVcJNDJL21BDaolzyxuuZpOfvh9ZxHcmxzNYlNYuy08m7KG4k1kq
qEm9esmq759g8ebyZ/iEqm4n13ndxVYmayxwHCSpR9sUTZPN9eawlC6rEeBzYf0DNHrt51x4FbDH
kGVGisovA7a64vm9Pas1GGdV5rtXXTUYkwJw/8kwnXszpLllIxlWVGYFaZ1jtt6PFcmVjoS32k49
8v70yau2KTYIeZJT12PrxTS7VwecePP2CWe0d9jhiIcqshlgV1yGp14ngAIq7NfL8d/QsKF7yBLk
mWLWFLMWOCwChbfngqP270j/eo3S3RjKvo7tcuEdd3Imw1tF5KpFBks7MbndABhFMhzKgxdnZXgZ
cMkIwsafuDosu13hjgZUDdxiSlc6JaaUky56qQsPyKUb+nOkSPWsMX28oVopa9J3Hntl5hbmd1m4
0xnecf4vUY4AqiZ0AmLby24UrDCoo1gl2BfZ1HkBvP+cUxhwgstu6X8JuQTx5Dzx1/6SMap9pKTn
dcBKJzBl7ZkfJCOeT46UP7PJArJ5w0FLCR7BK09dldE+J2PAlkvIZnxHOTiqGUSylLk3R2N3phia
GCraQCKOKVVQJJDPL81dAsljVFI2PilpazFmAhfB4aWuF71kQiQZcBLv39tRBt31AqEPnEU1wu1C
5YqMMy54WtOwU6PfCBtDQoYidQ8S9lBmuDERtr7Wirur0wBd/5g78QFTufbBAC555iBzZBMzlNBv
LXVhSM06b84y7dWiGB5/nFxeQhhtzqSFYnogtAnBWxeaO1zeLeFYNEoTUyP44F5hMpIDrHbEze69
0l7aX9hzaskzFpKDCJvLsMcfLgBI/usLwQ4X6ERd3sgPuG3yI4MsSMgDC3XRGHOPiQazOWJGSruY
/yBXgv1H6cwChmgQQwxguuGkvu2OzPNdxuYVg3ajHkyG0E1PdtBN13RUr8mMJFnqlc7ZUBsWoCCA
eXtg/y84nb/6Yyb5zxNUzgZsL8AGvkyRDdQIaQuno1MoAqqNRLLJaFQnqJOBxDhhB1Wvz8oWY2R3
bdkKX1Hv5+joyGu3c8aT3jwjKX7TswYMRFV8EnXsTDcm0F7WYITwfPwJNwRim0P2aFHmKTfjj9af
KG4BeOjnih9zMTczNmqsd6lCrrzUkauQxJCTibdOMhm2SCJVoVUCzNIAOFJ+Jp6mnHFrEcX/8Vsf
tS2Tty6bVd1ovsj+yooPxZCuYPUUuL0a8MWUsvpelsvTD7YoDvYEtUU6bH6G6RrhG1AOTaqoXhb8
qimPJ08n82xa9v0T0KextCCJJHD82HEzrZdKbmfzE+ds0Hvkcmxy03fMbum7RVHzx+r7tYWo5vfN
kxQHPwnZRuyHSgBBEwqrsoouEUTN/M3Yac4UD9uSHEXHc5ideG088I2ePDISpEHlhoENfsrANmmL
eyP0m5yfC59/rI1/34nHUMDiRo0Q3zizCXrbQ2MsziAU7jkPcZapKSS/h/RO32qmbiLxnwLskzk1
X3qrOmRdCWJrFeNNZLBYaUEcsQHgfCBOwa6i49/+m2g1VUgeRIc2xyqlnkMCLuyuFmHL3vDXGxYv
19OPqq/RLzGEtjBdeC5IWOZyj3wC1l+oz+/RLuCGAodYNPpU+PnpNhDd9ZsSit/ZKv+FjITB332Y
Nwi/fKf9LObFZDioJKJSZGX6t+1YfGfEo+rLpZnlylRoFDLfLvvxl2gOsnn/3wUmw2yeCq6Ndu7q
fpygFzPpSESv57w3cGFFdv27m06zg07xpZhSQxOxzsMCnrgfND+t1XZ6cT0lJpR2A9zEcxTm2LZt
dWUuKjq4/gkSAKYTRm1UeDh5+XF6eCNBI55ETziLeGkYLPKfKZBdUsH014fRF11fahCvlgfqy2x3
LtraMeBWam7pq8o1/9Gsc7swHlViWvGA4kVqzCDmWZQdhKYXDDVRE8jETpNmLYYIUq5ld9N2s1rt
4QWFS4R0n5p2LYp7vCTz8tOF4M1j+uzq61HGIBHggtn3HDPKG4zMTlTPBSf9gMs7uY1LUY6WicIY
pcxCiOrc+ZBAyFlsrYs/K3xg8aw0WYXKQY5nyAtF2Yc2VAV8MJV3skvQrgybwZYNeKhYBTi+44wH
x79z13zz5wH52VzRart9WSmPxjBrkVhaUln0JaOBZivRPotJScefHXcvb22L35BEXXjT+iZ+8mhM
B0FqtOHgrZXYbeJk3HRUxqHGwuIlYsDCWvPXiFO2AfYSAdzaZI/6LNQ7YGWY98nCTEzjr8M59sO2
Svxm8HBNH+WJS/w87SDFWx7oNmM5s8pO5mIKdRQQnS7/RA3ClByK1NkhKW7VIiQ9BmJ6gTODJV0Q
YqrwVJ7Rs60Sxynn8Vwz1BDldAJBaE7Csoys3sHH0k9IPVr12Zw2b8pgXCVxxYHuTjdJoohMQ5IE
9F794iWts7ZQvTPD32GaYFaNnSyVla50BFQiLLQY+qNY4jinC3UEMjVtBx068gDTKf0DAxRpOFIB
98snJPOKo8bE5LO1KJfJSHCdFah7IxGoEJmUuaS83lLmKdAHacCWP0MaS7exzjo0NZT8kOa8hjOo
DlW3cwDvrlJDhobKAO/l/CZt61z0gX/WQUafUskV7Ei6xWI9vx8yJhyf5yPX8clzjHwpTaZWZNZ/
bUOP/c7VjGuiTkBArzpfk7NMT7hO0l3UEkIzLArurq5G165o91hetM4vhDX83nfBlUQXnDxnVNfV
+026NQvqjb0TUIMngWRNctMuAMXZAkwdXk02gleJ78aEIP5O3xEk/VYISAVPyXwYzmWVCDANl45e
D2RuL4oOfYBCdGCyke3O5fZ0QlfoBufgKqUyNLfrnA/EUnLZlDL4fqCmOaLNtRCDZ0s5DDJfFxP/
msQMHCcf4YU/vKBii4NyFDbKq3zJ0uDVOYIqXDiHL+eIMT1SO+dXe0G30Zw13wbEcOAwPCSIYTUv
p/53mYgNF+eZd7jnAZwaXH6Ya7X2KL+YG/4wna8eeTDCENX3qIo8TyPNnf8dkENzdqvOpeR89pja
l0SEpQ9Re1ggEShGxrHppEjlhXpGKVpU/7FMSUWoAb1smJ1PzOPzU4eKILIP6Ha17B7EybxplU0F
Ko24mQFixJvp1Yy1ZOorZajJucsJpuE3ld0TecabOWXFEhbyV4VOmE1bd13d57FvC+Qs/AX1xYF2
WuSDfZXZDw/5MMGNeSXYSSPg2KgzjnaXw9gUl5P2EQhWyMj1dSiL8FeJjxERMHcidP35f1sbGpQv
XkZpNNjyGoWaoQYIJ/mdQI9Y1O6/H0qU/ZUPXTXalw7u+XggwpImriDITAfVadvhnB1tgQMox1k7
tJBc9zOifAuzeQKOtx4lmEJiypy9wBGejIIWQElP+W8v6Qjh+8ChzTlKTtwN0zTmiBC11w5ZCpvh
+6xJJW5lfwxh7+8iD22VE4RWtsvNWLikAAFVSmC3KkwBwgRdeA+lrVjgctGZNH68Dr9j773TWhxG
NzAA+Ctcu4MoLBM4n20YBZuFzhuNSNCo3HTUgiIcCCiaet5izhftutzLB+EkJVacKB0LdwJbsdI+
w36Abwr8pc2GAowhrk5uLLRZYu5/JKaRiTd52UhhW2c3jL9p2yZ+VLkdtTybB/Jxn0zlj0eysoC4
55ZKp/tDRXEBbngN0zEtFN6w67c4xWQwVLrQzqkVKtuuUQrt1TLAt0gOYsoT1YOghdj9BquVLCs0
bATX7rZwu8XvM/YXiVn8L+hm1vJWScdyNd3sHzAaREDcAGQoNzHHeEXryfb1/fBYdqoQ8ya8l56s
xE7tIttQVAFCsQIDAmnX0VUaNpsNjCnF9+h/qmdoS2vzKw3G+FPwF/gh2mKnD/Mtnr4oZRP8yNVP
MnaT61dBd7kF448mQvZtPNubzepiP5bAU9CoF9geXL6Yh9qc6bOe7MHzA1vhygxKwZ7XXzacgGyk
3Q2K06Sd0eCzgPy/lUSt7O6nwsu+i0tVA/gUYMa5RG7g2nYKnUibaLjKsS7xMMcwBEpZySi0a4Gu
JNeMe9M2KNheniWiRznCmrZ+2dXJZYYsJAInSlb1nQmOSxE1ZAunxO6qpqGKuAoeymmJX5DO8Ho/
iwZ/QpKwplOoI2P+vHiN80o9Wyf79EFcRO38Ne3DvQ/Igm4Mm0Nz7KMQRqiFOydAq97ud1JC7tRS
MbYFw60kbVgaYwNx8Kt0PvmWo5e0k/r/Jjg9xnSoIp5225hBvvqkQ7QBPAof57doj+4iM1OwyOly
EfPPBFHYZcLobNEKwpVRBnVuyIs6L6WfYU0/ts7BDFrzaJin/uZ/8qNNV9RVccDUpjXwgGDEncC2
I3Zuv+6FQXXhh+pIZL5JDrZRpVxT8T10xVCzpfmXad+gkGS7vg7FgTxZ68IQMMrls146ifXZE6IX
p3jkcDT1ZUV0+OJUD5XtRTFnAFC0yUwuQh4LEC1Zp9lVe5Io1AyADkWVDdGv3DkU0hlyeG4j8XLS
JTBhHnJSmvVJ3CZzCLycvc6dpGaFHLygQUHREKVsuCQ/h3w6W/qBEdlG8x4W4d+ly+XEhp+Cu9cO
n4kMByXnfdLA/4yAyNQ9lAocKKe2KtSQ7+jtRATTCmBW72GmgldMnJ/KZy5VyFd9xtEZe/gKwvrX
AWWJn46aCKY9FCIRNwVqQNhCqwzXttJuPAByZ2MF6MAMRPI3aJ55GfqoGmdZ+IBevuvyLlqi/XsR
hSUzN21l5ucUEqHx0mDZy+Iqurg6ygxH2yRuVqwusdu7BimsRNIZn9mdGnQ0tjj86IDVx0l7JzAM
V5AY5I6zlo+SxnlOjw5dYdWT8+XSJWNQ1dK3dMGnsFs5z6w7gKKCGe5vVcLuqzyT1fTtdYuEYKEq
Sw77arOe9XHfbOV7xaJUr8Bj4br9TNmCbzfYU4XC23Dz0fmt/kKQc2GGh3KTwKZwUHbHEbEyKtyL
zkODubEE7X1Zd+S6Sw8q7K94dAZU6ffQDymchdkIR+YBc5UtaJdTOr3fALEr8BygQMkWHp4tDF/n
FE4u8vdJsyyPXt+XMTSzFODt8V4XiYqrcKwsfmdYzsS71zBwuRg1cvhys6hw0I9EZ20ktPcuwaLW
lWhW9lhW6VzyQYnWZArGwEiw+s1WGWE5ngUCig5a4y09aoTOOen2JCaoySrcxcYkh6fs1uBGcqAJ
6QZegQXW8rhBI1X4hoOMejvAa688iit8gDKy4xnE3O+R9rRm4lLgXpgz4I0gTwyteItMBZ17FGNd
FgSVoeqOK1zymVKD0OmvbdyyUfIHhCKNr10sgD91+jm/5ESr9hkjMBsVC+f8BjuZ6wWfzwbu+qXH
ZMQclzRz/M04LxpZl0bFshF/iBiojxPa/GKf57CS9T2sQouprNI0uhNR+IRQicHASoQo/pB8eEtA
hI1cJFcjtCuHmPOwfCdyph3GDRzdHvjSQDiYULyhKIOtjBBivyeCCiJwk70ynU71hfUVOI5lmRZ4
27YqOSjxDJgWzqnEhpusi3kAE3Wdn4weqQk5ja7UMW75PgWZDJGkEEYS0ETGFp8z7lLuD+vxXIdH
F/fNq7PR8dBg7TvMhCG2WGHt3Dipt14SqkIc+0NTxgGU+5DuHEx2BzoLOPP1mbgYz0xFziKm176Y
jvqQyzIbE86LHvb7+ujAak2NC6nlLVe4D9oaRdz14aJHcdWrPl4xj+3lrQs1qb7/JfM5OozBTFqk
kNnYMYaUKnRLgHRvsIR9+rYAAe2CFhF3wZWL0nIDkQEFSeDhGkaxvO45+Q+EJHVS7+8qJA5xf6/j
NQaMOt+vNjHLm/EucYMImHhGjt1Qal2k1JjUlCvTDhgjaL0/pbgoEa6TSQWhav0epC5pr198msUO
W295UN8pTO8nz1TzpgD1TvaXN9BpnCjY81TiETwsMpaSh6CvUa+dmhmRkFn8kGSsAm2lWqn9dVJz
nIZHhHvI0iSLjAizPoW0QpJo34hfhAIS5OFN1lRwM5Hean4cbk4Jw53xTvyriybbIqMz2SyoKrgT
nm8rA+qaGeCy19nJ3BCNHLP7rVWmxdLJGXhO/ZKgEqOKlyiYJ5AlUU8tZAa/u81QGxEvYEisIKZQ
oR78pIoDPAqS246eqPFemlBmRYIp9mNk3cypwFkbiaNjbzBOIv0+0WsKJVQaxa/hhizZdWxQSzFe
icQAf3+28MDGmcsWRB9eN8AeH+tsV8ySyfuPxRM0Au5Lqh4NF3+e/JiT7FdOO1Lpfr4B/ouJzLYO
8FN6hgrDcUhyPSldseYHEa6x315lFLfPz28f0ofw0UDbahS8ES7BiW6oeir+7UWAFbKVti0oleD3
4IUhJnE+3kuh5DF+QSzZtUAbfpvnn7MNS5LcYZkvdVXWFctbwr900Mli6vXNJXNm97ywOgF6MeTZ
BTadj+uCfKEJ2/0eiW4pAHFlv0+Mwic6bpzOA0EDxOeayo9WkXEnIo4wb9XfTXI5eBk0RXfR18qZ
1IibpgZsUw6/BtA1tJ4Oe5cUyboDlcPlYhwhUhqVcis5eQmqHyqwpANGt0nVuCBH8sedTJi6zV30
4QPHGAQUsehop6+IatGqmMC0/Zx6C/Ldj6nXQQ65GRXNd0XpK5KQUr0ykNTueZ4hODBJ0hbA40zL
5YQlDsH77l+rMvFYfG7/T0a8mwCSRAdRLOPB2qDJgmR967nKEd/gv4OWcY0+fEyJZDv8neifsOY3
KDDlrMpwXW5IknWrp9oy+J9zNZ1vAsC5aRk1alKFtlJK/1BD4NRR2WnqKkwl7lJc0/1Zosm5+ocy
gcImMLWHBgO0Ngf2h/DNRW9PmpVv01jx9aWxDOaIrtGaCM04cSJBDfuAT+EN+lpU3fozhTbth7M4
Ai/KLV3Z1adAeXSSiIt8HWFjKm9wbnvLBtlBFLjsrjRaCBPAf1CVcHCsetkWUYebJLdsYIBR3SGV
S02K0RzWfaNo0CVW6mCkDicPYekp7DgeDwKgX0KwTSS3XFpyWfINf70Al1don5a/3VctF4gHE1TW
ClygPVJopo9+FFPYdW60d8L5vM5Mtf0qF85pkTh8nWbVrPy6G2jO7Bi/4h1ZS5xj9gRShD8ZuZOH
f+SgoR9Kr48cTt99A3C6XRB4W5n4m5GYNJ8VhlQpU9uGaSIVzkauFYXwl0mU35X1qB12ejwzxBon
zC4CncU5XsYIeAUvrqCzJxnhaGtGWzR4v0fd1tmaDPnXq7J4Pqiv9W1QI1a2a/EInB4dN7yp7WGU
NrV5xCQfBwQqmw8CROFifEWeQ1A0i+Yb9KFIOuHUsYmEEEbYxm1TsJgrzPEng6nDgJeQC8QChNvl
OtDGKJOwFDoB5PCWHcfKYQmhikIACgqEdSv8V5bqEtEpzUtRZq88cZJklJymB37DwU8gGykMHNQT
BKx05o+AKH0UvQUhXx20nJ3BFMJt1rkQYfFhrIg3qVRLJqXbttG39NM9PvpoGsx/NBB9tLTIsl9B
Hjlhajt6rztvwXmNbZUGdF3iivMS7/PJlyMa+IXb9iswii3kFGOlRF5y+FpnqDIPpu+E4/XJZ8J3
mcjvSw9eTotgtiWrU9/ktXl0c/kDtbjCNzhHzPo4UlFPVvDeUjh+6eF8c1mwulaKVTTjqk3XA8aE
sZBst/iZ/tX5bB1ofloUc6u7ttbunS0jbkczM3nKnL7YDFDvbeDycoSQc55cHXSyhPrVxLcYqcuP
iKVa0dN6KrZH/Z0SfHeykPyNhvpeWFmXVb0MQjEgXev107CFOaguMTZ2VfeS0rtnf6avdKxAgjOy
jTxVgzwmmCR3KuRnqMm48HYM9dZSmQUxDnlW+z0zwm/OWtAJ2f1NFrYkOjoshRXqfctg939byQ9Z
xaOUpaE4PTzFE9HJWeL4tQ9EumVCv/pGNpAK8wE8HNGTuRoffJKEzWO5jLMQs0vqGWZTlEuwfflK
zyc3rBU7erriE0M5+0fqYMOotCCecUCtLoDTFV+wNaUDQx7l9JVZrvStrbJzV/1s5UIXZk0FdCz6
2sIhM9lNdzUyni+OVwK0K8W+K+bY3woBfNJOM687uej8aRiqSmpeuzJSCwAu5+WdpxsRAG+XZYHX
MIEXTkI6viPcYDd1jImW/A9qwQJH76UHtZdA2+qUrZ0YzntMxXKJ0wNKvpVDu4ybmAEwUKh1z9Q4
slhvOqYvPIn8rDPcp0wbWh/OEF0OYJGVfzPfDOaCsUhgwTBtmN58jWRZgSp/zuuG0uAc3GmRTA88
gqxSEI6q3/3q3rt82rkwrmHKVdqSSRu5GfRT/o0reB8sSoS7oK46+95pK+K+8ruuL0HiY2SfrF7E
pgNB3PHnI21eMeKbhXdXvHEdMH0ZDxONFC2WS9bUMgFJq54uqL7MEwVQ+rRe64RwpRG4p9xQibDZ
muuSkNb4vSGaxqW+r7DZFkEPPuhBhGcqmBdsSwUap3B7V9nV4Wg4LGKcTTciLinLKHGYmO7CC6Nx
Rc7Kh7basjhdWeyZCq5TVr3g4k0vWlw88NO7ZtBi8RsrK6RCJyi4YA7/Tns2kPXwpv9EryP2ndqv
lgYH8SCLTO7G8AYaSFOzgd5Tzx1/A+DZLQe4e3LlDyv8IYKXWGcTgRrg/xFxcbZddcNWasl0fVT1
neyhnUlxDr9mNf1Eg4wZW4W1ponAJobNsl3PQJ2yNbVVgSLEG/p3C0s8bJ0bU7D5LSb0Lxa9XdcQ
vLSNFp7+gY1jMlzHmWAj6NDyeVbFCkw0T8gOLDCVN+koAqmgE//Ac9NydcZigoSb3eX3QSpGTP/Q
K6a0joJDQD8UX28K/A8tztpeO01XsmrVvtW59XMPJbpy7IMCnThFoViq6cxwrrGobGEnsP8YgKBj
/EB9HdYQOsdCSIJopNxBzN1/CXm1sPTyYd3u15rijFPOyHdpvwTpZB8fdUQaKQcOD9C8KTcjijEx
mFE9qfvLclCS0bMoU9G6icbTyFnW1CIPHonGs8sfUrE55y4O4eVweU1YzTPMpA6sV2JFm5zeukoQ
MCtOTfO9gArJ7fvO8x+W9ep17HW4b1wH9I46fHDOqcd9MRNN81Ar8UoIlNw/zveymG3bh1mICRFC
2NTD/4xHBwb0dW5On6HddnjGW7/i+2fYzP4BbixfqDuv4IzxRyjGyaH4hxq+kxjv1WutRD1tiF8t
QLDcHlvnJRZNVRitTMnrqho7BsjT9So3KWVHCbPt64ACJMjGDPlh/xhbJR0fmdkqe+oMNAiy7YDF
8PKHo0Bp5QvPhr5VsvPF0KupD3xr914oyFSvNz+jzDO1AKKOqQddybQmQIsMykeuItTPdK13JQ0J
dPBAk6NzIDv5lYRW9GsTzo2ULAJCjrUinUWOvSIp7vY8d0QoQbJAHa2Ar6B2qjpAFZTVFi64k5m8
7hraI0o4AKZSZOin5fHXSaiiMD1uv/t2Vn+Dw/INsvpVj4a2r6NBfSEcIsz7QlFgTjXjtOT2zysx
sdw9ts8wunmh2HwB3SkishaeggfdXr2bEM9DOUhZ7/YKI/nF/2V7UuwuPagRBjK2Tn5Tbuym9PBk
1ANrKMuPGqnPWZKvIdqEeaGM0dj9r444/zuZdRr29dRlgk/FNYKFXfRp0SBwlua7IvyjyxQMvSee
Ojwdwd8ncP2/GqOF7iKmcV63AgWAdvMG1IPlk3qhYbXh4glp6ERYsodXIWR2nTTODkdZpTPj3Mmu
5vABE8GqA9q0/eEWiX1G83uq0qiPivSIzE6/8AagLVVu0lp4WVf9lNGkv8gAQqFKmMZjV5Y2jySM
ckHNg0tTA0A+kN2hW7sPCdQ7Dd6bjyXxZ1hDPi8zcCwiI7RKu/s4UPsR4TClx+JmSLwGFOasBwIE
xAx7fFeIGCRPkfSrTueS3l7FoSVORiM5fOB2GODd6yv9MjIY9M66RahULo/nBRWHNJo/QFgX2N27
KZG49SrdfFd90OWhppBJkecZVMlroAKgjDyoHtdPoOnB5rcAWBUGc2AIfs0UFZebUc1R9SPA0ZwU
HykYYsQGW+2ODcJkU30TGikVl7WP24a8rcyaNP3zu6SuIkOyZd7lH/Ic/rWw+JN2tzvIF31XAwMw
v29RDRggDcGmlYwg0C/n+nzltZFg4e+ue+xjdEKMee+GbfnpyLNZkQUoKFIxKWXdA6YE11kFUZeA
oDvqnOotf7idmx1iKcX/OlafjZBP5nGLnbMlJik4N3jvXhqp2MaTpzgG4CT2EIPGH+BUjcKGNKJo
h7A+VEa0PhPSmBilx0m2widchrVHwNNGhvkmbiHIqlg6a2NHunD4UgrsecI4zKIsYM07h9BIMPZe
14LLO4FmGBEPXthQjFDSf1Rj7EWQoiYRECpkgd0wXXOTa6rZM2I6EgKx8EuFeOANZqJ0gG4g9R/1
GA0sE1j9TPGqdr5nElaRkORlC5OpH3kfn+4u77NpugDS7mrCuYS4xKBPItATU5FahJlE816c7ysI
1zs4gGjiihV9wx8AjdAR7EYj/MKQTS1yob7lz2fUl2HVua2SRFGzGACIQe8PCfCWwHFbPUfdEiYh
RjJ2z2h+GgqMbAqzU1H3914PoOCzZsfIpOUrxXFcg3k4sUuqOQ+i+BDg8VsTC7CtHPO2Xeg+pQzx
hgM/zN+pZMpVdaMn/YXGEKiK+8+m9Mp72YXOotEBJrB2IQJFwx8C6eCZf2D79Vk4Xk7KSiTHUfN+
DEjgM5DwZCnOcDdz/Ug4r8Sv9XuNtUgT24q63kXDSZ/iIeqy09r7jKRafY7VR2bi3zN7emLEVDwT
bjMS67mbtMpBUj6JNzum4P5X28EjeFrQLi5wCJYYBoKG1citIBypRp2/HqkV6egzoaFd4IOPijoV
MDJbZ0t6uX32WL+XhawqivWxb428RUsAYtOo8Z/s/tYEgTyRoDSEsdZesEiAIsFIftiE/p+FfnK8
V0Daknsi/oNwCdTK74JgZBal/JyUfUCVcqtD1c123nVGVaJfIXW/t5cIOKYxA33tbrjTsIsJUxLR
aC72ai1CCHmM8pHYUUEWGDNZ5v7sSVNWIPSVLUUa+Py+LPCeDZvwTgx2FW2Y9AMX3/YW2fT1WWk6
O2DWeTZnyDkjxRc7OCaegYDZqQacyQaNYCkwvmR4Oyanm5R24kWD0ok/Cq97qIh3WYpnNkbQef+k
lqsV4smwAFhDx2F8XUk9XcJihJOGWT9uuzvKKgCqagoU3vzgPJP+MDufjbKDRuJ5xwAYpQPw1OdK
I1l7UaDUfc1s1S3KZdEFrUHIEmGn0WUstKufG7OvCWoj8LpzLeNHTk3N7gIraHrzIBtIYotpMYHI
EGTWCsWmEPwevTyfezSD+k4Xcmp8zr+kUR84ImqEotge68lTw2Hsvg1JCLGK5rIEf221tGgXoee1
vr7XYeQZ4GIt5mNngGJb3o2b//T77OYgLmOuKGBCTpSh0cbVs8ycLDf1WcCREc7PuZmHRrHOURay
1F7XC8nnHpCkDOhsYWQn08iNG5zDOrVae6ggveLVmf5iIc1bhNscN+A1qhowzx5HROLfEs5wwxfO
ftJS9evBD21NiSK8wusDA09otRjV6k537odqpqVqiFyp8GDoVxTWK+97Mp6jZYx2PyHMbyu+Pb9N
JdCyxc5xXiEBIn0KAAvhb6cP3wcMSsGaetdQyXluYhXSGikR8lZem8zFfWmWGXXjTqXTyWCtHJV7
sU9luocqXJxvPqnuWx8jGFhuZv03oPsrWKBY4scoPgGlOm6f3GrudAPqXVoPJVHAv3zC9OA0PA7k
mpmPHXGkOrp3U/cDBJIebZOooWW/YeBkdEkgGh/3nzZhYbK1XZjdKQ0R4Aas40C01iYW0AMpcSD2
TQ4uJUoqvJAD2630P75t18CqHgc/u3xIFcWVWOrV0sRkx4iUUTllCCIOZmi+wd1/bUvIUMiecLMJ
TUshS/MX6EpsRN428ezmZVSz/WKZFnVSjGfVjmZiQrt51Eoh+7DhXYX3KumSzPRC325PPCu0fINH
BYUNJ1/5bVP2F9ej+scP/OvHgoCyTuIGJxu3Wq9T7r/kX6K4rCb5r/zENVCHwzs8Fmn8/orSkPv6
eoJTj51FrSpCUOtV/f/jvWm/+P0pXcRdUnTdLGnUJxLup5LyxdEwTz30uaRIRu3LsIvKIrHubnmh
P6o83RmMeu9aB8Tf4IpBtEX1zqrk6l8I+kXHnfnf3JDH3R8XdiFkEJoAlxz5iv/Yr3LhhH+w5WI5
coHFt/Q/MLC/MooOEd/9qMmup7YfdG8ro8p3aQ1Gqie525G2LUDhxvPrm+GQAdrW8ZkGSS+yE/f8
YMZzrrlQKH4hHVYvthv78dvMpYhpTcy/b/njV3BKLurc70mAgWqpSM6gnGeFAIbW2BZ5oV/sIneA
qp8vW5RgtO9xahBYmEKC5lPHGE/Z4LiNsDpf9ioRZKCfl24uImuJkmtXf5cmAEZ7lKGvksF7O22j
LL4zUDJUNcswoLcfAiTjfb+FysY81Izxiwaoa+21aPGF3rFi/gWC3dkMDis79ongbik+jxzMAVPv
7M4ve3RIzxdY6Y5gVlvj1gQrcSKYpblY++O0NufN7yEcO0e1PG3TYUP2Fe61CM0zL5Dpff5dhs9F
OE05+r14Bw15mEAgvj81fvG7UTE5x6j9q6hYu+98UTnQkHu+7KejizEUxIaK0jNqSVjfUvfLdqQz
8LpfDpYmCAr6HPtQNRLWjaldnz/RH9areSyQLv4zOZxFykO244vDXGLEk0yPy7L725T21X6in7BD
MxEu4lDI1pS97McnmnADNZHlcPNP2Pa0bN1skLtnAiAZQFBz0M7W8qAow5/kWEWE6Xn3bg82rXTq
i2RMfPcv4rgM6zD5j2aQ37vfln6e6Y1KAdg+Plua4OF2EPxSKieJAsdipi/1sLzSJtdVzYPL6MQb
irLmrH21qWOXQ5Y/hrT15i1onFEq2C8/slgzxcviItk4Jc8W+Hby4+HqJzq2wH52kqVQXkks9Zo+
VJ7rHCxrGJGgsK+catzLm8ItIkzx/K5V+AarlKkTfHwfflyGIQ7WqLIj8huBtXUjj3RvvKlMrXoR
8BcPv5zhN0rq9UR86LI81NFQPFdjHH02JI2+fHLm8Ji4VXPML76hCpU+i4EJ9gKDG97V70ybN6b7
FtPEa4HwLamBmWq140EoyM7uQFhhhIn6BHeuQjur8N9b22NqGOZt7UnS+0UEeXnYkMT+YP7BiVag
mzfxvrpVUln+8ZwS9WuSwK+OZi6MhsiYhwvSmkqIoQltHripICbabhFKKpDTeLIKouAd0+1Qbkay
BRheve9OuXcQac0LYlIqYzM/Qs8JGMJ92xPSkipHRwmBzjJRUFSlS1af/VXZTORAfORRY8XteN5z
OpbSvOd5ibFGVgoSQ/Tp5GIOH69JtJ0I9rL4mQaCDWCmbPlfDG/bRJr1lkAhU/JuS8puRZ4rSBpN
pQcAuFnnEyhrsFUPtyMrqFhBfupZ8JuTNmKLyzbt8rqG+mG9YCpIEM+URwf1IXwJVrtgNzUhoiD/
CdJHxjCDzUcx7HRav5nL9EM9FJcLpPrZ3YX3aTYd/kTkvy+6V78lVKLiFJmWd5Y2eT7ReZyA6rCU
jvfKnxfPAPYahXpplUgw2jozdzqn1Y31n1aYK+Fc/0N7t7KMfTzBN8h11SveNrRD9ckqC/PTA/Di
gRM8mue1Q47CFxpPp7obNInUDBTzR9eOmT/o4N4TnkK/Bu3IwCNnhq3/bPTvcqdQNMADSVY0xe27
QThBRtXbk2BEB0WHUhlMFihQlFkAZn9RS+mPg7LUo84pQIDyHBF3OHdCgKEpD8X5zIoQxztvkxmT
WzXQRmgHp6THv7Yaz4Zzjy7dvK1mMBMvKcT0xImpbUJMAp7V9Ax2JpQckf+vuB937B5LzXtcAr+G
GJFugpuQH1PrfRn3CpOkyAXPzhoqAC2dS/PUPQFcTZRYgqqs3Lt8m3lYEUlm3d3xMYXlTXYJ4JNY
EQ5kTiCdZ7J8hgqgiEXUbMuheRtlBjXCzZzJa+qkpYLsxn/ZlBNbuOhKibrMVktndCUdnayxTX8D
LG1mVOVdGNXiRfMYLFLs0wda2wWkzTiGwdiazUZyXQdwL36co5EQJeFsXikCvSSbMlvrafbJetbj
F7xmmvjIQ/MT4SCXkdeToldy76jwxkcUjJW+7e215+khSrD8iO4mcE3fUWH7K8Le+JB6Kvjc5/o3
ZrY+WR0N+nr/t5ZCF2UluKbXVoM2P5Dc2cs6ba5801O002zelhwxPPawvTRtbok/o02zMfcRvDwA
9w0kPQdk/e32eR4CrS+sbbS01nMI+JdzCG5IieThDA99D2f5k3R6gRGPKJdg1DbIqtGH2jaZhAy9
GjgyM37aqmbbmlILleqeBRbH/Ss03f/LsmLIWpbSfKkBxfN6yNcsfvcjli9TTyJJrpX/cPfeF0wM
SXjiX4iMD38blc1MrkyazJQNl0D7yG5Y3Xnv5Qj5/lFho2cv3P9gPMTYp7rhOn2Z4yhN/Cn1eCYB
nXFuYR0rl4b5t3+xVzgXAtIbkAVeV9UR68S0bbSP/aKDTGASzyMe2wzP/JHYw5kTm4rtRdpYTjAj
MFG1aPCzAqN0JqODZZitgpQFsIfk1DRUDN2GMPuCkp3vU625ban8vBfWSbjKvDoCk974nYW+EAO3
jKuJhv8aGXmt1P1QNnHExnhOk/fRo7zicBP2ynmOlUwdDxkrmu+Uuny1etTGeMw3nCISCD5mLXo4
sjbk4Jq4fH4z6s5s+yEvTkdulQ+00wRodUXK+6Ck6zZGS24B3SfBhjooa5ZcSIq8RVV/YPtCCrIP
5XHfqVgvlJZDCWyVfjzgKC1rZJyx0ma6vmPVsLzvUTiRVzS0WeB2/4ahD36QJNrT8QdKkoLSH8sF
x9dhqVkApxnGPAvuIQOalVtmaS+0EihcWIlDWjIBUiG2tCQ1WATPqgcfMufHEEK3Es/cAwkjcWom
ubVyYD5gTjxmLq05qoakoKBW3h3dvgSPppEFkwLX3FyqzRoB0ipIwdtk3h+8WvqXve77HiCC6daC
e4h9IMJKHgtVj3+9wZSyvrY7Mp4IK+yvv7Y2tiQMjSRn6C3TByIZSrYz9/6ZkpDQkgN0mIuP5pcj
wIXkNHvLl9DpzD0QR54lbNO6MMsWwqyYxYkWexkUbZ3Kr1aN5DeSoDE85qrU8BA0I9y6qDcf3kkW
LWK7CfCAYjsSSbZJ3xJmRxBGok/KETzpKbo4/3ECS9ONcJOxRuZ8HpSndjfW7hQ3qvVa7pFJv1/M
7QMtN9It/Dkw6RWCF9BdT6m6zFf32Mx6QQY5FDdvKnCqPRFUgaGfN3gcfIP2oHyPEpDSpd4sdOSC
0GO9+LhmNMG6d6PByM0d/9fIUI1caa9xiXiZSw9zTfV52LYWQklhyGoTPEeNO1u3YFJKpYGn8AJG
7myN+upGZfeUBKsLJO+Kc/oqQTFhyXsGDqAM8jc7PZTOdvV14YvuYCPMpXDbD8Q8MRXydOFPJ80m
iqCim/4zWCSTwy1YFj3tPviWM6eWQKchybRDS9Y36gbMgVLRFCxzP+gEN8NAacFFLiVfPn4DM4bP
RH73C0r394QqZZU3ebmqGJurJHVDQwPVX2eB3aWOaXN2wXJ33F1j0Z+S6zpXmPFBaGQHw8KzFF4r
/Q8Xa7EEVd2qnaVWSlB5L5jzwz3yr+Gs9oHYt/ie/w9zB7cua+TBFpmxR+6Rm7g/Fkh2VwznFM7A
tz+VwWjAedR/FEmnPEwFZnIUY4zezfS9SYYI6SvvTQP4W+uxf7XLHAGzAtro+DlCwMCSdq9JVmdY
wDFf1y4+Cx79WlRywdeeTAfgStCtj+aaZlW95hF8/HYYBcDSpXEPoDURbuul/D5doQYwCXNTpDbj
k+geeQd1UzGw6DoQpAluiN0SIe1sbpbpYtHSGmlBtqSUej6etV0IzSHwz2LhjeTwh8HRAgUM4LmQ
Y049IYL74bNGn+k7/evG9RXtADJ1YiDsXEAfzEjyGGdlf7j4v4O2ySqeSoQsHIcSLJcyrHZ7MMr9
zWgXluNRicr87dixXW1ITw3L4iLtxItqLuerqpBuaBZU+Ktrh21kyaCjLS1YD9roJPSP5K6FCXQo
MA72Bk+xqyrjblphgGk2ZDNsG8DTj5iZT0Z8jnErKCWVVnAZe6xO46UgJ5lKa/8OHQkJrTbvxzl/
+jdVkZRT2j8nSVozhZhstkGuxMVFOSdOl/W2KeFEiTUlF34ue0GrmRh2pMEgRJzcOBF7TbTzTWQJ
Fhsn3GvBdAkL7qvEhuWR5EnqpLEY8b5aHd2+1HTJs2OCx/PEdXtFN2MYJXoseAa98oymCneDtUg6
O7RkFZq/RJMHBcBsoL0+k06ujYx3hHRamkc5bQ6jBEcY7uzXW+3h3MoFuHKlLY7hfuTyO4XfaZ/9
6Eyrp3G3hJlOif5UteCNzdgvLifqCtKghedwVsik51BByWEIbVyAkGJtk3AaKlJ4D5XvGFCxuYvZ
Ogaru0EwQV2egBQjLxmscONDWt3WnGUSfxGYR1/Kb7uFna67zBPcymPS0YQP4dp43mEHlmw1fgPZ
wf/dXJP5hrSB4/MTsPZ9QZaj0RuEc9G/QZ/OjM1yGGFnQ/leLNupdP54zCQJTiXwImZ5/KaZ+1Pw
DFEJF4N7Xtavhaex4vT19K8TK9J6MgO7uK9nW+nxf9Z2z9K99rPQ0yqjwE96pEpToKwp7BdCKSOk
tMYF3PS+y6BhyxlnN8nv6eM0h7LjVZsbg+Bi0IEGBiQBO24g3NHnx1KesH8fe5PjrGAFa9FYli/G
2HYkuUQ9hUzE09UNOp0H3ZigwZ1/r3iBNhrNgXpeq3uvR5brssb1tXya7cKnF2IJV7DcYnH8A3vp
2h3qPjGFAth+ZKhSRtPLZb2uhaX2CDNYihKZ0fu5yOlGNmKTSXaRlyHFz6QH6WZkkJTh4wwbxuYk
7V3R+S/E4k21JaoneWGM4M9/hG0zTRCAZ/SUcH7tFu7B5tLfHCsuP0vw3SX4S/VfzVrVX2/yw6IO
0wdp65IRXXZexHDufXJ6u8vjgneabCT1Xr5H4UaG9YK7UiiWwxRDg0A+PwJTjnISPzPpSVnnoiYt
4fVB6qz+TXm/e2k+O3ZLT3fX5Jgy41wJa4Bmbh6GCQyqnAZlCHhOX+hlWV9Aro40Lp2mLmcBuWJs
GG/aqiHb7SsWPoj9syBp1OXBBaDbR/qKgJRAQs6N6LnYCIxdmShXBk7J1H/Un5nP5r4S3rBQtP4C
A8MntWC3hJN6PRrRE1LBjIYqSjUDCxeDM/7pThNCENLCuy6wr3c8S9R8tTkp9vsr6mw7XHMy3S2A
wprSkPcoY1/83rJsKrBp/9akQ9HDtLLKmAmZGh8SB+M/DGvr1L7cZBQdmKeVY9RO9IBplKxjgDQJ
8+noBPR2NiVFD0AmCrBJuX/0y4IPMLQX5X94+01hQLXCC3h5A/YcXWe0UCZKDU/PgGNRY8HniMNY
YvrNlPMy5R8RLz7QPV1ZiK7038kUVTYVbo2vthBvPApNm+6PLtCce195/4EvLZrBcOj7DuF2QYpX
WER5OU0uP6nbXSn2CeBAEcZhElBpdzVPVZQ4sX2WlAIvhokNvA7T9CLVXyhMNHdqEM5lz1YXye7t
dAm/LdgWd7pCA909EoXJkg12v817ipsIOxRfNVq+sGVWzNEKxfnVqtXEAJoGkSmCcWna6A37MDUK
qOmTqDCgOGGu6VbGkHTyDAVkJBQLsGCyPAzIjkfCVqJM3dMLqAAIW9cs5I4i0vDAP/7gNddfBqjT
ff1QwRbNMunwi44i5sbuk2k4JM+jCvmTTfHVoUXOTxcHs0O6Ql6GYW+a3VuUn2I2LbxxMqyTuuOY
ZFPOyH8PHE13LuPMssQYs0tb+m8OiXzoaXzzyDGipgKKMO0YNwnBH0HJcZT6y4fia5HmS0pQtvOV
h0ClYPCQ1zIFwZyk7kXb5Qy9pdpFVfymRMXJOY61ImiYWDln6mkXqy+7GmrTjsqa+GQiLqVWuO28
shnLxPK4OH01mh9OEHbsD9lGlOenhEGsYDeSY0Rbzt5TQJK6hX0pCdsbfpfutAJ4gmzRNENLOKr9
/4xx53huX9vj/Lb+w6UKkkNOBcYwi6UWhEYnf6nT36TfV008mrj2JL4EImRwtyDx0a/ftUML4p7m
6RMPh7TwbDG3eIrX8K2wiqSom2hwTX5S7o6OACCA/RiZw3D2DYc2+VnBizWEs/G5DrB6codyb7IY
k6JJpGg2nTMff+bJ3RxgfSvnvzyRJNLSnNdB3G1kshtXrGMkLNq/Pd8nT2U5FijNmEly2b2BG632
zQtgRhZ7Pbn97fRl0pQSc6wrXwYFTozq0HSmaI3WKAYDqdershOxzDTHvMCRivcoaK6UY1O2/dAN
hEj9rZRIPjA9gjQ0gev5w2tn6OKQXzikdI8x1lbAkGdCT5i8ahTQBqW7pgZzJ8PQbR8SE7Fu2Hjb
ySCc4bsAo9zxWUrpNbHBr4BMP1VPQ2wSjCNO9r3+vWyYJq1bC2+XrFqRtwrQqerb6yQyn5Y9n5GG
FtLWsRl49WdFw72q305CY7ZJVlcZfR3Y/pwkJRJBEmv5jCUP6rtNEY4zp/Q9f1c3QLEQi4lm/3YA
Xdt00A+ea6olN/NCjxz6nCHNzZPcr070X1Z34zfLUSKxwa8tlam59eBAo0wRu+PAFJhJXL4kRLmc
QJrddcCVioj+QGHySCiDo8bgj0VZhAh5VPXvmAk34Wex0ymkZFUz2cV2Y25iyCEA2bnbXWKHxdi1
V9zm1J38kQG/YE65SMxPR+eucD/gNaoOYzR9ib3KQ5meD4VKWJ+jLwRgHMVJIh5kA2A18IbRFttI
hL+s3uKkLZNU8yGYS17txhnDcXSezBy5qkngC/fP7WFl6QAQeri1o6O99LTjPCKMlMYWt7IbDEle
zPJFkH7VPI3Ku0br/DIJnLN5OZz3RMSxY/hL2dqsSZr3J4JLe8jrfUfUQ6bofAVuomc52gqQOFCH
hbJPzupIQJYS/ES3T80IZikaiv/Ev4bx0hk5kkIiidGhltKio+vUuetcu7SyT3LzcbRFFUCJCOP6
UAkEjxgHoowibkxxvZC3IdtkNIJRx/Hd4CTECK3fIphQ+KW2lbgBgJ02G695XYWtR0QSI7LNs+G3
1wTxAspkYsHHiOjBgH4ukKX3cgyJbSrl6ch/Ik1OCqIyxVl1jPB57y0XbptRPnElNsJYt/j9RPFa
1uM9skYoZ5dlNXGVoi8FavGE+tuRIa0RyBNrz64YTV/xUj1kMR2tISO9UndVZJqwgKMpyeRAEqWD
LWSCmBh/SumRwnap8b8c7zjHRMJ4qmwHd5W7rSJ1YQz4NMVDp9gQwDCE3ba2vs2q9Val0BUF53Va
jhgy+noZd4CHQZBauXfuTJMR3m5mIappnuTnhB5F8OayH6Yl3xJKQPAFhytq6RBJaMdhesmlWGuk
IeBGMl4VQEOTbzihCVckwY9K70vMtyfUhZEXrFrCXUEm58pupPwUhFGrhoF1vv8w1cdnLpUsD+2z
ZOCwP7rW+3QuWYQWxd7x1ma2SYck9g312thK1GgTDz+jLPUbI7+H6Exfg2waZ524A/8fAWbnsKzF
uuL67C5nG99LE/40aIyn/LeXGLy1/P0afY3R/Ujg/3e1BKGz77xZob7RPjtNhxjJSdTfjKsvABfc
eC5WVHqV6Aa/LS6ADMfYrsEnljx5eFlXtb8y9RCwfyfBfinI12QQbyhkNoeAi31uDWuD1vlETrcJ
TQA2ESK7/dvpcJgw0WED4Yj9fDPF6gogC3fl6EBuV2ttyhQJpnv4xgQRXvGtL+lJllmoCSdiM4cA
hm1j+pjtdyxlHnnRFywucQJtoE1MRXXx8uEIFlGmPgMj9L9Q9IX2wnCs9d3Wxa1FXS14PC4BKCCw
OK2ugIFDGeBwkZYR8u/rxYMyxjavprUKbX32d2WuYq1W2fLoa2U/6Y7owr1/dEFTROhlfrv3+3V7
/Qg87UixnpFD0xIzEwk/VC6K+YbUsuQP649Q14A7h91RdHSt4ZxouOXKn6ccl13GZ/r68nu1VYaB
T5X2ZvQCgc8/ovH28PfunOGWiSknJRjEobOOnIIiEdohS4DNcYlGA/jTJDwOoMPaaUcVZAb+4vwa
9s5z+GjqWTE0ykZ3MPNhgUFIUBOBkY+6iwJfYPEhUrL7FMB7dMNZMwKqxCebSyASs42UaGY764dE
t076dmTCYkwwVK63rL41Ot3uA6OMYGhfNpvdxQysX98MOYj1jMUn3EnMXRxFxeg4viOcoB6LcxC1
lt7hD5WuaICDzjcq9dlNkUCowxBJfQhWj90yEUs4faRjEsOFiaoqGrfbwFDDeeL6B+9Ralyfrjlc
1d5yL0M0CyaDzbuptfMSJh1diPnReaKxdYvb9EeULerLvMyojs6agBBk+Pt5aoXl0A7YWIHoPLdF
cIohHwCAITrOWszjHcoycyv01FRFlIBSiTjEKO2pYBTpVbXXRrsDfBfYT31IuwerYs0JFKrryVPy
DneJApelj18aDm1r1Id36qcbwapORKA4pZKWSZhZFGo8P5U6kInYwlkb6ka7CEvLQhSSWzxJcno2
LM0LM0+TGWd6zNfs+VjZHHBy1ESYkbnstEUEoz/IMWnF2K7tIefZaU5M5e3O6YiovnIxJ5wvDUa3
aiw/x7JN+JQVOSNF51dkiiLWL0hGozDUfC/M+LFo9I6JPiQ3NyJc0RVNpWP1cAy6tX1jx81m9Sx1
ugQeKkGnXc53V4v+U1fvI5Fej1vpI8uj6PrVLBLC2uRVZD7+LKP4CKQOjGoZKV7JJxqOvEvSfS/7
Rop5l4dQFJ3us+PPPyZpt35rd6SAmdFJY4xxBYHXSO8Ps7dW6mqmhDFcMV+6tF1XCoVhdcqzYYX1
j0gD+fC6/UkwtJB0nB+PwnuX2xabZu/o4UxSyGskREDFqt4FE5oknlYuejRqHC2OIj5B+yaSU5Pl
gCcF28TiwPEkmp3mQgQxaosQzJxvN1cFgXJ+ibqzWgQcDrJIBSirzlBPK+RN/KstSEt62Ym6p/Px
1WutK+p7fjtXTTEvCshOLf/BTkLFLisafQF77OTJSs9z9mhUh8CRD64G1KCXA9LCdcwy4iZydIxN
/JWNVTpaGmy54X46DFt9UitUvFbJe2CQ6gkNqi/vp8zvIyF/x/piR5FpIeOL6Ymyavu8LsVH/yay
NTrj/f/LGPXi9GyuReNLMxh3FZ7MfZxkRMaT7u0tXmK1zel8QIY+859nHgL4+s79MhpylgC1AllL
mX28zf/Dww47FcANgBJ95aB2gD4S3MnNlc3TZ/GCdKDIAjY7IGGdMVOO9AkGs8Yjclznjw7cn5TC
4f4e1Z45ESEkscjQ/8D6VCb9XQ09XN0DnhnlrUmR3xnS5j14+GXIWlTt0oDGZv8R/9FUhP/MiaM9
8sQ4nhHi1lBhOgH3OlhBm3wHa8iDLPLzFYsaWOdyd/TFjflJZzLfkm+o6mRpZT0scOSkoLT98QQF
a1U8JDEnoREl9zc4LXUFo3kbT+TcQ2AA0mXXbnx0bZR+xOauAF73YKbowPtXtDn1SO+nTi1SAtXV
P7Qy8g0FOxMhhdxG8q0/vvSMnNVBh4q6joQHN2vO7vMFgbZQgLDa1cpazQAKcRuU+fICsRU3aBx7
YSITPyqFRlVpuGBoOf620l5HQd4L3GIqaz6gZd3Avq+XT7LxEostICemIuyr0KTsYVenuEbcmDDE
fZBTuQ6r3NxlAlDet7HqcRn7jWXcdguWccz5iinNX4+6uyEiXVii0P2SXC3YbeFz1pTqyAu6enWj
oigYpmElH94mDiZ5QdcdSyTP7ZD/NGxIwCJsRTNKEbUV4V/Ay88f2ryVA5QklxsErHk49q2rS9Lt
317GA8DY5ayWgScL0lQXHILUgahYqGZYxuW/7wnhrXI/z6oKetH2HTr6LZQJgQGXHHXFNTq8rUPe
9qj5GTYaXnoWD7XG46IGCXCkq06PB/4vpSFDZLOotGaqAyzMGRifmFv98nQLzug4T1Xaf0ohu5r2
ING8aNJtiCETQj7Mb7uVX1Vm+X4Y/KjQcx4M1dk3srRhA9d4I5ZAkafRXZRmFwGYC9SYFyN0QtUy
EVzJn/MT93RMRRDtXk+vclHNSjPuLfnY1xIhSoEkB0B779S/muOYQCp4Zn8odA9PaIRf3fzm4isS
cpA8Q6bFgIUifAWSj+BWibBc3AfK2KWROA07qQwSWhzSNcZ8i0UIK+sIh/bSjTHKWlCcOU179xqp
zo9YrAKHO9SiZYRkcT9/YxCgV+4RARDHZKr5Zo8itof+BTZ+SSstzdBvHjvT2emW7q8/R1FHQYDI
3WqM5X8LH2vWttuZNENHL6MWOJwNAfmv30Gftmkn2eERcJuDzHSWvUxdYKjpO4dgWTCLUh9BzBog
vakbD1KcDqTjkuUa2jJIaTSB/BXtF++++Xpeq7qNskV7DHYF+OBoPhQy8AcIg/QgIwEiI7DrNj6v
0DoJV6KNFossR9QEX9J2BZuc7fqfj9boks1lr+X1HnkYfmb7AGNCEH66aJKkwfN5SCf6NdusFPaK
qWIahiX/Aguq+TBwcDJr+K2ShP4QCtRVvRx/FsTEf31kFz+YNVyvAfY4Gopcmca5cmqjsndEO7Bk
muPByeqnBss7b7PEhjgmhVQQ5NV28l3cYcc7KBq0l5UwAeJ8LpO0wfNH03iEuyqaXUQF06R64Dv0
B4Oce6BKYi8Od5YybzZuf/BOgHCwrvrlng/BKxCqyikImI9jS/gw6K9ROjZSbwjri/bt8jiP5EFu
LbZ/teq6ipdSN3ip7yMOvzkLSzDPx3lmJDcOsDizCaLEW+mfelp+dhTHC7GxQLctBMAT8yiAG0+j
0X8ClyfwIwCrZK6sbY4TlADpMDEi70QL7sqFfnxLzvxQORQbQP4p5fXE/a6bzP7pEfv8kE3pORWY
YSnzraY/xRk21QTnnOw5gilKlv1+oEu6m6jxO5TNPF/UvVTxPzEADliR79aIxtlyoGsLQssbdSjF
MY9PyUWJS0Al2OEn+uOuiTCNe/I7c8FiyFQTdqFZLQe6YmgMznaIvLw9GswMD4IW6PJ003jPw27O
1C+b0n3Puxi9f01qvKifbYt8eeW0G1K2xTPwlDre4YELxWFSpMtzfYR8VJessjiwxYs6VNRh9rRA
n1b0sdzo25R5iB8U5i18tSAybsackQU5Vdl41CpiVGUrb3KbmTunfZiFlx06fMQPZL3RAYIhEbCt
RgbmYRQsVrtFZDhIQLJhb3rD/PZwmtNQ8UoZX44BQjlq4LS221rB8RSuK1TJhHJjhv/rmeqDX9bZ
yaRFA2omoMjYgRvsNhMDAJVqOuNcrVF/bayb9cU6dBdXRKYf8tK7uYHNE/tB/+fTe8bCIZr3OGys
K0f0/I0kVhCl5ji0LKXjWpCrWpw3F+a2npoglSSWqc9vPxnwWuwEnpi1HUfB/0SdTk1AGnWUWZgD
C2HfbtMXFL2ZBj+fR8wi/wVSBPw0eb3uWMKBVQY1QodSQQ5m71DLXC8hKU4P4WAb/9hpLs5lGoEl
tI5VkC9buVunEcjvFAgdSnHCv8NZO6YD7dzK74O0l5RQSXwx3LdlvyGQcAwfKzDK9eU3QYYdS6Lv
7tiLI5QaQYwJds/bfgZ5orWKR2J1KFp/LPH5M2cT4g3wrQCpfdj6wm1RCZ/7hvtMDJ0k46WPeOVC
sOWEzj60ikkSUjsJ5Ha2PQOX5Q4SZ8vHzzwBCqC8GbKpC82WH6yNXw7lXkLnZ1rIFMsNT1h9U6WX
7bRqnV5gFQhtuMBDa6h7m8Z7eHiP5zS7DnLgbP4e/hBx5KsVxuPGS+u/Ha5XUrseExy6+ZQxPoVf
nPRojTQBX55nDcI8HoB8GW/0uCJzC1tg0O95En1w6a5CC9n2EtAAI/N8Co8cnfmXIiEzgDsAPamf
ppWlnHnAXNOTbuVQId4AlKTFVKHK/NSL3uWFJ5DUHB+2+3No5l9LaeuDhAdMKx9bz+KNpDTIx/ki
Qr8wx5FvhD6hW+JCk1dzS56YckGNnVf5ZEiPCie4rqHiWTgk08ImbGzrA12IbRr7BS1z1F9uCQDT
w2UYOtC2RYkt337cYhiFjDScLvy2TSzNr9klWyj/VC9ZVISSWbV1uEYCK4e5aPh8THBH+COy/F3j
QRW6n6On8wAKFLj/ak4PhSR1ZbPSjRBdSbE2UtHsolH35Pau1YQjTAd2rmkYUVCSvURD+aqn3JOP
kGlp2Iqtjq5AV7/DhPVs7hiU7WXwS+moZ+bQSzc7ai2zGDeztXS7ZA7w8dytxrSpT6T7rcUlVIu2
qMzFY/lxO5xXzyDtVsFxrpmo7I6PaVSHnsytg6wTTGfPzXNB7MeKRg0tIMPLO4ZjaUoYNKrQpVlu
tCi+7MT1YzFFJEeVgXYRukSbyJw114rOGUDLyrEXH/lv3KmDA6bt3g6bD8TwLjYHgocL+CSuqKsT
X+ykgZhfRl62fFep51O3kDs4gbP0EhwDalhNx6J/RpPXMp5gmn3P6UEA0RZnZrVtoREtzRa+BTde
dwY55JHWKUaTTWNd/fAfYLXPyYDAbRuZP/TiRTTPWa9xsek7gjavlHv/FyOgw6oqu6AnVc5kO2yF
iT8/ZrpDORnkR6gUNmJ/cNZRiJA4Cfhdp18qa3axDnDSmrqonc3vUBY8edp4qo30qneCXHePZdCf
w4HcjHsP0hCLz7DxFR3rJKeqFn8FXq//7Injqf44xNhwyK5MZ2u+YP0OZNxhEhR4eFORxDUnnGQ7
+191fii+7GiGR99ze7lpKlF1twfbpVV/hE6cEwszY176YiwURCGpT8mQQHPJ0j0E8Upu7OpRICFz
a178Mp2ZjRlVYwAGY6QqLoQjFGw7EbZsz5AlHzAD9YXVHOqUR50L8dFDWTDSxztmuGLUnJl2ejp/
QRsYbeAS3hKdKAfjYoSdemKBmxApyd7qKXxXixGyjs90foyN3CW3PoP/KSjn4p+kNYfBPUNiICcn
FK5HvbJgxxEdUGELNi5l+T/VLUe1VoRrd2p/BfFLN6AzH/JlOMoL2GXAk1mv4aq+ty12GUaB0rN0
bVwWrKHY/LhVoioPFpSBRP79kG3DyKF0fvaGiDaD1yW+FLH/NW/qMhhI4dBqnCgTBSyRjpPEgS7j
tiUaTtc9AScI4kMtvwoypvenFGaz1PerJJex7kplyoh7etUhv7W6kl5mr7dS7Ig3FVWFlYo3bqxq
9+Ee/ytndgr5mGsdxQoX8a2TNTHLwZCPbX2NvImOKdwuI4P4P+BoA/jphYmay6mwIVOgMX8A7bmE
pCIWGJewckUrh5k6/5izjMPJqzz1e+PF7gNHwJpr7IRYxvtt2Yzwx1Oe5r6i/PxvLpqQF/OiISHq
B0mi3EMe1kmN0YTii1ddJHSFqAOW7vNAPak7Pjwf2vDXRMNK4+20t7H8BGRWgS4JJyX4Mq/RHt/N
U7FlQhhGsiCYDiF/AvgDOw7ND14Y+Drgb88H5dHYg9QNEzXdPU8SW85aagYLcAKPtYY6cUKToCSR
tnMn/ynZSwrnBnyWxRcHAdgc546ZdgDoyb0HY3MbdlwmmD1BWY8hajyJihfIxaJ6q1tx8CBYe+DS
iJZZV5ch4To5Ndfm2mLB9GWcZeTpfOqKJ5ZqFojrzOhh8XxWQHueWI5h0cy1esjbj2RHl27P31oO
0akQCTG5jCgru3dfW56jUW3G9umTLSM1O6oOJOS1V/ZSk54CQw85KXePFsKqq+epYLxEael7D9DX
YNmdlnWMwitz6e0Mvl/Om/bCaZaGOgwmW/VQq+Pkm0VReiAmIhuySW9JfR1n5fugmGs8oIWFHgd4
u+QCrdDKKEThAdbVExLUtdbvi3Yaoss+sn5ouS9UMGpBjdJ0gPczZzzyh9inbGTe5cqxruVzS3kX
o1086Ytlyvh+GUc/vzUA40V8rMsyayYVUP4r8ofKsOLeYRALAgGinw4wsG8IUBmRjaUzF1bgPcuW
ZZ6iMZhckUMpcRzEhNk6kQb2xJRJPOxNh2Lh7RYyHn6xPa+vyL3VnHtnb8xnw1OPpCc7e3n2YlVj
+TrzPET+Q6x3eJWW0vi0lOod/b0wv/bqOML2+2sPIHVyfQtUHllSgaSSTpOOZcCuwFPOc/uwUi6q
xDYPnzKs6BAmqx+QlkwTFVErYn36H0mSbLdXzCR93siKWNMJdhpDgaG7ElhRAQLkF3Zi/Bqao+KC
VIVkaXldsE1qkfBM3iOiX1nLD+4ZawdRpg7nLCcqEyVHmEqkupCgNKXWBJkIuAkI4V3RjsBqgqmw
xzIqhmgx8UZSx7SE7emZSaG7bOby8BpTfn9w33v2qUn8SX4HM+QTJ58GyzQKReNA9DT8f5cBWSgu
HZXLRNo/63IwCU8gpxzuCcMzVYKneYbGn594VqYSHWBpSjj/SbXrCo3TJKPNRewbZUIjmjXZfpP1
bEzQwuPo/Ubj8KGdHyjD0C0CHv+XnqJGDNwUiAupWoFbX+4flmSer1xqmdT93X4daQTGDvTUPCZW
VwarIj9q6ZYDUL8QOj+JetuwN05r+tg45XyshWvPHsvJGjLal5SJI1ycsxcXTzej5zLVhXiiCxck
s6A5ORkqRJFk2JeXRqpveOs1Ac9pdjSaffxF7yJ7iyp6nPqSJhU8qiCXKTjoK3ZqQNmkY8VA51bD
DpykiiEGS8Qb0Ll+JeObDbYAcw5pS/JnfN1ltrnL264dSklIW7ai7lfQynCHY8KE8iAORV7vvzXe
7pUxU41gvwtiQ4NcLDalafpIBpCNUh4HwYTKtnlorqvMxRvt/qLqjio1vbBoYendz4RfOKB5SOSv
GnaYP312wty+zdmiScLF3UJ47t7PrbHg8ZCDuLMrC8DZgqYLLL+f+A4sy9Lvcb1QMsSrrafcz3iC
wh6U5drWtj3W0WWljHzg1hNY6R+pQ2AX+U6ZWm1+1z3dQMIiu3NNjOmENXYQXyQTXMtbbCpmnoy2
46DqrhRWMZ2xL1hQNRDZ674zULgSJqLvolr8hRonX2d+WZ7E5zOnh6l2WJw6rnQcO9RULCWBpDXq
okpwisUfY/zsAIhVuhDaY9N5I5nasK9h/XubgwRZkdjrcYKNTdQTj0WeR5d69e3ni/JMXrYZNeoL
DALmgQvbRifGt7OMvVOHePqzddyAJIF6AZsKTl1DU2mnqMdKaLSTqgXRliHxQhD2CwWeVQI65pAp
8gyyvFc0OitYTv4jKUFcua+2deIeLN6j4yaKDIZ1PnVRoxumhRJvIFlUmKwPXablcmwNRaSxfmSe
Cs98dJHq3EjZCvBukaEZrUhHw0YvDN9swXUWUd6BQgm2cwY+eJBDHkySGBq1+tCc4jrpLQwMdtjr
8q6plvOurVmvNFOa47kMgWUOTJZdsB+Q1zEN74e4i/h4EMorZI/2vcdNUGjGc1rBcdAau/eZXuLJ
SdYDLVK1yPCLx7V19uHbI30i5tThyvLlB1K+Kusouc8KSozhHGPJLawl5MoxDEN3W0qkONcvCQMR
3vaQYDJhFNkAWyLOPH7Lxbd2X6wYXTnw2sAiSmkX6hMf8+Kf09ugBE3GpUbFUeH34+uMe+g/pVGx
2MvMpHcN3tXAkvPzeyIElsa8n49GzP5tbe0FBFIjFGbI41cXifIRNGHdwpcygWIflKFwf127hEGw
2uMtyPoyWT13qdGr5Y7XkJ5CeICtzN+aYaP2Sq/Qo0t04dIJf6W+GfpXj1d0Whkotd3wuwduJMBr
fzj6hdva++1EXG7Upg0H4+WZtdWHAlJNJ5xT1sd5IYKZG2Jm7mqWzmsTBmOFH+M/BoaStCr6wuGz
Wnvm/L8aHAykrAkunMFE88OGKOIxQJwhiMQZ1fb4DLk1AdVRedXCY/6yQp5l4p2aBFNjdsGaW1BG
w8MfMHGMz+yIBSQKcB2UFMMycREaNeJiHCf2UmdbpEDWvA7c6FzV/jYM/CZ05AGS+WDTAwFRJSCp
ZDqv4E2Il5lApfTTKg7FhHBgOmOU+rpm5n+CYnU9YEx708Q5Cmq+lkuBXVRhW24zg+j66XQxpepT
4IDLw2duc4kmPqxOUOti+TJhCm+NXXv9Hh6dQ/J+W1ZAzdmJhQOBb/Iig0K0pyiWZSoU7u1z5J4w
iCSG0uAsEkRJzNItcJrd5/QEu9DwBqTomBkDvy/OkvRG/+iybLTtLbeWDnlH4dF/SY78y6l3yJcZ
QWslyRLEGVpfg/v/zfRybGmcm9fqPSO2aXiZDQVOLdJoUe2mrVaTCv/QxGe5XPcyXZHt9U0FundR
JoEQe74d51oUmup8sBh7gpWSrf0sqUEH9c5EhwfFxNi8LDOrjy3Kwp1049DTp3flmia9KOIsm1Fa
zMLmgK6i6aJKnd8bg2f2Lwd0+Q8kGojg1HT2M8zBVUclQD0YUWCTor/ZA4IStvTMAuR25+8DR1nz
XPjLM3+5NI91a64kOqrK6T7gxVsx/jbfsfkSG9gFuTb/Mf50/h8BDSBRByNhoa8dJg9WJHhXaXWC
I3oWg5+Bnnp92xSerm1Pxn2Y68B2hmIhSCbJMes3fDKPDNUXI4oeQmUApLRMpqzMmBqzei3zYYRg
rfgldRmjLOw7gJYk3me9xwNx78xuJB1xwIXvRd3XC1YiiXfzzk0gCjRzUd4fPpoq7TJV5tG7/kQo
g9BC8/MG3bNQpq/ErU1AGH7VLMWV8T67HfpiazfEamjcptMYNrwY+A3rtZEFuP0+xh7+aj7Emm9x
Bxt+bR9l6hiU7KDWUk6Ei8rf7m6c/Y3+jUth4XhKP1yNx055U4y4nl+NL9t+nJyqW1dceAQ0R23y
H7KuqNmpD4974dXmO/50Fzn0DPwp04xoWz0D7VU1bNF9iPMikUZn99yWyJzk3+j6UdhsFgtTUrdW
d/aFWjtoTWfkEmNMoPrZGw0xim9khyjaAb3GDFG7ynr9Qa9mLxKjRK++NxdJGfPRDZ+1qTxTzQ46
+diot2knxGSOOIM8GijCPLD3fQC5OF+zldK1WGw8mTxDZB1a5MwaIFsIuEVOMWzuXK2HyBFkC5e4
10LQtcjXKJ4v6FHKtgbZ7b663vvpvq9YcgGk/7fGrO6ArU0ZIAYEoLUkJYif3OkqLpjN5LAwmyw7
KnOKuWwnvKiv2SdMUqAGPNeU8MJIAOD1sAjYVxke1B16j5mi5ICCRd0Tsx9PSLa/vw1crD40x5f+
MzQIAS8MwP/srIKeqS3vuV4iQjAug+chb3wjoNsa6Xus20awivA4RGhEsuJuPUmoDIDBrFTReSCf
Doig0G9pzFOwcXft55PiNRSTOZf8k/9QnhaNDDzW0IpFB2O1zoS5CeTlW+yvzbnWVl5JWvoVv9Rc
MnZhzdQS4XpTjEa9jBLsq29uyiwQPMjiRQ+mWO2frXHrMKVjnrgKlkVnfOggaxDdfOSsFhvSCYPB
yov3rC1nCDxnXpt2BFIX7e5pf1WD/hDkNrGWZSyOEmFD02NSIXkI5b7Fu7xh3Cb5TAEMunQ6pLyc
OBbB0cRBMa8NNQ+tvC5t0yacju//OeXERVYlRj8Y4CA0HA68TU8r22TF4q3QTz0r2ZBqDVuTHGS1
Bu7oZKTaVXDM/eRdnmj4RMVzz7snmdtolV7GDzr7Q7an85ba51EXgK97sL34PORfmt1qKbh5pald
QDdCGyL0ZitDAmscPaOWxo17DU19BeMfE4SJGbOPgMJQKvOyI3V0HJBKRYBCy0ySJR9iFHKm1pDg
DP4YPh9k2KRiKv9lziAxrXZOHH26ms4BxNPXG0yWe4Ft5KI61RYqPx3dVQjholanRY4IeNRi7N27
uK79V8d7MXq9Z5qCgJmPtyU8XtbmUuFqanhOIXa7+Vo/U2RAT7yATOXmVUFgSnpdND6jMixFMLdv
ez1xcz02shN10x952yt2WsnPp2VPxywzI8i6b7Ya4h/Jr+zJajrlo2Z3i5LmFtGqZtpXaWlQmQx1
jcxv61R1EbIzRte7jqrBbALu4XndxQHVsfH+Yk822ywbcAgZ79feaKdjVq0HPup1x7of2RQDwmn3
8X09nKpBOIeD4ACTgErIrCMlpT5+gzQi9smg2I+Yb8SB4OBNWuuC3SEKEuK7vhN7Y7BjhKRdJU/V
F2dPomVnk/sytGDwk54kTurdQeuXac05uznafr4EmuCabDNt/AExjV4rr17iFS9/CvCZ5T272Svo
g1a98UtbHPfIe0XTX0s37aYuYwW+aW8pYTJYNgWTPyXWtEv5P3dR2CN3zfQN5jXkVqBsGRexd4HF
Ko672z+Go/qHjtJpci8UbJ9vCbpZX0/nN1aaFD2BhI6tetsIySgxl2G0N5dUrnyFMI5A0qrCXpCT
MWJuCcA/aLzwpyZmrHUXB96L965/WOZzyiUJ700N10SATNh+1Refk5ogVi8VKUvCKGYKbvOxjSeq
91G6L3LiNfVv8McXE54nR4yQxEUkZETz04s5hHOlZoColJjEoFgqQjkakzbjf7vKHQalZ+kvQX0a
Zxepz0OUdK6pwBPlAjC4H3UpLx+G65tMQfUr/u54uezrstxR1bWi7FHT4ZFlmujLDOKma9lQKlYh
0EmhuhLjbLAMXrFMhyQdHW2W4KoPIiJKGnGst9Z/pstCflXg+vBgFaute7QOjULVmrxX/rBL60zv
RWup8RXdFKUIfgotc4ews0X8jAeEJyTQ9bqIzNnKNaFczMyIwy1yPCYPhsjERSqONPtfeGJKmYHE
zRnK4Gqe4Vn2zRZq2mmCpifiA0y7TtDzHGtGh41UGDntlwZNJP86mXAcpAsaUdhP2fs8icq7b4dY
PmLcjbEAbvHXOkhL0cLVbUe1mhqlnnr+qUr26gQZ6QvS8pCEYug0cVuGPW4COOMnL2E9fld7Bz4P
LSgs1XqxKbzfuKMw/vwjF6fAb+DCIKcVCduJSIv67LrMqAbrp08tHonnnoo9hWQaLjl4wnwck1M7
znBcAbUz2mHNbQcvtE7jasgoSDQtFLFXOs42vR/vHMJhaZ4k/1GhhdH7cwRwy+QDR1E5n46VOuIi
v6r7QrnEiFrCqOiv5Um1XRGKm3ntMys1x3U0xzrzTUbHIg7OoCpvBH2hTUV9LIGKcp5vUNla0Bcd
Tk38bhLXmQHU2tURKFFkwD/WBdGF0oT7ffl+BNJmQ3KoHkn6W4nKljrS25xG7G+wNb5MbbFqXwnu
WYDdMt0/mCn39izTadT+mCkzsP5GV5++oHHbwXYmb+iRE/YowgdBC8OC+bT6U/kJpI8L9fKCjGVx
gFtTIsbC0b+7CsUUOU1YAX9HiTMr7DsM6I1yA+JORk7jtjprCxtbwhzPA7PYqHfNG4rGf9fW3EhJ
tRqN1DeRW4uzp9s9gQT/wR/RZybE7TZydu5uFZBMeVRpbeMFjP1N+jG5dBGMQnluSSLlIWNA/9uL
XVhBviMxhYOVdwyI0x5ZQnDD0FQ7bKhTK0JkKJlCJqWTwRG/HXju57JIAONyubbYCb3WnWfEFKfk
loX9BzgDyunrwjxYF6KeYRUlmVnsjw3QmoaS7RdPT8kQlbaCixH1D0gzkm64f14EFw/w0aY4wk6f
qtREJYZzBySqp46i7YR4SDJvimFnAOk8KRLA3ChsR2Lm6xg3FX1dCKRSbwoasRomgYwxMs3Nr09u
Af202ApAXedLhMDrE688mVSlnTT5oypJlRE8RUDfFoFkL6qWNfkMoSYkqXPaNSW8J088qqw0Jbas
92EQt5KBXWHecfm5FcaeaTCoOPFIRKnv6A5aGKX4Os8Rxb5S9ltSU44ozeG+gETWVC5QG+l83JLb
2jRokTRvgSWJa4lfU5VHroTctNtqt9YKL/SgjINZpQRcpwfZDYWPIbx3La5DX4ykcQiDUNJsl93K
WSASDpC9cCe5mOQBdtZOBoeKPVZYmfp5s6Hp31zDw5jS8c4c7oyzn7BW7QQkBWW5BrtylbujEsrB
rgxYX7s0+/0kNLO6MAlZb7XpDgs/WN9mkxYb1khTj6eT6ZA21MnHPl4+DvX1s1QSYgt5L5ocbrun
SxQS7WwQqrR0QuT0CcaUyguNdz6z48HhE+gMP1/rj20yp6Z38AaP31R67pQWPVn48kwzBUADLY8m
vbViN6UN2xJ9UmK/a1TC4iJEI9UpTUHQKFKmgS8L64a2ukbTU4JmJPbeV5k9YGAsil57b1FSgbPf
UH52oU73uDT2ppt9H/TYZ3Z944i4UpdGDVRuMOz0hMY2OvYWbAwBvsMmulQ9iGZBlWAnuTj21rwX
Jslbjc9UBZ8NIF160Z+dyuR+PQCj3xoX4tGvY6SrOrn4COVLUJKq5vPMQ+vy6I/BQclB6DiNyTZw
sYhasmI4LUVpVjPOG+365I1Vlb3nRh57GEztnsmrTqHnuIJJUCQELpwKS+3Mea4C0eKQSYZAWuoE
jxKT4PJqHj9m16l1VPz9CWdN+mSdKv399iYEte/lhpdSkqCmOJmD2OVPa3/lPiK3oR0Qk9SIVedQ
/lkzPF+S0EBgpaoyzLMBv9nndYmAroMbe01cIjG56ittVgu6A5d8eGk2OKMlURwcHzmUGPoTPmgo
h8zKz70lTlOd4dElc42DBCC4GcOIIfLgxLjvz+k3OgjNrHKu/g0qd8G5P4PqA3/+JbvPphOMX9jx
VEnkS0WIh7PjXhTWa1+EdtVyj3VfSOPgqVhKbc7Z0AqjluxD6jbBqkHjBgr+k46JceOSqfiB0yFg
Hxxekv3qB7CSIepaFdEWYllKVEVduGR2A8rl5F8sUeHwAmOuiQpCWg/8uTupKSvbUq6sF/lfPMrk
qR1s/CzQIxkH8VKCZo79/o2Dt7XixxdnOLYqVyf++S9k5PlaRFiMxgiwqY6SBUoE0pDtc1i3LKnG
olJ1BjlIDgKIZ3EoonNGnaL/YbffrNC20fjPcq0uvWlLgE5eMoSsh5hsnyVnqTvB6N4nJHvr/ZgJ
QZzK3zmKQcTnXbstz89IJ0ry49VN1RaCA+IxBo2NM7+11EPpoqby79Kcd0cejVGdJId9AhKt5ZDb
6GQm8V8jBuhEiC+h7KR9gutHZFN59PUlgaRUCfp0ZKMTTLfxl+gu7BZWTly2jlcFuBpZpWHMT9br
Dbwu9tM338rZ859+0ejynHbZ0lfQZmCuUOAdyjIUrazvv2uwx62Bt/m+mMOQtXfFn1MVdlIUu5Um
v0ft0Fk+KU3DUJyrpKKlIYtRCPmCiYQs2rvdQLReWAcGCEgOPwiIX4R84/inKtMrhVZAiFrjY2NZ
rBU7gU7O9OYbwPUkcRiyYVrs950UuGBAhr/GKI122B8densSzrtGrgtOWFbE1CFsS1ORuCF2deCw
Dx1a/mYOjch3u6EBki7uXHMXC6B997p/jbhRkCfF8oEMrJaUXnh6uMGFWkkgezT7VSUmpEbH/TUK
8HiHvemMiHrqnN3JN+1W5c9veMXEJUO6XQrYRNhPn5TBopSqJgS0Fn9DXvLryOA69YOmay3qC0ew
w38WvlAjEySf49L3I0U22EAYkx2ES0iVtPcTwd7t+x7q/viaCpxHQwomvhVApqZIhCP/eus6w8U9
iO8g6H5j14pQBsbXAzcGfixCgkTFw57skSIzYSuYqW1DU8i1evkxzpEBWbllbwgCxRkYvSgK/7rk
Qvo/zOnRxwfmQbx7Zaq9ZIy6Cdg7AgkFPDMk8c2Yl8pb+zTuKilLzzQJ+FB7kUVK89xIGlT6j84j
zo11rCDeKYspUDCrnFIu6qRjZ5FNoLuidfpWH0O1rpIoz/DtQoj5JmB1dd4AmJ1DLF2wUsfYJgP6
OlAoH1O6QxgzwT70vlW+cQ086L+wcxDNN9MI5s4TDHAiN6BtpBx+qntjw9x/Lo4TajZU+Ec9Q2J7
OJJmrfa7Gs5/Doza4Kve47dwApbwb8+0ZSxx+FZWHEYjtNBcOItupzj/LJ1n40OgwdmhCs56Ua8o
kZogdFFs96VkqL+49EPsORN2dqvx8D9kA+5BjwfF1fkHcEN+NYhd/D+56gDHSI/up2EyqxAy0lIh
o+9KiP0Kpw5CwJDYO6fRilVUIByUSwKKs9wDog8DEqJ0SwUxJIbu0eT10M70Mzpmy2hAtVX86TDL
J62OCcZ+xj0BipDl4f0cuugny77DuDBk0dYNsTqsHabYZ3VMIFJUTsGEmsC5C6HahtHPTox3gtA8
8unNcq0xnp/fklR3kRw+b5Vq6xfIoRHNilBD6MmCITMIaiH/x23D1fE9wUFf4g11Y+tj0t4FKgCN
CleK3Wj3ANstLVR24s3qOgER/AkCEtA63BvaS1+GPIJG/0F+0g/Y9Lt1uTw0rbNokBFSBLigSoKc
WscClUha8eRGI0qJq0dC2h8RBWHPfj8PTsXik3Py2Sz5s0RQGo9xSjtLmWEgYI0RjbhyDNjgAg0M
pTOy5k36i+vBXg0wI8mXVjFCMe4GvsMQffnxhBXfALp5/WakXBMwb8KMnanuxBuuDwSBUbPH37cg
Qaqb0vA42n2DgRGuTzFpcpjEWOL/UseHrIRCkn4f9yWHXlmsyoy5LFhUfcTosR1Wsel7Qh5KiatN
W5UPY/sV91OvHCuB/68n8dqVIMC0XwHMvDN3K0xmDwI9usP3QHqtuyvUKbDzW7m7nZnPJfVn3c4A
Gqg8/YvsC3KJ3O2DURGu445/WLTPxV6TY3PVxwOyPpZmr3PpNXteOH+kcq4Oi9s5CpY5o6K39mgo
f88VIs3PyIM8kJ2gcUsLSfgUS6uYykFC+xP6+uwTct87yd9JVKJyWhtMgSQ0W1FSGX8MuiNKtAz5
QLiR5LGdncYfl7Upr9cFy0frJxusPLNPJlzJEjMZBfZBURjx0/FRTLTwPpCZD/JLWma4QPhbGQrf
6rB5jXA3K+mQTA3P2AJzLQ5VJvAioZ0SljxVwwFMQFVYF2m3HoZ/BJnIQmzc9KuqasYEd63eReRH
49VmPuvjnQWSJsuFsVwU70KeSf96JjNLUGix7bnK1J0kTaYUbif0r0urPSP38f9iCAleJl9gReWu
BrDW1zq29hXeVwjZal4WTmF3RTLZdFBWiQuI6CV0Beq523/385G2Clx6zP2GWf7YmEN4md+RWFSr
IJoEAOcg9wGfQ/PfIrnDVBZ8qXpDOJJHmixsXSnjHT29OfycWsHpJ9a+RVD2HqGujgxiU+rnFiLJ
Ybdg/qblwwd9OZ7XRxWWBa5Z8OQnRWsfgnTA8BP+i8ey/gpEd+qOzPqN15e5JU/qj9zaSqa+1X5u
bs1bCyMBdkmy2SEsnxGVUCmj107oTKSh/hZ2VdxAT7vDNIiDJidQ9+Jyc5KNefslcF2s8SemH7Me
5UxuCkeWDoiKeTaTy2xQkQ3raX467PTlp5RcyfIAN4iAcpqYKYGgxX4lSPuznz5+4IG9AzgzXTJB
YCV1UZ9C5OjIau2AYeih2AspDnKJxl7Pvg+5nAj8oR4c+OlxKpLnc0EcCaHTzsjyoJA+eEXyU0ZN
qi+6L3tuu5V97xDo6O9T+MfqlxgFQ7MNtX3HGPwsVp3b2PMsWUNNwT0R59mra+kSexq8qWWv/ygR
IRQGsZG0E06IX77WpaHNLOH2aDkAvanU1A5Reu6EDzOWvRUcp4QqaFDaRBEsaZMRXpXLZ3V33Avs
79YCWVb0mB2ZNmJowjUsxkGTnQ4Hkch1v1MKO/fQ9BslwRTCrlbSebXafk6YhiLxRDIf/+BM8NIQ
BroYG9DSuXkeyo6EsI1QvFlOPUZ7pIfv8cH7jGno8qggBnvHYbiTRwYx7eRPIw8a8B+cejYqF5au
jgWtF/pRTmsEItn6onY8ilLjHx2hRbdeUe/J2Oz+UVTSEdE6nabQq0CgIIw7XcY1jg4RwhiXxEex
uEGyUHMtCRVia3DUU9ctofO3d7L6XMD/vgCmdmdFZ2FhfzjGrMhwig0Nc39N41J3LP8ep+FExkVj
jELSq1tUvN0Kx23CBG50qAqhdWW4/ykZo0rhG0eW5BTFjfA5Wnz4atPFN1qoXmwmY52O9Avw99xP
/yDoL9QxzWgl9ZFE8Rbjkq71boAmrqxv3VRuK95CEurpT6ocfkdjrjgLQC9zCWvtKhZ56athXsAY
+I3Z+NCKqcLYRZIvR8wjsdv4wB3o/rDzhNOF9KBSY1Lpb7nkrN4Rtvtu2rsP5SDWMs6F6rBTgjTB
bL+lz/myCYR5j0Uugd3DqL3po7mexkV40hXfX1f00m4bC16Ci3l+AnNA/Z3JlGa0dyGmurjT7Aoi
ZJuoeNmC9U9AGd00IYmFvTj7mANldyypBb2l18PINBFQrMv5WReyk9akaBOjf7N27M0wqHJHydlm
TvSVuzvA090c+R87ZmBar1OFQVLkClxaB9ZJ5q3D0KvyFMxr+Y1L0gLEj3LVDl5PjYaYohArdtFa
Zbf2q07gJiNxsTY4pKrPzGahXaqK/d2HPST3ItkHaTkbdZCNfdNuaDRw4YYMeHxAySOY4r/oPZDG
Qlr4Tjw55fxOPY3GvWfmfgSzctrxI3CA4/75hQGx2Xk9+gczTWP4wSRAgRmNP9ltzEGwLM/qC2/P
JWb4hwm+E8UL6HJvDxlVjg6+ysDcYulWKa/FxtG7VypnvN6OP+gBwfT39dySfHADwMv+HbzEw+tT
gU8Dzs/3fHBXIja8LxftPUJYjJCPCucTknPSdXgoXK5NCUOXXdd5XSIYy3L75r5N+uVuuyr14YxI
6JDU2pqSaEqJsXGyND5JY0SGfr1zATNM+ETVnRfYCA1ZaD/Nh8FwZUS8/Se+yE3BpjQsfVPOMaZI
jBv7JGouB2M1EfIWjnRVAo27bQfl7jlNnFGp2Eyge+VmNcpfsw1MnbjdTFyN+w0MSh6D988m1oHN
Mp4AOt4pyEDaYTmoh4Pfy1fbL1vkmRDjEZffCzhv9kDK3qUBdxZifWU69NLdccNLtqFocBgnSymM
Wh8N5ipo66FqB0xRjwxNcThfEgRIhsVFs7L6ric5RXmXGkMOIz1RPBeNSzr3egM94F3PBSQvJca0
UhgdYuP31hK2zhHpHLCNDKlKy06Ob4I5rjjsstTiIHMms5dX/9Xk9sBWp9XzzLMZrVEpLoy663gl
yq+DS1G0SE0/XqOGzSwJmvi41K1cBHLB4i6fjvZnDuf+BZwc+k5zmXq0FlPsJGS6fyn00zdudFpC
oU5GpG19Bkpi/vPGZ5pa0G+DJU7z1a9Rh+DPvIKS0wh1lExsraFE5XfTo2Nl+gP6H1Ry6ayEQId6
5m8kZxrsuGBySZAoLn3jNSkxGUwL0f875TkP4GqGjjC0N6qtW4thDnuQnpMX6U5eDxaDT3K7S8rY
5c8czppOdQjtWdlleNmmzeccifs75PmDBZzQY6pHFPNjd6BR8HaXpdo/KaMWSYWf/RqLfkxbUFWg
Ttt5BhmZVt3AACnRWjyxUzX2vSQipGDbP+JLeMKu3/NVNNCRONbOiRHX9t5MV2o9P60Fm+KNQTUu
zEU1UIRTzXdefKoN7sN/6iCgVaTkv4fRdi7kYLqZPt9Vt9Na+YGjjbjIASF/sQgC4W5sLRdJI7ej
W2TMPaupB8kE9Hh7YA4vFjFq74Us6lTOpVo3V/d0E1Vi9+q97i6YMGdg0AuyCLRv3j3DzRr4WsfP
XlbZ5/1CmtfdlYC0K0KshVDrFuARHoTJe7/Z9oSrLL3Uc3EKmp581yTAU/DSKEJrXslnFSLp4hCp
BzbnVk+A+6xLJ/UWPTbHN9TFzAOhgHe2NxlfzDVYNPg3F92iAsXPDnQyahBs0DVI0hNuchBAYq29
s5xwIoVdZvg3Two3EgCS7gBG7+9YIWftSO0b3Wy8NbpswRoKKNXHL5252thLjNbDQsjf+X5bCeHN
FctB+VCEQyt/Xku1AGK+neF0WYnCCDAe/OBM/7EaA2i3DBuQeROsUyVirBwSn9G/8cZainEL/1Hq
I55zvdxskkx5lmQlpIHuwCj1SAxovEgg2i+2uExEwZYPVMX5IEtvS9W0e5kanpbA4CyHXbnlRUAf
rV+Cm+uS9xLHBuvzgwWsThLxs2znV2YEc519BC9wPxMCk8o4VDMx0UWa/eN5d8Wj43qMru6RMJ/V
xULTJuqYe6LQnZehrjZtr0GXzNvwTSUJhujtRsamxocY5lD9Y1PBD0Y6PP1dVRZ548Hxx95ODbM9
kZ7mpDLd+J84pf8fEzzQYrer1GjdM4+VUM27MKAkUFCZnorPysJ+LHvNbb2MGG0gwDMla3fCyZVb
/z+Y0twY2uc9FvFZyDWZ7xj+qPiUOCaoK4AZbgVJO5PCMmXbBcLl08Uu8VF3Vh6Y5wyEoBWRT90a
y3xPxqgR55UidjJrPyi7RU+S61iQta1wP7IyOoFvMM3NV7z6a+wDyN1d3n6WIfcEaixG1k8Vx0+0
F9nlGFWcab4NEIkE+X915YCr/YjOB2oSh4k89YtC25bromgy6So5mzmPR2qrVrNo8aeq+FEvDRNE
IlDLMwzB4FJdVCLucFcLlzZ0g2I66VTZy18iZWqQ3a3xaQxq83aVfD908BJaCqxDkPeqTSEdyq/E
Cs0JdLAmcjwrigzcJxIXu6D3PA8QrUtatq7B6lRzD0UDz3GSdtdrM9xslqN5ZWcg9ATAcQd6kc/H
H5j/CAk32dvR4+NEVPlo8m+vC953+fShV57ArxEb4HeRlQ3Ixax/fuKwWsfa5Csqzo5SozHasMQZ
Gd62dbWwnlh6patMu8g25+4I8QiihkKNCiQ+NilMKKSVp+17CuLAYwq6PkhOtc3O+JsqMw2MEbLE
U4GI4QxTs7TG7dPKSqLrn1QhlgAEGx2o6c5pgigB3r1mL8AJpD5awzdv3YuXOfmOpkpxc4EqbJvZ
YLZHfS6STOfjFGfg688qiU0qjfp1a9Mc3E92VfokmaleojcyC26HzB5fe+I2Zx0b+Sb4FRqF225p
dbg4H41ENmojGKW65E5ik4N1kbq+MeTh3Y2Bv8pirkYc9g1QVaN6L4o4HcP4APcOx5ljRJO8Dzho
bkd0A0FxK4n9ZKqK1AQufeIVod+jYBduRm5kEvhayzHw3OQayYINYaKAJ4GPR48LH89cqV0lHHpI
ugchAu0awQpgFxDmguWAn9r9AI1nHqEbAdquZxGm7RPLHDwhpjp7nLeNqQRw8lm+1szIgRkMx9p4
iOGE4nnl6sNa6gXwEgt1YUbuKw5pbkycuK3J2ODUpOWrjIHP6xbjh8p74B6+pbVwFKBnWCuaqN3X
jxB/6x//eQ1eAtmckIRnO6ypbkChQt6asactVE4AKffjribL8aJa9ccCG5oLjF4gT7/Pl68eAcNB
T68ExvT/6YyAiR7SdaCKkcouYfajM7B7Kd2DOGqQKN4OaeST2Vl6m6Y27R7t2f9LuBWm8Wmlw9c6
hRXHJtVaO3J7Q6nEwJmScbDG/ApbZpuukpaNagcxXkJyYOCu0TEaiOYz3TdhM13f4/Q+yJsMkYv9
JabMqP1aqitMy2HPNLCLSh/jB4sWAQHyus5GpYvhZm8IN+SEey6+9DVutZokmZ3rf/ZuDc26bHlz
tlNL6eSQateaqYPgvPbxaLQNVPYD/jaf64bANaXPCOR6NlpGnz5Sw/Nz2h69eaC0ldLZugDvCMJG
Ut7py9l41au0SZi2W8YwWqWlghxxXyuspxvIS4DdHEv0QsfCX1Df90Fao7B+FO+C32rvTwzTrE1x
LbACf9YIX4tTszGrSnJfvf69NOhkh4AEl52yB6Mzi77127tVlQN4hN/THkPDvQivTcDOvZltd8kS
yHeI6kQrswmirpzyhqHaUs+wHBj8Wn18ZpNjDFtIAE3Gjo3clnK0tNcb3D7K4Oq3gjjPYsOJK+mT
FP4/xCtDH6A1gMqUY/3bAMbZZqPBTQqqedl5WgABTd0OMu2zODIMv64Cqt1LTd2SjUNMKulNcypM
mRT1qbqtT2PNvSQ1A5jWclLy/KDUbt/trxTZf1eQ+3gOYDSycO1suh/+UEdYY1VQNEv2RwVVE8px
Y/D+BswYqIGL6qzEet6NnfOnxnUT8spvk8rP/+mICpr+G+cBSc8XgdinrYTrknTJa5XCkAM6cUuT
/Fvrjyx7l8iJDTwi5/bSlLJcoFCwdUag1WSuqY8svGoxh03f5kkm1gC+JnAqovAN8N+gBlbT7Vvz
J0CkwW8ZN5VnzSoJ0+00Q+x2m+EWwMAb1oK9a7erU+SYkLMzV6sSjbxsQ6Krv42bOyc8QqoEZVH/
qbuVJsezFbL5VxggEvUnIrzySBBw8svV6zV/phkD0DsKyLWMo92NJE0rmi+Ican32KRb5+jq7GUC
uH9ZEoAjRA747tzPRwabgP+levdneiXmHN91KS3Dph3QdYdBWrkGcEU1Hr63XSjpua3jcABvBWNW
TlNx4B8Hpc8V7JQA8T8Cmmb60slnlB7vLoI8fffb7YszpGgtrKaY7WPIp20d3Carn1W79qvqK6GH
RLx/rScnMaNYrs3sNsXe58h4mVLcppD78myGXFdDLQsSDRNYEQ2XAFfCB+Tvq0QhVrgmOvaKIqkh
K0QJCLNvn7YMycWIFToW5qsf6soNjgKy9ChgC8hrLu33CiKXwPgH6hHNciqiMeJmuhM0nfJYxqoY
eNxksS8h1D6YYEPPZGOVx9vTlZyP3v9iTApAYiIiIYMS34WkfZGgYxFBbwKiklYuy2sZbv2+2CH2
I+ONzaB3RJPiBNg/KwcIYJoqrR6uVd861I++StA3jfNqMrOf6aq+JYmhE9jyEv4dxyN3C3uPQe3F
MKdJVEq0SiS9VQ2xXSQxiqqmKaHsHjdrIW/uvaswWiqbufEbr+1FqPnbHWw1fGHYMweIqtFzR2Ov
MtcE8OVRiBZ7UcQwReF8CWse74SIP/Nm+NEPOz7K7LV9Xf4K72WQxlwLIspTsUPNbPN+vLQub4q1
znq+BEUQKV2JVSgMiJ7hrqqddagcDk2UrvpOrNX+PQTUVgPRPQPO01oju4aZdHEJZo4j29+YFdPf
cTvfFgq2O0P/4EWXqsLjSx5xQVmX/nTeKUpXHHZmwdhttUuignAKK2GR2TkqPWCxdfEyYDyM7eDV
NnzQN6m5w9tuScfnjHCSPVJ+gc1pLrJ6B2Ad2/bxLT0KFxLhLOy7hHe/E8NbVOUTvcujUuhBq500
KYFwdcgylwIoAKr4hxta5+x9KyQLR9MCervnvZTScS2JkdxVNGxu6cgvkPx5QcQYMoqm4lL/7lhK
eCUu6fx57WbR/AWFBwqnD72sTm1+AKJlhjo+eHYzktX9ndRjyfgAQ2f5UUg9S7ouOG0G38rN4uwf
f9PfU6too0EAsijuwS1XfTN5PvBhDpqTn5k2Au2h7KpBmEJjsRDICst4zxtTrEPYIU14gvlL3XfX
7oM3PX0FeXMyHrAsVlt6fySkMnM65IH5BhqjirA9LM2Fv11bV7b0AkR4CuaS906wtrNsJ6uQE8yF
M2eo6t3O4gAaHWXGf+2UHY+xp2mFnvwULyNYt8PTyW90wwBo3Cuvwb59WZeYnyaWDhh+PWvdT6GF
ld43RuUocDH2xDriDLIECOhRtdb/SieQv6ivGus5F+1Lw8a7GFMDN3TsSOvbqTPJNXa3ysUYaTro
TobzKiKJgkc6rmriV4Ra/xiRpliPw7tEoaEkVnDzQDPiz6oCgwyW61CBw8c6jZ0da/WqbJHQjZk1
mIYamPF9wopdglUi7CCVkL6F8EWYBrJ7XB81pyDRJToai162u5kwFt+oE58cbnToYRNtpDiuy6yJ
cPatUnwdNHkf4oAueuSxxaAB+HXG116JAfH8cP2JhQp9sAZgpb55DctsDGEFkgx7NmKjTvmdotPg
BVnjQAXJDNShd28EHds2A+wxBC5Bv7sr3nGghknNitOAR66TOEtcEqRq61pdWfbUoaYyzhdha5yF
j6QSnNwu1BgytS10MVjHTfuxe2KwaZaM+4MR5a7EpHL94vQfeI42r9noWsZig0n9drQFnbl4nI4Y
29UqkVZ0OqCJK0f2+DeiomTqNHIpvYDNw87EnlOM3RSasx1ZwBQl/zdBMJ9F/Q/KaPjFRnYKSCL5
4dS8/e/DE0WCeHACNqQGCfz0Aa/uTMZRKUL9X3T0SeD4iOrTWnDubboLcEx8yqyfqPeCQRMtS/Wm
3HttEC3p3d8bUmuzoYwIAzk7111qI81CnHf/kvF6Smr3tpVmNpWqwRYgU6vuPsqqVYslZlE4u2VX
4Q38ezBB2eP1p8VGo06BIjrjg/rQdu0Q+jINZ6awA+59mrArcaOuCxMzuxFCuoVggDiLVZumuPQt
hzEr6LTAzjXNIXT4JvhWLfLYAuDF/NN6VEiTZSnlPCazlPotcv1h54ao+A1ZdfVTnDp0pA1YPmkB
12jfqR7ekv9bz+irvac47IUG4kcd7td7iVJWsTSMOCKR72aGQxEUxdwUXZYU/Bog1wn2eQe88zd+
kwpGkgEfbKOWA9n3WqcIuB0pzSWW2fh044+7sSoF1Nwfd5iE6spbOewNerFpc8/l6J7e/2HqUDlc
bpbeo2zgosYD9suKeGYEkfvWgEvwuRsoQNBoNsrgFpFGSlGzIBrd/gsZme3su1lMbOGHGDB5P8da
NVu64QVqIgTGKsEM1UgA6SXEy8pdyoAv8E0z0Wh3NLYKCCUteA6c7qwn1m3E8cuBb8w3S8E6NSSV
CHx8UyR+XmaZovVXlntWGBt/rej8eFaYTteZ+zPnajGVd4OM4pe1T+yw0hBmKL81rhCLFWqJ2u/R
LcD3B7kvlTKDupa9O4eBSuWFG0A+0/FWCBilHsQoFXnB6zd6yzb8G+0yGkFHYlaaLULayNfN+II7
s5Ka3n5m+IAC+8XSSZqQvuaeeLYZ2DVb23OkDZeiysUEXPWso8tzHOSa/rE3IEY7h2Nbq3TBmMGx
7XKKDzm8/BrTf9oWHmX+yR6P7OEYauXvUu1k831oIMwUDo7skQ+FzDbvMUeDtq+OXjNdnQ/+cbb4
wP7iLap3WtPQhG2vsEgGkYsOfRLvdPxqjr7Q7zkw8j757RJYLZofExs4WquQSUo+8PQZTOO2CW6n
gs9g3JvcIIBWKSwdhFJZKSZ0BgH6L21gtrUuaFg0rK0uMY7D4JaUyDkNNOO+SUVAOb/aIZHrAzCN
Cz7By06g+Ms7b4kq4zKDuK16dtDeKx/5eHd1pOJ8iRLa0DWr12sBai44Lh3y7eDMOspATCXWV5LA
dBNJv2Cx2n8A1nYyMpdgs1NFbQzR0SwRm5nl/h5kopG9JGUBAAOP+fzFGgKH9m1yHdBruklO55eT
9VWYsdl5j9qXijt/4tZkF/LzphvkcasbPRASHyWib0BXJz14MHhSV5CXxmx1y8HFbgFmQeVftvtH
ZmhXASQHJCwdxbUPo4DlO4WF6jkWim7ju0qJgu5wxiMiLnEqEdNbXJdaA9KpJvIS+pj1FLx13Fsz
53P4aFdzNIbNqFzr7ZFa7u5506HZVmMkKaYzI8WAT1yJAhiK4pBlQ+Yg4yockgTcJo8jU7BjwLwL
Rv0uQFWO1I147Is8q5X/54dTNdP9OL94Y7zLWZayL1S6dQYQMNIdce9KUVYBpKPFZ/0P0XK5VA7D
tS2bCU4UxQQTHrCqLrby6D/4bafb8dmL97r1T4OZSmAFWdqd9P+e9MijN0ypHHDErh+3IqQDb300
teipfrV9IutddBQdwWOnqJ49G+WiZO2nrSHW95ulwNKIg7GGg+Sjbz1FkpBRRzPK1C9JizMPGcQ3
iq7cqu5tAlQ3JGZmWDTgkOSdyrPGj51c5h8qp+1An1AVR+OOq5Fvd7EbqnsqqWmlfkeXDxmcvMZ3
ST2d33+V00Zkoz4hv+qwhxgsMKoR1THg7NDFmm2l99nK8c0Q5SpcO60bPdcl6g91RcriruMjFr+N
w/XXT4BGuGAXDQ==
`protect end_protected

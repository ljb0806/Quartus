��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�M��T-dᩴ���
4��<8fP��K���̌���j񖉾�0v�]\�Tibo�|z8��i9z����]���6� Duc�f���E�3#$����Z��E�1�W��µ���
�ﰰ��pFCܨ�	%���(T �F�~���O���7sQ��4�I�D�M�ǣ: ��e,4������x^�ܹ}Z��R�Hb=��c�)�k�R�
��#�aYt���`���M]i�1�(e���*T��:p�^WԴ �e3�)��k7b�=�	ֹt�b1��(=d*��v��&��*�9�uj�j6TLP��"-�\���偹�-�ꣂ�Fp
�[!�!;]A���z��Έ˳�ݫP��hV�Փ��Q�|鵘���Qz��T=3�J�6�x�A͂�w���� �j�փh�̾�Q��{f��)U�Y(�3Ե���w&k}%�`z�@�~��mj����E��c��v��Y�Iwu�"���M�� Q�?6JL�5��ѡ{2��8�nRW*0z�X���MeEq0Դ4�����%�뤬�"I*df6�;?鮣3G@�UNˍ�v���$CE�Vz��I����5��=��'_���Mj�YTǅ���ƭl�}3�
��paEh|�df�$!�����]p3�nw9�"����z�'���i�%��-mk���M<��:��qK~��y�w.B��=�8Ci���k�E�����1�u��ކ2�^��~������'������>W��;����be�_��J& ���v�׍%�<G���f}�l��|��>�������~4�ڕy�����,�P�n+�-�l2� �y:�+~����(��k�Y�\fa��5�$�]��ֶp��J�$N�|V���)���<b�nlň8�м<�}�N)�P5m\��i!��|4���K����+�)��1��J���tE^D�z
NT��8l"��%%���j��ޗ�o�-����Ԟ�ȯs��j����������c"J��,��s�4���Ǭ��Ǩb��Cѻ��oȟ�T���f5��Ol�~��S�0v����r�K,+� )�m��&K幱�"�W�>�E}ד�S�>�Ym$���l�6>��d�v��������fw�j��~��Fv�F�����:ek�=A���'�(�_�f��S�,�)��c�����Ĩ&*�*WՃ���|�0�CFcf�n^U����5�H�����X�<��.�R�ZC���`���*���E�ɡ�4�:/�-�����Hő��c������1w-��w�8-�,,r��[L��������jQ����(?�iZ�b��
�PU�a����Z���9	��m`q��W���ر� >p�g�'���R����f�)����O�#ɋ�����f����٫��b`���|��:�-�_f�a�^̹�SHd��SxC��A�t��oo�0�� _DE�!RJ�F���'ņ'X�9�4�5xV3�;��bqy9B��M-s�$��X��-�I!��#fs����vTj���  �+�W��P ��P3�5�ȹ"��~'6<e����=�w`ja���wmQ��	�R��ߢ0m��9 Bu]j�q������qۈ���I�1��N�7l U>G�����e?u�5�t��MiU��b��'���g��8���@TYy&t?~�ϸHrD#��C� YKy:���֞���pA��v�&P6!(Z��1��|z�N������ұ)I,]�V�|ץ=��Py	���K�J|��N�H�jMP%mq�Wg�"��|�+��ے�=x�!ɼ�:ʭ�7���4ϧ�=�Of{�������E
;�<�7��$g1o�$���/�KO�ko��8�c����%~�!�d�tp�[����[�,BSt��*>�a��*�JY��6ͣr�{W��k8K)����f��^U�|������Xݨ�gekK�MM��^-y�B�+Yc�)�)����gWs���fM|�OM'+����&��~ٶ��d���d��P
��ϓ��y�NIk8�`0=��.�
�adaC�o�G�Q=��Қ�p��Z�Ͱvd��NW�-{�wƾ��:)�j4W3]<�}6��J� Z���R����T9��X�N���p��l�� �iz ��h�oP�v�Ȍ�bڃdL�(� �H���OZ$=oY���U�:�g�b�y[8P��2�c���:׋
;�5O����j��)��k�Dw�g�J�ɢ,g{�!$���빏�B]�nq|3���u^5������-"��:x�E 2u���$�Hݘ�w�1��- �Y4g�!gK�CͰj��Da�X�c�4aA79P3a��	�HQf6V�N;��Q��o{�q�/GܠԀ�y0��)����~"���5���	F��v���D�1֜�U懃�
��eCS)T-5�� |�b��>�j��S�9��-������E^g�ޯbN�XEa�Y�a\= �R��cx�N��;ԯl��<u��p*�R'����Wc�]��9{��6J�����Y��5!��&�f4X�8!�EMU�o)-B��e�_�B�������^��X�M�(��p)�H6��D�D3�j�:���3s<�-ڢ�uXN��m6I�+Dٺ��o��%
�qD�����u����4�5�H���0���Һ��τ%c��Ѭ��1hm�?��mӚ�aet�L��K���G�K_e�Yp_cg����ݜ	kHp(sAV����$�VV�{Mm��0���!6I��g�ip�bvpG4��p0)}f�*�  <�Q�@])z�b]jQ����b����7p23�$V���� kR�n��p
��ZG�Ot-}��sĪ�Z��"�<@c��E�ϫ�;��w�~Vbc �7�p"������!nD9z|x4��.uWa�a'�p�wM~��W;��JKI����P/֜�C�<ࡌd��C�gR����gm~w��_M�_�`����N0O�m�-%��j�&u,'���>�b�s�@n�8��|]r�V���>6�x�!!���x��gF�=��/w�r�ix�Y��婒�8�j�$��+m+�����r%!���Yj
��˿g�N���,o�
��0Ԁ��?��QEH�/���P2��#<ُT���jH ��k-#7`��_)h�S� �b�)̬&k�ʸ��h�����y�1�$z��r!���+h�H�V��R��x��,Ɠ���]���t���]������@π��✻���4����ZNY����4N-�6s8���C��e<v�if;�k�T�x{�>hl���hB)s����F�un����<g�ڤ'2����R$��"Ԋy�P��#�6��;YO,����t���#� �V��.į����:=j/�����"\����&MIΛf���ad9Jktr_�*ަ �ڻ����C��]K~g[�(0�E-͎�}e�)f��>`�|wi/�%i��Gl�m+#��~S��$)"e`�V�N�(���/� ������#� m7�7N}�������^hc'���]���Y���S�e���cKH<�4��<�cBF4WT�>��!��w5���ַhRpZ�G�j�1����16g����]�C���t��_y�6B��)�	���G�G�q�G�*�K�c-x��u֧S���38�jҐ�SdM֯��pb?3�~���*"���g��2$�7�_jG߲ѓU��&�D��(�Wh���Vgk�����Zt���w�����FV�g����7`��b}>��<s�k�O���܄)M���c��$b�Y��\値I�k�dq���s��-�Rs��t�n�}���u��Y�}��YƑ�$���b����Ҁ	I�D��k�^��=k���{C�#2�&�3?s�A�bB?	�f3�+�6��l�8��nV�v42X���N�ۇ�ʵ�?���j��r\��!�ϑ�e�@4t�=�Ղe��ϧXᑬFW��L��.��^��=����〕�b��V�?��j@6����AI��1�j��KŮؔ=E�sޙ<�4/Fj��Fl�7K0i� �bE��V*H���N�,aX_4C<q��s	w[�W�|��ܨW�=�!��n!�S�Xz6�  ��H�m#E+'�1����S/
x�ې��v�P���_g{V)�{ T1.NXclS��f���|�^`��f8�
⭗xtvUm��������>���ˑ��ȥ���$f6w$���b�q��������Ao'�s��4Cǯm�`�af�ğ���<�C����q_���Hv�_������:�Úe��%M�0~5��汊vG�^#�yt�j����e�0AXEƓ-��]�;y_#X,"�6o�N�au���'�nйep�y'^�{�q�/,�b��/}X`�߭_�^�{7(��*��?`���c���mc
z��C����ҩU�/�qVʽ\�R�uq\���o��~���:���2n�E_p�eVu��m闱� �m�m*J-R�+Y+���y0��k�5��z��To^�9��3�ф�o�Ԋ�f��"�/��e�6�%���r�G�?��}��,�YC�s�Ck�sڃ�\���=�$�ǫ4�+@��:����Ͽ��#Iܜ�a��U��E<s�nm��|˛�j2���P��m�2I���@���+?R��)z�=�!����*��!T?s>�vk9�w�Ƃ�VVu�A;h`P�Z�ZH�|P�b����и@��V/�b�R��\�1�6
fwz}�~I7�pO����"�����nA�f�� ���g�����=2�A�z�g|�[p�)V�L�^[nj�qe&N�9(��Gep��Di�^�.i��ǭ�,��(2����\=-��oWtΩR���.��><�#���+Y���F/-$�Ԁ֨��+�>�u�c��C��T�s����>Z�Һ�F����؛��=��8�M��DHc���Dԭ{�	�ğ���VD�^��iuо$�CT��	`����2�m4͛0� @��A�m�`�f]��瞋�)�'���l>ѯ�X�Lt�(_ŊEB"M~ǈER�\:+�	.�B�?\��{����n_�'pT�ű@t�oSsOV����߁��2Y�����>������N2V�ߢ·K���1��aj[�����-���ۀ��+���Rn搣��:�+�!új�w1���{]2�Y��l?�A�JD;"\|\1K�K.�$"2�p��I.^�,A��}�ne0eQ�(P0�W	�yH�;e����/��#��3���W� P�渥�>3���L�3�B'����e�Юue�U�4�_�<��s��3�r��L$�sL�U�g�&�{cl~�y����)���mv����$+2� �Ji��$J�vȖ|�?8JՁnD��$��W��(&w�7댦V�T*�8��)��@�.��h�����|d��+��V���r����3��?�s�����+w�����&Ŵ8Μ9q���]�}���ׯ�����?-�����dl?��AHXeyx��M�ۚ�	�Tړ�a�[?�[zc�uf�%~/�YhpN7gt�л�!��=Q��S��]��Ʋz(X��og�,��!���­�Mp;�A	%_|7Хq\��2��Ql��q�X.��K>�iEѥ]�G����V`��c����M���AE��a�&��=g<6|���#��f��Gy3՝�\�̉�K��;�ob��Uܕ�c.�0�+sH&X���_^!�4�X�l/������7v)m�ZB}�@�-�p6>���Q7�j��0��L8��(�>�K�J���,�;�}�6�/�#C"[P�����I��GUa�7yz���m�Q�K�؀uꪚ�}��+���4�|@��J���A2[�M��_0��M/�⼔�bӖ��dI���Ksͨ	�	}\� Z�UQ�����K��̂���};ק�ǂ�I���i�Avc��q�{ڃpzdeCv+��]gkЌ�I9����8�	x�z�縲�ķ� u0(:�w��2:wU�_�����F��[��� ��k��}�g+h�P�}��%�ah:��⁪P���Vu�Y3���! �B��ذH��u�+���`$�}�L��v1��Tc|a�0[�����^�t]GT�D(ñ�j� ����kj��+����H<��q�C[8T����c��]^f���;*���{���P
-��h�K�T�B{
oj$��bK���Ϋ�{F`e^� d�'�S��֎$���e�*���1�D��ŕ;�E����u?���"^~z���>D�;��	ON��!M<5	�ҥ�p����a��??_�b)G�83}��m����RX�u�N��Ǒ,���홐��h�l�NNP{�x6�T�[���DX�*�R� ���1�+�/$`�6QG2	�󌒛�o����&0��l�]+qg8�����Rw�&�'��7�m#��{��^t;\��cA�(�gm8,{����'��	~��n��/#c�{LW����3�>v���a�1B�Ek��� ��@�`���&�O�[흀��g[�����ٌ���TߋD}��5�����K�QB!�VP��,�X)�0>V�+��;�[6@S
Ry/�b��f�-�2"�H�UpG����*��g�
���d��>�80��W1E'��������h+�X��@~�J��9�P�>�f�T&�@u�sd�Q [O�X/�ٝ�h	&4����N�i;�?���5O�e�������ۋ�_O=^���\k��)�F�<1�
��q|+��s ,�O�R��,9:�߭�����)� �*� �JS�q�§��c5���_*Osz��4�Ah�����9:���(�� y&	�q?�7�-��],�`��pSM�dтF�����\��2P��\$���c+ooympU�!pc\�ٜ�Rd{�Iy�7K.����E�.��/����G�1�d��5w\?��Go���[T�/��v:��Q ַe��f�Б�½l�
�p�K{Uϯ�P�3�M�q��5��7W���ƺ.���l����T���v��&!���`Gؕ����V"������V�:�%�g�HKH���Pa�R6�LƃnBK�ٷ��d�rTă�_m�j�Ak�`��YG�K�!�R�ӱ�g�ܯ�P���Ԅ�>,E��߃Z�ҝ�Ŷ$>�|�U�2
��tj|���b�)�_5	gx}]��;M��س��Ap���$rE���y�Uj�m!��c�-��� Rh����y��� �u��[�W�(P��&�]�@d椔v��9r�<����t�L��^|p��ϴͅ�fV,LQ� ���Xet��ۈ��.��7(�z֏W�QC�	X��l�b�`~H�/A��b���TXQ�=a:����Q:��>*w�_�r�h�sf�~C�9��)5�j�Z�\�"�-4�)�J���v�'V�&$�rG�fIHSseƇ7L���6 ��ѫ����G�*��w�(��V9Yt�ޙk#�7��f�#�3��l�#7�#�Ϯ�{ٚL��#���4���B���*�@��J�b6�<+�����&�L���J�-���iz�ޏIXk���A�42䍄d2�$���5)�.�)p!�d)P�/J�4ӡ��!�%��$_)�C��ZLS9���ihKE!0��6�<�����y[��̓�\��x9���Fcˠ�;��"!-.��~:��wRZ��;9)���g�W���6U�剐�g�-be0��
�f��[��쁰m4�jb[�����x@��P�r��E?!ɍ���O�������y|�Έ�<SZQ�O0���y��'B�BFW�3,�Hz���R?���;��
�B�5'��O�s%幫��(����WJ]��,�v7�w[�u
#�ٷ�z�1�����%�h͚<�z����yb�g�r��qi!ֆ8#A�A�m�{�?������vD�ȉ[��.a앴�a�_��V�$f�b �58�l1*M�P���bE��N����������|G�ط`���z.�iJ�s��g�>K��,{����¾���SS=��Y`�B�V��������S��B�7��'�kk��v�b{���9R�~�"c:q�}@�6e�N.z�j�4Yï|j��g�F``љ���T���2��	&[ɏy[�q���b~1�;�k����`�O�x�{�*ߊ���\=�^X�C��"�e^�RK!emM�!��h��,{�5Z�� ���	Vs��w���;"mg��f���u�@���ǘS��R�E�\ǕF�)�b����b�m�:׽�����;�DU���/KgV�)���ƶW��dCl��6�6N��z�Tt���� H�]�Ė�������Cx����5�X���e��#��=� ��G��:գ 9�`�4����Z.ܽ�J0SDؤ�k���,�-q\X}k>Ճ?<���������!|��s��|�z��T|9Bo�2T��u�?��.����"I���˶	*� �5,)=&�2Z�J*�����m� gݒ
�b�,҅s~�w�E�ZDZ�w7�D���P�D5P!	��V�t�S�ԩ!�$�}����ܫZ5�^�d��" y�8�a�t�ۨvs����#���A�t�i<~ n�Z��DԬ��қ�� ��zq�풟"��j�jՋ�8WYz���9�/����Z��#i��	��e�#����@&Ϙ��tϺ�&!�A�ɝ��dzEH��$="��h�T����f�i�? T.�"7��8䩳5��	�(�����I<y���A|��4��[pv��Z�8�9!����>T=L��>*�OZ��9��1�csp�,|�/��^CN �.�aK^}HB�k�8Bk�J��dᝳ��q��-�x^�>�φր���=1XJ=�c�(�#����Сͣ�3w=9�:�/��i㻥�ࠂj����ͬ�fFj�4���J�����M0�b?~$��ޫ`~�n�$q���޻A�<2c=�-i�}?u��
�ʹ����X�\��^8D��d�G����^hI�����@_���11lg��}���񯴥�K{+O��g�WI�q���Z�e\tf-e���Pi?T_��a��gǐ��FĤ�N��2� ]*G_ �դ{�s�˅��:�Wi��5^(����6�g�s4�xl�B��=l������tg٪��\�+Y���R��ҹ��9R��H�'��ob��4��É��|�F��5�u�Ҙ��*�����o��B��ȓN�!@��H�{*�E�*&��ԣ�������|��~�]߬�1�0k&���U0K���k�6�"z�ke���u0��ËNo��Ǫ�^wF�c�{!�l
W���(A��aYmѽR4������fjL �Ԏֹ�ܘUHj��/z$��m����m�
�X��e7� �����۶��anoP��J�>��
�?��7q�,���m�����Ѱ�c���g>T�
�&�H��ͪq�1���*x�Ԓ�&a�Spfs��F�٥�Й\F����O���<6����������?��l�M4@.X@<��r`P��r�E������:{�L�D���� ��Y�o����t��m7���:q�Y����X�}GN"�p]i {��w$���ՈĹ�)�JV��h(�3��A��vLen�>,sv|F�����L������ǲ�A�k���D�'ћq�?�T>��Jg���CcrL��k}��=�o���OnɓU,����o PVɆ��(��z�C˱D ��r	>&˷� ��~��유ܬ�y>>�0<]aK�9�[��f�#�Z���,j
�����c�	���N�d�"��s�;����kFABMr�w��N[��Yx<N���
�u�K4n�hXdD����?���o��;n�Ahʛ���Fr�ib�}�o5�8��D���3����d� ]6=�0<��=�΅�������+�о����Vv��
�@��Q���D�� l��ԧ�Z�y]^�ͫ��F$����}3cnb�΢�T�޶ŏc&c<��G���A �R��4�R��M���gf��q�*�݁V���(�W����m+�KwA�9�L��Q�v�4ȶ���
�MΨ���Ŋ�1�1S%BVwȕR��}/�$��Ɗ���H�+M��ZY�d'�}�k��KI_4�q2r�����"f��`a%���t:����Y���������C�����M��z�кT����bu�.��4;?c��hU��XsO��ƥV�nWq���{(ӒT2��BJ����	���2Z����Tۦ���* �6.��(<X\���(�����n��5ӽd�\�j��'-����	N��_��_��V�7����Vl�F�'٘p�9���5T2���8[���Hb�LjM����o��j�/+�j9g�}@e ���@<JD��iJ�''JFsC�R�"�:��9z���	��U�q���]ǫ4����BV���v����������#�rV��8�;��"���k�C2�@��c�`��1�G���b�H���X�Mn3�{i�(��x�T4��b�B#�A|+e�P8{/�P�������L�-̃����Sl��qw���Z�n���������OX'Ьx�b�[Ew=�>���{M��Y���f�I�XG����c<��/cX�&�d!7 4_QFi�v�
��i��M:���"d.��`K��6D�_-�%����+3�`ґ�1f�8Hw���@/�e��w����m��|,9#I��qla;$�Wo5�+�/``��m���8��긠������~o��u��	
��e*�_=	/�S������t`��t�
.GS��0d��Al,䬁+�1{��9p�/'D�J �S�O�O����y �+�vz<\��ϛ�q&��JF�u������a|��f��E�߹'y��x��ﲋ̀�
���;��L����w,\	&1�i����@��S2s��R(���-X��|��G4��^�$x/�
ގ�Q"�=n0+]S<��Z�����d��B���,\�!��N+{@p��D��8-��VU�z���I`������f`�3�����ZK!�{��CR�3#>���3�-yI._�Mxx�՝.���i�}'V,�i�v�l��6.m���.��B8�rQ��ڤ�
�{v��F9H��b��:0��x�)���2q	�R����M���S�6b�'q��r�zz�*����\Z_���usQ��17+��#]�u���+4��v�U�ʞy�fu�h��dd�>j��Ok�[��+�-r��:����l]�o�"M�I�]��_�*C��+��W�*�F��mU�e4�+WUM@n����	���f�L�b�������rS��P!��)}���P�W)3CQ�-�a��m�J:����$�Cqo�<�S�#����jA�E �y� u�3�t1KRJ� �����5��i���$%��4��	�T�K���*�[���s&b֞I�������cH��O���C8�%.��������6����rH��y��H��j�3��o���I	Ʒ5���=�?�޹������du��!/
7h�o@(�篃�
w+�م�r���k�st2���3TO7���b�u��zƞ�)pX0��d�o���ε�ګ�5���菞���6qN���h��א�2l�Bc���O0K����>F��i �Z���@�Au5W��x��NH�I[n"���R:܊;�z��
�{%�c�I�U��)ů�A�Ƴ8��cq����O�f�E6�
��`��0��]]:6?F!�|������~��?I�{C�����>C��J�?�����:ɑ�������7Yc@�P�No}�&�D��-�vU��YEf���,��n�44�ת}A7�3�G3֍;6�R������_��ϩ*C�XS���.-�sB��H�J�Q�ѣ��5�žs������4ؠ.+JQݶ�JVpl�:p�n�d���H���~��V~�������Fqr�4�E���Zԩ�5'=D��Heӕ�PD ���i������ï7�gW]E��N��]��'Fa��m⿁���3u��a��Hj�5����f�W)��t�QH.0!±3��w�s,*�`JDw�s\��~B&�����1Z��b�>C�Po��7����ˁ�7�]{������$��t�"}���)ɔ��#�J�����͆�4�D��ˉJ�^vh��k��QZ�A�hh����[᦬�8�>��^�f�u��<��)*ہYYoyї[�J� �b�d-��1|(v�;������T���~ն�]��nM�G�mx:���0�]1Ȥ������ځ(�|KU��-����b4������]�|.꫿�0�'��E�F?����١�,�*O����	�4
�E�'e<ϭ9���e�}1,��u=�+1p9�<��,ft3�D��t�0]�e���:��d��<��HԼ}��R�O�v�P���b�<Q�L�{Fп���~�r��z�}BVH��D��!RT�M޼�Oh�A�\��@���µ|�睐�c��Q���h���*���u�yR*$B
�ȽP��c�n��W�wV2z�1HJ�,��I
���F�'����������0[�E}�D���.ޤ������&�����\��v�͂�:ű�q��>
sr=(e�N
#��Y�_�e:t^���ZQ�9�c�t枠�"��;&�k�ɴ?	��i�[���jΚg�]\��4{!f�x�R�)ekbwW�W]�3vϤ�2~L�@/J�ا��Fk�۪U��+
L���?,+��=1W�)���k%__A�؎�X�e4���^�2����9���\�s��d���K�<V�%d��6*S�k�f�\yКe�cfүQa!��[��\�����oG��7�����ʄ}�C��m��b��$�+ g�9���c��a`���A�2 ��$��vV��OJKe�
�>����0L&�W���V.�fq$���g���͔&��K�Pt<�<��Į���*e0O\���G��UŌ�9��{wBC�&�p��
�~�6/|�z��&ѭ��1l�Yy_��#�J��?3����P�5���)�@����="����ªV��S��m�C���{N�}+v(���9��$_�z�u��5���+�(��oHD��+^�(���-�H%���l�0D��Er��]����(��3��yX�D����	rBY��ʷ�C��'(��d:��%.�b��FV��Q(�rQY�	R�ʎi�V#�����?�VHG�1�7$����3�����^8Y��]���{���#[�҆�J.L��1�x��r�7����UP�MM3M������ȯbh�.o� )DX��0<b煤�ITCFo�9��O�4��yCc�l��ga�/|���S����6�E���9{��nΡ���F�1����=�����}���rmq��⺕S�5#f��J�7uj�����#8�V���&^�������/ ��.�QX�X����^L�a�]���P�զ��wn~�j��Э]�]]�=�U�8��M�נ�������,��pg���4�j�������hrwt��S���
`(8�!��М� �*���}��`[�yN_��0�;��*!�� �5[�s�Ҫ�Oce�]��l�S�C�b�����3rҴ�6�M�4pvr��q���p��}(���F�a�'L�EY�59��n�\5��/�"a�v��/��}��Bܶois��כXׇ��w�sB�P�<0�:&wY�Nع�����H�����`�/�6���.��O޼�8�e�~��٤��x�i�D�1�V�E6���;�h����"��׷.�bQ���>;�9��m�r6�5p��Ņ���B_�Gi�k���8�����SZ��;#��q>����]`��Ϩ���"�	 k��ay�=k��ޤ�3�/
"$��A6ׄ���@�<U�,Amp��|�$�]u�� sl������H�!��R4���A�.���H��[��dN���/��q�vw��VL�f @x�&~~~ wH� �}�븭��[�� j'�g���+����K���YX_7�CY�6,B��2lb�� ~B^3ȍ���Yy�1C�	H�3�\nڎ7qlO�T��{�E�Ԭ��A��:՟z�o�# �E���8h�=1��6�yPP`v�9QiՆW��+ef��Ӯ�K����>W΍�V���!��0]�A�xmN�����!i�&��@o���Z@��6��Z�ȶŶ���(�����z��ZUR�K�ƚe��{Eٮ��0�n#������cp�g5*�������ܦ���GO����x��>. �J"���E�LA���i�v!A�23���żm`ֶv�e6!ns7��˫����-XM#e�>5*�1���M4$�u����7h-�2@vz��4#�������W[����C}�2���eBR�� �]��^Kg�6�sj�Y���F4�ņI���&p��8�e�F�C)O��#����I@x(*�����O�I���FZ�shd|��i���yz�U�\]\eYtDI�KQ���d�̺5�p��8��h��ĉЌ�Y5	= L��\KI9��[�'�/��$R �����Bɶ[u���\]M^��|pz`x\#=�p�����q�\���o��8N	��=�z
��[��H��Fb%9���h� �����3t�����k;��:���ؾ򗠉�K(ј�i��ќ��)�驶�iןa�3��$}�vx��Q�3��ND/9��b�&M�� 8���}f�m3*\�u4J�Sz�����p����\-���<�Gd'��izj��e��IW !FM=��ڥ���lѬ��ݪ�!�٭gDt8�q���p[C/W�c���z��!"�9�ȒHE����˘�*�3M����{�)�G��m[,���	�O���}�������_����5���֌*�.�͛�Rȟ�[5��Y�.N�fJ�ST���dr�xI���<�{ ��q�� +��c���Y�:�<u��(��YV7�W:j��]{��(D��J��{Ț�(�7-�H��n#Ò>qڱ$>�J��w���sVq��=Ê�n���w�� ���e��#���V>^��OAK��x(D���^�Q�0���:����.Ɠb�����j8��&&����e�o�f�Q-U��؇t�v�6+U.Ă}���#]��ᣕ���k�����j��O�e[�˿�s����	�7��t"$�ڦ�i��/w�f�a���5��[�Z<��3�K=ZXVp#��'w�o[�K�2���g��"9I2�Pn��(���\Ē��ƭِL�sL���M�jX���d���5���Ѱ�č�H�Q�ɂ&�;v�֎>�XC �A��G�N��T�i0)��j��^���1w�R�q�vQjx]y����+͛��V�G�JPz�d�ߠ�ި��Zi*E����^���'�r���n_�20g�5F�j8y����.�
i��@���E� �a���ĥI9%��Wz?�D��ICjn���b��@��.����d�*�?=�0S�:�r����+�j���}"_z2T�[���u��Oa6���T���C�]�����v�f�pw�qJ�I��'���ۅ�k�g<ނZO/������3ʟ}�����(�(�&,�T��2����~{�-�ЅB�ٕ�Oc�����Z���е?�M��|6iB�g�T�wĻN�5}�L�@��|���6��������1��/O�ǚ�t�'f�;S�Iz���1��Ѭ���\�J��h�zo��.J������5�7\#Ciʵz����>֖,�M�I'�xj���kV���\y�5j(�/��e	pHK���
��g�B��X�\d���A�?���&%7�G]ID���7�=���7i�ߙ.�*UuyC�
)a�e�'��j'�6Vj��E��(�BoXT}���M��!��ʓ.��9�B�o�akj����sP+#�*!��/�'��V��o�K;k��|ٍ��Ԭ�ᘆ�u�]zkl��tS�,�J�D
&��0�t�zq�q�������n�jh��]�̯�y�dm��&�?P*2��G��y�jA8�/3���:��1��E�Н������9�Dڇ>����V����N	`�j�^ĨHV#߅��'*Az@��w!��O��Y���}�������@N�ɖ?�"����s�����W�V��yE�����4��A��!5�3������b�^�[&���}�]*��	-"=ؤ!�Hp�#ʷ�NO>9ж2�zד�*@>5�2u�V���(o��^�#�# �&ekwAt	
i�t�znrW@-nv�S�$����P�;�.p��B�)�3 ��?����m��Kċː�к��Lf\��plA)��-<I�rbUg�Z��]�1�z�ea|E�&UH�����~#���V��\�������;)�C����Xo���]�H+�l�^�.|J�EV���_@�y��Y���Z<��R���>#1t-*��%��2/�D!�E��`�M����0Z�e�/[`X���m,?
ߤ}�J�ʏ3.�{6�n�#Nf���2�4n��'�X���V�P����(;{�"�R[�]�IyZf���~���c1<���<���u��������.��1���ڨ�jƥ�[�M��;����q����B��S;��@�Dv"EZk�U!��>Qxe΢p���z|��,g�.́8��c�X����yʰ����E�l����t�c���|/"\j�H)���܏���?Ɂ
[�8>5}�!x�U�N����>H�Ú9U�Y@K�q�å�*W��[�?]�=�"P���!�����>��KP�.�QM.�XB�����#��yr)him X�����E�C�p�[Ur�{Ͽ���7r^���+�3飱u�7���T[�:���ݸ�`�Hr~���lr,��J�K���H�8%�Z�,(0��y�4��ၪ�V�(�m�s,	���u��dO�!TW���kT5~��~ɐc@-˱�
/�U ��HT�;}�Qd;x4�1߃�w�{ǣd��&����I�F~���ws�Z�$K�џ>v�+���e{���V�t᪫��+�
�&:/l9�x��������bZ�8�T�l�ug(y�c҆k�z¤4l�F���XY�fφ�u�Ѷ|�,S�R�i��`�<�^G��u׬�����*y�F�I�@��A����~R�� d�GA��I��[s�%�P��i�ϯ�j�j��2�����]��χ}��j���m�������F����6,&UX�g�d��7u��m����ݕ׋ʊ��%.?t	��9!e�z���zjg� X���Pi�f��,��#�&�bڠ��O�����k� b�l�ţ��bx��y��3�� !�
�}(���n��f�k	��U�~A�3�rE�B�� ���G(J34���W~а��{>�0�k} {k������uk��U͌nY�J��[@ug��YƨZ̓Řg[!�&�����b��3�}��]Ka�p�I9hp��lW	����T�@f=��)z�;�G�7ڟ��Eֿ�"�~|	�W(��x͂���^�p���7P�1�"�o+~
nҋt�9w�rg��U���k�.�V:>����#�Xw��4�_Iy���XO�f-#Ԭ3��C�M���R�])y׆���+cF�`ˤYgj��7���-���E�#�bߍ GZ�1�I��(%�[�fت�.�@���z��9����XoD	D���, %���~vG87%���.��>a�	��+�e�j�Y�))�ڝ����v`�f�k�o.�G�38w���6�<�4	֩{��+�̣Nryy���1�Ѭ�����`7U�h&��d�W�<�l�11�M?cA�
P��V-�@ڑ��ɭa��(eF�^,ݝp>�3tnT���#�|��cm�x|rD�)A>�K���(g�)���4N[�n�kU���N�D�)N(�P�7�,�}���s��H�J
`<X[;���9)��K���j��όUA���6Ȓ*ngA�5�|9�"��u��f �l����K�
�{L����	
g�@ԟ؁�me��z�sn��o���+$	G�&$�j}�	b��5��D�^�<t��_�!n ���㦞X�����Y�L c��g����e-%Ǩ�uO�Q�8�%*B�?�%��p���O�
څ�+.�K���ϳ��:\�ˋ��GK'S�d4��>�u=��R�e��>C����`�.`݁�v���}
����E]$�UXs��#u��+,;����@�� o�g�@���V�F4K 	��R	oBį��+?�hsE����U�rBN�0�;�1���JR0Q�d��R��H��A�F9�)��]T2��RX��5V�B���"
*��}2��'`�|g�Z�Y����n��*u����㫬x�)��d�
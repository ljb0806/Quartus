-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pXVhQ4pfQ2nc9l/Es0r0UFvDeq2/3wqC4Tk6Dp7HOL//0qQ5hABnovlUISsN73ql4msATrdceBBw
W8Xvv/BIe0T5u3+5FcFIIplv1MsNR2B6w7pFzlXYpFV8x/Ep7JZgFZy5wmVD/45uO0gZXEeViUAq
79i2WNbnfhMB4lirG/C8Dc6fbswgKJHBQ1wuLCDCw0J5MDdZ3EMHWm/vXnooy2SE3Id9hZ7v6lVw
EuSCsuyQmIp0IqUygGiGy1NG1YUGoTF+EeVVMylE2ShIwTKinynaxm3ONlQVi6ljxJG8359kYY8M
7s1b/edOYStLCOJGnHCArxoh+4Rpc3ZtXj9roA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20864)
`protect data_block
OVApJ1I5wjJxCCHYw+XrN1fIuLZWK+4YI9ddL2XpNFRZmO5U9n70n8ehs/uwkSS6+lgedesdtxYw
LYVI2PmLnMmaZ7Ib1p+R1YgFP/rJ5W6MEc81bBLvz+G4MzfT5MGzdm4DW0sV0Ov4IrjjZoBJb/O4
SMWNYUbvFAWT9WyntdBbQz6R0ekBX2/85MED32+/3207SXhl9OQ6ewfEnPkcL6GOfZ5pIY3KiWNh
Fh6uxKLAJtasp0dRaZL2US/BqiiPuK8TEsBPT0U+yIQEGFSE/bqdRBZvDFcWHAtnCQR1k7bSpVJ6
LoaNQO3afiB6lmiCqJngZC5QAxntN+KyC3x2qVv4NudTiAQK9PcLohojOGop5B1znYa6JnrUbylA
yUkb7aMfoXAKPiT52HhKW9g1cA8UFNuuyx0foqG0Tk0uxepGhneJMvxqvcs0EDMbcoUWYEkzt2Tc
rDle6gKEDLRrYITKcW6tPME2W9lAYg3eg9Tl9K5oUz5gTnWkyPEwfjMWl2o80BcIFnF3TmQITpWe
djDP8MXLyhXKaDUhzCr+wcT9nj0DNJhKuoy/DOvCSxIsMjRJcygwFWV86SK5rZJTqcqe5D0ImH5v
waEmeSE+5E0DB/FXNZex4+IzozxhixEhZxvZ6RM1OQDyEwhc/eXVD1DYgk39XZFwDyD5cTxTjVcD
YoxyFwI6jyWcJbDBdRPKfJ+0aWDpTAu+xlTnnRH/Jgm6Xw+OoSjQVix1h4kHpTmPfDvq4XR7U6IK
h1vI8aWQuqjPe5E51tI9XJDlgyjTJB+xRYflIGsY4FcqMpyWMYMYLR/JBy9uY9sPPmwBTr4VVcgS
HfUF8GGT08NSVYYMNuDA4jXey2WJ3irST/Sgd9tOAVuuBdhNUVrL1H0KS/fY+2uQhExsl/7GFria
lxlhBD3CTfexrcOnwfW5wEgenpMp+qNB9420QlG+xDG7xOiwTwb9GescYaQxgoHJBbd9rq2K8inK
Reg/6FKzoBAyOiMJ0YU/UN6I3MnFb28hq7yOX/xLQOf+QlmLjXrZApJtpBlLrf16ItrtJnVXXUkR
BDa+P29TFnUbncvIBgbYUHr0hWxruMOS1O70vTOByfij6IpSS7/0eihuhZqMmir61+OcepXn7zxB
BfiiZT2C3C0iH43eBAkrDGA7IpFanDkeme/ir+dlwfDX5sRwTvhm/GhT/EEkTqsXpbWHa+5G5NzX
Ku+VfjzRRQh+43h8FRPQ8O3yKh6W5+GXF0OR50KNsLaU2matZ35c0fTGE+KT85r4G4K3fiVpzvbR
JfaWh3Z0ynQuZOUCSK4YXIRA4Ilhakp0YWOAxZIQC6WkV6TLM0TTsn2XGGdKaLULk+T4r5T4tWjh
R0j56EKlAnrlAEW/wYX8hlw3tjOPJB3DKSJmHMZHur1WNvI5jM5sHZOvoWnuAQfH70obHf8BSFg1
BBSnK901jawLPVZPnKzAPt+zS7aXar009AGt/mrpBElmFbFUNKTyoQ1zDxMACsWe+ProCwP70Ikt
5B7VZZ/3dQNtYNwge+xoPdOJN4IllOBorKoJ2j4+qPNP8OmnQReFNtQzK2RVrudqXsBZGXZCfwUN
V3Urn20sRV+WXRkkp0UMr00cLjDl5Rutrs4C0P4UPxNDMKEUXDZigfPKXQD2OgcFOlmRpMp8hIuB
DzEZDw0qNc9uP3p+os8byP4/0hg0CJcCmNTbQ5u9pyxaORsz32qabAfmsyOGP66hn7i4H+GeQ8cn
SSvbBgXjtYFvJLyc4rEhXsdjRrvZw0dmHgx3V4urjhb4CFoJA44sTyXZtgonMRdBKo3kx4V2MBuu
jsNbO8J0wiRfyjj3MY2+57Y7yuUhMCYhxnmu8tEStr2BVlkCWxwSvqqvEcZy2nQDw9orBMJeKk20
2O492Y3KAo4i8wq9gx2oU4E2S6laLDS+l54yDz4E5k7X7vBBbNliyRYLCF1Q4Cl6K453GftKyhMZ
uZokcfjgdcSLBnegDUzEOxq4wyv1zblw13GgcI5rrKxnqI+b5O61T4k0utVJE51bseqlH7yfGkh5
dGnwOkOVjlByi1luTymcdHQ8OafpTqeLXaVQfIqctsagAOJ65CoW2zVDtMgKpbrjfeB3NYwmn5N9
Z0Gvf3ylmxns9Yp/Sn4J2ix4pHrGsgEU4GhBgEZ8fBo3j/EjtVS9Vt/plFJNoQQDuD++7rY08BgS
ZTvmLGO+vQAI7hZ0r1davwzVoeGxiFdKVFgN+b1p5ZOaVG+lYWQBxeyM7dAiUHtE5YP42i1Pt7aP
f4zwriiA6Po24BXVjoeN81iHkwDsGOROrgI2fJdZBcDEyQAV2G9nkrnUEbl78eBfi3u2QiUL7vxF
xDznKUQVR5Uh5MjazhTZgQGMPlrJ7CADl+tkfVChSKRLwnlyXDp6HbfzIKvFx+Oo2+7Lk5tWp8Yd
/cNU0ZhHi4nVQoU51WIRfHKZ8sAXDcLU5eZZBWEN/AZubTM0yKLhfaWkNX9XEP3HRrK/5CDQ56P6
FyNvojSpdm4dsrQBUeuqWUmyBAh3DYA8h+uS3oe54IHP3VTrFfdkA8zyxTXkgQu4emlfnzY+9oJd
8HUycjgkZLMjPAmqCBb6+Lj2ZbynDa8MqroetdcfW8lmVv5nvYWv4UTiJxg29YOZRkoEGuBCZHht
gZvNQJRezr6uRAbesqmeKA9kaS3gRLb8cZhhgQDprdL0MQvbzXl/K9g9EPpz0DMdYtV5OKFKmvzU
7y7c8FRuhlbIpy0K5Q+c79F/BsyN+UYxJgjL7XT0LAHQezOGR3iKOipPzxTSWeFdwTt10ZOBhxsx
wv8XZXG/9+DL+XPvLJ38clQzEAPRxZumbkwJPYOyFfekJgtuAIhOAQEouHSL4qo4iPog01aG765p
3duFY/1GG9skFkc4VaVHtknjiRWLGh2Ua5V2TqOTPL+xHtx2hs2BsviCxlXWNV1+WjuhGfC7b6U3
jnx+k5PBH/pfds2TUPT8D/RxABx41UY86lUdVy74YVWxbP9kIkGEDqRjCdx4TNEQr21V4I/eazDP
2YVKiaNqy/0D8q6nggq5am4hNNmAmqKdMIJxBNtNMqyXmAFqM1acYXkt+j2l5NCqzXD1401yy4Pn
jfCUIL3Tvh2BCAuk8Ta+LN5lGypwg7gEuVnL51niss2LQYE9vze4UPvK1WHyzg6nnrjZMLkBGGk6
yPHWV3KKuAfS9YLLYNK2Tsp9zUnPkzzr4/rHQBYMIZZso+M1jFeCj66yYf6to0Lt3fyf70us1L0B
xMlxRJxnC7VRV+EXlgna962ufpb0CrWieXNvj42LTpIouIqwyKZg57ygoKVDrAyjexgqH/4+SVzb
Yc4F82WMuH/TJcLKRAlt49BpteEJec9plljYQoUJepQlrZTG5H1POe4zsRMybWNjNnD+MSC3jPaX
3KobzB04qYNxkUnbv25B9pJVwCOqXFE4cgU9HOrGvgH9y2c5hAhgoB5nVn6LF13dmCfDiTSf7REe
3dUL2qGJlXRXu2kMqFE6LgL0hOOUZBPiCajBYqDuYS55ybxwIaUzEIo+zkGnVBachFBBuCJsA2bB
GEUN5LcQXki6/8Reo+Cy+b/qa9gRIbID3OWKxXbLJagAT3e+1FA972XJpFAsIdFfTLXibgDNUQuV
l3V/gzHHmTphG0OthiW9roWpzN0DAih0A30lySFGD8Lphgb7CE8sX+mavIkqi8xrdvK4DP81Hx2J
d9sjLee/T/dZGbN/y7FCgzfiactjdmIltMBp/zSv2rIAZPzb1Cbjvnd7x+cnKuQs+Y7fmJJZJPWM
alKIaU3EZ7uIn58AuMIk6+tmYYwENPfX52pll3soZQsD4dHgVTVXPob7s8iETzm6YwYXmpeW5Efa
QrPSAeR9YN6PEP/Vv10sFJs03DsfkGdVT+gj35jkQMpBRss1+aNCrj78rGzgZIp+D6+agSMFJoe8
Ch8ScxWSVWvEBzfigmIqcQpYj1YDp1UcuMAJSjC5xVdPaplyOKRo+6Ya7dN02LyMT0mbvXs0Sjhi
1rY/Bx2e79edKL/S5OE9U4XSxv0icytoU6oR4OHyGgMW/jojFCyDI8EQgcFNlYow2WaKfM4vz7ia
l6vcj0c4iRiBl61MGlaSF4/knFYXeKddRn1cZHarXQTqYgIQssa7Ebc4C0dMG05Lao5i02uKvpY+
5xV1zU2pR+DySrx0PB/0YOwJaoJnOq2uGPORdZ9RHloaJPHEjQbpWlnMITofBXj35HdjADaNmmpx
hP1v/oWOr9/cfgfR0fJEh4frPMf0MdbunqTQaR5iAefPs4yBkLZIC7fXAgxWBVFtUGJ4WwSKJ3vP
jU7WzXOZdHcmvsGCIcz8z0tDXCI3Z1q6wvKUywkRLVG0j/0faSiZycSyAaDMYxK+gdfCfhvf0FxF
oeADa/9Ht8Ewd59sTU1QxfivmgmQEiF1BudRk180gdAZmTEUMLR9pikp3osFYkVUwoDef475yTA+
hdFBBrxdjLUdkFtp8Dn1fMeDlqUvV05jkzcWGUkvGQpTDEgtCnxrHRocvh5GRFVYka+mTM0XWMDr
qpcp2VNPpJ+AAbDQR75TeHYiVCeVtqU/KQ/jQAFGvBysyQUcMX1R+Nra88cJnc2poqRTButTHv45
hUZsJGRNE2j+rLQ4m0rmzkH/Gp5I6El9gL+fRmmGhDX9t8ZgCYY0L+LWYoEyXeSpJZTkR5+LiyGS
aHTLJgewJo8LN+FFNBRURdcljAyiFHGo3Go6klElhuVVyLtfBxJRDZZAcBErbIUrA4VNy2aCrs1m
m/TJuy7VB88ib3PGM8DADVrL/pPE4Igjho5pTjDjEAAl7FiIY6H6PwSI5KwrC6y05foOGlFy8cLD
Vxr++am/+jc4ayyN4rdwvlW44zX0s+TFcahrLeeznlcC6q+57HyjTO/V/Tj2ZEDSjCgvxzCNKdHh
c9qY7IgYT45H1UooTMZ1jPP2IDHMiaj7S4CuAiSySQu9VrXxRbzPjyjVwSp4tkFojQK8vZpuAOjO
tq6BwCKF35TfCAyi3Nl52R1yvzivbrF1Rn0waZ46poiZ+CVTpQnE068oMcL2aGse+gdef1NU1bo8
Ih8v++t0AsiDfNwAAl2sE8jrHkdV6/P9EwpnimijZ7YOWUsG0v6AjGq+RSwYOxS0gXVDFoF64yOh
4R3wIR4FnkFReC/B4OXpj+OXW6YG+DLxgLbOOhWAjuxRcrPLihPSDUzPIIStCE3gTZCUfmOXlT1v
VfqUgaItaJOBb71ZhUNqzHK7IrThJ2huCuWdvXFlHau3kdwp4hH5GRqUPT2M0dJQ2Wq0f0+FAl/t
MlcuU9c9OQLoxCCSIxQSU71Zs0Lit+1zm/s/lHi91khiIHRJaOnx75Da6n5zJas7wOpydt6g64Ou
4Fs+antbs4crt947+vcnpsMhawIJ0iuhtFvRMKliM+bAO33jVc/d4JFg/dE9tYcYay9kBQoanlq6
R1hwd8CVqj7ARpB8yEsFr7n75KEbzKowAW6ckx7X9j0gH5pkqB3oKiYSWP2c7LOhtfGFLmf2G5LO
CsJmmQwkjJAyw7gUEPaPa4fscBqq5zGiWMlQGIT9/yoYhZsUKbmxARq+SYmN3QuXEPZYgbPjVwIR
GywyplYx84Ru9odMk/Ahx1c0FIJBgeuNr+gYqomYtm83EgPv3uZjn1qeZHGKyjgDEmz7rwei19cq
7La5cCAStH9ETFMk2sEJP+goRtLsWrqx65esZc7wIZHqdW4w6HF58MOeVrtDQClMtzrGohE2xzqb
q/eD6YYzNMUQ0/1BrVbjYGzfYcAnZfhBMuMh4/6+/tSP/BH4SBxb3WDhzuzn8QTgD43tZusv+6Dv
vU3EQunB0iA4QMGfaiVRsfoIW90OOOlb/RYKyiccS9trZaRZyraIIQe/+NerH9JIMPqAx6q/W7o9
f03okr9wB9td5eHhNaL4CcF2lVcGUYalQ7Uy2O39+umTCMktTPNnnxJ7ucgVwUrfg0rzCSvyJ2ar
Hs0o9BU7LHMRpMc6Jbfma+A80tiyEJt4l0eid5GCkQbg1gZ9KyJijhIZu+iJN0ospDDIlGELH7Kr
CsTTvmJmup8Ktjyd2mrOxdB1k084/q1I3nTTmlXrU0f+beQ8A7uAocNUmpSksoCVkkS1ivF3PlPz
1ZN1RGgYZopA0RBOwSe4Ho9G7Z+98nd6yN2OKuKWn53NSGclqNTcfjseJGa/QQxrAMqxWpvEsvan
DfNrhU8ZRZZ92WCDRKpZBoN5+LsQEc0Fu5HufS54htr/nCrW7JbKj9EYpkYWPISqUcJdKxHSquri
T+2NDu3kipqtvn6cswog66qH0YdwLh+/9W6SJIV4EGQyHL6l8qxkShcFLqebv5iYt96/dXqTaEp+
3VXkcgTdQxBhJ8LWiSrqfBbwWv1SRXVbgh3eJhvHT0VCtFL4w9RTme1HRCNUEcF/rfyfmS4D55LY
LEr07Qjxv0GAyYWkWBp1tqGOjktd+ecbIlI27DV/V1Uv0aShTyXPUiyiw+gf96dLlGPkylR008wX
4Pil8VyV1BVwWcDcO7wgs/oC77SYxIIcLwx/d7hlwD4rqAfynLyPZ7JspP4oYYhjj4sUIX7qlfdy
h1oiat93thp4pOYL+0WNnNFJ0qpe+4weh8MsYVAdHnSWN5F0qDWhvMIEzUcYCfzPJGLrR9x2bMbK
65O30EaffttkRjfFoWhzT9OlcdMaEFiRjU1S38+APWtwPU+HDDmOR/98gcdlJj7FCeOsFofyS46+
s6omZkiBW2L0315ktUtAgAwlyFdfBtfYAh25r3O0aaeOfJuLTXsykScy7kcJtDhUYrwd9pmNf2pg
HAJ1u47gxtu0dOtPN7X73heY6HAeNTs+hsu0ZR/nozVeW2irflL/DXQjQoRL6gibnYZ812PiIxWF
fAS6yduBW6VXW9wJ2BT8FyPxnRAuB9spHe5WYA1Gc8GJOtjrx6MOVAsqeZTTLGKcxnguD87kXkHC
RSpHj4M71TR2qPR4WCj28eXb2x8o8lwe0t33Yp95e4QWjdPcRY3WX8BSAF+00SZxMl+vTM5xwgeC
twRXtVOLdc4HoToh7r0ZKMv3N78Wx3dDBqPEQpIWpqaKnI4EQNbg9XdW4CU6VUUdOFZOForMFLSh
dNNgphqOQqTCshhaxT0Mip7+SkrzL2V55otBcwfcTSeRuDIwdkRanc/1KABHw4xpMbFrvDNELi0P
Dw7f/uW7xSTGwEjnuMM9spczwk3tCt8/iJuvYXU1POKVqaEiSY9SnDQxA8wbASqjiL+PMeLWVURU
Yh2A4BLl66ghBh2JJpJhNNRxay71kSmRGjU1D/70JLkzi+CJjn5qs8yxJy8SXqJavfigR9KPzKqF
2QBJnmFo77vQfJ/IRSD3+szhmKcwMsUNH5HAATHDahtSipX1Gw2Mick5LPu4r88NYSfOoMTOrzeW
dar+kfQL6QePz2UuHJQ2LcneWC62kTHutsX2E8vDXfYKv0MVjmLKXtOnJ1JMNoBQA53QfoocTcFg
qntqoSgPlxr5j6o3rPmn1dRmx2K79FsyAwkO7KzsxYJmyejxk+7Zx2PWFldAhg6UbU2fQfdRYQoR
/fj5gMTCNvClEJlBRRjc2OMKoe+hwRk1AY9VE67ro6Ovz7o1koApjLSLH8AlnfaKvJBciIJJqcb7
HFbkNC23z43x/Z0QRDgVUhUbMnacGr6tHlqxz6/BZi0Mhp1aYhZXwb4xJQMnvQ2qwu6XXEQbk0UR
jFY3zP0DaG39wfnINzMAkLbsDP4N8ajLvbuHBidHL8cprJDJLZ790oiyYjrXvDcO1EBYn3ei1sl3
4hJKHyKf2jlQZCntdGrp2RHcqLtb7zAwwh86aeT7IzsTmaQbr4ZFQUoD0t5+FhZNYlCiouR4RjYJ
gextNa0duNi8MoKVMneI9QX27NeqGG0uTO+aRPgJyLfJMmIfB+0h4C0Pr0/DEbElPK9stZlsE17z
dipVRWFcqfPSOTcD56Ih2tOWG1zq6+Zjfro5zlNzNHzGGmq0CNqJ8O1uqV2ujHvi40CTCvk1bPuP
y1oU+PDua3FB5L2C7oTGXTnwfGvYwx+sh0xcIioVYkHx5I/k8PbdR1pHtbRQylbNxud+fNi/iM2O
uRGos0LoEhjQDDfCM8a6QhS+55tR0fXIRQ3EN2AXoSFT/HWoTIdy0MsEalfmAIRP6U06xHzZ3cDb
DDYUByQrB7HNvFl2UWN7gLOHyOYBn9t25jaTIA6u1+xmavi8OyCIHTXSnMl3B1Jsj5I3OMEl9KHN
kcm/r0dNruhuOt5A/ZGwQA2exyHApL3tf4QUZVM8Ppepyuui/hwo2Fi+M323aJZtUqtjhwh65PKM
kNzXl6gIFzk5bsNhiNQnimiVdABmRrdA71lKG+p9wFZoS/ooqlZ6iDYEStzNnZ+P9kcjv0TPzbOx
+1woEHhX1D39zm6o6PregzBXYrV9dumvaoFqnZxBlbJZQbi3UfEUWk6z4JORNGkdO8ASe+ghBJKW
TG+V2j2cr09DyzXBmYwVIv6BPvgmp7hENgx0hvEQOx7p8+TXcAqeP/6hfzyv/9yFTWmFJFcG/9/x
cW4TbbxVxsWBl5rQugSUdP8OJS8E96JnjcyV4fTZ8tlMZ/lcTWwBEO1fWbmk3/bm890rgkhwP3rd
FDQA9nebgs9flMXBJ9WnSRPVO4dC/A2R6gJyuIRH8Bxh7xkSMhUC/k8Eyp8ul3hNZIFs5C/oe5/Q
hvrGFFV2wxzLLFsJCNh/ht3LGqeVZ0z8u/d5dv4LIYfm0ma0+B0P8ztm5M+ehjn71eOc2StGm3h9
DjHnr6o6ZG4T3JHNcLGRHd8Blo6kYYrHwKxKuSu1IOy9TQPbc4LOR7CLBL8FHrBWtTpUmelluPSQ
dgl4oSu3UoAeK7MHHX/E9afzRl9M2glmY1XzLmZYqjPux86KhVy8PRjWbpT7lNxsTK5x9TppM4qM
fin8pmfGQ/fvBNvP1hhs1OmA5uBHxxwc02+MQ6pZm/ARBKBcSB2noSyXPAdGvjCAamk1psO1AmQu
RqG6B2WrVlcySOJIHHDnYM3QJ4SUj99mmCe+YTVbH23PefvwREWykN1u5JwrLyaioZZtQIqZkq+s
dI9PmwJkfORlQ5J3yYf+L0QZExoserAp+eURa561KxhDBXh9GbUkmLXnh4N0olZZ6jET1hDbyw7n
5lX7PJV7MLMfFp9Q//MBhJGBDxpfaqPR7q+6TVb/477jPoTVfI695nYCjgz4hBdpOCJH4YIf3Tp3
f0e5cAVvEz9EI/RqZi9qIy14QkrVMPjp6FvST9yWlbgly+P+JgJ9932WhkYpBwMveXoDuQlrDbyc
Qi/Zq9JGJjnOsFCLlr7bUHqSEZ8CmwLfAw2KarRwAA61INso5xPi7tl9+tPzeIB1ty+behEcFauN
etTPDZCmSJbVU+MyL+ZT7A8djsCyEjX9oOHB0d4ujrs2GckTm6ERDb7PqLRz/zUBWAs5yJ/kadAy
qpci9H3sERTfBZICurtipvzG5P7kyOpLhlk7khAOZvAr25qgPT73BQ2TJMsJ/b9oAI5udtLX+qfI
OtFBYwOvkGxb0stwvAmHbr8tqba7XyimCvRRtwuW/RXA7q+8tuBSP41ZL0XjaI8K+fW8r/ZR/0QK
/7fFA5R5+qv/0omNU+iyxOc/AtJXd7YXNPDqp6P7hqkJ4PYppxRTNlH9CD/eLUjlLUETpgWcGpmz
2gk+U4rilXqKchwdNKLpBNHfYcgLGNK3QDJg/QMRmvlRY5p/iBBDUgBCJCHoxuJkSbs1/y16FCD2
KZZ0CQYakV+Xs4MpwIvBHVGlAKW0eCuhnWbpWq7MttTnHs3DkhHYg1kIEcLj+N7/xoOjwmD5XDvS
AfSHbTpxoOIutCzjYy2RphUAQRFrS+oZmWNy3n9QRRCAHDanJU0dhrUkRCxLqbK0kZqRB/bB9Soi
rtQ+0K580SDwy18bHGBaJDYOQ6QDBX6eqyMpWRYhmZS7p4Y3vqvs+08MuuqNZFoUCeWsI/4wcGvo
cFmHbBORRqHWtB65Fe0EKkFBFhRaFF0SEuIqmh+3GggKz+PGlbG+LuopJQxI/h02ogbaWwUaHsA8
ejgGlRN60LHqQm4WidCOBjk5yOZByMIbg7QHZqkFzKw87GBrK/FEEM+2jPID4BKCeyk/CEj57uNw
j5VKKE5zfrVb7oLMCK2l8GvnhHI+jWejoyjVkjflRe4WejWFLEbk0B83dDrasF8vUr5gBdCjO3Dk
MmDzuSaVYVNcZMouri/6ddbu5e53Rp37jGxzDqfJ8w8XlZoqajqhgGU/zkaVCWVqKnzRatiTm0eA
28kqsVWRReUGI/w6eX2yCk2CQGRJ/g4ikcxywSvdl1afmEQmk0YK8JR7I4w1JRBtwasKNVaB0SVR
l5UQo7cFbeQCzY6evmR/wm9a/P6G7OiUxNAWSJk/H1XIPswaQ03bbLxmisJNHrTio7ytU361sdGN
xhAIoxaloLe/n9elxwVumPU8OWvZe0CKlRZBmMvlG+CFmPyTEzO6Vpfl/vMXdwKi4ZZI196cHBse
VeL7dF7uwBSb/Ov8CyjIIv4yNzaY5uo7R0OkxS6VTXWC2vqFgYjs9HFjDMggHyEkFAsnmRe6cuX9
dccsegJCMkETSRaDXsuuU0Zl0h93JktLI1lCstMCg8dwKtBdP8sJkBpSoC/jTGOuTrq94ZVt10SI
u3gmT+tGGIHuVyNsdaKXMECGPEYSEv+vEannYq8qOIr1/WpSGiQAiJoVhcIcDGwgjkt/prGeZ5hf
zIQuKL2BlotaX5FLotXQK4Ob7YDW/d0HP4Nhuu3jqTkkturjIu8VaC+LlCteaSeCkaETV6lMUJdo
DpBut6yuqb3+5s7jwa12o52gvR/2ZtLXPX73PjtQ3xpmUKd265ixS5domEtSiUyEA9B7jEWV7l7N
LIFp6yRo3Qms3KhND0l2YYr04DUVhCfJ5jbq43atVVr78lZTTN4pxVdp/9ywsE1Bdmqi036SgDy0
k51Plk4/TfINdzvl8DTUwd26h4oncfWR6NQXEs8u8FdINVmHClmUhagl7XA2bP2l79WxTqMqwaE1
2PEXmCGxOOEnhiF6cbDeZaHmUs9RmwydGE/XkM9rVMKaPbHv07TWKDgNI+g4acJ9h2cttgB5umfY
AqLtb6nGEiqyHgxVC4nEplTKwNgifM+/Z34vGeL85LtgZiU8Yf0pyfAxBfsRyWtawTb32LfWG7LJ
DSD3DgEliv8Q1VXPQpJi901mxbP0LxotpIwv3uo6YrDgnuAPrGWZLW4f8jx7WWwVIpZE6Hbg0MEs
fZWLr2t55mbeUfobSveUvCqYLZ+KcIrg7YSK6ekKFuFo6y1RCt8zwxytyMBwoZY3yCULJIGAZmnj
MMdobG4deB1ZGnhkY4RyKpTxzUMO49W2eUajIbioCaaOdIhc4iafvZtYEgXnKyRy1cPJk8uqI+4+
IcEBAMsncGqaAGXTXLZ44tN+imqvM1aZzl5LUfElgbfLkdZjQQYZ7QIuP8lZYvDNwiJ8Lo5PJ9Gr
olEVTyhDbgupNtna+/xqcYyGVOSQQVSVCKSj8H8MRLlo6zuQa7qXSrznHVIsU0MKshBEXVGB/Nrs
Opusk3/kFUB6BNzf3lWH4+93kCrhy55mji+uzZTzcIFyTzoYpxQac9GB2XvEOE8SmX1e7hi0bkLh
Kx06QrREBT+0erPX/MqDnyD34h0LTiVb2vWNxjQ5Swak+4jYu16b/09Tvntn0i3UCwTNkb541+QT
Qm+FzAQzI6fKDNIXvWEPVbFtEa34f61+NKdqDSW43PY7Vl4f3f/xdiNjRhGzhOgmj6XJklYrJVcs
3Dv1km1S6HFk0jCLnmDAAGqvChcgzo+3FdVvV6eqFXsJVxzN5RxjNd/Cpa3tp7nRuAJNzvwtAewH
VyIueCJS4uQxtx9U3DKIIObs3+fsxpPRO6HmFzRl56CbSUllQpGGQXUZ/kdBCm5I6tK0VpSFlX6G
A8VwFPx8V6SB9Oh4AupBvZc+39ZtGxEWM7K6N4SJ9cAuPu7erd39y2gMvI6rgHtIosZq3GeOAZvJ
hP43aQVtC73WbQADc+KZZzoSLXpm8egFPHPoj8ClnY4zN6sGt1p2nXMWJC2kX5dKMWq6V+U9IBiG
t0LrA0qtid/EwmGet+NnjIy+04rdbgteomKAIyrNZrlUyJF2X/QRA3NA6uCFwidQJm6tlNFuCPB2
KgN55J37l1fJpJE0E0XKBFYIDNKHa5f/vNfQJifi/kl8m+QVJ38tLvAvKUeGKsewHU0jl+Flsju9
Jj34b1TPeVC+opH8AFYln8bzWMVSj6UrMoPPvBpjslIBnuyObKpJX3aXWKeg/+KxX9tl4WTugmQq
uW1xOzebLkTYka7nETPx82qE9g6VfVat0YPUU2Q//9IdQOc+5oalLLAyVqvoX7IUu62OSHsF9+5S
C4HARPSN7nJG7gNEVhLo27AYY46i0WNTHDL2+y7vps8cG62wHo6rkg780InjQCBFM19jChwH3UdZ
t3haqD74PY8tRnho91i0IjZz9IplPM7tXnAeJEpCxXEo4m+8COtHyaEFKhcxBh2mjFjl1gB9g/wG
5v/tR5hVVDzHLDr4xu1/KuXZr62+g7BKbdcN89X8foiOx2kkVBfGlEHv+KcIj97QTNIrGxiYGZXl
LltPtqu3OLorQCK5UIyQo2slnTcZ320OZRnfRAFWhMqLNPd6x5kdBGzivmcwd0KeOQFkxIzdnVEU
4Dh1smpWbX14OUOpdzWU6KQGpVDlKnp9fr6APmVqvJPLhhI5iyUKuh2Gq45X04mYJZK/ueqhAbil
fWBKSKoZkorfFweRfoXv6QbEMXbSspv/C126DLbnjF43BYAMjH9pq/LTHKFOHXl6ZEIcB3MZzauY
h7PQRAmVoZFK2Ql+ocEDFQMyOS8FshRQ357oRHK/ZFGq3rv4fttC/Ko5GIsfxQUVVkmiboahBSQ3
jn13VpKtY0KIQfcdHeNbRFCA8mU1dQsL7ohs++l44pzvv9PwW4BoZmkQlIBuv2nYfGmL+doK5ZAX
e+frCa/JPpjROq8Xo6p2rfxYBZwrHyoCaq+6sserufztN5UaEBk2Sux9LF6JwpVkx/nZvw911s5z
CDWIsmyB+gLn1+8x74uQ7AUOJ2jCVFU/zCBeXY4q6TwYrkwUcnlCGU4j7UwZM3NWY/itsjbSa156
91LOTlca1a/oSWOHeZeL++BY6NC85au8pKC+XOGreM5VVsq2G7MIRrJjZn4N6SyD4J+UWuAjbZT1
kANo2mpklOamGF5mgvw1js5Nb5SMuvQsYGWSbo3dvws+ixbT7wgK0mnfu9g+sOBokva1VJ7Ignc9
fwh0Sgn6XGHhBuauY7CKo+7nR9/5SPMrUnJ7Z5UdzELMMfyP+UBtG3QuNIFza4eLjWBa0u6XlgOk
yq3pOXq0hz8EQEWudLxtIevn8FH71Zk4KzDipr6lkRsv6DKlOzeY7BFPbXmIa+qy9TGOxcxe2949
21EEvOGO6hElZ9iaQxpGpgRq6P1DMH+PeXHfRjT8JMepgmnHKiE7ras1aYr16ioAAassfTCEsUeh
rzu6eDxW47bkLxVBuwVPKVdq58DaDyF5zf9OQ96hKTgOozA5df6nG5E+rzQuiDxNNPoC6Ws0v8FM
SdNXyfeDLTIi4LO5JN1GkJspWWQFla1K6jRPKibKK4L0I5QMomqsypZHV33gaWnyeioSqY9MzvuP
jJLCNq4WFbaelnD3VU6HSFEbZHWbUKK+gbS3DZnGSn89bTFdZJv9IErzOFeKo0kHsN18W58FIsqb
Ggoh/1MIKZGxnA/yKxD765gRxSlhO7yV04p697DapPFoT6/TORn5fa+ASRLdVj7g7UVDFYHNrOBM
wDdqvkXgdT8WXFRs6Drhu3wLZtudf78XERptujfTiw5BAnWodaH6yWj8OkPLMoETpSObMW/ipHy5
tkBb5GWuqfe0Zbewc4Q85P2ggQWHEMi1V8fh2MTENU1Qm0NKaz4f+3A9Vq0iqKLVdZWPusMSXpLD
LAWAaIshPJBy9Ixqy2+3CJmgiv26D+WcLWm5mb5FngHQYP/b++zC6kfKp2YJ6I1Xa3ZcGEhycvX+
jxWeypDCgvNMITaHe9oliVBULa8y7sSOMPLEUj1S8iFFYGq0OMYrLtJXfilLUlEgP8FmP30gUNoL
v30xlyplPmECTssj28qH1a4Zb3Ba8izb4vIJDR8WICjBHb73X8aRpSxujmathUovwZ9jY5dbWgIB
XLEpwj22zkaC6RgLwOEUkzmraAvxB87d0r4DT9+FixYvfVKcrY5ppzo8QXISPnBaZzZGuU28IZfL
WlkNuWk3XNDEJ4+zSKK1mAcJnVhhcobla4frgIKWiA5GCVSi166COSC2Rdhv2UInc1uazu5ePTXN
6KpWi+6RQjbqr7sm0dqgDZADIeM3XKQrgwa0GbzkUB5wnLbgkwbiYPFDtLP3s42g54PXENEN/VZ9
PEHFZ79kyzyakmgZKFQn4Q0qf7RXQI9nFYfzOXoNyIvT7Ngmx1Zl/SXCFz1wABU7Er5sgntoERdG
E7ucfoNSIqXg27kFighjg1cIV+8K3ZQg/Ec6qUz0OIgkjle9kcMW6HepCTJ6jZSHu2JLQEuCKhw6
V90SZRNbi5jsjcS/DKIGz2LST6wiFObVai7XOLdEqI6pdDynFZmwFPwBX4YVWPo2gfyFqIpmBLPh
kJVXRcraDBaf9WWfSy5oavAmYHGrf5cCcH1VIesWuokIrahut2LnqbJEImaJN+rFbZ6MpjuEyuxC
RSBte8H6ULwBB3bIsw4Ll+n8aTrBR3bYK4jtkAChHlqv56uSM2kD1+XskxKlMdMghdmmIbWjWnVP
6neBfgy+ixHc5trlg3aaoP9k3T7UqkaJeC4ma1h1cC8CUp++9SdTfTJd/sZoWa89tP4zz5tqs7z5
uh3VGmi+BtdceKoe1yFGAGFLGbFjh3/gv61SiYaLBYBPG05C5xS3RGBmF4u5ktRX8nDOUBQTQX1g
e0zsH64O16T/+AfxTCi6y30FsDvdyVXfBdb2xYOj+q+K2cfYvmLcjEM5wjAWGmYqxabPoru8NStx
c6+M5ecF762Jhn71AoAhcOX82INvr3OH5ofT+AgHet9bwqdsx+cdmKBhVMZ2U3k+F8f/J9XFl9/Q
AN3YiTdJKvR/ynQh8VIYkirxCnGHn39vdwBJ65tmKiGo2Pux+571shEZ0OemohBFuRxev/V2qwFA
4weINR8vuLCP7uasfi9VNQm5drmAe5fCYry0viYY6+UwhaR+8U3mcKhIBnNGlTlYrMzdqybfcgyO
oOP/aBio4ogK3bCm5hyf4IB7vZevOX9UEyL4iCr9LqwccY8UnaGfcRjhaeDjexy03NFXNW8qQHNN
FGbk0lKNlG8RtboGw/UaiFhBhu/JIb5Me27AEUGyZ+xt5L9vuVE2xLQvsyzssixBEmictXYPwztj
Y2ghRQYLnCmo3NoEKKVLEFJlhkdGpbF1n5Xwz75bhDTnMojoOOSfHvrZER/PaSOMcViBzqVVbwk+
UVVTHlXYXoGytjkbgFrU70lopma/PcV7t9X+nHvVwlkk9Jmj30iY3VZgpUgveDIz7+PBc5KTLy8l
Q1P/QEqaqOMpmNKNBM8/AcfRk0WosP/BS0yX7lN+LLUGTPrP17Ipa/jAt3FQyX2HERwLqy2gLqSH
l/1IfAshzkwfocQl+ARCcjredqoKGo8LaJ7cvyGcSkkKJXIkJ0PJJj29aj3M65pAZuT2qZLpAKzJ
X9DlFpzsqPQTdtUT7CjUA3THl9zZrkEdckHYdssEsK2LSV/+w/KX8vyKDsJny5ZzaJOh2pNjPDYO
00/jFonC8ghW3lfPhPukYR+fNoBJALkWveBiArqT2gsbqQ0GdkXqS3GEZv6NftHov4Zx6mVHVLIZ
6qIsOkqumQFPjv7vRvQRU7vkqCyfrR2PyqYFU0X4WVEUn98D+Gm2KrnLSQIVhUy/NWIOKd4re8bW
2gf4h4foqVM80kL/qSnti/OhbY2hXUJvUrvApYCMaihrq84W10Zl/XrjOmaWedKJ4lWaLr10Je23
qRsi4LOtVtRaVPvjPUvLIwy8REpSM68jHlHnebbCHSErW3MYobk7lhW9URFydHcfZkv3L2dYiIPb
ZeMBEwVrQcGgbj6Lj33UZC0UbfFUiKPvlnBxefznDusBVMN9J9omyrt5xTbqqnaz+W8dQXXjbCk1
lVocX7WjUoBZ7pLukGCqc2cV3QqN04XNG001cOOaAUUM3cLG2+F5cA6zrXMJzkMU9Cc2WETcQ4kF
QDlt7elESRUYIgHrALuUlZyeAjuPHH3SUnONB6g1Lf6bsL/Ve3BxG5JqiGhLMDYWsGaF8cH82Wsd
AVaYfHvYJTCXZi4NCrTG1lhVhRNqtHpzVqcquRhOkgMqlKi5YKXWei+wDST1kISte5SI3GYy5Wr3
gIKkEGhJptrXdisYCZ3I4jRIGku3dD7P7fz47v4XV0IyePqVc7SAGS8+X0MuDyrRdgHcA8sivyr0
h8BvnNjJYljLyw2F/ImPeakj48yknyfySRyAKOHLu93nl1aJAepk64Y+YfdC63tBVzolS8qmUAhX
Gkwv6LbaoHybBRDKm4xrSBx0Lfdx0jJVh6m7aCfubuokGKIptgY6hLrTXKH9WEPtDtLZtgsPdBRN
2hGKgCUu/6IA1yWEWIf4IrWXoPINqAaQzcSRKbR2wBvu3EeTdpQ6jaMKisBlKRhCaYrxV8QTRzUo
iY81xIjWLrKj8sneD1HVoCXHr25emXiZ9KvuNrGKgpovms/hxMf1SXrMvEexDq109KZsoQCFRLmC
4DOPx4qu/L+TOPXN3lSjmbTXFSRkmFhzquJvchO0cg6lE+pL/XbG/isYO3+N8UG7mGWS66ixDgbC
p+BjzahpXUe7tnHv8BDAHIOC9Pn+s+XeYd8SuuOFTxd6eDkJvx5DVMXAkjgOCq/pjI/szdt9BYUD
sD8Qa2YnuDfTHbgK4CD1tn6r0ez1ITdbOeN1MD3CNciOBcGPnX+LehgNpmzNlSWsrc1y0im49KBn
HTf/I7yMvqUsm/UP1VQO7e2IvutollyfDu+kD0PbkG+eK50UWmZCkET901QLRLex5etvQLDOIhMB
ewugz0AP4wULaDGF1b8hq+MVceav8y270Ijaq4L7XVotCknt3Apmr2RAijs52zQdVNxRqpbhIEoE
5EFAPnOxh6b9j8E9B06PnvWDIR0RlWxGFEvmqyxY97GDuG3lVh7o+lI+AMnowYCnJF5SwFufZcrr
qzRCXmoYXES60CPdmaYU9rvnsxCSqAi7SjuPsw+SqcFL7bQAErEBUrUm/3Yqu0fA/Vo7wIYuj6MS
nD78cVdT32Qw3UaG1luxPFkEz8v3l6l3rRDHtGHs8jaV2lPffZGCR1xHpQBzK43D9CN7jYh6OmAI
Ic5obYaQBEFF/w8Jqj2f/CIXUfHuYt6nEdnjZTDzRoztFc+TgZT0B2JNPk0+cyFjrt80OLivEYUQ
T2w4EBOY8UMV4jkQHLdBQZ6LsREDxsDUlTKIigp5o+GPRUuBGu5O5XHa/nuUUmvFf86RNWoYNXt5
ZEv98R6iQE9n3o+J/1uwfKi5L1SQ62vqOeUQ8fmmLyZqd5TxkTT74MAuPzM6CFngAjdQ5ULGKrex
/qa2N/YuycGNxSbPdSr2U86s6TSbjqXc0k8E+vsg79ClFFT1hwhM3fqmLK8FZDNrharA5rbU7imr
bJNQXBPKkuHs+5syh7lZhds0SUEaHENZq6bkbQxTW98RrdfSpoeYN/s3MntUmdNiy8kMRipuC2nn
W9jI4DCi6TrVsnK1Af5C3sq0GS/8sW95bfUkVJ/cHcN0WO2AwOUBKti7JhI/76eBbsjCpeLROFbL
SrNEPaCsGZf3/IVGxPpcGl9QKwOTRxQL27pfozakAzrqMbWU/xLC3WWVVsYnSj0h1iIpmUfTa74t
6VCykOfFiarO7RBmfEQWdLHwTuCJQXKOu/v3QeLLI5DjWWqNOCANbFZrbBZRgGiKnaWbPqlla3Cw
cOF1AaphZLBLSXDtAJpBG+Zy+vYxpO295gK3M92M3ApC2/JGUOwDx+tjCcUMkeONXTtx5mN5XH1g
AcR7+dtnzLeGAps9Nd8jRhRz7WcL5g63JqywEOQZ38jSuCDC3rRoSLje71CMmNP0heWun9Gk9BpB
bkaMXdGntVLP6O9J84GR7HUmQownH8gw45Hw70ICuT1bsjQUPZ0eJACs9aEXyMfO/47i7T87UEk4
X16aJW3NGABJ7heJ+vxmQ6x7fpVXGNdApiHVZEwAru9xZ7YzvOI58pLfGWSUcTYr8UhO6kLZ+ZTu
fRgB9KJR69+Ss0+oaxUpwj7ToAghU+Qq8ig6Nnm6rFgSY7JoXclSUZlyUH59OVQP1/h51wdx56Af
C+qL2eye53J8V3+AZg8fnIyoe/MHB3OPMJ3Pmd+h8NJwn7BgUWjMsKmqkMP+WAVCvnAMKmf611F+
++fztOFv/msXzTnWskyWdlegOETUf7d832/SKvvC63vAI8RkZ6siloTXyb5jYpWSUO2W6xwa597P
Z/jRcWOmPACihBfOJG0gYIJhSglNX1ZROOjJTbz4EMIL5fYJ/80CwJkX/cS1CV1QeKl5cxSmUSkC
uFKM8zYsEvLNrKWEepvjmyQ8uDZ+qyVi5oJ5kmIWuZ6fDT3YSc59ltcqD85SZThD2cISbDzMGe6I
uHfd1QFO02GSte8ByxOkGbu2s8Wd5jwnpDBCn9060gb83kwvmqrd6rk4Y8kBgmpL+repHEspGKgU
C0ju+z00lr8RbQEDuk0nBi5s3P0olrIXJtTP5TrPc7fd1+D538FpPU/QpnXA1/XehpBfakbq6dJu
zejOZUbuWwGISwQy0vAOR8P2HH5hyHlfBB6RIbXHQLhnOJ+0hr6kgv9SrSnGeLRY6qNwb8zET9eJ
xJvMNEHRmSxTLFrmqXkb0t68X4cNinDMUMysa/WHDPa6EAUycjCCZ+cOZNotTlyoa6jBe7ksrgVT
N9H75usNmVrP0xwS/5foS5REZJmtC6rT659fJogVK/D9dhj7WwT99e7N/T+wIISr+FhjDr/UdBr/
+WRIs96w6kPsfvbma9LzglvBy7PwTbZ93sieekLXtVvXACqi1N8hH6aMPEHAgqgjEsWGnsTiv9nn
106o30NvT3lQ3SRQpdbzymjOU8XgZoOPyYjTNsh+4vUbwjqy+FSuN+0GMx5A/rwfxoriRzADQwD8
nN/+mlvH/35EXXyOcrisayPtu7pPyzeRFeai7VQWW3uVrNieTyGYpLtd5hf8mhDiknhUf4tld+Mn
btv3uKkWrF3kS7MSHAoTcsRoVUTIOQsROopX9jM/aBzGG2BjwqVkfs5LH6D3cs5xlNWNX3fk1IgM
XT/Q1U8oygNQZhEmuOvqTJ3aTuQkJN/vyg3xS62xbIvOypvk42SmNIeH/aLVPDjTwSvRr5C1yqT6
jE5GUiJxTpL288oZn6/W8N5OBKMUObQkYeYbbUuLDJ+EIYfiuNGaQvoMRLdi7cGafptTqEP9RZRR
1brtlbmKJQKQctYVFoyTXYM0GWD7iYVd/gEetOzxTVG2bjDPYPezrX4KqNSTT+EYEdz0U0N+2bvn
twd9FRISRV5A/EHicoIxZAMfisK3C98jtsNT/sBIT20Qi8D/mOkZ8BVEERUMleQ3Wxv9Slh3Fi6p
dj19x7HLQcatZy2ML6M1CWCNPmVrt0VZHdvpLaplHtmr03qNxHPVXyTXuFG3eZz78ahz7KynqLmN
+YDzkwUjLVejGu5Ivd5FUjEyyjuYGMzZWo3lWaGe364QrL1t01eQHuxKUFBl4AQ4KxJJWt7ANSsb
OJkAspVAccptdAonxc3N+moXP8vln3Si3M67vS/YKYj3hylqMvu208by6cR6CDO3/NG4hu3EVkJf
hr27Trgjc4elTdflJji+rAt3PvnclqjIQQ8DmWNT8sbgRbcDBHOBIGTOAG75sNhUMDAj0VXJmVpr
vy7uu87Pun6Nq3DyggQe6DL0/VFq30u+O5TpeUjQdcCvMA/Ctqfb1xbCzLfbFCK3GfRSeDcVS8QU
VAtghhzkS8Qa7LJpvH9J8E4T25ZJpFQlkL2KRtmmmoTltWDGWn7gbzYnXmCXv6cxTBoPFBUKmAGs
uKM6yY2/kPudFYrRhcFWIC+2stBDgPfIM/ITcBTOQXqjPZEV+ZLNj73iYWn2v1fiNewlOJ65sIT1
oOX9ff/LXCaOY9I3ee+rdJrDJKFazxR+zTCY2gCNsZl0UiW7FS5Laoxfg4p3sWzG9Je4ZZqdDG34
yQfc/eN3a3nJO0/rPs85fcNRcN9ikXD02OqBS+mUuDc0OgsSJN/BQM8NIplzT3rmXaCTMRs/fJwR
W9ovi0Te2AEiHbamOQMXX9YWy9t36bp53aQDgoQZs02tFvuOC018Raq4kPK6BaF4TluLJEVsdY+0
hh1jFOjglKHWzpcn/uFsIKax8tXDsgnSvPwZa6kk+gDfLMO50NdX2YHhpgab0m2D/BaorOs4lQEv
YHESJEpoAJ1cnhSilByEADP5jnH+JeF8ffZ/5Z9qihWT+AbrNQFNe4ZalVPYrAGEidSO8iVd47CV
lHZBswepHsq1nojQSzJGE/UKEUQ4hp3O9Qv7NNZxYrjHxTkI09D52TPjq7f+p8ay95IOLTKIDL2V
/0ZZgAbFm/ZRQtwIT5RkTuB4kwRIu4eRiURi93Jcv8Hyp8FsE8tHm5qSsRmjXVep6s4HmAWUx+3f
UnzSpE3m55EKCZe7ZZAN8oB8uBqsK9Dfuam2btDXBDF771scDCBItIbAv4D99rgmBRg9GqP/aP9u
66gCoTY1jHY214ECfUrG3k3SvulTsCkDY546nxHPI+Xdfi8O0NdqmsnzNzn5x8BhoQyXz55YwRXs
tIbmH+1yGNyU0COCoVB+6bWL0Rbm4tb3Ft8zQufdqrNx0skFmbH3Myx7CSd3d8t7TAkCAYXwK65L
6NiLTAvhUxE5lMgL92vE2CMKCumLxM6zjkrAWpjxLwtW2jpglFx+cg25EvTlopeTsQE4iM8ZoVQ/
Qgd5Kd0fDtYYUioxyvvvnoUOrfOboBuKeZAO5Z0cyYkEVzX20YGGTzJYxfVkndg/3SWH/V7WapnV
ETjg7CHl1ml19xlokbBc4RZHWmG/jBPmBUzunanysEYFQ6R0X3RMuq0qRUluDVkWKXo9fiETIZg3
4XIFsx03UhROiWi0xCuxHWqmoyfCRCa9UFjjEsB/btcv0DaZpfHnFeHWDh4AXJwY5/G2Ez3WcYFO
yf5iGTECIrGowujsD/PympdueWAL+VmHk17c8sIxiPtxYUQ+lDXNjGkEUzwZqB+aDnNczMlRh+f7
SW4yYmGhAsSgSowB+4T2KF7AE5fLf5ddFbt7xfR6XqqtmQOaTVfkhFC9N5Bz2nIpUSHNUljIS8Su
cTdjFRtqi21vO7VlPz50iTrk8B9zXlQzfJ+czz/akhg1Tgen98PKisG6K2sQWggGf9I8N1k0Na7T
tKOuRuo47UNHvbKMnXG+nPEulzGi+o2KRLhacRj90+KumQM6srZQw0JOduxyvrYuzcIJga1cmJH0
EPklWoQLPPmaEci8hwgrZIf/hZkcSVTLa8T9u+RAk5myuqr183YKlN7S3luq+uqy53cmV0lq/uUa
ZCgzxURE7OVgvLbLkkrY4c9T/fqCE4fS/mVVtelgDNqiTLH498DSZjketvn7af6z0NMmW2SXv+Ca
AnxfPyOYw9Qc5vn1U+cbDDmqQCFOqGuHKrgk4/ayAIsyoBPBQSL5ULJWHKtvSMnpdtRLc5pK+IbV
t9soHgH9QE+O1Oo8HykSjStADLA1eaOpYo8fTzCtYvFMghn6CPIL6DAIZe/zBcxBtWjatCbiTDV8
jaqlAWdtu23MAfpMwx9nZ1nwve/jcbvvCWw5xW5Dw76d7ksiqdmTDLx0FmUvdlc9Ez2AETz/eZjw
gxSmMob8bRjaQd7tFH5rYYLl8rXivmEvybOTUDoR45uwdRuBiTz+41dZ2EfSHR9kOxqPfOdbVzQS
clFarIiYpjgQ/sdyXmDGBVHEeocgQY9ne2SJNfUbobqDN2BXqur3u5kUJxfwnUWKkwk97KioByQo
o+fi/rtLxnBS0pH3G3qt+aug2mXWRlj1kpZNNypDt/ClULbww9ysdltTWJ23BEemGrXuVR+tQ8nM
Hbih8xNFZjdmiQCMEDstXzxThNMIetYZ1MG3NzUJSCPITcWJdRxuQDnJJZcLSdes9ZHwVzPlqRA7
W9zt2TXMreiEAdBfSJofdbNSV66g0PkJmvfdCLRS3rv/l4b3C0hxHyz62V4QhQY1OC/ZQOus3S53
C48SPlTph2GUI7p2GaNpT8xYHFx1VZg1X8S1664scKzorVkS/RiyqagCzih5nmZEN+LTLvPzEbw0
oX3Y+JEXt98gkS6bq9MjMGav715h5UY2GqOQUIC76CUTouMXM3oslbZOR9PLHcyl8uTElsYt85yH
yOr655FFebUdnbiFyzKrALcBQmO5HVFJ82a/tC2CMBJcfl74DP4Qpv8vdH6dzByvGiAXSflGd9oP
jK3B+CtVfcZdo9hBsoOFQSCjaM14FRSnJmykHQs3cEgnFY7eaK4LNT7aAT7rKq30DYhGxCLhmffk
Y8GLh9bCfeRZECYp2G3HRcEBbVEwxp0JdeIIokrc83+X8oeEit3AOaALfRKdPLwSk+pi3WUzxWpQ
KwXAK5SE1C+QL3hEXrsNv9Eq30f5X9C8kgUQqnmQBjjEf2GIM3TOftRrTLPWm+IV2A/txgb9tu4I
XHlnkTruBzgEXRdvYil25zNJOrzpPsZp2JiBYhleiq6yeeMRbnswlrC+Y6ylyVx0NE0dZ9Eskvo4
c7l4YNnClwxQR3o5jKnxOPTcqEr5xHTjlegR0AKK2ZD4IQcXzlYCTpYICmYOTDVDa4ztQY5NBDxa
NF6yiFSL6coDjHTybJ12q+P87hdvaSuQ2trmsZpTrtaF5MmuoygOzXLaYemP8MLBUqvVwUuXRJQu
DMndXBWu1SwAHX+cAWFGj4ouYiXSUmzcBnrSgQJtuUY4hOHeRwMPxLUHAZOfUQiOmBD+WIIML6MQ
FwN8i9Q221ePzf4eyrSk3c5ZGxoXJ983lpLuO5WkkYv6RDx3T4hf/txtbC3EPtdI5LLlBLKFYQt6
J+1ZFVDiTtTwKLj9sz0lyrkL9LR/7tiNvu1vEvsD7wPpbIiB8TOCH3toIGkqX1p0n6L9/Q6SK3lj
iIpGctWLSPrh/6A2FnoF/rV82NhqiuyUGZPwzA+aUL5Kx0ABvL67ikdj1bmaL4ZsPt0r5ro5azf7
tMBv5yJJ0OsK83kfc6BdWAHSLxYzx3q3kz/c6coKkPDzcQkDMWpOfoLzcsU6ppxH5B4dVBJ1kUiA
0nlIJvhthEaKls61MUYGLnXEGVlSJ0UVz3cYrGVqNXHV+sEv8vLfOGZK585AfJVEeknoo9lfe8Sx
dtjphyAyHLlhohWMZAkD7L1bJ+wTyJ7tJR0ynSn1xu8YZtsbZS8zfzr6E6sArEt5AojTy9OTUFnf
f90OtlDaW5DtIYVEn/C+HWmvWryAzRoxiKvyUHof/cAWnWH2pcXCDuOW5b0mOYsmd3zj/U/qqCBR
z8IRylXp5Kw9LoALlfhJm1VVTC321FdEDkpcwxWLaf5gqKIK69xUnLy2qqshr9RPwEYXXg/wGJkG
Hi02X4msevhK8yIBjWDHuqRP49anZaykqPe1YclvCq5H7NQpFII190cH5LHu6WB3ETmjtN011wRv
AoPm0lNTRfNvQMN9wphbQGaiOzRNeX7HFokerL1GFI13uQ9tgHlYRgDK1HHa9JhMimWylb6duIDa
CxRi/D2MViR0tbM7NDyEXux6+ULbUtkRGylOIEpmL9pb4al5e74Xz6NvRBxNMwNUAEFceJltt4S1
k4zUVcfLz2pXN3bnzspP7tggw44y0m3mn8WBAPtSdmRAHEPV/F7VLyVCMRvhl2JrXHGC3oiuI1U+
LUi7oGrnFbj8K1zC27tnSps3X8aRnXSjpomU2xramrrIsK8zp6tXmD5GUz0t7qPBpgTDiE1bvK48
7h7XziVHvXv2RH43tmqyHje+bEsqCXJo6tDVBgUklQI1Vc+aZFUTML8mZWNZuyjffMtg2wX2l3xE
DGWgyUo7R3xhbQZLQUyWFZNp7SK7pELIxwwoOV2+WZSzShyBkAItSxpj40nY6jqhZHfcZYWYWy0X
yKmn2NxqFW4LEsV8D1qESKv0IS4pN4MQoKDeAJGX5Kj9vm2BlZb4VU9Ifwlb8fkhwUu969XWOuQ2
R06MygxhlB0bRVm5uKOulsQm0k9BA4oSFxMHwon8nT2P4UzWu38rnKN9m1LeYY4IjxzGS0O2vOiD
+52tiJsuKrMMwdJH/2OlxoW/YJABXy8O6Ba7qggL6Cnr4tgzPwSZgLPxiHfMn/SkLdKXJFK2cRL5
LUNbO9GuU4CQlA5jfDobFD034sx1+9aih9cVJVkCy7MKADe9oLrVmGHOolzm0eLkmyeKWsW5JET/
6eovSaRY2g4r3tdCErEWW/QWC1JlOdt61iizO4nghPQTCM71YT9Yb9/sLpK1Y01fMlwbU7lSBBPk
gAmZkrmiWXjDLdPC3l0Iexgg4Rk8bt96AfVxQJK2A8PE8KLuxxlDUEx1VVQ4WbizZALeTtmK2lqg
Up3F72O+bNeNZqZOfsZE9thM6VDo9qCroZB22QzPiR+eFgQ52uRMVZza65cjVbYnS+lVU3vaRcNA
+rJcoImk2FIflEl+kL2t7QkYFrCRPG6h1bPssHrAnAAK+ZquAv0jexwkh4kcqoxRZ991G2bGEVcU
BNCalQOgzp+8Kf+wuaWPQGd3NRFc4PCTGAnjWq4IcfSqwHNQ05VN/IpJMt/2evI3kSJmSNbCYRc9
/6dInmCEOil6QRnjTjRwkxWUiIa3Mtc2hVv+YUJEL9NSkFQlvhRwH8N+IPOdx9IYM9aYzigfVhgt
CzMLV1T937Fol3Xn0rye1zeXAgMBXh9hjlFZZ2DucvpRhXUV1mBAwqEv69PpPNgNqBXiwxr3b2RD
EPACN5C9Rp/wp1pbE6OhKv3nsm2nN1npK1lUqZ3B8pY0KkcUCS9OEftBX3O6vaeII5a7SoHHELPs
y9Oa/xr4hEeKcIFXM2TkZVjXuS3bFDhLhwR2NIfUT+pU3dh7dK6Isrey5HqiSDqJNcTlS9AzFU9k
PuB+ppAiVmuYGEKhrlx8HB5YmBX7H8G/H4wGNw6XwgIcVMqTShtaEl9vY1TcZcsrbAjg5Iu153j5
S1M+tCLxOXmOljZLC6pCkLkep4lKPEYT+wfCyNeT8ZLN+4ijVkmXDYLS486sZ4BXlC4nemW9GqeH
qeoYPrOVT76iFoKKL+g8kPIBse+k7Y17AndpAL+k3jMu9ML9ZT5TXHTcG9J7OMBSO/PCuAlNx+dm
56Ugyf1ArsSf+ue5BxAMFsMCKQs4Bd/+UtIhZMwc+JsEWrHonksvuCVjHPx45HAbZVp0dfhbf+0z
BFL+UMqG5YkVedwScUPU0mgC4ovjMArkrp//9lYV8hwDcPbXB5Vqt9Y8jSPj4Rnbi+EqjPH/pyG4
pnkKCyw6peYUesC6/Vc2KMp1x1lq26wXM13nw5Cl5JmmBOfHe/js2iLOES9Cs+Jt6ws5j/xQGGut
bvpPca7nc5yQrF4Aqx763EWxAGOoP74rsqrzJYNpZl52N9SRb2NYxHqSZH8vHUm2RzVWPpzOjvh1
p2n//9/QHN8Y55aOfCRdLwhchcmQdfHb1stNySReeIq7E/jQjSYRoI+vCEtFP+KYzM1o9jlcbaqw
lbg1GXZOnsSi1ByZAId7R4LVx05NDru0m0sY9n9YLeBQoe+TjxDkw8DSfmsXLxr3gd55lVQPOEgc
/Rl7mWH9Znfny49TUI5u784KCguvDz6YHHeuL/87nBbd0TuEiuOJ6Foj4WMSXg1w89B/sJzPQ/E9
R+VRuT+vJaFET27B+WZRk23diw0ulDRRhH7Be36kOexXbjFiuUL1VNIcFDQyprV2J5oYX+DWrXhl
1jL4QtvspjrqIs34B99sFxa7Z5g3vnlsMN+ebG55TDtCLN9ZuEC4iXGMDya/KjKtL3gi37usBCiY
vEWjevotqqdzEPx6pMjdXfAgjkWNaGp8HG7zPYlQzLGbShSGBXcBIxyumxFwSwV2vi90o8PRQjje
Bao4ZfN0DvKslLLoL43CbUjNO0apxmU78RAUamOEB/8MrShGdGzsq9qZQ0HE75WgGjpxJ/qG8Ruz
sYW46VOW98UCQdbzxUQMQXErQNshSW54sJejVeXL7/1emF9FToKi+IniwxZe/oCqCgJiUGFlcaav
2AYqAPcFzpaLFLUJcLHqUsbbuLNUBaaIscKqDJO4zQppci7QIWrIpxBrABNmfys6V7Lg1shGhhYd
DHWw0+dNsY/HtlIJoojI7REQHWsUM237phqZJLYtRIAKjNB2ELR/QD99qtvSjdUe5/AYlO3OjhAw
kgxmegL5xaEX1B9CINP328KKhs886pncpl4Zkv6j6PoVijvGlEqnqlNIrSSsmseJ8GD1hOKOVeRh
m4prgFRKpU9QPnTR3SS/if2G+HA76ku/sqiN1cl/icdiQmroukFmY0EjLqBMRDwBDXYm/gooV4tW
FNWlSimB5Fou2MYK36Y3qpo+KcmteK3yCh76wJqxSXb/AYa8pR6ULT5g11hwYr8REsi+RLoEUHoy
KYpvkMebnz6BApa1XSVbPlrl2VGByWevsF0fJBgZEEFaruFXt4hL8t9lTTk8D+cG7zYgntrCiX90
MNQ9CqH4q0LdWz316/jLbN8bA9X4CqLmna7T1PnNa2Jy2D6Pc1p0RmqiGcqBHzI5mx6tPIf9kF8I
YzrBf4+SzEC748LhyXYzFJAdH+3y2pQEM5zRgDikk2rjhz7d9D8hKC1XnF13EiQO1m5XMHtj4fxa
RNA7sdM1i9mjCq0O8c1L14dftIqMneuJuFvM0AyRcySCdq1AqFWH3lGgeRRkRU0oMJP0i2KgtRZe
ljEJHIJK/mOAv/uKILZVhl15zRDzgFLvzy7pdQSvO2/3r0eNP248HTjr7+KsW9sV5ow26y82mU2j
cFsB8682s6o8Pue/sbK3CapRnQdtyInJrfdJVkQctsacH78rElegrlD0kgMdG0CGAEyzhO8wVSae
KhEo1vUgQf9WWE/NxaJeIdMHHqTI0uT7EUvNhRiVi+GOi63eZDIOBdgkfCRXsnN7SdRlZyWyr8AD
ZCJVVUisGV5l147rvJh2k488Tj9LLvIBqbbuJrC9KJl+RqzdOc/W/EwTcz578zfrhLYlk5bBVoma
7TyTGVIr9Ug6kjrSL2c83YrtCMfNYnhcPpuyZwTSnMLgWb9k8pOgPigF7BEx1IlIo6V49metKJK2
jKrS/Dz3q+Ow22LlqrgaRGkAajnqs4+a46AeD4LfYZGVER0uo8EW0GawBTN3CQikaxqU0+OFS+9e
EHqxBsmphbUIUg9/QBG3Xjqo2dhmk2cSLpFgFzEmjwAgtknj8JemDh+a8KEJxBBiebOh5+CIPq/0
fCegr4g62d6KsLMw8qOhGHVb35LUdc8sfalAiPougl6rlmu9B4ZnqcuApKGA5gli98wVVuhEaDak
5SScifdau1Q8OqzDQxPK4ATtdDOd/ypJ6x1bUpEr6bYS4wl+gi9VGbteN0sewiGj+N+cy8SPtVYU
qJ4=
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��F��g�#Q#�Ⴛ|��0���)¯=�Ә�$P[@�T�]��V@��W�D�z��HY�lHS3}�[�zf����c܍�øvP?eؓkEы��̑Q��G���F�3r�3^9Ra�"����������J�U%ra���xc�Mu�IIM�6���JJ�ǡ��c�BAvmo�`����Hb�l�����E��W��!���Gʡ���4 �L��$]'ͫ�8.k��P҃X�h<��5�^$�i�����R���Au8^x�����q��7G�c��������k <BnF����j6�P;i�1l��1^�����m͔H���O�k�L���X`Lӳ���5��}�Z��K@�U>��c�j�p���jme(�Lassx\α��E�����0����k��98�=꯳JW���������&M&�+�����-��QE�oH�.���V�� �j0m������fI��ɚX|��yW��_?|�%�N�e��,�&ݖ�P5��>��;͐�a�8.'�m��_]\�ǹπ]��jJ�5F�&�ON�������|�V!]��f��Ի�p�1n�Z\/�1	=���}Q��հ����-�w�v�VB:�w�\�#:i/�HN{�8�J4묝��I+X���^
jG��U���"�%� 7ܝ�?B�j)ȫ��,#�	в�2͞�|�3��M�M��f�-\=̞���b�?=�$�	nM���܎�A�h饟��[ی���OI��U�U'���'}����p�ss�ږ��*�߈x�o��F�χ%2��4͂G@��p7��45�%�AXX
Լ��є�Ơv����)SC>��q|�5\�L�:I��ɽy���5�`��BU�;����dI{�"V �F��atI����<m)\au��ɮ������T�<��	�"E��&V&*�&Fo�U��O��5��xt�z	�ԡ&]�z��hE.��e<"��*�����o�o���UD�+��J��W^�Al�\ɗ�� Ξ[}�&�M���P���ι'��E�<h��(nL�n�]�>��6ڜ�T�&f�g�͡��3s�;�����&g�1�&��Z�b*��FR�ۓq�z*�J�u9�P�	�':�$���'ؚ��<�강��VK��D�Ӛ4���*�"�K��E�H�/�BJܚ�-Y�v%OЀ_:�
�O�)���Ot��qp�*�7�U���t�����W߲����}��@�M�l�r��@x��z����&�:���#v6n,Nsta���	�.�;9�0K�U��*�K����I��`t�Ab���G�i�xǗ)f�n�S0~��5DJ|;�� �}R�T��K��͠KO��Z�"���܃��wp�SM�P C��(D������]$�Ko��'|��"O�?�r�b4g8�5��,޻�4P�!���מ��:v6�T�9E0'QWjubdQ��q�hV�����3�7Kް<�l�`�ʽt{[���_�N3��A3�(���d�j�lh�I��q��!�I/��D��]-#Lb3�����ׂ�7.Av�!YV�{��=q�c.������ӣ3�U4��=� �0�$Zy�r8�$��{�eMwrP� ���$���j8�:�����waQ�D_S�UDE�fm�JA��Hw�0�|�����l�pE<?�Z0K�Ss�����f=����4�g%�S�Ɯ�Ϩ��"��%b,�ξc��-� ����]�CK?�n��h6��p�9k�
o97��
�?D�Wjy�3=3z�z=,�-b���	@I0��i�Il��1��#hp�\�43�U��[��BV$ZƑI�aچdؓ>��)��2�x�>c�A9�J��>=�]h�x5yX�f�A����D
g"�g�	�L��TP�ӭr�21s��1⁰;�n�L�z��hA�b�ԍ��$�aZ����0�l̈́a�Ng��0�j>͍<��H#<gi��_.2�b*�8�J�9��&�z�.]��	u���"436�=��ek~��n�5d�<,t���#p��o�!��%����D*|�lW���F#�gS�6sW�x��M��.4X�Q@QY��HSC��}��/G2�F����?��|p�,��w��,�y��Y���v��c�@������9�b^��zh�����'(d���w�)���F�&�\�Ob����1g�P���֪�4)�� �R2��#�H�Z>�PJ�Y0Uca�k�r�3!��ZE��4T��0�����-D���Y��[6����k�Q����MI�h�
V�����r-0e��m�l����vhC�^�úm��G�Տ\�"
�![�]U�U�[iP�y)���{�@W~1%$���dnoA�Jvǵ~���G��fə����OB��b� �Q��Mv��QC!7)����s��$@�ztn[�E� rJ��F����8Pj1c�<�4�dfxk�5�.�'��Gޥ�Z (n���x����]���ͳэ����\ ��ʆM�s]�܌b�
����f-o��L�K=�GDu�Q��j�i���(1�v�iZ'��ūm{�w$z_��m/>F��Č|Bن>W�W|hle3P� ��LYǹ.�h�k�prVK6v��+�W���㍉�B���è�
b�aDR�nF�G]E똰�Dt�֩�sVr��^7��'��?�f�^�S�������g�"Y��8��7�ԥ+��Q��eri۾����n�Y��";�0��JЄ�~\��k�S^G�t<�pP�=%��n��S��e̫�vI�5{Mg�`-�DM��Q�I|_6*�0w�.҉w�,z][i!�ʹV9��^/Q���\:��z����_qwUfCۈe����p̎p$����D*�w�ao��Sޑn��@AI�@�2�;9e���jI��!�N�[+��[�d�P)�{:�e"��*v���M_�De����J�޶c-� ұA���Ә�����.�4��h7��j&LL1z3q�^�gxWq�\�V�Oi�"��hG7��W)nP��Hc��سވ�L�U����ُ;��D��t�MtԯB�4��*lbV@	�/�#�*rt���u�?����Ӹ���u��|��J�5i
���8dLa8>��ǧ{�S�a��+��h�΂��m'M�Ho?q���:ņ����H���k�����7���i��,ɣe}�׃�\�"g��{�h�g�Nڲ�a�wik�V��4ĸ���
' �	��\FE�S��4ܺ�B��#V=�4���4�k8=� �f�	����|w�xąA����ePZ9k̏���6܎{q�I�*M9L]ퟖOV�Jک��4�Ѳ�xI����A����73�#Qt�yeE��iY�@'p|v.��?=���U�9ki>�|�di��8fK� r����	&��a���;<Dm�
'?�,]QP(�9���M-��p�O�.}6�Ǳ`����8����b�?�z��/v!Zs���p���E?ɴW��U��&x<"�~�=��:�S`��.��5:j�{���K�1&��#ރpY���{��?!��{�?u$p:_�'� bPv���/�U%��`7+�ÖB�a�"*���S���ȳ!�RV�x���]���2�8���*w�A�R�T��'{F��%�h�L��"R�ˮ9�8D��@Lq�GJ��|�Hƕ"��z��J����M;\[��¨�-4��.g�2VlH�7��욋v��m	��i%����;�A��ւo���{�g�_�Ȼ��m��]n��;����U?�!��|8�t�����O8�)����z�|G"��S�J2�&�l���I_f�P10_7�=\s�#�� ����o2�8I��Z�ΏK���;ā�*{?،�B&�o�D�#�y�T�gA�"�-d����ԇ��T����L�F��N{0r�N/��w�Zn��B�$y��Ջ\�'��4���S�U�q��y�V�Jznic����*���z����j&������թq�N��(��`2T�m��fP���s_�]��cѫ��n��:��D��{���}'���q������L�,�Hb�W�,[t��G?KX��"����Ae�Km&s�i�6�U�/����a7��D���O�(p����#�Ns�Z9Jt�[�|ke,!K�򈃱1Q�sO�SЏ��I��j؞X�p{�`�0٦��%&�}n��"����ie��L�|MՉ�j���yVPO?�U�NtB����G%�̉�$u��QR��<��1����gly��m&�V��?K�Yw׹�TDok`Goi��
���/E��1Qg�����ث��C�f���������DCS��R��]�s�+i��BIE�}�@/gǗV�'l]�݈�!��E�i�Tu�j���Ň1����Vt]�&|o���Mj�Ռ
�_7~�<��E(1h�˛r�W�u�֫p���T.��$����i�*q�R�`?�zr���h���<��!E���fϗ� [Ʈ��1�u��켽�d�J?8D{y���� �l�d����ZV�f�Ȁ�WUl��	Ih~�L������qV5Ig�qn՘S�Q����9�1Vs�3$�@�4ь*^#j��B����!�����]}�
�c6��TJȊX�!'2p����(�@N/Dy���:������s�;�{M�@�C��{�.^"�~­I �h8p�{{�42_n�*�����p�o(�������h�,QT?RﷹL�.TS���N�u�m�U޴q�fx�l��u�|�ـv�j���玦ɮv�"/G��֠7�����V�	W��v>����!j��V'�Ɖ��5��a�������V�횃=-TT��B{p57���Ջ��I��d҄H�̋��Eу�6s,��6~�Q�����vy-�\w�����tI�SL�86b{"�&�����-��0�&$��9��Ѐ臺,1��-�9��ؘE�q�q��R�^���~r�H���Mn,��`��]�i9�h��q'��"��(��N��H�lsG�ױ+3�v�dn`��!�]�']�aG��]��t�ʤ8��N�rF�&�'ؕi^�����b�v�2�J�)Rlmv��'�@���Ud��+�D�A�ە/�/q˷A����x �$۶��m9�[��u�2/��&��MIKE ���f��>T�L&g.~�Ngu�]�Xp��6K�d_���b�N��B;:D~�8b�)�����z�+�d�]r=�S	]02��=X|��.���<a��`b��%��N��a�U:����=�3���������6���y�|5���������O��B��k��-=�nv$5�Q�R���<Ϯ��	�]xr�5����뚾*����sqh:����9����y5r�BJ/z�)e�̴����A'cW���,Z=�]W�Y-�2
н�`�V�ϻ(ӑy�'og!��f��W�pX�x�<���)��2�zn�9���wp�����q.y,��x�;���"��l���������*�Cu����;*��&��f�7Y3�`���c���>��9Sh��<��p%�Y�i�Z?@K��xlU4�=g<=m���ER�3ɡ�zo"=I������'@jRG�=.3�eD��M���nE32"1\�ވxEH�KԸ�r� V�|���u���r�>�K<�^���~���Ẫ< g~���LL��NM�&?n_�GV�qօ`�����):�w�*侽��%��npN4��v�#�(7�w���;���A����rW~۴�;�c�k��jZ宝Ii.�7�gB��n���O�v*Z|��L�^V�����y�u8{p������������g�A`>���RΫ�Hd�2�C�8
��a,�OIH�ŨbdB�o����6[��5伹�kMx��8�	yU)�4J$�������S ivEH�=)��;;���-��dh�O9��D�ٝ����r��\*ݽQ��u;)k<|�����GgSx)h��,������-O�;­VbycdƑ_�9��f��¸�n_����k2��a�u4E��ņD I��"o.�k�5�z�����)#<��̒�3��B9��x�m|�&��U�|ng��/��&�iY��|��.�wz##��X�v0Π��Hyq��}v�2z�,^fA_<���I`�1/b�:�%��T$�����P�3-Ϫ ��� K�� ����<3��a)攻�܃������!ޫ�ILS�@ǻ0�ԮP�<0@�t��]-� ��.-�F�]}�k��}W!3��Q�CX=��u���+Sf{�����w�h�}f��+05����<;dnO^��F`
��Q:�ǂ�~���������Uԃ6ES�d��6��,��4ًS"^�v��f�U��G�[�*�:��C�Ĉi�-�w?���`/����P��j�!mB������#Nj{�ǲ�N� swؒ<��>:%�� �z�v�YMPK���=�'�eA!��\�OV+�DH�O {^�.��|}F��-];��<ȋ�"�/����MLIu�h��y��~�5	�,���\%�h��P����S-B_FQ�sº� ��CiB�4}�_�3��,cbj�)����O�l��!Y:�LHƞ��y!��Ih�x��Nٿ�YW�z���1�� �adE�������wq�靐@d�m��Խ��9��0|"��;;���ė����nB{`@��E��r����b��?��W�3*9	\���9ŀ���w;��`�;wh�ӂA��6��$�`�\�Ǝ0�}�������zT���:z��h�/�/S���^������}Z�����&j�9A��wW罾�@��z��Ōq���Ykª��B��H�I9�7�9>����;�C��z���<�����4�|dHr.�۹��e�b�d�u�c�U]��1�H�mL�Q��e�P���T�T�
�K�]&�E��]��Z�s\;$��>�������S~&Ǔ	[�([J�Ca���'Y�&M��j��!����vd4(�����E��ǝB	ThZ󊯓�*V���I�ƕ���7��鬽��.ĥ<bU�tlң%��R$L����*��4��� D}�w�}C��گM: �'�(|=V�|���7���1�f�ks9 ���#�d�ep��7��`��Ajo���U�i�pLY�;D�e��P�Ű  sۤ�V�y?�?*R~Y�[x!�9O�32���Orq޳�;tSL}��|�
*"����-f{�W�ѣ��Ͷ�TS�!��vW,vB�*��/��L+�LMLab��l<̴�q(�Q]u6��\$2�O2�R�{.�g�9�4$�]d}����J}~����{�Ʒ�$�=0[^���������;FD�1�b��̝�4:>n�2������	d�aL���uu��c�S;m�ƚp�7��\Aq/a�u�_�DIc��X�/�S�3��&&�2r���~�9�)^Qg ��V
�rT8CF�xƹ��F��&�}�������ԍ�6,�Z����m&���*��a�\�\8��&OM��5l�?|T�m�X���V����`��v���Z�	-�(jf�!�Z�X�JX�#�Χ���ۂ]#�L�}U[�tO�F[����-�k�'!�R���p��uA�7�4�>!1�q�5�b��,�*�:���έ�@A4��Ғ)��G��Ͷ�B'% �Ϋ�_�Z�
��!���'[�u &΃
�0RM;���=eU&b>�u{sP�Y�Y����le�i�`��T�m�R�K#���ڻ�6}�T�
@�F�z�ɡ���jeH͵���'s�%P݃�*4>�� v�9��> +q&�1��Ѩ�[{V˓u�Z���o	�b�d\R4��ͯ�[W�A�epheD���^D�J�'��V�F��}a�I"���7C{�S�Ԁ���mF�+�t����AQ3<=�
��'�L�X7��!��r�V�&�CnW��e���?W�@lR?,E\T�>��b`SV��XP4���<2��56T����f~�5Mxy�H�}����ѻ7�S�G������d�/
��0�Ⴟg[�5�Ja�O�˹��9^�͒D��l���Т*0�p��%�
t�w�����/lP������8JE�N!�̇�ݨ3.���|ۡ��#p�(�vơ��f��,!����{�	��9W��<���r$���o /���,P��O�0�KL������e�ц0�3��)6o��`3�"�1Ř
i�� �f�Bg��nZ���@�$�¤U�9���L[R��5M�N��{�����8N
L�u�G�{�$�W��=N���-G,k�҅4�� J���P��������a���:)��pE�W!�'V.�ŞH&D�H�Y�����a�W�62!�F��/��#2'f�up�C	XS�'?����c����z�ު�v �.��>��Z��q/��w��i�5��3Ym3�*0I7ĢRf�N����N�b�O�f��`U�Tˑ�2���\�M�߹xُ�Ҵs�=br��I:6�����,�?{[���'ۨp�֫{�U���K���3�B�rP�
�`|e�QZ�Mir|wf"[��
�?J���*�A�@�\N�[ݕ��A$�����L�~d�u��79�Yұ ���o���vu%���b��6�����i"E�,W�:��z�m$$���)�����W�&��=���������ڰ!���7p�]j3�3pU��+��#�m�D��3�{�bkc@�wѺkq�5��N��1�&��/q�I+�o���̔@�ۡ������E�ޝT.5sjs�ڔ���9�����U�8�6��}*5�yx��/���>�Pp���5�C�\�rI*�Tv�������L�_� u=)ES�� ��Gvlp�hޥ�]1p�����a�C�5�(}���41<VL��먡�����4ԧ~'���f��F�j=Z�<c~��]L����}������쒗����,�$�@�T��@MFG���tWOM��εm���4�X\z��g�*�+�����t&j��8SMzU���8���T�Aw�G�v�����0#7Uc���r^�eo��t������8�cj���k��[�Ʒ�^`�j�.�/��.�LqY/�It��0���J�M{�龼��kN�I@뤢�\�<H��hh�5��`������k��a�x��(��v���k$!��(�O�g�f�Q�ki�p� =�߸}��F��x7z�DVa�|t0����}E'�4i�����U���>5��	�J�kة��Vs`] ���|`�3S����Y���"�����%�}���X�z�FH�	��W<���|��J���^��N������_x�H���Q��K\��}`b]N�E��pA��]&1�_ᵧ
��I���.vm5t�鱨�c���E�{wR2p��o�Wy�h���Y~H��2��Xm="�����R�<!�ܦ����������o���Ti���J���6�>F3��Ӎ?�9���3�-fX��[�*S W��س�<1�v���E/��3�=��S��s������ϐ�ԗa��3��	���S;���P�If���LyV� ��§�i8�d�ZL %�o����
�ߒn��L�M�"��'��g�DI�;I�\���T����{a;��]=Y���l�U^�&�M��Isq�S��5.\���׌��Y��9KB$�62m�M�;;DhX+�uy�Gٍ�U��X�M�q�~(����8"�zא��%*O%��ޢ�
s��~��B�2�� P��{���M˯:򅹞>��d����@�U'�����{��Uo=Qo<N�6�Sg�5t>d�A�d���$r7��>J*�q�2�#���͆�$��tq�-�}�-�Y���6�eg�l9�J�db�+�t�	�> ^�� �A���}�^!��G��.���z�/k�x��Y���� �-�Cӊ��ڛ�cԀ�v��y�-$a�YE)$ tU�W��F���U��d���S-�,:T�MVLԞع
���ż�a����&Y<X5=*&H�����/q�L�򱼦�gp�����@4�z�E�d�SnDh�n�`���H���"��b�VYF�?Rw ����1V��#
*m�ؓ�NT�	3�8yu!�e��4�&[�RF�P0���K�q��бZ�>ԑ{0T��k:����.��*ۮm0�Y��# |���t6�W�?)��.1T==�2S�hy�r�d�'���D�Ltߜ%Y�� �i�g���3Z��A0|�O]��m��?����1�3�d�*9ȶK!2w�� {�����j��oj�t^�k�%;�J^�P�t��)�<��&���A�{T�=��њ�n�/?Ai~ϭD#԰�vȋ�Lc%
����^L%\�/�ER<��ccE3W��� ��C�R�'8��@�^����J=��[m"J�f(g��>m�;&���R�̳ں鮾�"��'PA��t�&��^�����?OoO��ż�S(9�~QY�P9��H�;�2�<�}b�ж�#��<��AB:Twx
����k�`��m� $�5����#TgM��;!�N�6�ҡ4���i�C|�	<�Ӣ��L�T�^��|�H�LKn���Rݐ�V�|������b�e��ɀ�ya�!��MC���* +���� �~�z�iI�k�Đ��[�D��!(o%yX�O�Ɗ6�]��UV<�3pu�O^�0��rզZzS����=r:6���-]M��$�Ro�f5��P�^l���Ea)XMT��k�r3�Y��� gIwU���vK��d1y��b��'�ρ:X��͛�:�ܬE!���d�nu?5�������i#��/M�Ɵ3��#S��u�;�T�����d���������E�Srv;BP�=� ��e��5P5`Vy�Y(С��8[�k�G��t��j)����*�`JxI$�x�HL5�ЬnQ|�;/o�St���SC
�KJ�����s�q�P�Y��b��Q�ťU��~��A= �V@
V	�o���gޅ�:�f�N�� ��[;aU���e!Np�>~x��l�XnQ_�\���|���c	��^�z2���6�=����@�]�Ǜ��@]f�6
���v��� QO�&��S*��ᗷ�O�~ͣ�g��J��S�_D�og�<;R���b� �U�_�I�\<�`���Ix�Fms�?��R��ZJ�/�2)T�a�WfD�
��ߛ �6+n�>yN�ƞ��L=���v��3ZO�4���'�cHk4�l��YNd?_�ɰ�VO~:N��Az� u���ap���A�찳o�h��VoX0�c��E���{���Ά�4GX�����=���Pm���K{,�7��⦱_��������Iz>C�1,��q˳nE��,4ί�����r�C��[��y����vkKk	̞�+��s�.��'\d��a���
���"��`}z5���pcn
� �6�O��9�T+��:~�����i����w�ip����gOy��`hr�Z��Qjޓ5c�Ft�X-�#�v�9� ��A�#>���p��2Z��L�cTh�*v�MaZ����@��f��?�^�`�����ҹ��{��
�wC��}L���p�����S/�l�I��Pc=|b	dɠ	�����br���p9�g����ծyi�h�M��G� *�F�v�^�a�+$�}�؋(�F@9QV�������ә����_�U�
+T!:&bt6/*ʎ���]hv⁢�PFE8c����2hN/�2�v&����D�M;%`��j9w��fq���4���}F�o���֤jtA۟vW9�A��9�j0��g>�2إ��j���l�Pg�mP�Ի�G�����7�N��D��A��|3pda�'�A@sdwz�~��O����;-beh *�w�^�f��^���<��VD��7D���b�~u�R-(�{�c�vq[�y����F2-ZC��L�%������բ/J����9qV'q�S��ci�`Ia̪_�̮k!X&���Ii�+��;Ag�2~N_b����vU��|�v� 	���uV�2��	��� w@OW�D�"��,��ʫ�y.�|��P�=���Yn��W$7G�<��rB���H���3l~���Xv��*皊��l�R�l�2�Jb������q�v�<d�X�1�ٖ�h�~����Va���{�'Op1k.,�2�a�T�7�"�;�i��v+3�mƋ� "�>��E��U��`�e�͝�񳁡���<mv�b;zl��*'��-؛zm8�Yl���׳�#��g}Z���#���rV.����'�s ��h��G� ����g�X
ı!�e<ڙ��I��X:��{���fi&�m��Ѳl����D���@�����R}k�q�u	ȍ����;����^=ʪ
$�1��������H�ʟS1&����d������ib�� C�����p�c|%S'���7)������T��=31I�D7�S?D�,j`�Dx�~5�N�aC{Zm��|�b����9�h/	ŧ��I��	O� ��O%^���~��`�$�:Dk�M��;�E�C$T�K"H4�I��V��]0u�鰯��Ͷ[A]Š���S�+�_~C_O�%G��]Q�m��r�n	s!���ͯ�@�J�g.BvDh4�������RQ��aw����|������sg'���fȹ�:}t{�m�X0�xbN��щ�NZ� Z�J��9V`zJ�<>O�rFQP�&Bn>x@�>��֜v!t�����uZ�u������yU���	�́)�9��)Z$�r������$�=q�uKʦ�7��π�33,H3�X�c[O[�6���f�BZ�A��hC�W%�m?�t��}XPC����4�<E{�ˡ\%��$�2(��b{H��"��ߖ��F�2)�uqa���m���.K˻rSND�su�\�:�b2��^c�'3��x���`��?�Ii"o5��-9]X4��=E��w�5*In��b�N`�T!��;���m��O�
���K�}���wn�\��X�F��ה��ܡH 70u�Ko~�y4>��zo�󍠇_WaG*/z�Z��f����qTu��(��ԗЂ�ذ4�3ɯTk��`�[���Vdʲ��\[3���;[�}B
�8�q��&d��k���b�j�N�)ҽ)`�9c{��/>n)-�Ew`B���|2"���ւ���LքEN�w5�Q�^D���gcZxJ�d���أ�٪6@�g,k�qV5�_t.�G:OjI���yې���a#��j���[�4�!tm��,dnE&kp��[:��f�Z�"��@$J�Ĵ5�M"{��M�W��R��gXC��w�����^����Mr3e�'
:%U����4v������$��Eu|6�W�Yk�05�U����y�~�4z.��$�Y�u1�3�%:Ȗ:�/��+��M�kA���#l����Z��?
���Gh25�g�4�q�`�R ���t_PA�cU�L��%��ߌ��-�2���$G /L S��~��wnc<�As������C�['��	�;iD$7K�mPp��,�rעR�G[�'��ʑ2Eu�o�U�����P��]��/�l���U��)�+�}�jb"|�P嶍�Rw��w0�MG��"��%3c@����d[���~�v��o��4 .M��=��_��z��Eк%��g��s}�~�AE����q�XC,.�J�Li�g�y�*ͷ�'��j�U���O<P�{R��c/��Z�q���;�K84�{��@�q5q�ƭ�	ͳ*�G���ϑ�%�_��S��g�����[���b`��	�l'?�k��Gj>mj,3X���{t����u��8��7>V����<<N1��V�~=�[�����Â)Bţ~~hy��.���$��9�Xv���m��Նt��괞=E�"��]�l���}�j��N�6��T5�X1��`��F�#p"��/Y��/��ˍ�t	
���~K]O��#*��4��(�[�&�ַ^�������O���Ӊ2߁���F޵����rOp缣�''w����֍eFB2�L�rO+uJO��qP���?�9�S�.[RC9T*��/E�+8��i���ŉ��$E8jXR��W���+�<�3/ah{�������	lO��I�`�/yL�Ɠ��o1����g>}�/jjg��K$�o��-G��Z \޷\����ռ;E�r��կ+bP�*u��Q�AxfB�j&q�s�w؊�0	�+������s���9b#4�lho˜>k��m���S;\��#����T΅�'�����Q���Y�3�ͥ�Q�^���l�z;�[b��h��`jp7�Ku�VC�[�f4K7�v~���؊�(�T�����6�~()�<FT~Y<u�!��8�Z��e����G����q)с&��V��8Ū�W<	*�"�&�ʿ�[�Ȁ�����x�IpA��;{��0����6_
��\a�B�_���8E��j��z=Ȟ2�����!��VS��؊����qԩ�'��22�s��O�^���<�w������?-nxާS����9��� �Ll�R�2y�n������������V65��퓊s(V�Ui�7u��;��ƨ84&sR@�UBV�M�)��W���8���3����n���Se38�h�Tj�w���n�Q<��fZ�丸�W,=#���Td=�?cdA\�ɲs�5��7@�:��韲����"e��Smӡe�_Y�D�	H�4V�(�����VG��92�\*�1& �R�ra�/,�Wh��gY��b���Ʊ�򟞙4�B3g��F+����$�6-��,4ˣ����Ж[���򿡟�sn�$�Y���K>l�up�o��ǋ
�F;�6N͸U�<�C�qFX�n���-�ڜ�]]|1��(���8,I��l~Z[Z?� �Bm`z2�D�]��	�'��5��c��@��;����ֿ0
Oo刯��g��Z+$�ԕj��H�t�=�IU>��-�H�m�x��%w�jڐۍ0m|Λ/��y�b8w���Q �t?Dٟko~uE�4�-&F*6�m&�T���w%�r�Ǯ����}$uis7���'�n����ίq��#ݘz%���ԏvgr���H�
��J�ݏ>G4g�s����,����9u�X�L�H�S������T����N�.l1���.'3W�>'';ެ�o�F�;8�4#�k���[�F�/����a�e�����0s*@�� �6Y�W&GL���[PZ�ox1`U#�M|\�g�_�Q�d�6��4b���.љ�EO�e4�G�[�6�2��h<M�<7���v��w�#���I�e���񘟽φ.(�Ԉ��FX��$�=S\�x{�)J�BZ��}�?eS�+��F�k�5i��nӌ�_��5WKR���6�vSs5�2c�*�ؘGJq��i�vwS�����{\:L�ެi�<3�Yu(���9�ƛ� TH�Rtt	�Z�4�,5��L��J��:Y��r]�P�c��^LВ�.J��ξ�3���q��w�+4�/�#�)�%�j9�)�/J|����}M��������V��"e��U�=��P�p�Pա��t��,g��\t�	
ȟ���s*$�>��ؾ&�ep"�ې�ψ��#�Oݶ����+�<�4ҭkU���v0������)=! �����N@�J\�YI�>��<\hN�=�
�-���g�b�@d���}yƼ]�f��g�e'0�~)��v;�q����&f���H>�5<�f���_zV�w��SX��Y����"TH�Y�je��1Zei�y���憁P���bU�������Dz�-(4��	V�Ԁ�=�"���9��������́V����3�	F����Np���A�:�|�>��v]c�E��`����ޫU�Mtz����)zt�����(N���I=� ^����*:D�J���"<i�2���	[L���I9��<�:6�j�;�ܨȑ��>����&���xV�E��_a����N�<Y��إm�����,�{U������c٤C��.l���_[<��<�x֍��D��)�.��nv&uu�?�gsH���Ѡ�,���^��,�P���5���f������8쓈�a�� T����E3�/�ѱ1��C�c�ٟׯ����hD��@B)d��pB��)�����b�(WQ-�Sb������,U:m��!<�6ʀ�3*�Ôx닲	c�㍦�{�����b�*��Ï�8�����Svj[O�5b�4T�O��V�^1����.A���<�����K�{#���}țk%�7�˧	��K�f70�{f�?-����U�k��	�&��x�Ega*�R/���9,f�F���f%_�@Y�����`�Ni`Ui�ktZ#���S�é��ן;y{>/T?>�FPw��BXfI�?p���R�+�0{,�P1�C�Ff$j�Y��	&B��v����̲�[+�(�y�"�0�[�y�h3jP.�ʖ�&�^�6�U)z�fߺ#]]+Y�J�6���$���}s�W̕X���;���p&�V�����~H��E0V�ɔ[�~���"ޕ��%Hg��4�g�V�c6�!K�R.'P��~��E����
�	v�<��5�!�GlD��`f/;�6(S |�8��r����g�/>�):Co֙y��V�Xj�;T�B~_�p.�WFCÏn�\mp�����P����}�,Lq���>��mX�"˝e~֢{�FtU����#M�W����o��Bw���!�����G���
�Ǆ�_��P��$�D�bA�H9,�,��@�o����ݞ��[Kٛ�D�l�Z�p�.�a�[��>���"^G�j�)~��YLH+/�5��V�m�U�Յ�P[bW���E��s	��R<��ߜ�;���u��x&Oy��������c�����@e٢�/S.��L�ýR�H�^M�N�+�+�"]c.͝�b��˫̡'��jj9s�T9B���p
!H�aiu�*s�8�j�i9�ٽf�=�d��2��qN���5�����D7�씦y�^�sa┟cV�L�.Q(m���/��Xع���f�X��D��u5"����Y��L�`��h3F�Pb�S�����&Mv��jf��i���6��K���6��T�)�E�;7n<{���P}��x�p��7#1z�I�SGa�YsO�Qayˑ�����X!3��~@%�X���� K� *�Z�kX�( ͦ|O�{�uV
�[@g���8]}_5L�"֌��q�٪j��R��O�utS�d3�d������%�"�N��(��{�Z!����ߒ�����:Z����l���d�ŗ���6�o/��C�B9��O��b�b�Mξ����p1{a�]{��Z"t��Ł��ͮ�`P ,YE�Gjz�=z�s ��~-ַg�}��	r1����A�K/O� �e��K�qy�\N��ɇw�eP�8��k:�~�4�r��ՂS%� L��®9JrU�~��i�p� ��>�� `�4dx"��DMs�I���Y��~�W���煕|��+	^�*!�h�#5���!$�20y�����&��z\ځ(�?90�x�_y��TeJ�����_��ȓ; W�g!�+���G�r�����HX�S������x��Xt�����!Q׽>IE�ʺ�d"���6�hrڠ�z��p�=U�'������Ņ��Zvy,)�Zt�y#E�2W�*���N�6Ao��Y%v
�[6�?BX
��P*�υ�f�B��L��Uu�:䫿%>h�ٲG\��F�����I�L|�e��\�]�t�[j����,����(��yx~G��~e��>��7s� ���5����w֐�ح��L��̲1����썃�2�h�R"W�u9��@h����I��fDzV�.�y%��.��QM{$�ޜ_�D1?�ߊ���h�.e�\�w����kƓ��(��w�}���_���qG�Qid��S [��(��ƪn���޳��z��吼s����̩�;ʒʺs������#5���C�$�'.��&�|x�8�Y�R���n8ɍr���4�<�2�ٓ��s@�5+�ݍB��0`V~�-8��T��Cy4d�-t
��_��ǸK��^�}'�LN	�*��R�߃73�5�)J�>�(q���힥�ET��^� ��F=��_���`���l�e��(��|s���Tw����U�|��@S��xX6����HU���m��_E�l<��S��,�?]�f�i%����D��!�ʈvG����V�Cv�h�{�A�Qg-[����c�W������8���нH�Ɛm`^	{($��J��Op�<��ǝ$�>P H�b�u���o��wBgb���Z��9�L�(J�5����z���W.B&n� ��1�.���n�8�!a���@DHM��`�iR���d:Va|�����}_���_�^�.�8z4�]��i�=h{_�Kl�%��)�IV^$/��4"�+��;�h:c��/,ת>�����;���Nvr�!�>z*y��?*���C��	��XR����ҭ7S��7�K/�cf�}��?�z�Ϯ��t�x��ċM�1V5n*mo<Qݮr�P�%�<o�<zV�#@���	����[��\�x�ѿ�@\��&~_�E�U�il�����?2�V���k�
�x����� 3���2�e|mt��1B^E{#�7����\9J�.ks�_N@֠T3�1����=DL5&i��\jNMZJU�����wr�9��ԫ�3�,�4�����Yɡ|�A���:���J�g�I�M'���`k:���w^
��m*��K�5�M�xm���q�HmꞄ����,�F^�O��$<j �shh�X�ҹ�cA�9�o+�b�BC�Uv���%�To�W��$�s)1+����=s��н��'�ɼ�-��G��c���q`*:/�>@)�
���:�g�����z�i�	��@Έ��)8Wn����#K5p��w�ʖ�<�Жi�dt��E��%, �x�2�5��&4��Z	s�4-�@������a��UL+�xzЮ���,�YZ�0j|u�eB�;�ۋ����#�7AQ	EX�D�k6jU7Ƶ��Kj�Y�۩�>*FaG�-9ʍ7����J��y�Z4���0�.�h�=o�����K,?�K�ȋ��}�'|J	�9���q0S�=��������_�� �}yO�����!Sظ��g���Q���D�*�6*�nY\YY$�C��us.�x�6W��aF�Jbo��Z�I[F+j�[տ)J2=vZa����my��숏t��7h_Y%C#�ܺ��W��16�+���p����I93�N�@�~�k����x�!�*@}^̌�cv>.���l�Z�5r3�S��q���������v.K)�z�C`{\�X>��_��E�� O�`}Ͷ��[&�A��AK='7^�	V[�"K,sU�;�.�3��a&b�j�h�����C
��Rʮ��NZL����&����g!�>: X3�T�i��\o3�G���7[��8pqn1���[�CP����~�4��p2�WZ�����FI�gމ
^P��O&۪���P��I��|d���S��>�Ox����H�H�h��D��������1̿z�բdu�Xi�k��t}ps��p,7�]?Y���y<�0�lN%Ås�������4|���@�Ai����v*R7 ;5) �T>�1&�Q��N��0祦���(2�d��s�k10���:�׍^��Ȧj6���=��v:!������k�\_ }���v���h�7E��9?��WK�1���O~d�#/��p�cw�y�e���h�O�Zp��:BB�GR����,ўJ�sp��R �(��[Ղ9�5z���4�X���<(W��H�b?�_�(wP��������#UJjk����[&$�zr�O��&��ڽ:���r"�Q�|���{x��q�V��܊���˗A�U�F�m�����Fbױf$>�t2�rY���yG��%�h�%bt�}-0��^K����Xm�8�����r���g��@�,�T�4��˱�):�R.��(��O�#k#��+���}@�:�N�ч̚UV����0[G�P�&3����.�������݆#�'�!��.h6�c�|ҥ����&o	z�g�zH��ן��9����E�W{�t����yW�mj>7��h�La���ֈ?8v�ůS�TM�k��2D���|�B6�1 �-%�|w�� ���W���X�T	d�|j����є�?�x|�a���h�N��w���F�腲l_6���?󶜂�CqSp����A̓��w� �KA�@U��P��=ܕ���0똯�#��뗍���^,���{�@$I_��?]j��?ξ5X��$ѿ,�P�d��ׄ�<���{�i��N�	��M�"0�R�it����*�z�A����tq?r$�.T
lS`7�i�����ݴy�>.��_��&��7������������r&�&)\�C�:�\�y�I�iI}b�T��Yw�j����*O��4�_,� ��H×|���)�sA7)<TO�g����x������ƌ���^���C��W���S��K��������ܼ��[Y���ec�����,������:irlp��u�O�G^q.?��v|�����H+G��cgf�;'��MF�T�h��w�cu���+�À�?�=;��Z�+f�O�!]�6'c2�e�����'..�}�x/M a5u���^.�.O�g��cX��g��"{�9l�I����k:��}�Y'I�ΪA��2w�MTPN�rp�i��]�ώ�.��'��?����b=C�,�N�����-j�Y� �o���"���r&�|�Y�0�َ�jϳ�&�Vh����Ѣ��v�:��<��G�躕������V����	߽�}�w>���b�~��]4:<�rdsm�>��1�ch��-A��G�>F��Ǽ���!`p0_��C��U��+ω�e��Q�T��)����������wc��A�ys�����[x�$Ҧ�ࡤ*��դ0�j�ͫH(���F��C2R�E�D��zT'��o�a�F�� ��$��<F�B=�w���cO]R�Z͞r��^���|k����>��ag�f�ѐ�9wCX������8��I�:^x2�5�X���깤D�󏔌�CKcS@�əM�{��FX��+�ૣ�����*���w��[�������q=	$O��Il��0꾀6e�d�鸝�� �Y�n��Q��HYa�|ٸj�������CQ����-��hi��,�b~�H�.%��xW��}[h+�9��/>�b�]��`��R'g�Tg����mH��e$��dծ�t�)��C
��MX�/����R���,�Z���F������P��6q�Ǌ��c-F� ��߸������pAȝ��h�e-~�*��W#<b�yT&%�{>+Ms�Mj?#�`t~e(u� �faA�����}��kR��R��1^�����5�sK|�ǭ�g)d)J����]!�%2N`���']%q�G�<N�~>��,6�ƲwJyr�P.���gi�7�����cwǤ��<(���h���j�$�K)]��m^ �	�i: !�k�qt��r�	�NU(��'�5	�i�?:����J&	53�F+Q�7�)��LK%���6�n�h�g�'����M�/(�[
	����L�!(�)~�t&"���ƽ��I��/�,E{7�\e����K��\��S�C,+Cs���iF�ʃ0����ɑu�R&e��˧_8"�[M�[������jf�hE4hJ�gV���m T�Gn1�iq�[�&
���,5��)xR��E�CM)��7g+P#Yq�x<�'�-n�w�3+��#e�hL*�G�)s���������2�ٌ�����Vc`�s��;�O���5��T�s	�ׯ��'�[��U-0��?ъk��b>d3G�w���x>8Z��(��&U
LdR��n4����	h�x,�e~1����mYyqOD1��e�q�Н\����2?t�pB��Cpڦ��x,��Z�'v��N��o5����:��H"m��f:�olb�q�HOxg����)|�*d<1&Q�����[��{2^*_:?�]������l �#l��8�J�)�����ٮ4mZw�W�7#�@�{�n���r�N�2{�l��qWO��*��O�I��;�_h[F<��߈���ĆI�+e%�� lY~�stO��&���R�Z���ӟ8��36(� �	v�C�1U&-262��qz�y����Y'Yۏ�p������G�9��D!.st� ��pg�l�'0��!����!���I�d��n�?���[�pų��[�\���e��v��3��`�t���P���\n�ݳg<�(�Uo�[��ŀ��.�-,lIR�_�6�Z/f�Op�<��5��m��O����sW���y�^$N$&!J�џ����h˽
�L��'��Coޕ|��2�V�)�[S��f��J��J���;���q+ %�0sb��G�F�K��.��e�^N e�2�G���C�6��}�5#�"&��}�xY�m� �ހ�6�ڵ��ƽ8��҆�JE>��'X9We�� �.@�}�e�~��R~Q5E;��܈>ZM�P&%ahg�#��������W�]�me_�ˁg��b�V:���L;jdy��m�Ux��Y�yYB���p%"�q�KҬg�� я>��Q��y�Be�C�|�Tu/����F��o��~��e���J�}��b]d�C;D�b�}��i�gI55����9)\��\��x�4)�Z���d���>�T8!v�VH�`@T]�}��� 39.��9.G�C�Co��[yXxn�Ұ���� W�Ȗl��_����ؖ��K����:]�!Z�J|F(��ѽ�~L�A��n؛�&u���	��!���帻X�Ѥ�����`�g���ۘF�*�[�F��t����k���pQ�r�?�M����^�� ��m]��E���w����s+-W��߱�U�y��b�k�����3E&tiYZz���咜@m�VV����k��ߡ;n��s�'M[1r�7|��W���#�f�\���V6@E�;��pʡ΅*��0��t��
$���Nqh�J�#oE����e�1�`N�e�9���+���,F	z��T���gSH/V�t����)V���՜!cr
�F����M%��i��L��`�^k��g1��L�= s�Vܝ���(8@ׯ�>�݀#$x,�����#8޳Ɔ�<�I�n�̗�;Ҽ2��U�u�7��X�Fte�_�%�~߷�,vn����'��)��VĘ�T�i5F"X g��GD���ћC�6k�Qd|��{ņD;u���Ř����Y
��ۮb�ɐ@?g�7�=7��2`��fi��3��_ g�-f�S��|�<�y3|��S��%�PCOi�G��#G��c��B��!�s�g�6*]��[�m�N낡��>�SѪ:maC!��#����;z�LJ8��@��5@�,8�u^���c+ޅ\Q��<�e�L��9ކ��#��~�����T��q$0b���XFT՗����,|�2_҈xn45�+��-O�����J��s`)b�&V�,�Jqg/W b�ޕ~��������ջ��ͩa�����vx%Ylb�xHڃ�����lf �cI���>��RwJ��U�9#����c�٫�������T3A���MH�M�p��#�� �KV��E_�#@p6�l�I�t���i?�c�1������qm4g�S������Ĝ��w:�h���4�����d6��?\�5��N���Z|$�U���n0�(�K" hX��[�u�`΅ҭ[FEMoj\���Ā[ֲ5������	~ $�L�X��.Sf�"���
� �8x?"M��Q]�=s��(ݠS.ÎQO�jkdg�,d��a���)/��F��BԹ�����J���|+�!���U&T���ޟ�4<p�A !Cb=�
T� �&��F@�##�:<���.�w����[?�߬�\X��>�EkNwF���r�f̔﹅�n���r>Э�վ8�����8DZb�������}j��x�B�.&:(�DN��ț���^�ہ���}��O@��e�}S� s�=�� n�A�G:L<����'&�ޚ:4��+-�_�_�?���P@[�w��s�����sI|��0С��˙�g0�S~�}��J�H��#��s�A ��0��1��e,/l��$L
��21�p��Ր��Ӥ��ɻÜ��"n�!�������f~���L��]!����,UB��W xV�Kg�<���92e�g�)(�6�ZO\=7r���f�Lk�{�[��]ռ���(����Í��pX�=y��-�@'#.W�wno��jɐP-8#�=l�ԫ/����=��H����|���5�5	۲=XRf
�OHϱ���J�w�&��}��sQ�O��_��*w�#�� ��{F�t�pŽF,"w@�x�~��mPƵW�K���/��UJ�{M�w�b��ڸ��ə"0DM�^Z0èX
��/�y���=�=��,�E�,3p5��9����6' ��)@8;�5b~貑t�ܕ���8&��0�x���̢���[��C΅i�4V�<�������v�7z�����e�ml�b�f��"������	A��Z�!�7b�bP��/��l%��|������gB@(��"�Y��p��dV��VS�����Z�lX���5�h*���صݻ�~X�[u-�]W��	` \1z<TH��5m� ZC���v���������3�:����j��gO[�p=�
W�za������]W����� b}�5� �E�ͦh�
3�o�q�tlҠ���!u;��Ȭ_륃A���D{�1�2��+ղ{�� ��6��&Cy�ԋ4�^�F� ���G�B�ͬ���gK�'�}���ճz�IĞ���Z���R�������@$B��2,�xF[	!���㵇��X�s�t��_聾&���,���@ɿ�v����÷��Ax�'ce��m�����0��݇*�*�a�f=&�҃N1�G����S{��o�T�B�x�_�k�}I�u8�Ќ2^�KM$d����`x�`�~�xZ���`F�;�� ���Ujle��8JCfv7�3��\8��'7�l����>�a�XYt��>H�[��i+��w4��yQ�(FIs�5�Y�79����!�لmMD0�WKG���4��]��#Bl&T����aV$EVsgȓ�啊�@u�΃ݶ�����#>�͆��N��i �tO�9b���4@^���
�i�>��d�[���?�6r�͕=�X�cqAN��NO�Fc�vY?M��� z�V0���Cq钙&�3��}Cӝn菋dP��+�1܍JZ#�C��L���0Ӳ�_�bg�,����0a0%y�CP$x"`
���G�߯�Ա����Bm$N��֖x�>V�xm�3�k5�-�UZN})�����~-���Yg��_ƣ�Ξ�<$��J����yOuo�����|�R��e��:�ɡ�F���%�䛖�v�%�}V��Y�IRg����O0p�+�Eb"��#V��9lt��iT~<��G�*Cݰ��\�E'��_զ�n��H��P��᢬��~%@H��Z#�͈����k���~�����G�	� ����:.��
}��Qn}���ڵé2�aw���G�����LY����ל �D�v�c �*{o��
5E��Ԕ�
n	A�ALv��෰���^δɯ��Qc^�]��v�����&{�9�:c��T+��b/��t�7�ߗ���{Pv��?(���@�[8��D��c�����a��b\��4��Ўd�P^u��:I��i����h�[k-$kV���w�\�5���VZpf;�cWXD8mQh���^�����kJ�)8̿!lA�����x�y���ު���}���-\(�x�o݂|���w��\�r����1$����?mf;�7�Q������� Ic��,3å,�O���ɶ~LX��C�e��65��_� >���Q��a0�Y�q��u�ڦ�^�_�2�o�@�u�ú8]bg�e~&M�����{��e���yӧy4~��=O��(2�2Gw� 7x�A^��7jU�q.�H���󊬢PL���Nt���/yL��\x넢��=�Q) �ؠ� �3��� �/t��T6�[�11����T"��NY�/�[%tT{��4�[�����Fr�'糳���ZrV��g�=v;9(/��U�>�i5�Ԓ��#[ћ��킳(�C�gy?��	���J�4��y��g�G��"�W��$�Ϟ��8`�11Uŉ��EV�<<�&��b��~B���askM)
�����Ry-�K��}��SckQ&���װ��
�ԯvEWr�=%k=8���Ϗ��#:�-F��CS�.'r��6)L�Y��3�������e��G}݊B����:�d�e̎Ku����&��ܺv�4���9����||w���G)KT�/*$ #Y�3���z�bnI����K����'5�8>�<+O��s� .��*h6��ѐ�5;P�m�q�5���a��&x��_�eў���H^���<��ؘ�O��#�T�~��E#a)=���m[{ϓSj��T��*h�`J�B�>��.������Gíw�P0m]���Y[Sv� )s$�3$3{V ���l�4v���ŕ_�1W�bS�p���GQ1�eU������rO5Qc)`�$��N�b #�b=��I̷��sV�@=��I� b!Ν�.]�F����c4�Lk�zl#�WMET-�r*ݝjO�3~�Ak�V!g�{Oɫ���p&���W��kve���.ܳ���@��%4>|:4�lY@#���z$���Ѿ]��7��s���$J9�H��(A
	� O���F���rV��e@y�P�A�*�K\�d��t2��HS\���!�3ۭǨ�K�:��H����`�Ѽ��dqg��Ir{��ipL�t�����$�� m�ҧu���y�h�Y���dd�)_���:̾�0�3R�Z�����-=\��iJ�^�J� yP<0��_��5l�}���t�
�dv�m�=|�$�;��*9��M�/�+�,�6��v����"�s�8
��P���ч���z�,7���}��e��dRHs*�1����~�y��^qt���+^[/�.�5h�s�~����a� ƞ��3�KFY5zu�a�B��$ќ!n�zh�Φ�5���Ç�QȐt=���R���T/�ߣ� ��~rc�p�U�Z�&^�U�������xx�_��'����?��]Lxr������5������QY=H@�d�v\
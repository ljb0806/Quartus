-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Gpm/v09PwJRtHXOX+DgjgcKYQJJfRYGyj7S2DCprI+3EYvwuUfCLLs+fU2RfZwmmPylv6cORCTEp
lWLK9Qryf+JXDG8xhS5vu6Dhx1UyWguLG4KJZdP+Ae8LF53f0oTM6ESr2CpRVGLgXE7U6hlpvY5W
RYC4iBvgOVptNQ+0ZOneibsRsTnbnt4sX9UqHI88C4Z/hJGj8cdFMgKnuTgxDBzJ4HSaxSbpazVS
6tX0/gpJJ7KwkI3g6CPyk5VQQtHCauq9zbPZcS4gH1Qx7PfAAbEkqKmF5SiH/lKHvILRArC72kc9
ZpHMYys/Bhg5xaHrZAq7PHiMSZjUHL/nmX2Ulw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
QQJshqpsKROZ0V9NTnbMcgaS8VPYm54/JwPbP5geI6pWVftQjDgOBBB1fZgSTii9UpJq+9lBl8g8
pYuffkLA5aRmyspUIcASYDNSJGWcK203d8VqTsNcxEkGp1JTsHiD3EnAhoQ7ekuNfabEU8MNCu/W
atlJujVFDVuwEM/CQ07EnkeUJm/JHQzfoAQtFRAxURJdueWGHhN8eTrOECMQ6UElCWE/1WBVCntv
h2Ta/G/xZQIErnejbGMx44C/Ursh6K2BnvHTZUCnWyGE445wZdEuoT5cPcE+wQGwFYl4yFBWjiSb
/CXoWbfAFP8FMgUlvcFl46frg5TKEYZyKw7fMBTuiZ1PIYk2fLWNUMkK92FoBD5NL4vjTrerc9/G
6aOsOwKKWgcYuLIGAtAVTX7nJJL9FzTE0/CwPfe8juxaM87EYHLoDBKz9adcHy8zVunWDX4KXBps
lZJrBKrVyh1aRbGRuoTkbqVLfHiO/B/GHvperKODZZS2lFBqEk4Jj+jCoYfOFbvJDnVWgJAvOUA3
SDcf6CxPYNYbOG+MasHfCU9JzNko89Em1+k80Jf1IQtFOR+av9UaVfkp3Fci7vpBxw2KIN6YELs7
V2DVI3yfntvbqKo7uLsdnKUTh6iDPruwMqnNvGAx/Rvp36HpoSVuJvc63+jo3fzyyPN7fGNBbRm0
wJEA2LUOoO+BiGWY46UhcM0Uz3BsCrjV9qjDWUAQXucy+J2WJ2HwrkmQ9ruE9rym41Ln1eeB9Iro
pxdcUb/RYERbYR4eWcsqhzB3gQh3IWL4e5fQ67zoaNjYIHvUIWLlEeNxVA0K6DK8I0XmeGX8DPar
KDAxf1ffqyszH5QGoTIBdCY3dZNffVmKYyksij3K58J1+C5E+OV4SSllTIAuMQgtrZXy+oS91xF+
zyPPcq2p/Mbgkd8MrQQTU9IPYzjAQEBYnz/q8cfUzs7hoa7VUEM1U6XYy7ZL0rc6fWrd56NxEvZk
TjLRzsN+GPF2/N6qJT99/M2uInhWObCmleVDSXAF8u0H4AI2LA6CXgr0791tVaX4cZnJzg3i81Z2
7vEa6TRLo5JrXouj0NnDZE/7NRzHKRK8mFOMqcOLrbezIEa/P9iSnPAnZegomrNZ9fTAxFpagSoU
S1EbgyZhTsMDVRbcx5VxRnhdw6Sjt+l++P1t0S/+4TXLJrXIj9tzjUiDp+TaZHW28qSDzXoB4wq9
dy6SShm/y1pjbw5VLrZXVPlm+y7s3pXAlCJ4sqXfmzG+TORG3q+NKYZy2JZsXPTIo+SdARDB4xKQ
VLop7pB7LBAFjKuHf1n4v3g09+b946p7gCkRuGgCYhoFltnFWuCNUumgEJmEJNcaAUahVOggJNbf
rLdOGYEsTfh8QHJKZllg/XbZ2s3wT4qB1gBZ8TmL0Mf02bGzVDbOnwADkwPVuH7nU8tCe+Py0VFe
uMAfdFPeQGaw6fh5j3ZKJeRYo5OhEeiEVvsaPtvIkVDfhaAeX3hvLOtyLJcqKph3KE/3H07G1ffP
nurviPXVj72SIx2FbJWoU/bKxHS1dvHOqzZ9KkIrAP+2lQO7TOvoX5wD3QEf7LRMos3WOapbwZ1R
fnZCBfD5s8QzB0cCp0I6wK/ZJyiK+QEHjD+qD4nD1s1XgxzgbMFRuA7tH0CTEFi1vioumNCi0r3t
uh5f1SROEc8oDmPVP/vZbjVF9UOaPWgMhMxvFBKWUzfZmDYtzgyeGFc+prbiRVb0mJgD40kdpu94
sI8LvNo5Lso7acV/3vP1frJU1kQG3D7HfbdjxEQsfpdgoK958VeKRmZ1JB6jfiJvzM1Kk1kmWFtD
tcm1eqrVQrkhBiaxDqh8tODnuYtdY+wTmCNGQqZVQHiyNybZNNQsCMA4GXWcL0L4nip1Rw4r4kW6
LQttxunBurrhyzmLufuQTRAbeLnb04Xl2bD8fFU6GTl9qaEtCQt6ZWJoeDde9S4DP9eQU6WoSpTH
fqQ4OikK8C5O045BnuFOoCHfw06pl/IPPr4Z+VDzNLVHAGBHDiieL6bUeT9rgS5St/lY+3Orxavt
p81y2D0/VjARY+qIfJZizKetI34ehhVu/QfGb+WBqnfSQpOGhHW0j5rv03WxpLQEAxoB7tvwBDjg
G3m6i+qVtU95SAoue4bbmoOh8Yo6KYK6GrRrfA6LWE6+xJkcquDPQLXibs0h/KBSnVkC59r8fkXN
5Fxa0XA2iQP+hg/l9VLw1b4w63PAUwzV5U1dBfX0QdctZ3yM4wu0S/MwRFklvW3lRMEBEYA5zLCE
QE0/lmk6LTSR7QNqvnG5W9+gXc2rVf/P46WwApq79V+2+0dqUSRV/lxzh6Q8pq5kKKzcXP+rCaPQ
X95CXBNZn3ywt5YWFceRtJMuF77DTprpDv1/ddNQK8JII5I83g0+U2RRu0BZMW3fyZ4Ohcd0BZqB
q5V244Uzp25Zg70LDFDEC6VE3hA7xfAT5zBNDOTNKnxI9EuJELl+TA8htZ4J1QBgCDdblogYQwdi
KwCNADuEKp4mk3G6VIlvpIGm3+fB1kZGH94D3j9O2XdzrZttLcyvUWXEbZFFozTIyOF9pVpSs8kv
G9FfogkxzuoG65Qnv7anE7IFVPqiymVFCzKqqUq32KbP4rH3j0QEa//264XEOAX7gHYJ6qZNkgDL
xAoi6/9ACZ7LUdQ0wzkoH10M0+GFdz0e5F0+TEtSs0ufHkaOgKgtho5Kg2lMbutNt4ufVkOJVGdn
XsrmaSn2o2eqFLcUvzZ7r9Je4s1/7rX4KgduDHmSkIugR38GtUHm4EGQyOXHuCmgmjHfwkVPlxkL
Cy2XxbriuTvAHPlKNZChAIsH/R71ZWOSH4IfeBbMMuR13hTkd9OmHt8pWB3Mj4zvizxssb5WgeGe
T9D6IiMWhN4tHEuWhPoyeLzGABBXZoY08P8l/qGrIij29VZc+LebBeu8PM/b27BrTrF3p7brG+F7
OOeP5UDMF66SyEvM0xhHr+HfZkUDoX2swf8lumUfT0Nv3REFWzCHdneObOQVVOB5eRfzwDUfBGpJ
J0zm2uUf4yfXR3JGHi84KaaCxJcahu2bc/WoabPzWirKIqhPm604bKpB/61GreOYop0DmPRUPUX9
t1EsiqrOuyZZoIYE80QSxLm3G3fWpk6huVUkJdpMYxzMQDVPYvtF5F1u0pu9WtO0vBgQTRGAC4II
CXieeaS9MSERJDv94kpyxn9ALaBYemz26eu1xqB02+g1qMzYlis3nqOvTSf5lZuHPT9mi46WhG3B
YnzdpVBXMZWtXYj1WBHffK7abji7ahM/0+QEID1mHheY/cxWsaZQo4q6CMEi9kRnQTQ4CkIqkeeK
0ARXicZ9u1iaGyr6MdKebmdzDqB0Gve/u1Bvlff8TdefwVO6VF1AjCjcy0Vhq4ed4U8d06wkAeoU
x4RNGrHeKX81Yqz98lbMOtCErOCYHePF3VrhBFu06SzH/eNm1YNDhJJLs7Tpas1SfUGwf6Rkhycp
ge3kUM/VX2/xC2S3JMvZKgrUXWR8ntejXO1nemgxVq0We0yhjFBHVI0greh0Db4gpI9JZ3xvPgTS
1Rf4y/+6SExjNs6Pc1q+jjh+9tgMYupDHyIoooUCG+Z7B9sxYJbBPKvOmSjDbGIqle7RokRv40ij
hX7bMn2hN7mNQUlO7nL7pMAjr+jlRs0IWdy8rRahRNrpv2AQl6FaDWy3ZTsma/04m/dPIROwhXKP
HwZUR3KR7tRdC1RKut4RlwFmDo/n73Ai+ffKajzCoL304GRvJLu/KwA9D3nhxzpcMLVVMXSsxo7h
91ERzyFMR/ia8/iFooxlPl6V9ivcY/z7Xe32qJn32NzzepZ8OkFB4WyrFQpZ/Ig6XPTawQCpY+Fh
ryqFoUiltUyoneLUpOD8QPSvsSLOCrL11wQkBcAE2ihi9T0febTV0iGCuKOx3h2nR1j1bi9zXsRk
mA2QuNwxhfJ3fQQ3h2O78NOI96wvKsFitRs3C2K9jgTHHkWoLpiFjkvmlNEXM+WEIRVtoMvYamur
9RaOIL8SoohWQdLZYC5963Vi8QhQOGFUMkRtHy5XYdJun5JtWdvzYn+XaStIHw19NsLmz7QOuS8V
DT2o4lc08ppNiX16dQDsjVKsrMSy7y8e8BwM3NVuHWcFRJcS3mBC5ob0iplPITYz8RQ49ZnHW298
shA7YHj3b2/ZaujMQ9sgSSOtmljT5SSPbWQfglohMFc7DrIpkmK7sw/ixSb3gpSR8Z9Jwg5Yo2C/
Y51k/92Ecx+CYbj7IMEumxwoteuPm0nifeo9TRvuQhctU7Gh1SST4Ge6/RiZB8J4JLirKCHMMQdT
eCMJgYv5SV5wIoxGuy1ld04tFWC0Cwrlb8SZabzAeZ3EOhswqJY+ZyfJNWPUizSuygroZ5DUtxlW
3HjCNfSI59v4VDy+8txNDY01GsRxM2CzRn0nJ7rOuTmtuol6gp12rCMZV1ylVbhOxFUTymjNug+d
Ty2AKN22K2TbIfyetW4Rbgv1bk2vEFLRnBnWqBy3xYOJEJy2uYkUTlHTd0azK4D4UcB2Nxc6EJFq
6A7JD9CRz/eTl3b2a158hRt4pQ3QnXNT5LgcsFRKfk5e8hSyNQHNNSlpdRLW1IF7CH3Tylt82llo
T8lV0LyBXMsZv6c+2ROs3G7u111ZRSgAbnuZ+KAnrTusa/vNxkWSP1/OuasRd8q7VzugNhM77orn
bmv0sABliiQDEuzsgGJ3oFeFIUQKrf3AVOpblc7zNEnPt819Rdav+SbPHWkj0yiCQl9j3Id1kdzi
lvEIQvbBIz6GYCkjt5rEIsbNJkePG773m+Lc5NqJWJrYI+XP6Krkgpm2EpcI6UhDAmqmgc2QhUJW
XJ+b/T8edJXhTKmIg9zu19j7MpvfV48NtKmGnGgjuteHJ2Ij6iwXnqOhmzNJa8pW5CbykI3Pi6pM
PaVnQ2wDtcnhsREvDygLWOc01JYBogkRu/TldGS2dwzOLVrG0Uqd/4aesNExDEsfSaKfaC4xcsfX
ZKxDm0ltEwlwVi7GMGvLiy7sII6CUF6paPzmqMybvyzCyJ/oFE7f9tAjai9js9FocYbmDkmKNjEv
QD/EWUkikSpiuaymxAxUMkEDrfZ6/NRVaKOcCsWxfm3+N8e2Ii7RBJkP9u3fxOabr639Yx2n7+Ie
cnkQrrk08qIK41EGDe4EnSGET+ESbmXD9zpbYiC76xmUwJe/PjZ72vNOb59WwyyoLolbPvSUhTaW
iD3lPlxLQs7Lb5AmF4hsJJLT/nDttL6qLxjfv4zlJgJyzkU95ZRn42XL95PytgXyoz5jEUg9J4ej
xSeoqMAL2LVN0QO4qA9P7a/EYhtUxVnAR/PpjtqhXhGjc3JUqU4+s0vDOIBux0vABE/BoddDWfIc
7W8XrK+E1kbZd7ulaH/1DF5i0KbBXxVNaXmuqn6srTKehfp9DlLQS10eqtziCohKJPbwZ12RXZGO
cWICom19wiB24/AFIn84pFMFHXJRaI6vxBRa/uZaYx1tVJ7CSvXuhXAbXYtahECP7zOlo1m7zfRY
4s0Wuw76SZgrKDqSKjODGlytogjKxBUCXbNVgKIJEDgVop7PThVFKyfqEo+fBh+JZNuA8OcZcpkv
pVNb4haaLO2lDSFmay50t14TTzJQwKfqdlxWImJCeUL2KbbV3sYnM0BqZs3W8+jYOZWjnFSxj3rU
tqES85rqRdsfmqUT1hEGkC/E1Q9fHFMUCEOltOXSSDMSwvZXBsIlyAuYuPVCdWfiK3Tnj/rJS3rK
cACYrGgMGvnTBdkyeVP9sbrdh2ljoivx3MdhgqySE/U2nNhp+/udFBijPFLCnu8jy45PzXTwg/GA
QNOiTBNeucicZVj9seVRsM9+YsUrmeVEbeeTXVV84ptfXilOoQTln9f6WXLX8hUQJBNxKy/zalWD
qDg3AAC7T719Xr++xWsjRGTg0St4+1smVHM9Y0sFRujIid5oNv0FQItnsva+vvJKE+BfZCiIOxJf
ZFIy2NxiatKG2mYzVDjBMKYW7x3ZkpO62iIzE3iaquCZuLn/HK0gPjK/zs1s0NvMJN14Qtrl+hgt
drQSjinlYypS50tq2nWxaOZ8VCZNZJQDTmHMOEl+CVcsLO08VUKHrQ5OTdGduVt8UF4ZZffjJbLe
gf8CX6X4ah6o2s/EwVGKFV+RlYTqoPP3B50D/ECNZfD+tzezaEAvc8N6L+Wl1AFP4u7LENE06g==
`protect end_protected

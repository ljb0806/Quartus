-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
G0gIPjTfek0C+jMLe2wuuJ7ijEBBgbHMabh3QanLdYkwIiokG9Bqs5hudp5g6PdbAHXJ5vPXcl4l
2D4eyEjkz4Te0Sxha4urjtV8Kblf3uH2P6gbkJYPKal11jaNTJrlSgq7U7XG7nlJxvVzv4EyIuVA
HHO1zcEQL2nFZ0MnLg7WH4ScHumrqD215Mlqm/VC2aKjbrv5CL0FAqNQRfg9BFOt0qyujgOQpFVJ
tQlfsRto4XJHqbpMqIhGk9IwkBvuSNNvC7ELl/Bdo2ZmlXCZZnCdlp425iawPIH+zlpSJVcw7fkn
Z7pU60TrvNL44EqAVFHrMMSjjHa45UX51TArkQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 50592)
`protect data_block
cP0IpzgzGzwP42rQHQWE8YLZE8wwUom97qXttRxkqYZnhIfJKWV8woLyUtVlCyvhCL4DNe1WcDKx
ChR1FlCJVUjPq3ZxIiPx709o9avLW5Z8p2OdC3gkm7ERzb0M/HQJoVLGDTo23b4rm3GRLooEsvXX
LBQVBDSqUFhuYV/JHNpy9yccDqVm89iiboEqmiQy3qWK8l9ozXb/FXqQ+/NOiDHbItDbSlNxhrxP
HWO5NA0fFCnGtw0VMcqTKNC7TU1BnvUe75dM5I43mb464QCq6XJFFDIdzI8e0vYIxWen6Rh4qOfd
xCEel/tBoaP0lCT4dovJ3yuVpfh9Jn0ttcEnQ8tIfXsktYiMQO3EvF1g+T0p7rc5Ryoe6M/0DtSw
si+jp5vGpY7e8vORjo5HJblNPogCudOSpHmty4yPuFSrSaIOsctF6NK6c9aHLYxb6ut+c1Ed5VqT
ycNww17RU3jhFIqDpzjq4xVahYV2w2bfEmS4zkiuI3K+9zoX3onekYjTyFZwLH5t/oeYGOxKjKTS
DOtiydWjympyP4dt9+tZEXIGiem2xK60DqcnkCz+wNvZzRJ+zIllpdMwzrsiVljOO1jeM+6QIHvK
slo9pAcvMxbLwlaDfRmKEjlU5eutEi3McvOebsFTrmDbVTSCgbGI+I/ZjEnYaaL+IJVz3fHEvmtY
MOKSC7UUsIkR+jhtqLPod8UWn4k8r7ZfgnLlXylm0t5/At4vbgO0aE13iM625JHdWAuO5GsfJwiV
VKFDYa76g8iMRx9Av27bhbuP400HsBO3utIcPkHgtrnVoJJQ7hLSZ7AK537VPhO8cCh2BQrJGXiY
aV/ZYvp/FNv+zEqxkud+JwaEE3HB06YuC3Q90DNW6GFsEL4FWw4qhGMSCPDAoBl+JC3zfxXie1D9
KX0banZJDmlim102dv/nmHoKJMZZEyGXSALcmelunrriy67G2Un9x/5qDez0cnasQAbO/NDMTqwp
zO5uWFPWe5uQf5LDPj6EzVUVAh9yPemv9eb2e4E60nX3QwNan35vI6+7bKjh/Tu5TyK48MYBvavs
wVKy/1rkGSMXG3o046MyC0t0jeNYKPcw/2O9/1ZSW8/U+iZk9yKZUPc5EAebNFpOGORYjje02Itx
FeD3lvP+jn/ZSVq2zG/xaqTgQQyMFb6KQSvthcrY6S+cWeEfHwXjyFyH5kDWXhiIkpajAdKmkbs5
HV1ef9QfznjiKafM3QzMhNfzzfw+6ML08QsAfjhN3dyOuPV+FCV4bEtXGGczBEsyoYVdlJki9Xnh
BLZ6MrNBEeSiJvAkWKCLEzTmnL+BJVAhHuYx5QfMZYxXjLW8tCNV0eSMw5hRTIMv32maL6WSHmVU
sm+1BDaWH27lirGR9vgBzEI3ksUQ1TwrhZgxzLTSHN6JIEwqnrObS41IQdOhojfwX3lvwaHhasPT
epB8z3PoPyPdY8/4MR2T4Fv87lGh8J4yoIlzwo11dki9pCi4NtQogoBDhS6Rbr8/9e3LByGrBhNP
xLN/pC8AC8LXzn9yTu9AHb7X7YdF+fx3ESgu/L7pu3dkE5KCYmL33/RLs5ee36HPQvetXqVpHYFQ
tAWIa0mGz158FS8yjBXPH+P9ysDkoDJwxDrGyJ+dzl4xlAcl81NSqy7JY9rIBoyu/ckoCgaplcq1
FD5v895PSeZD/X5iuvK68mqLgtNSylzwuX0vuduQGLtLD5T4L9MnhIblZz1h3j04DtsZjb776lqi
/Q7MqkQ21Bluhmj4rx1miHDJiEMiLvPu288ttOJxOKVRnCtNvWA7ySPEGUqul8dd57Ockf8wImMM
/suMkn9PnJObVlcI+4WCN/+9PoLmZrXsiOFNUhU0lvtFDS3WK7cIPD8Ru4tuzcRR2XqHXC8pyAle
j9KOjt2vEibp0PF+lwin++bI6Q9bEMVwpPfkpNtBwJQWJefTNJkz1QKsQydgC/kirANeJd9OLrBg
6JHkyVD/tZdT/U9txLKUCXHMfghk/9LMYdJJOLY3StzlQywCJvT0rV6g0xA/1zw+dwCHmqLqZZdn
QGWuFSoOiSergLBsnMNUaExNr/KpwnWuwPvUPojKhmjGHtt3qnQsFs5YP/U60zxwnQKuc6eyZrQ5
2By/auJufm16/itY5DCzNeYhYBFGXe26fePsyXH/S/ZonY8hLwblqy5RaXP1e3gMQPL79NOjn5kh
i1kqlDXu+IDdXqgpvpH8Zj1OZejidEPGrud+ll/bXHwLHds5zT34zJXirw5K4CyJfpAmk7aMqG4A
aENaGJI+dpYpWCfTC96RPbHm6o/HGeuXdEsq94DQESuF1+PAv2KveEGuRTq/OHNqoY5lvJAW0KLi
6PVsvmQ0qFgxTueL3zN33BaiTGzYemb/Ev1wBJZy9lkf4WMlQNZMSYUOqsIgBBkZ/cltXvDAIIn6
zhJ9PvvYWMNiHwAgX5WxMAG/K5nnJPtCqKStMvE/bAi1czJ2JlY4oiDuSJqLXDEiTxnPQzYODjKd
JA1m37EZAYGRW1CCBu8nVOyID8Z2Tqw6yx4NsyBh+eHk5HbL5R30H5OqT68pxpwmeBMbKjZUgjG/
jCpJLsAnjDm0cLqnzKLmCV8AldZIoeFGTwp62ygc8BWjF90/NxWSiuNRyDgjFK93np6wXGZ0jpGC
ub8Iq1mZ3b0O4JGAZUEhOsUChGlCESJ0dzVyzOMseONJngcJ364GRqOdcBtlPuhQhuI5rRm1bbG+
sylbZOZO295zBF2IY4zL3YuymFnUzXQ0D5Vzmadf2ou/r6ry42hFOCs//9UNBH9004Wa1pOYsmVl
bQOjV20ZP/v7YaV2tmIt3v4PrmF8jo8aaBhYRoiNnINtNs73TjvdV1cfGD9b7nWv36sY77OHe59K
U28R7E9wVieWHlseOeSlOJ9DmuUEw/sJGUhZ2YAu7EfHoXhTmXMCf0MrkMNp0XFcavjN4MtpGkiT
VorzaRp3VXpxPtrfVxA/hUZspNr0U/QNbsHq7hKmSRvfzHpXNd9sFYuaMPDsolDQ5MszD25nkzKh
pcHFGM2aQrsW7hPGb2Zxnv1weWxl/X5YLNoRbKBwpidN/TncKX3cixsFZVesF7JQgctO22TNijSk
oIObNDRIx1YJfEz5AJt5CW2lw/HK9ao3akLYxobUpSItCAtCD/kHf8lRrKqL9ZEZ1OK3j9LgZSlP
3ancsGDVYUCuMZR5YsinUss4P3mrkqqHrWYXBJbRJWQbG0D/UbPeoFi9uuV0mDf9jW1Ig/wodo3A
YAadjpwQY+1QDRat/nnzZ/9L2aYOQmpJ5RiTHjbhy+rRkmgAZ/SGHOm9RuHzOISX0IAw9c8il643
riyD5MhdVoOwmPCd5MuvUPNkOds82/EYnUmqhySDlz3XViaaUDiu1gH/mzNg9DxL/q3sppKpZaHR
8kIR8BHtO65KqXZ1mL+wccQmdp0H6WlNaKetILhxzAyKeU+hmFh6wcuP9LEvwcQqtwOgoXM9BmAe
m18QKOKi8gDlDgQFFk8VEM1OvNoK64N6McypHhztTjZuRLfAy0m0YAPiq2kMGs42N8kYLeCFrhRP
pcifPSsJ7VXYShihB1R7fqYrysNXceFiiL9hYMXIMEYgxrkgsKv/3MysY4iSCks9Hb/dLEj1QMTH
Sxuo9lYfItb1o31Bj0uUWM0zdoV4u7i+TnwcoNSBDpP5MCQjasxxx4JWtBVLkG17Lbwys87I9RKf
rYkJQQ0qo97LjCfUxf+cYPbMs+X8pI4O+CvvKmUW5wIU3sTlXF/S4RjpMFvvBEPI67sU3XoVEnBu
8nxRCz5yGqAdegRKx4vO3DA+8oMykdqG8JbE/+9XGh6/39CdBasJB+C0iC4XP0cFa+GgpCKpKDMg
HTejB/7lGtmOP8y/6pKBa6rwoT0Ap+ihi/CJ8/rIbGyvTcHuIiTtEEq3F9sI8hQ3Rl0h9AjmwjNN
v/a/KK8JrBOesaec3byI9XM1Z8typszmboD2FwYAPUsREBq041SN9ddJ4QeMsjcoI9CAbZGXaPSy
J6ALNDRFgu+DVE512N0pDt6dL/EDgtvbjePpp6QatrLJ4E10/OStkLlJAl6JW451tcYMWQEPaAg+
/PPWS9NeoMuRIr77SZbCL36rKV9PtuNW2rZul5M4EwD4SrXYFBYaHqAueu/ApNze2m0v93LhYLq2
GQQ960rLcP/XB81Lg2ifQkn5iNF+oIOguiQYR0hscFEsgR+Oe1ZU/YMM5JYWhh2pZphqbDPnkc1D
znDoA9EY6RbpR3WH3JbKDe8439F0jmKFoEvRXiOI6ow8zgSdoOyZzoL6L8POS8D0zFEPldBFo0m6
b6QCYuZ5ZtA0yjIOLUu9gyGftzfUf5oI+6aVPiuWroWq9O9Ew1aE0DZbuxTt+nylORT+z80RiOKt
I8rs6+9cfHeJhWVvQsQlhcHY2bDYEMrBB3FRKS/GGXfyYONCY9wTFDALbEH98sX9/MGJ0yK5UihU
V63Wld8sZE22fSNustX5xX+s0uXRLFFMR6XriMZ+NLIvxRlP/1JArvpYctjr/YAn9BA7ipdEXyxU
4kXX2r3P9mYxisvlxjFmNSN6KkCJBlKXwnSut62O9XlmhJ4Kzk2tBlvCt19J4rQT2I4rGwkBg8cx
vT1KifA21/dY/C01PBQ/y19ugidt/TUpi64QTdYFsd+KSxAJJVGjbige6FFObwYL+5KYUDt/gUmZ
ClbCUBqXMCntSIXilVzRvn0IgPp/bf/MMUa/DKZFPKAmi95M7eKVGxcgAUrIG3YysnQ7Rv7PKfox
/XzF1C2AaxAM4kcql8G7mQANVjyNXRxdSDvauyyuZu9NvUnrlA3L+PdCR3cTwsNf1l0VO/6JZWLY
wLWYkOXkOevU48CgAMhMrVn66F61/G7VVs579MHnWPMXGZTuLkin8k9KAF/d3n5ySdIRSREDL/uf
fYKuGXVd3AaiiWTZ6rOr5fbmjh6EkDIwA5eis3ezYI3ajztqPosWYpOvB6WwfCZUrHuevGHrvL6v
IMFgWwSvrYSTNxDRB69e+RSZLBWXz1/MIJSiz9EuiWaTGJ8Cbmm/pq3hfhKVpnB7wrQJ9/8wtVX0
y7georQvBmRoOXO/A7XBh2p7/5C5ZgxqSltJcRDy7+1JIKYI7NCovpgQlcZL6v+4i+MxdQatfOj/
mGkBgiwo36QKy0ARtLUIpyo6luIw0WAb3rsTHFLjg9aGgyCunBVfesDjhac3VdnOCyQqgfKBh63h
+puadtzVjmMCsHCrWH/3qA/ACVFUbVUdqtlLT7Rdr9IAeFsrn6d30oDFDZBEt/aZUJsWcNL4KbYm
sPTQtcTMrWGvok/yCODqknZCm/ZLgtmWi9mYU0o1avKDHWX1FmHXzvnKcsAki/iQu++TW81AQNjq
87aUeJhnCqvqM6dP8SnD1usZr2uCw3nghueVxSzSi2/vwi8Jo+YIEgnhy+RVFJ5QgrDc91G+lb8t
xcfI7s6aXUheiyjiDN2XKkliSZBwcnRUBL69/pH3XQZR6+cPQiInCaF+gJUsyJ7A9cDK5uyyAZt7
O1qal7CwPAAdN6wAqBzKODmutYFvlsDPyLKSE2jMrfQ77L9DSuSdIuFPsB2njmG+25H/hU/rI5bR
XEtF30GwHjP9UgsUGB5CNesUPOpVS0vgP8q1ugRvg5YHnXdIO+ef+DXUjO9EEO1/Ji5wJTH2hp8C
wlV1M7LmYHdKhEVQQSdoCJTsCSxHPjhkgIMAy0ulHnIxLwqowsp2T7TFBIlSma70IFKP7THTUtPj
ePxCe0nVnmxITYMlR2FIUxcGhZTp6xKUATcuqmhC0ekOfedxe98JRLggNhjyoqOcWKMg+Re9WE7Z
G26otsiOF6rTW5VchBSPmmOW+4pcTCpZ1PHXvRWlC0FSAKUfXyp8n9O6xWZhlYaqtDLiTTj/ZzGI
s0b4biS8LfCxpETl1aaJkzLKbuZsPvtvpGQzlfD+a4HsFuAZKXY1N3P16M1YRakpZ8cwph3uCv0V
t6F+gqZabuFSyIj5QqqS/TfBVcMaGPJP7Gw5m9wb4c7GfL8PhJcUxuK5N1nrYGZK2KWkF2JayVWw
06Biy0jHBW9kQg2wXj4NTpLjp7pvWVuyE5VwS7E2lGZvOJSJT11OpXUKKGuSpFWlfKCyHycTzVLZ
KjPWOVt0z7dgQXtRs7me3oBdhXuJp8YGDvlqesqE+NQ5Pkpg6+R1QzN1V6CNWBbMP/0OSSNrE8w7
vgbWnUuihXRM8xpHAW8VZlBh1AdtBn0zLH7jmehHgvtibi5d00euDHpD/5pNzUb8QzDe8hlBYJXC
aDX3afvymx0d+d67kRXIRqxcfefikUKlRMLEdIInw3HctMK0eKLccgXPoRA4lVzJcGVHwvPZHjHH
ZAhY5rYNZLKp0/9fTia6Hx3zbUL+2zJA9UpXS338QjZxhlX/vTRwZvv60lPHf3uVwoH9nmxXYp39
/jaOGvQxNp8ZN4EyS7OzJr0wDNbHQwTmChyIIEBaFsBGiaSJ9aq0hPUAEmYpLLmndA62vnM78I3/
OOapv8pagc1bqClmlg1f7u6cc9LfG3nOgD/I8+ZYrTmbzd/INoIcoGm85R+hSQ61X7AGY7U9mzI9
HeJawXJe9iVGcGYIPulscT7tpYUA9lV8tXw9j7HGjksXTte1mjv3/WCyprKMKb+fk4H9GKWORPIw
yAadyZM6csuhN58Hm2seBaFFxxTbJpnlB80VvTxNbH1+ikkmtlfa8pPwxITc0ckjO83bVGLNmmg+
iVFOIa0HzLT3HDDM46Bj0+VXf9AvGjVUA8XuUBLksI1rZf2wcp84gREvmBRouXGle8SVdNMGJNj7
+tU/YA3geCBQYQByh+zXf0OHek3s2qVM4yEHUm2K+V+Tqu3tgdPnHMmhk3HMG6yRT9Anq39BBRC5
+p2j/MO1Uw3HPNgqXvk5QEaj4F+xaTAo2MR4hPqJzvvISSjjz+v2NtXrniTLtysVyakretNx4OYq
sCLQo4jldEVbwjql6DvOzBMdao63dBJxsYel2izLyt7T8rCmQTQ3/SIhdR10xfQMFCsRzluG5VCY
QpTTqUfYARqGOHb5nTIoI6M3qUsEKKWG6y3wTIdAVkgLrzaIofp1Za7NeeplP5X16H5F5C1QhoEK
4o/ZzY0pZ2j6PqMPBrGWjT49+e4oJ1oFwM8j0JO9o+RlCgwP1g2rvX1aZTMDWPNyT/DpStwcbxmj
oXontOPC3qhmAkrnRZ2EqPWrTl8JyLukyadWgqdVDJdN+XaZuIrwTbVok/Wr0+GBs1h096JVCIW8
Jc/2JxiyGuYw5TOFW+37Xi5L2GaFEz8vZ+viDbzJhTpUu4f0UFozRA2PEx43IzHRsZrYXhizjPpA
5+NEXNv2LeHr9AeDQzxHYnn1wOm/rp9H6KO+h+RPmSIS6AxHRIvgPLQhwveZwUljY02AFCZ6m/wk
+G6uGvmCzKi6Gg2lhKyFZGLGJHlHCvtopzJMS8tqvTZpJqLfVuZBsIfTLf3HOUO0oGYySUl14MMn
B6mIRwpDLW4ZwtFJqDIxI4PpbRrWc1IV1S6b5eqOg0lxCiChvItZvnobiPldSXe3jK0JSa+myQY9
A81WAX/JaTaZRycmVLijMEVFl7A7Coi1igbVQ1jqOLb/nLctPjym4eZcfUoAvJXB75CxL2QIe0ZA
y1JdPfJIHeXCJSqi0KwwYbhIJzFEQ7alYvAfuUTYQVyEpU0tvLr0G0CFiWZA2RaemjwOgRrjQSN4
WOviMv1l6WK9k6vTSx7sA2JjtlGRi3OisBLCw/5O2/zhQFuhOfumDDd4Hl66GYEtgpHOileiGEvl
MKXVBrtTlRTxxWzdD+dCX3cbK+Y5plabcXB4YURgBaG0INmvtlFg907p3sYjc7oDtCaXqemQ2e+0
GufX7/t+5z/CL9+6gtUEDO0qF62Y6Pv1w3KBuxhbvKXtLzzzh3EZgu0FHfbEa9x+BGm0WQCGVy0W
neAsjx75xsn+P2lOWVLSoRCXubRgLea/8F/a1IC3gShNF81YPPPD2P4USnOxkC8S/NimLeGNXY+3
lfBg4Lq6p03kE+GJtg3h1UIRpXj8PHNlQNLgWvjcqZyuGLpLo9pWPr46M+rls6iPXPZGyp69GDKv
+MmyFxOQ9GyDTBm50iaKCVVJsyIk7jyM0AZ4IP4lC6JUAE8B/Z2zzhbXy/wPV/Ugcm9PGhu2YiQ9
GdAx+WO+/K14eFFT5Dpzi5rOqHVdGNWMdiuBqgTUqKRU0hCjbg1qOII3E9MY4gUPr675bN6iLV1W
fjxakTMcROjwdPBk1XWzCbQqJZrVAGylct2vh6QQTwPAvhG/PafuOxInFKxvhcnk+8XQLP0LyNPt
pSPgddgkJ+3094L8RndyW3EpizaaKUC8T095XjQ5iuMWSnETBwcalbrrOKa6EYfAXIq8WFztbHQ6
1yQtGcMEuvWhA1MG5ZR9WPdjm2wB2hvRuriefaEALrdxol1UkjWcMyYOPvuIO12ebSCMX7qATfru
wxT8r8KDhdx76vFhc+zeOuWIJyJR3Od47bzYZ5La5MtdRqXaPSeN97x2GtTQo/z1+M0+8bKkWrGl
mMVsmjqyR60km5ASxy1LkefCqzn1hAEHaEhY1HQi0MhICz7l4XGAqbSTOgy6/sBuGYnVAERNlIZI
VANrM6mgRRkwildccFFe9mdqVIqb7V6qUfVuuZVRO12cFmy00NMETJepqyltQuD1wHfa3KwZWS6w
AfzTsgajiN/OT8C+tbQsE6BdNxt/mHN665GAeI2M/tp1Lfdm7nKs3sxnOSwS2J0duM4Sv66OrdsO
nc9IaRjUSSCOvLKHSWAFBxU9r8QTEYg+J7qwaEU2W7S3Q1FRi3WtpwQRWeUVxvfDgIzTQACicsmc
mawYUOCNuCDL2vdBhvc9lR6xQptXevBmBaP2QL6zUVxLBihWLTxjPhiobQUBT4ymjeKIa6euvxvU
T4s4Xpeil1vS+CCRdxyH2hbzNucv3kUAh3M8r9/nKW2H3Jpmi9GXqQKysqrstPO8Aiw24EPVa6g2
r25c56Y6OyD8OlZgLm9fF27TbqLEJtSZu8DdR8UD/eq3tvJTRRMepBWW3jDIUa2CT39vxj8klHet
LdweeGR8CQEzRpx5R5ltGVOtRUg99AB1I3CQtD3tGllNuGQoYlVWLWDlsCko5+0CHFjdtRkUjDpY
NjccO8ZYm/tf4RRVGwhcD9QR7SFAjjGU0fZ1WXdj17BLMxVG8ObGW/BNguBSQupKRft4Oz+IQZUv
Jq/5f/6a+IDbAK3Hf+TFEZquLhBaf65ctuDw1ACWmvF7CaSOkYlnK5+2uv9wsKxn+IFqnRrdkq+g
Bb2Ef4pnesSn6S1SLvlyca42O8/3NclxFGJyfmNiUuqAJvnC19pisgB3S8OPIYumb4vEzdOOlkcp
TIuJRAA7rvdRmZ9IjB/lUI8pLFUaGEMSN6650LomOicwvFAYFIqrDkfWQFrfBmwrQ62yi1TnJEGg
bpFZS2hJtwfWC1EZo43GNmmwOLWr1bVdc0SLFie50ZbDjTZKmy6AVhj/0Nf8GOlR6ZtcnudDJUCw
XozLxP+7viW+B5ELxvPiUQ4oxSYa9HrOFWvVo08iPZr1hYkAE7hjCqJ9WFLxlVPcHZSI6CvaAvEi
0sxlWSOw1xsgzoQZO+CQ8Vys/egxqRe4boyL0inZj33ugMq2HmcimFlmAsSTATarhy2lGvp+MTEZ
aBKBA6TvOKXR8pE6CkOgY2YYWSTeVjs+bU8HML1R5nmXa1pMe7pjx4d8QZOi9WT6Z/G4ZIkj92ml
1QAurs2mYP+gaaEilbWrLEGtLCAkzL1bTMVfVyuWx19pVNPRtVUVLNm3kFvUu/9utL0Sd3vwiN4w
JVEOGmmhVcGthYwSSlsxj/4yGJWvgLv5lRy2oZolG0gy0YXdJb6SwJ9sIx8r91UZIf0V4N3JYfp1
xT6E9gzMxNVOSxtJhleHBZCHTNvrhbCwllnXFKtQ1hhjFXL/hNZ2teRd+SZq5az6Qvle1w0E06ev
zI2sxzToeaNCd6Hr1IEta04rWt8T37ql5TJyKgfiD521stuRlxJVwN17kyjTdXIMdRFBQjcT2a56
5fQBmxhk7K08ESaQBv9/ZqTj8TkVlzDrv29BVF0KS0d4JkLkxDZ+pS8CEkQH8vERPWlnKOeNq7lm
1wlAUvvr7DRLzSq0C1O+R5mHy/1esow9+Lq2SD1kH90B8KtIP3bsc8hY/uCRSAW6cltdTeLeG+mM
1YIKg1vFKPlBcC9WyLhNG2A4b8vL8wxiabwEApNNVBVa3DldtOiCgHpsdjINngtmHD1tZS86oy5p
bfIwi0RmCQmRMWjrsB0qxrBYI0TE3ZktYeBDj2sQzBiOmlXFwKtdZeFwUnY1+eyug4PwcJSrahvd
gB3Nn79UiCltwAC9YlLC4/8g7OQJhgkDtRG3+UtxVAwpnrszd64nDAH83Smc9hBZ2XnvM5eAfIHV
m+87Wy5mZoqnCX9G8VNxpBzK4O8L8I5uslsNNHBrf/+27dRMDYIfW5iQTO0euc0PxVJlm5oDWtFF
9M35UtnzpRevx4atlj3GbdEexXKATuvMYyDZZmpLusRR4VQIFCasHHCJfYkJah/iiD5uSxiP5mPJ
JOhOZ4sg3820tsHTsJwyF4UR9IVAEy5sc5ozKp7DDhWN/q7dqE686e1Eyg9rD3A5924Bt0cfjuPB
uYyouF9fvKEffwv0X7VjkHyZsZrUZHDtNM0iXUPDOg+rMgv+/BQF9RavEjykRL6x3dVZAFIyzn4w
M8LBiDyGyHXuR1LML53bbh5DSIGjxrnPdiQ1XjImaJqWCXoGhetJY+cTWMWjEQ+ubL1J857KuOJ2
v0F0X+TXMRpp0uI7qAb0TvHfLc+tQzR+ra7AAvn0hoAvsiMzXGiifQdGkcsQFA8+u1cphTpVfVSM
bSXr5PHKgZgL6HyXqmfoBheWyGgoPy5oxs4XvoFNCMcbM2x4oZy068EIPzAcN9TLxbPMzQTbhZKS
uuJBOROuJlcr+KpBLcYR0RrbgJqav5IeZgYLtDyEKUiOmQt1KIak7xNPPHNYFQb/lMdj9ddHnM3O
fbBmFZ0lQyi+nIRsEhQH/J27W3UaDvvrDV7tWo0h2zGSzqH7/AtmaiQUkAJSTGPn8PmTQEncqfDV
8MShEzuzaMzoQCr4OuyX8+7HKI4pRh7FOX5tYfCgjgK056mm7dG5yiacnS8Bj9xQhfI5Wa7PMgmC
soaqqn7uxnpnUytFqoLxL++4aSdqF0p7LpsK9J6oyY7HoRUn6qXcHSzaWvR+qheo9PE2zgpd/29z
Czp4tVKcgr3xqTo/gjR1oJfIeOpy2OXZfj1OaIv1Chc76gcUQgxO9VsQio4RC+l1RPcAzgcVxlIR
YyMDixBY8Y627yMABqNCd/+tBO7+a7lmrFjzWsBK5WT34CZ3iqqyysllKja9u6tqJBILgdWDyotc
0hJlgWF1jIlwSP4v2i1TMK4jdgImOgf5/tqgdYQyVcFdV6muma9BJXQtLRPbstX3YcsvsuqHU7Zy
RQ8b0VZI/z7uDpK7LU2+JztlcYYsWoU5pXtUzJWq4igK7zH0dLBvsya1BVssaZH18qU1UMIKGCph
5Cl9423IVGMhJvklpd9TerbJKkGFqbroNbeO8F+RZ1lgayeIsWviz2WB5U7/OZeJIB78Ec5stvxp
4S7PrpsD9lEXeewmOCyEruU4oC3rrDOqn3x8xuUBfRCrWnZnRt9jdUZvsPTJEnegzo3bteXXdOWM
F1fRfg0BAUuLcVtTq1u/dMVrYKP5YPgqG7XerBqAR3d9IOWSbpOkRXhN5oBbwdU09XdAu7WE0ZYl
m/+f4btAEpu7/o6AOVrWFfHsAizk/q1+kiLAO5iI/I3r8K9wxmbTjtIVhLBQS2mOFASxXJtgXg2O
FB2ihl5yzt4RU3lELDsClVgT7kF9Qk53Vziprbn51yAyGGcQu5UTDYXzHuSyaQ15kS6uChW8p33j
hPsYOx/SAgFrvzTBO0kOFu9IsCftd/U5hwWMW0KySdLdrlctHBBVi67sJR2Tv75vuVpnt3jhxZB2
ljnjr2m/jmTxSxf3CQGdrMgi7UBaMlN+yoHjiwktu03yZ82L0Gbk0ta/3ApkhjZOiH1ybfMRvkng
tgSALRGhvxnegkr+TXzWJ8yDyQtPjk+XRj/vQs1/97macXFj6WHZqIHHyaWm88wjz5eVtGuXvf/A
atW5WHPb1nB+utCxm2/EzGkKHU7khJv8MkY4cp5p47esL+2a3vAx/YsYq/3kt3ZN1JrjBfznz8T4
vrXvCgbsxxaWUeBzBSwUIis7HAlBVemySTTrYYJTH8k/D4iZJ8LbRwFFfGSnRfVgO/EW7F1HdTkG
8izm20wTf0JuzAlRpZnbOjwJ19O+XlBqnbrQrC/KOz9CgLGF85IIYKG7TQXm5Q0iLCDsAgTxeCf6
wJx74RmciqYM2X8Q6ITNgs9D8SJRJB7ckH4ewQg2byVTchmYb0bc37QiDSL3utrBknG3S5ZSSQdb
ap/RJgtsn8swAsL0To9oJQgm8+5VOgwFMjfF7ir/xM83/zCMD37YIiwgfwlsE2MCYecElqOBTfXR
lyIgHXBlGGWym+4O8sSQfYvNN99mC9Zkvhv1rIMpCmc+VxqZo3FeuYQEOZ2EprypZXH+yvIcqAbb
lH5qDdsBDxkG5qqY0tme/fhoYlKCreLHPb3PdboJufWJi51xxPK8AdTmlLQnVDAzmmLHOBTUWq4E
J8ESaP0dcL+BS0RqV7kqH/soUuEHXybdm33ZWG7oz3Sm068SVH8lc/vA76lR3amfiBVdKKXl/cI3
eHV2Oj5mS4ugICzJbPWA7bpUwR6Vt1BS3w4vsMAjD+gq9zEagvrAGvm5D/bK4s67xjdL/2cOYTOs
edn9dxdbDG+QtzzhLPWB8bREgE6Zg2IvE2OdmqUN/7uYBOuHOpry8wMd4eNz9kiubL2lyLYRCnkx
50dnXhCZXLpnZR9ckqoRnj1tFMhEQkvqQpVo2KI0hs/JEJrzB0Kzymufx2MdjlekOLY2zkResZvr
uJgQrnDXuXFJe67K4TvOSeONSD3wr1+3YMvVLl8x4rM2H1mzxiH/Nmu9VvtXLEDxS5I6gPTbnWF/
4e/34uBnQKIL7BfRhBI3DNWUNygBOwtoX5ely/26LAVmGEaVviZJOywpH62xRG3kcEZWEDqidzsq
es5+5u1jyfPGTnKwCTCtuYIbVaRHSI0JBlCF4wgijAeEN8zmwvMH4M0djEMhP1yhCbKNG1zelm+b
U+suvbHp7x+bxP7r3XbVV5e8kP8SrClhc69fBvzRNkvVhUOCjH7PSlw2R/QLUbsrHgYhMkcZN2NN
raQ5EdaQWLDiM8JW0LG+KW53gpmhs22bI7TGwlZOG5Xg7YFh7LF1dKpbWn4pF41HctO8c4qtyBPV
Sqs/COPxePGiGUsARnoUONABpOSvTpeBRQXss9JStkbXGujlHHVbo7bfY116FTOquVAka7vG2xl4
V2mpG+njBmdrqAr3flzEv0tW+v8/D4ssuzIkizrt9p8XC1ylnL2raQBf21OysMbnBdbmR3fgVlP2
dwsw9rNDO396SXDDoyUYsg/6qoRG0UKlEAvfaXsbmlfXUlBNNBr3vGftnJOeGHx0+y9snaDeY/3L
BHoXOslBkw2eZPONZc7dJt2IOiFuDQUBMKDeIiGI8GlLJOpxIg+WaUKfY6WwK964+KLjbDdZzIlj
UV1qOJMZkleM8zG0Mk4F+MVCKrQ6gV5BXgU8AQ5KjJANXVbHB1k4V/yNAuFGgLqwYTavbYGca0SW
io/rxJLB8E4wCTDpvtEabk+PuWx+lT07/dVmEtK/L3zTIscgDaNAS4SghoRukbqGthhNewSxrz5X
oUWzNcq/fOCyXJIh3rFn5A0CcmDeUm7qBJwAXVu8/QxwjiY6r/dg+JMs/cJxnUQBP9oDq+SK8wLC
OVvzeW05Kw1JDnBGXorBm5Vet5oiDazh78AQTlzeIvpKdkPLKXiIjwVNHsaS8nrSTYI6VUVSRmbV
15gMk1rs37eupmpMSJpKyyQXeAZVIR4w2q749EAX1LwnXt4+vP4/DdBGLi9tI3p1GqxNAX5y+F0n
WRyTxCKICZnNMSHpb4kEnCXbVbVQBa0IYgeORKsdb0qbybsjn68mnsIZ6MX505F7/TJ9dLT9B8xB
g2dQP0LiyODQAKdQq1WjOXCH6AnhOeazdnlPXErOJxRjbg0O9a1T1hCjUh3T5TJ0pESW0/vB5ARv
Yugerrsx1jUXxirbUD5+pzlgGCgnj9Pox1p4sRy8bP/IZxq0i/1YgZecNXLtUcugfWrkB3tr4xgT
RQUsRUL3oopgKkoI4siUfZ2+M9HXqis1bV+0iGu0um4Bq3Wr3SA3D3J8hKh2O9781OiSNlbLedN4
ohGUK+P18DJjrkLgMRuHSzV+BX0809S3SHdrWN35A1DXZjDPdUODjfSck4qAi2cU+q1ShWmUMMtZ
ELxUTF31Py0glDD6IyQSLLEE9DSEc15CqkbHwmgyKs64wxE9qkCXuZIZoMIx0zptAuGleZcV+MXa
Mgk+AWHPBfV9lIVxLpdblF+8YhuWG7iRBHz89ckTFcAeZe+cri6ScaqeHkwmYjIgexEF3j3jWWAe
YTU9X/VVnj0BT+I9TCnfSNAwNLvUDPZwu2V1kQRoLy1jJRrvDSbH1hGbyOOg2xcmL+NSkf6JTPVC
bCIdFDCfawW50p9LB4BKwZ58CLwIBBSj3WY1Vjiz5/HlG+9nGdC2DVpSjxsrVmxe7cTTMt1Y5fkQ
r5KuVgyC2N+G4GN29EdAjZtYOtyaXlaBaZ84B+SPxHXV04jf79LltNvp+tehpoxWNWg1JigkeMFz
mJlL1VkNSdUIP3Yq/+WESY5MqqEGuw6ERy2N/wEI7IPO36qLVt7WQXbpPgMCg/9DtDfa/btuzJJg
CesNVtJb9d4jniuHvSVVoEiGf6Yxjb0dOHbqZ13Hvoluuo2DDDg0C2YB+eB3k6LDW91IbjYYIg5Z
ZVZc6oS+c1pAF4tE0xLQ1E3ewkKKPEqmYPoIshgi9dMW7KVS342jqR6wSPVRZUyJtkB5LgFK7PTx
3ZDhVnDGbJHipFO8mLpd9Kc67iIcT6WDkXx+xTh3kegey1C7NdePvwOdq6amZeb9D3A+zg5ZvfL5
H7ENYZPUjFChP624/cipMDHNl2SRMaZhkpe69JxISxjSnjG1pI9DoIe5deiRhRAwsKw3j5w7nj5m
MjyhpO/Z3QEIsQFphjJAXgShyPxzPmIIxEE9LWvT70iv7jLGUkxMRd4Tfr2Xf8Rcm5Dm2aTqiKwD
J56mIidn31R14+kylcwE+bBPu8pcqqp+5t8y0yZwWE8+z1nxCPjaASvL1iqT98nGOyCETXuBdX7u
Io+HjqAEfJFWuuw8GWj4OZpD9mp9l/E8AAKLrU0vbM6YreatJ644y4sBHPI2bWH2EnFc2AtfvfUV
kci/+ag0Y9V/bcF1Sd/j8vXpedwNWCbrGET6dOgD+T36aQ26qcb9s5NbUnpRMZ6AATpk0mz2znrj
Kcj92NnFI4b1BATVzmSKmA+Icwg7XHm602dj7PWqzMC/BasTQi4l0/bRkE0XAV/9cmW6qFbaDFdp
W8RPKjaFDK+g14LTknNDWTFoZNdJ/IPOyRPg2z/Z09UiTGVdr4HN7Azxh7fIssOFeiArQNMALehv
DOtuC5hkxgd2/Td173fzKH4AXQZNw5Hff0IMpK4QEejkYIDBuc+iFfM9+SPjB8v/yUF4tzlnRqyO
FvHQezjql8+ttEHenGdnatdQCUvFfgVkpsTuisMuQU9vy605tOWRoSlku8wVdNezSOvkNSmz5yKL
JWrzYslkTFEmtHztuTZr3HYKjCp+PJQRlnfS8issyV5/+7QT2r9L94mLnKVdrcX4jHH5HZumtLcp
lscuOyeoepFfGI1F4Y53J5It62d5FP+krc3xbW3bnGcEX3z6YHyH5MiNSqEcpEIGIBZihZS/yI9O
knavIlwIXf7s6coIuUevNjqU4xTRTHjH23xc6gt2Ku1EzqKf1inG/obmkXaF2Q/KSwGwIu6mIo5X
3InFo5odzGrJAdQREGBbz+iSFCSOk3aX/7tuHoruqJI1f+9c2IGfhc16vo0ZoCkuLjoKLNGXVnmV
fmQx2S0dcVqCXDvhVw+qayMMfUhzHv81ICu3HAZOEcXsrUFESDIS1o+hbOzfuPW3hV0oBZzXSDSv
0ztJvjysRD2z04Ua0ba+FXy6hYEh62pEuOVHmwSAEaRmK/nw7sD4mlnfe0DMRwih0KETBSTgS8S7
X/DrEjrPENYs0P0z90Ckvq3s8/9KgU0yt/BSshHLM79jfhfF6l299Q+ZpvrpY7kVOHCfdvKOjeeo
7q+xQDbncfNqgFXvoGbw2kaUnrNxnf1YtmijvXGopqW54lBo2EgFIwjl5R6KNiu1BydRMe5l4Egc
AEJwsRa898qo6rgBZYo65jP03tLVqghkov/gmhNfcCQ5w7z+xvSDB+kR3fDfly2rYUEVcOzCGfaJ
MO6btTCCmU4CEncgihik1NPEIed66F+qePn7MXsxZ3qu30euP3gvJ3AX/UsqS4/03Wp7DT+Cl0a0
nIFfDei9ouIRmapCpxZGiJPPSbpxlkNh0DB80GJiUxE7Q5aP6doje2PPLc9HqwoVCU+ZKWGTDQ2/
um/MdP/4RNVKt/o5jZStDGJU8sQ5bXcaKHtz40efqTGZvL7THi5OuOuqZf9nUSh+hBnaXlaNqm99
xOpNpPzhMxj63JLUyVyn7gFF/Q+awhj4B2fhsyWYmLxNmO+mzAwzIrICBzgPzbBUt9C7BdI+Vp1b
3jTN6zDMPIibCZuG/r42zAcQYFc8c6OYxnH5hkn24JoJ7eYzrTKmnAiTqNmDI+2dxXaSD6rYiPr9
gX9KR93jKcpxXd3g/JQt4sFr+NIImdcnMMdHxLKYge1+Ot1aETiTL6813GCzRluJyZgmFzDCFhAM
qB/PiXfTYbZtTchIadbAZSoF7i46CvjWF0wchkJ3wDT+PrfLbXGKwGNC2R7OuzL+Ddii/mQA2i/l
GDd/UbUh8smIVS88mhCS+ue9cLT2H3FcRB6kNW/VrNO0ItCzqPOeSo6iUD9on+buFRmdbC8vVTvg
Mv5zsOad81MHXPOkjai/7rbUDpJhHyuwFeDVpcJPK40dYfTXouFLGDfjHDfsh8E+4Ms5IWs9LUFv
nj2v2e1jKCWcRub3yK+fzmmLaOng0FSlRapEIK0uqBJTyBI8yHsxuPe0Vwt/MDPfejige4hHtWwg
9SYug00T0nATSWJDdiueV6yU1Zu4f07a++022qkyg6ZT+tE2yiYV/eiQcLHenpn1FaeXuAGzP7er
3HET+sS/bTwFe1rktUpP17yWFZnoni0UM4MT5H+MWMNU50FWInWYBlNieUA3zxIseEDrOwtTZeEh
H9EioniysWajFw5W+MjEnv6QZJzNwrl0FwMzgKtodticnbntslLKPalLticG999gJD/eq0/8+azH
HJfqWdqpF7O5rDWmyDAzuw6WTrdjllm5bVfIhy8AG7jwXkCU65PdtbE+2FMUSM02kTrPloh44rIi
WEGTRT1yYpUArADpwaP8tAp2mhCaxLwgtPKoSKDYYlwE4IL5G80/SlMR9VGPxq5Of+dx4JoSFhb3
g3y+GX2EZ85AxxTzLDjL2mXLaQcgp5OdEzb0gt4C/UTiVgXG3zVHJHOLmWgwQeDo0Uei+Q5tSQiz
ENPH1ERbqostObnV7I5vdwx1f2RGC5AHc1zFvhU+LY8O5EcLrEDt+ZczkVuiOr88a7W50T7vv5Mj
YZppSdngY5QSKkhTiVsM5lcZQB5iUSryo0b9ei1zvGgeMlSiPyopp7yck4wkhE7NrADhmafHJwb9
u3IyowXtNZoIjHk7tLWim3r0h1iAriild8T2fj/dERmnZqDfOengSwwbgPojxL0wjU+MLR4qAIZC
OXFJBJjMi1xL2AhB0yhr6Jzp0Ejyati1glrfEStjznmBWvhcs2eYmiGAwhD4Abl5h7G2hj7gW1MK
N7UCNhDk3BMl5JpAMr0Fxp3kVQ4+EUouKANJGl8J3seIMJMrWh84ZIPOW1R34AG5qVKfHT7BTIFi
sV6iOAeu5wibIsrkgKLD+9J7HNORovBH/LzJwiYZkGccFTKG04/dAzNwMEtyisUi5pXwCz7S4DiH
5Mnbl5rMLLdJ9XT+/VPbPSuzyWneRJs3pwywprzhxV1d9YSRl2d9XTYWB13PcXQguJbccMZAPFij
2/yn++vT2WMxmkSZM8R9vAuzAICvmn4gAQ+MHiph7X3Hf4X8LLlNe0652p+t0EPRKakJyUjKh8Qh
veY8WQ3iAm12HeLPM4E/t4n3MpbTz/LcW0Bpoc0JbAQSrJADrd+73dzKwK7yYahynTBWX2FgL7RJ
wai0/VEBQUEtbQGLvW8z/dLS88NQNVcHoQBNmi8I5WdanEFTuvCwM0t7ZycDJRpwiLayMBfbDhoq
A5M8dl4aPLMgGrMKJI6su5czhawS3LLecImPaqAfU5leLUnj/J9g9I1okMd4C5gc42XXyzDB1bg6
w0Vf1IqonX31b4aUY7uOJ/c1yxIc1oUdPF/p9gCXKZTuvF0r5m2/B+zfoX9PJ+Mc7AE9wwZRPozD
WyQbWztEYBvm8A+mmZr3wO3aefJj3Yr85FOulp8Im/03FEhhUZLh3aVQnC+PzilWmFPIG4+utfDf
lxVqQcwIrzKz5wjRv8ZNxZly7Q5JxOC/SvisnW1K0gURmgcWzo1nqqA/3CJqaCpagzucsSkuBLeJ
+Ve5V9TfbHoOALgwshUbrQkLD3iXOIu8yiWPLZ6EluTcCdF6k9hUBAN8CdlNqQK24Alc8YG4CmNY
ZtSGZTc1mI7AynJh2/AS6sYxkVhIGcfqFfjZoRpMFjrfBSuv9P9S4w4iy8ZoCfCMA5y3OHBAy0lQ
XXMt4ucNoeGMyFF1xPhJ3nbIMVqPinbvg4S2gS2jIA7vS69PHwADrUrVxdau1jsNajPQdXuGi4x9
p88iR1+8boaJaw/sFoxn+p9FhKQSbVsPID9tL051Y+YNEK8wFURgvHGoqg7aO9i57VtEAxuafyG4
LZ2eM7M62ukI2pMDybeQ/alFuvrdBXQ8md/UAP3x9ai7An4ty/q4zuPapK1XLhSM3IS1XspC6vty
2bKCBfUE11paeGj/DgaYJD78qEzIAU0mJL6diDJBqEJPvRfr0jBaZsPTkvvLKR14aWYIw83Wm7VT
P+V1n0umsVKdg+P5r5s2uhIlbEf/YXftT0mf1VCExGpwX8DkKnn500duBaX+gclyZVhodQcbdTCc
OTCOE/EbH8a8ohdxPMlflPho65pZJAhu+SXzkHaiJLwBR6AeltjrL5yKmVuk7s54bwrqj4JDXrl2
ZkazLooqwwKocD6Z1CsPTpQwRLpjm2vHBdUKqg6LB1Q1bC0aei9WnwiywOdh5jpQ8LdRfSZdaVl+
1udbf8vCC5LeRoFDcCXNakvrnUODFsiBRlxTJD8UmNLWkCrYuIqqaZ0B3Edl+xMMlNbp90VGBYUv
sSEqcO5xwPpdP2DnjNkorE/KE7eLCjS2zsAVWPHPPbB36DtGtl8w6kUlUK89WoCwQgBLfQMGQGq8
V32xkuKFzBIIxArQ9TQZAkPUlg2++iM/BRqz7m+MRRWlllWL6q8mmYAWTYb+obUzayMyCMZ0tmvb
En5PCLQb/fu6Gjvrc8ux4fTWluz5wDEjFht+FinWo7BcS+2bGFXR/Z2ipT0URD0LHC7wYBEgMsex
a8sa67mBW+/RAKzoPy+8040v9eOB5vI2lbC1cJkh1ypkM4/NP9Xf6mpDwFNZQKLofx4jGLwTJcE1
jjST5pCZSYkmGoNQL2R+pYnMp5Xa2PQVRP3N+lcSS6cHjYmPCo+QFuhiatXQtHH7sKKKi+dOwb+K
lQ4ERAopmwMSK1MzMsExOaq6YGCRmoYKs6xztW4SQK0ji/TSHyzTv5ETJnU8pdY2KpQlkhlOQZAd
LUkLnU/zEXloXeo26cpZQNILtbUfzxeWpYu/r3ujr1ccsY/e3S2IQCTfMhzDt95XGbm0QtRufXwF
Lxwb6dTdYcXCNVyOcQWajUeahog2QQHb/pfalHtojdJ5bZkQUgffjNItlQJ5OfWg+fd1VtXn9kPB
QylzlG5lXdjnbW9GDal2KJvxVzZgmbZCwu2o9AHmYLdIrGxUX13SgWjWeGfew4kMUxTNTGFSIbEa
8EYL9bhliWC1jLjS8QBZTDU+o3wuU6Os48/e+i3wIMQVPM77KQ4Kvaj/4R1RTBTXN+xU18bsvdp/
auRUtJCdlHKEelcMHf3M5UAC4zd7FNlas8lh7vyxIZ65Ra1uKUrFuNxsiN9VVhLQ56KjzlDFMPBC
feTCrlTubJlrfT41BRQp0fc9TtXrEJxNs3HKlewzRDYHd6e9XrMcgiUhMSoXlGnFV5suWr3FzlVg
OaNLBEpUYHq8E1hVH5nlR2dRV43qykKgtIqE7bI92W377DgQa1ILDDUQL1ZMSUvD8NqmDzYjaom0
939w6prokkESXb9PmTLcSR4Iyead1f7v84bLGDxyFaLb6JzPdorHFeePinbFuxRzr2CxAtgnOBl+
IXJDJgtFccJILufIC+H/5X3wugepQXVNsfw7Lak+4+H3/6oYaRyK1ZdC0Q4WEeQ+V3fpZZaTIyrb
poHlOzUvPEd/izHK2wT3Jtxeb32v2zNURtWMhyh4qKxjFVRVvBrdkoBl6uUu+xdpB1VtKSYp0aOS
IQiSkgH/vQfk+VVJntuGe2jHyp7hjdj46zZ7FJzkgBPydPI3a8sLmdfasUw0i/R95h3sWdWBPfNI
PM2OxEKmTE2WywUqEa2iGzCbufjU1pIQkqWr+389WHP1oI51lL1eYp8VYklk3UKmUp/Q0YqWridV
d3l7bJcdHpluwrXpwdhOpH+y/XsUL4P9Ocdr4JhdZlfrq94bxhR/xTv8QZpFz0eZdz6mbLQ7Yw9o
bPqq5F0FNXJpAfzKkQfLotb626B4j0fWvZOM6Eo2Uw8blAyCcWgNyEyz8bpE272bfWYXS7AOlmuj
qxtzoqmpnboZYN3xSFXxR989sPj4gf+uToc/FlwCLmqQ+XKophUiLPap1kZLf5fg0rd8foNvE5T6
CJMbxAUO+myHlGVletIfiboDU6j2lxNMyoHRMunC/yhoF1xH3ktYTQCpvNFXFc6dzY3Tns6VfXDB
dSxvr+xJP9il58KT9wn9FcyYW3Xu0YbqhyWQLjQTHjTtberWx7eIyXsrzm0Td7Qsv03mzew66z/N
I/xxGyc/P89KZ3TE/F86rV/AtWVq/f6PcZgR27wF4DDV1AVqQSunkEkZgmmmPND9xDuwzk+3nbvm
eDMZ9//bo2LhGuqJ9M0wmMu2H3qHSV8CeLOT7j1dEVupK2V2yYNrkAkrDsx+yBTfEtqnf1Fn8mpq
XQw1V251t7LmSNOAOxxIAbFHprZZtnYDupyjA5vbBPKBtZeBp8X8aUZ95c5ev3ZPogLwQLJpEMby
EH9T+YuWof0DEoCFE0SGASDR2ffdIc9gBDxKR6VLPeVntw4W7U82IQc3ph54+YiNJipredm4CwQ2
LQuRbTl0AMxpaL1E+xeF8+gHsaU28JddiQ33ARa9UnZwj7bkRfwCMj4+n1WEDqHz4Mc7MbPJGG8m
qEd75xX0SPJ2yWI0lReYnimD4ZSfXHxpLgrkpXSpsZoMcuC+fkf/yyBzMCzg6iirbzKzJds24crX
GHK434Lc+xBmMFxvSRefoEVF8qXkSBGOD9R4zweuzBci/UilIiWQsSPqHnCfZiFOlmZeSfRg/SXk
k2fZvFyupTJwMOQRknc91z5JiYm8fjnlQkm7JVwwQBxdb5npaBIVYLxa+DCA8vW1ojK1Joq4lg92
FwqQC4WuIichHe/p6G7ABEw1vGt/ngUEZf8+nKGtF5M09rK4m3a5i2MKHlhLH8uzurnjYa3EnUD+
wRj7Md3ANb3UDzHUZgLK5wuNMC293pQIo8lKo2vMwgjaM8BdLWLC5E64TzWjIZpTQgjSJhaRON3u
wCPOyuFpKIJQ7EmnLAt9ndjqzxhk/9jldw6GKzMOg7jNHquZ6I1fFGpM7nZSUVR0JQTkc7ogn6PI
BG6lvl38J3GOSpYp76Q4WADKiwxEzbXNpL9ZQoFEyRhSANLFJObzt/N/sjTvvk8vbbjGivABTPgc
zAdV4byb93AI7t6TxI8PklDq+4qS+IGnn3tE6XjpXbjpeOqqbh5yrlCQBeYJL/aogU9AYnM/YMPu
LaOoIxFYy/nV2ooGygqIsr0rIr4VwQoVDzkt8gCfCgeqXMXzZn45ZmLPOvhv6jywNuhLLqbPo0vk
kynEpTkjvWH/uUmap34+1iLfr9Idl8mczKEGD0Gh3iIFJhmyVuULPuxVODdnCAxHpHZA6ln77t4f
UCAur8QcrYmT47QDzNPBIpTg68Z6FiJAUT1/lULXe/mm42k2jhflUog00JjCuwRiNYOqpIV7yyVH
3FqRPYqdvjLrIVBEH8OxXTCP1ufp6ehRF70gIaUpOsVyhAcXx5AUhNYaHkQOBxKWlBnvrOUWJRVO
/dkpaFwYF/n+BRzNyegQhdS4yI0QoKepiY2xLWQHmK6KTE0qn45tx67LGwVx4dtAPAY/8YAO90RX
7QvxCuqyNOWvNEYDXmym7F1lsB/bwvNYsxR5X5TLI3hM1LwepFpdXRs1lSsf1vMqx9alG7ztd+xR
QB2E7gta/fmja58b3tDMXYTEXDHrLrLR4495Ryz+aiwazQhFwbCKUFhuZ/aJyw/ENhQcGOcAk8YX
qi33F9ssAzvLIvPEGvePTjRwTaTzDVeVcuiGmHtqhvkgSkoMlaYszKdiby2E5mukDIiTDtdRLVhe
cdHjXMD6wj1d3plvkHaKNEXNWw1buxpahMASjyJ9ejIAS6Iae7Dr9nCophyqz1O6nh2Tw0Tlj/8o
80uV3qjhF2w1wlrm4lC0ulti97SNOo6x/+mcvKYZVkULcC7SkWFQ7KNfenrAFu+9Fye6NHlxjUTb
6U1FGSDqz632nIOx+s1t/08SivW5F52cFpHOi7hmvpv+3WQmPSPf/8SM9vMh5RGM/q9HbwfPB0P9
0lWur1L1rK9II6hGp+PX93kDDK4O7RCHeqSxdAOZD/Cc3521GxH9SK7wH+u1fL3/J40Va4117OGT
bG0xEILvLksMQyanPVxud7npWf7T/8Wlf8kgK9dC96NxU3Q/biPdG3fVALmu4x+i0EYB+T460Rkd
6tSCH1FPXs8UlPeTpoHJm6ob1CJloLXGil40MVr3e+Zz5pC456+K4nW/IBvsDssIf+m6NJ63CZEM
yRX8XnMVD7AuhDQiWWnQFXQvRDe9+e/32JjxhsAhofE9mCRiymzQ694zQSfrbU/X1vHb1KYS7iH/
I0Rg+ONDd+x5wWEOWbyoQhf4wgE4WGLf+JY0j/04IT8aUFIxaG69UNyadP8rN6ACOekf6pgum01K
DCxFunolt/B+P2xXNIO5f7LQmFDDxyuY+fqWrQAhhGy2iqyMOOruziicSnZBZSuntx1pXuuYGlHj
sd3NulOmtpQfcLJzB4ltrIDh2kTjFbELp3VvxDTt/KWjhpqf+45FHd+7INYfcnKGvXJdy8KM5/7x
apESpK8Y6CYQcYMOP2b4FegU9Pw76WCOuazwa1t62E8RuF4plmKqeTNY0Kxocx79SUX2oioaEwmh
yma4hegDdsKdL2hBYT5sUKWU6VzT1/ckzXFBUEX6qsyZz4zxq3uR/P8jz8Yhyx33XyDQhcuduvUO
+qibo3L2IrpiNXaX/6kiKga4nr+XLMmHikUvgojq0Pd5DIKWJB+78nd4DkQK4Qcp0pF3nBxLDrZG
2wafcG0T6QesroWpfhycE6WL9rx22ERU4fA8+3iiRRm0G9zW3d8CNC8dNiksCWOw3Otl1RBksmIT
YJE1W4+BH6ufNrjfPWsU2M9bvz61Zgsi5bhk/Vvjsm1+tPEUFk6Q2Bb/dLK1LJhH9ajquZ6k/O8y
9z1OJmcmj3chQb5MOvWRjduhOoBVmnFsyT/XOQHH7nkuDZzDGohN/SuMeHIY5F6L9ZJ7xAmlOZEd
B+fvqSEdYOigTI6nCVsSYFxUswtG+k1I8PS1MvdtI9brC2WIdKDR7obFrVl7z0SO3eU3NmvkvOJ/
vUyOK/xH9/OqdtQLhdi4MPPA0EA/3aADFhhBNXmqmyPghf9N3N2UXRSdeItHy0B2wITp+mmqst95
eHAv9BHsIYfBaxJXBjvb/aeCxBM3jhWkNnQ/bt/+gzcNLSBNsoK6uZVHc4UixaEc5c9RboBnG4Y0
H/HdgX2IER3VCoyR+V7JXikuYeeCroU/3jLCJYYg9T09yM8/0zeOjBCar/cHAsWiEDA7SpPjWJMv
t3pcGjqYXakI+hbaLA+/a7rFY6rCCB8QjotShZRH0oPJhJpWVBAX2N0CHm3g5pj07JJFG16I3J1b
1GjQFoLz3Nyv6HNAS8DV5kVcJE72T96QczOOhp1i50f8jAcBlQU1M0CZ3LmTTT7fQG7iI0fLkj21
ebv2BVfNgs2LsMToE0jlvqWvwOH7CtFe2EWEBwQ7R2jetKE9Z/jbvWseXFy0QXGGoHMzi0tsQcMk
gYDnSEpWeoQAtZK+JHzPDeRORW4GjinQ+1x8rz89dsebiSB5fb9BKF7/43DzmwbLRusiuS6t/O+q
YHDHL4RejbAx7XzpbVmgzvljwmsHgkTdwuXNPJq5f89ug8S/UkrsxIIPP6IBm1d+Q/7w4sSF6lwT
7RDhYcs9H1gUfMr+LsxaY/OkduUnEu9ZcGNxKDJzbQSrhi1mIDXPDBqD+dQkmcF4KWeeOEL/938Q
IIIE4wasv2DSYon4GcIJ+loX9x3YrPdwLSL+suCFAv6y6PdYL/JrX2zaXvuY2ekyhMYMWEvbdyhe
nl2IAklGQ+hyPjmPrPWiFYp3pWiscK39CEM2eleoU4+FQJdngETEGpAQpKqamIoRHopNj1kavyi4
0Q9QswOZlEtpUJb2gQ6HA14iKis9JU/tlh2WPB2EcDqgOqosYDdJwaTWcR243J9rM9cS2NM0VkJO
QTG98cqTgkQa5ZGKwjTLEJ3WX35j0f9QCT08c2Xcla59bpiZKV2dVC2bExlv5oPSihtlejlxoCyH
3jd8zj+zr0I0sXwcpiFJcN7nIHHYivofrCvmyXuTUMDrY+XOe18yX3Qp+ZPBjfkHfgRy5oIWe108
g1nmkewfRrtJc+GSmKLXN4hb9lMPFwYZQHzZhnLxuWrntf6GNEX0E1U45yIhIcyavTnOfjWNcb+p
dUvCZQRqGQfnXF8y1iL02E63lDDdHypfWB7aXtJ5Hs1IlLxJ4bcDsYgVaQ+A2bwDT82Hqlx/oce8
6G4jeUFFA9Kg9vEQA/X4dwumEevYAowRECO4jbsJ6euhoHb4rtb0r963d68Azl1GIrVmNQRWBSor
8vfcbzOmVLFeiM5y7hwAW7NTIApgJf3Nzy2uOsEWf+557mZ1u/eJbiSsg0n9GFoI8TKZ+AZblca/
3IzAaHNQtiKxW1yjyNqRZGOcsd0/XC0B22j5L7yXonXzQ5kO54QBR0+da4et+a7L5WhIv2HDCYPP
3pE1/9NUYW413V1jAMGECcqZMd6XlhDM0pOPKJQCjTLlLiLm2XPB19PwX6Mf/Ecb7t0Kvdo/0aPT
R3PgXU4EiNXoHhu3GQMDj0MnCeN3XLVypk1skqCn44U/2VE0/I5AQUOfaf010bezWhsMh80o9zTx
f7yx0LAeTd5LKm0mQN9O9ihD5nUG5q9thJJsySGrG/aXB9rInLJNwMK1aFgZi9YLT4M7Nb3gL8Xn
cptaAbaeZgNDzgvO8ilqc0IS0BphRRanMeyyYsZadRQKeNP+3r3lGTlvYNN2B+CysWZqmxImzUgZ
K8zrcHTUU97LQezBTqusOMCf7TwHocXuczkBUwAc5T7tqfcKk3pMhWQ7QQv4kGTs3C0J+zGdbUf/
Kh4mcX5PItehN8BR1cJrrPd5B3OvQbXqKFeqolAI0oHtdSTe5xyX+fVzXFONKb0+vQPJnxRVUNdE
42Ovprp1yPIeGWRejU2txbh32eC5IenMFaYfZj7zFrOxfWZzouosBVo45+c9lvBmI39xxhS6MyCo
auTf+6/uoVk9O5JdZNU1CDxxTygE+hPjD0TtZXWCSr8bK8FfSi8J0XQR+QpHWtht7VRyDGjc6UPi
/x7AAt96VJS22LqcH46vETMVdgzFzQz8+aEMS8A6LAjgGV5R0MGqyb0ieYT8wKq2Mo9IDHnTd0Gi
iSVP82011PLSOeoCnJxM2fcLCmDnNmfZxZ2jglwgESRlSaYEOVStORR6EIjlz+NxcqB5wtMb14AT
Kp7Vfsc+88Dw6R2D+JJXJ0jEOMFfAx6UTwSzG3qVRewViv47KIFOj9abCGXpXjlCNWfyvbVkprYj
+C61S+UTi8sUalu9nu1GGdnW5zi4XBVC7SEuC7medYttIuYRl1ayT0QIEtJbSXogiqGgT8ARykA+
PpzIPjBkPbVTal8/pnxN8r3lDXCw0aeabsYM8yn2yEQnlLJQ7pkRwCwivyDhwUPKF3qKyjBPqcfv
aE0ywwb4cNBU6wAFzbPIxxVDGo91PaEJg7pPOAd1odHh2d2SxNeSmsLYPyvh63nNYXfNKAnkdnP6
iPlmv5DXNujPFAqs2qVPQ9hZxDyQHMfQYvS+EXSU7TPqKjosEm6PoDq1YcTRC0eO26cX60A6gvFB
mpNzINBYr3MBcWj7cWSlEw7ULoDmroUSFw86qlme1im9Ghk0F7FeQKito6f2/6l5iLpdctTQCHx1
SSA+KS404hgTbxc7CVqdrg5sTazs0hCDZpGfBziC+XZLMHgIMsw/OGg5Dbqci0i+IszzVQcyD8VL
1TGLfYS/1hF+5Ysrqxmf1ttA3f176RQyK2FbhOkvV2P2eULEMgQt7+pZl8u0SoplHt867zWW4czR
iZUgSqlU9ldbFGiWcneUniwG79TmeQyN4z+2Uienq0G1zF6jcma57p/Zp0L+CjouZ2xulg8ZRt09
jkG1+GK4Vmqw0rFKr5or9Pfbgaksn9NNp8T7EbfEH3St9aWpBNgRu4PWtyvm5peYR+pEqorkhcij
P3qoEM7EJgd7SVSno6g6mvm3+/ZRVFYD1HmLwW8CHS7Uc1BYNvaCcXM5UGfgj8w3qpFMM6SluDCU
Dy5NpKSjRrIlmwbd/X3pcOz6T8D39f8sGZvkYVbfuSLcczF6NaqG4ltuIkGjoNcjamwbowZEzJOA
oGYUJ7bEyBcpVkVqU6ciAQ6ESVFERqJnZPcHJoDgAIa9V/xu/UB9eHslJF/PGfoncQz6JY3NB3Oh
JnCdZSp8v7sqJ+zZ56j3b7wPgb3p/+OH0X9rYZA6qhrEneXqWYFNUMC2IRgCZhgDWWGPZslOy6rN
nd+cfLRxfhIg76elvIFAAGzBGaQ+0a23AjqRzfZkbk5CaWibC26cvh0lL6RxKNVzjPkZpsdsqk9T
j5mfItz7L76/rVERVwCKYVdLvpvuGS36almd8GazYo/gQ4eWsX0XvF/FvTt/xNGWlVTaBKD1k6KN
3XcMO1UyIJgyC/j8vxJ61skPPTeocjaChMoXIbIm1NFPHQIjkq9qYF28TO5nEJ08WX8bDyDB3OXY
2iW6obwTsA4msczxFcjliZYW+yrASiI0edjE53iwGyzQ+XxfhXqZegi5AVVm6EqgRjogPkxqdQwE
qAOIbXDvARju7J5kTYmFhCofUHlah5bBZ94R4rao/I4dLo39xK96Aapj3EZVBUeIwAPBcIDMT0Zg
vUyWiReGWbazEbRLGXghg1nh+Dk745EZiO4RG2Kf91kn81PTil8SYqG0R0s8VqGJ7EphXRQWyhpG
y8nu7hNvKNgbF1QTOvMcQ9ttaHdILuqrsCBefw8SzMkpg1G0tp1nmf0d/47i/+FuNs5dbgUc2cEK
hOb3DUG5KUnYc9Gq5uiroZWp77275vlGhTVm19JUQ/Ca87bEAszXOgC5NML1PRRB1M8FfsKhH1WI
oVWBaf+3EmtF2YOEqroe8FaQBFVKST3jXPKHmdugHzKa7L6s43HwbRWiB+vR2KUmlyr8C9sdya7Q
NGRdnM5dJ0Mn8DSpFfeXdQpae4MoFV9tBtLeEgVSPmnyYaW+JzV4ROHMdeocHAqxVf62sxQGIeBh
jDdONduNmoOlcsYuYTAg3qfHxmRioI0VL7VXZLHKo1rmHBVgPB13Sf8N5ClKQPGr/91fjg8jWOj2
cE7GMGpC/q6NITHH1T1b2YU545AhV3w5I6m4LV4fzfRhYnQ7WJ7U2zvTFu0Qtf9+UbheQKyVM+tf
42YMvlOT4Lf3+ec37eCxk0tmZQ54zoCenliDEqmyysQEESeNzuOySk8FZPbEfBSOy5qORHGtP9KE
Cyi7KQl3dKmXvgW1yANmlrLMy4s+Xs8DOOHa7s1MmG5lSLrOhr1TEAXRI9l1u6uEGUIae/4PoQPH
wvYQtvzxW4iPawQ8Om1387Fb8AkBq51PPaTcM0ehGVH8PTL6MbkrGq113S3tzJtm16TWXh6xPZ28
70my1f658phlAqtbM0L83iNexV4meqpc8fzN7xWuRpR+jf0p+9W3y/9pxS71dPV14nZB5LmRkdfD
LZModpA6Gu6Rd9Etqyi3lVTCkB8f41ua9l90uV/UKIkJ0wagFTV2DIx7Tw6FGWQG086/iy2YakM5
394eWAt2t8t7XPlortkOxhtyMGo9X1fUMTtU+XNGn/n/7gN8G5MsNtvSZ3FjNlC4yzoEyfSgvZNz
fsaQiEBHO3XL1IrCGL4k601L8jSBTTzS5qOaF0Aces15ekELhacjSOzdIPZCf8c289hrXmMn6P/g
fr+4L63DLwhb2eg4SOs9uROJOii1DPSsVluXci0AftnCgWjzw8NjqwYwoFr+bfrephpULJdYBB8h
uCGx2n2XqbfWC4qH9OebDwU8oEX74K1Owz3ml4Vaq2Lnuj0Go7MZwKJkDwsUIsQ3OsXvOqMbqMWA
rM3ruXZc+ppHs9o1yKqrt6A9qEp67jAByMj2PxKxcLckqFJI/DSykvAj5V1ofqfEl86skKt4vbiH
9+eXV9uB6CXfXXuvsD0ecy+krJLnLpo/JuVnVF7zUzUBF8bvs6XxpJY0QB+OCx0dG40uU6iplUen
RWe/IsoppwlH0z3zRzlUPIQgHEo7icW6mDHZJKkMFdrC0J+S6CgX5R9UN+slCko7cKr62jvV24Q2
D7MRqLHQfRPrf+RB+oSHZ03foJL3r/8PiWiCNCotB+1tVohJwyZr3IAxE3yV7qKndzOnT8VXidWE
wxmkeACiUwfLraxoH/IaX5bZtd8Jwwf3pfOvp8gQ3HLm4fJA6eprhMI9Gv4J+6gy1/QHYqKYcCBS
wSSn07lbcpvtA+NS5Ll+X3tIX73dqOJsF7awecmtR5ZWgBsKJwwB3UWYIdHicZM+24EufvHRu1/Q
HLE57dqaYD09/0PxORKJRhan3OEqKpV2BEJ2X4mEsmnIjKdM/62zFKawqaiDJdpJqV0qmT63d5k2
qRpRDDS3irSeKOJnluBP0HbtgY5A8/xBAR0a0/hPkGjsR2aMc+cTjmx0o0uKeNirlDyugh7Avrka
uO6UlyMSw2X7Qh84ZXMJBQWI2EarMmMh44rBJwMPqX+W5iYMTYO/nh+H+EfCmuE9ab4fh3LqNGGH
9LZynMGMJhdOSsO4kmGYqpxSExkrvsF1Qkre15m6zkZmFOr8MxvZjiDrQ48zfbch/6B8HAQRgnoY
JRkyeb+8OJRhUvDt8WZKchOGnJ0abBoBdCXSBVtCcNQllTUkrj/hnFYUK1Jx9M8A2FpxZAFf1g49
BAfyQvnWfnA/TeSFRLOZ6KxaqMNJYfbwFJZVF8Vi2DjzpgKmRuZG0ONJdkEC1rKfin7xsnk86ulA
7siupgkeLT9+ZvpCU0jJBHeBDpY1UGyiQ1N7k9KmvfQCoOJwotTTrZz0XT9qtzSGmeCBp8phk9ms
O6ykEWyPgkoMecl/OtMIIC5izr4yIWAToix3yUILSvEQ8TdNnwoUUULeQ/4tTFADzEo9Ao2DBqDa
PWk2WLRUxC2tOple1pQ0wapfnLeXnqFh1+m/1Nkzes3Sx+epG9sTT+0LpjU8omqs4pl1jU/upEPN
OjLvTjQvIUe/3642nATYAtEx+pamOymTV3x2ekVRaLNVkYyDHQ46ETsSi4ruEqGiEi4ow9yab2X0
koUPTbE9xDHm77co8xPx6BP631nVcyfJztuO3TVS8EZAPYaFYXHFS8n320ZQrHjYOCjFxICRWgIi
Rr7syHd800myUD8qOG/s6AeyxsglgW38PteM6hfL+eNgCGC+gVdDo3AkBwF7qdyN4aBHy8JicBfE
Q1sYAtoZRCA4shVleP5EPbOuVZiFwCAWMI5MW5IpPAccEK6+pfbpXh5TU14PZGSnNL/6je+Iif3s
ue7fFxBIHT9qLY79V60sDFSnu2/R2Xsg88Q57rpVwJrwKv9DzO1RgQHFaqKU5CBMhIXCfgZfqML/
qsym0j8x0F93CcifRrqG/z238cmQyXHT9St1aFdj7TUAQ2yMK7NEJmqpvLR8mPaPNP38SiZ4OALv
GKMadt5h0DQRM+f6d+RThx3LOQcc62vf0KjxbIrc/E7/Ngxt2lqC58ROntNumkXYBtv/ewmCM5j8
c8Wn84uuHjtIgCbY60zOkd9cvLM/GAFG+IbIAtbQP8j2duVuX6ju8kjZakM6GYq9hHbC1qCvTFX3
U8GAGv5peQkvgTpcPZvl/BFnJTTPtjOfWuT6bAAnfn1WA+YqW2/7Tu7qLnW00W4Tl2aotewdZxPM
auBICO7sz5tZMxtdiSthx76zdqZHGJw2FUWVf9ooHIjXJUzUBnr+aGQeEMImgm62b4xEOi/lOwt4
97Xpsou5c2kmMC+9diD7ejD+AagKMLdGjpgbmERZun8qNaJdKxjOjyWoQmqC7RfzLPnHaXy4Om9A
3vsjK0KDOmhaf9GYUT19GdUu7G+h/E3cTLJEbvemFv64jvyx12TaKnZu1V+g7p78mdeKw4yZYnM5
TzxRXu//YM6EZSwGAbjs4OlCU/9df6z+X+ORakszs3hAPikQALtOjn0xbEqPo/nGR2xBYEhMjX4R
63dyqBFRwvX18RGtW0ep/lhCi/vGK1F08VhkENGBVv6UUd53QF80yNAlxR2gY9b/D0YVTN6fyvvH
/MA0wiXu4HKcBy6gZc6Z5QvPn7TTQNmJI8w8n7mWtWeMod2QVqbWK1KGwf9xC2upuvlv/orImKwM
QBOmt7yTs70TqlepnWs8H/gxoZST3IQmbdgzd73IPtXAiKMpAC7LGHFaS0h9DbMJ4Q9pnDABv/dE
o6gjNgY3JXEju0noukCdli3pvs/TGZ1KaxyXW1o4Zi8glQTboDilv59YligKTwUDCpbOmfhfeN8d
QUcobTQqjgN49DmQisyxqBqzQUiBZiw6hdOXqdwrbC8WDPasGaVh9d/13d7sTou73v3sdTKR1ULc
XVazseZTLDH514lT7oXZzEN6vbQd65h/Y0deXrvXgvAvPtjTfbV9N/KoELt+nlrlYwG1aKjR8QSR
s/OCVRxGomYYVxJ4hU6A1d/Pi7f7p0lhmr9cXFKP0xMF5bDbTRvt9JoEqrCozfEgZ0NsjhX45IHA
Fvfpug8MiX9KK3jozaiZC2sES+bQ7QCuagOIgPOouKWB3+EWlvTBhR6L4wpK9+F/6OnZdsJ9FiAS
N66oWkd4d3U8SSpMDSzMIheD00hAc2FRQo10KzanJupmLWacmWcPtU+a9cUnBcKzzD4KHBm4Dvvh
rEwBfQ+ELGjkVe4e90Gr3ie+gqXYo4ioGDYH08VkkKw9RSIirz1v7TJ1Lzo3yVclA+oEGQ3vaPv3
5A/M9LR9C7WAag+XqpxT4FPmwX+3WMz12dCIHohFlMgsCvTokswXcMz7aiv1vVoqo9a8qH24Ifk/
aMDO+FC8Dg45juMvGwskN7QoE5/Sn8eKd+lcIFuZhtKnmNp3uWDpne8w1pAhfFR7iOU9Lg64qKe2
BJs6plR0t65LCOK1mVo06m8+BB/R1y1R9R5xgw3YLyWh59vmv1tuS3uDEjx7LbTuqCRp9C8yro0r
t4vowvZBvnCyZqEv94gVidIS3ll3QduYA/f3IlfmqONa9dzBoyvW8/9HVRgXLpW0EZumekBwvL+X
FXG6qE+w+u+ZQdeTufmnPkLZkKpLZ7O+22u5RjxOUT2LQWKjNFB55bAiD/PZXYEx2pZDivd6QPqa
3eBz8H6rwiarz1V7mX+1XhsUJ5O0l3xlupT2jbP/ehVJlps1cX4vZNXUEUO6VET33p/0T12IeWzc
pKpz501j/5M44n3cUN8RR3Jl9OVE3IXWFdK5ElyIuuOj/n9rCJeB7oyiEFHkYErPZQUBGy7md6/5
QX8l+X+gApyXxAf27PUN+uFrQTKk7TBvI0T93GQKal7YVlrH9b6NOl4QFG5Eyy98ogUnQbramKtp
Oy9xnPCdVeEUgJgCJe0IKl31LDsdEaZuLlmL8gAVvKOzKf9mzFxD5RBm2IngFkYlwzKAufryuMqW
h0ELxT9m9PUCJYZ2/b9VF9L/kRKqlRSrYxG3nN0S+LMkT/bHqTChsgwY5QT5mAMw8q5M71S2jFe5
3Tq0mOZGrqPda768DfgpMnY9QLn2iu3n/4/2q7G5K5p0P8jjh595EaUuZ0ueRG7mqws8EN0zS8AC
hRJ2kwMeC4V+zcyuFKu3hHQty0oFl+9XJIQP5kxMpBnKeQoXFP4eow3Cy9gncvRfNecd9Q4vycK8
w4jnNbAxRXSI6HYVD4JeuRwPbgw7ZQ9qz3BMiDFt4GphF80IkGd53EweRxlhsNccFQFeDPc4gr6/
1hSQa/774XxGXJ29gnOhpyNetK6LReP+qlh2t3jYMBMxtP6JSikU7BKWlqFmggjLwS4fdXWUM6t2
UTV8l4C4CL5jw/bmXG++2yZY85DwUW649jrsQu7K0m13l9xFw3oMKFmDGF0PPxR2xbqE6ThMPEFo
L4/E4WumidomHGOno9nJzZH7QEICbvahyaRszSBXpiAE8HVUCb8n1QkwhryfYLakdzlxa+WcK4/7
2AI2yOYu054zK+XhudyBkhVcuP5HSQCGpb5rE7YWxhseoZJvUiGxFOc6k1gB48ZZtjFRzRr3wJN2
RqijnYWLWQmulwuuDB6pCkrlNHvbJ90cRtAzRhvsRU9icdZVAS99Skuvsve5ciDBqbK1zDjqJJV2
77wtfyNW14Uo4MUYd+QUG5LioUtj70uwSt83lcLEXh3/1ai0l+RHFs5aTZwmSbIDuf92FRpOUzcF
BJYETPAbbNn7YkZYZl4r2mzJO/W2j9gB6ArOFm4U+rFtpWGXqNl+3X5FLNPDYg5KJtocCh5l21Us
U8Vxrh6Ckpge3/4SieTafY2xjrBNGbUzZd8vrv7+rq9zRPis7gMy27dMI6hF+j9tkq+3St7tdIXI
72DMv4hgAht9C3eEPtquMrk1amNsy04jnQYoUJC9ik0nkqd+Oc4ro8uJ3E+7P19xlAlmYUwWk9Cl
k1ScJ61D0GgBoCfIAsmgS7dLtBFNyem2g8QzDVvmMhSu2/zsfp8GmvxIj/73DnDlxunMiYNChscM
2oJYd3xZo5JcTaEOu2s+R7D5hMTfVgrPWcju8pnaqW/sH7/QUMdfPag3QhOwUeHZBc+CHbeAiejA
qHAFPs3F3ld3Q33VvGRhBKiGJEjgDelE96ner/7tUhLu6wq5hSnpLSZiFhjPCqHBLlmurXxi3WSw
d1jUPr+aVKNwHEGld6fFHr9W/GBGOkU12jjAQDKXPIu7UNB7/ippxjtgBhUWvUvqfbP3vK6yKLxS
9ntezoV1MA5Y1WYyqgB0Lo95mxFPiRc9R2Qt68Y/8CHZRwOY3GYHFStKVIu5bQOZgZGLIGGtoElV
yMWvxgXdtOMucZX54QuH8nPyD5IcVJGBxiTcNn517EtB2A6x7Dtb3IyERfbFvAlDtQaT57kddAiT
j1JXWc2weeyV/kOshONPRVQBS9CaZ9NWUXfzvoEo0aGixQInDuXy/sHyURjhIpKozXFf7Y4Ginqf
7MJEPFos1UofWSZo61rWQVfnN2MZv+1a8yG7pvn+ZvVIFIHi/CD8fDndzxVNrkbQj/QcTFp5vrLI
8wnRfW0BmIHuTp5OkFgp4TESk8p8ikRqyQ/MczvG5Anu6SiU88MpDpqpYMMutD9AozTxHv0ynSIh
Ts9/yzMM+CyS31BTgW7rdw8AJCU/QDGL4uElnboCFXcYu3ZWL0XkB2hv7LMzYiuPL1chVKNqK+5N
CJKLQ7NiOLye/zOthJB0he9Uuclo1CpM5yIRjK7fvpOo8L2bYmPz56FsYnDZcDf6dkYR0YpTKKLf
3SIvRpBsUDHvBeZ9RCcpTAzjq15RLWEI11lgsDhMCCGEG0+yDUM6/fqe5BQQ6K3lb+pQWVEhgWF9
cQvoAemCoKipYB0DVNWtldMPrKZabYZ4Hf9oOoo3WaDrTlg/xrca+zPrOcFsa7AVuio4hyjaAShU
NVFjtXF2qJj/qRTQo3Bz1BH9ACWB0gJp5ofJeiXJIIXgW6U3f0Oo/A9hyEvjD8OovjpiHMLXTO8j
M9Eul4H5d57sNPQtiq4DdMlEQ0M2yqJg4NN/WzYcpBabkz1Bw+tst8Q6Xoe6ajpOED8NONUywNN/
ZSNH2p1VNyEyaUCaDUI/n8s/HY/EjpiRsPbZBnY5wJzR6nwQfCVsHIYW1UewGXgRc81/lRjev52l
HqqzGqMksq5SDXCJOEMIpWax/Dm4ighPWSPylG34xgVdYUpZH0hHDKXL8XqDRMet03sQjvyxkzxl
5El8T1+/YEhnnLYFI54sGvx5gMNUSSksbEaZbXJp+QaTdTUEQpUgPceLewM5ogpojEO9RoFV6HgJ
5b4Q01xPgdR5/X9To8fjpaumQ1kx6yJYqZUJTrG4KKc1Mk9EXkz0Zp2pyGTVzKTh4a93rc7mzhbl
aRICbKmnOnPvbQQBZQJ3984HEX9kYsY+fA5rg3FOBv06xuc+H39uInejf92L0ay8doE5SkFUEPpP
782r7tGUrdwas2GPYgdRC6ROXT9ldL6iyBQ6mQv7F+bKM7u3G0jhFZdtA4eTheg15jcSQSELyFp6
6rPOJ5QNsX1Mr0bdq9ObOQjE0XOcGfkfqbDfh0JgdbfLSe+TjqfkI6r0rjsOfri9krzJh+FY6Edt
fz+7zDl6vVHieKxgKhqJrAUOyNLUC9Pn4fggpAVa0q5a595ldkfWLosp3hTVxzTQ1fsVujibTzjM
Bj2Z2FUQPP5uVqjZrJLf6UD9m2mi9DkuWLF08LrH95ClOijqlY0XcqzsZNG7RQqSEYEge1paPj4D
94FGRngv/NtDx1fQO+R7WbTL/DKjVLzMZM3kTIwrUvLWUUmUJIw5kprDU+Beq0utfU37bSehyS/4
6mvWFT4sHFveD2NmmdI3l53qnzHpHNM7NbDl7w55RPjd/Nxi4FTdm6GGH7XLxUUeKxo0+Z2n3qtg
wId++3A6GlSzonDcNm8oNFhlW4hpxYN5bGfB+4iDmyNCsstRMId0aAd40DiJNFwugkj3F1Q+G9v4
XJhWmd5cW4gerYD9cljKoQteZm8uf0UDfNnKNHwpqU0DBReeesJ0halWsQIeNT1JmVyQQAKS/Ebh
B/NasRT2KovEGOP2qHssS11PqtFZwEUxSjgs0BeBwb2PNcJOAPnwruLO5x7vTJr1/4UD0icX1pk/
IQkzzb3PY3u4Dly2f/INNa9PSXWRIRY+rusciK65mVIRfqUEwVbBWBLeSCG/xVURYSEBHW1zq4Df
L3bzqiWpRlEUtA7RV7DvVN5aIu41CrLhfbN9zKKdz50cZocshOLWxBjNBIUnkeddXhYqODy6iDeU
kjkg5eHBL1ZuD4RTzpx4n9e4vVlWkClKmPBtzGh5bQbEsTldEizqlIUhITHbI0qrZXCCVDeblcvB
aQsLzY9ECJG8yZY1K8g28ENa1ah1yqWkq5MrtoQunrk8sjgYpCJJTBv3FqSqCET7TSwQWNLMwPsn
Mxsv/ycY9NxMs2+n+7TNiCcHKyn+YWAg6wocsUTiGeIA0DhQyi3AFTvxqWSP4J/QXOwfd8pGCcai
PC05hmhByx6uElXR/5UdVIGBtkJ20IyYH+Z2jaNrltVG3vzLinkpKkaNauZINHn/VRdJ0/Wu8+bb
V39UBmZslixe3hvTcszOcXiSmSKvaP1f6HFFN7jF+1anHZO01i1K2E4dxkhJKVxFGNoL8f2BUvur
z1baon7Ajxphew/8px5B5owsAy3gzSUn10v5P6TcuDRyhL1otPfSIjsQxWzxkDuUyPQC3Bo2OrXT
YZKd5Vb/hKRPIOWgtzkPGv052CewCNttqoVCmKS6W12wvocXL7oDxpx2dbImN1GlE5oF2/2LhfRK
Eopw2Jr+y4iCn8QoOxI3T95INWT/jiIh7M72+u5YXRg2u3CUPChwOJnYhOWsHA/tX0ByMkjjZdzr
3wT5YWNgvOM+D+HC7hBhUcfPXOs8vWEFzZkE4B08/OkfQdHe7v0yawuzW2lnaco6zjHDRaf2ISqC
Un6W3Qv8xK8Zf77rkuKoNlsqjf1nmFvNCV6oD/X/ZYlY3Xl0dqK0wFopaaqQPm/L4Zgi9UGoNfhd
4VWGbNSFdyXEDftRGPtNbe2kkjlT1ufUJkWAGe/x1kmiWUF0+FoM0qjezDMh3uaKrC1BL2KN3sgE
7iOkICCpRWFL0hCZ+overemC57ZFCz5F2smyB3jpB9Dp0wAsGrEUoYdeR6Tlt6zRNqK503fXr6pa
Jwhp13w5jX9soYBgzhifmmNxa7RMjBBZeoBLez8VsZ/5yPuBjCfSa3upmImcLrlrax33xPkX4qYB
2gOKuVCKIkUs1U10FHTH/juEyQ7xZit/CKQua/XJGjVNm4RZot89VR3kf1YmvUET8uLVrpQVHQRn
YuKRMHAu5WLS39dj465EcZzG4x/q/kUAC+/s9MDBzkfRZ8+hCsNnz12KZkAxx8Bc3wX0PPCPWYI5
5jPdIhHQ8CtIEk5ieIUBTWZ6wX1LR9xi+6YwHASjJ9uFSEPk5AEjhPDDwNMWMQmwoBjLggpOaKDq
9PYitC8da7jM9QhAkk5AwuC3F3O4lKN0IrhqAOs/anQQ0ZFxt/m7xu/9b+xh9FI6vj7uQ9gzCnTR
bEU92PrDqMe1VcfSlaXqt2RqSRwq4pS7Q4dI2ItwXE1v3tST8ZXkkLi3207F0s+e18hLImBWqXfd
o6BW95ZEXEwLWU3sq42y6wSOXAA/9xjHC5pxWEcx6piu0x/37rS0HGuOVUytyJ7EtAL1iOI+ldlo
sTF0rfoYdC7op6Mx1sc8Ul9so9oTADmdnYw4MhE1P+4L9cG7EHmOLK7C4lRrCKz9chP2xiusoqTs
r8iYJSaF1NjrXzOoq2TkUrQE8yuItEahDNbZym/oNFKgNiHflTscu3wQFjmicXGlHzw1mYliSOXh
sD72igdkW8BVH8E7oFVC4NgLtf0jg6v3K23xgolHTRH75vg8cNE+fCLeVU4wtb3gmmtXv5KdgJKS
FawmYlaJQIPJZ++nyZeN/KiMoevziFPJ1ubZInBXg3V1vCDssBowy6cb4RIOMoyqtZWOsg1cvvbH
B4RkjTmIPSP6J67XI9FPmsvJHY5DKAbMQVhhsILQ0XpKaU1+ld2nXTqMlope7Pev5m6ev79rYrrb
fAzwaJVq+0cbOdA3qUNp6KX17nRyMs01qKAdUti2J77erGx5GMB1MmXc0WNgAGwUcDHc+hm/i85e
KJ/AWnPFmIL6WeZIqbDwg3XZQ5D7h3duPy4+PfQRnVvXsJFEQwfo73IaXbSDGtT/0Lj4TRjFyGwN
sYIKsEvtCnq3jjQRwFEWvhxjuflH0Xgx9GKcMDm0GnQswDVw3EbS7+68bjLKBMSVdEvzbaPvOxyr
8GibaDd97DYXFsOxwNFj/C0cxrVa5QKEX4bA6kPAsFwBq6fsZ/iGoPec5488//nU3dsvqFMjoAxg
6ixoRRxuwO6DGNZjdE+Sqk2EMCEy5vvHOJ8V2UiGWGRnrc+IzuTBFjT+Yx/NtdTWn75VUF3XMfap
ZrtGSCH28ivVSAtcGU3Xkq5sY6vzlKv8aaip7X98BqoLH1ooOkZRrgtG3QbHEj42YeWuzV9gJanY
19csFurMn7YXnWaTcQHkgDJNyWl2Jgwfsofb/na8RcHzuDs6URNSEsem+MVitC39XxkZQChATot2
3Q86vKbIv3ELepRrO3cTkv1Yx/Y9PJYRZV67Jg8QWt/utCvEIIV6ELvl6DBOzcMpbNmoDCEIryiz
1TdStKZHeQTo1KHak/FGHyykHjX/ec4AC5KfC8UA5855sy85R+0vxbuvtGiddzETAm4Dbk1SPRTn
gEwJoUs1rSkk4B23hsiyeQykM6NpyT64M88C/setSwH1nTWtxEg4TeULKGg9sX0uIwQ9qrB1ho9K
49rtpZ/NiB5CDXG/pYhxLRgeiCCNhDItKuejl3bzW/3/xEGI6PlLK12YL/MknXxfLzVxc53WaJyw
0+bHGF31AAoaaV6mvxhxG2AZC4DXk5YTcAl4pVMNxOAWrN11o7l3tYaXZgexyRq8fWAyGyZHB/G2
xtlqC4NKeLGOJkwPS4B/K5JPIjVM6b9RP96PTsIrnQpZMbPeTdGJDll/6jK6N0/V+Lb1mJZRMpI1
v60KinXAPYhmRdWYN/rqM/4xtVUVUpbuKJIdUrL+RTj2EjP+Ok3Woq7HXhPN08W9mDcS57FzrcOM
xqyUGhLi1ZDGYl3dyhECQ1nnsFrArZkwVupmCryuTvxbU92bTYrYvZEtcfD/t5ekor1JQx9e8/st
6ptcRYry6KhbJmNzDqMCu4ZsL4tRbmvKHPIdocKOOLIphe8GhhoC7wui5mPS5Mg9qjZStHcj9MqN
WV0MMNMHNv8y4KtwSU8zPtI3TOcO4dY0D39zVD9JZ+rGO9mA5Bp8CgkWOtdsHU1ZBQyZWYl4wOI0
gJI9253eQsKukEgW5RpBx4yZFju6ax2UrFHi6IIgZjgkpVH7BVFX7ikRV5DdNylVVghIzQucS9X1
RiDx+saAmCU5V1ayGyAoVtG3A+cnJNaI8QS6vujnUw6A+75Ml8iNjDRGM+j/xrbKcVc8rAsFl/Ow
WvLJZKS3kjBVECRqdPIBLTQnO2Flsm68vKAGkos7WKUkiOtsn+44DLw1rKSGgvK6/9GaAduTirCr
DyE6A+oXV3qieYY1H4SjyejQTz7yIrZ5/QI4PNHPzXw5fHmBKVN+wnoNNZpf0BAypoECZ/dLttVW
ThxzHkEDAY6JTdUZHkxDgNIERJNEkBk7SPgyIBz7fLajAVIG+qIQKZqJUtPUyF7c7hBQ242Ky87Y
7gvTINi2PN6q2oCovX9/wLvqjCMQY81iyZ4yRNYnyRG6DeZxbJLJMrbADwuAChkLG0EawDwb3t9O
mnNecuQ4eXujWVKqeqvrwsV35TNP8yMoeElu3u9LT6A6Hxd3sURsGu3bET+ZIUlGlVEu0QgFH4lX
9/2Ul9GHVnqNtdkY3OAcE0ZZYQxGhpKBzLg9M+vDUPER/EGwNu9RwKUhmfldC72ME1lk9Q28Y3RM
Mxg/anG8NZJXjduf4QoVI/94q5l1SLoRnPwNguG7MXNTW/SNHu5A1/v6FksLZz41R8GeN/6x4m+n
GsoZsEgu9f4Zf5yEIOSlzg29TQutmmKNUBF6GpL8la0091tAGUOZTA+4XJNhXQXlybJu7m3+Bx3a
g8AwXOnGFg/heOxvo+lPLzfROl2q4CToieUa2+Ry9bYssK7HWqQvBMEqAKPEtXco/qMbERMo3cVN
5EvkK7p1YHr8F6eJ30t36xFZHJEmcFZflXgCihg1qnRC8EePpyWsJFMr3D4rFGSNOq5GpQrfosYw
0JsJ614ljprjmA27pgGTa9T8rfPnziGYHDyetmeJNkJ0UlD84cCDSRPBVxuFNBIewZWmEETSw5L3
dgcSBKFIoF6h9xK376CgzPQOFaM72jZ0VIZfHugPGRCr9cXjWwAcewwvpXGuW2Y0kQna+O41nBvU
hNJhmVXHViQITBERDegCdtU0+EcC48T5g3CmiN/TbGlXVvOII1+MKQq5WIucjSe+twmHYUZ4vdHK
ZQfuKN+/Db9lJKLyG7U7gaflCQVBAJ+YIrz863PyHIDbvJl8xW5XOdl5Jl5JO/46YFrlXjsjuZd/
/KSNk/P6aHheeoZH4GHaOBoJ//Ywcq1DfH0p0HhjFTTs/VUcw5fvGC7kLy3WLjNpvG+sIPjZ0WiO
FiRt+o8g0jDzabvj4rHmZRPs1DSHlA7f6Z/ItbW8VEE/32Cuh597cXdNkCfSL/9+ezw9YqzwtuGo
0qNMUcbKjD1KU39MQid8McCxH1EqaEaTAne8oJTQVoZKiYmGl6xeGtAmuljHX0bIZfGGPf3mTY6D
gXa+LomASBGhkQqj3dG2EAnL5WhiL9zhe7AvPr7lYsxcqu6+6pgIwhGtm39yLbegC1AZnr7yKl8V
cszCY0mTtNEtDe9PAl+oilNqG5Vxb3ssSkgaTLwT5o7DBYZ95CK17pyOhzVMqkhdIL53I6Wcbz19
wiuolgOQHqrkQRBPBderLvfCX2fj7m9kfgsZWxXVvJBZj0+Y9fc+JnJsT264P/xJP+osB5t4x+Bf
6jKNnfi42CGs1sbngUjR1HLj69Mbvm7OeXRd2EFOWNp2+2YQXjEFIJ1jFHmV10GcBl6kcz06piQe
lFtNRVsf/7iSpxxAKiLH3S/1sWI50eUzEoAxxLIwLzt4mUZwdhg53IkWqXBDdCyX/7oLk5Nu9Icu
vT+YuVTIWPwDE+vdLnjLKwaoLLNsvt8+j1/uxr7KuPC9e31BsZWTtZMJAUpromj3nY9HqrsKXlr1
KmYQOcqB2qNSkS79dTVrI6HugiKmvJo64YyE3KqpSYxOnhYSI/kKPxUh+sdWYCtHnD2rHvTmHizB
VRi4h+/l4izIVOpE/Tqbt7nfi8SO3j/VWNHBqfXTwE4z3LbtV9X6n4eUfOaFurvzRkvxHbNLx9A9
T96l6DxEY5nbbeKmM6Api3aBqIkF1fNMNiTzv6rJPotQNxBYzo90i1KUdhhqfpOJv86LLszvA5MS
47xdyYF6rcUNdcRWPghgQWQvfnyW0fAzRMJCVhyAdunA1Bum2Ofg7/9/OF0mFCrEmiSNbVgePHNo
VCy8DQbDusZMOoZEPhpUaVKBwKXQRGwxoQ1sCV5GQRlX0p8qp5m6eXCMiivmQkcsT9mcDJG4K/T0
nuAywsZTYeHaKaOtAFQxA+V5kNI2eId6OmQvfdubHPFQMft/9LFcFJhceKQRs3CPVrDdmWeudhim
3bccdTMp6BRjoZ+jkbunLCmJU2OerflhFtWkYz8TuoEO+w6QVQknmCfe5qGYJc/7XUWe4JNPXWTQ
2LDEjrUCdv0M01Chg6SLnbDJ0SnGDgTJncF33U29f1wGpaQlMsbbKDIVF1rZIg3ULfpWvXwwDQV3
xOjqOct5zWBlY4+4klkr91rIeOEDTAP+yj+0WNd3FYl41Zi+etVuNgDmR/3fTODKWKG87rjagG7c
Kfrq/MaZIFQl2mWlybCaCZ8z5AQXqr/gj3K8V8AWU9CU2ceoHerDYQ9MDOXIfwmJMionODxohbvT
LpfEss1pTnwi3gxYfHQNX+X/KaMkm7Kl2OpAT/rCK4YTwBWcVmdLWq4RaG+0IHRv0fJdEAO984OK
Y2IcxOR7FcJFBBl1tVEIR3hGlSuAvXaO+K3jpvDGUOY9lBfyLcR+h1dxjbRnKbjvdOxXCw+HKJw2
Sm2TAYigkyBjZr8g+9Eptq++IyDg9ir32lf/9Fbc28aVBZhIdZhwu6iMVBWHvUIBZirmOfD5KyPp
aK5yH+NEoIE018NURCOJwEWAtYh5Dk4UDJACl9tz6VxXFSam71Z/d4a/gnaSgB7jWrkBWL34sWdp
Zb/PU7EfW1IAqXD/vCXe8qtRZ8jlxS4oufw7+XW0GEGE7i2NXmRFQllaCT5FNfL9tdkkFphcDCti
gH7YM1asLhNVy71sGm/lPD9XiaZLPRM1n4dSHpdYNMplBQB7rs7a5UPj5V6joFNLt+kmLlRawPct
ry1hhwVWkj8oRbIjsRwbp0sykOgwzPKwo+r2sxBAYZcjiLUyLovw6Lkf9QYQ5eRui/dyC9z9iVaQ
Ag+ISYatjd6ah3i0t+1zTH/1pInJWK7NI6TDP8GFX0zL8J4HufABL7GKzfXfqdBYIPld1oKxOazu
+sOzB8OLPmMw0LBtN8WAZPh2Fe5Pf+BQoQhZaHMbD0fx9TjV35Qm+3Fwz/LOTH54pwgWitq62UFQ
gfY0vncmazScqQwt6S5OVE/j7Se+kXuil24mqiPRaE5DUXrUiX0C4R5s2Se1ElBTnA1YNn/q1bdy
mGwqlijQE1tkX4nZUsHRtxPcmewlLJgj1I5dQBWP/4gwhHIC16oNl0mhxdCrMGRnawI7rU9m+Xb7
PpoSopYnmoOOy3VlpZa/8UHtFoVF5CipdyfggF1Z0ijaSyxLvg8hM5PoX7WcF9wh4nf8DTKRBNn8
GHAfKt+fdVXUGYDsZsnq75Kohkp+4agmR7+fOC5+Fb2VvydVdkdJtz1A2O5y8tPFqN3nQaZxJTup
GiFOe6/XAoSaulK0iOEvxIr2sEuK21899dNH618YIm46cQ7wDvIbEivV0L7azkl//CYUDHuoTha2
4/obKP/oyUDQOTPGr58Gga+muxGbtVpl8kHxo2zcZZKwiM4GHqgncwEbIS9zfOUvfulC+cpbnQe+
2BftsGKYf3XG1KbBrblgsVWtLauTTWu7O2SslXAXT0QNPeeWR+Qq25bXCRHIqyXz6YJlbdse63z5
LYaxMm+zCzDyMigo5CZ6QaQHIja9Rc2ZIW7h65O9p6mvj4OgXPCe2UK48NwY66t0SKOPg/kNrVVa
A4ihY+3J9fWQqknfqPU5+wm2avSdzJXrrxSdSlaJcTZqJok3CrfgtNtge7izyVbU0ZZZqxi2nHSV
pKbjjxtKmpRyEe8Ls7+jxQOXUA3+1qNBf7zjqk7vZ6fw4po/CttBRzBhwlsw3/VOiqrC2qbhvJyO
0wp5Fg9HJiu7w9rvU+TeaOhglCr/QzZ1zDJXimfuKI8acFnWAg5CbxIV8WRYjy2NbuW7Qw6WIioF
/NfdTDt6q4p8aJzWLjC0C+8mUf74IPgOAseQZt+fmFQSFG36u7Orpz5BrHHCFZWHNxE4Hdx7RCd6
tsjnILSuzLQ442fdNQeLVUxfuvLqdJhYQ01jmmI38m33wqiZrI/U61B9bcpaA4amQdumYTIn+nL5
4pxsLxBsruwZmlwd6iTRR9WK/JoIbSJRXaHkIAuQXEMCNOEBqJnWSIp6fe22+wnCNE7H24fGRuUX
yPm6MC/Q8MkXO2KNLHuyIWfHjYH2fZDdp7z4o3xk4wIPhuzB1ezpxWKmfoklKtRKaP23btdXc5HU
yilvSKdaqtbRL4rrCtkRHedgkS8KfBMSqaMNz0KjidRxx2a1frZb7glNYhnmOWKi3ajbEX2xiUzv
WkCkfsXNbazwwIMYJji9TIK/NqmLGj+KcCx81SJL9XXSqqqxGFyYAVBEScIjre5XqbnuvGXwO+yD
/3k5cHwp1tk3rSLMCBRJ2evp14nEXfGwvWhVXOyETwYZkhxPX7nzNRLAiKzEFlxvr6WXfQ0NwAMx
xn2hd/rxVvnMgyxsGtF1SiOQEIoStSwKqeaFkTwwd5bPvTDy0x496+4lPet3Mqhc3ZrUrZQBMSLd
fMNoQ36/YosZKTboSRFoKPrFmHKWpqj4TGRC36PAVa/9VNZlBshQx9D2jdtF8Y/6HT2bZzr+QGmi
V2rWc3mLesZmM2fPeRvI/o3e9X3OCTgX232VhaTzlMiynekYsUX5BE+Cc7PAqn524/cqlKI38RRi
oOCeUwtBTxwP8b1ybrw03eX26AwUEEozrM7SkmwvI4RCzI4D6AJkmscxtEQ/fr5V1bbYAEgEN9IU
DI1Q47HzKzSSlO/YGRXcmU5r1IBHo4wMSoS4sObIubvhmlYsqQU886N2YhGdlBDY+O11wgF81VXg
pea/rCCuk7FDH3RLfkFEaLmm+d5U/DJFuFNl4ILyHS3HeIyAH7GNS6U1g3XkicvBFe4s4YewQiqr
CFxX4wqwRnuYl5ln8e9s/uFpK80Qd+LSkDxUNP0TSxPMkeSY+vdKvQgXbfD5/S0u6LZ6fOr9oLG0
W8lVzvtFKTlTrJELdAmRYtqVF4KKfakHpzBQprIJSg6ArOBujTY0fsXdl/4kOAkuNekoRAlmUbJw
RDYhVW4wsvTFVg9ngXwHyKRLDAuxq1OIF7QojW863qtQff6ys/UG+YbM/sw5ZY4sNP0DmftLnzGp
9XyHqi2qHZ2O+J6wcx0mNVq1FrPGqfNwJMdlQL+l9zWSzt3OvSy+kobZ53bNR9na1JzI017z2GtF
6R27pJ4DEKUVbeEaf3oOmnQCgRkY1XvIUV7vFIAfBv1mhv/bGsyoCN3coPXrKGl2sAnJiFf7EHXJ
pyRgvg2Zx/nRAFMtIVkBXK+nfXoPRhpTJWhscswPR4n1qLWSzBMSJ/gWjDBczebSqMDr7WR1LTD0
dR/W2re9u8/OwaDrHr8FpJeZ6X0eEzNedxm4hzuoCpXcbeZEPCsZX5H6wynKypl1RmG0sv4vxokX
4U3ydTzZQEC0QgTy+FkXTCSXIZCC4WJeu5PeDkGQ1v3BaEWnYW4TMO4Il6dv01oiiNruV5n9TBsb
tYI1jrNeORuEL4xZ6HpFvbbKFVLgqvF2c2cKEXhrzmLlxiXbCJL6n7rM2EBjPZx4KheFeq7H1aaY
whMiwXDaOmrG6Ik/brisc5HyK6l15irW8OXjtzB3jrs77lrTdIrE6bvwxPKQyl9OaWEwnb6WTuko
5AFRWIBsOvR2RSi0yQNbsbK1ZrIKvfNSwZb6lTCgzqm/qQdArg3oeMf+YuJNbIMU7lz77SfOTYQZ
ppjeR0K9lfOTAMO8Qler1CXZDqkxxTvrKsVkTuiIuloC3WKjAZM4m8nAzDc3xQZ9YscYkocCbQbv
z96gvef18nHDZ09IMnmLsbGcqOVuile8OQ3pDyMpayttq2Wp7rWSLgjdMEML9LYgLXRlttD5e/bX
8HlfkpTpHOGUWFVKdstX+znflYbZ/swtGbBQxt9gEMnzoaF0fSMyYr1JiZTtapc3vOslrx5Bx2/s
rcVXmzzGZWNTRiKMea2p85m+naGUb8e1/vgreUZnk9X9DnlCW4EGmtmTglcUCHaEDbwfq+PajKJ8
8hfXW2jb45Ddyrzcn5d58e+QcriAxgh1iWsMge0E7eSRofStBtTX7lO+VjYeBdZaT6tGJCkfdLdp
WDNrd5bpgkUpDZfPwiwl1a9Ua0yt5rZci+92vAaAHmyJtXX1Xo6RLs1rgigaGa5O1Qk4ErawyXzm
5lRHhMk5Vj5RI/ywFw8Tetuo5sJT5y1Xeatl+nHlAGTxw4KqVBpwjDR5IROEz1iK112D9dih9TID
7/RfG1EEe9QEsmmIV+QHiYXIRZfOsFMbo0ZlgwDFYOLHC2zj80wLD7OyBnHjcDnTQCZrqZIfhudM
JnoevIvny/HHF5OA7JranWz206v3GhF4Z+XqtU6lenoCnDKfA7DRxu+JEtgwqa+AgHFHbJYXPSSs
xnEwxLoKUou1tbWqJwV47cU9GdHrkfb6YUU8z5hg6ZpuR8C3f/k9dveMeOVYRz2DQbKXfvMZ6MiT
CnldZYjgk+CAwk+4/ActsPBzdKB4lN3U4JXhaze6GAsOgpaCSBi/O2hsvZqVV/jVkf4nDm3L4qqF
NSYkY7ISBSiBxxPcJwDSe3e6jnRO0i+O+gL4B4ZosSFpm4YuSDz7TkLgDloVT22UjVnS+HFy7P/l
/DaPt9Xr09TyFfEKXHxSR9uoA8j0PtTPzJ1hDYR6BauS7/BQiR8xI/UGMVslg8cyZEs7KpNFbOi/
cOuOiR60JKg+rZalcI/kEV49RQcQNpkzLroOY6AaE6wMa+TAG6T37Vt23tSVCGcW7GmjCmZ9VdQm
ME/Jt9caKLpo+vVtRpP5s6m2jnabRUt4VzWv01L6ZjEjgCnFQ3C7Okzm8RNEjGVqML/O5liLBpDn
hHImzbWGoDH0QISSBnB94efuPBEWmfQLqJxbzWTUKMsYRaNCZS/wudfFAUFIjkyg3+bEbZ/ZhUlR
ARFBMiGHLW6WHSSj8q6RGHLdSDHcWn83EvIILKhNRjWMcOZf9daG8HJDqcxuH14R0uhWu5+TLPUH
paWa/47cBEHLhxGZPQjE+2T3FQE44cAtItKfYcxu5faus87jx+EYSKQd0ix/F7fttXK7mNJF98eZ
R/mnU1xSr87iTunzJ7p1GHaOTyoCaQOROfmWRVcCd5QQa9/KZQAiK1QM5PtdXSgD1m56gAhif5x0
ALbdCE+OgWDAXQvIj0XkCnMdFiP9gbrwd4GVSooVSVx3Gp1wttOz9m9gttxV1VUMNZISwZ61B/CK
5Nk8xPYwt8UouWz6gbrw0IAsEtqRgqEgXz49vlRUkow17o5fWRL4GYKfMDBoVRiigyslxofZZm4s
lkyNzQTSBTgiZED0dx8LheOv4B1xKn01htd0U19g6c3vxEaUr0hLW+PRUFfdoFwx994HAQAokNHk
bb62JH0neb+w6O7TCTJt6fWh9cx2PN/ilF2EFzv66WwQMgGwosmxfjXysZOP67bLMJuMUodRS9Dc
6gSQjKOw5nfB0kghPAx7aJqy1wl48z/fQUb7Nz9Woy7EqLvwF4IwDsKGV/W5UI9cN08NbRMXP/rc
rm/42PBOl92Zhs9/WG2w8dEVe9W8lwKfPU/NKjIH5XLHmVHHij3Z+4YHxgHUhiOugM2RHUjeVzTW
4VQwswE/ohh3IRT1Cta1sMG87tatYgJgyIadtFlwxgYVPgjG1V36vyqq0BEECrYySP89VrNfd2iA
o6TO4ajANXaxgL1QtMW+wLkniRzvMOjttQmghP1kNa3XBzPWkzWaWn7arUnj/ry/FWJYmTdU95xE
z2pC4GsjyBZRcQuXHzeLevrK3VvUZvYsSgssGA2s3HlRBNKgbt9yghR5DPXmUGKiN3AqSRf0m5K1
soinl1AejDYT1i8GPiUKBFfK4YnB09HDbbvSOAeleom0R4UMpLxq1rEIJ5GZEn97nbr0dREmXQ6K
ZkQk3nDKFAu2cnBEpK6lrDjTpwNBEb3Zq5uOSVwdhtQzosoHd9dAaSmCQApR1OoVH2NI5h2e/D4r
oX+SCPnZ68gdOheG3Xl5bdA9YtrvK2/hGAOCModIEAL8hjdqLvDy9gTo+j1dP4mcAngmpXUL+QCs
8sNB/9XTdBpccMnLJUv7G7IEJZFM0oPRtse6XJ4PGYye3qyCmYw3kNj15yELf6Im+VXa/nIXrqla
LmVkS0iqp14fnpyVrOxdeZBgnjD//BRi2wNNuhxoAKPWBl5O5j/fSq+sxUVEE/AdnED9BhQRiN0u
J1MDuCAKQpGvfTeWRfY72Mrg4oUEzaAXEqzAhz6nUWuKKhzG5yriwynWruQXpYwPp6tskmCEeur8
sx7gaMn5QaspVnzzkCuJL928f+DjCWh8gk6eDqdr5XEPALevAMxyX4HlESSIioGuaHp+Iuxg/GRf
KvJ35j0mfHE2HVGzNqiW7fcV4/QpggmIIXyX87qPlf7GUy7JOpHLdXxKwzRO5rN2q6o+Z1NhvfmS
LbDP4PrUFFsGusfXrEi4Z6xt59M3Z21mXxm9pegfyvXeBKZVxPvUCP/Nhakt0EXVEbWtNjw8g5h1
G1W2LZkxqvL9wEJXsz9sgNFVdTgWGAVHlhjaozKIh2hpleEQucwd3oCNjhW2zXzN2ZhwqenGOQ50
CEhlG9kFWNwo0Xtp4n3qrsMu+CZZFj96N9+CCMm/H28M8Frq8xwgm94RcK9ayj7LVbNPAl+9dg9v
UdzOSA60Mkg3OswBFlrAwUrmN94bSnQkWCIZ++H4vuiVO672hk0aZ9D62VCUUZA9AB8A6StUEDps
E6mKY1lkFEu/CHxV3qG0a5k5z2ffmH9cJrgBn3dva/4A/rjIFkJlPA10b+4PbcqYHtCylfqikYWM
FeaSEkq5GtgnI2vVPW1TBaLMVmBaT7jK4ool2n2WLKUdX6zf8H24xgYUuJ+BbD+zBto+ipJGEhyj
6aA4Il8URwKkesK8TEfH6X9LIJLYEkZWJ2d5QHGybsTlCA4g8DuOLX0jJ/IgB//LOHgQM4TmY9i5
F+SY1z9XjxGEOXRsX0q2NSEUNI/U1z8A0vu5uDb9tJPlhaM2/i5N8u0qgzHvRqrN/MuxJsKpIPwk
6o/YeAJywMwO7CvWD8aQ1+I5CRx1zgADYyUEYgXNvG60n32t4PifLdkDDvGa1dTLrVe6rcnBcK7I
OJrxAfQyWyEOBQUg+HiRlEmR39JS4m0ixK5Os9NMqUH3+Rx+ucdvdIaOmknTQHXUdjV8lTwazBZB
bGEl/VNugmPe+ionNe32F5t7TExHbBgArrrCGPU0CEKoM1YnKFxT3xWZCPhRUFHwcJym2iOHQ1ru
7vVW3kL4WWXMkzw6bKMkR4n4KGuU37wJ8vHBZYNNVkbeNqbqrnVDWzPLaOjurO39AF0Zr6nnLX99
IYUSA2wkzEV1XfPr+CEq+a0aLswYWsitzivClfsM1Vj2I8a+NM16JOntxG4kyjp8dNZASX5E8h8B
EDro7I8mWTb3aN1cSXyTG7WYQ+kBGPqURzjQ6V4gwL1oK8JsGZceZWPBJpNVgfe/CDX3q4KtBl4F
SD+8dvmnbGE+UnNBlvK21oQ21/D2eSjE8Dwp8JBdrVt8iXMN3YbjMO7GVDR9+KYE34cdzDsur6Xi
HH6RuBbYbda8ujC1x/wK66GjDCfQqXBVKHetBdawkfxui2ZjYWYaJ4XQs7yNi61vTnJLS1Bz7eND
mENJCnjHiBPr8w09g5EY6S5I9Ck+S5OMLFhaG9UmdoMZh31aU675Jcr/fjqlCt6z53bMnNdzPvuS
4F6a1SKVdjtb3llLFPOQbCQVe7lZHtAG9dbBlsZuvPvwA+OuL4qrnlau7PYNF5DJFyOGLDzVoAmy
Ies0pW9hr8du3Hf3hSrREbofFvCJcmUc8v8Ceb+Uy31Y3WzyyaPckCVuJd3NDk9Aq4ij3tDRZSHw
474la/g3N3kvqMwaduWB20Uad26h8ktlfqldR9uxGXp0mNjp3OdY3A+tbh5jAlB/8ceAKDGr15le
8zwl0im+OoIy4buNYR0MeLezbnicn2CdoU0tVZlUK+rQY0Xmxbebeo+M2PVApgC1YY0N2OzgSSPy
QtblZkn/7CNb6xXRVHxzrLRXImoH9d0fzbiAxTykXL8LtXORe/DUZldENmwAEe86MLaE1Ts3PZim
bKDHsqzQndBKnswitFrejSGZAS/o/Rw7t9zWDbmuEEfAXAnQZ+zsTDWaVnHVmjNy+odi8KwJoS8s
81z7mUIycK8a6VQ1byWFZeVw7XLV/iZ25L4cezQyior8PU/B/wl4a0y0NzOExQ9vjcGEzWIcSDl/
urvKVhJIdtwFXv8LqPD4BOybYLXKcpGH+UwD/MH2PxO87z1n3xhPKZC47IxkYbiZCIYWy1BJ2xy/
uPtNz3CqdszPeJ/3VRXDvOyO1w5yvgjRWXf2TcJfnF18RdrWGkyhYtSx1b0+akX7Xm6pUAqN1uM2
ziqpCTk9+l/LD6bOVcc5/RLefuQjTSMscTscLTMRn2nz5tUzbxeIUbM/xbwD4sMWhrrY7fA82IPM
o4GpLjqkNkh5eMhYOkQDvB5hJcJNjLZA63GwvUg6v5G1oBANxRcJnHRWUsrir61frlshl5eN4UGc
EvyOL6G6cPk7mQDUQoeFNokpul3GXcw5THSNjdepYCgHqh4rdy6VDR0VGG/ECkExOH7Ou2+K5CTQ
fnIhm6Otd7E+gKcpG0ZMJC4B1UFwHlmbGQQpxtdGaQoX5x/9enqtMH/rKKSFq6jr/vOd6+/n/bHH
uSF7g7zaiBW0XAxZF8e5maapMJVwngo3Jwpq5bBDzeN5yeq4lmXE3ooZbpsdBU8/9UOemxo5hgjU
J1D/Bpq5K9bSL4xLJbC2rf+SPG8/0hk+feo5Lfqjo/R1vC4C5rDUuhZJPdy1WqN+WnTM2E4xLFRK
U8PzdZ9Zzw3NKlkG4d9JekxaVmccOb2e7uXDuIdMG1Y00AQozyyR7guhSSFkz/VskerQWJZU3FvR
+Yktmmi/thDbc1XPbbaUhymDvuxrOw6SwBleez908pQviYEaziggGt2tYRFPm5gzTqWoncuePVR5
9xnRBVaBXQpbFrHKCVvWiWCOyTw/mMxWTCYQga4QbyDKJ8Cc26aKNxLUP0UM5PNlIQpK3sXIVu/D
zc39zsNSCQr6pvd0cEh56HXvQxIX41urMSzfvSkJ/ZjDsoHKDfrfyJFsIPStJS2cdM7vY9aE/28s
WNs1doI5JV1StXfbWLSPb9R6lV4C2Z/BO0L3wwAVXN68PnXEghxcFdE4GzZapgRAf1ZMMHpXMs9C
9tUq7F39KF6Llx5Fp8AB0YjWkIWYLz2unKpuc4mO4Rrb0F4O4K4E32VwRrpv9eIahq7hlAtxYQa8
bArzjMg3699dN059VM/2OS/As8nIE2pGDIcIMIl7vwsCbCSKFDhiI0al1eLzlGMkSKtCZAW4DW4F
bUa0ik6fYsX2D7sfeHONWxgv8/hbmUNXF1tdQRGf4rVZdDMX5lNmRcabsxUbZLapuYAXe0B2ZZco
h2YUdysQSsnDG0AEoh/NdOeXScwTBO3+RPraGJ5MC6J/2mKihzSqNnSZVPPGdhenWZe+7MHdoSv+
ZdXDz7G9iVB5iETaqEVtgiNSjxlphlt4u9gX0oxfVNlCVxJqKHY+EdYXfv4GV1LbP5H93RT8NymC
ycOk5Vpik5hPyxxZudxfIH9n9ey+c44BhM9nRl09nBWYFB7UOXTzARAdWwHKUjvZoF7n5ePm/OHU
qo6px/IcNFiKbEZMEnziWmNr1iU1aK1jvIFUMf6AhZ4KU2njsSDzAGSoDgf+xl5e8BnEIwAVl3Lm
myZzHJ2VB067gK8COo36bMRFrJhNCOs9DX4TFsrcWceN5PVFqc3mM0AEOJIHcNv9G7YrmoAMyqvb
PjY20OwPrf6aa2x6YDYLIdCS6WPF1vtPUPdPofcm1DjCyQxhxX6TRRKdbn4R2TRxfJiFSFP3y1he
YosIrCrBLx+6ID9iB16cWblfPr3lG8KqVNzgMbwgeQenjaioZZZrFIIlDm6Rd+6/0Csv6799hayH
b/EGehbtd9FtVDcxZPZtDjBXADwndroOz/4bE5XqBTkizODo+YJaVLWHn97q8SzeTYcoYL2hAgIV
dbCV5VygG/wFYNosjIsgnVttzK2CympGOmb6pWXRgB5FRncD/E5ae8ajM6r+6nQp7L74fsqVjjlQ
OZdUdegOiFL53hP+Fe8RSGP7LvmhorRIwZaJRPxosIcsrkYuHTTUB+5AxF59NOnipEyFeSVg9394
EeiSv3MLZFpl8bzPVyZzhtXZw26YQravQZuGIMXjV3L1GZUCAwJvJczL0R8cEM/+HstLuxrC+mTk
JM44vM2DUS7oBI4R5hBcwovsTNs0s1fYIxzANZ0gUBIpIjZQKU6KYhljJRBFtHKZn5zoOgrY2EtO
X0EiUCDfva13dtJf/yhAlMHxUpoxNb70qBsY2qn0BxBLIeqIVGTmZ14bSbFF6wM8jyOmgZFLDEXr
xt/9Didl+L19RJz6X9w+SVa13QQ+zvd56nzx8zkpWHUM/EDhC4voKw6VgRSMmkjY/09six0FTcNL
WjjH7FOtOKgjGrARCJpk4yaOYZOimoS6QDVS7Lly7aJsZ009NkUhZvqLPKNZaRkj1GTabb4UpXx3
Vl13HnpPG08nDfouk1EVvphj9kTDAnANMuBizwFmNFwdBMHCnw1CZ2scW/x1m/NjCya7zq/hDIUZ
Nw0sd+KApLsPMY35I9m154ZHITDw4+FH9SRRSLKxj/xzxi3PmQEfy3gb5i63MWdzUhyZvyjaltf7
7Uio3/XVapNo54UgWkcX01clXfA9bP4FjRqXuCnofTn/ZIXvtx2OYV9dlBhzy/4BZ3Xr4CQLpOox
g0Vhzlq7+iDhLgmE7c3eYEvT6mmV8p3fOerOJySBdr0PU/73BHr/6qZGuMmuasUkbTPbz4da6wmg
Ha59ZMZT4uer23WBdnUlptZxnQMo6vX3rj5I+Y+suZG67f2SKAg5tYAMjghUHtEK8XxNNjwJE+fF
OTNwakVbonOL3uGd0tnvhjUmOo8p0GHDkdGIL2EqXOj4xCyBKRbKuhBKtaAviBLuuCIlo8ZHruvs
+qxfRzx8Np4aKVOMulYzIGNuAHpkgvPON3uVR2DemW4Ozix1f7XeoJXyDx16j6dBftOpWB6d4yof
3oQLWiagKCVcIzR1vwVfi6aL1pBhJS7CN8azLIlCTU7AG/0b2h9+eN2t/hWsL3+9SCAf9B2yVEew
F8TFVb5YQBrYTWriDKvlQeTsZrGqChaGftOU19KiXUXiu7UA1+u/+cTybkjNgSkaB4I0Pyon56vD
ot1zN9qFRyy0e7okK0jHLpuM4ATmUxBYbYpn3jMoAAI5kZAZUdFrx/OzKF6fCV5pDFp0qOUMvZ36
JyuGQslgUP2Fhojrvqks/lysyO+al1qOCP5fbQNZzs05G5a+y1JtzmvTeihE0MfzVSWjbvjRnb+z
TD/P+uw9h/51op+czowpX3nJhlraA/6qavD/XFMT1l5TtFnuECm8er/arL1tpiZoQbWfpWVV1585
kK5+ZUiiwm4c0Lqcd+WfnZg+u+h2lFcx4jKCaRqbPcPaN5E+NtsXOthmkumdmOq2HqNdi16Vy+ic
LVYUnYiZylO+U7IcHGkWgXCrUf3rskcW3wRIOijNZzYjgh0F5v5Nt9OjphcYrql4VWLNlT9bWdsC
2BFclmI6p6ubN6ziu9xML4Ajg4yXvLQd2vtTCKDzkzA/j808VutrgqRvRZJtNMUXNGz1Kjf2B6Qc
zZEfp3whZRm9WzuB1aKfXxaDnWtjIr1yK77570A1fcsSAaCRuvwnpr9Tg34rkQomIwEVh9iGExj7
ac+g1H/rEwc/HL5ACEVqijYE3OkxJm3lGQBHS4FCSl0PJX1fx3vhPGtPx3rSRqN1N3Hr3VCHI+Si
GJ4vN+p3o1gT3D9syKG26pgqUjA7thBmX9tLJun7szOn1BqFMs9FYSO0jcBG6IIgjETar+xs+ZRC
nS2oqzukK+ECni6Zpkr64JWWyHGHdxYrznIE5F2PrLCETqi/xJUn09IG0LGhYUlPSCGdUN1Yic86
Pmy1Z+h5BQpflwlq6ITSJ9GVN/CdiCFBtdvHU2t/WArQtU4u4HkZAuUZ9vI2z/fCHBwomuaHZKrg
Q4FYYbO3ByuYAQlNZ2fn/lW4rIbvwuNcChQoCg743ARYY7RZxoyCzXlgCg0jsfnHmkRzJsKE2dt1
lFyBWr7EftwoLLFJoSoEwUltsnabySpbDTHVfrRqFvBPubsz8dyBjP1Hqg44jxTpsmQ3kpy+4oX3
0pckiTJucL/W5cMsVI7Wy8Po2G0UNQvfJCT0Hlaxf59wjWv8UZe+DCakXuBEsR2m+N2z1VwZrmRS
ao6tLQmn7uf54FhT05ZljjPd9vnmBmDFBvKJ+rEcJ/t8LNQmxAx3SiuUYb/6Mxofoddkjnq1fPD6
eCQKSqZwBYv1LB6xuluoD/2S32BSQ1VRqaukQgpT+FCFQisdPi9ZEa7g/EHklyEyKv9fW7h61anO
WtLtHET1otgGuc4W/h5PVxjYF84zADBYGVT14YTzwVkS1y/ukfkEe50fIyi/u+lGOPZkORGjhaRX
tM2X/28Nfa7m4pPeT9CfDYX2unNXfvp/eWVmY5KGKAb6qS8DPieWRb3DHbNSk6VvDkr9YzTrSrsY
q+DufpENQaaTDMoOWegGTgm/Dn4Ni/dIvleZwlfLUntxg3Za83Ml/15D5+mUTy+slgLftwwOdgJZ
42J2QSodVd2g6u1rfbakMZUb9Pgi1/ojSzk3Cqs8SQZusLk0HknXg58bJ9DXdCieWparleGD6X1w
xF4xrrfnv/YQQo0443qnAg6me4dhKIFMhl9yTsB2FifcyTMvNGIp5nufXpURr051eCeuBugP6ndO
kVtQPhtvgnj+6Bncr9h51EKU3O9u/RrziX0nuvzS7HS0tZHKXd8TAtmQ28C6wLkaMsC8/HB1FTMy
TXMMPYJw6T7ctoP/kCyTw23JotXLECRYn1BAkYrQUVih8UavMKthGxuKv4PuimYU1OxdlaJy+BiI
XqfBZ9yYPcQGIKZ/mKqLfBKvXK9Ium9FLL3Ay9SHlcTI3PuRikhcU8AT+tccKB1Apqdp9DVgc2SU
xYOaoE6QGFvF2vSWH2Kg2dDf7Nq5ojHbXDs/XQ8F3vF//UMoY5JtskxM2vJxg9xv7k6xTfGrCxNr
edZs65SqMzcKy1P25oqJFNLX0gfq6EqcB/wz2UPcSf13p9eCSwKS9VzaDFRKY3Hvy1uS3o5FSfDG
nTbYw0IWVSTu1S7MTYAi+ByupSU/A5Kjoj/iARekfbXou4qmRdlEMc2MVrwGIUbI1NRv/urNXODe
DWSRB1h3RI+VxUxPlE1TC/t2Uu0T3e12fM8QOVeHBMmO1126RZCd0b+YyDPt3wkyuFj8ncDfk6G4
V8iLenlbfBzKtLgkrvnX+tfhu90V21+pJnMDCJyPmAGQ+dnEtM15QOiQePZT4M4Rf1VgDI+bcCQl
ZeUeAsX8Ph9oxv/0axiZwtcELZfuRe4xQQCDMHF7Qbdebedysw3KwvbfdF45QxCgkLa35wAJrbiy
jF1o53C3zgr3rqLZQKglIJIWt0AdwgG1+8uYnIOgkL4GoPODCWaV2wVjJAakVYcF+F0dHN+vG6j8
Ismf3jYrM3lAmkSSnSMIDwTD223td68hDuWZrlxzqmW+YNBDu/NecUx1GxIZSwRzDZOOugpkCvkI
Spj9vRPNQRmHyoWfDGxQSsS1DEYDd/5bF+TARREFQCzamELEiucibDVNJjr02vLyUIH4OGQmYNyc
DG4k+BDB4jwdWOoboLERZFQRSp1N6x8MB0Isc+TeJGI/uym5GmXTE4Iubbe6rVqQu83C0aSaR/Rk
Hs/LVNFz5NimRmw7QHu3ScQphALOe/3v4jJlyWxE2dIKGZMjH8LaJFueleiNJv6xny8pz+mlRctJ
ckj0ElfjWv7F4oLUzTWnCKQ9+JPxuxe55XOQhpi8z1S8O+nIhq7vf2zqbinjroAkdIMQqNelV1m9
i5YtCwuBL8lhAWTHvADUbPLRf7J3+tLNGmt9uNd4L3wHKK3YY9XwrwgUcddKq5ysI5EX+1+dFY3p
ufzX4+824hIQMbJtl5m8iwVr7PfoW0wQGDfeNlHb7rKeU825p79i+valS0I7YpthSTGMo9knm/E3
vKzA1r4Ab4xgcaWqJI8qxHmGAcNwHxZlu1u+RpB3mxK2Vgwpebjb1ozKzXY0ToqbZ7V3Rup6LHuF
rBc4DZEWTv6GqMfxNVqqgg7Z8sLOqZn9H+RDKM9oHhsEt+z4ikXa36+3cXrwBQqOYMyUybJu/zgk
9HEdmdT2+ueURs6IUbezreEKLerthcWQPOardPAXbyfDxC4H7WhSFUtKV7ZBmqkIhzsR4NcfJOir
/1hneFUmUpzL6j6u4Sn2dL1X75rjj0wRKNqkNFZlmEfceMJTuxHHxOXp6jiK0DyWvV0bZGtuA/97
yaJlE4KRja068FpvPL5ErtR69y3UI7B9rdrsuZF8XqAaBHSO5ntTVIPZLR1ogX8QzK22D0eNi/UA
7q1bhpctaAKkN0EV/WMlUwE7tJbm2Ik458QHRv6xBEuCDWZi961SkmIKA+jYlSllxzeTVGv6S6No
smOFryP4sF3FPA2t57qQ6RWDfppyDrbI7c87tcaf7QxKbgHRd5YYxL2MqPnu08I8V7cwy56dufcv
7hzGvF09IHgZ5X3q6ii3F0rXvSrp6F9Z83y/qGtGNU9enaZkASHnqPs5Ju0mY4qNzYRmBljdYQMg
6a/UbeiNuO78G5UZOR03RZA5Vn+XmLMB0jsbVEVaT0I/ytowHX+YjIvSsT/jN7TzYsKXfvjjvSE6
6gwxq5GWg7X9TTPwugHnuFuRqrDbvrdTKHBgUsST76eJcH8Coi2NWkItiuKRyH72dyp5mQSBUDN6
wJrJKL69haEiYpj7cHIXUI+Q1Qi1XwB//QvZQ4pSZykxpapnT3VRqpesQu8Xwa8MyEQIb58AEY4z
qvMGdGB+/IpYY1BPTvxbqMCBmqc8Zexj/zwzRSYQxfC03KKUEmhepSHEPm9KR82l27/UGoZTkciS
yMRUY+WS6d5kGkuRTMzfp9hrZPObL8UUflBLk9FHPKmx8gV3BPPSABxepgS/B6nzUOZsEQO51IFx
l/XJQI8oHDWwGyaKwSCpv+vmbBzEQX8mwAP4ccJ1tF9pjngDsGRBj/+Lbd7NQFavQRW2SEaOOJdX
2rdCwdq5sUnhlx/kRgSwPmVCt0PpcqGMjHiO1f84Pd7oAnyCQPKWE0MMTB+cufvJFpgmgx/PG7rT
BTgvtp6FsT6VA6eKr0vlPrIjEP4eUn/jqxUHLpPGd+a6r5Dh0szKKVrOIai2bJSGQ2Ai87DS1ikm
+ig1lZaJhSyGkI8thRvzSX0FBFo5S90o/1P/8wlhGABkXqJz4dH4/+pmEt+f+A7CJSAggG4V7qdq
n9lWp75QV4eVHtDCJMhhSBMTlxsJT0UWc9BhLjPGogNcLsfBhG0gFOQtJpdMrQuSEvJL8exulLps
303ZN5PJAlzoP4kmOjTtmmMGUSZOCxUnAA2+PsfoJgDJoe/wPQDE49d10Qcl4O5QiHPPES/BJX4Q
EMXNCnSm4JPuWge1cyJp/b31vUwWlL1LhbZu0x6GLuOBcmxUsjNTICCe26WpH99He/xsoViXu83N
ZuP9jnrkQ64u+N8SSHD77qkE0f17xCeNxCl1RIg7In5NXcVWyaFISCN/RoSfaCxCL+vzeuFPUGdH
BpkEzsnbY89jXylJTmFVjUAZv1IVisSMLUwbBDWssmyWfjI1mehmPjQeBg6/WYtSt4ZKWEouDJT8
OQfn/Gm3iw/Hqtu1OtnXtNriCue08S+avuxsz6kItmTWt51e/xhcHIrqsdIT9pAECmhRTHRJzcSC
gE1/jY1G/PV6OB3IR2y38M2P/oxS7QZy+F0YNGyBsA3ZQ6km6cYqTF329esz1Eg/Lw+li1jiJr7Z
twSyy7TUmaKIOo1p78CkqK8EUY8Yi6KO8iLJeeCgUuTKI6uzKy28bTsZx1VkoxvHZqvq2KfVq0m3
EfelaEIRniq8d/7qJo1aX9Wx9eQq7tIiklmbe+1w7DPWRSuDHokN85J8Nv3wEWtXOGsIY9+iK7+Z
4RAKx+6ObhH+vKhobAEz2uv2hm3xox8vqnxNwUYQk5Y4r1wOm4vXyOrHxazCa2/dGdXTTB1wK8x1
rw2ZT/Cy2/pOqaDsyOG5i1lzuRp5TT364QnI43Iy2EZ4aDBAaBll5ucQj6KRgnKnUDacBILDOD+T
qSGcn2pgvf63lYYQ5ze//s7XGvAj8SDBl3s8apc2otlTsuULFQmBNjPwyV0PyA9U/yCOu8RuXIel
WVY8yCcKA7VnmVTDAyidA8djEqEII7qhjMScSHYuz/l22CAJVGhI7Tj3gldHccny+EAwncC6BSCZ
lUXXBFK5mNsZVSlC8SJnbikKn/1DKyaHxJhq8mrUrvuzPgvhCfeevI0Bp5qrJnCXG6DWLWSImOFO
FqoIaGhwrTIhLBXvtOQF+lgwHRVpcAL/bm7QGEnhjZc8wWq4aRTvXQyjURIW9ALyUDvq9v44X3fF
GYcd8QvtbGwEecDUYv/0E5I2eYWWQ42f41Q/ysmy6qlw4BTNHzHpErfh+zV8ilfgaMyXA8prYPnJ
LJ64xxofEczB1BWW9wuEnKEYxRsdCSnmWGjZ93I39wczUUyZBN/NEHVlN5T7/pW3nYvd31TSmkJj
AqKofn/cPiMJ4e+dfqgCawCcSuI356KxRpqymc98hKDdEGDrEaBy8DfYi9CrReSqgofq3Z3zpX5O
Q3YEpYllQsWmua4EndtZ6urN78PEASu0NlWkU8igOUCIl63hDA6x4gao0uCEYbNYKGwYz0A39W44
Lb73FRIgP1hJaac+/zj/L8q5PZwxehmot5zqrFVB3kXrJXDPKMMKJmTosFfWsFYWgmFyU2CQKWk6
2ZlG/wI34yiFTXNHQuDhHNZl9Cv+5rdWEeAQXuWZY+JUFGF9CN1pSsBdS+Gj5FTipRGqh/j6KFlC
WiXnKDijkrAnOQElKjsc5kxlQ6AmdX4REJ9cVRtCeYFf+yjGUoFdHRFQisELu6M3TM0XT4pGFocY
6CLa4puwZHKeFnq6WzBMAwtJ6Jm4HEXMRZirZUhxwqub+KwgtzY6/yi6jhsUfnX5yvwvXZzKIAOi
GUG+fSJe5jUl+wnWFRu1XC74Gj2il9bvY0aDtML1wIo1rHLDvg9X+HyQhKQFQypbEVdIJsK0o86c
/idGwgpQdTU55OanEFnFCz4de0gNrDLP/nKyX3MSjp9u5vYZOFltBkgnZlo8Iah/ClrT5Jpt3uR3
6DG7TW2XRqW6sRSYrcleokEiCS9jW3MygRvMYhMv9tSPvCP78hcYOTnU10PJdqa0ZsVOpArhN5EB
hBsv3zcpCBQmvqcF/W1vpqoif3EbFpDR2FpQjb3lL1AO7C5Jh56T1DakAoT6i3sfmCLPUoJ3mU5v
OFWCdYRnR2qtZ1SE7adawY+jMzg+HlIwOSb8OTbUfBIQzsqjysvbzmrIiizNZ8oHb1Iz4gwQci0N
+XrLdEWazX/sj5+lNO0vRRLzs4OGGVMJIP3O8qCZ6UBnvTQGtP22xGwAYm98BnNut2SpPy9zOJZS
L/v/MVjN0Jr5EsbsFciOXFA0hBkDfhvfTBdBASPQjOA0uopvWjfaCETnmL6ljvh6L2Bq37qEGccH
1mTHl+YA6myl0vR3Pbt9IvVm3eHbrp2VJje7u2SE2R9UA8k3iexj1/FjIgh88CB+AIuzgq1IwDkv
BSHyAJMb92187n+Otwh9qqwEvT3nS/Sl0weUYZSKMQozJ3riZid1VoInWGnzJgL2VfIeQZrcC+vY
u78NkvNfeMCxprIt0ZkJziK6sjIoy+mGTHu0a20xRH7M+bE0oBB0JQsZ9tMHI3gGTXoh7AtulPMv
mNXiWJs/jd0VaQPEc3XG8TEaUboz86oUPCJ1gsZeswCsBQLwpyZWF8f4jwUAYra8ZV1egPkutD0c
dmuYCYaV2PECtu1sA6g2gvUdtTP2DdJBXbVBwcUGicEWsHlH3UIZIOyyTuLYo/8zoGlN0+86jgh9
DrmU16AUMA6ncqMDMhHMUN59IrvQxVQNb2vEcuVCr1Fm+A2Gi/hroBnVUCSabhXOLPai979BpLJY
XvHdcC5VXAODmdftFwQaBc7cS3ptGNGRaLwtrJNOubEGFO0hiSDUdR2772GLDj8Dz7hNcyVRZRgl
I0EziWvpKeEgGoFJmkQJvCCsZ2n4SviTmKtZ1HyKzhagMWzzFGXX+qPjz6o1/V7yEq/AiHz0cQ8o
XrDAFi/MH3EsIM+ofRv0Q+A5z4YBBrMJ2vhFV7aAmNrjVzaNbnsb9qWUURJJDoCv/S2/gnNLdhtr
7oU/yXsRZFZnlS4Xav83NEhNQNK3pzzp7SvkgUtRpqxC2K3wkblJ7fW0U4lFaP/yP/Otku2kNuX0
ndXpbgf8VLYL97EX8c/wQKFgMxiA9cfmBKhuPoU2teAS8e6UCK2zpuflZ0RDckN5jgARDPKGy/8F
V67qu/aL8yxTjimKBZZCqyYJ4O8gXc1Gif7GOsr5QMQmGEvYvftODv6AZSSz4sK7Zk0cOmVcKrin
KBfAqe/6NEmYGK/MlImiB8rAbaL2BKfEMorK9NEBPkBXP/XZHw9x9y0Zv2T2/88Ze0TMZT0gelDk
lquDNIw/4jIFntGcckfB6t9YEio/7FCFb/1WJidxY0R38ObbB5Y7dHztFhXPS0aMhiNmkx8BawPo
PooOHsDIPR7O1boiYoCscq5ZgOriRq/DZLxzzM9e+fhW895hQKa98Q4+F7c99Yic3EhXoC5DCrG0
SRCopHo6r4ZXjehLIlTs2B6GgdKhCdZVb6UDk+i1bI4xb43468Qca/EGViAyZgoFQvFqcN7JfkFm
3qce99UkJGWPQrcU84yKkd5vcCzsmg2XENRVghPPoxOUcEUzn6N291rbnpHv8cwaVCjlCgiagyse
jpOtkrnTBroIkz1SPPZxrYcg47MlASv3jspkUvmkYIqABVTi4rbu//1xj0rN5lA1b0znOiE8JyMZ
XLg/6nvvyn0apil7nc0yYbXaz/EDiSTFijOrhTGUpIXnWpV4p/Mh8d/25ys9OdT4PLhaT/DINJRf
WWH0ixpmJytmcndyEmfnxsxgP66Re5gnyxgpWaYbwJvOG37BHDIwYbTJJZHQsJQEgPB1+IkTzfJs
9NdIPEEczBH+s+cPP38Wdn75+bsBx49qKhb83Tdd7WlnEoebSVNHf1Yl3CiCjj9VNFV1xfIm+gRQ
qTKkpqWRsxjNjOlgIJ/iT6erfDekMNVAjw9+FA1MB8THx2DBYYpqdh2973TICgZT+/jwSvCZztjg
sV/hIfI9sDZmny5naiMXTfhp+uUL55/Hu9v6xWrRzBUEpcxEbp0TFggcHZLHEjLbrePxkJI+N6Mo
inVi/UmzbI5wmxXLUciar5hDerYecFiyJQeb4ZhSSlLNj4Laoj+0BR/aMEMfECmmgH2q5SBgjzIn
iWSa652AYJoU8gnD3H8caA8jrU0a7NhMIDSCVNYme7el/731eUiUGFUBERv9c8fy5JV8zA7r1yuH
RSPfKFOCZERY0OfDYPZiEVOma4Ku4hp3B/dFNo05m/M0yK/qIjocDc4WJCe7TTDaam6/doY9Eug8
ukyGf+FddDgS6m1wkrEMpyHN8SoyhyjwpIZ1TbziUmOwxPSQyrJ5joE2pGJucdah8hZKLcW+R1gY
s4UJlpk1T5NP+d3GuA6z67Bb1gPGG21BSVCIXeQeg1ACy6wfCmnzH/KcOUR8N9MovyxE31XfZsIF
bpH8T1U10JAFOy4i8GYSJm7+MM9G8HwJG38TRXL/cQ0DBVauTQU0rAJ+vEXmvGBrW162FAdE8JlF
1Q0TleWmWI+buUiWpCbi059m6WxfzihbgSKq0bgRLeoYrO9UCWrXiRMTOGkcvh4JpdiKH8xIvgLr
IiLT0wLDl7QVetbjmPKQcOOE7AyW6QlGNYqgphreTkvsASwSQCJZoGPj4C2yXPwCM5JXfQASf0/O
NBoLyROYSM5p3IFC7M5yLr00ciWKICWinHtElbP4CoO9v27HXfAV3xy5hW0DXRevJVcH/yTSB87C
O/Bx02ilhb3skMsjx38SE8NBkVDeBO21NFyMOgK8nk7/QqwwycWm8UAF42uHSPthhxQjtg25DkF3
zgh0oMMbA2UBiPo/n2hvI3da7n4h98jJ95IgAcr03tJCukbJFae4VuyhpGZwaOlsth7QsumXLHlp
DsR5i99ozQFRf+tsYzNrh6Dt685M6rVA1nkVm7vIVhCVfFay/Kndnl9uLkR9LiUBl5Pwyx1C0zbO
/mkjhSlKlDt0h9g4B7FSET89ZvBS+0rOOZc7Roew0T/UH6khgml2eYh4QnrdVAIIgV/tJaGotM3D
kpcW12QgM94/zXCOfIg3FGCNFuDLSuJPHwn9jZyy6J9KtFzJMyvlO2OObIJFg3dqMVzyuQsy/Z57
AVAi2j8uJaqfZLWi8sBggwDOQvzcr08bhaQnS4bcVzwEY5790vE7+GZvqHLlfnQNvRc+DQnIbF1s
+tEFU+lqBObEXVnYN/7+c8kB2WJ7rJ7cUIwx7/RR8pIXyZV+wETukYeQaHRVUZYhLDIki3aUwto5
SUueJwj1hrYNzV1KWbFSTmLfrU3xo6gE7ZolHhqgOfnLxP4+O3i4s4vugW1Fk4QJCD8sAUwSf4Xx
sQ55oLqNz9F+2k7FlWYG+37iAl08YTj4PfgZGnrGwdqYG1loVEfItHFXV5XqTXisPKQDAgVAiDFd
/gDxkT7mwiSA5iY6vBl+7Od3D/2iXbrkDppwWvUsTi7LGDlnSioQ+0XwAZVNpybqyW6pzGt+PZcL
FnrGfvmFGER1CwmJvfudE6RQrpRAOO3bJ+JCKnrAvEbUHyM54HXp75g4W5kPkwMmV6WtIG/FDSGe
6bWkAMuwK5ax2Lae8bBPxoY0WEo/oTNEFb627IlSvnPC0+rwG5uVnoFhsR+/QHMDmFEndEWSoTP8
S7R3I9Xg5RGeVshVqVyZbnWaIJpqcHeFECd3iokBrOdTqHRJ5tsKjdUHhaoDH8hzP9W/Y+pzTm54
fekFFFIxxXWZOQHiUimDoABTkhipgwheW7gULTx87u2x2l4UscYxPAyoKZEFkpIYE2ftrJ6TFFQ4
g/SZw8NeTg1QqpdWJfVNgB1pI/peFwXtZgSFt70xzXH1r/UFvxmil/jA5gx53BzxuisJdXxCoh+Q
RAjEbrRiI8k9hjuAiTgQpZal6+502wlfTOzBrRfrqpSpgW37qqHrI958f4fAb6VZQjB1OZfW6cN5
ZbHqYS1uEbHUHIm+k6HX44rupA+oehjYwn6M0CU9vI6064jDSDrzc/PWpzynA+5JJK+3OD3COHZc
K73JZlQgTgXKQ4Nxqvs//oH6s9l+xEE1aWsoBAzfjokLcI/C3/GB6AE81RKO/q9l0f8Lvb2dH7R/
G4r/dDZ13X7JDg3YLj4whm4t+goTBM1VDdLXbGDnj6uUb3F7PamJyudW1G+cCXp7ORfJMi84bR++
n6HKkCPZiVaK57MDFG/gLQk72LKhypNr+6UQli5GrZrtHJC14zTcQCAQsE8wpjmm+psdb5DKJuMw
+lH0vN0WfYVtoQcXthkzBrs9iGHg5unScR5iIbnea+LkRA+eZa6sXn+GzhFfU4TXkmlQdaJf+D8g
L3pGXUVAdPGbC5voczz9WoclIJ7ZIdjHrKtelK1R5wn+Pg17r1WENug5Yml2xpmt0/dYy9OdVFSS
Ye5FdHe5oUfUMereDl6sYADABcZU6ziU39onrOt1YMyN9pfQDfAt0DxyJRvjpnWId9Wiu7SZqlS6
j34KmdREmNK9+lynQSrp6/p2kz3WQ4rPJdgt9lsVstCx8f/4vReO6xVyV68atC47UE1Yn2wc4rsN
wYdSIGHWiR7MX6U/HEFhyJPVWGEte4u1HWGOrTEiStuvQuQFgh54H0ZKgU0Z2/X3GqzqtivWduuD
8y6sSRwBZaU/zWbR+FRcpJQpbTi/6FsMTbnX3nUHEHuGPAtsbT5SvdjX5muW+1D6Z7igwdL+05kA
1o9UH2Ngcpf9KcXtTxvdU3+hJzPfRRhxBd9YGNFkYUio/ydlHJW57M2OUu/CgGEpdNjidvntPg2i
9JxeK8tNpFq7V2CQTeBgXjMBrYLwgSIN/7wKXO8asedPxBYvnhX3yP3geOiIRrJJILQLY5ByCtZZ
E2mkrlYtwm/wUf/G3PWIKY/6v9Mf6qSjPE7JiQEoT5QO8mJ4hoR1MoLob3rO05XgzrMMRGKbkbQF
UjAe6FHKsh5ypIOqL6r+AM+wj3W5xQi7vvkPg9rhmXVQBiwu5S/OmwY7aAeVlF/4zufBPDGV8E/u
hTyNCFBHFW/LY/Bdy43NoucBdEqrJ2z66sWTtnspZ5GFd1M/IRvhkFLrmGdonkHhSZcKJRsZa3LH
n6En0u7yPLibjqoc+aAWO3SvwPBDUAUwmrTvhqHpbEYFALLbiaudNrTyJfhospSPoSp2ORv+wBmW
CRQaHtOTid143k46XLGjM1bbyL8kUQw8Vd3Fe5QpHfKYr2p8vNIsFLcViSs9u1aBbezTfKqLkQPB
EluLQOI+wpyUcICJMII/KlHhggZOvnf0lHyUw5fIHpDEW/6LbpX/M+OL7NK+QUC06ne56g1K+Yn6
JmvWOsboUgWyAk/PuC5bQ8lUxuAqdvKTsBiKWWdXt+pSOnmbA9IHq/Uzs2jTvfvblBP7IzhGnWfN
5RUR9mZWJQeNjWZl92/WHJZe8sAVHRvSOw1qO7zyquwNjePt1il2QCsYA0RlEg0oorbxtYRzeMIF
iiTjqEhaE+9t4UuoMMizmsdFPOtUKT+cT3y/WorJfv9sm7rm3pYbH1p/iLKzcj8khWM+R0MIyl7l
7gGOQKPKUCxGHcCH9xz8nfzybSa05/oshyMXfZb9M7LF3fqwRBuoRL/EYIRi0LGPN5N44SNJILEx
knzCHzJ/OLh9wPksoSyrRcpuEg+AHFTSh/fe9DvHHCtnvySSV6bjJ0iwjlYtZJInzrQr3TCs8OVz
kYFG+f1fzg7BGfYFbrQdn2+PWNpWmk6+sGBlwF8CljwzhSEYQ3XdiLcG63B/Xd9o9yLnd7CZTjWw
7Ct9WMwgAF5dgKe3BbnJVPTw0tGxVYxzjIICCdz7wlXWzA8XBQ7Pku+btKndCLqcJl8zHFK6GAcb
UP5+KOa24/GcX0s9fUh6ClAEBOLfvtcteq2NkWSRs8CXavswt04RtgRlnx9i0cKlxF75+XroThtM
wjCU2CNiiO4Emrk1usjbvOYM6dHtC4lIhGbAUi6oXks2CCLI0kpoWXXwU4cbyzZVjOPMR2zm9tGi
0tiDPCCIGGQA5PCxV7T4vqjKF6aW9yiVSP6y26a592w4ShJATOVGWLM4nkhbdzKuh2Sq5hqBimS9
73f3qvQ99lRL5COeU1zpDxInQie6FsaRbsjeiDztwbk3pGhm12iILcJmRLf8HvKxhtwRkUvvgsXG
4DsNxozaUGskKDvoMfnXiUO1yV0j6EpfFkMeyY26stwfkASau+6KAP4ixG8k56wXc/ViIB9dFXdm
pJQ2S8RiTW7Cws9iQpHPDu0suX1xoLEmHv7TOeKPTcOwZF3O2GML6ql50r/qkQMNyzjFPn+X3niJ
MQ7uzUgLnl9tDRTkRPX7w4LIsmPPPKZWDbWJChJ5BkmD5QRkWi6e1VaFDdDGcskflOlQ+8glaGgf
wO/zgYZk5FZgXWqgD0OciTsmpPwadQaZ7a+9yRBMsFsphyf8HCKRmaViowM3MBToayfu3yqW5nQ+
pQd4SjPz7RJyCpqtfcX2BXWO5zMkoHppuT3hhwHYKAzradouQ3i38iR9ak4Rxf8eic40t4AXi+Zm
I4ewDYQIzOcFurovMlD2gaVbppG/Xqz0pwkrcG1mdXlnNEa6nWVQqiCQ8xPQn9CNs7ckFwoKr51Y
/9Mo22FYUZytIgKC7hChIKdM8yxuVdkSSCzSTYABtP9nbFiYHFJ0TFPZ3UwSRrrTFkB+IjarbdZQ
SB4qNHeHgdam17r2AsQSoSqATyC9js7cAjH+2+vQ/B0qKGmt/gspDAewVkmbsmH9dYGoha+aSnlK
rhXB9E/1a7188FGJ/BZmrsrzcyHHRb1J/7wtaZSiYTcN81dQlpKPeSwtb/99CI1FXYvBVJ768juP
FTdPvrx1TDIy/fpjF5Y/Tk70RtZUaLlj0oTgTN8m+wyCHtC+/oVcU61KAyfOE9rH6MQzSOeNwMNH
4qJpwNqiL6SxFfSjn3oVWV9bl8zGs429Jet7P6RNtRRgFz4M7v3Vt/r2Hk0GZSnKpHjqbsCugrXp
QAiCE76NVOiZqUqBV460qu5NLfN6jkYLduOiPmDwXEM8KxxcyrvH6WuFKWSsvxXlaa75jo7DJPvq
TzgBguvkMrdOlRjGOovQz5Tl8XaBzizqpw1G1GnHnaAjSQTIupTP3IZGGMce3SuZm4nmHi0lXxoL
AisPOG9lXtwFRImGPxSGFsbRNAFyXJS8nucGwJKC2xlUsYYL8n9/K6oevAoDNCpida/+iSCxpB3O
Kq7W/7Q46ME2xH7uvqQ5AgNwzzwKgMpvTj0icuXxYhdKVEzkViMOp5q3/uxpCE1oUeOiHV0kjm/D
N3/cOm+dQSalUGlPsh03wZGCqJjx6v2h8LL4xEIVShB5oob/jp5ikzQPtaH4OKi+QuPZwww6bVz6
UZqNxmlB6S7RnmmkNWKGOfuYYwPczE1TD/h5jcqkaJS/o/rW39R91h4yyumZQDp98UZDZzvf6zx/
7tngAz3cGfhANZrFT96gtp+HZMMQ4cqUyze3Uik4D8uEod2vdfC/mMwoNRPyDMS1dd2rDH+GR+Wd
Mk1XsjuQ6Bdjw8XzGVpUcGAeXByCbmiNJDSGhnfrU/TWEZwI0eMenzQCIDIdgo5t0AsDVR6wkQQQ
dRzfdy0twMaFuxH08reQPKtb4MFFTsGeQsENvB6vtt72WgD2Sm4urn0E1qTEV1bCGBFJIcB3No3B
U2jbFPlXR23uxnDzy7Tk+YqY4yCg7gzjXJ3k/2+2jGukSjyIQRoHINJKcIZFT64EEf4OsWmM9nsj
akTiUGbwZmCSxS50hIlUSZZydCj6P2/SByh4TaQ0aqD8CxWAnxtkNL2NlqVffVENprw7X2AcxVkB
26ObbpN3PvjAcJqfPrc0XDJBfkLqn60e2ESmWOVU1iajtdZhX67M4eFe3vXA80zM4Gu1hdNDfSF2
QpqySCD272lj260afOCtUDEoXdqDQcUo2rpaep5fh5vTG4YyOb+y9nnoU+xYWLyU/amOXImNN+6X
vX4HlC4+jpvlpCtb2ReNHYwHNZjB3AxpYaKkn3aGbgOEgPqbKM9vmW9GyycACDbh9pfx6gD3XFsu
MYtMB8EFtUINePZdwbr/hf4pGoRGJq6Eh0xGsPR5sYXmqmS2bB6nLuXnaR+zsc59XoAuQaW4WQ3Q
6AQtlEQ4j6rH+VUArtAblU2DTGTi3d1FriIt2ycD5Y0ay9ksEGrgffZatC7tijg7HBsLiUbA8PY2
pZq/jmqMWDMpG+QqhG8o8mwd+IJR2F5Kqu/ZxpILfg2GT+FzQBFmVMK98bP5DzyhdAMxpSIjcBfq
F/N+fA+dbJorKM4hgPdfhs+/PTv4TKqZCTOrB2NiU+seQ74H1XeKpvjNHImpXRX81W41/96OdJ1S
Jj4yyi3wp7Ndv7r6Mt8S9jRbBoe3+Xsoov11MJx6OMGuTvddhaoo4469G57yD+rmzEHSYdIhNcZg
luAuVzAncJN0BZlfh44/rbwvobGEyzIf0wSToe6DuCXQCeG7HNNXc1RZPE/WW0gnDI/FpCQhEdGH
w4u9XO+0dgQBa8SYq47Hbizn+/rqV7um3MIiUgTDJANG
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
trQQGtv+2xFexFpsY3I6b16ZbwVZDJjdI7bQXWveJ2Sj0LiplC9Bjl1Gd2NIaVmrQhjhoVUYM0bT
qWcAfvFgwiUCxLZqMwJlgqRRUcUfSQct53L+NuCg7/+hmr2SzXTQ053G8hR2c8eZmC/zimCNWQBW
pSEqjQCluFZaW68rjGNZ6IsB2TVmyq3j1zDgQv5N1BGPC+1E3wILJjN6x0Vy/DL/yrByjk45hKEK
LMCSdfifpohW+XADLXSiK+Mt5orAsafPJ7qFWaVmgD0x7c+pi4Iflk4nYyiH3L1wU4Yh8MxzQbH2
pceA4GxjhxRiIlZmShnaZ94TDbS3Ie1UKBE/lw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8880)
`protect data_block
aP8Ldc5bo3MWtWTqBelvpLWpB+PRNJdAa54SrJY651CI0/6KtEYTBhAkDo6p1WDpOhuT+5tVwANB
3cmI+Tiiou+BhObIVPm6dGLnncfPAA9PLX1hGLqMOPrbKAUJO5Uj9YkiLXjSplB12tMEV9jGWhQ0
ti6kb/APSMDjRovdI+TBuOjOVCyQ+7eTMD4ij8QFqXMjn1mn0nYLFD2foOOSVcUZT9cOH6GgsjcR
2iSZEiDza5aqRiDoYtttr9WIPbJ9oGWyjy85Z4EjkhSJ6UL0dZZ8qj62DJ2fjze7NUc4P/qtHzHn
HXdiM8URf2+9PaioHChSM3EhYGmHBvdAyYIywi0w6EyLe2IILMlPaevw1KOfW+mS9odvdVG7irwc
itDWFNbg8E9zdqUJTI5rTXHcibxTqZ4utf3AvrIAgvzqkXIh8vNlKdLzdGhYtOFAT++0U2ouZNdt
hseiNyviuoPJQnyESLVDhr+RVEefW2dV/HsSBq1UwNHJWGWHEPwcj/Xw4sTN6T3jtvZ50DDyMWXj
WzUjZnFKXN3Lw1pdCVN+zFh0TX5h7EcNwBpTXEL8oFwBFu+04SAl+XcLImrAyoxWFEljmcbCV7bP
JAmbE5Tb+4IScFoJn6dkbl5KVYu6AjLkC4IiCwT68Mj5jlN56wYgwUUxD9HrSupa3Ok5zLN6xKC8
cMc1W0uDp8f2GUsafhjloMJXolnHECN5dWYfOrlE89/2cax7KLuJEVVC5G5s8he+DLpc5eOcp3qn
+RxeN9AGPmuk5jCU/z+rkylCQHgCmWk2lAjVQQ0IhbBqubDtOzLP1m9On1vtHaI6asyhfzZO2Aha
4RmNzHL7kUwJH+gbNnkM6ZXxx3lElEauWSuU122kvmXrxJIsXme1tAufYKKSc9s/dwBbRcnIOely
cnIo94Bu5n2tyEM8mAcbxAnBrp+VEhw//v7h73WQNwAoulRcBeZYFn9oKqMBERvj6hAs0CcXRxp4
qzJ4n1aOyEQe/QLINDNPaW/7VYbKYXmSTaOUM43nNLeXdhpMk5i91vfEnNjPWlOcUP7ZRN5GSasR
bKI1FAQyb+3eDYlVxFEaSe3agzceBkgtApHRZFDzDQgoHOsm/rsE3WW0OZeMbqeUln2bTP0zIp7o
95AFQ44iZ1Iij0OxWMR3YEBgdl6qWSyIriHLLia3DyVdMrjA6SsKl92P2weoOxrEBjWbCdjNVT2o
D7k7uPpeGEo610K4pjPT/wfRUS7g8ZFavpwouCTKUq1Tl9xBrPH6hhEr4jBd0O/HxdFRhnLFXV76
ST6epxZ9Ov+/Bmvp78RNEyf8IZHiKQQdzC2XtsreLaoCZa2bWTGJAXOPCzqLFz+/e0RKHdBihx4E
dRk2PBg99ehO3g/+S980H1qvNwRJDVG2j262pIo0oDs1rhTKDe5/ZkYpnkb+4jIcvE9g/AYRHrxJ
Tr44fXJJUe6G1WERdgtQ186FMsTGBg7BZDGpBop75uNul5RiWtlSLLdVXZEHnEdxx6iG4ALepq8o
uFv40VKzMjM0PO0VI8uW3xAo69ToUFlNtIeTch2AIlAids/wPaXV1lcF3yGaq0Lx1vtVrRdp0OKq
YYrirZApZzMcOZzT+BXiXoeY6C/JCIuOlgvdCFT0EkxlhgJjzAAGu8nf+Gr0udsAfml82hgbcd0/
wlcoChkdaNEDb1p3Jmi99TH+J8LMaQjFkbiQtktDFxZtHa7jA8dwmZX29YCgtP7ms+kS/lEa7K7k
a2QSt7LLo/XlYFUDBkdjqvNxsEkBVsvsOgihYH/PZI4jry2VvrTm5/J0ta/RDCPw2pZHJ6n7NT9y
fVtYWCm+hoTsZia1DOhaGg5/ThBY67M+WBWD7tqt/L851P0QbAfPaBUxxYnhr0MZ8e302yiKhKTF
VpJva0q9mdxEw4XmeZrfclR3lpGKwarOTHmgR7D3Uban6AbfcT+hmIAAtRMLP/oeVifNUvXkjHN1
L79YPadsJHpJKD19tytZpLiawUCZnZLS0dp2hZPW182kj24kGgidvWEWSsAfpWQBMCTEb0BMjptE
WbLJwVwm6gozN9h0xFIH0u/Q8CVjMIjeyzu61RN7MH8YRiA2C9CromXgg4DLK6fM2jrYTnlzYzl8
OC0UQc7trFoS76jgxLSukzu5EdQlXzRAZfjWwqnphWA2alaPKGQbxf9Bbj3piwFMBdJKG6/y3Xxg
cYDbVfkfPGnV3/+Eq5Qv1x740v/Gj6O+CX+BKzleL2raEZ8uV1lVDGGJY9J2QR+xmE64qb7s4cXC
Z1j4K0smGoLGWbtXoIDoByisB07+Lvu71UHuA3yO99yFVyDVWlApcUqCd1+8OHQ8yr8IfKJNoCWq
hVC/nWZHdvq5q+9W426z6m98VJ0xNifRwToXQ8q5zoY4VNluyNVAEfwpff9dVt4WyAIAE6dD+tVv
21Dpz+Qtt9aJIYDaUoRmjhN+2WUOBZ6eeMhdLxJh+krEbM+TJ7aCraeCLCIRaoNbn7BVb/tzXd0V
HzVMe/5e+ygz3OMOYkird8l7iqTEEw+tApIQjtEBtZxu2mlHhc5oQBx2Yg7GzQbr4wUGpEzdn4uL
xk3eO+IsdCTiq4ExMgV6ql/xGU4yz3nwhVXzDwiL0DQsmtzoUfGoNjhb9OIKl2K6EhM4L+mv/p5X
YnSJpfvsnLndWd/yxynGUIQlb/lYRMdgYIiMpNqk511p8UWs6OnjVfL1hYmg8USG+AGliI3O0GKw
5b5uyKHFkwzpdvGSNhciaBvQ1mbRpj+0nLC8600gVd4wZOWD2MTLcviVpVfyZComOoQQaNd83ljl
1ROqU97crlLD6lEvKII4whob/UZnFuMl2JaAhGSZsTU8NYHjVEptDlHS5Qg5vHB/8CfHo3mGDaS4
QQrFIi7aHLK5S6psUpM8UMZM2QkrruInyDPgpl4h+6WYU0YaGaNT2XXSRQct9SUyHfnDgqYncFmQ
oZD3awwsElPRvfzj4x/B9EjOg9kESYT7leVAq7IWCLZFtJM6xkzGF9hkAFoOP2/EpwZR47vTQoOY
Jkszmqjapnb5+o5xPinHjG9BOzMdB0BGs7IY2ojX87k7oBIKJNPfYUbkinhGmYzwDMLfwIn4sypE
V3TkiEPK5LYIGvx8eVezd/15e8xr7kY4qpfX9Ie4cE4WG/yeDDYlpxVVfJuPfz4ZV48J8pX31rDz
gmE1ZIaqiCIQ3RR/DbxnWTRe5YQzQHwbtHtXrs0NIRqnncQmOHGMDrr00C5Fic4TV37t7yjkTvL2
rPL65Tx7+vzOvpRk6KfTxZVF6oXMLaJHlUFgE5ocmAWof9Mkgz3LgD9UPHCrXT6RPXDxSwykF5aj
9XoALNZP/ON/dkhIwgO1yeIFpbK+ArCpeeT5R/izoY++Qe2nGa2LVdW1RBeC0XFcJiqLde5ED9Yz
Bw0GZ4ltomkqNah9BxhRgsIEZzKWSaNcswe/Q+tqsK+QPDGRyAvdD7OlTa7LoUZexo0GiX9/golA
QoJGpvKkuMEr00WARbAENt3m0pbmj1uUWGGkG8zfQFhSjMv0CgJiXqlnZIcTktMNNvvZbcp5QHgk
gFvnCQQ4wvnMi+0IVGB7KXTMIeaZ4VqjtDQ+y4N03asT13dTeqlwoDoTwY/oCkpK2eE9juIE4MVr
Z7sCspk8A58PhFSayPZksfytVB0f1ht5/nJ91xrIS7BL59jYeBK6d6+vg+PoXucSqTY2OdlUhdGB
WTPAfoEYLWBqIgDj6feCVCbzS+eMdy4g9nHP86XXSud/A6zOrFkxIxXyhtKDmAGktfsDvrz/l279
MJ6paDvxqmngbSptwCjEVMSC7DjSGYJqnnuQk1b5XrDThZaCCBRgRdpcN6lYkKml198x0clGgVCl
CamEwZNx+C2syozZDDoT7x4LqrSfQhgWzQYtwti8FhQ5HN1wwlADl7ntGi/I2iMT9iCWIRwNG1L1
ftkjjXlN2VWKlWkbdTu+12zs4rG0zoq3coGg3eMm6Pr/a3ERhwaT+lqfbsVmoNlOPePYy3BDFi1/
a3knrdUacdgPKg7qMByfwamrjlgJwmE77b+WQxy9wWdWYQlcP5+U3eB+HFm4ytZQmG6lXiLWGzlw
FF9qlZA7PtIPtsMWr518Or2CssHyGrPJ8ewu6OG6FbsY6YkiMQcxths/SzTSKWq9OwVt+zszXQl9
al/CGm1aDyZQaYSJnb7lvjdFGgWEZR2Kdh5Y8VbxQRIo0q6S5pmX8N++CiEr2xsYMIoZuHkIq2ce
HRJ9pJU2K5yjOoHXIKD6nhXyrSlW7O1w4z2XUZQEA0TBMHhNSz9uwhmAbf+fBZFUFC6ZNiBkdsmd
btHqAmCJPk4LpgxuNw92HlXxbqKXT+LR1Aqyf0XLNyQwjMHCv0zKFauKEaJSkBZTJR+dJh7QROfo
/+ovFcmlJfN2ltSmfuyehTF+frogwJgxe3vcMAyDM+NkxDQEMTYvM19Yr2oR7vJgGUC42MOHrOMK
zcq8mRNFso5AHmjLz12UDUCwRqjRIbPFDwu0FnG5Jof/6VwvyZ1KryFTr/PoKuF2J6/8y1lYmobR
qZxfGABKcytBr36tAYp5Erb0vJ1NwreOb3GW6MH5tsILUrbvpw6K4a+if8+TGVncD66o/GJWS7No
DKZSgMRTjwxge6xr9BwkcjjXtmGbLVNtJadyIWnN9VW77aHCWMdVcioGr6AH0M2/QpC1FYAjUa+D
wstBfbSrWKHvnLHOm18sXbG4sLgzUgMS+TLy/i8TNSgFeyUfpcNmhmXkGkWTN75Hht7teN27Lkxr
2CbCLXIlrM6MMhU9/P78nIizw1ZKDQfGCuS1XiTFeOi/cRXP/GX0t1qMF7rkJY+L3O0KJY6T39tN
CRKiT/fzqJDGEw+Q1CObesQ+mRCsMPxd8yRRTfe4HIamBt5sbGeyAYswWPME/umXwVL5pvGNHhcz
H3J1QV2JTE279yh7SHyh7p2I71baJBrD7qsCJ4V1cIbqWflqLOuD2nVRCGdgSB7rSG12sdj6eKi4
5m1S+xvqshPfR+7nqbY79CujoY2XRMg57lI5krWwI0Q4M2YwvhBeSwoE40UGvSMip20p/R8L76+Z
wlxnTd45npARAoQXBIpCUiF+Os73gy35EJ9xKU6YJSiEeAmlw9yaPeJSGh+fu0oryu56so1vho8i
tn9L3M89/yyHg9ujty35nwjqg1b8a6uzcUV698h8HQyYD8HfVBVtJTjEtJpk90xPMo9+KX1JPfVH
GvwVyb1MGURR5RcnvkhpErUVTBBkQZX6zl4CqZ0wlKg+WwyVscKZGD62+RWuHudgA00+h/pKPDKK
imxKksAim/qmk0vRvuNOV2lz21XEzN2A/AxzGzx97XbLEW3VbvytVHoQT5OM7wlhPd+bZJv1uk5t
vHgSXp2zXlKvk5sA2NZj6Hr7LcfAuLLr9L/ahnH/LjzFAFd4XQRH7EFmrDToQ8ot0/PSnNFAsraC
MspxpVC184c0QyC4eBso7HqeLyvPG4MqPeYDxCtxUwMSiwirwKeYPdcBWhY1nDNAH02ikZqzNBA9
vJey9NmtvWe9SbAZ3v468rWwuh3J55i3fLbxVl5I1Mdsed2f2Ry4OOX6KDWZXqk5NNj2fuML8azZ
LYiFlu/7T9vvhRBBlRnq6+bMAbqOcf+wJ5sKRG7RUFBX9nPVV41LXg5bIuG8eJ90VLxn/jCpMUiI
rhnbqya4GFeFJSNVw8a8NpLshSFixV+LQOkJ+M/TlBfyOSEHAFxX93aWTteeW1r4Cd2GtmDjRNVv
5KQtbme4not7YbBvoipoyM9QqS56xI92FU8ZbeI8Aq3H/hSmey16rvB2ql3AO3aVgu/QaiJZJ6QH
QTJBkwPWTrSzBqnkvVMZgwLIVVl02KBGuDabkweuuEgk0LrEV8rwnp7j8g005vvDb1mlOEA6s+rI
/MCpIvB5Vd1L7xajGpvrKOpGHWKizWJ3/X7DZrI37kAX6qOQY+HnlJlJB34egcffNP+KffZuO7Kz
f0jvDeXGaG7NETfxRby1933Yk0YUl4kqolWBFuGJj6YHCE2Ulm3KwiHt3nQL17/FxQcTEfn9Lcea
rDy9kbBlgGOXmvbfKv7rpfy3CIQOojFCJ2tv+VnqGAoTuDgJgIACbMx2ImDFotx52EzQae++rZaw
Edysk4mVwry4SGOf/it6Sq7rc0Jt8KqNG+uRJOXKI7IwdmAN49mdalD2UldVBlG7aetKal8rvKMc
xvPm/J4ilU0m50SaBq0bRAZW/uGm1OhJKMoSRabs4rSwUzBfCl291zIwKKKlL9zQpTeAWLRoGg6c
9/3FlGZ9coBQddGcIz7zfkrNkUH67TeYxRD3Zf/RROrJ37vNplHeklXfzQhIEZ9JV9LZvDkliKv9
+C0+do8QVw6xRCJYDZjhXHTjbA6/4+qabEkgl6oVhnFTQpvM05XCdbN3yyGLpKooCM+RcMgNnx85
R5x57+dWhfUn7yGdKgmLGe9j3Q4kCd17sR2Q0Z70SzjNnIfXcikvHhyLM0krjrq2sUAyjbwIBWpj
YDJRGjLtaagqTkuN8g7A9vkp6iEf7FimIIG4qLAWd+aknjd40eJvpsjZ1CCUWX8jTl5nkWp3FRDl
mb5lguOzPKwpKZ84daCoqkMPh84442rtPWdN8sL4ncSZIqUWfmvyi3x5vPTUM49n1KZZNCU4iNCz
oAtcyUff8R7ZdZ0hd+5Emln/kkJNW9LGly0XNbqG6JF8SHEQoi0YVxRmGMYwbSwOkISmT2Uekbj0
liqttDJxQxf76kvNdibUAZ9Wb9nZvqPILMtLryzct13NoncW5XbFSULF3oXuK75bLRm31hDzS3UX
3WtmpT/ze/O/9d/7p5h0EviLjmN5cg23u77eu3QcBbQ2UBPseeh7svdPGJoKtuGkL4gRU7PNr6B3
0E2MLEgx3rUMpatuvpsuyJOEUJnAkJEd3oaRiUNIPwImbU/hkbxatZ9OCF/Cqomb4+IegQSWbwcz
bii1BZrjNnNP9eYXSPnd7QXmuGbGzOb+QA/bp+KNj8RSL9skxtsGKpemxPIJPr7jLqvsfKvJ0Ehy
WuUmOwDBGQw3ZSrSJIuJ51mobtj1/9CE6xiRckmr2dmHTqTw+0M7NIfsAjmj9BmkgzFdv/1GVhDq
EAmpPIxCAICJSfrNK2hbAZOyZ/YgTGdWmzEYAdTzKpf76UFkK06Q2J6M0LFR8JSrZ1JhC1avMkz4
2LVJZ9AWSMrbubJUyJBEmBMV34GaVyzH0rXjhsXfdVB9AflqSZ4fI9CReeHr3ddIKDKZk2HWppr+
qs2gz1dnpxW9kv5Wf2HOnG85alsjyKVBhc0Pe1uj5UnlUHsqD/i76TIwbCi1405Pri8ykLXU5EIB
lwPQLW9VjTh/3biHYwdgVvmtZIoZdOgSVvVhFrnJw1b8mVdn7vLZpoPeJecPCtPgKYZz22uR7qf1
96OMhW3Ks8tEreruCoYRKKPOTamLWyCuvCBIpqKttmgiZR5vBm1juZ7L8tdtDRJ0uQdiBWzVKV9f
BvoUqe99/5Tv3J9snOVwpN6g/Ne1bds02F3/yAXAoiKz3+NrEt9htsgwaohGRQKtL16Qkckf5H5a
U04+w3w+7j0NAQmdOzK/pq24LgziwoTQch3lP44Rzi2hQ+nK48QfDBG4zOWFiJF18Or+M09Hbf9G
HkIcgiSZCICV85VCGZXpQOcd8iqtN3OD5YUn9Bk/s81N46jvE/saGk/trt4uPQNn/d5saJHY30P9
hL0kamtc/P+61ZBO5/Ut38k0IX4AzizFgdfvijn3vSgdxwPlqCmN0jl8GQeyX2puv/tts4pI8+6C
QQc+u56aFNbXIkru/xyPNS9le0/GuK4gDa+odDCkBoTsSb2zQMvyuOJFvjoCqfg/oMZYa03ety+W
wQ+e7hoaLa+aoih4gM6VcIdPpB5aNjrgYPOkb28+RHJfIA4nQ4aNeggh+26KLT1GrOURJUA+fLA3
9y74nzwOJZqcpQp6yhja4fvkUI/zo8wCTINZNEU7n5qMvJMYgE1NWujpfNI5IvOu/v9h0Ba0L4Sm
Npr8LyLHrs8fL8msp39q+3DrsR+MKT0dsbt+uHQz+EOPE43ZEg+8//J2qndfQ8Z7stk8kxNAHZfC
u9IoIXsxWOq5qcnJXYrDWoqyy+Yyil8lVT/LStTufRgoADUnzs5c2/kAUmTcJBUrSMt3IOsrp4gd
5apiIGqCUBuvsaAxehGFDDnSLah7CTpN4Ge9tmrMwXFIMi3NmOF8uc9L9dit2mWjFTQB1r/+cNMn
TaJYa2gQz2Gvhj3hz2zsUSyG2Vd/mCj5Q45Xw8siB228dyzJS0bUlRLiGvcLJdDRg4dHPJWjQaCf
QK6yf6qCTkknkT6Bb6Uwy89CGeYa7/xJ1icLR4C2YFWkr1SuYmMDdMFnE5j7jpR7u8X9gTDYRVLX
fKxgOA3SUuuLwn536FKbjl3TG5PoAnt5fINRWw0NViK4mEZdmbTp/NU1attzxhqrdAwLvC3FBD/l
FzdO0MXMxb9spowAdYvwMUUlNFT5pakyTEwMMicDUXRqTRo4mJx4kDPqnS1U02Mh5tx5hrIN2+MI
fPkDU73NS9hlEfw90E/GXnI5jLztvB/xdgtD42LtjJ/CJxbp8xSzeayM3WeWJhmhpM4uHot8njcx
g0O8qRgmD/lcLMwl2ZX4AM+ACfS1iksd/9nwvywG8DEeWoexgQnTrMjmbnSUDD+vYwVrinkClsJv
V0Xpdhxo6x31TRMbkBkjR7y1vhQzB1mgrW/jWocBF17USiWZPwILj2gFHs4v2hLCNd2qVkvimKPB
+on4we+99QsP1vGcCouqa0HsX4iI3D37/suFTLyuIybjdxF1lzInqLpnpZC1XOUyjVKMDrL3Qd0L
Ly8qNTTLellQ6a/IeqE9HjhuQi1wQTDSO+LI85lf1TbfCPKySYfqEwAInqJ/sGPG4IVNMO487TnK
e8UUXzXVEpPUPj93dEosdWUFltDdzViyoCigRlm4a5rcnWypKxgNsjvWq3DTBZC+jfSQf60HE0Md
BXtnG5oL9le8DZ3A9kqj0bUWRWvkJBK3ZtE+HOQpWxwdp5HV7Anfm+/6lh6IaEQRIz7Narn7MGLg
pwVb7t7dynHFgNSeYnynZRYKiWi4enKzZ49ZXBKXwfaJju/BAQywSynKHvlZagSd6NJblDPxa5Lz
/R46cS6AhO12iAplvMlbdgZWhNpD/B5iQdUxseczIm0RnOpl3iBWU47mmv1gZHGdrtqTimf7EP7S
/kjAfn7Uqj3vufUPSoVCo3BuqrCUhKZuzJThwLCq1mYeG/2zhLDuiJPxFzpxaLbdJ6nXzQeDLlGt
48X42ar7l3BwEbH82aP474B1eKXWcF3eIPlvmX1B9rb49RvQjQKSGaTLaxGQAzl8mj1SyChlkEA6
AhQ0PkWyryXXGN+Tu8ai2mi/n5w4nuMFD/Xrs3uxjLbFrSYZhfLOKc3+sh6MkokxadYHIDki9Upy
nllyqwcX7x65rlYKScYaqyC82VQf0+/+T7zol4t/V/E80l8NWMeZTqzI2+G8zznioXEtGSyIGFa6
lsKs1OtKA2WeUy/aLMoCGVHms/xKoGmWK+OZeqQxIkaMRiU/4DDWbHFqLVGwwG5mit4FQNMzljyG
uEG/MR5CryA+bV0KuysAa8gX/Lyo0QTA1DyUxWFgtf0mar4dYgywj9jROT1QYGfr9twPYfPGQJKR
1VOqSyF5Aryc9oRXR0FNGe4m/VAhAc3nGXxbEL81KToA2Z28Bo3GFdkxcJZLU+9RNhyyfAaQftdf
kpPLibwXtqbqIdb1UYYzEPgAiMyi80TrI/VxmBYCed0uOv9NxaIzpYHPwXqjmV7TX5WTkzojTuDc
bwVQ/w8uxjS977k8FiDNGMMAkvORfDEM41WbUySCMTnhAbIo+bOIM6HxlamxQoEova4BOBOFH9d8
Lv0j/4lBSIrgTUg2wSkCUsp4mECSaLwkychVzn7rdgDVor9jcg6zKQeOMirVJ690rgS+REXU92mV
p7H4t03XY4eWoJHd6DUWd3AjeJUvfaiH6GrPAXj/YyoKJIBznnefCueuJ+JALZxZOp0pNEy8G/Bp
wkODGJMMFCsbHsuZpi2P5qXhotbvTt3Ect/WL38I92bGHOvwfngpk0xrRu/XQvXoiN21bWR9L4MU
29TP1f5hcEtyYaRycItn9WNY9Sb/MTpFPF3IpxP9eNTABneBEKhvuniQxfSNJEh/VJAnnouPNcgG
gyoae95JL1fAtEA32YqqyXCWf9KvUwsYYCJ+dTsG6IoCrNauLw6IYgJNBuFwdJOWNJaZyM9KLuRE
ZVaQ8DXRNIZ4j7IRcpDn71EzPmlR26+3B7gWnnEsksy0EzLFWO+IzdiNkQr75ZzxKaPeHE57DEXV
Ppmw+HQwj7V+AZVABV2rdMiXlmgNi4Si3ryVzeWXz+KRSzoV2ooGYRCDFqsjUMBLw9oyvLIEbLF5
EKmLriFDDIkIt/8yMj8SOY/h8WvEHfDdXjXzv/zsEzlZ7GqrdngpG+d/ADk+AUymTLz/Uzb77zNM
DUDmTxGTv9fsqKxRFh36NK4SIaKvi5cIXUx9cqFZZeWeix3qCOM7MKC7rboNd5Vp7yl+6hJNZIAj
nTsxCmJWH7cSgYSdOLBXWH1PddbU/EEnHRDIzCiH0Mg3Z7yQevfWhj+1O39Hx7x8zAqAardQGtld
gjbhht56k3ZUG2/F83IcU/tzZ/T94kJuJ2oIsWR8ASmD3O8o/U/spZ+CjX2jvKNXOH1M8RkrVuzI
ALcbF1TnobFn4SzWJwBYxsLor4KyjmukhfHQxL6iWGDsr0gTWdfu13l04pSkhHDEb/1+ZLZ7uSgH
Bwti7SIpb9cuLXDoUlvMTPinhjCDQpj07JCO8z7hFxFZl4R5QuTHGXEZ7+cpDnGYpl98chkcb8zh
YOWzfJtphrIp24otC5sOo2kEZJP+HmqdOKTiakLXLRNtcBf4wUFJrWcR651UR1olQxMxZGjQBHtF
eLUWR6Uboc3qNWFVCg4l2IQl/uZGzBL4BlZMqxmiOd+l/pRlytI7KyzgRnlrD90W+Ue5tEhahRZo
NnHng7H4o4jz8/wL45ut8azJDYSj/2W5CwR3v2D2yYSAt9Sg3z/XK9KEOZd+5aL1POGkNaLGxO2X
10c637DaV//pwoLY5m/OP/wLJNcORTCeieizcNF0au5YUYCA3AySFvEaz8z1sx2VOER5focihE8Q
QDbVOKeVnmxW0Rrd9HnBXqGmUur3A600NSBjXGRyHdvgAFEf0WFrVeBqdzemrNbwynt1eiTsGZlw
Igv0y4q71OTiCCBoNg0A9R0mVIXlrTWy23xqmMITo4WRFCG1wExmZJKtdiywSb3KkMliDeOPo0+8
Tj0iMdVws+gZI5svep8goyF9KfvexqDpX3PVx/CvUTtDGs194wiuUTzULVXZlLXQbaIsqpzGA6ac
D7S75E8w6esg+QkQmLxTLPJjeK4cG5GHQWMcPOvUCwcqgQqZKdvU7uDkONlGJL4BzcHO4767/ree
mkzrZ8FoJ1USwphux3X/PS7S7b3015rcsqqXAOd9arVokYZ9Jt3ZBBjj361ecaaLAm54AcNuKE15
KVtoVyCQirZ3aHepf+PQ7nlZ/fMTCS0RS6qIF0FubZfStZsIrEpSQAnDpy/9HCEz6KuxMr71jYT1
eLlouwYGPyHNysSi+iGuHC43jwr5frXuu3CCoY9sbF/oV6ShvPfb7RnT5oqPKcovZlQs39FnZYuJ
zPZk5rxxBW16z7CqoBNAig9gZQP9fgBxh8TQarlrU+/vsoo7OSHhqyQIraFp
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y-=^��l�y�x���(� �c���Y:�y_�H����@�	�D��Gs�i�{�i{�Ur�ʘh^���63^'?�Ϭ���� d�9�u���&������Q�{�Ox�Vpk켐�im��W=V]B�\�h��r:�x"	�_Yc:��l^�#%������ETn��tH�9�>����! خz����S[($Ѽ|@Cv:�Q�õ�O67g���yJ�����%��lj�by_�����߭7���һj������3N�<r�\`bL9b��À5'T�����gƔE�Q[�d��f��b"50K_��n`��C��
��<)U�.GF��̓���Ǯ�Km*���Y�!#U}�McⷬK�a�
ÅaW���	��T\�Z�ȵg�3Q����ã�@���A��u�����F����7b	��x���pÏ��W�f���NJ�	��v�����! ��d7�~����U����/��DQ��@I<m���������b1�E뀴�i��l�X�����L���I&��q��w/#��	}�v|��{80���ϼ҂��?�b�}ʋ:��@9tR;/��(��B����H?EJ4�˶�����|?9rP�"sv;��P35��\���9�/?H�`b#3��Mܧ^Y������E�u1���Eҕ�u՛a� ɼ������O(��U:-M�߫g�®�(����Z���m�J�<�D��JNLc~�0-�`yw(� �W����_G��I�!R��+e�=:��ID��:����iO$R�@Ԓ��^��t|�~F6�DS�:��騊�Nr;6�+[�
��Rxs�p&UJtz��H����ek�zf2I3�ޭ�F�z䭎���(��Ot����ҕ�u�@Bx�څL��	�) j�2ª��M��P+�JaT�av��Ī���)�oQ�Q���P�i�+M�B�-FfRE�@K�e�C�cY�)M��a����}�^������:��Z���pT�h��f�"� ��*�Ʌ�[E�����&�Fd?�9ի>0�>"�(��}��b�$	<�m.�ى,l�Cܗq�{��)>ל��j��!I���&�}�����WU�@Dx(��������t����VP�8�,�VK��x�����'��Y�]�/c�����;Jj�FX��%˚t���n���y����/�
��:����FQ���N�y�0H�̺�Ku�;�+��IHb��ȁ2
�%�w6��x 2�NM6D�dS��7�S[�����^@�;{�s�
�K���c{bZ��x�~�Y�y�Ɲ`��{I��οy���(����7V��lٮϗ� [7��>搣,�6.o�!�HG�x4�Mgv�;��U��{��r|Pξش�C��7�5z��q�&2i�h�G��r����6�PR@��A,��5���}y�Ou�v8zr~	Ԍ�����}dw�P�[G� G+Tpz�n͊��2%Z��	Ԥ�o�� �E���ڊɷW�Ǭݒ���Ȯ_@<6��E�ZCS~���ɳ��Ȁw"H�G�e�2Ysf����DB�I����B�� �X/�=VT9&���?S`2Tw��g��*�XÐX@�%}��{|.��\��)π�T�A��qT}Y_�Zx;b�����]��bu>:���k"�DOT�{��i��pm��_��}�ψ}��7��t*������C�@�kv3w��0}����(_gD[��l	>:��{\!l�4C�Q�LK��t#�QV/s5(���0,�ă�Qt���{e���o�>9��@-�R��y|�a�fR���0�[���)���	8n��/�yA5K�&�)�	�sy��͇������T�nM��;����¹�
���eW��{�6�%ǜ��%R~�F�Ȉt;N0�h˩�K�UN���}�t'�O"٢M<G���=�jR(T�w�p{:	���
\��~��e*$��d�$Hυq������;Ŀ%"ʨܖWM.��Y��Z��5Jv������O�F���'tV5f;����;VP]t7.��O�F`���T ���`-�ӟq�����/{Q��E��^��SX0�� 
v��C�:"��J��k�4�������~�7k��&���h�:a�k� �,�w�E��啳����u=�{�=��'"N��]�����O�^ߖ��~�n��֩�e:Źq��2
�]��I�.�2!�YZ�wĳl��*�%�J���c-��01�3"*Tx�R��R���@\[VlQ���3):�	���K�ʸ���&�`Rˑ��P���(�pu�3��R��lW] =Q��⽮��s�ٺ���9�ߤ4b�Z0Wg%�3`]��dd�B�KCn㢔`�V���愧g{*�!6z�/d�y<��I��Ͱ'ì�W��j�碠��_�C�17Y�P��`\���6(���0s�4�u�=�:x@<�?�Zx�'B������?T�Q�t��9��|��-�RW8�E�����ɱ+ԟ����7��պ�/rcYB���_8B�Z���p�^;۴�ܿV�<�PL�Ig�x����,�em�
�n���Į	>����`���6*��J�:`���H�hy���⭍��&�/I�i�vG��L"���y.T�#r���l�$A/���	Iv����5����c`�}SfA*�펃�b-�D5� &��.��A	?��F$	)Rq3D5f��^˜�hl�O�$�����+�lHy����e�:`Y��f[��Q���HK���?�*�[˒�U�`^�аh�#���+7 ��\d�R�L&7��(cݛ�WX���D�g����@T88���ΚȀ�� &�IۺesV��ޮ �����������~������0)�um�*(�<�L�`a�R��Ƒ^}��5�}����-3.����'����*��y=%��<B�0����J�Zc tU�Fs �"} mL��Q߉[zH�ǿ��Z�o��1��ƃo�Qm?�e��?"j�����jɔ3�^#� `D�~d`�D�E��.i�9�i�*=z�f�D)����H�sJ�r�GHi��ur��V��R[O+��]0�<�ؖR��>�y,�7�-�� q�}�җOlx&�m��$\��vnَ�8m�ԫZ�j�ݽS��]l��<=��r��)�����dL?��,����f8�pb&�@ �f[  �1+���u&Id�vӑ%�2��b�޻�{z��+���V�MŁJ�ҳR�	sL!3��6ǉ�X�>�w��������R&׸Ŋ.UzT�^�|�U�Νk=
��4�����~<�@�4��a���+�\��fg��L���)W�� 6���4ް�����xe���F�4n�)l{�-޵U���A�,�]�l��'�����x��<�Y�f�U�c2%����B?��(-U@�'ԙK����#�<�ūpܾ �#p��NV1�ujG���j��o������0��>���F�oOv��\�E����׈1o��m焦M����4�9�afٵ�!�=��|�|EJ �M�Q�l��_&��������п���_a���^fO����W�����V�*NkC�,m$�
�[�rx'ɂ.���v��у3燻���3pc�to��h%���f���*׹1O<�~@�k�3UQ��i�"J�����`k�6��#����L��t��.����	���x>��ۓ��%;u��I=v�HK��9�t���r+G�m7�W�,g?zk�w1Y�!%�p�Q�����zzD�<��wN�F�� ևgt�]^����������,e�-�f�Eh�L��"������
x�C3��'<5�����(v�oV{����S��*������ϙU-�I���wc�W�t�E��(% ۱�i��"����'G[��/�\c
PW���'<��Y޲����lH���}�oޚ�3qF�صGy_���%/����RS��Uk�	�dk��j�����DI{�a) ��#���{��e~H�V��P~s4�Q|t��l�r=�X'Li�0y���^T��¡4�%�/OQ�:���S�� ���O��-4���n�ϻc�£��[	�o�U��I�����(Ը�]�eD.��� �!�"U�}�2|���6�{8�k��W:r 4ǧ����U\�q6���n̉1�ޛ�t��pR-�ٶ�Z�c��U� yv��P��׬�J/6is�ϭ����&�OD��J�%�8�+V+�HQ��2$o���f�)ꦝ�K0a��B��-_E?�] �b��B�Zm�,��bUL�(/mlZܽ�b�(W~ ��?������&����0NH�Pۈ.�H<3���7K�o�*Y�f`~g\։gH�3��{G�  ���3�IAR���;�v���V�ǣe�?����f\�Y��6p~f������&>d�)z����vU~I�6��OT��h8��_����|C��t�L�hA�����H@��1�\Nd��[-k!~)E�*�_�*���r��I�hÐ��b���N��/e��e��-m�K�+��ő3c���ѡ#����(�Ҧ ����r&Eav� �C�lP
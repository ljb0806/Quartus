��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��$��~n�{��ICw��"��@T���f#��a	5F���8a ?����Q����(���o��o ������e������G�����Y7��Op(/~��+���䏫
�T�IV/��}��z\8��3C���^軑q�K}C������a������QS q���he���۞	�J�ē��J-g�av6m\�b!��d�!Ax�3��Z6L���ϑq7���@#�I��C�����[ik͜s6`a�Bƶ��@v$�8�����>�2����l��.�/�p)�/��`��-�g	�cA0�!:�K��~�ݵ���� r�&[�;��'Ǽ�]��GɎ��u+�ܤ!����. $1.��`3���7\U�!7�S����%�tB�i�<���T��&/�'���h<��s�l6�BvM 1-�t�gh�(V����»���7�iˈ���@W �1�um�~�]c��������%t����2�-��=-Ft��c���;��w���y��
�X�櫮u��	���W[��}[{ghJ���8�m�V
�O/'�oO�1��M!�"��;~�%{���6��A]�؈��}��D�>rE	�B]Y�����Hp�Y!
���`����p�2�o
W}#9<����������8r�wI�ւ��LI��#�hȗ[�_�J�?��}�#�@�-���Y �`*�����o��d�T�P����m	�(�Dv���E�d�V�$�.��A��w������f����>L�����>�q׷�M��������IH����<�c�n����EԠ�7���tr�h�8�l9�m%�ڐ����UQ���o7�Q(���2S0��&o�1*X����Ϟ�E$*��;�u�I:?��Ö\6a�0���h�|ֻ;󏝗=\�';Q���.*�װ��q�s��ŃⅽϦ�c�&��CCC/��p8����i\�?rN�+戩�Ϋ��3�u;�N�]'$��%Q�ّ��0�$g��U��j��L╂z���-5�O����t~��V,�Ui�B7W��e@��)"4�J�����Yw��)t�8���i[lf��A-;{=�gF���*3!����6�Fc/\P����U���h�u�p�&��2����(SG�������:��;��1�s��$��ȣ��@Ȗ2���7�sx]?�,A�5lF��o�����ѕ#���G��漵�3$M�����q�������&|#"?V�2�3C]2�u��^Q�l�jX�ӼI?�ɷd0�� <�m�oaS���c#�m�W�Yn�y
A��<�Vz�{���IH0:g��j wo�� a��b���]�㉒�~��"��A,��}�T��$sr�H��tPҖ���GS�"V�M����;����Y�Z��6\�&�
��o�E"�7�6Η�o�L)+�x.�ى
搱�1���i��+	3E�k�0'��jf��Nx��F�mg�״�굄�{_�����JG�f.\;�����0h�����V���gx���J�
ޙ/��g+Z[��c�����Uw-:G$L2��?Q�'YP�+L@�3�F�k��B��5��	3��׎�T�<��~�ߴ�wMkTd
*��$i,f�t�	�˥:�e~y�h+���J�bC�qv��=Lp=zj�`�DT�|��gFOR.�\˰��GB���n�^�8x���ݜ��WL��l��(�0`v[���P��o�̾ H��͔ؒ!�Y2;c�9~X�k��^�\
{+�l4��Z���l9�>c��k�S7���R�[@+�ov�����Z`��r�9��\�C#��0�c{О���4Z��zlW�����ɸ �.A�fQ��4dq��a���Rl��R�ZRB��<�&fu�v��(.A�S��$slX�����J�<��R����fPxP�Rxe?Px,�sS6�V�7���ty�x�{A�g�?7%v0�	���W�U�{��f�b*!��(�^��.�oO7�fp��I��f�J��/e�OtLb��!�G��3�|�)7%�"Q�F�H��c�n��yR��JM���$�D�U�uJ[��w�����Db��D˔n+*�Ҹm��L"��P	��gI��'���8��?.[� �:1mM]<<%�������yS���]�����M�OL����{�@�h��bij0w
 9��5ߣ��qp�c^�H�H-��&�q�rߵ����2H1z�7�ƭ�q�"��O�.p4<��� ɉ39J1Z�&���mOi��Xۼ�g�K����^�V�����:���9��j]-S�%��n�j��?��8���2�@�ރ��JM����`J��`H#�G\� ���4ճ��vh��HT,{�2�EJ���qh�2DS�_��V�R/d�ۂ ������̑P�����Qt֑R���UP�8�l�>қѭZ�2�����`90�����T-�Kr�A#�%�g@�0�X��կ����3�/�?�M�.*�Rn���B�����/�|'2e�젬p��B�DC�=����YPf,E)�;�P�����fO��}�?n�7;��
a��AMѶ� ��t�e�úیTv��v_>����q�d�r>�}�2W�+��z���O�� ϴ�s]�U� aW��᲏��@ҍ�L%��M	q�D[��Vj��o�N�q�\N�Z�!��+�Z������vM6�K��]d�9ݴ��?F������"��z.6R�KE��v9��K82��N'q}Q�V��w{{dLm��[}k��!�����7�K�^P��5i��ė��9<Kͩ�p�=����N͊�ِ�b�Q�1y�G�5��O��ˑ(��s��Ui�Cu�dю�]�����<(��%�2��ҎV|��2�'��@nP��3|9�_�I���? c�n���w�@@������9���<<����>ƛк�K�<�I@j6����KK}ӑ����ZCCp��ۊs&L7����r��>*���Ŷ���Tڃ�eTD����P����czf}󜐪���b��\��_�{9�g�k��{'�ɐ��E~� �0���Q���q,��!��٦����X�q#��X:}��s�%��L���S�o6�ꌶ7��X�$�tq���~^��eH>pR.2�ʈ#3L3�􈽣�ox�j�:�V���%^�����FO[^��P}�� �$��8b�쌐��D���:����ioJY���H�kB��0�Q���3��]�����l��H��߽,��شy��������W��T �j<g[#T��N��C��ޜ6��\�sg�/e���{����'���<p'�e0�&�$�at�gR��H" �N�_�إ�m����j�9Ο����])I�ދ�U�4�8D����h�`3O� ��X�6OK8��u�W)�#-�w�	���NH�/%��zΦ� ���jd��i6{Ƭ
Q��F�����&�Y��3EQ��qt�̘��gU��ז��%&����"�ކc���=�[��b^�Uzg����Nw�N�Y<�U)Y)�����]�/�A?��Yj���h���9S
Kf�6���`������i8�W��s�y`��e��j��^|X����Jh���β۰eli�����C<�6���A��'��k k�*�X��Y9�64��q�H�0#���v��m_�W���Pd���_P�Im�U�J�RB��$��F΁�q��Z�(�()�r���ԕW�^QƣPn�g8Zabm/�	����n����u��-��n�ޮFz@��ٟ��D��|�tgd�<)�Ob�Z�F�������soNC�Xr��0NS'�"ʁo67������e�M\m�%b��rH��}#�$4�I�g�'=#<�Y$E:�[=A�"�]�t����+��	����:�H������0A���T�Ѹ��!����Ȓ����q)���Mʗ���!	���}�x�0V舭�@���']�rmIk9Q2�z�څ/+�2U�R�Y���د�]`g+Y��G�؛|&�F#�f���.:4/�>��#��,Q���ZP������z��8�6`h���%�����8�b:㭱M5�|X銉�D��`�f)�(&?B�ŕP���,�՟��:N�(4�J����{l���ـ�Wf��������~�]r�xo�{h�Q4g".�M�����۶B�H	�øO���:�q%1N�RW���e!H�N�E+�
�8����ܓVRu��H~ܼ�TJ�y���wwE4� ����s�isa�}�~��$pXP�`	:2Ak�sK�m&V��l?,]�Z��U Xמ�l�D�1� A��J�;0̚��q	 �W���$�5?�@~�K5�����t��z[�x(̀�M��.p'uV�U{�{���j�~��yY��51�T����զ\[���k�2�l���QW�٪
���4��sT��E�P���&�,a��M�V�����9�S$v�o��(H�����&���J��6��z�����B���&�Ҵ%h���E�N08�d�'H�I��~1^s�i1��0��Q�$XqCV���1AY/��^�b�2�A�$(�zy�_�3=�G�֢}����ɹ ��W]�sðWY��U퍠P���n��1��}�P���t�"ُ|㟷͝�ܹ�r]Y�
���Z�����n�X$G=�����B��WA��}�����Y�>zV��y=O��$�*~����?��4�9(��h�@!9�����-��|$�n��Ʈ����@ɺ�"ѿ����a�i����]��5CU]�T-��?!�Kd�^��-�",dƅ����r�ѧ"Ǿ(����l�d�(����[�89�M��l� Nm��MO�O@�{p4�}f��&�V�O�e���J�"�Tv����F�Y�	N�^uD���Gh��~9�MHA��\����W�g��9�|����^�&]�;��[�bw2aZ��æ!���ژV�Q���wo���vѓ�!8t_���jY�Y�8�il��bI̧��?Iɚl��B�4�I��_|Fii��e�6�7����*�BVgS���o��;����֊�h�WbV�Ҏ~��W�x�Q%�"E��21�ӎ�K�&���i�r�1�����/����"���A�P��l��>w�J@ݰ^�7�l�ta���l�������A�&�������1����+	p8��nǡ��ȧ�ei��/g�0ɰ�P4.hC.����kK���ȿ��З���n��2 ����fn��]%x#4{���1����`�66���.�|�
��>|5�K����+�LG,ZOVq�^���FC��M6�g��.�Eڲ-���f�D1��3��X>���h���]qJ�� ��sqٙ�Q�Q}��|�7� �)�L�T�s������2��f�)v!��28�_���/���2ɔY{=O,���1�V)�Ȝ$6��yp���g�CTK0}0���TPz�����q);�Q���ga�腽�(&"Eyt����1M�n3��1{ q�=p
��=r-�v\^��x��S�N_F|�����遛���:�xUtx���47�ۄ010Λx��+e��Kx�I�[��� D�:[G�[�_�;e&��A��L��c#�"��@���zbR��Й�z�����Ρp2��0�cW�t^�U�|k�5��J���G=�q�r�0gxi����$�Yh)O�|�����qx'��(��zDϢ�G�ì/�C��/�V��RJ%��,ո!q��W�s��l��t6��~�,�)��H���+���2�wn{��X�fR��W�����݇�Z1���}.�!�c�'��!a8GZ(��J�����c~^E����w��R_��>jۀ+��l�o����׫J�KG�꧅D8�@m<T��=�)�v�r�:�$dFސ�m�]�7��x��`�Z�e�n���nny�G�����Q�}��b6=dҿ%�0F�ʅ���pZ��ѣp4��^������<�!ީ��y���Gk&����usC_�{j���{C�� ���4bcr�8���,�k�+$�C�"����⑂yǶ�*f.�Iq��S\k]�A �	���{�G��8��j6��i8KD=�)����DW��@�gٺ���vI�����1θ��q��e�'�����a`""
��5
:���W3��۴�DB�M�Fd4�S�[���������	��������j���K)B�ʬ��)eaA�՘4�qm2Hq�X�r�<�<��΂��}1��ی�9b��=�K	��Qb�s�TC>0Z�����)I��������i�U���l����}�.�SL���z6�����=<.xE����3h@���>�4jNC��XD�H;i(w)���H516��"���������Ik��5�a0�X��pYY�"��Gb����M�:��L�����C.�iG)���Ĵk���9�գs�;���>�]��M"Ҳ�V���'ϖ�$_��mm��T���Wء%�ݶv��r�nB����;`��ҏ�FԤ��G�ga5Ρ1$M�"۾�l��a��Sn��q*��a�L��9\w.ɧȢH��΢*�q�����e�}�L�ⷵa�3�2�
��E:����Ğ�vW߈X�J8�iM(�K�#��`2�4��Q-N�Ë����cOE%MZ��L�N��M3�1���J�t�ͱ�\�ӫ������{��s���f�R�����AY3J���@�ށ��*�(,4�z�böu^�`�R;"�/S&�&ii�0;j�.�u�Q%ݡR�� ��!��3�@�>�qȫ���]��M��E��2�K�3�'+j�/��ե��Z"�%��(i[k@�('澆u�T4���6HĿ�	1���]q��)�U�n�C'���b7����2��X��pɃ���3o<�2NX9�[\�⹃��~�c#�V̊�f��v����`
�p��[��t�#��}_ɐ-wH��"��Ӿ��"4�*8� [�`�V�4`.M.�K{���_��v�1.�d7��M.ß�"�D�:J���|Y���6-3(���R֕	�mH=Hv���|��m �Τt�Kaih���25!G�~�/�({�%�o�S�z����" �"��zdS&/���\݇�![/�_gT�C
_��zZb���II;�R�t�5����J�P�,��2�9�.�@�Db�h�-�
SA���2���#��%��*m$��o��my����,3U�[�b��M(x�+0�DP���l�^
	�O��m��o<�[��IĽL���S[�p����^��E%�%lbs����U��`�G���!Z�����q�ϵ�A�g�1tT�Tzu�����p���i.J���gAX=��)��[�"N�� ����06�|_Z�f�u�����Z~)�Nb/�/��Wq��?w��^Z^1u�VǵIF��I��c��&�֭>�{"��k�V�<ɐ�8���L�K"<4KvO�t�?p,��&�y���S���q�û����4�Y_�e�M`\ �����08#%Ԍ�Cam��5 .n�
7�3�-|��"�� ���	��ml� j& <�K�x��c)�G�[�p�4�F��J��z��S�y�()6�G�'��ʈC�c�)V�8��E����]�o�o�T��^f�3[fi{�P�؝��$i���V02�L���rKk�v�ߐ|j�´֧B8y��>�K��n��4�T�o����a�e�o�'R�(��H����j
��SE0����q��8���+(N
 X�r���Z�s�Π
����h�o+��C�HM�V!z�z�� �ӫ$�-����Q�I�[����R}:1}�Y9�;�2{V+��'�y�x�K,��ː2��Q��+�uZU\� 5M֭�R��Tt6c!��C�YL���Ŧ��NUȍCT�?���lI��y���ᑌ�H�T����߅��ɓ�S����Y`��J
���3�4��Z1���m��;+��yY^����N�cs�>�7axm�{�@�D�>��]k�6�"L[0{)�hC���@��-;� $�׿�q �4JG��l?w��A��7FH��o�L�`� R~0c�)u��A�_����PWud�#�`��Op|Ԝ�����8�B	�JR��ѧ{�$RK���}Q�~���m�Z_(��A��V�$*��2�A2/�4X�c�Z�y�}���������k��?�����}���>����8�fY��B�z)j�1bp�7��uK Zp��7���[7 補��i�#0>���-�#h�ޭ9=����JǨ��GIw)�d�<�U-V8R�+��:��9G1t�C�<���v�����H�੯"���"ݪ�Y���n�T�q�D���f_��^�'G�C>�	�'�N5�o�E�x`��d�I���<4�Ǥ�Dk�v�rQ���Dl��U��ړb��Px[L����/�\ P.C������V�"�eQ)2��=ޗ�倗�z�j��t����'{��H��'���i9���Ɩ��N��tB�n�@�Oqۆ7����c��mH���վ��fԈoj��J-��8:�������ԁlJ�E2с#���^������!�Y�m)�ɭ��K���fX��1i��l����Ѱ_�] ����J��H���5��s<xɦ����Żt�@��,�sH�I�My�u�Ю�׮o�x֒	s��Z|�Mѡ}M➨�Nl��d'=��y�힖v��O#�/�v�-ނi`²�~fe���B9I�d����y��I6 �,@%�$gF���S6L������t�� ��K�➁g=L����K8[���՛?�|���/�Q{��	�Z���+r��l��	��)�� ��M{�o�X�v������"8�̫MCEl�����6�5⹪[���$�`�1Xc�Y�-ՉT�O&�c��
h �L��(OY1|���&P$|��A��gG�&D��x�8W�ay++0�����,�w�em�0����k?>.ͤvJ.Kt6 ���AJq8., $��#u_����D����\�u���b�P��B�hC�D��hx��Jū�Ⳝ�ȕt^���_���$��-��Շ�MH�m�ݸEW�uwۄZ>�yZ���T�{oy`
��,^�N���%0�3<�b$��s�̮���`lr.�b�t[t��֚���<�||	S���mp5���]��K�e$�Nu��<b���tp��4[��Q�tI�.n��"������LË�Br�9��/YB�J�Bv�/��4�ka��%��4��Ԁ�4�gBGI6�K��6%˅_���xˌxb�;x�	�V��|jif���z)L��ś=�և�#j��*�Y��Hgs-�;<��M=��k�8���@��F6�y�԰~ht���c��&��d}�n��|���]��x���u��-��v�5���r�
1L��������7W��13��/�l��k��t񔃱�s��X��oϼ�1Y,@g�|n����+U���vq�x�X��|	�C�]t�Xi�w@ӿ`��Uf2�ꝱ���h)�Rd�d��+е2��B��2i��*�f{������ţ�p��8��π��Y�z�h������um�O ���$ݴ����ĺS��l[�?�(�Y��{B^K�F֭[9���-|��3c���En�7+
�Q�?�ʡ�=����3����L����{�0+"��bƢZʋ�EMm������R���i��1=�X��P:����7I�V��X2_����0$�J��w���V3ITs��o%D꿣��p<�;_2�6�v��%�lz��h�E�i@�T�
<UK7�s�U8��9#*�O�v�?��F�6��x�S��˶i��~�T�ݖ^�0��7��� P�G�}�LxEh� ;"���o��d��K�u���d��5׿TN���S`�p����e��ߜ~7:L_B#��铢�����{�8�l��c-H�U+�?J��W��RD���y�7W՛��[7��#�rN~=c���Uߠ���Re$uw�Ej�Z�B�Nly�Ͳ#���`!|IYn�4?�fw����WS��%�9�~F��?�XzXo��<�$�l�W�CB�n~X@!����s~���B��U6b>��]ݳ��iCo���#��'�	f��4S�Ԯ��o�&��V�����י���5�[x1�:�}���}L62�q�sYS���qG�W�C�c!� �1CJm�1��/����]�;��Xa����4>GE�iC���\3�=[�;��;!��m�:��y�����)�g��I�|W���L/%�Yץ�x�;�M+���(�E�։��v^�9j�hf�H�Z֡�b���m��\�yj�=�t�~���(��j�s> 4�"��h���:to����=�߀Co7�I}5�8A�a���<�fK�1k���M�����x���q�W��Ρ�(١F�-�����1)x� #����p��?�VZ����+^$���n���*�_�q���x��lG�&�-�y��������x}�v��c�{���f3�)�[��7|!	k���.}�8�=�W�"O_�[�G��t�#�����9�ќ��u;�)��\�z�����*Y9��+?�������bL�
f��(����-��w�jtCA�������Ÿ~�p/X�J��;j��KK�z8����y'�kqs�V$]���'����ƛ����.s� ɤp��`
˽_�EbO�=]bi�{f]�٭�L��h��A�T�ke'wu�!_���@tE��LI*�"rwt��'��Y��mY�C�9��X>���]I�*��]X=��|�2�[��D@/���]��5���R�ë#<���m��~�"?h�;�=�4��i�+eU��+RDw~.�*��%��-Gg���@�Ģ�}��Oxf���d8��'�UT@�(:�3���^����B�����`
%g���6�t���e����߷���@��l�� hw��2-Ϙћ���Ь��p�ulA��*���nEQU{�G��rU�",?�CQ�*i��]��]��U��Tr_7fS��(�L~�z<�d@�O��էf���U���t֬�����:!I�j
�QˠJO�j���� �o |l����w�$��l����՚����5�+:���C&�80	��E�|��4x�ކ�y˽�ZU���RrQ{q��_����� W�E��ߍ�#Q��Ӏ�ͻ�9q��M�UvNu�ZNӸUA�%� M��|Gm��{��Bz��S�QM{���<c��|&��:2"��}��p��Ws�to��H�;�ۓ��eUηe�}�c^_g��ͤѢ�J`�q�Guf��Y�r���M��o��Q�8w������&ᩲ5)!�&�6���� �*"NR��E���@���a��9�� 6HI<�_��U�5Rℵ@�rM���~�>�Y���`��}�$��(;�/�8�30�f��ݟ6��CyO�<�7N��ON\��DE�����7����.],�f��K�H@+��� �?l3� LQ���me8C�~8�dKVeci�DL[[TJG!�?�\��_����p��|��x�z�l�^g��/�%�+�r��OJ1�J�4��ڊj{�&̄��=�J������6�N 0�8��hcQԣ�t���L����oQwg
�e�xc�{�Ll�)�,��)J"c���s����?S8g[�Xm���QX�'z�v��(
�?ѓ|	�'2��.�l!�g���P�K�+]͊%������!h/��A)\m������B5lf,�B�^�=t�s�1�fw�~���>�N�FX)۵U`�����6�вI����䦱v�K���<��^í0/6LU�9x]y#!s^�˄��rG�cK�Bn��dȧ�~Rt��2[��,�lw�?�t���iF
4S�*�����aJ�7���p���XI���"W4�_�g�bK��e��5|��0(�"������&L����GG�D�����K�	�M���0�#�����|������YZ�ǺP�C�6�2a,ݒ1�����£�U��z̐Х^��h��]�6��>���;�x��I�j%�V��3��W���b)�8���Y���1�. ��U�� ��	y��`�Ӟr���R��"�,ʺ�,P���ơ�S��?A� ����İ=AaQ<*���3FDq�J�V$ �~F9HB3�g��>�sdj_N�)iHM@j˯�B���9Va$]��ܸ�\���1���i��j��0�EH�Q��?#��<���߽���=��9��xW��k�%�����Z�q�,����7 �2H�`)A�cY�g�4�p�Z�Z��(hEpl�����#�=�E�A�J����z��JKvn;�\�S���l���-"��!�6���UԠ��U�F���#��9Ӊ'D`,	������rwa�K�i��[�j�����N�ay| _���\��CU>� )���L����-���B���At>����P�b�����}c��ŉ�}��T2m���|у�*$�Ǝ�᤾������z�����I�X���J�8$�m#�q�s�� � c
f�J슮1�5�X�]�4�S�Y�7�+�>�Q��9�������K�Tv����]��2ޟ��Ə}�"1�L���u�<}a�5|��H��[�����KK�(^+��ćT��Fc������\>/���v����ZbG%�Հ��h��8�sP4�r�g��*���-BQ�"� 0����>�u��4EĽ_���RW�Zq6�s����=��Z�hr�;(q�Dxh>t��?��))�#B|ZV��r;gS̔����������C 0��^Wn�W��J���F�j���D9�<7����\I !���L�u�m�T��.!4� jYn��
�g�L�]^TM�/�E�ق�3ccd��b)�{k
���/�w��T�&%�]6��u�-ʶsۘ;"�醩v�<���܂�s�?�mO"�O14���G7���)�6��_��7A$e�3�������M����Jto���Q`6Z�t%d.�	:Ў�)�)0���&�nƂ؇ɓo��i'zaJ6/����$9"W�	w4	]?"��e�+���/]����Q��+��"me@H������� �9�WoG@���#~��Ƌ�^r0Bd�uE��YZ�3��o�[�'�R�ŉ�u��cpZz��B�/xK��Σ�z
�~���+���2����L鶮~1h��{�P�^-w zeHf�Ɉ��NΘ���iצ�-����.ˈ�=:;y, Y��������k�J��}F����W+T�"@vU�=�C�cO�Ϥ�/J2qD����+�s�m[���3~�żPOG�7F):
L�rq�8�v˥�`���f��Y�T�5�����ED��O�Ȍ�\2��9�����p�q��*޷��t�0�D}[�R�?5se��%..�@ԗ��k"7��x;���ҋӬNU�J�"7���-t�ɠ�^�>�f�ݜ_�'����(=X�y��~ݜŇ��F����'!B�DQ�!�t���[L�+�rM!^=B&�i�]��x�:�;vu�-��Ε���E`$N�"W)<�E��T�� ǔ8=�s��������|�xC*nR��p��=��LR����Kj���h�����Lx��O8F��fH�s��z� �-To��vS%���:�t��`��w'w'��]5�?���> �K֣�W�]\f�kj�c�A���S(�����1p!9�
�g�A�N�� dR(�}ynϞ���Q�^�޹�����P��H/ �֫�jF��aI����isH(Scq9�f7�9U$j\8%�ll���@�����= #H���4p�ڙ%"� +6b*È��p�6�(��^�� hk����Ɲ����gp' ���
�k]t ?��-R�=�<,Z#y�Dy8�,��^����4/8X��p>�:|��=qU/`��!R%��Yq���,�?;�(+���3d��N�B�n�Y�+���ݷ�b�G{o+��I�-n�<!v��ÈKg^�ѐK!����p0�3�e�'�>�o����u�?��agj�9Vy�
#B%Ҵ'��J�;���{{Sm�}��J�����ަ��4��qM/�4�^���~�>�d099`u���b)M�/�����'�4X�ԃ5��nM��W��/�DXy^*U�귘\�#YT�ځٺ�2����x�~��Eb|0,��喻��C|0i�p������e_�ɋ�O�Y�b��!�)��չ��5#do�g��4�N��u��]e8<�VP>F�얚��:f�	�|���M=q�Oh��Iw�$��>4�h�R����1>��L�o7*��-c�����J��I>�t�G1�9<fٸu�7<�����>J-ɺ�����d�H#~�850�kO�״����A;�����*��P�=Bt'���r"����;X�p1�o�2KX>I�D��`��6�5.0=E۴�{н�yߠ�c�@��^�nV �����>m	H9��M����1�y�j��L#��r��� M��v]�y~:�3!�^��4o>2����˽xU{��!�q������@�����vb�$���+*f���@�E�%꼫�9<j�V��>;\�4�r�J�F�T�ǽe�8��KŅޑ�L�}�B|]�*��1��)e��?��`�5��k�Bn9���m�J}Q{S�{^N��"B��!V`߾�$��?��K�\�=_ v��k��n��igI6�r15��M�N�T��DR�����<c�1��Pyd��;���u�0�3�	=HE�n��A�D��-��e��G��U�t��8}<���V���!�h�X�P�[r���ӵ��d�1�ۺ����N��x�:�*�`ka)�ȂT͡qw8L�>ޣ�M}�u�<Tn�^T%a���g�O��_!��R��jL.�X���A��9��k�ڄB��2?,���g�9C�������n��w�%��p�����N�Ÿ�W���@�-��|��\Z��F6s_���&J�v�E��hH	<�f����nvQ/��`~�Xw�Zi�չ�=7�ƋG�l}6r8�Ɖ+�r�wh�9���� �g��D`U������o�V�����,�|h�������`ŏb�]�1����DX��ct\�k�j�ǗB6�=���$�G#��'�����q��8p�|��|�zZ�	�ꇇ��ȥ|�#�����l��Z
�cgE�ʣ����&�v�n���M`��7�.��ȃE4��q�w����Iϭ�,��v�ћ�<<�p��Y!��y$ƌ!g.��v@�� J�Ɗ�V�6n��[xh��ζ�O�QM6����'���/3�1�e Z	��:��=w��*���;T;E4�?Ֆ��D���-���z�a�a/�?(�_�#8JDEc͂Lm�\b{��%H�މ2���}��F{��r��ng�^ ,�ϐ�@�s��F��Ky��V-7���_��By���O���}�r�~��e���j0��ԉ���I�̼����FNu�/�'������IL��Xz�DM�t�N���b���}�Pd?�-�T�di��� v.k{Ӎ�s2m)+:0ܫ��E�4�Ҳ�1̉v t3���$~���	�k8*R���6�=ZWQe���䚦�&��a��C�Jh@��n� R��n``A$�]�7j9,�����E���6�׵*2��>��;	�R,�"�6�	ĝ!�f#e:��W� ?��9�U&�C�l4��pWJ)��)g`J�!�9�7)5�6�%�������{���D�Is�^�M��B���
!W����J[��a�8�!���:��ăj�0��,:�������_o�����e�Uk}Ie� ~Nใ����������?b����ο��v#�sD[��Et��fF�V�?+9�9�H5���4��~��4:��0"�U� �*��_t���
� }�s{�1��(�,��ჯ۰��q��MbY���9�ԭM���R�K�6A̟�T�S^�k�$-7�'�3Z=�����Fu�Щ�U�*�~���M1k<\?K�@z�AJ��k���AF}ӵ4�L#_�����=�%�θ&�흴<�i�}U豀��B�����E�.�'�kG�/z̒�e;�\*��no�O��XsN�f�-�}*Mf��`_�	���!�!%Έ�&������x�������$�r1R�ID�{�i^rQFn�~���)�t�5ڢ�Wn ;�lBE�F��q�����	��F��b�'| szN����Q������p�C><�KTR<�|�w$�_���m���3Θ�Mۖ��;Ņ��Jp	���7S7�Sz��G#�d�m"�)����(z�jX�B3j�C��'���%i��[.�!��H���u>�(��p��ߪ��ձ֧}ҐE�\h���)�U����"~'���d�ŀ�7?���N�����������{����W	��z��0���P9)�4C4����h*�d���Lu&��w|�A�V՟R���}�<C�#��Ӷf6�E�L�ľ-oP#%����;޹1",k1��S��K�P9�R�q�cn�d�|
#�Ί�@,k�r�6���q?���λ�&t#~�R�`��6 ���6�@,`Y$pgE�,�LV��6�e��}/�S�]|="~]�����B$r���İZ������(4��l�!�4-Q�@���-�۴	¥{�&�O�{S�-�"ɢ���5�,�@�ʔ���e�� 
\+� H!�m����������MsVo�F�~�v:l�]��GK�]�!y�A��_�!��9�}�1l�@��P���iH��a��+~'ߞ�y�&8NS�n|���E���K�H��)���F@�;쟣V=���H�ӻ�+=���i�&l@�-j,��Z�9ޕ�q!c�>32������X��N���x|��D )g�CS��+a�Pb��;F���k\��e*�F�퀲��RG�f5�n�W.p?��_{!�=z�ES�̚cT����A�=����6�l�Tby ��dɩ��IJ�(�5�fl����N�/x�IQ$	Nt\*�&�" �/7��v�Xa�8W��m47~]�̙G���B����p����s;p��d�	LI�5蕚��\��[������f�9����-������X�z)�3���1Ƽ���Z����K��O���A�:;@�4�ovʞ����={�D��w�39���6�ω�9)�;W%D-��G�YSu)��*�wm�$ڴ��a�߳�����x�1FF��]K��^~E���t�
�599k<;g����3�hJ_���3�9d�U����s���8�gom�(V֓�½dW�7(K���\�GC�� M�${G<��1�h�F/Ao[
4�
J��k?O?��QV�������8���.�B�˵��g�R!�����<�>h��b�P]'��� n����3��m�OG�u#G\��� �����eK��`}>�soK0�q�+y.�dKH�f��@l�m�[	$䈐sZh�)*N�Wt��+squ�ښ�f���͓5��IV��B��-���!�]Xs��b*��wK�Sꎷ��>	0�M��������-.�U]�~}�uں6�>��D���gw')���Q-�ُ�3�������<�#I@��	ҿT�j�o!�LH�ޞd׵0v�z���NKr�%^+P^~�]dd�ض�ựjջ�2�d�"' 7�VqxS�ۥ�3�%k#+@(��nm�R��h����gW��=�k���u�����!j~�r��za��lc�m�/lxK�G�#&C�U��6�:+c43j�|�FI����%�V[�����T��]�h��l�����GU8K/5�����B��B�	m�|}�P������F��{���5�+���(N���5"ݷGFQ�.�ɺ
��RO��e�H��!�)���8 �׿Ŭ�q����󋄯�%�+!t�%@�R!��b��N��3J�eQ�e�
�ڌu��\,��&�Cop�ژ;.��e�A\��Zi��� ��d8�L!о�()	�X?�=y�̟���j��V�\Q�������r:�.;�.��_��ҦX�	�Wg�3�[Ff%�%�hD��v��,�zqF�J����F6=[R¤I:���J�وX�F/}�T3{<����o����nc1!�{0k�
J�Ԣ}�O>CQ
���{RT���
+p/�N�3L~ �` �%� ��}~K-��^%����Nc<~�77ZU���gȄ�[~U������d����JQ����]:oc�>|��3Eˤ��T;҉YPX��c���Z>��(����մ���I0ЯY�.�Ou������f�j������b�>`��q&)�����E,_й�Y	���F�~���n�rQY�D�j�%�%�IHpQ�Q����`��l�%OV��(��u������-Z[�k'�ZU3��N�5f{ӎ�$�?�H�+�,&��Հ/)�S+�B�s��ʾ��3�J�b�!ҹf��/@E%;��Ƨ�������lpy��K0[�s�՞w��q(������f�{+ʒ�D������j��k�
{w�g�=�����o��5�XqO���Z5T˫r:�S��a��Vs��m�6�{�%���~�#ݴ예%�ݎ�z�w���9���+���~������1s���I�acVL�y��J���9��C����ٞ��|����N�E�g��^��;�	MH?5L�o�2T�V�8 �3ҙm6�c����C����AP^I>�)ŽM� M�M������� ��=�t�(�~Q2~l;�z��� ��U2�j�ڛ�J�ӕ=��w�_��b1\��=|^g��-��ʌ��=�}:ps581�����'Sc<��!�7�t�ύ7)���83�ѕ���!qŦ�U�1��0Ԛ5&���鈌L����!ٷ�?{��Q�|�xZ�������@$\���d�5�b���(19I��V�ʶ�$ ��a�4�m�)�D J�;��	GI�5}!���9y�"͟����� �_���so£_;���ѐ�I1���'oL�j]n��?�Yw� �������6>��x���9+7�| �������w�&�X��ƕf� ���D�G+�~0[>(�q�[�ħ�_Tq�O_-y������Q�(̗�@$N��3��v�#`�c���G8�����zً~O%c��"<����v�,�~|��`J�)KXq��!�VZ;�g!B�_ ��P�y{*��7E�k��1,�o�W!��i�:�}x�Cۉ����x�CN���Y�����R�/P�2	5أ�ۊS��"�b=�
�B>�Ѝ;�k`u��m�G<����cW]�<��;w���t�/�5yIMwr�5`�=�<��rt�uU;K�7��6��|��y�R��
�;��M4S��!k���}����	^*�h��``�iV����v���LG�A����Ȝ�;��4{<H��>�e�V�T����Zo�a�$�*����G�;e�#0��~�R�������yJO�0^Ͼ�/c�������zE���GU�_� <Wȱ@����VyS��л$�g�IvአA��� ��"p9〭&��գ�Ee��{����r@����Wf�V�R����������$2�����#��0��9��wo*nu��?��m�xaɈ Dѩ����y��_ǤE�ǡ��Vu���,Z]�aY�Fa �$��.ҽrT�������|��_u�QG����(U1��<��2\li`V	�0]���a�b����7�}tM�&v��l�Vz<��FE��"+�F\-9J�t�z$�8�GUWՑY�B���Oy|�q�J�*��vuT����L�[�:�3�+���Q�x�V1���t�&)�O�?��Sw;evR��v�P�
���JAQ�]!q*�dD��ֶ��V��9Б��M\�(9l��9huJ���XV���}L�>�����pQ֞̗�|�53�@ߤRa��#��]W�h�}�84�Q�R:�o��[6��VEN��9)x# 0T1yϜ}���O�	��⨙W�#:�p��R�݋�#�,^E4x�>�[�	6阋�'��W*�>�K��!���A��bH�OX��hd��y���ܔQ�),��[FC����{z_����n�$��b�r*��[9�}Ub��,ǥte.�:�]�0�{LO�[,qL:]\s���V��	�D%g,=��$K�1���4��q(H��J�ī-�iX�(;;��!�4�,�3J�G��VWM�Cf��h3H�1�n:j�Y���Ϛ��G�i	:��R-HS7�������d%��0ـB.�d�\7Zra|�4du��& �5���q�g����):!����Ag4e|;�|bi��XAJn��_{�ʙ@s?����/C��%W������s:ή�{�Vo��� Lϭ*`�Z���O��Z��-y|�����fW�v�R[+!��w�}W���c�
�0�dH`�̱|f�촕mL�H�����0"g/�ڑѮ�u/"�%h塻W\Jk�-1\�֋��MDz�=��������������[� }&� �y���ہ�=��[�]$�{>>���������� 	�j�Y���xѸ���)Kɬx�@�����p�ǂ���/Q64{g
���Ǟ�16���(d-nC��F�`�g��%ӝ[�G̹�>W�����L���T��A���u���	iaf
Q�eJjD��jǦ�нGd�C�rk�_����lY��]�RE?~E�H�s[�oD�� ���n��`�Z�4$�0���3C����\hC�"�ÿ�EE�a���)m��Q�#��_�E2��}�/�]s�118;'f&9uy�}Fm6�{��k��F�!�etV&�"�e�Q81'��E����|�m�������B�;d�������a�<�}��Of�����!��;}K�2����f�)o�z�4�Er��W�P9#+��m>Ѹ ��z�vp|�qwor�3��4L�ee���#�L�Yb��G�H���k�-���
�A\��3� ���|�S�ʝ����ܿ�	xg@G>]?���S:���������(�Sz�=QrR �mo�,�	�c�4S� �����~�-럎��2�OEԻ��R�׹o;�;��sS��@�����M���au����c�3�FY����"گ2ri�z;ADb�ǳ���wȵf�7���Mj�.�|`D`Y"�b��gV_H0BAc�܍��R^uvO8��G���vG��J韧�W��j0��"��%�YJ�w���%�=�Y >I�q�O0^x�Y3&�Xa��H�CX�p�D�E�5,�Gc��P����Ve{S�2�|�/���<���T����3wG[��'ǚb�o�f��A��A6 Cr4?'W���y�J߀�:���Q�*�%c�g-���T����˜�4�xo�9�$.Z`�p�k��R15���dr8�C��=y���,p��x��W�ףٶ��ALa�N��:T�D%#S�g '�h�X(xC�x��,�[.;�Q͜��o��T����΂�D��4d�.��R~�|}�_�����UW_�ހ���C$V�A���A�T.Q��j*��!F�,��Wa"��P6;�\P����wh���������Q	�Lsf(8A���u'9{�U����"l[?Y{��,��A(V27�S�:{� ���\���ى�O�-G!��ew�qlሪ v�E	(N����ם{I�D�z���L�
$�ws�ݪ�b{�ɬ����ή�z�[4/��g��m�����>���o� f�(�ò��B�Ľ��<��i����a��٬IM�f�.�K>��dh��u]ZA^2<�ۆ�HO���+WPbx�} f��AÎ�f̢量��������#vRW��T���L�jHs#�-e>�Zc����N*o_�Ik�U�뾫~�>� �Ҧʧ�3N=��KR ����a�%���1���~'�eGu���$�΂C�"%�AԬ���>/�E`��S�Z#�1�z�"�70�(v2e.Џ��>_Լ� � �A2	M�09I F��I�36y�1�CY����3���F.�	-�B�slu*����ܕy_�g,:��M\5�RP��~^N���Ef�p7���1�������{�lD�>SnkQU.���e�?8&V��ͨ�}��W� ����FMɂ�̪b�R&ҍ�r01�e�����#m�v/�;�w@8n�Q\q���:�	�I���"�r�G��ID��O�P�$f�|�vl�K�us�v6cK+_�����Ig��^�_'�������z�l��H���wiN]��kZS�z�Y����{N�H���������
'D�/_!GY�,��ݍO���N\'�j��L�41ӱ9��%ߪ�92�����e-h#�Dnx}'TU<�n{L��"�O��V�VG��RK������ֿ����	욥�\�@��#����a���a���bCJ�īG>}�(��@�ށ��b?��G������ΰ��K� �ܿ-�yy�}F�12�=�]�9/��>��T��3�r��S^�v�Dl���E_��y��+��7�#C03̗������ٕ�8U�7�L@��S��>j�UM?�Z�^�w��.F���;��$'ZF!K��w��J5԰>�.T��[ش�]G�U�Ǫ'�;}��-�q~��TW����:��cX׃��y�/P���
�oRϠ�	�g%8�q���<v�� �W�<���C �&�˴�(P�r�z��p����Snbp���:�}�,�]��)���BĀ-��t ]�ZG/0f���j|1��m��meN�	"�_x�^��UT�D}���֕���"=E�ٻV?���q>�W-`F[�Ko�R}`�ymD���'�4���pֻ���yfE��t
�ˣ�oD "��^'�༇�KO������⛞ƭAEnhye������ڻv�j����=@�^K�ƽ?����7��a�]��}M!p�ܣ]�H�� �/G���@v�i����=5���_k��Y�!.��u�'�{�U��J �\.�4�ڒ���`V\���s|_y7�6���AwYr�7��^��ק������{yS?�xV�<�w񶕿ۅ�#Υ��^��'d��c�Χ�*�f���spKͅ����M2�	��<�`:��H�������r�}b�'�w]n�R+�6Z�� �ڭp[<���!3~������VX�vȑN+�N�-�x�3."u���xsw%���U�ac7$(ȯi�U����s���H4�;:1����ǦϻU@mi�\I��?7CS�ה�d�'�M�-���γ���̊kX�ɮ��/�������E`��Y�����v��ޤy��+�����o�K&I8��r����Mkeu�rs�O�˶�N�;���W��y�r�W��W�$ި��+�;�]5�*
�Զ�K�ۂTA˹�"��k��5����7�ÿ[b����.�7�Y.!� &/����.	����������F�q�Պ����I����w�O��YE#=Н�@�u;R�]y�P�zvWB�M[ULYx���#l/hw��K�\�Kcu.�������%��rс���&�d�3�"H����7 ���w��:VV�l���N���dk�8��Y�H������7h��4����ބ�t�>f�Ǔ&gv�nQ��v�Mg]��=�p+��QA=�q?	�����n�����+Rh�Ȧ^�2!��Չ��d����[VĄ
�_5I)=����L��ܑ���6��|GU5�RdW��$�6S�Gxo��Q&Q�_��A�Q�j����������t�_9���ꎩ�̸� �C��󽐾1�Q:��C԰O���j����D�&e����B.*:*a��엪�����C	g�xB���~�\����H���m�!����J��o�v��'ŭ�q_=_��{Ȯ�;/�.U�>�s��׽4~��Ortr�	��[=���0�չ}�����@ޤ�!)�~\�þ�(��8���Y��<�"g{�G�/DJ��kқ�:�-���'݆�l�L�בS�C#h�;y�)I��[~ц��Lu��(׾�O�%RI��F�`�VFn'�
VG`�:�h����;�!ǋq�(@�0�$�����#+Z�sN�lLxP���J>�s�)�u���A{Fv�+��*,�����b�<�� :AX j��dЧ��P�$�\9��TMԥs_�-���J�*�^+���Kb*x"����<S��>�����)8b���3K��H�Y�y���I�]n�E
��S2MUX�du:f9��Xϳ��&P�U(۶��8�&G�,5V�0[+W�vE���z?�?!�u��D��!�B^R�� �M�n{�衇���u�����e�
�	*� ��H�C4؝4<i�X_X�Yq�n��zf�#ة�SAf`�/B�榟���\`�3c�,Md�n'�Q)��̤����-�S�fa��\p�χ�*��H޿�U<66�B�-
�A�=D��#>zO`�Z9yη�;^�.�l�=���˱#H�p�I�SxwWW����ܒ��ﭼ��=Lt��&Sߑ�lk��gة�༈�(R�>�[M���;�p���E�&U|���T0̣D&�p��������a�����Aމ��qr����v�'�����i�إ�dqdk=�H!X��B	9�01�w�d����=n�k���ɗ�u!�*"��?�/�����/IJ��@v�Ș��1`_XǑfF�$?�	��qo���
�a:�a�e���Gi���vV�7!Yz�݄�������3�ܻٯ�cןn�`uU����s6*y�L;���|
+��H��sZ�������Uq���W��w.�vͲ�"5���k�*Gr���Ć�W�n��he�}��c��p����@au��.���XL��wU4����� y��η}�E<���S#�ӑ������y�L*+�ب���X�U��d&LG
����>&J�pE<�20�}�?��0��C�W"/ ��u��LSʢ�� &���[�uE��B������K;z
��V/�
i\{:�Y��)ѹ��C��8�)e3�����j9k�\���}]� ����,���� `yC�0|z����ky����b�i���(�9�~˸j��DX�"�O!{j��� /j��A���b���C����P�R �	b����Ur,�Enݤ4:���eI|�¤,��BRf�R�67���E��?e����AH�>w�I��h%�wr.�#��w�a�Uݘ�n<�Zk�mY1FT��6��4�L�ƿS�"�Sh�H��B�ۓus6Cf9�w�O��^CS��e."�j�����:q0�MY�f�1�gm��;Gkͣ�[�|*�Xa������&~"�����F�F�ٶJ��j�����LƩ�=�7��|pŠo,03M�͍d�&�<s]�r������h��mZ0n����G�֚G��� ԛ=��X6�$3��U�Ψ-��l|�r�QQ��
�lzI�ATy[�5�
���ޓ�� ���6�g��H'B3S�uL�4����D��7[ �Q����ui�%;�B�^���>jdA��;:�`R���I,�>�"\d�3�ݫ=��0m����k���������_��*�����Z�[\(��s��P��	L����'o��3-O��:��V���m���iB�%��:�6i�$�7% ����r(l�K\�� ��M5��6�*%�h���IT?ƪ��ټ�V$�J*u�N�֡
�������zyM�7~�5Dvʌ��npM��.5.w܆ocFڽbM�7��/�X�Q3��������w�JF��߭w�<#}���eދL^�AGG���k��^P�mRj���з��0g���J���?H�k"�l�����HFA<IR�j�),^�&+�;v���Bk�ÎW������;�]YfJ�Ep4Xl��x����~"yH^��H¡�mڇC���R�.E ���<��#sÌ���v��l��� ʋa&z��ά[��G
f����j��=�2��G�˽1�b�Y��m)�-뾔�����[�kd��B^L�`*�/��p	���|8=A��Ctl6�|Բ&�f[e�;Z'�(tce�r���"F}��I�Yr���kҌ�|�@�[At�od���n^H�-iGYW��ک�Z��|V��nL�/F�]d�+�YA��ϓ�E�� N�U7K�6���f�����ͤ�I휭+f�z�o�%%�y�?�RX��2M�:}��_v���jA���;���[���d"?���4|Q��3t��,/hD�0Z�
�*�2��Ds��8:픇��n�*���e�mi�6��|���(1t�Ћc�p~|,��3h���d�N�H*sY�L	+��Aͬ\?u{x��}M���J��)��2�\�W	^ $s�<�PN�
f���j���P��w:�i��u,z�{w�i3����m��5�	�A�/Gt��N<'x�'����F���xw)��3DMX>D4(�Y�A��䰐��\u ��U1[�V�����@�8I4����֖��;�����Z�f����y@%t��\�z��YEݔ����^�x*�_����iY�$g~��)(_��8�9p�
2f.�����%@L��1�S	�[7���O���BCK�\u)x�##BH/��H�aro������
����+��a��q�ɪ����E��������������
V|�����mV��)������I�~�/��������$짙� X��6: �U��U�MOFJ�$�xIJȌ�U���g����yɩ!��1����w�f�W��`��B�0Q��8���p�z�r//�h�$K���i$݌���x�x\o�jꚓB���uҘ[a��Nf߸L�EE�Yw�(ۉDYP@[��swK�J��A�=� ������_����՚�Ƃ?ڋ+!r�4�������Ȟ�ه.��Ϛ��92��V���Z˳6Ø��Z��e� �RЂU�qe�4v2h ��"���ZJ�$�6����I�ZRf�_��������L�d;�3$�_�HG���=�w��I��0PNRx���_R$��V����(���S���ŵ
�4X@�)e}�K���SƷ�\�ĿY�[���8���cD��;��ǿ��q��eJz��C<Us/��X4!��C��I�k{�W����Tj?��z��\�Y�p��[		&�|ȭ�D�;�l�b���D�z�*A�e�N�t�?����O����u�3�;iD�;D i��!+��P���ڼ�t��8�<s�B�O?֗����*��v��Bb[�	g�4���~�EQ��^"������[n�^%��G�#3���"�k`�$c���:
z�w"Ԓ��H��-����;��)Qfa������Q�y� ~��QT�B�	{ �!�/%&��UI�+wXy��ULy�%M�~Q\�p�
\����u�Q���u�;	!x�9{���b�X D絗��'g'R�=$�@6�##�Re ������Ʃ�l<$����A���o ��.�яw&F�����2�]]�tά|)5����o�A���JB�r8ĳ���Q+�/�<x�y�)��Y"����-zS�����B�N��-��@�X����z�+ks���B	��-N\�y����[����>�Ǣ I��>��XX��1?A:ts�=�[�H�O���>TA��BE���i�����������_
�9�|���_�&�NI8P�r���[1���TJi!m��N�CJ: qɣH�%�䨷���O���f�s�D�<�?��e(2JC�,��{�I�o��K�?˙����\�y@�'�UX�P���YD������gm��k�i��4�<�xۀ0O1A�}��Q�Iz%!mT����}x��n���.[�W¦G���Hp,*c1��\_ X
��H9:��b�"��^��w��yraN&܆�����e��G �8�T5@����k�[�~-c��]r� ��@b��x(��5H�	�_о�b��1Z9J�Ƀfi�[��Il��X�C�����{8��ʪLv����(,J��[h(���RP�����*P`�r˷]���36�	�]$7j��U���]�{Εz�e�X?�C��փ��0�l��I�IOjG=��<��I-r�m�z7u��#@ğ��r�㏇\�8��b^	�xL�XA���ή8x;�̎�C����ǵw ��@:[�+H� {��-FXx8��s�����ic�b�wp�����Si�}4N����oy%n�c���a��l�����v1��*�dڍ4�������?�c�Y� �N����&u����-l����I�L~v���*J�#@E���(ދ�C���ƚ �dk�����'�ך�%��q��\
[șC	�^k�K����j�D�w7���Rѥ�Z2����嗐5@�_�� �)�Of����y�W��}��\$��[�'ͩ&��d�+�϶+�����0T7BvT�uC��B�;�M��./+Z�;��?,"�%�Q�a�T�o���0#�6�V\�~1���["����.�M�{y�����1�q(��HA`	�uf�H��\;s�	��=E�kv������<��7[�������d��Ơ�o7B�BK|��� כj10f�O��/66x���1&$+�ǂ9���tZI����q���a���90D�#���ݡ���������ZG0M,�4n��+��B��/̔\P��K�:'�'	��)��H FU�EhR�����ڭE�:�Yܙ�~�g�y��\�m�:�b�.���b�M�G����C�JR�X/�z��o@�����p UD��g���T���VK�n��kk�}�
҈��X�b=i�^�n�WTR��2�J�[�U�x� ���t	��2e�G  b^h�����X�P��鸆#��{v���J����*���^#��J=�Q��rB��˖�=m�x_0�܉sAj]av���,���׍�}��U��mvN�����'F3ߏu>,L�^�F^�ʉt��`m���F�I%�� ��H��OeD���hr�@)�,�H���9�-�g�{/鹛:��t�9�G����U�}���*�hA6� $Y+�̣��3*<o�~q,������,J������Z��W3uh�+���g��>=�����m�+x��]�T�[��4����l�<O�-��3hT�r���&a
���؋�d��#�C�Qi�����=��E��9���z(<>��&��� t$�1�AE�D*�zs��%��gѝ�బ	�,\�}�6r��3&Ό��{}�L��Dy7�8�/l�@"���
v���ú_��b7��_F�@V��E�|�g�죺�#oP�<,�w��d�5E_UM��1�Qg��TP�\Ri|���ϧ�AԲ�R�j�2nf%%1��޻�DE��h�t��d��vE6���o�3�x������l���/L=����o�5<�,����JfA�r��l�~�T�x/�b>��^jdg�N���unSWX��]}w.�p>@p9��!��N��x���ps#��������1I�"v.t8�V !�.�_C���+�1��F<dҡ �����@w����"0��������o�
��ȵi��������a%k����e͙
~�J�.wG�WxN�ʭ�r�g+��WY�ah�������FP�8�z���� �[�=:�ioC{��,���a:.5�]]unH��a�.)/���>��5�;��m*�@�T��_s4p[T�f�$��1���g��� �-wX�"yi�y-��#�9C����&�E�d[���c��� �nww ���W6��J�n]��D�9*��l�:P��hb�&*�0�ԩ�4G��%��]�%{{��4H�`�<���4#n[j���	�w���/�͏F�i���''�����O\�%�U���of�R�u1��C��g��J�	��$W\�T+��Y��a�&��i��-σ	z�p댝�����bzj�-3	2�����`B#�Z�$d�8V.���j����h�� JT�t��/���n��*�GĢy�z��p�SX4�D ����<� �+���T�1�>&=��Q}T�Ȅ���ZX���,Cak�a�ݵٓ�.���h̹�6˅sJ�i�-*�F��S"�|� y0Z�&=�~%45qj���*�B�~iE�A$'�h0�yܯ��945䨦� ?z�����w�`z}1����
��F�����:�3'���CJ���/��p�i�RT������d��0���n��P�7)��,�g��*gZ�W��z������c-����N���8��%o�� ��k""g5�|<7]q�^3(P�1?qϡAcLe�[�_.v����l���@Or�G|�������fA0���3�����i��Y�4�#XƨH��ãӑ�.	����6�����x�VDZ�ֽS%�Α�+�*���
�?bր�X���'����4�����B+�ӊD���B��nnl����Q:�!ZD��ՠ&����"����K�:�'c�!u����D�PD�	Oa�FS��0�9L��.�,C-Y��>-D#����%�Yk���l�F����	f{�9!��PR��\o�4v�}	���Lm�J}�&NV��\��Y��,ҊϞ�&�bm���
�~�����Cu����U�����зUN9}F����d}���$��#Ei��n�ܻ��E��l%iള�������v����b,�J��V}T!m�3�|�Gx ��c�=ل��Tڝ1e1���a�	�cQ����qk{��K����?xE�����U%7��3�~�KP���mNa�Y��+[b������'~�Gvm�w\�$8p�a�����$���u��)�����M�|q����mFϗx#_t��a�ıM$͠�EҪ��/��B�%�Ȥ!w�������a�,A|��cT�լf�c���.�c��퉟��I��)��)q�5W��_��Y�Uw�+:�f����=��CX��NNJ8���go��Y���3K\_��s
�*F�-���R-�'P
ڴ%�*,L��*��0 N�)h3���A{�  a"6�r��*h��L��F�/�FQ�Yn}<l������P��I��+�{p#xC(� .�T�ߘ�-�q�S�b^9�D��O*n.,��@	�� �_�腹����eCL�b IcY��_S������v��s��$�\�A���̷�.�䬹D
�qJ�n���䁅����\&���Z�{�p
$�����mi�1�#>z\�Z�/isb���n�b?��3��X?hD��Y��)����aȘ�?&������^ˮ9	��{B:�����7��+��ע����5��uh��D6�d}\����P��. ��r:�|l��e!������;�qN�y��F������gW�*�$��j`L �>�V�l�a®���}ĺ�����s(=uI�݈��@am ZĹ	L��f��l�L�wà��+o��@ټMW�q�6^3o.~Tfc��a0=��@��0e4�,��YsH��;[W��d�?��u.��c%�<n]���<�L�@�*����#$c���M��^xÒ3p��M��d�,�C�F��=�ټ��D���g�W|���mv�A0^l�H4[�U�Ǖ�!� �M�׬%�:H{z[��v �� }��|���St� �
36�r%�{ʄZ2罖���21���RP���v�y���/>��L  x����a	�eA��ym�Y��TH_BXP�ȧ�ރx�35.o�G��A�e�����]�7Vo(���>�����a<Iw�����x_�$8ݎ���[N��Gx
��.c�	��xD֜�Z�VӤ�$-/lj��Ќ�}�����J�u�*����b���D�ޯq�k�zQ�}^4���J��8����S�~%��H5Υ���H�<S"�6l��r�)ۺ��0��*E%�d����lY�F?�â��|{��%�${'�eFU�>�y��E'��g��pR�C��E3�Ϲ�m�F�����������s ��-l:z�[19�w..���i!�hX&��g93o�=�&����.⫥�1g�V��g
xX�6�#VWf_�B�*�)7� �'�󀅬��f]��X��7t�o���EÅ��L&�����<�d\� a޿�h���"�@�&Ɓ��*��N��ˆ_�u�f���Y��O_����9d+�*�#d
9Nm��(�~>_2��ݾ+��ڪ��3W���FG�:�rhMԮ~d��NN4�G0��hJ����&[�a��j�+�UL���i�^'����{�6�Ó���4ی$[�W"���1����'��rE�O2
��dĦ����h�@�g�0^�U�zzg�f�mt��P6��C+���`yk��%K�]z.���ը��PU"Ⱦ��&U��� ���J@��Z�x��P����RӮ�¾X���%]�/�,)��;!����3�O�����=���z�3�H~	FѶCI6s�a�ϳ���#���$>��H9)�
u͐�옑�T�7��0쿤��ݍ�.54���d{���3I5�w�c���E�zyr�I��j�9����|��KZ��t��܌f�0�7SGF6�	� W���}`��eFj 'jTZ�K�|�e�	B6�o�C���b,����� ��z8';����U-(~�
[	� �`�j{b��s�Sg���)X�26�!��+0���D/-;:�ʴ�P�lb��_��R�}6h����r��o�F��B�9�Ԟ�̺.�	��T�U��^=S��N�AJ��#�̷������7ݟ�>���9��Ǖ����E�t�4N���o�]��=����X�+o�P6=#%�C��۔���3T�^���(OTqơD�9�2O������������5E�nCK���$�Ƌ�����e�����@!p�y�Bҕ���(��kAzM.�M�	e�a�p;m��Ȣ'$�-����O�`|ۆ�.�;�m���|\�f5�V4�A�+�Ǵ�4
�\a�`��_0�����ꌨ���K��]��}�_��W�\mlx�,��`�VCm��H�����W�� z��`�ٺ̩b����5�'�K�J�.2jn�� 8ؔ����vk[�\U��ۿ�s�U�;��"�˴�@�i�OٱX���LM��0���mG�p,R�3BM`��ur���T@`w��({�z�������T�� �&تZF,��� ���r%��|S%�����;a�[�u��c y6�Ǝ�1�}Jr�V��"��ڂż�P�<�	�dE�u�T�If0�opLv�S-��̣KPjp��Sw����J�� ���`yY�Ր���./C�kS^Y�LOK��}]���7Oó���Ze�/:.��k���qs�I�����y��H+ܾ�`�M�.�쓮�x8���=<ЪE�+���b�/O(��h4�t9-9Ӻ#���):����
�JN�n�o��d!��O��Ή�'���7��B�n�A1����ج ���q��n@�`D�8"��9p���7d���QA���7څ_	�����N�m��wDݕV�ȭ$�go׌���2�:0/eq�b)ʎ�+x�Zd7��Cc�_La���%2����x�:mO��@3��[�Bԗ��B=��]��=9��M��k��rP���!L��Ry +�������i��A+���XLօ�h�k��_izŭ��P��8�-����/.�A���Hz�59.г�CF������$σ�?����A�)p�%��q��|��g�� �j����+%������w��QӢ0�s9����لPոu��+G�\�SVg2�Wf��k U�_oM���Q4���	{o�LEI���mJ�%�MfS�����9���a:L�t�"sU�~
������I��??}��IqM�K�
N�8�i(ʘƨ���]�3˻��:���]�:�^�G�~��ΧN,��^MǞ��C��8&��QI=���Xd�ND祄�߼����U���~���}1D�7�\A�C?g6�	�����@�0����#f����<*	����3O����/���?�GtC��_DuC8¸�%��G׃r}~%�ԇ�ʧ]��u�W�����LI�a�~N�o������]�6Zg_�g���&�!�".޹,���*fy:�)`2�D�_���
n?��{��Rw~�&
ζ�{��=D3�0������%��"Y_���^��
	�6n�x@��q�d�KՈ�H��"�D@(Rq��3��ӂD=��Fk@����n��ߌm�FdPN�k���d��AZ��2=�L��Qn�R��D,3t�ڋ��C*�'�4y��Pj�-�b�Es2�H aU�9f�ü��v�#��
�^@*�cߥ��S����*�HF���z� � �6�*��+��D�V�6����p�U����n��}�VlW�V���1��7�QDWM���e�"�	�`A�Sk��RuAY��
�.o7��
�����_ۤ���+� R��$-��_�;�4��<��L��2y�,�L1D��%����cK�'�M<�,?u�uh�X�����7(�Ź��mKR�v��{��ݒ�
#��Q{߸��|� �(��Q�Z�_Z��Q\�/)�#��&W�ޥ�H.��D-��(���*��rC�P��,⦋n�&v�L�)�a�Rr�bA3����ރ�p�ڈ��&3_([��z��\�����n6G}�s!�7�3�����)9� �][�l]�q����K�ܕ��U<f+��{��-K�c+�������yAA��G�t'	}9���a')ka�߫��h�&�h���f���c�`�F�S�[��U��|���?]���UD0�3�G�V�����9���ؤ_O�1h2&M�yM����[{�
���q���dGJJO����Ir�E�r}����7�{U���j�6� ��`y�*a���z��io#�.���&5������Ux*a4��h�+״nެ���ֳ����T?PV�
�Kac�#�OPb Cn�A4��.�5�/�x�
�@����7Q I)�2�������	;ЭNm��5(�wK^�窆��b�����<�4S��a�瘞��N̿c6��lkqO�3*2J��_�
��o�w']�R�$�>��^ ��O�	vu`Tl���ϴ?������C9�q@3�����Vn��:���]�9�K�����?Čf�[B�Uo����js��T�������pP����\!9jCg�dH��-Q��'�7)�9ێ�A=�ve�eۏ�]�w!ѭD�`���H��;Y�d;t���[��xp�@6X�KտN��P񓵩` p��v.h���9��,��4��H�)1/��K��at��A�v�r�6��ϵu�S�J��C�1��y�oGc��	�KҦ�Wa�$���X.lL�jOrֈ�BH��K�N��6�2��v{^c��1���r���ޒD%������{oՅ|\���i��D�x����$
� �̂��CG�#"�|~�k��*-������5�T�ynLhj���Ao��Ɲ!����e&*i��/ۗ\�F��S�GF$��+NW��_��2�v����x�(����g� �Zt/@���$����Z A[}����M�q7��:��ڱ���oۙW��z�ip0�줻���8�
_�4]�kj��Dd	vP�c�΄�P�V����^|��{���Vy��g�̔�7�
!B���M����͊Xx�n��w�L8��g����>�"���,��Y�`��p���9���t�mRNM���M4�Ӭ���ŕ$���Z�V>1���M�f�`�wZ���'�'7��wO�}�
�PMxVB�3�m�>�z+�F�K�I�=�ޜ+m����5�	=��TjF������9��щ���s#%�M�|��K>���'e�c�
z0Rk>�3�{�L����e��u�5�p��
$Ht�Z�H��a�3&�b*��8���,���*���'��<MԘ1�k�������r5����Iͻ�m�f��z:�s����}g�s�h��~%#b
}�gu�p�9g1|rq�W���C'��{�,������{���ꮂ�<�����g?�{����lp�N%����O�-�s��`~	O��s�2l�g���]�>�WM?�
�B*mCp�J��+�m���^�c�=}I�;������f�AEJ������P��/H��l׳i 3JL�t��,�v�X)W8�.�����K$���( _~�)L?B�Au�Ƣ3�J�������N6V�2��u���D��q'x��Y98Ǹ'�O2�c��IDf(�;H9���P!��%��iX��� �v���щ�>q��
��k_M���Vd�����_����O�^�m��v�>�H΋#lI� �h������Qo\�k�w ���7n_H�E��
�i�ۜ(����{�_o�����j�r� ��Y�$�\�%�)0��� R��b��X�u�NVc7���$c�����ۘ	&>E����U�3�KF�>��I���.� 窠'��� ��T��<��*�X�8QxT���8�$�+��@:����������檄�`|=g.ٞl��(���Z���ix��
T3��1��kۻ�������� �sj�^�oeSaD���z.l;�Gj⦘�ZI,u]2���)����o�,*-��'�(V¡��v\\�d�������Aٖ0�{?��(�enư�m|�*#�Bd��S[��s�f`n�t��!/#k0yzE����2��Pi�^�BW�ڂ�kY�e�
m@=E���asa} ��Ȟ��DX��Iݽ�\������ύi�MQ��qS �(��ӿ�h����7�I]nr�r1�?��/���#������P��	٬��:�ȴ�d4F�)�Z3�G�_7X�Cn���8�_�Yn���>����#���3w�ʭeD`kN�Dc����`���.j��d�^ץ�,�?�=�sI���Ƅ;1�Y�=�Hvŭ��I�>��F%��p���sՉ������]M�-�jt-i9
�7F
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB���jSAs���ݤ��aC��U+7��[Akv�Eދ�-(��(�N�fa�zm�#X�����8�@���7X��qV�i�J��0o������2�y�z.��p(�Y��$� �`2qG%N�L I�=�<�A,��mo����(<����_��T���%�͙aY��?�oj��2``z�9o֔��~�]����@�����(M��W�f@�����h�߭���AFP�-̈��C똱���Î.N���%Wߍ
��d��{j4-O�_让\	�ّ��zMN��{�
~ţ۠����O�.���/�iq�q�p��OA7ʆ�B���G����f��@����W���܈������l׼��xk��L�DE�q%��,��P�5~H�]��.X�(N�Xn"y	�����Rk��fi�
��9��^v��T����r��Tp�L?��MC��`����O���N$ͻ�r	q��j�y�TsA	�7L�K,�(b�$� ;�RK-�V�#�翑iu��d�wnQ�#x�]6�XP�B��P��p�C�h�����۷�
Ꮮq�)}�?���v���?!���+~�:�H�B��
�H- ��-��ǫ�;Z��}mİ��~z�͖�D�,�#Z!Q���S�%s.�g��3/Hڮ��pL��C���]$y�Ѓ4�A�����}�����v�2(7k�<�q�{\��09��~��S�u�D4�Y��%��&���&	�����[�K����3��;��P�B�]�-.�L'��5W����������hv!�tujJײ��+���T�����x������{Rr�@��ɍ
��4��?�%��D�p���:u
q���e,����<��dC�è\�g"��4B��ΤEj��
t�C?�3��p��#j9�؃T�@�~��Z�(�t$���C}��0ρ�K,�&>C�3OLew�E��)I�b؍�K�6�ntH3ƻ@�t��٣��|�Ƙ���g���&&+f�V��G�?��Q�1D_�*tLh��
�~�9(i�Zx�@��ֱr&���8v�K;c3�1h���g������z����4���Db��!��_4B�Ѳ�[��nE�y�3!I1��;�3ق17+�r{X6�����W.�lžh����m�si��+��( =��8>jj���s�ǻsy0�%l����HE�{�	2��r��F1����Q>I�;�m�HY���ޑ2c
q�[����	�!ң#EVg'î��4zĚ��5��(*�Z����)8���d�4J�0z%fZA��A��I��D�C�B�����y=h_(��P�2~"g޹��������%��`�0�NX2M	:��
ӻ3�eT\)2o��X�$I���7��W�2�*( �[�E�Y/r~D�*	���_7������дa�Ch[Xmm'MN�ݗ E�����I�J�d_*yG��`���~:G���)|� �)?��g��E��@��[dF�2�@c+��cڅ	D�RV�7�
_�ߢ�3@&j]"[����cZrUQ��/�k��?���ib�zpf��H����\�H�?��l��t܅}M 
J��+`S�9���J&�wb�`7�)�,��i�����	 �X6T�I�H��;3 ��=�.���9��)��]���~�;~W��!���j�vо��Yo�n��M��qA�6؁�v������C�	M����F�[�d��UMjx��a����$p���
Ƕҿ�[���i5��.o��l���P�?��Pxf2�/�D�T"��dF�������m�O�&��79 yؕS����j��ύs�S2�7K�7����0�"�!�`J­A7p���R>p>�Oi" ��L	<����B�P��IJ��Hi}G���/@�I�G\z������s��L�gn��.qD�#X�)��a
���:��>,.~.��E��%E��!��-)$��t��It�"�CP�1�
maoK	��N�k9������n�O��� �}������d��������Y�x1����i��� U�5٫t��1���r�ݜ%u��*� ?� ��p�5~�8�S���A����A��V��R GI�n�J�ꔾ�g�}3_�Ko�~��Ǽp�a
r�Ϫ��@�I��Ϙn��u9�g^��}Z	�:�+���*${Uֱ`���_��˧��	�O��L�(!�5�t:���Z�W˓x���6g�A֎}�9�6����'f{��W�"��b۔�6�O⸆߰$��<Yپ��_A/1�}�w����ӆw�9%»���5�����_B<Xٚ" "���Uk�T��c2�v�W��K��ӊ��?e���F;}��b��	|�U�+:~Lp�x41&��ڋ�8�R�nH�S���׵B1���n�p��{�%z	���h�ĵ�4~��בA�S�����hLT4V}c�Ԅ?FT��)�fk�"T�u!��ɝ|7��N�ܯ��(- 6*�^�����u�3�G'�Oa�SE�}�zŘ�ݒ_#�
��kڎ�й�]^F��u�n9��rT�d�&p�'`��}]l 2R�b'�߫2s5��	y���2@�L-� 
�$*XaSB� \���q�<VҸ�P%��ao<�L���������Tm.A6cȇg������}��'���c��Ĉ�����������^��s�p�ՐuԠ�35b�ƞUf�Vi�C�-Zۆ��L>�=Cs�96�ML�ӆN�������{��-�,\�"�� ����Þ{�>%���,��VA�S�͞-��R��P7�����	h�Z��:�fuP��~@���FGz%�������/֍�6x�!��>m�������ww,��}FV�vʡ�!������y/�V �;	��N��S4�ʝW.��������h�98��k4"o,�s���$}fd����c�c�o� �͍�OmF����ԪWڶ���DLD�M�9�{��q4|�����C����� �����E����j�����ã�=��=hM�5�i=����i}�}�w5�3�6����Y�#V�l���X?�I{�WGq\P�GB��M��֢/E���yi���q�����
@U�;=p�tfv��J쭥�Ila��(�J�%�26>%�0�CQ���.��'^`������o�M[�n=
[��3���dE�5��8�Oz/JhGA޲C�&�%C���V�k�$PJ���XL��O��dɰ9*��3bW�k��yi��Iȋ�IzTr���I�Ws�)����u��Ϧ��-���H�\EKx�S�۫�Z�7��V2y��ŋ0^��
��� é�g3��%�AM�ñmoά,�S�����yw�v)�u=s/`��,���D�S[v�U������*��(ꩠ mx�K.#�5�o�Q
�Q*���J/���Q�\�͌�gi�a����cL8��Gd0��Wj@���ƛ[��t/"��Ⱦ��*��Q�Cf>�˳�`x���o7Q>=rڄf���2h�S̶#v�*\��c�f��I~�)u�B��ҡ�\��u��>e���gC�0֧�Rڰ�K K)�j0���S�̺���!��"�g�O��{L����Y�X~��EA��`�fq�zK��:rY�bXV"�Z�Ĥm������|Qb�[Y�I�8ߌI�����	<��6����_���E<�㮏����~����nd��?6Gd]�̦~ur'L�(z$���,�ۮA�FU�2a�#eش�}�Ҿ�M�*���_<]>كR,�_���րК���6DB�_p,4iOd�~��~.�o;o��枅�x��������������M��)�FVRp�� RV�S�Gn��LH���'0d�7�>�+��	�;��0�>v��m���N ֹċdH��:�U����N�z[�m����+������2�������s� ��Ơ�KP���d==�uL�򍐈i�A�Ć�x��E�o~��D=Jx��v�([��!c���=*>GvjYfﮱ�T>�&fC�ߌ��R����۲���d���-�`-��TJv�����:�C�8�c��Fj���'�RP�G��G����I&�ά���O��3�H�a��@넊�iC��*҄P�^�а�Mhx1�<�RO[;Pd����no)Q"�_�"67�h6��َq�<�����:����$@=�x���@�2-���$�Eô�G�Mq��X/e����	bgMO\�6?�	�0��P}�NNfK���~H1�y"�p��G=�㵳Y��#�p���e��W>�ƾ�lc��y���,G�X���]����	(�.���^C�K@���T���Np
|�.� )�#˫��,:	�F9ax�V�V�%|����+�Q�L�WZ��[��^j6�sA=׵�Eb��L/��_�l\����MpU�ON�E[/�b��^i��`Į��T.�"��h&�� �TJ-�����s0��l����4ã�<�>�}s%/���6a�����{��Gp+Mu�a�g���R�|%h��_�=����y�/���}}Ah�E����ZXx�f'�InYȦ[���}���=��vw��T�%����hDSv����SHں�^D����K ��ݠpe���%h����(}>f�W�0FU���|
��	,����Lf`e3
��ђˢ4���:��dF'����e1
�}t"�r�S�L�B�-K�ꩧx�i�Ƶ=��A��U�DV���rg��鄒!���Au������*s��(#���vEG�I��^���V�^@ؗ%�T򮡟�'�OR,Ko�L;'u���� �$`�����,W ����S�Փu;����N���I6�A��݃X��Ɠ����!�����kg�RY���]>��O�Ԥ�u�*���&���9�'qD�����f{���� Q}r�	3�)�O�4w�����S���	��j�Hy�6�Q�Wx��g����t��:�	�դ#B�v��u[>���p�}�F8�6��}Ď�����C�js.�6�N��� GIұ~SUE��;S�@!b]��k�*~������}}�)�>���0$ǚ����F�ՈW�����{m}@��}��-���s�l�TǠ�m�0��<RiyA�ݼ�ޘ�:�����|�a���Z����F�����ZI��:y⠐2�]M*�X�.�3r{��@� 6��і4 ���$�	F;��[�o��l"��n�P�[{�|6M�y�V;щ.%��)���|0|e���v���W;�,�Lv٥�>�S�S��`:���	�rʾ�M9>��e<O�aо��c8n���9�N�N1b�����vکH�
s�k2Z��i�����m]�?Ta��q[-��.mi���$dk�xRZo���}}Y%�⦭�f�˝�������j��&{�qH��0���G�KC���xX7�ݫ�E��}v����a0�ѻ?�$�l�~M`�� C��?z08])w=�������_��0��$R� :Δy���g�P�F0|��n ���۱�|:������[<�Xd�9��b����D�I����!��\&�ff0���LX���⩥?�?j�G�V4�:�E4�i�E�d���`gz�=Vr�d��<�(�Áܘ��߮�z?�lC��K���n
���3`ܗ?��<*�:�B]
D�.㍄�E^\��Ϝ�$�qWz���ꥍL�7Wu��Mक़΄uw���i�q� FЫ���J���VU	L�v}*ײ�/�ط��[�m�W��o�є��4�E&S�$�3��Y�˅κVx2��$�N��F}�TI��贚T��G�`�S�T+�g���闇A&:,ұ�	G[u��E�Ҿ�C��V3�'DU���m]Z8����8�2)D̪Π�
��%�3���>�w��e��]i"���NJ�9'D�Ph��ND�0,��SG��'�av��iH����aVқ��U8_��>�e3nCd,mȦ�w���V��?n|~2Y�C؟j��MӍ#�$�2�c��cpo�9�[2���v G<>��������\@�,�����^8.(0x���(���/�S�������fS`QӢt��[sUC�`FH���5-o/_��Ǣ�|
^Xf���#]�@E��5���b���}aKo {*p��P)A��,�[`�[��.�'�r�Z�Jɡ�i꠽��ٱk�P�Y����1��cӖ|9���O���j',P�7m`��3��!ɕ*A�����Uֶ:�X�y=am4gdC`��GX=j%??�H>�^t>`��)9W;U\1����B������,	`���2<��#X[�U�3��G��ƑѵalIG�$;�`9�i��-�\�m2�k�VD���C�1��G�*P"8P����y�$�W�)�rR�h𓦫��(	��[z�[�&����r.}���'T�?
�U!M͉(^ײ�bA�eɤ�5eĉ��7#�3�0��M,�SD�T.C�%}��1�I�Z��i;�v0�{\7���ۇв+f�Ũ�ڥnkn�/��LH �ۚlqa�"[Lv ���Cqv���������L��Q����������"�!L��"�w����d��"C��j�[R��t���UIv��1V�ɒ+�; �J1���[��#�c���`8TH��~�6>�:"TZ#�R+.u�T	'v�A��ZOѶzR�ʴ�~Rpi�UJo�TёACg4nN���6Р�GnT���t?M'n���rG����ЫO�Kcj�~�R�� Q��fk �h��ݷuBy�CVL�N� rY�U!l�"�	b7�t3H�0V�k\�3a���������)�0���j6�2��s����(ǭp�Uif���nn��h�v���A����W�>U��J���p!����!�5��ck5?h"�t�Z�����raǂ 8�j�7��$�FM��f��� X8��6̓π�XIP/�j4�c��4�2Eٿ?���&;��t��jCﲜ���	~��B�lf��T�9/�r����0���V��ؼ�&���rq�0�@v�%� t�x��0�2���>2T9�[��^������^v/��8O{���e��O_�����Z�:l�`��R.A"��ųd�>��g������)�(����Ӽy���\����$��"��.�[�o���Ӿ��a��M�95)�&؟�o��g�s�ꮩ����\���Zx!��4���*��$��{�g����$�V�������c��x����5n��%!��Q���RsSt�b0jV��[�t'�y��Ӑ����������sJo����w)�U�Yl�7����OR���x�9�;.ʆ�g�Ϭز-0ۏE7.�Ck.�r3�a�s�3PU��s#%x52e��������.���'Zb9ϤE��zh)��6�/�n�c񝌥%��l��2��D��k��t��)�f5Lhp �W��3EA�Rh�.�U�Z��ᜓ`�Y|l�K&iQ7��7��O��gܙ�W��LJ��Pqﮯ�إe6%N���.�������H�5��� ���Y�.�P�T5p۰��䁖\�+0їLJ���6���w�ƴ��z�)q�jҲ%c���<T1F?��+����:���È�e�Id�En��M�	�(=wW�˭��n���@-&q�^�����c��N����^!M��S�1�@+�~�("��̃ӭ��f	+����Xeł}�"8AkӹW�W�{�?j>'%&�L�F,?�������; z����H�H�~�&L��>bl�HZR�~v�``
�GƻV�=շ�>L��W 9v�>��6!�H����lEEP�����yWs���2��]��L�?�Ϋ⿕p{��M��R�������UP��~����E�2x���8�n"����`�8���g-��i�۷�9�3{�)�w��c�W-�j�]��2^�V�ҫ���&���尷o����.V<W�[^�Yx�
oD!��i��:~2ܝmX��^����?����8e��l�!N���:U8$�kl�p�>�ZZ.��To��
��Q�#�U��\�`}���\�_��?yupE���Єs!:?~��	y�2��@h)�=>Y��F���gq�/^E?��8(_��S�t��M@�.��ͤK�
]��:�����wH�{�q���H��)`-S�$Jb�
Y�l�k����I����m��T�;�e-Η���0����y����%�,&J��K(j쒛V����2rs�a�`�\̞ͻ{v<?�}ؘHc�C5RY��Z�^�>�r��T;��8��� ���$yIlf}� �#b� �y�8�adz"yJ�Y�C���כ�! %"��Az} Z.�ԣr�5��ƴ���"��y�]�ë�n0�u����D�
�}*���r�O'�O��q,�k�G����9��o�񽕺�:Ԇ��׼ܪ��蚷�ZoZL���Ox�t<��5��e�
ɜ�1����A	4����8�:a �ZFDTpj-���8ڐ�e :�<��lD�)����kx��v8�5�?�K�	qo�Wn��,��ҍ�BB�(n5x�!���H4V#~���S�]�)<_ ��	 '�����Ѐp��!�$�}z�U]�1��K�1z8"(ʧ���R0�D'D�2o�<����T���u��S�ه� �	M��S
Y�2�:SdCr�P!njp������)ڨ��|�?;�=���L�(W�GD��4�\���b���7�f��yz��@_�O<����{o��D�������#��,r����Z�Eϼ +ҁdo"IQ�^��V�p����" �\�<�ŢT��U�2�iժ��_S���n�cRW�KR+�J�#�.��>ڄ
k0KNWW7׫{m��q1�T4�hr� ���c"�h�Q	V�|�>����!�b�8�5�(-� ����Ϣ^�Y�_e�lo?�s��D�J����xs��v���=�۪�'�OR)��^�b����b\�&A��񒙋�m��dϑD��r��R;�j��A��\�l�Pأuo�]�1ͽ�?19/M�,� �|-X��+
��!��'�Ӭ:�n/��B.���Aޭ��Ep���_�/K�^lC��'����o���¥��K�?+C(jz�K�K�Kg�]?8����u�ld�A3��AY�×�]4�>#��*\7�Kumx�H2��,��X2�RT���~`�6�Ihl�{��S3�-P���M&�JդD��i�q�P>50)�\(��Rf�������	W �W���_�`���p�X(M���{n8!P��JV�kߺl����)i�<��Y{Dkt{Z�7�z�r�9a)������$�a��'�5S�G��z6I0R�p�L��$1�:6W9{�Z�ʏu��!l����t��8;�jp���9%қ�猊,�P>o��nP���k��G�9��"�+=�a�}����
d�v��������@]�Q���g��j�2�ن=�M�}�m�y���Lʀ^V�n�,^z�a�K���К	�_%�i�[�����5J���7��p>�����.hk��A�G����v(��%�P�@"������;�_�Fgޟ���=�	
���"g����ð�(;�8S�t
�#Hf@0�ѝ=
"|�TR\��ZLv���Ch�5=t���A���F��o�p��_-23�~f��"�4@h9�P$��i�?��S(O<�1Us���.2Z`p6��P��îv�s��J�-���	�7�y���Fʝd�x �1Ǚ�~§F���^��@�*I�F�ث�@/H���7���펋��F�pD�'��v ~f���'8�i������i�J�'��_YΛ0=��A{O1��IHV1��$�VQ��Ӓ��6-����X[�e�A�6�V�p����STl'&}��"<h�^�N1u�[�ҳ���r�+���'2�=a�>�X��a]b'��&o��M �k��9���_���S6n5�r����i�	�#��4
c�c)h6�{ Ͱ`��*�$�.\K8������t�)wk�+a/�_�&���%N�.�[�����x��hz��vW�E�EJLm�bg֏� ��[.��YM�f�ϸ0�*w?*bbO�e�oٍOH6����h�%�{GP�Ũ�'�	x���+�#}����Fp+hd8�	�S��+���,�(���v�,T�s�o��*�� �1�1���M5K����>,v{��%��Gv��,@gf��ӵ}�黓s7v}��~��ľ�fs8����ɨz�j[7��c�;����V�l�:�,% ��$�v\,�b=	��պx݋�1�]G%{[��s3�qn-�֞&6�/�h�LE��:�e�ژ���Wj����gi���z��5֨����N�o�#�x����8��#���j�E�4����&ݼ\�
\��/����?�H�g���&���c�������2��0H�ZZ(II���ݕF��8> �,UaⳊ��3^���J�aV���]������]ً�(�����$Gs���K�����N����}lʊ�k�u�v���[��f���[��F��83*�0���u��x��g�6���d��]��_7w�d�3۴ϱ���i.���>�Y�*2�L<a��s�i�ݙI�vv&m��NV,��r��^l�0
!�/�[K/�NąD����p�K���-6���m*���B��X�2uх�؛��+��<��EL�VuN�����c}��[����:���)���3|�m�HE��H:"B����$�<�¶���wV0��H4�C6��@C]�~�Tb%*�+�d$%��CP�A��-��s��2ݳ1h�q�����*y���s�ЯwL{�J'Ge=��9>W9�����g�s#��\V����+��L��)�6�M(p�����j�'�0��7K!P������b�Uk���P�q��.m����y��RȳC���*-�R���w��O�����*�Y9CíA,�w��%�"���ӥ��#�6
="(N�0�Y��_���qj�p��yY��H:�8�]E�x�T �!u~7���Rn�0�����_�Pv[g֒>b7�}Քvs�����o�&%�'�%&�gX�u�(�M�L>���,C��{�КA��.�u@���`�����'7޽(�#���ܠ>q�d1}�k<~{�ߙy�>?x�Ѱ^<,���Ӕ,��	(Z����={������C�_V��/L��&'�j�w4�VGP�������U?$ڎ��K�;Pc��Mv��ͷ��X ��*K@��V8�b���
kL��˘�Sl)�]C|Vze\j���1�#�w]|평\)w3�U�=���[�2�5%�mαi�# ^eɑ��'�G'j����\ae]�G;��рK�=���gŔ6�x"<$ߓk;B5�����zrK��DN���s$ "0{!��"#��b9U���Q�����^%C7�����۲�N�����} ��)������ +���#���H������	��x^i�ƩV�tKa��vM�\A��!	�L P_�f�e��P}9ַ�!�e��hZ����琉1G�3�N@�|rT���2��m�EY[v�3��X���3������Ź^RK
k>��0�8r�����Lc��#�<��XS��؄��ACڞ֭��{�]W ���4� ^#���I�R
�ї�tv��X�+�
8��+��_��.���dehӫ����(�,��:bF^��N%�AWp�{^|P���<g��`p�� k�ЯK$_�Ok+�I��OBt`&KZ�j~c*և����i�p��^~:�(�"!TE
�]';�3��Z�����kv�&�V�5�[������.u�<wr!	i�����%Ja�o��`vp�pm?l[`�J7�{�f�{��E7V٬$�5�\\s�5������c`���Q��߮ޫ�'�a
�uJ�]�����v�����1�M�	]��9X	�Ȏ3�/,��ɡ>�\@	��:��3<�x�������ْ��M��T�u�J�pd�����4G�6��1B���629����̤���j�W�����I��$ڷs��,+c�r>���..�*Z֧K�o�s��]*���ݮ��3�&W��4�9�>Ge�w� ��{VW�YS�k�؄��ޞN���1�y0�_0o�X_9�������d_f��F�--ߪp;Q����tZ���h/zҿxe����W��U�|A��WZ�h-yi}�#+���6ڌ���]D�V/��Z2qĽ�dk�&yEqb����5\�ZU�} �Zh]KT�3���8�B��ݯLZ-�`\��n�c�rḾ�q	�պۀ���Y�-��&�����|E�'��ދ�*���� �z��wd�dN�� ��3�Y*u�u�Cξ�}�uQ1�e���4���nq=�i�<[<-�o�a��u���l�&\���t�c�s�N^�h�2�|@�5�_U�P�1/�~�������Y���C"�pW���vӸ��;�3���F��g?�3%�h�困=B�}��`@�2d�p�ξ����]	Ruje�`{m�LP*`^ZbϜ�D��� w�Y�� �M�VX�%�=)]��o}���+��̨ؒ���/�S?� ERo��^_\�F� 3�2C�&}�S��e�/�K��Ÿ��u>W����K�w�"��Wvn�cS1�P��A�!������x�(�nh?6ؒP��A⡎?���Q��+R����4�i�Ǹi�@yа��p:��^�m����5�_ՙs�:y{���#*2�~���bl�޷.g���k/Zw	 >|FG�I������1@�.���ё��/[<���n�*��1^R߉@�����-�v�C�9%��԰Օu�)\�!儑�� ���>>�.�:F4&����&����<�kwkx6�R1$�mbO��x��r��ǆ���1��|��(5�\�W�~X�>�;I�ų�X�B] ��B�`�A�|�̔dQ�������3����.De=0��R�P�4�S�;��D��-�Չ _<�돨�d7�9}%��W���b-��� �<b�����fR������?
�S��Fȹ�$�O��A��+C����ķ<����X���v~J��}XC��ݿ>rJȢ(/�]��3��O������p8���Am���SZO�'5F���w��~w����@��4�贀��h��>��a�c��O3��ڦ|�|���Hp6
�Y�w� H.J��w���AW�ft�0BM��,��O������N7L�	�4����sp�9���*S��ْ�G5"T��u[Q:)aHԼ�3�j-pϲX�9ڵq�v2��a��XM�ʠK5��j ����WT�nU���V��&�2�H�{(qn�
�=���6��W3���+��:�#1zy�S{'�U�g�	�7�'� a�~���A��4'�4��~���a6��:�j����&�������V_�&�=i^/�uǫ-N�+���C�@���O"c{O\I՚G�j�~�ݛMs��Lކ9�j�%�h=iZ��j�~"@s͜� vӢӄf���E'nX*�Z�RX!l��)Ԍ:���] 8v��o�����o�p��ƌv��L��c�H������'UL)/��V�C��|�W �����-�d;J}/��9�X^�n�3n���}��ym�Ꙥ�ř�/̳W�-PU�\�[uB�Ƽ��#�B:�&����L��9o���\��F�G^�{@��fN��b�~���Gi_��o�?5�x�tDXD�P�+m|,t�-~����]��h�6�@��g�述�*%��?��I��73yz>�}��r�r��uk�@����n�}r��qO��?+����2{e�c˭<~`Z@J%�jP��l���aq���
�{�.�����8v����A�g�Ul������F��օ$Gn��� �2����l��N��R�!�;6,G('ѕ��LY��ӿk`͉�W�7v��wgP�-����F����`��d��%9��/AH�Y�$7oF�Z�H�����.�G��<��_�NS��֚�|N���<�b�w�:�,y4�	Cɫi\�KE��Z�4����D���Aΰ�Wc�F �]�лhP+�⥚���+�{:�R`pL��f�$���f��}m"�tm���./��KuTͿ�m9W�@��u�c 
��r�� �U�9$���Xl��~�t�_D��MQ�_3ڝ��S�
�S|� S��P1J�̬Y����_eg ���*`�ʿ6��)	R ]�tBKՁ=u������4^/g�}�֍��o���e�����r���&�Ui����E�b�ە~�c�iX ���/fvƷ�Ɠ�\Q8����Fi�����].q����D�ߪ�RK���^�	�ޛ1z�9w��)T�9;9�������?�ʚN�I�>y�'�����U�� ��.��?�D7 |�Z�����M|�+Q����Z4K���5�l7_����/�!�y#�|�/�e���B�5��M�e����=/ �	��E
ԤL�
\��nb�)RVP�'��T��=�X�l���lB��'�����g���	9���E�F.aT��B<�J�p"����L����r�(/�o.W*�'�^lW��eg����B1]�D��)Wo#�Y�(��r!���f��x��fk��e~��p]=�����f�=�tK=������?���I�m���=l��fT�$�q�pn����G�S}5�f���6����������-ˬ�~B��
9~ؚp���b�4Y�@/7�]��!,-3�Z��	����S����������dx���(;:g㊔�NiN.\8�ҏ@t�=�6V83��ς�vk7��>9ok\�a��_v��0�vd����Df��F�}I���W��FW�Z����de]�5NBv����H��j�@�j�b4��8�F,�Y�f�A�����k�j~~0��q�l�b K)�q�jE��%A��ft�~},���.5y����<l*�53wC�ͽ<���2Hѝ���ϸ3"�wy.T�W;����e��I��LI�#��ږ�A����j���w*}"�s�b�~&��]X:H����?P,�V����W1l�Y�л�?�#�7�)�ą�:ka��
���4�ti~{���F��<��I�Ȇ� �ށLb�wA�"�7��(����Z�9�~������&ɏ{�0a��s���!�-�Z���۱�\�����'�Ԏ�c���}���]�`Z{���.��r�n��R�jV�jv|B��o��G�xo�͸��Z��j\���OOW���(k�"ȶ�H�ַT1h���:>O�DP�V��XW��&�a;���)�U��!z���tY�͸��m�Ggv�N��K��i��M<N
3�Ľ�ܰ�$���f��>�'�D����í��~�����3�3�����+�IHq�����k%q�0�� �w`�`�VG���BK!��侫�/C)r�O8:��d���f
�_�?�#���#�����Tj���ltO)�t3u�%a����dv�Ş�g�\܍Zo^�ɖF��� �j�M�~�tN�(E�i|ԫ4�*�������T/������)�j.��n*�1��9
��D�b�x��éUu�cF�?�װ]�܂��+���.�/��E��!Q�}����֜�UL��&���A���u[���d�g��r��������y�]��pg˷ ���h��m�7bU4�)�84��R`�{���Y��T�bz�et@�=.����v�(�e��F4�)OВ���9�(.Y�E4���F���P'��ӓh\�gޓ�ki��;�at��F����H3{)n��ЁѩTs��]9EaQ���I$���6��H*�^3QL�>�)�Io�&�b��]B��m�g�P��Ó��6+Iۧ& ����
x}��NuP�8#}��#�6u�f���r�"���8g��0J�xχ�[sI��I!�`����K��G��ݬ6��$��ap1_�k�O�*WL�N�ɗ˖@��W_d8�(;�{�e�ۿ�r*�>"��$� ��0 ���jH��A��Yl�->�{���Rlu�_�a��k݊o=L	F���G�ė��T���V᛼b0��3R>9�"!Ԓ��4��1�"�&E��pfu(����K�<�;��k�z x�O�����(ޮ�9��>�F_{�q�e�s��aH���&����r aE���B[��_��q���L .�3\��Z��ˋ2aB\2��ز�Rዣ��)���^�6�'�#� Y0Sφ��
~%��϶�+����W"SW�v�u��M�ek��^r��t,3u��z��Ydx�~���0����/��k�i�W�}֏ͫ-b.�K���������{���Ă�7UY'��0��6������k���Ou�LU���,�
.􉕷�^��.ϥ3zqt0&��h6��O&G輚x�����y+��;��|��Yۓ��4�D'�ƪ")+���,G������������y��t��i�|�&���m�A�x�FC;�$PK�d��ץ���_m�P�S(�%V�UR��I㡖�j�νa0�HtK�K:�~!T{P�(�T����]N,;j��Y�;7csD]�r�ٸ���2o����Z�)��_+-+���ν��'���V �M
)�i�4ބM����:�Z����.���C�e��`��a#~����n��g����
`X�t6�:�2�)g}�֪dCaB=B�f 8�����Q!�����zH�oz2,�k�n�?^�\7�󥺲LXP;�v����`��y��� �R�KT�i�~�n�.�f3����!��H��E%N�A[�Npw�E@$�4>���	A�t���a+�5߀��Vh�y�q]�BL��9l��p#�ˮ~��(�:-��:����@k�kV��ϙw
3�}���/�t|��F�L��f��47����`����tj+��a)��T3����-�����L-��F�.J��L*��>߅2	�¶h�S�*�1R���9l�7N-����@{�
�ux��8�x�1��6��-���)����E]R#�_ʗn��t*��8�G�]f�����N�ޔ'�-�~���;'5�y�Қ�퇮ڽ�,�U��%ԋ�L��}"�D��Ω���l�i�T�Y�������U*� ޿������7��i�-�1�����*��?lI��4�(������v�<��8�M&�E�R��v{��~ӌ��|�~������AUǚJu�7�gK�G�����E�V���뷝Gb�J:y"�j��Ij��j�ٺGbm�c��h�e �E��֧x�x����Z�|��u��\�&x��$-ݪ�bJ�W�
�و���B�[u8R�Ã���`A����;9�+Tc�46j�2��.��0���^4+�LHI��o�
x���%SV}�:�� ����B��v*�P��*���=)���wV^m���&Z�O ���2��=�Y����xk$HRc'�e�]����Q�8�a|�N�ϑj��q���5��ӳ�Z������Б�UeY�'lPOc�`1�J2(�產"�*gc�].���2�.q)�̧@�fg�#"���RI#��Rs�A��ת<R���
ݶ3Vs�S�]�V����.i���Z<���(�AVٔj�Cl+a'����5@<;���3�\����/��teY;W	@x:[�&�6}��۾y؊���2�Lu+�Ji��#p�i31Q#yo'��H�A�l�H�h�*Ȁ\]vs pe���Y�s=.��l�>|2����z����y+�N���������?Nq;ϧ��_�aՃ��Dw+p6���=�]ӵ��4$FSg��C�x�p�q����/0�9���#'ob��sY���o!�-f�e7�����E����({�Q)�KP��,x�/���@q��Z+
��f�LmH`���t��٣Ek@A+HJ�� �SEW_�pK�=C��H��6��M��M����Nf]����������. �YkZ��h��nYS�O�96!�VWj8�VJ+��6́J�Y7�gr�x]��Q�"�R���	0<f8��x�gfK������զ9��z��o�?��f�����J�ı����ڻ~�C˱V�^����"�����'=r�D�1���m�u}��ސ�OW'����C��[l��b�����i�=��,��Ia��#fŪ�B���+T?��Y-�b��G&6׋ϡå���	=YB^
O�&��O�K�3�s!̫M���J�X
w��Q1��V�Щ�!\����2�(��g����p�ƿ*Ó��ށ����%���)�4��y��x�k�4�Q��>ș��k��O��/O�Պ�ɝ�����H���`�/�*��w;:�g��̛*�9�<��]�R"��+����$3e��0yǛD҆�u�aPM?nII֨Z/��3ϻ
�X�n�_�O�?�O�i�)n�4M����x�������;z�c���q��x��My~Z~l�^�Z8��'��<"%6x�O6��j�}�w�P�sj�c�ާ�Fi�S���~ ���K�I�@̒��I
�*� A�|�gB�y/��8�M��B9�&�v)-`�$5��xf�[u�vƣ!��U����7� �\�%���k룉�t"�;����4�O����s����^\@-�R�~t�d�食ȕ �H'X*K������4�_�b�Dbb�~��1�&��S�����/<���_ ��re0�-��_F�jK���:�A���`�[��P�W�&*�u}
WVV�Cy����C�k�k�oO�_xIEޙ=O��9#�wCx9�-��T�6�w	��qgt �iA�ٝ+>�[d�h�h���j��2\zU�8�ռ�$���	�����jß$ԅST:eh�y~�ڹ��F#ڐ�4�a\4m:���kŰJ��|�+�n���㴮I����L,�01�}�!'�x����LQ�����3�m�K��{c�xcu<DWw�#�V�y�t��s�8#���a�¸�v
��1]��;��}��C�'�Ȕ���ao���c`S<������F�0J�����Y�f�Ls�*�����vR���_�#6b��Na���yw�Zf�sX0c?t����4^jY�l-���Z���V�w&d�q���J��,P�?���O��~K�o��O��q%�[���N���è6B��v7�2$�0�	�5��8'�H�_�yM�䃮�o_�N0##�#dSR@��B[T6�<r�o��Z\9�R�S`{�L��LY	���=#��(Zvb��r��~�q�\�XL���U�QILxݨU�m���[�)yӊ�d�]�fhh� ������2��%hsdnl栆"��ɝ2W	i�n�zdݭ�U�.5h�
�B��=��i���u �JG�`��F�#��C��6L�x�x"E��GD^�[���j4�r��`F��.r.������^݊��˨�L�V�%��Dí����h��Qx4�N�R�f���$�G��9�rx���e��z�)^��i��L�8Y��2Ю��NE�q�h�ha����:TsH�hd�{./DV�ʹ%!gpzl��=['k��ӝ$2�*&.^��������0F/���ģo��k�X�陋�t	��݌[K�
�R����1�=h���߃!�j����;ExRňr�}�~�7��6����-�I]g��Q��&cyqP�OL�@���slg�6]��(���9�U"FW5�H�o�_���L/��>���y������ntf/^J��.��t@������=q�f���w^4��hn�ȹX�]�xY���$.x�To�M�ł4A�U��;����-.g��m6|�$�L�-{z��R��A�M[���f��MhS=+W&BaCڟ�ѡ�����S]k��_;X��o��I7w����؝lN���h}N\�\5�l'j�#&�JgBե���-�"�@c�?Ɂ�U�F#��w���q�yK���Bf���:�5�S�І�Yu����HɕH�q����ξ\cÞW��(�>MQ��p[��j�uAma�1�1���`,ʖ�q-�bdܦ���9�q
�FA�Ã� h���½�C�p�|6�ee%�d�wA��Gsn�Ab2.N7����N�/3�#o��&�G�?�����6�wDq����U�9���--)s�\�1�琼�셨��_-W� ု���e@��C�B�S۾d�4�E��[�:rG���3~3?����U|�t.-J�C�iC2+/�U�9z׍�O\�:�����Sd��Ӈ�-t����J�-�ae�)+�w��)տ������׉$7�̏�/�ǋ+Q�����a&�)�N��	��k���ѐ>$���S���e�@��^�ֲws����@z9b����&d�`��ƺT	�Է%p���g�W����>�4AZ(��	s1��GӇu��%r��LI+�]�X�ԋtD[��v�Q}>�D�a���"W�x�h.��9�	�"�o1��S���"� ���F�����GIF<�'�F�D?x{��JL�
�L�օ�X��_=k�L?}�!����˝�U��p�5�9�*Hm����j!�#�P�s!��
��'s)h��{~Id�����q�U��{"�`\(z�
�Q�	1��P�ז�麔<�F ����s^��PS+ŵ� �A�-�A��T�$O�Q`�F4{�=E`�@wOu���d}Z�3Uh��]a�5�HC:\����)LF8; GO�֛=N�5�P� *��(�70���O����� K_�+���hב�nx0������6�S�d������2m��a�!M�0�+/5���ե���J�k�J�ՙ��w:�U��O;�9��_S��͒ʝ��9�#x���l����(9��F �#]�]�V�����O���0���	Y���t��!(HSo�R��P
6�S��'���aAg��Q�f�������1����ˊkRO�	��R���k u���"�|;q��>�V����y�b&l��;����_�EZK,��0�V�!"��&���b���$yN��=�:���uonN ���d�7'}�iT�nx�9;�*����c��%�_VcW�4^�2Ч+�JP6T���xo�)H�Rx��	x��۫��E�7����	v�����wc�"~��PZ���!ى��E��s�����W^2n��p]鎡ڤ 7�������#��x}���u��	o�A�Ɣ��(U��+�$�g��Հ�#�7�8��m�	��DyT!y��X%j���,�;�i;��u�S��fʇ�p��xdiRB���Jo��]�[1��7;��1�i�̐����_GѦ�"P�c[P��P֎J�74�c�A)i��ՙ"�`y���92�Z�$h-
!'ȷ�m�y~ǃ(-�U� ۉ�:��-�pq9�:������T O�&-V��Q�a�l.��N��l)V!�vԏ�/��}_ s5���Rt1�������"�KvN4�wAR��}:�T�w ��v)�^��� :$�<&F5�u�P�q�0|.��[�RN]�k2��A40ڸ}4��^��i\nƄ��eI��R��t��R-N��*[@T�V�I4^#�~�7bl����mb9O	�v����?��HS����Q���5Y`�Dq~�SFϒ��q�:��)��0ӹ��aɧ���r?�d��3dR��s#�V�����ڙ|�q��z�3��N�bjV��&�S�T�v���+���϶� �L�Фk5���:&��KwHX��YDHU(Ag�<��u�>�vl/xo�I��-�ܛ���?�Y�v1�z�2� �fhb��n��r	[6�����K-�G�ͱ�,N�r��O�ِG8�M-�pi��	L��#�%�Ju�Q�Zg�ԟz��2_ȅt��4*@W���`�kѯ��gX��xߐȭ�]�
Q��u���
'��sR��Ǜ���+�:�jm�[|*�ud�B�i��fn�}�1��=�`cGji^J����<���P���������$[W�6�oD4�(�e��,�ş�vX�A�$�>n��Gѽn�r��1���qRCw�YW���A�$#�������@�wi�~BG8=s佻�ޒ�wO�4�~B�P����r`=k����T�O�L��PU
�Ja	'�'�6���q�x�H�6r��~�p���4�rھ6K6��Ia����GhsCT(�KX�2����雉S�����C��'�r��Hn8��1W����iJL5�I����^6�jU�WA4c�uZ��h�ە˂�S%l����5�1�	��'*�PTG�6
�F"��'�޹��i^�ى�B��0�B��X$t��h��}����1C,5���'6(�����RW��[X�M�3+��N�>�Ea�e.��r@�F����hO%�z
Ed!�
�Y�z{��G�DP2�H>6��UU/M���T�A��~�RP+o��	���M������W��,�ϡq{p����OE5&yX0�$���-��A�y�d��2&���T{N�p�5Jz��8"�)���k�@A��'�����k�/�[��6k��F�~�p57|��j���=6~C��Չ�	n��Q�W�@�/�}#>�Ə5�R�v�ߕa�
�5?mãܒ� A�2��(6f��qn�����h"�M5���Rc�B>�Urh�����@��,ч��߁Pآ�;���hpٹeZuuD�{�U%��Q<�O�����z�<��<��/&�SnWm�� �&�h�ٝQ�c��ߤ��63���w�Ꮑ��?��{�!w%gGUt������;k��&�gvZ�P�|$�2]��)����u���,�Z�>�$CQ���*q1�[��t��t���\ɥ��wR���J�؜u�����`��;Rs���ݲ�ڪ��v���aL�_B/'&W����2����Qu}p�y������$�.|}������*
�����ڐ�~����e�u<���az�'ղ���oJ���.�,����s�Wtٍ�U���j���;��S�^��6.���@��;W��7�����z���T6r;�����:�0�wxp��oO�cY�a���vv��@��c5޹�C.�FM��b�Rby����0o��֡&�
��d*t�#_��^6��ı9��@��!3:~�:cKɅu���6@���$���L�;)8j�	��a��C���*p�N��p#)��X��\��S���$Xt���RrB�rV��e5��*��Yؓa�[�Ȟ�ԡპ���t�`;��o2�!���6��v��h,wѲ���b��[��{���<�.���ԫX���.	~Z레,�k�d�ѾORW=���9�ߛ�g�N ��I�V�WZ�d*�'����Ikg)Mўܢ�ف��� u�o����,���R䔫�e�s'�d�N�ƹ��S
.��� 6�-uB�Q$��u0��pX�q;��I�_�ׇ��e����(�����fs�v��Q�.OC�8�>Ks�V��l~n�1���Ts���C*g8u{����J&y�6cӂ���"D�z�W�gh����
$s=���3n��� ���;���x�6�^�kƴRU:�X������+����������̐I04�gS�gql��N��L��/F���"�'�D�:����)@�d6~}_�݉e0���q
��pI�;==}�$��1��"8����=�LÌ=K`' qD$"��m�2`W���/Y����Ͷ t���B��ZbR6���rL�.XpKy:w���
1�|�G�C�ʭ� �)�	:ɓB��9~�Z�1*'ݝS��.RR\����E����u�5�&[7%�𤜚w�q{Ր6�.�RsS�,������8���t+G�Y��>�o����v�
87z��х�@�cU��t�$�枎�3*p�(�	ڼ�!Oz�S��C|�>�
.9�Bl�V
�3\�������vnɐ5�O���S�0<��5HT��p����t������G8)��#��W�8�t���Z��Ӵ�Zf��^���s��\ߏ��
r��sּM�H̠����yBV?eR�J̡cMV�ټ!J��IZ�����wv��}�+D7���7]�������mz����7q״%ѹC����^��l�`��V�9�a�L�a�Tj%��t<|V�T�y@�_�Z
2��wQ��?X=D�������d���s_0�G��n~��d��$$g$��b�y�-�Lݩ~��{���9����2.)G�8�u�){�8�)��5��
*/j�e5��{�P��OY0	�D��KW����iֲ�"� �:�s���v���3���y)Sj��KB(��8��6��,���)z�ڞ�$���B�u��nhՏ'�ؠ�L�	j����٥h����悟�����+��'H��;�$���	�Y��a��L�o�?��6$$�x_5sV�h�	�b���Rp��hX>�D|0��5��5'�jh�����>`�l��A��c+\zD����v+��Qԝ_�ĭ|ͳ�7�?�����Lty+�e��q/��sD��t�9ցv�c��,u�^p�ry� _.���r��Դ�^.�
���D�4�$]l�D��s�40���@��֓N9�:��:_�+Fl!N�}~�����D�55��Xa��og@S���8�r��[���i'�LN
 �O��
&�S���9��m"�vI\�U�d�� y��ܬr�P��ˏ�K?��*��B	ڸ�V�'6�(th���e��XWU�%���p畯E6ESD,WY�_�+M#���Yr�?͇RcC�Řl;`y|Sr?����W��uW�x�@����z{�v��n5�^��^kk鳥7n�Gx1nN�X��3��/̔�l�H�5�pP��Y�#�w	�k��� v�*`��;Ɏ���B"�VeB{rLiE�eJ�~�&N���*\�>���D�����8CW��?��'��¤��_k��eX�}��Ec!y���q����� /��2��ByNTMM��cRQ.���D��z��+���\n`V=��o���� �4g/ ��͞���J1P��U����62Ǵj��ھ xno%}�~�p�!��c��Η��>�y�udf��q`{<��Ʀ��*�t�� �i_���z�1��W�/0`�i�����g��������uPpٜ��y�/��7P%�7,{�(���+<{�u�d���x���W��N�o��D����u�O֠i=&;�K����y�y�;�Uoʱ��$�mC�p�by��tWZUD�n��&kx�2����i��Snߋ(�r� ��(�ˋIՓ��զ�ɓo�
��)v#�-�&t��^�����:�yÈB�h��Nˀ��9������I��[�AT��B�n�}��yI���>O��y�;qҚ׎�&e����s�i��Z���Z�����h&�kOK>n�tU	�f,�X15 �(���KU>{ڒ����j�u�]�YcPG"`�!�X���)��(�H2>Mo��hbv����!b�n��pfl��f��6DF�.�J��	1�c#���g���\��E�� �Im�,9�{]�\)���L�O�ڥ�a���>�4�f1V����H��<ԭȮ>�e�#UT��<�	ΕI���:Rg���C���)�M~�b����ee�b�/���ɸ����9��]�����^F�Y�m���4�c�
��r�����oDg��o|Hy��06A�ªY"`n�S��U�r,�����t� ]
&�})j��LK�k)#-���g^�m�w)�j��b{�Z��Mm[<�nk1�R�)�ai�`�Nxs��0�kX}��O���J9�)Ǯ���4�_/:��o�W?F�s0��2#}P�}[[�w�>i�u0�Z�h'�[0��{��p��tY��S�V#�p5y�!|R��cG���ne>s��o�rc^O�T��"���KqZځU�%}3��ߟ���9�����t���O���ANB]qp���؊u\�� ��'4�
9؏��Ԟe%��J�,\�<�n���pM��.�[�G�}�$�$n��o��+�-��XC��R[+u������錵��8'lq��p�a�A�%Z�<�2�S���I�Bq�d��`���wV�e�9��dZ�ia������@�z1�pdv���O&Hd(�0W]�2e2�s������g�MDlEey�I�v���q]������-L�EjYf8��+��L�V�ɛ+4ҍ9���1T�H���kè����Ӧӧj��-?�[9,8F����C ��Mx�zژյ0\R��B8��zB�}r��Y%V�����y\�#cE�f�Qb,�/x*��mT��;qq?L]1�O6l��f�ĈA���B�\��~��O^�Z�T�����`�!��(C{�Dx��h�q>��ݓ����Q�4k7�r]@���\~��X�êi�ߟS���!_�/C�I�����P %�TŹ�J�>��V+-B	9�
���n������񛆝��U�|�{��N��&{T�eX���s4i<�:�D�dW�k��뛉*F��o߆�inObL^8��U�$��DN���-1d�J*��b��ߴ=B!`mod-J��?y<Ք���������,d �d�]�S�v6�*�"�aX_9�dN��Y���t�S�X��BF���ٞ�R�;kс�Q	0ﲩ����Y��K�l]޻`/|C*C����B��bl�gf�0F6јE�ߝ�~�5�ʦ��	P ��q��a��r��G���A�(*�ݚğ��>al�:C+J��W)qx"g��kwz�5z���\u���X<>��F��oewF��O�
�:)Q��'���s̊1}�/���0�1u��pBMpn80O����9<�oFm�������AF՛$ʷ5���;Q'�Q��P��榻�(��$A�@�K;�I9��;Z��Gf�o�Jr�Ӗ\B:�"}Ԓ-��eN�3�Z�����"F[l�h;Xox�#<�qF\N@�ɪ�5׳_'��g��WK�\/B6×-���,h(�נ�D+��L�/�Ҿzх	F��U;��U*��X�2�*$���q�lNԳd�*}<留m{w�{~=��7B��M�3;c6��ާ��D� Z/���@��ٟ46�E��A݄��'��@�Pe�S��)�-:~e��klH�k!Dт5�cڢ�Z��yc��� �^�^��g1`Ƅi�k�Y:2�����Eac���@	+��7{�E��,o�5�<Ǖ~��T@��|���s˥&����x�[P��d9��0y�'=Ϯ���<��V�C�l.4Z0���^j�%���V�dn��/�5���HOֱ��7>����b�4�uk�Hd�p/�8_F�{�?0��JǬt_%ڨ~4È@?�}�s)���7R���|^�-�����%RKAN�T@1I�i���(��b�̖�L�Dg\e�Đ�T�d[��!�ޡm+w�@[��/\�^`泦�!��
���y�F��Ss����-tǖ�iI��T������?��)J͙of���r�|�L~3�`�(���Q�E ��^9�@�_4�+��i��5�l�s]R�έhL_��亦ͬ��%�&K#���X��K�x�RA!�y甹0�x�;pY��*����������:��pWщEK��j�/�i���b�]��!�(�d�!��f�w���
g�׾q�)��p��{)��=NƜ�{���%��q��c�%��9ĦVkr����1�4�%D��
�"LlCq�:�����@�z\�%Cu������PQ�M�����	��G��D�Y俸�]�WW�ٺC/�3��k�*Q~�
y�`�3^���.��i�51��kɮޜ�7� ��P0|�E)�>~4ђ��Q�f�V+d�FʸR:��3���hrTau3b��/�KcA�!�ſ~o�����i�S2Ni���Sߗ�4r�?�2���HIqXL)5H/��`�pM�L4���$������2��>�./��\�I�Hm�u���r��s-������~Z��`�A_~�<DF�G=�^��	�0�q�.�A?�r��f��N�D��b�]˄[J.�;OQ�BND�T�I�9tۧ�o�l�aB-��<(d�~ǭ	���K�Y��^0����v���!���J�v��$z�h�DV�W���]��T,�'=����O��0N�RF~���ItF��_��F�\I_T7<J9͓��Lޓ���=X!j�>�"�}[���>��/�����R��Y��Xw�UD.��]�����G��&W���\d�����с�Xevr(����W��C�&}W�ERS��L{^�;Fm���Im��hFP��\)@qq0�Ҁa�۫���uz��{,s��-�juT��'��N�v6&��u���9Q'�/l6�L�����S�Q�OR�Kx9%��G�9�9ߚV�g��@�����g��nǃ�P���@i, ����D�R�w=�18av(]R$Xj��4���N7]SY�ޗ�K�M�p݆v2���U��`c����A��D/[(�Ǝ��>K/q�p?��!�Uy���@��n�>��PR_�պk�E#����U��Ɇ�CB���kr�J�.�ӑt	�
�G"��}B���A�+s�`@̵�d���?��~�؞���;�V|�[���rFy��u�_Z{�^�IF��U����� Zw�#%�]M�&��s2�8_=D�T�gP�ˤ�GԬ���Yh�s�쟹�r��c͙�`q���|�D�O����>V˗nF,.����Sۤ��D<�7�J����#���"A(S�Er�:s �l��`<�,���v�*z/�*�h����No�����6>��py�eGlcN}'e�f�=ݡhz��������ѠS-y^��������7G��Hc*�Q��/��(�M�����<��\�h��Q3B"�O�"g]K�X){�ғ�)���G���T�w)�Ԩ�t���"�@H�Ϩϔ����_���`B��H�-�����[SZ,bݲ��ܓ�)>���ʃ��x�� �]M���lp��0�V_N��������q4UF	����Ն�"�1�g����39��$��z��D[ͯ\�N�'��]eE8k�����rHT�� �P(���N��J&;�0��K`�xJcZ���Rz���LԌd#�k���'\m�i���ē���~]�0�"H�r�Po7T��� �!<�q�2뫠�Xn�*_�[@l��¤w|��&%ܘAN��}No�b���zL ���\iR)�m�LD���m�X�$4>҉0�m�Թǈ'.�
��h=mO�[eo?�ҡ�',DZz���cG�,�bd����\�E/
�9~٦� ��j���.2��d8��|�iT����1ʚ+�՚�q�Ib!��dٗ&�\hV1�G��*_��?*�&�RZ�xa�u� Artض��������G�tZ�ϱ
r��,��L�KJ5&)�/1P5Zf!�qU>���A�@
���)�p�&�g⑦��[�N��!H�����0���o'�n�#��f�q��)-�����v}y�ݶ�=�,���m��<�z����_���dh�HfV�-ٝ�H��=���n~v���G>8)�	!:����8'bi�覆����b��j���X��������t]���d�7����@	sGV0*zu��	��̊�����#q8�8eyB&%X�F�D�YUc*0����;�~����g:��T���&��%�D�1�ert���$,h��ڦ�3��
s�TL���G��W[A��X�i���@=9	��U�����6��{q3��`����o#]�k�%�#BʙȷbAW~^�{�˿i$ZL��MA>�;̲����T�<R�Pwy���H�C�
�y�
@�9ͮ����ZT:% ��(�O}^�͙�� �I��>�F����\2]�U@2��C��
j��n�% 9�o��À��c���.��ss�5��| '�}i�=3?\'�dk�����M��Syi��^KkЀTfn��C ��Zj�Pd1$�|1|i�H#[M�"X
H�<��+Fsk��T?bv���>�f��)6�i�
V|Y���Z�#a>��sa='ݜ����W�u- �8h;x�,��M/���k���(D�Y�	��R��tҬo���b}h6|S
;zv�i?6Crͦ�0���.Ҭ����x�� �:����/cc���\��L�OL��|BrL�׵*�E�k��k@���1���=X�|� u�<?!���$����G��k�O���̾����U��K̿���B��;�f�w�G�m¢�Ox!�	rM|w��CΓ��L��oE��N�(�����߿�����6=.���>vK���F��m�2�#�G���qA��֗�P�Mn��P�GT��/�\��K�����H�k٪, ����t�"He���'���[{)�,�j�aau��(E�m²��u�݌5p?�E�����Ǟ��t��UM��V���s�Pa^�`�i�I�ڤ�d��p�e��w���t��ha�dK���˪� 9`eDgpIj�ʟo�2��������Hf���ɨ�n�42�@�Ό­����%��1�`RȞ$�uJL�Vٽ�_���`��ѭ9���'oOJ�h~mT��z�4ԃ����}I�5��'`v;��8�?|�D���`(�恵H�%Lɓpp��fR�Kr��c�LG�`���ܣ���������_��s!I]0(�I�%�縷����(���}r�zaLA�2�>�^�S�R�+W�(���*�Z�-�c\��N�@p�"�bj0p��-��Z�.�Y��`@ފ
���u�[��A���`z�dF��&uF�P͒#���EE�Jgw`'��y��zI��+�w�p�o��Z�Y�׈��6N:�F�Z!��B���{�u�>1Z�Y�(��D�i�c���ӭ!�кr�Ol�۾�2s?��<z����+�b�ۓ��M�������t�A�?;j�5�j��}��F������i���c���f�&��L�%1J��yT<Y$�,����r�W}�̍�����Kl�3�k����%�_�6��<!:���G�pc �����(b�v��p� �B���$X6�BDl�c��$����FRM�oܘP3�0��'s%"�*�EY$@�չE_+�J�3���4�����Xl�iI2��#�G�{��/�;k�'^afef{�#�����c�����,3���=�lٯ��xV�%��Rπ�9���A['!^Q�Ũ�@S ػ s�ڈ'���ơ��y8} z���g�w.ݸ���R83ӝv)X�`�<��Yp�҈ڣ��vY_"}\�M�.�蔿s����C$�tYP$��P�u',j��Ҩ$��|-^ѭңM˹XQg�ῤ�0�z��^[���Ne�v��U	�= ��R0�xk0�ո�f���[wj�v�n:7�B=$Q/��+S��q�z�r*3%4�BZ����/΅X���+�.;���%�e�C�?(ݡ-�V�Ѿ��Ɍ#M��»'f�q(L'a`#ER'�1�)�� 囓�Z�r�YJ|a�a����]|RY �3Cr.94b�����>��b1f0[�3~��5�
?0.�L?Տt7��߷���R�bn��Wb����+���6�b�m'Ө?����?�/8Y�a�Q<Vnj+�z
�4$Y��+-�&s��x���_�jX8���|��,��Ͼ)�_`��U.�`����z3�|��,[~���D�y׎�F0H� �d��+?\}@0�u�f:7���3 .k�ٓ��@|ǻ@n3w�,��K�~,�:�/g��{
��?�{+�4�,�Ȇv<̞%��$��4�f�mx�)���P�/TU��Ѽ��jGǔd��X��L��8ny�+ܜU}�\ٓ���&\}*���k�#��c��	�&�=���0�aث���ט�Y#�����{��t�B�������3�R�v���2\�v��
}�B�w8��U���P	'jj)�)���9CS
�z4�D�B�t�v"������g&	=���~+��9�b�n�{1Z0��ew�O�)��Ԍ��e(:��{�tO�1<��Z���bw���4=�h��R,��xkm8�����y% �3�f=������8юZV͹����{i��AҴx��[)�@5�,z� �	�pzf��_F�J��z,߉(��!��Ve�4���̢���Y���7A�/���&�6Wf�%��M1
�A*q��<k����cV*jG���>KmdD�&�JٛZ~+��9�,�F�*b�(h���qLsv�n\����!&��k���*=�Q����dǑ�!��V���\����r@����[i=�:�(�v��K�#�����+�����"��IB��$R-�B�G�Ub�K�X���T�5� �^9�s���N�g�*ԱY��[�]{�J��&uxW��ߨ[^> �j5d�KƗDGO��\���炀T��\u%�T-�O,����eA����w�j�H�d�{����t�q�WM>Ԧ�M�@�E������7��:���,�.?&<�����t���Tγ8���%��<���c����G+S'��c�cf+T��ik8���~TNhc�Z�{����Nъ�f�&?�S���j[G�O�&3$pY��O�ĕ$��"?�f����E��cq��#Z̳��oUV.Y�����8J�7W%���f�[���4ge!�:�	�_��lD�*)��m�}��==��*6*sj�B>�Ȭ�'���7̾�7x�%�?��t4*�@ {K�#k������:��������W�I	~��:��V���$�(PT��ԧa�'\F/6ߠ������ӛa{�UǷX�8���~��D�c��-j�&����H'�of������
*¼���*_)>�� �q��o~W7� ��ї�Δ��j(F�E���g3����
%N�Abi�阽Fѓ�IU�w��|طD�����4D�#"� VMG�}rmG5���J	��/覩��	zG��4X�W%��O�1�XO�x�ijW6F	\�$�~oܹv-,b�i��	�hxt�fP�5��6��^[fИ�t��y�>f�դ{6[�˂Jb��[���0^�{S��'j��Q'�d����2�w?�	��i�N���8 ��~�8b�Qmae%��'��̜S��+�CG���ɕ�q�6n&�*���G$��bU�����ÍW�B;(�9>Zy{~꯺����=�&0���x?m4,��8n�C���n��D$�;�ֈ�c�iYji�����`�SR��v&��$Y��M�����@8�uO�Q&�i�q[���s�$X3���Q]��yӐ��='[�b��uъ=?&+��*��IR9X�����ԑ�L^��+�G�h������1�Z+�P8y�8@I��L��T�h���o���TA���ۣ;����ζz��Y&d�ń�ZP��ϓ��ڀ��t�[��I��(��	 ���3J�Ѱ�����j�Y;m����~���kKS��=��s��B>1��<�~�n�d@0��k���,�K�mE�n�����vx?��o�D-����Z'`8�v�����9喉�<����]�P$�2VJY��K���sOc��|Ԏ�W����8 �naΛ�+��J��`�Kø���2:���iO���.�^Ɂa"�(wŚ�����t2���w� �/l�Q�Q"��f^�\�fN3%��>��פ�A��F��sH	οzLA&��V���$�ub��]L� ����33>�n1'�Q�y5�ݳ4$��g<�N������X���	��U_O�f~�;5r�9�ڔ�ɤE��(���j=�X3�䦦E��y��M<}
�>B����c�n�~i�2�N�qK�J���t�"B�o�\��.j~H��n�]��c�ճ �A��6
�r$Ø>���Q��g��`�uY��%�*��ѷŏ{�*6������/FL�a7b�+��ˋ��N��3�(�O�:��G((�-fn�U�	�B$Hҳ�r�Y���͆x���4@�����z��d����!�ZoT+�{�?� �6l�ڪנ��K��4�'�8C�SB��^�IH�(��/�}E�hO�z�/���5*�e�qv�܌K��"�.����)G��+g���� �h *��n쁝"y�۩��y��-41��isZ*[��RU���P3��3�9Tlw\s�M*Nc����xb�czg��w�TؒC�2¬�\�S�in���Iib�Ly�y���[U������u�:Vb��)�ԋ�U�^��[7�O�"F�D3�X�0�͇IUz�8�Dg�ؒ���T��v��#Žr.ϬjY��}�����5&�Kr,�~n�c����G��d�GE`���S�By�?^i2���H3f)E���Џ�j��3�$h��������%��]g?���_���`���G��sɔ�zJ�x�QZ��P�>�&uD���/Ġd���PU��gǾi��'�,%�e܍�jx���sխGkBCQ�{��R?|n��S�d��bY�uH؍�K��B���:r���'����r�~���@=�FMZ��2S�:o�8�ߛ�i)MЩ2���^�G�9L"s9С�pҊď]c��F|��������h+�z;�W�&�u�Z����c	\x��Hय��k�'���c��[f����JUƳ}���Bƿ��P����<-���w�ׅسW;EC5Hݰ0~`{���`���ߪ�!W�mW.��nU1��G�e�JE,r}���	��ʶ�|�)�!?��FR���x�$�Gƥ�+Y}�Vc�9��M	h�f�[��WRz�AN��f�������5 j���+e�cEq��Ψ��&�.sn������+f�,��X�8�I-��@���"�_�E�����Щ���ݗ[p���1;�Aq�,w���%J� ��Y�{w�	KC�e��D@���AY�[6��Չ�ޟ,.�͡���k��0�}�+e�%�8(�u�����������M�'�C+���:�X����٥�ߗ�oF��/���&g9T^!E�G��í:�7�/�2��<*��~��C��c� ���z�q�B
�?�Ć�.�&x9����l�y�82��/�v�BCَ�Y8O|��O|��6�ϓ�[���#h��`�8?�;������]Ї_\w9����&�&J��Jv��S��eZ����P��ڦR�儴��QLCq�������N��f%d�c�D	�� �vO�i������j+B��"�E[;��(�'����,��
�P[�(�����R����8��ؿ��~@�6a<t)Bt�lX��K�` g�иƘ��S5A�6��)���땷�
՝Fz�2�C$CN``&e�&䙨��8bCԛ����Mb�9l��$x������� �9`S�D�Ҝ�pJ����+��mu��)��z���Hh�qM��A�1��C���J뭛�v׎�m�#;�D:hTH�0Y�|[�������X�1�ᑿ]i\,�����S���g��ù��.�(�%���F�����M��D��]�{U�`D��y����f�������H���V�����?T	��^XCv�f�-o>$qpg��K7�I��!6�C���2^��+�t�]�лc௓��m#��;z�'��F�u���¹���|{qE1*��'(5��g����I�:|z�C�o~{��,��޵<z��K�O&�=�h?8՜�cc����UM��*�R���_���h�E�6��w�2�5��,/�<2��e��o��A�
pO�\��%��>5ɏ���~)��I��l	�.��@j�s����'�/�m,Z�	d!K\�T����G�zg2e���t��h�=xu�:�T�-R2eh�j�T���r�M%��-�RZ G$2��Q ϖ!��qnb�һ�7 (�_��!��T���Q�/~��$Y��"S驙�4MJ�T&�E;�R��;3Pcp�R/(�Y'�)�����
@x� ���\��`5��|��Bߘv	{z8+�FT����0,�P��q��0<z��OGP�ʡz*��s� ��ś�3��".���P/���7�s�eW�l�W�������C>�ֈS�� �j��C�M:��f�؉� |�~g���/7걷��-�����зD3�t�B���-�KjN���B��>��h����
d�����Ǒ#um��<��~��+�qM���e�2֢C^�W�iO���+�y.~��b��"^��9��=EQ���r�r)h�t�<���오�s�Nt��:�;���ؐ;A�(�mlT�\v��ns]����D��'��M�_�7�J��ڈ��*���W��8�|*�>bW`�9k~!`K�;�WX֕��Β�;]�)6��ӌ}��wX4Q�7縒V;ӓ����2�]�7�[Y,6�z���w����<s�$1-����
'�t1(=��51}�dO��T��zQ�!;�n�VY��l�60.�KAi�V���R4_�y��Ҕ����}��P's�G_���C�U����z����oGj�(X��^�ͪ�nY�K̥�@�����u�����V ,{�w5{�O������b�Fi�FI�A�3<�����c�Jv{墳v.�W�:�
�\�T��p�TՆ����x:4��q]��r8�T�z��D
&����S��b���;�;i���yV�!Y���:�9?"`Z�,��hCNM����p.�ʓ���VV�)�B����
�-Ǻ�H�q���#l�:=H�2������!�����5��N�#fzJ��((2�o�fKʳ�ĩ}F��q��
2�),A������b��)�����9'��+��ض���n���dP���&�ķ'Q7*8�"I����5����t�k��а��$QMR�n�Ym{����� ��?�p�Yy��P{�f�ֺx�U�����0��)�NY�\���^��}{�W��q��~�S�BI�u'⪰̨���I��ԽD�~䖒h�[�$�A��l�xp�J��=|1ep���G<������)�!�q��P�ep�%��$�\�i���WI�q��JL0�������=����-֠Y>�g�3����QX��&��{�Ջ��[n������]˟��6=�]�WH�����]��|�dr:0�'j���u��]!5q:̇٠5z'AZ�@�h�{�6����0��^���uY�$�'���i��=B�=�n��� �E��my��@�	�ɴS�P�h��Wi-i��F��L)�Ǌzhu\籫�|ڛ�<����F�j`����r�U�C�Otj��##��fRx�`F��2��ֆe3AK��SXD�����}�Q�+g�A�0�eZ�������M�1<piPc�'I�}�y=��o�p�l�G	8��X�
�T� �o�/��H��7�n������o�o,�Sy����q�\����@C̎2�+�;�u2���x#���w��KX���e�&wYs�`VF͑�H\Z_8���
p��A�Ct���vGc��cw�ڜ��}]��yMvJ\	�m��x�=Ҩ^����J�L�ﬡ�|��-2C偓̇�6Ѵ-� R�8dN�s)������.H�0����|C{E����Ii)њt��P�	0��z}��lX��"��.�a�&"F�T�����Җ�D�'\T%	�P�����	�l���,�>�N�6%�([��2FA?,���u"XO��!X��N�j农�3��
�~(�A��w���5'��)�����Â�FF7>�;܌���&�X���ZV(���E��F�$�F.�UJ/�8�~�j"����Y#E@����Hn��#�y�����E*����*�냞� � �g
�J����!�U�'}����7�4@��|J��� FVNq����⤭�@�Ժ�*�8lX��Hs��|\`(��?�-�V\����Ǚ��x���w���[P_:�X;�!$��~ C'��~�X�'�`S��F�J�V#k�h�؋>e\ Ru�8a��oY7?3�3릛A��<�s�TP��K:H���{V���[�����B;�6Ŀ	��GD�J��ƚ�� S\:��V
�K$�V��Fy�%bd�r����E�*ж2���[��rQ�ʝ�Y�m�q�W����5��X���%`�y?�����1�a���E�'\���F�+ $�)���<r�V����F�S�tU���N���c�̉/2��}�|*ő}m��r��8�4ݩ�EՁĊ}>�{�VZ:GJ6;��20}��φ�ؼ��~�O5���&��\'g��c�([XP�1�d(����z��$D!�K�0R�Ma%�鲏<�Ev�,�4p�Y��f\��w��4K���^
�=�@ͦ	��8z?�^%�`ۥ�������]._~�Ā	���堮�j7L�8bqt)��~A�
�M��M�ޒ��oL�vě3	�u ���h��N<_��8%BE%Y��f�N���5)9kz��7��}�����*
g�G��:��/����^⧺}�#��������Pm$)ӣ[��4aiE�HD}�Z@�m22:��n�[7�W�[�3� ��*]��5_D�31��`%Ф�4U0,��q��-O E���i<���v'l�x�!�W�+@"����S�p�QlUX�nUͥ|~�������$�Pl�j�2��a|�0�Jv-0��L)��[���D����9������y�["�)R��_�a8�~k>�����1y�*����+Ex$�J�������:d��ܺK�Mz34ӹ74��X��m|�dlxR�B�r�+9�ǩ�st���?Y��s=���|v+���bM�*,ѓ5v�y+t�iِ��z�X��X�2��� �r�(� �"_�uQ�y����z.�	�܉�;��d���Ļ<�Ǻ �
��Γ3�op�
�o�2���9�}7 �,Z� �c-8��b��0��tsˏs�S6ݦ&c����d�z&ٚp�<oUy�R�܈uk��RP����j����l2��ȼ�d��pbB[so�|i��Iޥ�/u����R������B�����u�Ax:3��f�����_dDWP��R}�2�af�d���j3_��Դٌ��r)�� _�9����g�=x��H�����3��BD�?d��/Q��ʎ�{/��o���U������"R�5?x��C�P}���P���׷JVy
�d^�eV�(B�u�,^�F��c��ׁ�#�&�YQ�c���dB��(]�:2�=�-�Pf���]��:',�ϸ�Z��QW���@�>�fz�x'!p5@ĩo[Ɔ�p��#�b��b�R���*:[�t��s��N2���p>\l���Šbѩ���d��" ��J }���p�1���|�)�4��g�����!q&�uf[b��I��8�3�^�u�Y0�ؿ^�F|9,w�@FH5!NV�@�æ7o3���c��z̡>�����Q�a|`�9�����O�O���~�)3ՈS-�n����ч���I�-��!���΀�2q�����Xpu�U�Ws��Z���N0I[��Ig�3.��[��}VԴq�CLX�ʀ��ug��܇���g���I"o\n7	�9<�g��*;z�QÓ���� �u)�0��Al1j���1�N���4�/�@U�E���9>R�ִMC�5��
��)W��^'�ƞQ���s|d�ea��^����Չ���x�U�b:"��Г.�[k��s�eNCB�j�ς���N_ۀ�z�kI#��"�Ksym�����~ov9*7^^L��*�%=�P�L�h<؏���fJxry��0��5�r���	tAJ� �HiqL�y���7��{L�I��A��Ÿ��!m9�=F��Y0@�=1s�Q�����V�{'	�;�)������X"�-���\W	s�0�_��8�����Q���Uc�7?1O�_�c�&5^6�l;p����u�FF��F���eC$UtǯzB��&��^�5���O���Q��Ew�v���#�}bF����>�¸]k
d;�Y��#|H>n���Iw�)��O�6Z�8-O�1�|vD?TFg�l�g�����|��/������ZS�e�<��e��
�ُ�1-����6C��:�@�g2(����g�}@��cL�KDH&���qC���?}bk��f}��GG�����	�Y���(���V�����G�ֳ ��Uy��Z��V���;�� ���~(k��OE���ExYoI�
�ZZ�p�Eʣn�����9����mCB���X~�Nr��:��C�zy���B��
%��C�%���KPV��J�K=}"����O�py��/��l��7��v h]����fm{WFpt�QUҘb�h�<��
st���� 9
{�*�T��i��za�TC�Ɋצ��2���ĥ�&w/XP�9P5>��J�O5�O�Z��*�X�Ua�p�0�Ɠ�*�ncş���e;�u1�i���������`�D�����dz��\BݴmY,�	'R��5��ק�1�Hx����D����c)،��)@A4w�D�l=�pEGҪy"5,�����d�qCj���Wl���L�j���Ӧ�D��t��#�4oJ�:4�-N�)k��2��bw�EC�\��U�S; ˊ��U*cǻt䦖�tvݐ#�������+���%���
�i�?�\�$x�\�j;�������E@q���hɈQ�3��B��٠2UcX��C�Z��C���Y�c���a4xdk%�7�L�7�y��m��]��}�s9@(@��%��z���7׈�(0�/o�"Y���9�jh.J�i�L�ac��3���XgZ�RGE�^��jg�:��V�^BI�J�xٝth-R|������8 ��'v��lm���_kq<I=�z;͡"SN,>9�x���δ�X�Tn�=+Lk���₷�q?P���6�1 =B�0)�sVnsḲ��pE�Kg0�%��Z��$�?6�
��;����c�vX� L�U�&��Ł�;R�mIo�`��o�kPo�Bs\���}�w��w�ʙT�����J^ռ�B�0�Vrڬ4�����L���2qWP��֙n,��	�en �8CL�4o�A��㬟isp��,N��W?	��ʂLUw��hRM;W��m���O�s� ����x�+27C�l,��ظ�H����_6{!�ˬ�8o�i����˶�SM�M���%��H�����#l�q�%��F���*���,s�w�aGټ�H>����6EO#���k@�B�W���i^��������Uo�!�iˡ��Ϧ����M^�dL���6%���lȗ��`=�{*l�i��-!�5s�Yz�灗f!�8WDؚM��°�P|�����(=@�s����f�p�QAr�h�)m(���!(��ɏ��ۿ,Y3��Ů����@�Kn���ĸO��qm1]� V[��:���Fnw�Fn�eFh��ߎ�7*�k�����BS�"}C6-��%�����pR� �k3'W5p���rd➁��l�-�C�8˦���]�H��l�t�X\�%�d2��o��:^���<'��F�o�5��2c�$塀�9�>�F��C���I"�����Y��ϝi�)_�{Ox����)�MM�]�.�j/c#W�|`9����L%����~��O������}��;�����7���SB��|�k�M��/��
|B�o��>��*h�pyx�ƛ���Ě��r}d �����W�N�B��
*�4XKؑ�9�rK����C�`���X@yY9	ooen�d>���(vAa=�f:ZR��nNͩwrUG�(��SP'�3-��͚���0����?ĺa�P��	��jhv�r$ׂ���:�_7�y ��t[i��T��j��U�H�/�:�t.�Ftf) ���D ����}?��c%L�4A����k50�/�E�
�G�޲Ƌ.e��b(�$���4�;P+���Zȼf�9���/�"+��91�%4D�Q�#yY(T��[~�7g���z����S���P��u(u�� �g�x��)�s��y!0�#���,\J&��@9�?��V;��>�ĝW}���d�\��c���E�|��u��j�U\�c���N2zoK*�fP`�)Z׳�q>T(m���S�Q���ћ����&[.���G�'m�/���M�%��0:��Z${����M��X���l2��'8� ��-��%��8��U�u��^z��Zicp�a�����P���~�1k���\} ���^M֙&�	����Zu!��u�Ǵ\<\Fh��ͺ�	69������/��fH�[	I�b�,�*:J�~�R1�z��쵀 �۰ +�_�Ć5 ����ӱԵQ!���Y��m���O��%��au��-��zmJԆһɅ�<��������`�G�]����R��~�o����7����bpsy/A��E�
iN6s��ȅ�(����4�L�X�{2;�,I�PWt(5��)�����ܿ��R�µ�_a�K�Ћ�k��%^R��j�݈O"�)�YeA� k���:�����!�v�9��l&�Z�6_0��X�7,�����d�+0y���f{��J�x�:�I�6):��C�	�N�-&��j�;Է,v4�g}�S&A�� �O�W��O�2'h���B�b�0�_�8x��D�ԑ�k"6R=Q�:�����<1�&J��}3��83�u��W�v�F�]@��tp%܃�H�=���n�t^ȹ� ��;��z�S������\�&d�����S:Z����Oc>����L���6�t��b�(�k����}��>��\���Z��D�!�22M��"�L�G~����z�nq���i����:G4fB�?r}�(�S���Ї��KVS�a���m*-�aM��*|kc�;��6PI��wGɰ?�d\��s��y^��h�|�K�g���l�BtA�U[�
�^z �eqJٓ��v{�uL�#�pdό�Ny�t��s�� � �L3�M�3�PF����;�w6�����I�6�ZO����{c3'M(�!�P ]�u�K臹m�须:���L�j����G$=@�",�hn	�#��CEe��y�?Ah��\�_�Id͒uUj�*�O���L�#o^
�8J�.�G��V����Q����U��s�D�J�@c����7�`kbLf)�ѵؽ���8���9vx���D�q���MUb�cMA.�/����9c�}�<4RA��c7f�о�������<#����d�hD�BBn�J�D���I����tvڝ�����-�ti��I��d1��g/��z=3+�D��5��ah�cd:�S�ȿ3܉�߈*����]��P���+���l�hO�#��D�.'Z��=C���׸JS��7"�?��(��B�Hw�|��3�����M"�h;��lP�G��}������a��(ZT��?-��͓�f�S��ΗV�Q�P���Ί�+[�a_i[Y��*��Ӏ� {XF�?~�Fxz�#~4��(X_ͥ|���		_$-5f:����
��J��՝�\��g<�0A��J󤲬����4#��a�D,���b$�6�w�L��Ex�ԣF�q��� ]����z��l�ʧ������PK�]��f��僻��Li��&���S,Q�yK��Rt)\]�ȼ�+ C��x!�D:�cU��dG����0�Du�ч�^�q���Z�֘z�q���h�=�Gj��֫7>�d�ۤ�};n���/N=�"M+���ey�]Rf�y�H-~(���ϋn�þE�Kf`P��	���`H���ĉ����zx�.>q��E�;V+�^�Z2-A�u�e�����ӈa���.��� �-	F��sN��]P�	�*u�)[V|���Y	&6������~]��}���f��}c��H*���H=�]��ZoZL# ��N�n8���<��\�Q��K�6���؜-��s-�e��^r=��݄-_r�`��4쑨Z��ҷ,�~Q9��&�1��Vݯ`Z� �B㫏��7�$6��
�W	�)~�{_<�y�wH �LΆZQ혶=��*�|�]��]/�!���u&7�6zcz�U��u[��l�F���ί�ak��̿��N�OU�d����/��ƒ�m�(F�H������b҅���h��A����w�l4�WzW~4�Y��Y��8���Tz����w���(��h������l�t�~�_��R4\�HeF�89.M�܈ �q������q��l�=ǎ�WU��\x�?U��?I0�R�C>�Z�iXq�����m������:oH6v�`�d�����}'��g��KC/�,z�e��ݦ:F_k�#�j����j�����+���C9���0���;��no\��ª�A��2;lP�����"������XZn����_�+.�J�^_`�[^>�k�!��8�5�33 $X�rK��Je���l븏����,��5�+��+Pl�W�!�oB�b�D!4F�D���$��]��:l	�*V�"�M|q������0�|��+P����j�_�t���V�?6C��*���':���n&��/��58!�E�A�Z��y���~�/�#zA���Z�	A%�|�G�*D1y�d!�~O��YD�����l:Wt7ZÌ_Q}
�m�ZB�E���+�����c��������-��9�Ell���tRsd �kF�v:�]Ƞ	�@�rt�I�X�=|�iQ_c�2��8�9H5V���)�`�Bb|;�c�"�{4:��}��z��"���t�X�_-G
}�fg�\wR�@���B02�B�?g��N��`�B��nj�
��F�k$�ݩ~��au��X�C�ۍ@���Eަ{�4���V2αp*���,�$�K�PU���n:4��k�i̚a�~@�u���\�"L2r/��wrIZӔ(p���B�V�Y���g���ϻ߮�a@�]ð���{��`�q_X� ╇�Nu��b�P��n�6mK�vq,Y40����Q��)P�g�'����������x+OJ����Y֥� �6���J�.������(���/�MX���X��l���{Y�ם ���`c��)�<�o�Xq�J���k���E�]���2V�	�߬4t��Z]$im���%���p�.�54�n�
-�D�|�PsP16es�0� �)&U&0��fR�:tT`�?u����х�L&Aכbusb�f�݊]��[��(���TԺTX�]p�o�*D���w��/Ĺ'zݨ���&њWt"m & gwǠ�t�L�ƖKoE5t��DO*����U��U�N8r���Q�Sx�Nl��ȚɊ"DB��6�H���L'���U�&�Y�nc"D�)�V�GA�k��r�4�Y��T"*�ҏ�Ik3{�N�?�����dFD`�p.��g��g��}f�Y�o�OZ�׮��<��@��9��"��x	�L|����~��*0��ݦY�Z�D�c�7�$�̈v�< G$@NJ9ց����l\C �'���Y�:r�������[�������(<�=���_�Q�ma����ǭ�������X��G��RjRJ��lߖ=�f�$���J�%�CwE�-3/�^CAFj��PB�CE�K��>��6%���%c5�l �(8_�0b8h���R��{�}���:{X��0��_��L)���i���<E�������VM��H����/��*泝t�gɳ��uY\��dҔ/�T�����TkS1�$6knI���Zc��2�<�U6��$Ȕ�I���Y��{nk���f^ea��(���J�{Gp!�e�O6�dQM����M��t�U!�@G�� Lc.����׺��;Uvn�I`���KlJ.b-��VC��}����\5y�}�{�G�b�8��hp	�oW��;������c�Kƿ��q��(׊�	�''��vR���}���gtn�1/1�U��M
z[)>!҇)%*L�r���1��\���Ғ6P�yVleEJ��uL'��'�%{W��K����(J4-��+r�U
i�\V��rR�m]6�Cb���"�Ed�/��5Th�7�����`SF���>�\����<���Sjohb��9	-���K�(���+(_Y��K:�z<�(o�3E_��O;��VMp�+�@4�1�v���"gL@"�N=��^��Q��ȍ%j���.*�O�)�CMm/����_ug�k?\�9o���S۰�����g+؛�(�M��/�U��͖	�eG�S#�iô��9��K�%lY%��&��[����P�]����KR�}�ɜ�мS�n	��#*L��3��H��*R����G����)E��!OV�����S1�������2:� �01+P���I��'��j��	��K+�����3�G~մ��Ɇ���ˁ��oB���d� �<��=��	�'���|�?T�Z���klNw��U5��������^��;գ-�f>d����R��;5X�gvE����J)�R��L�ڴ½�k[|��,�r7MNӦ���.�~�h�_&Voˢ���Iŏ[F�|��V�Lq�ȇ�p�BtQ�j�g�]��4�`Kִ~��L�#�S'���ܓD�z;iy �A�NS��1`>>�V�s:Jh�n����)Jȳ`��\�};iy�3|�7x�����'|�eؿb����L)�����ͯs�2�L9s����'�܊��>K�w˧cj��)���NTFS��d�)������I<L��S�_��� 6hpv���{>����5I�Db���J�z��v�@d� �8ε�7�h�~_�#��#� ĺ���ċ����@�Rn�$�u�8D�5V�/㕆�n�4�\ N�l-���V)I�mP���{c��>s#R{��#%kP+cL�Zy/�o8��y�1W�����D��0�<ep�P�J�NX/Py���؜l��u-Q�������B�-�r��ė.)P���u�XWm�;�?i'�%�L �S00���ԩd�N-�ƪ��k� а���_�������9��`D&��N�Q���7���W�`��L-�8U�ՅVρ�F�F���2�H�_P���&�Η��>,Y���Tȟ6���%�#h˃���u?N֧�/� E��UW�a�5j��S8��灁��॰0��&������9�V���2�(��E�=���[o�@�XH� k2�0���-I�����)��ø:��8?#���Dw���0�V��_��&�����	�{�,	m6ɭ�'ͰC�<�2�p�ΙD�;`��J�Z��I�"(�(�tK�˼����ǚ����� ?�\��wʱW�Iah��rz�̫к�u*�c'��;c��7��L4];O��H�M5�
��k�+�ڸ{�H�ʞl@/���$R�dUaΏ?Ym,�x[����Z�����# _����	�v���n����䧢PM���Ok(4^g)���W�i�
�WD�w��i[���Qc�gO�b+�鉞��"����	�-�
�^~S^��>Yki���\82m1���`��d�:ˢ�-��|�����߽��~�����Ӆf�U�)U�!��`=�i�z�	b[%/rY�b� ������ )+���L��_��,M�I�Z���ѹ�g��q&�[�B(�
��O��4n�K]�k���ǫ�am�����7��x.b����"�G�v�U{#����|����[��8���i^*=���v�C��[)���)��+;�}�L�C�'o��#_�"&sc�����b3�"�BGi	��U�����|lf
�D�%�asd.]����5�p8]q�{��������~(J�J��ı��A96�&8y��i��������\��9f�V86sRŤ�Oڠ��F��P�S%8�?Xvs�:�w�I�*qzf�.��e5�\R�Ɣ�0l��N�o-�R'O^���$����4�;����D�a�/G8	֡e����m�5A<��r�lA�� ��_��>4�W+l-��"Z�9��A)S�V��B�Jj�MI�7���30���*�y3�#7��__l@�[��bD#J�Ѵ�+�'�<���^F�u<��h�"�3���?�;d(�]�V\p�1�7g�л{�(I�b�b���b��$4�F��P�� �ժR�{�$��6u��d���&Uu�Ug״|��qW�KQ �r����e
��AyZ9>���Q��%�����㹿�E�[����C|fU����^6�n�<�7sDJ�r4gZ��ĄSY��.��g�3䘝݇���4�u<\��7E��4�ݥ���e�`U ����䨖�f��H\�z\�ڭ�+�?7�������2�b��U�s=���4��p����4�� (E�������%@�/�VxzI�.8.��}��%V�7�j(�:�`"0&6&;����Ӎ�SS�)�E��+d�+�lv��>YrH��Ս�>��e��m�]�RD�<��@��)��,-<���~�y����;-��V�1n�ucCa��`�U�1�e��r�\�~7ࡗY996xK��U:��hL�Ƚ����o�9l��S���+5����w�R�Q�wa�8�
�����ݬǬ�8�*����
�L��Bo���=�';�H�������jII�Q�:tÞ�
TP�g��]�`O��!���3�{y���b�0AǄ����ɝ��rL���+�{����"��
3yR�-�h-�	I"��^A���� ��TMVMIm�c�!��x�b�k�k�����k�����3>�R���b�Z�cd��Ҋ�m+�r~�8�U�*�U�"��|���Hz���'fW	j��7et�}��3"��@l���:;���x�I�q�ؔ��2_�qp����.睄�<,dx��S��������U�N�o������Af��~%A�����x}����;�MN2.yg����r*��/��נ~� �U�w�~�/)�ޜVzW(�7�M9X�S	���F˗�&2��a�� ��b�etK7�Fj�AY�Ʊ�M���ZuwU��w$\!�*���u[�^>�87k������gh�����2eN
�@Kj���~�ڬv���mM��;P�_���Qw=ȕ�އ��q�)�_�Y�����������/��zU�,�!�	K�Jnc��F6D,��w0�W�k�������R����l��yVn��ij�T`R�Λ؝w����R�_�>�?wU��dZ�O���xy��1�����R#l��K��џ����n�Ē�-�=�)����f*�4�=�Ov�p���@�2�
��;�j?e1�nh�q'!����vߊ��}3�*�q����9��
�HxXM�Q�#�G�@Zt@O���@��1r�b�z�b����ld�dd�	.��x\0�'K6� yX��W�\&K��a�g�&?��K�0蘣��}���I��K�{zjI�z�bz�jÀ�6����"��i���",ꖸ�dcN�Փ�]g�9%�7�栢
3
R8u��m��4]��ţ(Px�u�i�,w�gX�g�v@cF~�����R��T��Ėj&`�D��G+�N�D���\R�J��ٝ�܉{ґW>b����z�����oIjG7S�2mt8��/�Iw˯z�ՠZ�
�d�u^p�؍���Xa��ed�I���O�HI�,�k���'X���������vF�ė�~'���Kka�;	+�1T2������`j�>��[�9*�>~j��NE��9K�N92J6�������dȽ�J'�fA,����;�i����]��j�U�X���W�-⼥c%�Kjrg8&���hě�HDww֎��Ru1�`�ȯ#��� rX8:6�^�a%���$�/T`����fG��]������W/yG��-H��u�]9+�l���d?��)/���B�J-8u��� n����K�[��(�ݒ �;zo�:�Y��/��g�6�G�%�:��נ�S�l���-��R�-��"`[v�ը*��m`�� ��Y=��m�� Ƕ��q�W�"��?����(�S�we���B16,�c�N;+uZ6\v
�A�R��y	�F 4�8�ɦ�Q�� ���b���N���32�}��XD��2_�~����{ϓw挞}i5��c��&O��wm}^��E����Q��MT�U�6����Kn�,���Z�ti�?a֘�}�6��[��F�\�H%B��5�Q[\B�?<�T��I�f��G�)��������]���e�l*�/`�Su��]HP�����ɉ�� 
������uɖ�� ���^>;������H�ة���
#�a_�
ޖ�Lr�b]]ۢ�;0��H>� M��!Q��n�=�H��S�D�[]���% �O��|������C8EÃ�+�-��fW�xŁ�jݚ�q��G�إ),��;��w�y'���An�|��|A��/m:�c%�Vک����E�����1W�m�}�/�V�c� ���ĳۯտ���(�]�n����HS�toh��Y:��^��\K��kn�(�U��:��|���Hp1?�>0w��4�{-�Rп!�C��g�|����Q��S����>�f�(_���[|z�㞴�u��T
)j��ku=����5Mp�2�^4��;��w6��,��1Ͳ���m�#�7���3X4�p��g��^�I�21jQ�vK��C�?J���-I�Y�k��'_$����6"��}�7^��L��݈�؛p���i1	-�4����g�C+���b�w��Y�e����ʨ8�,bcp�]�Y�8�Q�z������Qu�?���g!t�ZC���*1�����zV
�!�C��ϗ��T���|�C <���l��"�q��q�&H��>�:õGq\��%��\��,��,����nE2Kx
_�pE(�.��sQ�
����qR8̄���K���t�Q̯M��=l
,�v��N�'1J���Y��J��J��g-�E��{��? �֬O�Q�	�/��8��Z�eD���mMd؛��(����)՛;m�E�N��Ɇ�c%����#��g1H�>)�al�M����̨��/5���������t�Z{�۹��a��> t��p/��H:v��D�&����ֈ� ��	z<�&���b6�Y������sI׶�c�Ha��┄ߺ�'o����+�Hs���deW�I�� �mf5R	R0�f7��A:�1|�I����L[�\��� ��*� �f�}�Gc�XOm����/ZT����H%xAd�[��7*�AT�����&+Mٌ��8 P�6X��@���W廭�*@�CCv��>w��gRl��2V򃯛6��ħ3�O��=r�-���j-L	'{Ɨk��	�/�_uw�*z��9q� `�+2�����r�q��O��5~���' �GIǔzؽSJ�hX�ux�t͔��]�Eؚa�:e�uO}�N�Wy� ����d��5B�6��R��n^��u��Hx.�˶�$sm�i�l�����hTI<\�����WT\Z2ޑt-6�dJ˼�����В�]�F�f�?��O*;��W���n��d��#�`񲛹�N�K���qk�z�Q/�>�1�Pz�O��Ъ�$Î�K9k����QP-����y����Z�.!���T�~�N��&�1��&�`{q�G�1u���rհ�����h2�r#q)i���&�8.��vp ���P��蛄��R�+�JP��>D@C� �׆�񟗀C,�W��0�
��G�����O�M�>a���80���F�w�����/B�]2���m����F�B���~�J�Ƀ�+��Z!�'���LМ�i��hoV�� �B�E�)�ő��u6�;8[P��΍�[�G�rv"��?&ܥ]}�Nf긮jV4�A�䵲UA)Y����C��o֦���n �j��i6<*���P�����N�p���qb��=]R�ҶR��Q��^�����q.+�#�v�PZw���#�}�o��r~�ޱR|q�ѽ��dc���̆N��!��f�����������\��`%:��tG�s\_��������B���8w����pz��pr&&�y����QR"{�Y�"��>�ɞ������]�6��C��"�u�ِ���[A����hl��N���给מ_h�)�憁"]3x����7�(���Q7C��һp�O2>���fd�g�UA	@�,�I�i����%�G�A3�Z�[���;�cȀ+�|K(��Xx�>��E�~��+G��&���\�&����a�����W����O�W�n%�����o����d�'9S<Nd�^0_�����T�{�F���_	6�s&X���F�7�c!�J��T���[No�∊�];��
ҭN~L�H3e�W^8��F��iʀy'��ް�_����%�~�|̽��~T�����׽��C�O� ��0ؔ�dd+��fz�p�*fj�>\Āx@Z�k��q�����t�����'!�r�n�\�HpR��P~��a� \T�4�f�~p�V�6s���8��NZ��-Ȗ��x��I��)懛_%��2 |#s[�K��h�I_xq����Jn�,�
�"���T-(��.����抓�0(b�o�N�DJjS8�(O!�B�bf�
�B�����¸�Pg (6����x��͠#��!��@����SJN��"�ԑ��[w��w岪��� ��0�5o�a�7oiZZ���I*<�jx�ߐ.��.�,7��V��ɮA��w���nw�>�%�J]�r�(U��ݿ�R&���������|��8:I��ҫi�l��q����;��zڠ)Z��l�V�?_����������t���39�79�㥄�}-~usǠ��vfv��|�X��8�Q�7��x��pf�:3�'�K���AA"��zѩZ���I��+�܁��C�����q���)�`���� �)���q�;�#��6Y,3�T��sB��s����;
�V����'+嵠�.����?����׉B�������X8������C�rf_r�6������PfT��n�ط����Y߯�2�b�I7�*�0<(0;�<�gB�9�_
	P^�L�[&���5p/�p���X�=Xk���ĪWxuE�w>�4|(�!Ӝ���D�cJGW�g�lJ���fLe�����֚7dغ��~`&�:8��=���_n���Iq�`eU��ub�T��B%���I��+ǫ����O|/t�i4r�6D�n+԰UK��`���G�A��x��f��R�mt���}�?�q'+c)�
=~�D�C��V��Yv}c'U������ꡙ��!h�*�bWkS���؜�]��TY�R�U�`R�]v�V9�&g�׀8���K61p3�#U��5h0b�8s�����~�
��:Z4\?�b~Q�ތ3�^�`㰸�� �0�_�!�V�.dћ��H���V~�t��3�;��Q�E�Ӭ {�V��~���'�>�ٯ='\d���k��:��t�in�V�`u�`�Q�F����W|r^uiS?h�{M"=?�n��u��M%L��?%6���IvyX_^֪-+<�Ī�zd
��x�k�V����O���}a�͆�9�#�n���,Ic�g!�L�8v��C	�^�yY�/	i+�8��ڞ6]�2Dq8�å)�JOtS��8�w��p#��H�3��`"_�O�L aN��6<�]�w� CB��)\4N�j2>�Fv��G'�4���lq�<�!���YY�iH��;�N��^
�3+�|��͇Ы9Ϙ���Q'!vq�P+13蚰��v�EF��#U�!	�A��T�I�h4-ϖs��}ϥ���b-~�m��R��^�Q篘����]�����-;�j�����b-����X���s)Ȣ�R���hi}v<�@U$м���gc�#M؁�Fe4��x�vd��.9����J��M���[�P
X$d+�2�� �ʛ���Ъ�W��+��!O�w�E���=�[UZp�;�	���
�['���<��\�@V���BnC(�d+�P��;�E-*N��9޿�	���;�&v!f�\��xA;�� yn����+/V�ۣ�郀��{��*�0�m-Q������� ϬO��ET���'ht/Š/��EB�����Y!`�����@��P�XI�?��a��AF)���^�^�׀��9A��ϗ��m�E��]��d����Db|UM�:�����HM=�Q� ���v��[F��]m)���;HdW�x#3ƞ
�g/<��j.OR2����%���OVbV��{��s/.�dA��;v������'_�vE�=��bƤ��լM5rEOV�]8.���f���CBC�UN�B#�z��3-Z��؉wM˭d���O��ˀů|�}�f�[�Fi�O,���U���#�u��0>]��S� �����[�e��ݿ�ℕ2^�t��(�SP\��@)g���QT�YP��e� � �AA��Nj{a�)9�a��=�S��>^Z�X*�����m�BN�̽`?;:^�xH�!l+�;����&5_^d��A�_��[̊.N9_D�o�t�*��^i�p�}�����!S��� ����&��c��`�p*xL�3�%��*OS�U��jlf���3U�C�9w�`����m~m��n<���ݻ�xZ�l����s��1h��-,.Y<�Nj��8�r���> 
�M�y�N
3�J���W��MSz����`��c	;����&f�hz��[�ʷ3c*�?�f�DT�b�M�v|�N1R�M5�XTL���/^��y!�����ܔ���[b$.N��؀�Wr*��ȸ<�(R��U*#��;�[�5��͂�	+:
�Dy�8Q|�
\��%ӺWޜېP�����)A'vKM Cr��m�)eƘ��Ûi��g��y~Y��]�o���뛁w�ï���5���?�� ���5$JfT��M�%�XJ�b�.6F��!
�iW��k]�ҫ}r��@�f[!|#��lZCXK�m~��4e*Jn�b��,��^�N��,�XP �s�l[(�T>tΎrM��������M`,�)�N�A�s1�<�A\�8��5?1�fp�������Zʉ��:t|s32ɛ;�v*L$��ז�g���`}�:�P�����)a暩�p7b�+��_n��trJ���A
��5{x��#2լ��+�N�*���B�ꯆ}��]�tF�j�6(j٨��:�}\�Yv�Ͳ�B�g�WjM&�^(�BQ1I +��g��!�K�Z��<`�pH�0O� |s����ߴ��	2.�`�.��a�p���)�\)���0����qV�|Q�����d�D1�����QAdZ|]��0 ҕ���iq"^�-��K�ˡ������'��]Y�8E�WFj�1 L����wA\��&q'���K����p@���y�p=@�%r}*Ð~A,��+�]��"���͂�+���vI׶�.�8sS�����4��P�e�z�������e�)���A����9����,����=����F����<wd)��n�TJ� ڭ��b8�.�~��{�1�/d!N���E���$���9��F�\�&0�zu��B�`����T��i��9����j� c#4E�4+����*���f<҉�3�z��+,_܉�+�r�{��*r�8��D��6\\��:�̺C�U��.~9ío�o�eP�A����Y%�Ŝ^��G<Q���1\�k�Of���.�$�����ib���d���oe�+fC�\�V��Yk+�b+Ґ�~.�z�#AȠ�����<)$F��T�T�;5ON�PF$R��H���xΘ�[\�zSƪ�B>��!�<�J*��	�]vǡeÅ���Kt���d��{��=�@C~`=�h8��?@Je��m��L?~D��0��=�V���7�d̖.��bg>�p���B�z���}xE�̒m�EN�8�U�8���V��1����(����`9�$�����Os:�Q�g�@TkP�%J�0<���'D�4C� o��YUf�[��fh��Ae+u�B"*�fx����ht��.M�s�<k�[�F��Eic*��$TÁ�$\ɥ�/��L��luP�������:<�u�����tE��%�3]t=?�i�Γ,/$աz�ӗZi��p�Q���%��E�nK�J�Od.�T��������*�ʅ'�٭�b����&�c�
����}�s#Oc<�����6_���$ֻ	�I�3X"��� 5��ʫ7Z��u������a�H3,�<������3I/��h�d�,�e�fU�je���k�Y�M�]�f�c�Ј6]��jpIʠ����U�������mVرT�熆�V�rK$�� �c�0Cf �ԟ�)�����; 2��o��{Ly����cx+�A3k"}V@
�N���?�(�xOP*��:G͗������y�\^ � X��2� �}x����� ��V���d���J��O�i〖�������п�9�.S��攡�`���������q�"��4�`��+���.�F�Q
L^��Y�N�}>��?�z��%�L��$����i���ɏH-f�h%� ſ��g���ߌ�<��g�/�cى�l�b���njpr"�Q8%�93�<f 9�uY�����ƿMstt{����>�S�愬eI�h3Q���R�L���M4'�v�?����3k���2G��J4VoP���g�w���We�x��z.�Z,c�KJ��\��;q΄nF�Ɲ���Y�R��$���:ٺ�
iJ}��s�0���7��!}������Tv��ԬP*�s����mȠ!���"��i����~�Xď���C(G��	�����l�_Z�]�%�$Aj�:��[�2Ľ��`�P+EM�(ml��b)Y��Pg�prVC�q�Q3�&�8�ݓ���\�qo��]'�8p7u�0�Q�k�l�H�����7�ۿ���U�'�ĺ�ڤ�T�(.��O���L��3�mR?8]j뜍h��<��Ƙp>���O�`[�K�Zy&�G�I�tZʕ��^}�lO���;q���p�s�\�@�6�[:�{4�ܙ�`���K8iz	ud��Gl����䉖i\�,+��!l���ͽUau� �߲	l�H]!��*�}
kN�
����4�Sd.���aeܿ��Ͷ%6�� �B���ѢB��C"��b�o�z��ur>����cq�e̥=%�X�(�C&��3�	>I�g+d���TM��v�=�ʉ-֪��H7��(t��9�H��ꮆv�++ɫ��v�+. ?���bW��b�(9 ��C����e��'$��O\-��n��d��A��^�M8��Vv��J�)Mс2"H��V�yn{4�4b��=�3���
v�f�?O�p�A�j�R�ݿqhM�*�"�ìxV oA`���;?�g�W�Y��_��'��y��Py�%�E~Ŀ�`�+%��t ��#�Rw��d�F�mӞ�Y!4�2�=�uqFo�O���]�(�Ӓo�_FJ)0U�� ��AU���v�wm�4kb��"t{4�X3�?I�����Vy��sQ��Q��/��/��_q�{��iZ��%�F���	��t��@���>��8��h�k���5��""%�Pl^e���Qo�^�2��}<�D\;�<���[�Y!v��^O���L�Ps���mݪ���\&�5# Ƴ%en��_NF�jס穀fR]���υ��&���������H|��T���llC��rJ��U�M��r�4��YdDOp�Y��w�xh�9$��cT����m	��9ag�\B��N�Q
�F��{lG`�X&����Ee'a�4q3�Z�ˊr��N��h���X�.�Ɓ��7
�`�3�&.��9�uH|���Ze\���*�$�2�*z�\t�,�:�t����J���*&.}k.������RG�V���dr�A�~�j�ʥ��~�쮖p����@���̈1�����Jnc����!���-����r/��}%qq.)�^�h�ZA�b"�\c@�"�$u�B��%XTAel��e��w+�l|��eX�����:Q6���;�_-o��z)=v���a
��	~?;��V�8�e#���/�P������f b&g=�D�u�y!��湉~��х�:9ڏ��ާ,|u
t\Z�2�y��3Z*p���0{%<K���q6Y�V-�'����b�iq"O�@�,����b��\��x�&�N���ka�9q���ц[[dT7���q���
ڝn�~�G�NA�tnؾ6˙�}�����<�a���U�:��鞍aG���/�>2���t!��:̝T6��p�<D �s\o[�c��	1DLƖ,��.��97�:�Ȯ�'��|��&!��b�A�ʥĨ�JdW��+�W�h�����(H�V���ZP�b��1�Ws;������V��VyS���.�-ˬK���a�TW-���	�	T�a�Иo]��y�|��Ɗ�}����� t~�=g|{�m[��%f\�x�����WP"�r@�հ˾�4P�8�˶Ӛm�C�)d���.��j��C��eB���訠`5��I0�zDIO>~_�~y��A����{-N ���D2��M���C��4^(��G�Ipd۪7��p/+�\U��hr��w��fH��La�=!���܌�\Zgp�V���@�{ ��ڄ9�4�H�.��KE|����.����À;�O�	"
�d��r��5b֥�ğO��~�'q][�M	.�.��%�{��3�+�� �a]*�����1�%�?z}j*���$�R������DR��@O̟������'�����4���T���5#L���2���o,����n��aaǥ�2�����y�ء���ۄ����.��=�[B�|9������n�[ߍG�p�aF�up ��j���ݮ��䣽�`�b��~2�i�P��c�au"	��Lje�ӯ��yd�^P�1�@g�(�K>�����|�:GтM�&#jƽA� *W;���+��"��=*�)����ȌJ�l1e�#�R.U�f#�b��b�iٟ��"���}��̨������P��Ƥ(���4��/��U~��e���xt�����^-�0�O@�ܗb����P&��6��� (����*56@`�\�iӉ���z!k�O��57{g[���D.�c3A������[{o�L�7�;,�4Rädd�]�V/�1]�>��]�.�����*����#h(7��B���`č�O��"|�����a�?�P�������]�1ϥ�5*�w�� 	ɷK��~@E�<c?�F��{Lj%��:X�Za!P�!ƿ��a�J�`�v<X��&Rᒓ��	>��$��W�"}/q�~Z�h��?,?x�so�X ��a������C��;��Enzӕ�U�����.n{"k?�"pVS��A]��Bp,���R~k浅�)~/�D�^ein+�7�;��g�8)��ۆԛ^��nh�-����5��U�u:��U��0	�LHA�=p�g.�4�)�*?��R�0���-��)���f<90ֻ3F��d=~�7E@j�?D�6�p����}����ȏ��n�����%�|�}�q=+����%�o�$�
d�
AS�Ι�]�Oa���y6�O%0�-�6�v�^��;��72#g2[�$ʧ���·����W����}�p�p����'�17�D�R���w�ڴ̥wӑ�a&�z�� `����뉚�ầ��UK����^u8'�/��F�q�Pb~�Q��s�~"x�ԏ�{|�%-8����� ���Ш-9��s[��x��s�אz�ڡ��H��U���b){�M�w*���i�e ��r��~I�D�L��`K���Y�m��gPpT{a���&wQ�"G���W��>좚&۹|�J�ȕ��v�܌X����|s9�D|㛾^X?^�XC�6�E�Ew�܃Y��>9�}��ʓ̝�u�j����oӵ ���nN��R�0�	�<��K&H>�{���"K5����fCf�����.-���n�޵۟�U�κ�nM�u9����冀�k�͑���ń|�}�r��H��ْ�vJcj?�Gl���[�����%h�dq����֊s�w�G������%A�s��q�6���=�I�̥�%d�+�4`�_�ǡ� ��*���hݺ�
4���|[b�@&!a@t9Z�qX�L�ύ�O [1��\>$`��P�-��A��	�{Y-&��=��om�����	��^+O}����	<�]p��BQ#$�<_������k�2C)�j=��Q|7:AJvB��sL�Po���c�3+�"4p{�����E+Jsr� [,}�Qr$�������w9��h&jQ~��Z��cá�u}��w���r��BS��Q����Lλ�,�N�P���d
~e��Cv7c!�%�Y�硙���^K��Ԓ��u�5}pgf�9�NX���?}��0�TI�|C��k:8���m��ب���/`y?�~�.�chKp\�1�i�M�u#YDN|�zyb�ē3��P���ׅ��z��>j��⧑����[`��W[�)=�N��|������K-#��$���PL�A[�&"������5y�Ѯ��ic}��wy�t^3�2%��f�GO���i��� �|@�����s�"�4��5[���Ln��Ԯ;F���p�(w�Ç��u����hO����s��eq�>���h5S��}4쓔rP����Y=,����d[`�V�h�y��2�<+d��L�T�"�ͧ�_�%����^�AT�?J�\�f��J��ڶX��� 9d�9%�a�GA�sf��z @��2���ACJH���W�o,p��G�;!��I��f���1-�QX,���rM+,@�0P�<ts��tO�)@&h��f+�rGU�Z�c���ny��������ړ�����ɗ`EP}��`�R�T&$kV�}G�ч#���iPz���ӏ��}-5��������r@:�dDJr�	���,�W_'B��[{���[�`P(R*G�-�=�[�CDK5|�����)�{y=m�q$���>���t�KNjЫd^�'�i4�V�	�8���@�<�.�\�^ n�{L>^>�]_AV(8�v籼�[:��_��x̆�<(b�O����;Dn�P$�g�d�h�;�v�E�nρ`�-l�eaAbv��9�zx�x�p(~��ps0H�ljI1un�����>L)�V��,�5��L�)(��_��r����И��>\n�o�B��h����ы����ڂGp]��fe"�K��˸�܋+1ؐВݦz/�c�]�z���< �=x�����ˆ�Y��\��@��`��7���������p�{΅���,��[QfIQ��ZXM�l��{[K�D��ƴ{=�O�P��o�=*�y{O[%=�NA����2wd>Ǩ�^�#����Hf��3ʺ�<�tɂ9w�� 7�:�ZR� �VH� Z�bX#�n��'d� �'���k�V��\f�J���榬q�,���9�ޥaK�AD�UT d�-���|��ٗ��nY,��k�~B4D�4;��������a��e��������I���\�k{�D���i�X-�Bf�vו���po�W_5%��W:����ܨ�%�q��Ok�zu;O�~�)3�No�S1VR�չNj���&ar�(��^W��NT��-]C����L��F]��b0:��lM���%ŪT+����[�������]p��`�P=�Sc{9˝Ǆ��Z؛Q�ϒ�狥�3k\�M�-��Vv�nX(�#�-@2'C�<�a� �Ta� �{���	�>K�!�O4X���=�oa��ޗ�!��PHkXfn1�@7�hmB�Q/Sn�`�nM��VQ��p/�$�Onp��<�/%^b�V�P.�RRrŮ洣&.�c(^���a���NϠ�#$�1k���UN�\=Qqx��2<Ļ�ĞU�o�������,�.�Y�U!D?�1|v��mn�-�VƋN�@����o&���-�P��������� G(��A�MO���ƧAp�	W��@��+j����ߢ�

�U�����+�}�὚f�m��W��4�6z>���q/��`�1��dQ@==�5&�gȂ�-^JV�8 ��!@z$JW?��������]�*˛Q��&Y(���]����y�����2�,��2u��
��R-���_��"�g還J2�E
)�����-qbX�1"��^�q�J��@sL�K����U:���~ŤQ���})���Ȏ �ә�h(�ڝ����Y��y��YZ�^Aa�N��;]�6o���q�*
�	�?9�H��6Hȗ$'����^��i=����������t��t�Q�l&�ۥ��1:۳�u~�.���[�Q�8��7�ފBP� �]�!e��x��DF��<[�x3��f�"g�ʓ���Ӑ>C l���Zi�Z:�V^��a�gA�q{�<cB��U*�/��Ӏ�J���GZ�e>'��*�m��I+Ԩ�fU�.%�6�K֊NN�T���8��\�sh
4��Hg��S]:�����Ŵ�؍d��~��M<�F�/o�<�4�l}��r��i�;JH�E�y�2�)�"V���}w���zI{����Ўby���α��g�9�I6�A	(~V��y�8�.}	DgS ̞��)(�?X#�ǌ����G?�D�\hɉDs�O��\��	Qc]��鸅zR&���2�{s�����<��]!�����
�����
���Qa�W@-�dVi/@[�Y,J�� �$"쳤��+�};�]Ԁ�ࣣ���x =��g&���o��<Kȯ���F9HOѪY��%��F�j�3#Qk�]XPw�uUP�d��z�KD�{����y���m,\�ϻV���0	����y�k�b�B�Dp���r�N�4�37��(G��B������O�-ߦS��s���O^u�l�ؔ��m����)L����a7�O9W(?�3n�Ϛ-����U�Q�聘�pX�!��l����?�ȝh�g�?��"p�����,z@�خ@4ߣ���۠��!��e2ƞFK���N�*�5	�g]8��-��G�֟�:��J�:֔��<`[o���Z$ A�_6'y_��]��3OCvQ��"�3_�Y6W��l��!�ǫ�w �8:���d�C�*�M�L����ꭿ���id)����}��E'��,R#[=�3���B�sd�[iKӫ�wb�^Ҩ��bG���qC����+�9�����V�
<;~~m8M�a�>�D�9�Uޜ��1�~���IO�
%�r��;~�� �_�T��[��Ы&"f�4
��L����p�"�(����-FHN\0<�9bϸ"����5S��]Үj��;�� �& KN���~�9l��%�+n��=<u��$��6�4(F��|?�o�(��Y�K{���Q��2]�0 2��bw0�r:�/����3�g��Z�䏊=�7�.L� hm�Ы;�y-v�dSKj��~�1����DqHe��<�?=�ud7���`�b�������YyoZX�̧ �&��O,H1I7���b��|�\a"��'��+�!V'��F\���Vư��f0Ѵ��&�$�I��Z��i�Q�4�S���=+�&+J=C�ܛ>���x�H��߷j�+7�NUk��h�7��o�r�E1��X��Nu>�]�JT��x?��}�X/5�.U���\�RJ』�Aҧ��@�/X��V�����S!z����_W�[�o�s�(HK�c�)_���A�G��q�u5S�*�����b�{<����ws޽;��=�H���ۯ��0�U�s��7�	�����4&��'��4���
��+�K�.|�eŲ��[� \����U� @Q'O` �k*�K�9bI�spRO.,��"2$�h��n��DAPo�6��Te�x׀�ܹA^���ɢM�T�0v�8�G@��Z�:%�.$�uRqz�~;�)�Y~�WeM찆�LP��@NK���`q���B��2�WU�c��|�]�,��<Jc��@$m"��zƇ����q�k�s[S�wWg�P��>���Lx�������r� wi�P��)h:�*��9^(�fm���1�.KC��\d�)�x}I�i��jS&��?��?�
����k~��\�#wִ$F%H%	Pm�IZ/rF���,@jg���@�0�nD��)�O�z ��|�8 ��1���}l�X�����y���#��g+S�͝u�+UG��V�yؘʺ�k��v�/���_Ch� �S��n�Ȓ�����A��!����U#�i�P�n���lw%T'#r	[O���{ ��b������eb_:W{�O.0)H}dPN���_���W��� q���Ke�����0��]�c1�WE�����J?4o�q�`~`Sxp��S�@�����I�����^��g��)Y�	�]��/�e�E����fU3+E���Yl+�+F�)l�|!��!Ȧa�+�ia�c>���9�����$�o43	��X9CE���/�xNϥ���o��i���mH ʴ�k�V� ;R3۠����1���C�O��՞Ca�p04f�h��ˢ����+�-U�$��X$�����fv��p��5)���&Dܾ�S�!vv5Ak�,�!�đ���vW$1�H��S�Ug����enj!�:K/i�q��ϗ�i�ś�5���i<7��޼7.��C�P�A(�j��0��Q�����j%�����y��h$p��u`c˭�v�B��>��G�i"�C��w�������C�dR�#c��A{M����<+�(nU��~<J>3ֱ�o��/ _��z�g���M�Cw7�}�+�����= Qמ&�����>`���ݹ�V�5:u>D)�hd@����Gl��7Ec癨�
��K��8Z�� !.�:p`]��E��SB6!UBS6/��;�s�J��ǭ&�)n�I�ŏ�v*j�����lLLQ�Cť���9�����������4�����S���)�)��u��OX�$1� H�T�)#�UX��Uvlӭ�y��;-��q�[c��k6+��ɗd��|�J���������%z������\JDKFK�D��"o��.M��+U�±��78b�R���g�(h���6���@�FL�/ ����q.��A���@*F��%;��1Dv��6��|��u%�TGv��A)�nc{���2*f��ƀ�;�C鉮�MQ�鹌��󴽵��[A?�4+��H�P�[g	"�L�x���i����[�m-��(�VGYYM'��u���Px�G%�388s�L?P�D��R�SK̢\��L0[.&u�{��}����/���:����Hg�7ql����X�����WS>�ȳq�#;@/!�u�-����;�_���o���6��V�^��b��U�@�m�UV��5*�Л�(�pY���K��]�K��7��U3Z^�/C��T >nM��x�h5�9��֗%:����$PAw5��z�RY�-%�^�y �{�&/ ?ĵݶ	g}�����qMӊ�h�O�(=EV�0����A�?���OR��Zb��q��j>�ǰ�U�)ն�����7E���ԫ&i��!coQ��+#��h�%%��0v�|��bPt�JGDTܝ��@��Q���#iV�*î���jhG����'����D\b �EnC8Pn���C��������^p����DO�|��Zod�.�7k^�a�\�Ko��D���B��\rQ��)����}�f������A
nV�����C���hI���z�)J�)�����cX>�Z^���%�c9&Od>;��(��(r�K�0*���Tݳ�-Qw7X-���7�����lɹ#1P��F�Jo�c��Ѕp8.&~Q�,��uX�~Mf��Y���!����'���}i1��CN�����?�X;�!�I*�9�J���GؘI�Թ��Oh�ӠM�)�>w��X������n�X��"�NT��� �$����ԙW���3�����]�?�]s,�7ۍH�P�e�<^ j��F��l3E����[�j�!�Ք�L�;��\jǝM�Vp�d��x��y����Q���V_
G͸�z�`dڭ����kq±Gc"G0��)�hj0V�EqH{���u�,���Wj��E����n�� ߌ^x��ԉ�b��<�W��=��O �k���8 ,���ؠ������jhn೻��R�8���|�(�������/�DR�b$�b�Z}f����3��v�IH]���๴&��	nZ��Ry+|�]��RЂ�� f���ws~��.�����˦�ত��ni����ɬ)*Oɑ?|�Ւ]��?v~������0k�8����o ��3�qo�1���,Ud��'2����R�`4�z;mŖ�T��k�X���U�A�s����N� �G���Py��&�*=�N�� �n�U� 2fK�h��Q��V}k�y��b�� ��T>���;�ٞ�s��lO��쓕q@��^�9�a8Y��,)"��W�$�@ 9L�n]�M`�r��шS�V���xA��ޞ��Pv�|@��.���c��b�p%l)˛��]�Z�ۂ���V��2����ȉ)�ޖ�6}L.�Ta���aI�n�ۯ<y��;e0��?!�+��<�՘�݀��)����� ��QpJN�Ē�X?!�Z����@i�j�l3���$�5���
������~�F@P�Y�N�ڴ�@LCo5�yl-�u4Q�/{�����ni�ip�r�l�iX4����Q��y��������\Ԁ�P��5s^���2��ɑxh�=�� �Y�2�Ua�rj��m�����NjԓB�� ��	R�z	O���K��F^����z�h맻#9?�Q���2�/δ�<�n��U�/������d�\�8�ș)F�d�>�fg	bhizO�pD�R\��L0'�5g��dƿY�����7�twh���@k�=X7���7z=��ޅ`;�_��*�f�7�Ю~�[�<%�3����%㸕qW<=]Q�FH��5HM��8�3��"=�el��AE� -�F�0�8;@D>ݍCh�R�fQ�Pk� 
?U��U��L8��D���H����?ԼS�����j��iਾ��6��W6 ���ز�����)=����7`�U�9v�� �C�)�'楣ۑ�2��淦�2#�M�Xr$>��� ���L(&m�L�����������R*z�=����R��vG��T� �M����A>�7��wvL�#�C=>[�9ב����A��()yF�G�F��Թe�ck��|�ڑ�iū�й�� ���o�,��{��\+Do+� ���-�άOW C���H��+��NF�1��!��>Z���H�>';���J���ع.��$�(�$wZ��ip�X���}<Y��H�2��s����l�+�}nNr�s=PDCe��7]������x��#�՚U1����43`��ƪ�+�i��鉎,�;U� a�� 0߬΢�� ;4�k�/XFX�p�j^7���>4���ȇ4�RUw>������w������j�����\J��Wj�+{i�k�{4����L�[s�⛈i{!����y�0&���#(��j*������1�к�z�$��z�#{ð:[2������R���&|�D4v U�ڵп�Ы��3�5�0+}cT����a�m76��x�P�\hTq ̓��t�5t�0a�c�]�ze	X�l%�L�����fDȪ��� ��
�ɦǤ��|o�K+�N���
He���	t���M�2�Q�^@Z���U��Q�мw�ff*�'b��2tQ���L9�r��_�}��8ha�NxK��n�`\[�q2ڄs��9-�>�9��7��}`gd�p�teq�j@��B�Z�a9<�A�d�w���	 x������'����Xm/c�gGZ��^��t�+��ث�A� �v�2!���=SM��w�'zՌ���P���8�L���6�����jvX���$�p���r�~(%ar�(W��Ìz���,��t,�,��� �����L;tT$�Ʒ��p�i.�5�}�t���BS~����i'�4��#�*�"��g?��p9��[.{Y��{2x��<����5eNW8��Q�Nb��19�q��׻K�l���x!��������C�����Qץ}�@%�Z�������yd��4��z� {y}RM��>�#�G.���نs���hg��2!=��4�ݨ���0m�L��s������w�1w�h�6��� c���MԳ=��vp�� �,�	�E�D!��4	3Z�BOL?zv�<�TD�N"Ug��3b� �nV<�k���8�d.ۘ܋�����=6�t��[�\/�L��N��(z�V^s��:h\jC�J2"��z
}�p�I���a��Dt��"z���y"��֨~��Qԁ�TJ���gS�:K@��?�pDJ����g;��d1a�s$`��^�@�H| �(	F�)̬qr�Г������+�������.�c{U��jzu���K�N���/�Fş�E��=�Y��{�Sȳ@������ԝ�?�[�YgZ��C��Y3��]+�������M;:�rssi�jKp�*���lD�L�~�s�g��������A��>��&��USV뮝��?<��^��;ـk6����ƒ
Æ�͛F���߰�/O/�<���nb�T�c�3�Mr{-�����/.\� �Y}�Tɉ+�F4��X��w��$�Cy-�x���|���>E��Gh�o N���Uy��������T�Z[�f)��{%�D[zk<� ƗHCu?pPRT
�Y���JX~ƥZ	�骇�
O����m,r�;1�U>��D8	�f��b&#4FC���a<%��y���D�����,��~wI]�wL�ؼb+?[gFMV�!�gy_�XZ�e
Uo�ңV�'o�S%�`�ss)IL���X�.L����b�妗@]��k�'���>Cp0{�KLO��ٴ�#�x6���w���i|�������o��Ȯ�x%�w�Zh���R���@��
�:(�<�;�܆���^�cT��2�51��`X�\u_���/bk�~�}���y��7\[���I[7w�.��\���J]g)���]Ľ�µ/]�cT��	I��2/gk�xw�������K�	�������C�`�:f�|e>�į07l�:a��P��bo����:RX���8� @)H�~H�/M�P_�����5����V��cе�78��I?��a|�h��g�tA�4Z6a?ң�/�]"EA��4���5�{+��$��eǅTȕ�H:a�k�"y��)׋��Ё�%t�P�Z?���`�j�g0�eɞ�W� ��Փ�������=83�n��(��7���K>��T���>��]���a�'̹^{�6�qǵ����uV�4)���`m*j �IH%D�����bh ��5���n���n�I�E��[�'��5q����7�'�	����d����]]�WD)� �S������#�u([����,Իm6s`�ƪ��z� �`�-pjx�����ta��o�q+B[�7��y�9E�����	��Ah4t��A:���Y2=^�eV���ٖ�	��ZF�=vHށb2�6��/K�d5���CH�|V��5�¤�{*]��dt��\u"Pʓ�J�a�T���S�M�HM-%`�����2�{���#[dPj(�\t�=i�S��qE_����9�)�iG������Vs�MM,+�j��P�qz�%g����t��i$.c4J)I�U��w��@�/I�Fu ���Z��~��1lK�5I(Z�JQ)�=X@�(Z�)F�v�#���� �М��LU�3�����x��u�q��΀|VW��(�^�&ԞY̶���|*F�����?&"R�$�RJE��wZ�Sߒ܃T"UtA�C���__��i(��8�}��	1��ܼ����AH�G��#�"h��{�i��=A7�&��ip�=kE���X�����7md�������yq@��P��4�P3~a=�.%�\B�!��NM�s��`������-f��F�Il����}l��/�z'.x5���oO�ு
�s����́����x _<Np�|&$y6�%�{{}þ���W*�p�͢i���(�>�e���~����#��C۷���>��L��b���Qn>���U�]Z���P�#�?t�x�,{6���
���r��?��1�q��G�I?ύ_g�DOn�dyY�k��v��>��"g��9CpY�����[�q)��	Su+C�@G"�� �Y��`�Œ��×3����Tp�{_^�m)�v�F
�\?Q���d��6 {�av�Gtq�/��A]�9N��& 4?�ASc9��Ne�I1���6@��&�$U�����.�K�\��+���a�Gg`�ڗ��� F�����){��B̜9iI�����2-e:�^2,�����ט�as�|�֟>���H�/�y���M-Se��&?YEZ��,=�X����;'~2r��*������=�X~��wPR��"��@o�p�pa1�d��[�B8�{|�&��qV�8�pI�M��ʢsI�Ȣ@�K���IdRX�q&;M}��D��6��y
��#�Q���v�L�BoTWM�)w�U-A�������4�A�����w�E��+��rÈF4�8����'����{����ֱW�r�ς��]n�@
��q��I	~k� ��p>A�|�%��:��]6SnB�Z�!�s�"
���]��.YaʧU����v�깪J���	�/*Xl_{�q$x�,��� �|*���m\���էءT��~\�����M���� �nQB#�haS�±^zj|D�0L�=8��nم���p^;�e��v5�����1ƟL֍G�f���[i�w;��096������:�jk8�����.��C��Z��=�袻��u�E�: 4ʺ��"Cԏtt�S��y�v�q7�W�A^�/A�a "!ɀ���&6b��.�>;Bq����ǃ�����et�1��\�&S�K�j����_�j�M��}�o{տ`��逷褉�L2q�-5bסCa�Y�#�vT1�*�#����M_�"���R��>\��몁S�5�MԬq:�i�ٳ��o�s�b�/�k�^��%s�Ci�N>nM �C�eU�"�]�JBm�B�V��{$�T]HnN�^�3˝{��[:gM_sf��k�o�5i�o���=�ƇXO��g B��fZ��4��.�P"�Qڅ�l8n�0��#?��Vg�~��%]'��:��&*SX��Л�g	��c_���>bq���He�o6���i�:(l;�C��q�9'WNQs�mQ�>!D��h;!�b*i�����O�}5�4H���zA�����D W2����Vn/6��$�VQJ,N�P���y���������:6�D��_{`엩����N���F*�bܸ�[0�1sD����X�`���,�q�<�ҬqR�DO\7R@��Ԩ)�����C��?�ե�.����?�����ͪ�0a*�.���h.��W��&GK�Ԍ��u�]�m%��8S�X�"t�ӇA�\���Ѻ��<�f{O����vH�����.:E��T�5�$ŀN��W�G��H�+rL�Դ�1�u��݁����A���j5Z�o^��Jˉ�YC���w�!�AH'YQ_1����)��u��9;
�$���-�<WXS�h��9�����}-�y�u�j;{afl�f}td�y��;]�vg�5���
���~M|󽣾i�.pO ��1M]�C�7�>}����KD��n�ӌ�x�Τ�ۮV�'�,�m�ޡ�i)_�д�1ٕ�S�Ut`�o�<P:�`�+w<*}b~�:�n�����&gW�CY��gV��i���Sr�"H�M���Z�BrS���ZD[�
3�"�Tj+�P�x"�tJ�Z����[��E4�1��o8;4�2(ۺ|���U�Q�ى�'暙]q{�Fh�NFe�'�4�>��n�Ik��{;�@كkW���J�"5��GHrG�3�5dϝr_	����;�BR�3��3�u�Pt��tn�qn0M�І����t*4&An��4�,Z��\q�j�_c!��������ؠ�{ ���ܑ�x��ƌy=�}�Ճ�]��?>���n����o��v��mj�Vc�:� ��&�t��#�M�#g��X�P�LV괩]�����e묄��i�s��Uǚ�K �ڋ#�vV�p{K&\ۙMz|Y�ťG(�v���$���! ��T��bk��tQ*g𝰍�}o]�������%S�y�c��ܶLRogM&�����|6�,�i�f�E\�K�T�y��
��|<�{������m�r�LX�>v>�2���������� -���s%+�P�DRm�Ў�֛� ��3�M����"!�?Q��2@��?Q}��v�\S6�"j���.���(���\�J
i:Fd��aa5o�M��VO(���Hۉ��*��
+�Rd6]�yF��Z\��l(�US�c��̓]g��o�g}	�w�����n9O�V��0��@K.4�]�n1�;y�%���f��-,�	!�a�2{�I<���W��,M�홺��-.�U��K�������Q�0��P���=��o�*f7�Z|$7����Y;�8��gw� �i�@��/��C}����a �ˁ���A��\���g_ �ݯ;���-���DKv�!��<���~7ӯ��DGm�$��*����u�4y�3B�6{���5d]�^>Ƙ�=rUp1ɗz4!`�R0�U�TB% |���7��D*-r���7"~:��$�O���T�$1F�j�Tr�mG��]|"��
�-��|�ポUŦE��>�O'Z������*�g�5!y;s\ �!/i��vN�;����\7����?u���Sx-2,��r�!���������П�*����fW���b�Ǝ�U�3��Q$�gJ�?�:uTu]*�T���Se��F`#�I{rl���]�D�p�\�7��+V٧T�A1w�k������'�F��#8y*<���0s��H�*�Y	���<�F_����?Zb�&a�n@7�,�M�7's@k%�݈�����9- B���79��4f@�q�`2.J9��(��a�Es�g�7\�	��{����S|�vK�'tCv��]����o�uX�쯪��#�/�n�a���� �A-d6e�f�f���٘�0����9�E�7�c\Y#�
<թ��G��:���2$�-��&XxRu���0[�G����1ƍ���z/R;s,^ô�Q�Ӵ�Z��M�?�	�Nx�[`���I�L�j�����bl��l�z@�����ql$�^#�E���k�:����G*w���pc�UKlLm2CM��X"%�\��@��Ȯ0��~o�q�i�����&����B��uEI둝�/��.�4�F�)x��Q+��q6VP2V������oD;/+��̲�\4�� ��R�%����0ќ�+�U��)��U��W��'���.Ko���ts6�	�y�>3Ya
2�T�'�-E�џ��P� �
E4V2҇��	���ܽ�������w�ds������3;�D m�u�xG@��37gJ�#H���n�7VN�D��Ih,K�HW~(�r����x|�����x���gN3�@��4�n-�"C���il�����hҪ=~��0`�mM��۽`${��RF�a�w__��ѡ�����[9v"�+��9a�����WS�H��%*��Bz�ulq��A�\��5��l���&e"o硹QD�󕞒�N���2�	[T�Jxx&G0��W�!�U�7�<�_Rƹw5��7sz��aJ��9c��@ I�<{Of!�p�A���D���z��{�K�A8TM@�o�Ef8 �����"�)Ћ�NH�� ���o6�驒�'�PFg9`��U���z`�f ����Ş�����'/��/�Ǒ�B�r���X�h���Y��D��h���7ʘr|�t�$��nݖ�����ˉ��u��[��2�zrw���Y8[�[@*q�-+�B������:L��o��H��q�[���h�\�%#_,7��:��Xb��=]� �ከ_0q~+f:	dn@�y^;��G��E_I�*�_��>N&��1N���a�6<���Å/��0�]-�[��sH�0S<��@����c��pR�R��I���uF��/�d�<������J6�5I��]��|�p�#��}_�������k�f�W���A��l�<��%?�dW�/���qN,r�8��%7�ڨԬ,aD�U~���t�)P�mm�������gZ$�J���8W\��AY�������σ�F�N�x���������\1,(�j,���P �b��i���Q�h����+w�to��>�Q��Wv���ī���o��H��%>4�A��X�d�Ξa��k?W
y��q�v5����L_K�����0y;�z��k�{|w�R���.�W�i�B=r����i:AU������ 6]_��_�ˣ�n�ٓ�Y�KI����zɸI�~��	x�w=8v���)&��M�{#���=-���H�,�	�h�����*]�]W�/8B���A=�6�,����t��pg�ne�XI?����F�j�T�F�Z�v���Nw�q�iԣ&�e8�-A�9�`�� �����m���Q2�wh5(�t��v�H5Mb��9��ӱ`�g�k��z��r����G������lK~<��P��{��	.�R�}+��;�!t�-���F�d�Hi M�������'c�Ԏ�8�g{؈N��R��^�����ch�1�X,� ���Nd_~Z1�Փ�6{��<\-�\� ��������nF��Ě��#>Z��E�Tit��Ie. ��<9�-��#�s�]o�<��3Ο~o�W����&[�YKxMd�?(Z���O=Ԭ���U<����D8�K�6��^tO�Ȣ+" �K��M�5�M�a*��Ί;�dYEED��!�-_�gA�� �[OH�{ف��e�	���M�Nv�'QV*#���Wv�C̅�jH[Z����݃�o�J99����i.����F��`�ٜ��xSb̓V�y15�&�V�+:��<�N\$Rq�xb���f�?��|ߚ�E�	�����vՍ���8Oj$�vT�O4�n)N���,��P9G%Kp��s���f���1��3���Yb[�]o����p��09�-���1j(Ԃ;'~_*�G�YlE��+��q�nEC������d_|d�{/�������t�Cc\��Nx�������x��$�t�ؘ#�+!�r[�쮤��U����� (<j��o�п�f&���j�B����7�P|1eO�3�2��}��~7
��y�VA^t��|��g9߇�~`���%j��8Pw%�!3%]_G��cS^�W�Xگ�dg��� ���vubmO�u,U'�cа/f�N�3�|}���_'�0K�t]��Z��Y7���J!.h`-��V���J��8\� a��>��ȻAQ��T�+�O�yu@��S��sqSC�,�EPF���.I�ى���h�Ag;cd����+�D h|��&���7��cUC`�D��@���ɐܞ�o>�}��x�˷���>j�<BR�C�x�<	�����[S�,\ >a.�B�����<?�<k/?ޣ��pB�-��|�^C�t�Bb!ۙ�ͭ��=�E�k���D_��a-=;[������Q>f�Z�)/���t6�����DB�˓:˻W��D�4N?TJx�>� 5��Z'ۺ���ˏ�n�<��b+?\��jV��O�֮^�N�A&;-�0���6k�0�$K�C/�GM��H��z2��'��)B჎�,Q}��z�Jȧ�������N�'����D�$�K�e	������W��c�w�B9�ۻ5���TUN�Gq}¹z�������%]n)������e§�u�+J-o�s��!jii�l��Z�Uv���s�bQ?6����YY�0�mu�\$��l�Y>=���/�Z/�.���&��N�3�Ğ	Յe	�<�WQC�𽥗i�ZQ O�H��O�Oc���En^ c��&��a�䲑�[:���[�?�%fu@��q|�C�42���?�� ��B�c� ���oZ�<hJ�vHҜ6X�A��M5޶�ߜM��S��\�sqc�u�Y�C����M+F���9�����j�,O�y ,&�x��ww�wwEx
�:��4����m���Y'}���}H�8/�����z�A�~�O�\���0���/����m�.TDUY�k��`��Η9}B�<	�	��@:Tf�����KA��\�^�_'��1nD�F�[-#��)����H4��6$Q��R�����Ap�k��M��pu*�����s\��>����fOշ	eUDi�r"K��p�^@���x�sʤ���k��g=�dR�:n����L�2��&G�u����e��r$��B�S,H�s��v�lg��P?��%�B����]M�l8j<*ݏ߂R��i]5��y��Z#��.��s�V� n�����R�ɍ)��D:k��!�p�b{Qd9���׶�
�io����Ȣ0�:O=*����u��;��4S�漓���^9���h��!� )��5�W!Ⱦ�������J��������rD�Q�VQޕ�~\�����Th��'�ԏ"M���i3�K��KWq�
�
�����ԧcrZ�&����9Ef�-���fṦ�SI( KL�����7a�&�6;N
yV�z4�r
&œ�S~%����+�nW�o�g�Ӱ�B���5i��S�Ⱦ��kj,��6=��r�1܇�Q)�<�ߛG6Nx+��O���n&��Q�xe�M��<�R�����N���,,���Z��p�O)�8E��,����l�߷M��|>bɶ¬������Y�7��-\<��C���;;�����jX������x* �5�?���Y�"����:.�9�{�Q�<�f�l�
V_��_+�u�j;�?J�ɉ� �?hT�j����Vr�����UF�5X=��c���=puu'��ݧ�R�j�FVN�Q�76�� ��j�g�8���?9{ø�T�M��a���� ��.`��t��HЌ�2��L+��?�3e9>����6JqW�o����w�����t9��C3��R���lZ�n*�u�YbH��J)�?���]�A�86��w-��\e�u'׼��w�~;�����K<�`.���hw
��xm6@c��'�w�xS���g��w���0��/�#�O]�Yr�F>lĸ������ڑ�VL�?�u[�J���;z��7��,�Yt{��%bWV\�g�-��K�2G�
l"�ߣ��t���_�UZ��@�~aO���	䞥{�J_[B*jTáD�x�S��'C���bb�,cq�Ŏ7���F!��m5F�|��N�;Z�7��p8�ѯ�7d��$)'d^�T�ԥq����jE�}�>�{S��ntҼ��e�gA&�wkAl�E�R�R;6A�Z15r�q
�!n0J*�F���Ԍ���=yC�14V.�0������Iє�t�����Ċp�o8_:�l蛟��Lm)����Q�	+�D0��Ïh�eY�L�%���S�.�]��)\�?�Ǟ��E���L���ǡ�=�<r����Er�h����A���>�}p@���1&�EC�<&��Q��Be���ːTB��d�`�ـ�cb@
���I۴\�ښ�7b+9QVqA�����U
$Q��vy����qe�Ϗ�o�o�B���Rfɱؚ�R�x>.?�Fʙ^�z�&c���+�_e�˙�F
�ߐ xK
����4�f1?���EJ�'z�$����)�|r[ �x�$���e�����9�mT-�Q�r-�F��-r	X��kr�1�@��:�$ �Ȼ��m	6�]�c���H�&�iF�S���6�rD�W�S��[�)�h�Q���օ�ȭ�T�� y��r��iY3�7BGI�^^�?d2����|Z�����Nܕ�(�fC�X�ۮ�$W�������;��*�x7�z�K-k��ʰ<����L@ "�"�M�� "�bj0����8��vZ���E1`h���8(w�*�G0%FC&��&��qy�tcO�Q�����X�ԕ"��2�������� rǁ�K���H��T9�|�!�p�(�>#/\�yV8��T��X��N�dkc�`����a:��oW�������Ak�k1���s(՝��4�EAϷ��a����S�x��Go`E�[?xN����e�A���9�g`qRO�c�.�)N[�!�u�`�
1i���Q�O�k�}͂�N�`3d]�b�F���iw��!�Y�_=Bm)�d4�!��{��B��:�
vP�w�fM{��f���- Ei:Ĳȫ,�~!GC݊��%u]�bTZTׁ�j��i���E�Gq<�B��ea�8��B��	��IҺ)��Yκ�ÕbMn�ᷛ��M {Ͼ�|�+/g`�9��8��	GD�N��)�Fr�Q�gh:`fk�H�3��!�&� Vs:�`�mG6���ɽI,��	�@ ��0�Ȯ�|7� Da��j40��=a-1�8oe�ClL��&��k�c7S�3�~�J�D!��q[}����@Sņ��o���P����<�&�j�ؑ�(GRQ����n.�ԯrsH| Jڢ�L����b�!���=�`�Y�aٖ��'A30N���|x��jL�V�Tr �����b`2|�3���m3���$��|�����b���>�U�1q�o��&2�H#ymN�@
칵�}�}�H�A"��6y����%Z�����'�w����	�;)��T���׮��M�5ԛ��!����?Y������~�>���H*^ڍ�3f�~b���҄�@�ڎض?jsX��u�F]U���4��c.j�v?�D��Y����sy��g�~��MC*��.k|��]~�8�*��tN�,{���H}��xÛ��{�����T��=�%��m�o��E����
��ͩQ �Jkw�P�Rd�}H�XcA���4+ȗ�}�?^��ֱc:y�6`��F���̅�"A(�6������[�T�qz܁�t\�C�x�� H���-/�����o�&��v=�w��g��Μ����PPlD-�m�;�/�U)�n�d����rݜ?�>羊�^^�՚���0�E��{���:��?�r��U�3+�y�����4�����G��qQ��[k�mkiR��(���X\��Ĭ��+^���g�yEUQ�_�/��Jll�s�MM�}f#�U�9��m7���P&�\Ft����D1�|�,��#BEu>���c�Ț߃�~��2L�0���$m�/+�p�]��:GM=l%�Xڠ��M�~*xr���05|���E'��2C(@U��\��W0(4�35+f	�8n��A�������bE ��������-��)Q>��z�2[���@N z��6�ܔ�y?곮Gm���ب��)�W�N��O��ǣ./}Á�R�އu@0���Y7�$"�8+PR��BǕ�x'�gi1K<IlnAg�<b�D�����h����u_QX$�p�����|�K�T{�)!2I}����f�fgS�"�����Y�ڂ�Bޟ2�s�pY��cL�U��Q�Xȫ��>K8F���D�8��([<����'�e]�_��~�@������ga�G�	|���{{�� �I7͟7a��\���u�K�tR�����>J��h>��|"�{,���Q�*�YQl]�)1��՞�Z!�+q��������\_��V��9���Ou@�������>��&���HP���w�m�iĮ6��BN}k>�5f^��R�^Y�C��4G-y�~ʏ�o�lK����
�N����	��,+o�'0ġyn����w����l������\�	HLi筑���@�)DN+`����7������A�	ၪ�[����̺3h�e�T��"y�~3���ҋ�r���biz�^P�7W�|E��#�.�9���]�97�{˻�_�I��6����k��	VC�������^�KD��y�8���D0���n�R�`��*��)͝�y%�|-6�y@r��xХ�@�H�Jz�w���[չ����\T�mA��Rb}#�����R[C��M2�E;S�=LxI����1L�D�e��U�A-��ז	���# ���eK���`҅>!�}���k�/���o��
��ܩ��U:B.�]�0�)8|m1FIs�<�"A ��%�zT�j�
i��D��]X(z<2ϥ���b�y��$�#~ܳZ-QD�{n�P�f1r00$��%�g����͖�lt	v�2�O��+��m��ۙ�t7�2)�)O��g���*�f1 9��k�tHJ�)��R�����g~7P�U���#�GEg�씧��B��1{(�1�T�{�jř�ݘ�ҨT���`0�SN�$�V�S�-�}� �c�"{݃�Q1l &q�;Ϳ0B�҄8n��o��5�M/:�bS�j���,��D3�1(c�M5��������K����."6Xz������r�x
6��D����+�tq�b�.A���P7͹v��`�2���Ǧ�ecu�6�ӭ|�L��G�ua���&Guә������Rc߀J��9�H�]�{���Z��'h����gf�[$v���I{�	����>� �d�\??�i��h97�r�梐ss��f����9����Ӊ���ոl���Z�S��v�����9yL����ĝ4_r��5�X��p���B��Y
�L7��WN�z�'�$� �鹕I�����F�Ϣ������$p�	=|�����D�Fa$Sd��w���}�[���8�ۋ�ㆪF:��g�	�&�S�F(�q3�� {P�!��"�Vb������"!��>vY�tK�W;�p�\H�h�fL70��>98���A�1OTղ���<�ڗ��x+��TNB�拞V�L�㥨\�F;D�4=�M���$�Ptt/7?��u����c>mK�2�J�.젃��Ks�
�m_�F}�{d�1��BY:X����N�He�'�#x��y��ӏ��&$�;g��D��J��v����z �x�P�JÉ��T��߮.'��q�����Y��u�쾦n���䈝�^�l8���؏г��`�Y�!����{�iTb�~FZMf�u���C&���;�� �NO�N2�7�[C�E�Ư�ۊ���z�oU@|����o�L�i�{�l�Q��b'jp�/� (M�a�Nm���4�/���{�I����L�o�>,G-R 	�uJ��%cűjS,p�1:�f����Fh;
`�tJ�"��t ��^ݮ
���r�C����dw7ٶ���R���KY�Z�LAKcr"��~]&�+:P�Ni�̆8���]w��ę��?g�Hݠ�)7��PW(u��>���t��m`��Y��鿡+PY�.���zŉ}�U�P?ݺS���i�8�0���	�^�G&&a�� O��('���yB}(%�T�҇Z�N�N���=���1��j(��04k��)GB&�f����PKqd��f
t��vϼi~@��.G�L/��ۨ�F��q�MX���0�t�gx��U����K䈎��"v=);�=K�9D��,�Q��ϩ{a��m�F8���Y��㓏�V.�д|�L�n�O^�Vt�����HH~�^�>�уP����2��G��a�K<��F��^��-cp�#j/)j�����$S�2[DBW7t	���]y�^�W��P�	�(.����c$����G�h1)d�����w
s}3hwS�*i�u�³�	����ت�9�͌'���=t{lU�_i#��!}{5Lp�b%e) �D�XL����Nɨe�
�X��
��ˌ��a�t)�]x����Cz$�^�d����L��_��<�kr�a<E�HH����P�QD��|��y�$U���Brq�3�՞E$X C�<��P4� �翆l~�����~a�%rx�Z�u���/��IJ�?���<��_���0J��Vm.�f�<gH�����֪�����9Y@�*�(ܓ�7�X1.����'?k��a~I�aI��]QLεk�aS@���sB�)�y5�r�wE�6��;�!�n�~W�x�$�:<�jت�F�4	��RE<�n\�9�$����kZ�?��~I�/r��-��k�����=/炾��������;�*,�}�	�U�	�4A�S
�(�
.�Y3�5d��v�Q6
���g�e���x߽���
-4RGj��孞Q�l��P'��H`ܲ�����-�`Tkxk1W<K������X >�*�]J/F�]�yS��hh�}4��_�2��z؇N�� G6�%뀀\8E�GJ,/�6"����'�|�EoC�Nw�?W�흜�O��"ZF-��v=��o�=�'��4�)�b���x����GڔBN+sO�\4�������ݭ$��֚����E`��$�P�:�����a��t�T6p�l�I�t�}hW~_�߫�֞����߈gs�.z>hb}�+�k���AD��s/�>�"JC'%�%��'�Y�-@4]C�&
���}���|Xߜ�8@1:��>ʒ���:�I���fMR@����@2{�'R�j�Gxo��/�����|��7��[X�_�}����[�,�fq�.�h����U#�G5֛�"���+��V�1ךVX�/p��6f�ڨ�l[5��Mg�[z��1I�A����c��j�ë��\�kwz�6�l�m��JI3t95ƪ��k
�N��)uD4����{�V���e0P�\��/ڷLI�^m�f�U
4=̜[�Cw�9d	$b��ow���6L
~�p����M���U>�tVk���� ���8�X�ޗ꫉}��I���"+_��{ࡨa1Xj>��M${x$����u?[����t6Y�-�&��)��3Uc���c�� �Uo|��g<�]*�Ӵ�ٌK!'����S4�Xӯ%w��i��@�����W�'�5�KQ[
j��:F�z��&�PF��H�WRʊ�]M"AQ���[�K�A�Ȭ� R�s�[6���\�mQ��i&�,�o�k%�=�s�H�x�绠�Q
<X��B0���BbUpGT�+t~+�1+�:3�^����*0eV��^�UW��ml�MoNގ�_M�*�&�!9�M���yo{%TL�H���`�O��Y%W���1�T�������N�{�"Շ����l�݁z�s%g7MߛGO�ѽv6�̈́��=�(Gc���a-�R�$_��?S�G$��I$���0}���\�SX����3��m����8)�damt��f�i"(әn�#���ty�(ŋ_��1�ӊh�qb�_���4ʌ��Kג\ec^ʵғ�����z��]�+ZX{t�t'ٺ�9�|��� �����xG������\��f�!�l�v��z}_}��}�+�MMH�ѰW�-<;0}�՝&��Qݚ����x5�3҈D ���(~�*	�S�^
hl�et�l�Nle�VJ����h�y�Sǡ�`^ҽ��7V6䙑�,�V��#(z�On�	d�r2pw�D�+L^
�0BQ���x1��M����J�J���
��Hc��b\ofB-����+�nb�<���%x�ң�*�p�QL�}`��U��f,�6?�`ٻڋ�r��q���Y.��^�T�:!"��]3i�H�����nsC����[-yջ5ɕ.��`���)��� ��?�G��/�@��d��S�`Q�߱��r�i�\J6JSǒ �,�[�?#>�\L�at��=����<�>|�#��^�����*��3+�۳1����ir�7�;��?HRu��KD"�����A� CB�~(�g�욒�� -�#�@��`_��a��>��H��p%����y���#v��w[��m�G�S8_�Pٰ{�}�# ��~�D�8�����o:�	��@�8z�t�H3�O\�S\�J��Y�*�FS?�QN�!��|c=�,z�TemoR��.2��>���#��Lm-�e[jd%�GW����]5�%0�����	[n��};rg�R�.#g��mq�@�d���0&
X&�:�zWz�C�?�ޤ�^�����$�7O�3r����$��^&�2�]�}J���y����|�,x{����pz7����Q3��Js����zatGNw��T� ����d���*U��l<_Ä�����o��i@�Z�/r׭W���直0W�N��U���XV����n{�4u�O��pa���R7�v�Կ'5������۬�y��}��W�
�t2=�ICE�0��-���;#!|z͵����8w�_ew ���ި2|>��j�)r1-��E ��>!���_�5�<�hXX�l��O��F|�c�>�����=d�F|JuOh���į�*��<G"��gk����`���j��9C���)&��&3�ݾ��S�
���¥���i ��S>%���◌�)�7�;Sjs�J�=kr�@x��y���V��L�=�ů�Y�A_�o��Ā�O�Lk�ܑ˯���f!>�St]�<N~�T��v-Y2���[���"!��9���_U���a���4Q*��gƅu����.mIM�����tC"���-�[	^cʽ ;�nL���ˁ��Lg�E�:s^���P��a���)^�b��贓���"BQ�T�[5��tHlۍ��2\�Ԏ	RZ����Eq�������+���Y��;�}4��b�q�@G�<��0���D]�|��&���R��³�Q+6
Àռ��N�zJzMP�����vn
��c��!ٳqO��ª=<�l���r8�Fzf�V4h )H���q�B5?Z�	xNc��ԧG.���S��T*'*l�k�q��h���;�C��y D#x�4�A��N�St2J�`X�-_�^�<�8x��_ĩD�Cs��
z���| �RP� �H�:�9n����z�&����n>�=�j�)�D�<�g�E�F�
�e����Iy�}��*}�/7hW�r�G�t��Ӑ){�!0�@����ƯR܊�U�q;_�1/H`.ʝ[�ܲz����^����W&���^�a�	�`4BD���ɶ�a�(�˝�l�w+��\�%�h|	���/en�<��g��I�*j�<S#���"�w��N���}���~
���5��C��ܿ�Ta=�dif&0#x�g�x�mR�Q�6^@���8"��>WPEl�@
�d�
	�$����6�K0ѿ� ���';��㺸�o���IDs� '�:M� B[�c1�ގ�F����J����ej��ѿ{�#9��'l�}�9,�H��?%ebXtו��J6���8�e��ЎX:�\��}����(U����	uTA2�Jq��r��*z��pVo�$8��%�G�m�U�E�� ��k��X�f�$�[��t����/<&\�h[-n����H/� �Q�kF�'o=L�!��*�(�Ad��1h0�:����c��rA`��o�c��ҹP�Z�fS_�#� )��o��Q��֤���������ߥ{��s]�Xɩ�gG"�N-+ݣߒ�H<�]KH�X��T����u��}tH�j5ᵬQ2P�c(��jE�`ÀNo�^���SM�����h��ѫVX#��ī�A���ch���e��?��2�Q���cǺ�k�jU���+�u�vm1�ȓ���nR՟\���8�$��'jB�0;�ՎWYgpREW�`u�Y`��l5*Z�0ʗȦ�Ĉ�q������bΤܐ-���)C{�q���yG���}�NsA�WE2Gf6|�sA�&x߃����.��Y�hQ˦X��!*��t���t%)F��s�#�)!d`�ٻB�<���e"��YܝW��J`[u�������OAt�Y�V�W@��(�uI�����l�t���\�N������nu�H���h�6]�.���[uG��*n����(ÔC�o�?B�4�v8,�([�bHE���z�:���=r��y�s	�,��)6F�$�s=�T��5~����މ�B<��;�J A*�S��v�����`�������wp�(�辆��<�!ר#2�Q{[���b����IS#<<^Q`� ��ԦH�GDs��|�����X�"�?h�0����[$)&���L��P!��k�]*�񞲢V�/���u<7&�۫���"��t�ubE���ޢT���W��QBad�~?��4��U�Uep��}G��K/��h��>0 �O�j���EE�6Nͺ�����Ӄ����wđ ���xM=�-�+}����2�N�����¹1����|;2v����b3�S���0H�ȵ!�Z��iN'���:}��1�;f_W��X��$t8��g-}
��O6�p�=���s�N�=&��N3VğN1qnJ��B��A�N�X��⌠["ջ.��z��%@�6)|��)�H*�c���O���U�';���i�"�$x ��v)����j�J������C����� ��������6�Afm	�	��qڛs�v�����0.n�.�U�-�2�?c�jE� vfz-�T�8�I�'�~k$��BC���rQ�?"CFM�`��<�3꒓�|�7ueB:��_O*v�l��s�!BF��b�:�ƒ]����Z����~5��2E������?"�iBdM86���EG.0p�_�^�L5|�w���cI�?Go ���6m_Fs������ĸa�{���Ѿ��g��}`���'�b0:EkО.]���Y��Zp���=fZf&�*�@��Ϙ>�Y�魙���7�\7k�b);���-6!�E�uzXDa��w���P�6��@�H=LBc���!c���<�=Ё�5N��~"T���B��z��;���j��M�؊��4�&:=.�5�'E~���N����M��6�F���~P:�P8Lzy�4).[�E`�!H:�����YH��Y�>��ع�4A{3:ty�P���*s��=P�i�^_MM�Ƅ�c}4�h����i7���\�*��赎�h[4��#J�޿��bC���7�=���
`u�#y��u�NH]�d(
8��œ���2J������1+���H��-��G��z��ϡ�x��>�W�.+36P�{$�'"����hNjK͏#0����ʑ3�Q{櫑��W�E��IPh��D(�1<�c8�kדu��O:�YI�.�0�4x��0$�4 @/O��)��>W*�K\G/~>i�����$��X?}����2~�>� �d>;��c��J���sð�ü>-˂~r���5]�zL=$�H֗����-q�0��B�A���J��K"�}��x�j<�.6���q�b�?^��_>(�΂�A�jK��+Z���
��ux�i
8�.�}F�g��+�0g����+j�1��H����������`&��ɏ���
 3g��V�	�tx_d��eԦ������FFΓ�
Sr�V��}�E���[��ZX/2���
j��5���C�=�iH��y����4��hX ��#���ʞ|P����2�Vy�<�*�1�T,�G��b�qN�C���+�+Aжc� �i%'�C�_�]��K�v�@nPSɛ����6{>�c�;3�5?�����n��=��7�oPk�G;b�?Z9�köF��O����G
)wUw�S�\O�uR>\ՖB�1/�6/1����dg��m��] 0�� ��l�� �W�5�+K`U�r��ӟr�Q��š���M�h&	�*����yצ�`At�aEp=c���q�J���"?<E����k
_�Xl�����+Q��u��Щ�t��|���`X����^8Oτ���s=�X�����i��|^������2s��_�8��}g����&vK��Y�jW>P`�߲�%�б����0j_��i���<���'M�\�(O-�Ρ���S���2�mTV��w��4T��_!�(zo�o �_��3��V�]/���6��YS@{�	M���ZZ��U���~V����k����;� {�g�������26,C>�\���H:
��۬�f;@.�H����]tl����^8�쟾s~T�2'c��Ϥ�>י\e���� �CkX�M�wŮ�Q+��q�y�$�iZ�W8�",	t0���^栩��s�^5ʺgZg��b�j)�%Ϝ�"�iŴ|4O�['�nCe��G#�/a�1��9\{� ��� [�p8n�'�'����|5M�In_�F�v�/�\/[HƮ�Tp�F����&k�b7<�;V(���/��{�������S?T�2
'萊!6��<Bv�ԭ�L&e6N}jI�����nD��ںx�e����������ֻc��#��BB��<&xڤ�}���qk� E�N�2��U�]V��hso��G�2[9�Vqz��)W��$�+�WZ������]�fhc�]��t�~��w��NBn�h�W慥���d��c�,&�ꂘ&�Q�&��D(��Ξ�N*L�,�HB�+�)��SWM���4)��kIm(w��V�������E7�U�:Od�uƸ��䐈� 0�瀍�$�	�	>��z{���zЌs4^A{x���K\�Hx �� ,�M�B ~�VdN�7��������Xh�>���g�<GM��`�O�ԧ�n|4>L��[@��|�&.�'�^]�C��/6�O;W [#�fK`B]��S�k�1u^�d�\�O� ���
����EL��o�/nM	@��)#�������l?�����y/��)>�� �ڌT����÷�8g��W|;Gg�P��FMwi�k]�Q�C)�exVw��,`���P!{�����#i���d��>�e�wYw��~8�YǗ�I 4����6 U�WZ��'�,�k�������/ˠ'�go ��>L�ޥ�Aq�ڴ���I�峄�b�& ։�P����&jق��UW>*�c�y����F�A� �;��Fy���7��ۿNG�8M3�y�\dZt]��Hg��5T�IrH P	gg_�ыޚ_�yܪ�W��K�.f*�R���l<cT��o��u[��`z\l7�F��lۿ��p�Ǐ�d~?#��>`�vO�8�t+:S�E�=��W��Azkb}�C�`|!?���9���#�3����o%HD�H[��Z�;l۩����?5h!Jf�۰�]
�4��=$z~|hS���G��zf?�~������8jn��m��ߺlk�J向WFK�/��)]@fѹ/R2��Ѳ�i���<4u�VLx5@t��E�ʢ�������s�G��)}�6�6Cfu��!b6E�e���:@���tf�u"����%�u�j�K�-���I���Q3gx1��^A[�.;d���d.���G�>P,��h�'���%ԽRnWi�?z$�o����!|���S���uN���g��_�47����}�U�假Uzcrϛ��R��ĸ_�s��`�g���Ґ�/��t$+Zk��c�/�-�F�i_X��7Dd�E��#O�5�Q��8Dщ6PK�s�x���̔�[���HԚ��*�}qE�u|���{�?V�,�=,�ih�*������i�s�z�#m��� ��[�f�`P�W�<�	���DY����L_�-K,iP���/�E��S���6UD��'�.���~#����9���)n���t�~~%z4�|�P���=Q�kj����V��Q��
'�b��@��j�q��ӻ2&LB^At��w�&��v�N�Q���J�J�3@ҷf�(B���b=�=1")B��_��=YG���Nm�r�r�6�?����K��tw�8��%�8Ӧ�X���c��w�w��J���U���iYLOe���-������2�eԁ����&�l���d!���6�t��4���aQ��e~�?��6S��"�~*�P)G�������W;z0.��w��"Ț~KVp^�Z��ڲ�~��3@�^�z�8c����T%�t��?|G>t4�}:�_��{q�zM,��lڮ
(��y�Qai�\�����&����Y�	�n�W9eB��35�������1��2&���z�u��[@X!d7����}� ���A���S1�EF��ʰ��9�G5"�_�=?���jf4�\m>�𑕺��-�$"�"��
EFW��)i�"��$�k�H���t�[��zD�I�|c���[�A8�ݵ�C�J���-j�9�9�B�x�_o�,} �U��b,�	��/G�w�nd����2õ��}���F�Ϭ�oƶ��<����Y���HCkm�O>���Q��dM�A�"󅣻�9C���ҋT%,8O�\)�d#�
M��D��!� �a�&-����NL�����ꈥz؉=�CP�����?�A�8o_m����j������j�,��<��C��or ��;uG���S�7ʁ�v�ˬ%�,�-֢C��Ȃxb����=�ܴ=2��!�Rρ��#g^d���#%@')�"�DP��c��S���.��Z;����;1*m@4-��a*�J\b�fAí�s5*�m�9����fqS��%Э�4�5�Z$�Fb�+RLj>�U�}8TQ�ON��\�65]n.�HD~�X��r�������GL	bl�'�ؠ\����
]��'�L�bUC�Qp��=���%Y�
x:��'����~�[�A�X��Y��7s��Eq{�ɓ}�gw��w��陇FM\�x�TF>�[蔢W��O#��p:mԂ�gMY(5�~KS'UȒ��vQ��߽�x�6s!Ά8���5��&%|�g���̖W�����PB*���R&<҅G���b�������Z�WDaS�\,gB�����`���ap�l'�Bz����ak;;'�T���G� �f���Z�y�˓M�%����-C��D6	[���{��XH�O0xK�eZ3�-�*�ʍ�=�/�'�>�D�Z������y���S]ꑾ�d!�~9�u�(l/Tr�R;���@x=���6���E2�'P��x�*��j��&��K�C7��[ǆ����G�2�d���3i�uc�qC���@�������"z����Z����,���M]O�ȅ��պE�~9�#���mf���l3�[8c�f��?����ň���y�,�)���h��<�v^!p��������E�x# �c�N������v2�x��'���l�w�W��5kov���H%��j�C���n,/�"���)<w���%$�_�!p���Y'����E��.
[YI{�h\��JQô����WEh�t9|`!���x8���+/V�$�{4�}�$�����v=`�ǚ,�Ο��"N��P����?a��o6׵$���+����I?`X~�_�G,�^�
��9bB���5�'Y�?���4�����{��f�Wl�����ݗ#-��
��(�4�O��:�w�ku�� ���Q�%x蚠|/Ecb��}��E�$�#Ҽ\fc{��Ş����C�"`���۰@�,>�bB�H��Q��A�gU)���2��Y�nF����;��"g���g�����Ӗ�5B�<
�%"�r*d;��c�X�'��<@�ҥ��ބ5���\�%&�m4U�
,?=pN@N]���yoP�I�z������_E������绮�� �P��'��v0s5/����� )�[	���N>A�����e9єk[ݷnB���f��<��v0���������GD�X�y�,�y'(7��>�]�>@M�?#U��T��p@�2�Pn��.v`�����|�`[�~�j�Im}��+JR�a�h�g7���v�l���mMi�5�����V/��(�+���3�|����J-��L�)o*��z0�	<�4��P�KϿ=*5��6����9���E]F��7�p�G�`#����lL�<��S�:y	��{S� w���S6�O�}��"
��n�U�جTx9��I�K���悧��S��R�
��G�5a���.f��y����#[��R�f���\mPt��׶k�F��u�E抁�u���s�Oo��F�����۵\�b���I������4�Ŕ8���-?B8�خ�8ޫ��C�,��D�p�	3�d�]�dl�ك��#L�����N�*��5�
�sf,�<:&��o�g�s0�8͹-�i#�\�|�I���Y��aݦ�WԄ�$�0��롾%���MFt����Ng����.�3��{�^,�������g��E��F^+�4<�F�~H��R�~�D*~,����o������W���0�"H�� ��N_1}G��6.����x *B�B�Qæt|�yqrH�Eư�� t�M���.��'�]Y'����v�lZ�ʵ�'�=R�������2�`5_�����b@{�?��<��
�4�u$�ة�=��"c���7����Q�M�(<q���6��G�4ҧ:��]\]��/�qV-��f��b�%�ex�-�ʣd8<5g��ARuM�DY)� x�,d��3�׀h�a�h��e���Q�J#'��97���4�/Oܹ��$�3�n�FT�����R�GNmf���ʬ��B��$��{����nH{�9F2/�v��!�W��L���Mx���ʷ����w>1U��ࠊ���Sg/�r�U�xۖ*/��;�1�7��7���E�q�*L��vTe�&��%���h蕨�A��eQ7^Ñ�H�ň�J_,^��;�%d���ʩPA����paZ+Z�
]�H6���~�o�� �ڸC�3�M6��<z�U1�]�����u骈�������3��ã-ca����i�`,�V�8�0Y���m�V�Ȥ�M+�/1Jѷ�h�irhx�HX��6<���H�w4*����s����3s�a��5K��ѡ��6������v��r�@�5�����;c���Ֆ7�S-�B��$�48\>����<^�ɲ-�Ƽq/q��P�m���+�����n��C`�iv��&i($���6�{��D}�K��M�B��^#����̨���v���m���^VX5A�j�C���~SR��4=��x�u}�Яf��]�C�H��7ѱ�:E��j�e �xX���9����d䌬�m@<JJ��*��X8Ӑ� w�V�l�����9YI!�S�_�b/(���f������ 1k@C�.�
ƴK,?$W L��_�`F��T��qa]���kcVQ�B1��14�)+Ȉ�����k%�AXĴ�c�M�\��9Q�ݒ���"�~1!����uF3`���u��aS��K�6h�S�����e���,��m̵z{�{�Vs��T�Q!�PN�}{�C�O�3���zh�����!��U�,1�Z�<<��o��O����k,<z8^�fe�1��cX9˓\�Hm�eu�9 q��g�f��w��m8�R�މ8T^�h\�ȅ`Ĥ���#�m�,{�b�;�A�9B��&!v�ځ<�F�g��9���p4lJu9�Dm�GVIC�-�x�ʛZ�1�}e���/g�]�.���Y6��C���Ge�B�a�uWH�!Cp^�L�f5R V��-Эr��#[c������f9�USȍ+#�F���D��'�΍9bl�\w��1O���UY��@�k���f>~�π�S3M��a�4����G��#�ni��)�k��7uu�ň:��3�~�n�Ç��\����(����%��/`����ݾ|�7��&ޛBR�q[�,�</��j ���˅��p���.1�qS�~�{k&��ի�AyQ,���W�ڇ@a��`7�h-�{��SdQ��h2BA�i\���P]����*���1[�QW暁����<�N����>��4�-F��u_���I;*�e`$ڍ5����L����UJq�3 @1T��C�尢?/�X����I��)�z�=�Ɉ4P��%�{��Mg��C���G%x��T�ד��Y��t�8��@��Y;�8���I����%㯕}M�HR�P�f��'�p�b�}S�N��	%i�P��l���b�DG���&H��ǽ	��η9�>�pH���a�uj{gG��H��9�Qb��V'�z�(����G[�y���f�9@n��\��J���m���%�7]�l�V��D�w��1���"��H�y?$�x.7���h&a'�iھO�?����a����4DقO�c��z����$�����g!�A1W?$<H��0A*�Έ������[w��]�$�'��0��bzb�xOfkݻj`�E�S�?=�p�b���N��;�G�rhŝF���I�s�ՅG;(Y�T�.2�%�� �c���'W���iF�@����>"�"/M��ĆevyX���2U�vԁF���v�?|�l�a�RCA���� &�VZI"�n��a�8�&�e"L�Q���C��uG�e���FsW�?	�~���ٷ�,��Ei�{	�kK}~�L�l"�Z�{��V��ܓ}-]�v����~�ݹ���_gm�J��u!o�q�bڃ1[�"l<>t�/�V&�&7U��iR���ڍ�Sl��Ho� ,5P?al���G�8��(�602��\{���2cdnjA�c-������#��A0��E����I��������]p�³�l�U>�w�38��x�� ����2��|��j!�.���6���6�Hк��FdPH(v�B7R �ף��C��w���h�I�;ag��AE�$l����r#� ��9��_�1�i�u�ޅ\���H�5�1�N�\+�Y|�e;�M�cX{`��T�M�$1q��?1Nbg~~�f�1�G/�i��7���J�%��Dы�0�<S��y%\؁S�3əf��T�#�Ɖ����"����;�����Fo��|������K�{�T�ZwC'r���91�����!WS��)�~�6��&sE_�	I �P���!��vX�;�qhW2y̠���_�����
^Dl�����@3�A��\ĸ�L�npp;Ё�w�<+9����U9D�ל�}���$Jz�;Ǚ�0Ȼ���D2�S=_��Ob������ׅ�dIL�H�	��;S(=' ��x��ߪ.�3�q�Ƌ�-�aûO��\U�)U%.�A�9.�Z�-
�
Q^Z�˞n���݈c}X�45��L*�^�ih'd\�1v��c���iF��޻ -�;,�EwF�ǁ�{�3O:ʸ'�N�ˌ��Sz9?賆h���
���`<����O��R�w�<\D�nٶu[T|�V��`<��F�5�"����|�r��ds�O��ٓX���>֔"*�e �4�A�G��5��H���S橊+������Pת����J��BQ���;&��Vu�#G�ǳ@��sqc,�n�ReϣZ�A¾��*��9���b������6�l�h���nɯ�Rk�'�o�;�i^�-�P��="�_yΞ
}�>>���L�Ȏ���j=�̀%�<�2+��źIZu� ���&|N���
�W%���9�/yOU����8��Z�ԢI�)� �� ��O,
�q%��O��5�0X�FE����R�Mo�ބ*�0�X�k�4�t��^!�(
q��Z����B���p����E�2k�����'��/:ע[�ss<6,��g�P�2��,J{W���aU��l�7�.Yr��+|E�~q�-hc�p�����2�Ы9g�^Cg����Ӆ����Yl��U���*NL(���;O�M���>��v�@�ģ�S�ng��*j��x��|`Fy�D���Dp��IW�s��'\{-��f\��ҴR\�����:��q�Jr͒9I'��h�ER�����\4��؇��Xl��8~�h"BS/$���L�D�=<6�X�,ΐD��B7T���C��P�)g����@�~�Q`�7�p��%�">*�&�w�=���Z+o��UB�g��G��Ec��H��|Q��h�ތ�8 ��pc�eKI(��񭁀�Y ��FY���O�i�3j*�Vz_��e:�����+��s��MI��9V�_�l�*���f�x���q����ȭ� $~�]㾧M��v�f��'�C:� �Ss�֞��H�t�9ypzU������	�.Ӣ4���R��22��պ��W�M���z�$9��w�dI�,��ί��~���w�s�[��<2����r�e��,�]�����a,̐L�m�����)(Z:�-���ou�о�]�h�lU�l�F��;P!�T	����C���Cԕ���c�|DL�Y�m�]����Q!��<�XS��⋭fS�t��h��B{�&���o>���4��>y^�k=��,�b��������
hq!�j��$6ݴ>�ԨV�^�BcK����
����U�$���ڒ얳p���T�A�d5�Hg]�j�B�h��#��F�F��l'Z�n��I� 0��z�|�5yۇ�^gr#��_��W��A}��	^����!��+s�t��I�t��`ᷩ�K���uu������5+�"�\X}�fm|�=�]���p	��B^[4�E��V ��]G%�[��E�L+F9�5^X�$& R?�h�ľq��.��dZ����g�k:�&H�@����+s�U�k�^�Z4 �zj����,����r����̫�.M����Хc�ɮ	���Q��z��I���~B���˝`�@c	����14�Mc�z��y�gv��$���5����~W�)oxo`�D��E�>�ۛ��^%�P!GG�EE�Eg!nX���=祥���5����(C1D};��W,W[9�sMħ�P
��r�v!��nES{P�+-���7fq9iw<�F����Fd9�5��4�ˎ���/O�Tq��ß���>p�K�^{胺ִ�S�w��n`�>+�@בEt��Ta�{�F=g�J��t���E'�J�,?/x�[��^a�>k<�*e�@Ggm��hFgp�%��%z��Q��Z-*¢}�����)n�9��_0�Y�&���ss��܉I$���ҫ fj|4K�;(�r�k���`�q���	�6g.1cPk������"� ��UbaD �Y��M<�2�+��� <á��,^�g�|�[�<R�h%�i����/j"G"Q��'�
g�N�8������q���h�j���$��;l�rt�p$Y�ů�o�Nc]H�ۤ5S��KƐ
�0}�8'�2��;�{�����Qᯑ�>���㓒Z7�t~9�*g��Y׺��*�Q`	0��J烿��Ё�Pi�s灜z�m!��b_"���w��&?��.��v��/!В����!QT��  #��A�����N"��<���܍���Yd�����(���×��]JX�TOZ���0��Ue/�,Y�iյ�9�ZQ�`����@�i�/
�7~�`[.\!���4�03U}-zƽ&8�J{�U���7�V��
��
��Y���)ɿK��=��հ��֛��T��@��Q+��;=�"���ߢ*��浝�d�8���H:�O\�$�`���<e�ǃ�AƝSf�v~����q{<���[�;��s��ާo��S*U��%3s�~Yc[�{y+�s����9J���,�m09����K5����7��f�"[8���"��=��;�{C�<�qP'X:܋��L}��n�D��_�rL���X�&�mƕ�[��G�!�HO�eC_��v��:��3�m=?05׈+�Ǜ�h�U���ou���Fe��C�a�ob7�{i!"�����hj�7���؍{�q.J�0b�&v�k-0�Pa+�"�n�;"��l�5��z�j��^E(�{i�B2F���	�h� n�۵�e�>�j�%�AﮉK�G�?�G�r�ȅ��F\e�;`[{n;�s��B�قUF�;q��٭��c>D��{���X٥���;P�HVDǴ�M����b�$xC�#�����y���1�R��h7��
��Z�8�20r��b�oe��7Kx/K�t��.�?0]�ʬ�FWs���7n�(e��"��� 9.Rc�^��Ttv�pP�H���*;x�3v�Pn�=4W�/~�^R�d��F=����@Ih勯Q�9�����O���\�S֟4Fr�/��Q��4{Ո�m�ڙ�=@�����ֵq>�l�	��>p.-��K���~��^f���z{�uo������8�Ps�^�0��v��4�7����oVy��5��ۜ�6�j |��1*뾛�����g�lrϻE�V�aa!�����*��Ƚ��Z+��vd��1��A�D�>S���{G��)�R"g�/�������e��P'ш���M����K���P�ڻ�&��*�/٘&�=�'S�Α(,��(�J�����9��"	ǸE�'�]�ܕ�Se~��?�qpˢ������.�0�"�?݌Wu8K��T�"T��S� �����G��vI�3��
t��C)���
�178Ԁ�,z��l��J\h*��M�B���Y�C/%˅�e	܈�%6�M�m��b.� ��3���"kr�!�U�2�Og�|��+̕���<eY��=�~��&"l�G�����{a���o�V?\�s�8`G!��e�%����Ck׳��X~��J��$5�����[�j����t�e��P�l�U���(�[|š?��so�|1"�_���.<)��{�_�f�c��P�q%拓vf:���CxdY�ٽ/�u��.��VK]�f��.�2ب6�2�9�v2�HU��I �9Z��l<Y (��՚Y�6P�'�Q� =��`�!F�ˮ?�ʳw�Uz���!��F���oT3�\�|���jmf��G���,#q�W2<pk����)c����4��+�Z�<��t�u�/Q��ĳ��ԡ��8�T#���j���&��P�2mL�z᠊�	hg�x�u���eԁ*��`͠��_�,�����r�>a���?(���>~�cgT������	��*r�Y)�����EL�G����ğB��UD����Hb"��zT�'Jb%��)_���E����I� �C2��2�zC��54�c��͙�e�PW�C�:7���9�f{�3�8Q���Ǫg��/B���?֭|34YQ���_���ļ��'��RL����j�K��&~�.��T�I7�Ow[�
�'DYٽ�Y�Eb���O!��ζ~Wd:f\\���/�F]���y��-����a6�x��x�zC���Q���6!@�gi�u��O�{����P���n�ڍ�qJ�8��vC�ȴ�����%l������%MQn��({2�Q+�*y-�uI+eI1?=��誛���0�^M5S�.B*�|Yt�S _%$���9~O�nq+Ws}�Vs�Si���I��}i	"���BI��Z��ks!��` ��c�	���/�
��v������~R=I��;j����|հ�k�ܡ�E�Q��Pv�)v��� ͬ5��o�&M�z��Ε�MW��m�*�F�ħ.+���"Ӏ�(���;˄;���@vLw>��"l]��r*2��d�(s�ڧ4�#f�i�%��f�Z��n�.�n	�)!EU]���3�pS�L��U#�>��S۷��n����2�O�A�o�/����
������R6�a�$�n�R�c��؂h�Q�M#��:D��xc!�ȟ���w�F]�d;ltD�q.���ïBպ�N����k�WMi��*�Y-�p�=&��O�!����]��Z.-���{�������,ɷ�s.�����C���{\�D[���O<�H/����6p��9�+8$�o����$��چ)��K��� ��i�}���:�c�~GÐ_U�=@8�a�r��ﺡ��A�E����<|�?C�Ьg����*�&h5���kA��¦4���?��3���_����r���MDeҐ�Q�e����~$��s:[
��>�����e<��=���AxCl^�C��EJ5^�é/w
Od�}t���ɹO]
�n[|�͡��&��aBB��ܰ���	�:�4���c�(��>���5L@:tB~,��pSB����ݔ�E)���9w��s�MU3�a�RCH=Y�p)����g)LOG�]���+�H�z���(Ĥ~_Q�����I��V�DM�r����j�w���^� <���3�5�ߏ��ɷ�C)o;Z�s����PAAck��9$d�B�*qd%c�94EWժ\n=P���v�E,�n5CE��2�����¸�V�@��\�#�$F-�����C�t�'zE�lS.��O�I�O�1O��|o�5�p����U�/bqW�\^
�;�9�P�a3�x�/V�g���PE�j��KC�I�*�J�6FU���0��i6�8	0)�7�����R��V^.|`�0�( �	btz�&�N� Z�����CT��Я�K�k�&N�&p��e�M`E�'f�2�qC2��n��i�DP����M+ ����{�D�ܶF��$}�R��(Z���A�����_LE��۹.�:s�<~�v��Y�Ɇ�;��W-�Cà���?_��2\��Q_�}���k��"�sd���ƅH�B�煊�%ߦ�����bg�c_A�g�~�!
�͞�VI�W؝����Bx�X�L�{=�%a��T�?�����6U��᪇(��|�UM��O�a��H�4Կ����@�A���T���Z�&#�2�� �Θ��{��b6�AY|�s�WKZﻑ��C�0�;�5��h�gk\Ji��@3q�Ln���
}�4�*�n[ �Iaw�z�!I��n,���T�$M���(��L��{�l'虩ҏ���������b���3�[P�16�"��Ü�;�7#�rim<e��`�����b���)���Iy)X�o:�{l�"��z��⑜��>��]-�K���j�9�4�����Sa��͛sr��* t��keC"���W��J(��,��i�����Z�x��	�����������|v��:K���V{�F���:O���j��]DY�@�jjډ��g}�T�[i�ht�&ԣ��k?���T�����vB��s��rL�X���w�RAjܞwo�LK����7��z�G��@XoDAQ����yOķ����0�������Y pV�u����O�`��c��֞���f�"��d�Y���ž�]k�J�
�5_B�j!l�ji�8fm�I����ӡ�M��z߰3ٽ���q]�`��4���aZK���8E/� �2��6�/�D�c��|�b��-rbqu�yu���"����d���pu/�d���C��<Q�u�q1�3�Ų����z~���7��3�-x��ʢdRb�S1\������P�b�9P��J�r5��3�
�]�N�%|]	4�Wk����l���?h��\G_�ه��"̲m�Á�6u�����E�f�A���H��2/��T�����ř�U L&�UY�CL��0cl�V�1PQ�2O�!��@��EB��2̸�U>%� S����l����s*��k�H�醵a�v��?���􄻅($���`G4VS�9�X��z�!���B/s.�F�kʆ�{S"�eMHW=�������:��VI���W�{�@I���i��ch̨���H�*c�������'� �r�-s���^���P���J���W9����2N6�Q'� �"�:#$[��l��v)�lkB'4�:Q)`H��법6�z$���}YtxsU�6�xIE���r�K���o�4�d:����5~��~�1��gF�{�Z��\�������2x^���n�K�h�Q;�c;�º��tv7��ud�9W��+��8����=U�le�f <�T8���Hu��kD�
V��2|	��S�Í�ѫb\bL]�ӠNf\B�X�YȽ�}�����U�MƢ2}q�� ��K�+��뱂�8x"�͎�~�)�p�������4{
��~�_��_�U�����͵��+r�q����(ì*��l��S����蟶�Q!�dn����_Q�:�Ⱦ{�T���ͯ9�hDI+r��s�
�r���-���rR�p<D�3����K�Y74h�њ�ڜĲ��VjvQ�Q�9)���?�V�O*���Yi����K�<�ʿ㰈k$��hm��p(|���1=�nF;���U�Ri j��4��T���0;o��s�q�� q�p��z[��_%�M1E8 ��j��������L�K���JZ���E�r�EA����A6ň'~������+�K�0���[�Ci�պ^�'��'�,��[7~)�V�s\����
&��������h�L�=;�S��T��b�hl��8�z���_��߷���	�1�����>i0�+���du>�؆VI-C�O���+!t��4d#p�[���3�V��8��k���Cb�����;�~��䀘*�������<]���=d�Ye�l�C*0�׽�����q_sq�i�
Ə��iy>�0N."ԥ��qY�q<��%Mfr��x���\Kz��ϵ9t�rջ�3�!��s��_�G�J��^��ٷ�]B^/F���̥�]��^�E�xhk_�����?�yoYD
��0�=B���7o� � E=�rS�4'?�	���:L5�	��3L0у�o2+���feg]gB)����R��9r^P�<���Ll���C�ۇb�SA��U��c�na��\�M���=��KǶ;�X/��]�s�r�،+?��_�|��
�.ID�N�e��2���Y}�`�2��&[�����nq�KJA\a�=6Z!�X?Q�9A�ߑ�"�-�$sF{�m���/� �$+֍������T�j��'Q��2G�f��htؽ��� BL<(�m���}?
7k1�%\4��eѝd"9�+`�:QF��6�ro�ތ��$��/im1Q1��/�a� <b-���3]�H�b�-�����lj��L^ nZ0�i�)���$�N��\"�gJJT6H�� ��{#U�YΚ��<�7:6WTWp��Y$�"x�M6n�d8 �=�<:�6Ua�נZ���iԻ�$k�^�XL��'%~񺭽USv;�c~m��Y�K%[h�[-[|i;pD�H�H��K�BV#_��\4��&�uor0�/�d�{���R�C�>�G�Ӹ����{nK��y-~��i+��ԨnW��ˍ�?�:�,���Ea{��rC�­�n�Lo>CI�W�KuJ헳΢���J}�ٳ�����8�~{=R�TȽ���&�>
�������q�e��Į}�ER��"TZM@���+;9FI���=(k��1X�����}�|�Dz\f���5y��_������Eൢ���@֍v�#�v�;fp��O�����|L=�.%S�(��&������2�P,3����}�̗˴}�n���O-O\���(ZNYdC9(geu���X��H��1��A��(�� �e�%m�A�Aa���H��a���2�Uɽ���uj}�XKq]*[T5���e���	��|�zqUAL�����C�ƔG���Wآ���x�VH�IѢ<=�N	$�3g܆�Q5g�L�jN�B�FG�ˀ���c�V,Cj����S��'[7�~\�q�n���H�^[��掯g���\ʍ�:��1���6��kt\�z�e��k_�2���<��z�g~9��A%\:�4����d��xn_Ё9����7X����$�j�F��ZNfGH�r����'�W���'Ͻ��˝�}���^V�����`b� a�ޛ:�ɝz�̴.�?��MYE?�ϭa�$_z�ϩ�ι[�=Hs�)�f��|�%�oG��Ic����(J�����1�G�fpJ�*�e��� *��rI�y�atS��w��Y�^�x��K�%-���_�n�5����bI�26T�f����W��"��7���b�fLA�	�:f��_�fvf�Ԓ��1RA��G�\���/�����d�:����F���Fȃ�cA�ߦlʍg�N˰{��Z�n;�R�˚I�h��ӛ�hﱓ�G�G��^�.�|â�� )4�DQ<!:�(��B\�o'����b�����-�_��LrG����l��س��8�H�;�<x|Z���60	��]J�O��.�Φ" �FqI*�uM-���Ly�xw)��>:h�@�3����%p�R�gr����>hI'v@Ӿ[��G�7���8
 ���Mӄ-0S�Q�<��WE���G�te���A@|���ό@H������L�L����w���a��d���'�^n�#C瘱ni�E�앖=���
��пʈ�����세.`)M�R��=8uϤ�.9����v�18��#�`ڐ�_�w��l�����*����-U�˃/Y�ǉ����/��Y�jE*m59fE@ >5i�(���:��#���^����L��.*Ҍ�)v>��������z�'������Д�`�����ͤoO�$�C��oH^O�!א\q�$���̿d��茮1���B�+f�ݨ}�慚f���-5u�c3q�h�����	��0d���B	صΎ�[�9��^�1m�vl�P��Hnࡤ�^�Qr���*�-���7��
ѱ�}ˇQ���ip�Q�O�����%�O�T;m��z�"Ǥ����4�}���@e�UG���ar�^7��o��Gs�]���Cٓv̄�^�]	�������(�K�c��,���(���E º:�k">^t��fW���,	q�����]H�;:�1p�������f���l��EQ� d�b��0�]&��}�A�Hg#9z���2RIKCBG�+*ڥnKH,\ ��{�o�Ɠ� �z�h����sA?�2�8��ʱټ���^17%��������%ta���:�G&E���>�1Zv8s���ok��m욊�,.������b}�JQ� �OM�M����DgtwJ�&3�ŃfZ��j%Gq:��s!���T�V�12Uz.��{{e������E�\r��ǒ�@'捵(��f?��_���k���� �e#��;��	�haַO��-�8���>	}�$'�(_G۳��W��Bݐ���6�@ʖ�-�?�M���q&��C��&'6��3C'���^�Y�k�K�����,�Hj��"�<�3�T�����g���3:mo���jUI��3�l���*�Y�
�A�
=�F	���g�?rlX�,�X|�ڰ���x��8�@fl���b�*����N	P��ES�y�"��+rqDx�q�I��B�v}���i�N�-}�p#E�U�E�{���Jտ#�q��TRS�d�h�E�{TC2�& �JH���D)�UH�
�WZWgj->�;v �����ƻ�[���L�JP�
y�i�@u�xal"��V^�쁡é���L�.X��>���_��휯Dk	�8=��.����TRh�""�o�GC���&����1;��G���QR�=�L��;� ޥ.��Z0F��|�?�p ~�ERR�Lh%˵΋�#(`d��G1odKζ  
-�H_B|iX�crv��qEtl�*�t j���@��%���7'�G����J[iW<S�~��K��d��2Y��h^�ta��ŝ{�	�C_	��*嘔\I�y���~�/b[����1cX�Ų�"T��J�-%�
y�+T̰&�ni��8���Et�lܵvQW��ϕ�0Q��)�6~;���J�z�_߮y�9
^�Z2��"lOF�Tq�����,μ���t.w2Fjw�^�Nl���^�>�g%zo(�ç0�6L��Vr�MQ���#�ߗ��yH��>d�+�,��c�5[����^�|��r���hd�d����[!��9�����؁���[񋥒�u��x�K��.+$$���Vm���/Ŀ�&P��x��@Tv7�2̭������?hK�Y�X�D�8��uAO9��z��ڄ�vIt����a�N����V%�F'd��1��э�6������y�r�#��[@'J)U��i�>�2�>b�"�~c�1]��3�!���K#�^v_��M��W�e�Q���=V���ܽ�n���4@m�fG�jB�$��B�c�S���0��nP�\����X�!sI<��%q�a)(]� y��{�،�~��j�,bk9��U�6̰w&��K�R����'�,!EW�_�&�+�W���G��Y� ֵ��圅�F��-Ҫ.�`��"S_��S�[�����y��i@���6��$f�tO����k��/��'Y�*_p�H�	�.��P�:��	KJ����i��G�%WbG��3v�D	� ��P�[��������$�3z1�P�G�@��j�L7|��d�|>�hO�&��j��._K��!������V%em��Y�YFx����K �W���s��,��^�1��v���
?0h-V@���9-���-ܦ��3z��%e#�~����~� qHc ����fU�>�Z��[l�M�8
ld�x	��8�6{�s	���a �󧛒�t������R��q�S\Z�Y8�#7�#��� 3 3dMT���R�K�媵LA?\�iϡ=Cѿ�;>E~���7��`v߽TĠM��H�d"~;��,6�{5�Ȑ��P�t�p�8`=r �i�	��F*;�I���]d_֖���4jAV=!{�ԯϜ��@���i�-j�U=��~���n����UMs���	Ok���шJ���޹�-z[M��������H2P�Fy�p]O��������5�9���;�T&Z�{Ќya���~�jۯL�i-HB���}0��\�G��C����
����;�!:K`i��'��pol��S�i��d�o8�ee7��?!z�%��)�6�(��<1� 44 @j��6騻�B�'*��]��m���6�Q�����g9u�����i��ΞqQ��$A�g���=bɰ~�w|���ݏ�	=BĐ[������x���P]N	�+��!!��o륾����nW��@Ә-%��@l�Ӷ^(~�?[��`*�	Y��b�����?�ʈ����F�W�K�A��QE�z��~2��֕V�`�$d�[� -D+i�2"�,G�����2L�"E��Ps60Y*����E��T%J/�L���M�6�v�L��cW|��ɑM����PNu9����H�JW���0,rp��Z������B�� �K3�p`~1�����O�Ɗ8�Ѓ�D�)C�#F�6�W���T.�z���vu��\�>KKb�C4�$�����~��܎B5a#;D�7�D���&��%�" ]��Z���%�x������%��7�U����<6�_Ehӣ��kD�wVFmC���*��Kh����C؞N1���\�8�o�-q1V&���<p�3l>����E���ݏ����7��S���E�q����6u"�!�X����ѣ�@2���JFΤ�^�$�_���)"�0+��$��	?n^��yI����v�@�+�bZ�� Q���T+�,E��h����A����5��ʻ;t�?��z���,̳�[�r�z6Co�@�2H�B�\�@�3y~�p�oߚ!<�୞o�ԭm�yή�է[8�qd����l��Y����CС*���^�Nf��$5<����8�<	��Q�*8)Ѐ���kI&�.�K=���2�s9�`���Ӳ����g�|*�a���wK�rO�9��W�����b5���a�(8�Vp Ԓs-�nb�g�SF?Ro.#
����]�|�w�eo>�LhW���:�73�F"U�[l^��wy��ރ���j�����/Y�T��(���C����Q7&~�M��摮���)^mHz�O�DL��I.�s.��@ʹN�s����7�6)W/A ���e� ��*$��M-��j;_�%QH�%�c�g�O���@�Ԧ����<�%�GJ�0��=��6'S5U�e.j::Ơ�]=���%��ý��Wͥʡ 0�Pd�^�&�h�(�}�'�$�����Z$ʭ>���|8���u����L���w�v�І:�&"4c �SC���A�k��m���Pa���+rXo{hN��Pq��QƸ-wz)_x���U����N�3�)�xh0MOXɛ�p43C��v6��E�vKA�JuSR�Eƪ>->%��j�" vH�p����%]%�Rbg�6q CFC$	i���j����!��qT���h�3�6�Jb����u�O�S�qIS�/k/xa��:ѷ�����Gy*ޝ�ο^�(�%���G&;�'�3����`W�ܟ�`�K�@�bI��(�q�.'|�9��t����`>1(��.�\���X.�G[�'2�i!x,R���#��/z�xͩ|�hzusN;�M<Jh���Q]�I�%h4�N���H/5^�8w�U�Į�Ȳ:f���@ a������^y$ ���Ce�y#�Gw�B����B��{��>?'QBA�D�m��{��@�DV����T��Ȅ�:��)\�Wɬ�I\[Ő�:�T����
�����c$��k�/Yw�mҒh��V� �w�4݂�^��L�e���Z�i��NүT��]�1#a�G�������rz���C���5�#�yjC��gS�	V��p��=|�v�δ��V�Q
�D��P�Ib�(�/�#�����f.Q���v�L��d��-5�c�d�+R�x����t"%��"c�WQ 
�h���n�y�.]��qָx����M���o�E��CqΆP�����
M]��s��o4�$Z<{�8OG�G+�&`�^�N�)��aR7�%�����TVOB)�m^�jD�zC;�#��%FӺ��Hr�.e��d9�\���pX�T�AŰi�)N+�е?�D*�j��0C?��I<_n��+@Z����~R̏(*����Mk�ӏ��_����2d��f��~�Õ�X���a�K��~2�Jt�w�K~ÍD�5h�����G؊<����EzF�W}�b+_�ʼ{�4x�U��l0��L���d�x��
��
��H�Z_1���5����+R��=>�E+���(:y���|�J�U��֋Ԡ���J��O�Y�Ü)���:�*"�b�'.sNl�J�
'I?��mC�&	��2�8(��z��܍?"�B@�L%�I��.W�xsǌ���0�p(=hRa �R�9lt�]�:IzHL�M}Q���x����SH�?�,JK�?W?�Ǆo#;-X��=�=��ES9�XH�`�3t1�������HArƿ�/+�}���5�a/�>q�@�Ad�&�3��R��1jTԽ�Ū���Q���d(�_��G���)�1��������@Ks�����ҬiT���K�[���`L��.��C�ߪ�z M�ݟQ�N���6�`0+^E���p�Up��#/5lf��"`���(>pb{oEV	øz�
{b�e��i�fX�0 j;�daFg)V)2�%�~wh���a��:ׂ4��pVk%9��7�������2l��.�7C*��7]8	��|���� DM�B.�� �&����>};M/�~����*��5�s�A�G��s���׻�>���J<�Wf3��FZ�j	�s6TD����ؽ�Y���ɩ�k5����]�Q9��Q��m'�i�ɦŝ�DkO�b�g55ZF|��K�s�t2�%�(vK��zf�brŊ���e���OŦ\��d4���KDc�-�[.����ٌ9{��5���5��j�bx��)�s��ܜ񤛈�Fڬ�ih~꿔�=x$O��2T�S2KpΌޔ���u`�u�﨟}uGx�p���WOp���u�`�����LP��k
l��Jafڬ�ĽV��W�l��V��s�A�?�-�Ҕ �]�M����9��j38A��F�����A����wI�~Wn�A]6o�o����ՠ�Ĥ) �}�r�=@��N�4��p�A�Ш-zgn�ĻT��b�>�Q$q���
	h\�v�`���:g���|�AV
�%�1-q�=�Z�Gc%�@�DC��"h�bN��ʟ��u�m��}��D��Aj��M�qn^5�탗�U���K~�R���2EQ�S�T�l�a�X��f�~<�/f�w��a~Y6�*�C6����w�;,x.��w����n���s�}q���
;�:���p��ۀ:�+A�����f|���(����o���c��ړ���+���^ώ|��R3�F�DE��M>vZ�Q��� ��'�KdZ~��T���q�Q]2.���,A�}=�/c��e?����g�@�oČ)��B\'��ѣ������܃�⑪H
������r��*o��ڍg�c�$f3DB�}�J��K���6�M�Iݺ'%w��=��I�&}���0M
gH� �[PE��xNvF<� ?X� ���ɻ�Ӑ҆+*����]�O�vZԪ��s(g�@�|��j9	g��F�}(���6	%z�w��\1��/﮷pt�4lWN�bօ��3��yA�ܝȥ�v�]2 �!�F�:׸p�R�J�FM���yc�~u@�7a��4�eA��o��#�P��\s�:$f�K��[=�62��C����B�}I$���XH��8��u-�$ ��}����r��];�ר�B��9����8?8��z�����u�/� �)�<����ܨ���tX��ghȥ��]�s�$d�>�8��0O{��8������{Jβ7A��|M��G|�N��E�[�����b�,���Ұ�����j����e��`�n�`n6�ӵ/����|�lR';mY��>�n�0�/�H�e-��?�-�����AH^R�P�qT��K,'��yX��E��!�J��{�wI�#����>��_Gټ��(��H��5Y�"v�!X���v��I��ȥ������u�NCN�R���E��D�H[cx+�5��=k�̝P��.~F��������?SoM��j$7�R?�@��
2r�:ELya(��3KlҲ%��y�X6l�G����a����x�;pV���,���l�,����.Qt�op����=c�*�m
[C�PV,p�Kv���*�wbU�c(gs��o�}L'%�v;i�_��VgiHİ����}�4��xKF�沸�k�_�	C4Ey:!`/�iRP���������ҟ=A�{?y��95��/Q4Xx5ѥ���^Д:�wF�����2	٤+rI3�d`F�θ5��Z*�
s��jyﭮ�%mF�P�.8�.�k?��Y����/�ɺ�ڼ�JUS���p`�OA���9c&�93L�M���+�[4T����C|��@�!Ǩ��²�	��h�=��h;�F7�VT�>+�On�sI(�5�A�m���.)���I����w9�"����4% �c ���ӋOyJTܙ��Bs�X�6��ZڷEsA9�$H0QUv��	03���	�n�(�����
}����՗��C��N]հ���+dx��g�O�l�=������� �a���<�t��irB�8�-�����%��G����\<79�锭0�]��n��{:��ͬ<��e��T֎lv�Dg��I%����w��n�ޏ�N$~@�+ApY����l]৅Z�'��G�u��8�Ĵee�d@����#�ߵ�I�@W��T^դ8�:5{���Im�8$lж��FW��Y}��IH��=I1�	ԍ.�����b��C�u>cc>#<U�V����>۬N(���y�	��U"x�o��#`m�]�>XD�n%4�h��(���X[4e�E��C�"�u���
	�.�b�#:Ȋi�9�s ��X�ҳYe�c�T�d�v�V����g<��]�G#CM?��!e�ˑTq��F�O+�Sz���$ucƌ߃+����:q�߿�l	�j>s���2ۛ���Q���ɉK O�rU�Zt�UEONf�`����Q@;�iΤ�t��{�_sk*�Fe k�4�oN]����B�o�[��M��1��*�;����҅��1�[�Q��_E�5�t@%U��w�uI~�[RC���?t�>��\ʕJANq������i���HO�1� �n���1*4y<��M��ƚ���LM�<i�I�n�r4���C�>���f�U�!�bC� ��γ\�C���l�?U�8(m���4�1W��r��%@�����kR��}�͝�MX@i�s#��$'�/���\$���-%��Y[D��[{8�/�X�\u������E�=o��e*~8�vnP�r��W-%��zW����ԧ�:� j��E��������sKJ��K�K�Y����w4�!u�,-�tӽ�l�m2��v�BI.�E���)�@]�����{Ul�nU�?��%1�AR	(w��T�޲���>��t��c�8g�����D@�ij(@�M44�7P��2)�� !G<�S�0�3%s�A �DxKO�v3�O���r�T ����rG�e=\��=��r6b��J�{�f�
�;x؁��� ��`<�壉 hk��M��61T���B��LQ�H����_zL���!	�δo�E�a�����L���{7p��kÔJ��WA�)81arT���L-���TO�hP,��R2ck!��5��^ga]��\G2�X%l���o��M��C'�T'�%F6f;=
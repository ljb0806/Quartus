-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zXCGafN3cB+Fk2tShV+dzo2Yhp5rHXJiw080Fw1Ctcr+vMawE9cyH7i9Yc0A47/93qwiJKJedvOO
8f3HyKh7ECbZsAZEJHsmduxZkEXa7CgqPC1roNCWPz6Zc/ymVjrzzKWA+E+9iQpOXAiRbh62UXem
57FINJPtQJnZJIXVQoPjh08wwdvJUW3KQOld3pNAQzXOS3CkBQRYuO6yENOMwkjNi+CtWUuuMoty
fm7goOe7HiY9xCRuXy6UGq0Xbbqi/M9jAVtkM6Ef9QEg/Pbtvf7nAecCCTVWNjvoicAQ2n5MZgPZ
oZQwT5Ui/oAn8OSFcUHGX36pWIBUvM0464x4Sg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7520)
`protect data_block
O7EtCSQKqKVH787bcwvPzdNDBE5r1TM5Vc8/9YkKf0i/UgBv7wm6LMqGgSxzqAgKzvJ+Yyq0aaL/
wQym5tWEXuThjGdMwySmjgT6IwgbCnwkHBh2TjYAHGA8sNllDbb17R49vma7c2jAcWc7ZMRCP7DW
1HQCF78crRs3qnKLv7UJioEPRHLwWS+Pfb8x4WZpwP16BS2c19wJU1jkLoX7y43yrO/PHVdoPApl
Xhc4GB/LMEfBpZVtnBHnY3DcRrpiG7LwDawUBx+DqnCqbIIj1gPyFV/VPL6yixQ5SwtnDJnttYUu
cD5cLZWSN+eyCkY1hREe3ZaA22e3Ea0ZJrERSiXFYNJNw9KEBDhKDeIfOw1whPxxMdoxx8/YTTYx
VAWfNUq8HDpn0BgwTeEeT3SbSfGlUUL5PH3VX+tnTv1I2GXYpbVJ8AOphdavwLX0RbErIDPLlUSb
t5iXSVwETc02n9sdJTcZW6vL8od7JD9brTjBgAnxXNSCEJ/uVcp3gzMyrp45r6Tbimd5x9zCUOXu
FtNTO7PQO2gC28Y+i9/zQqJPbql6Vbg2rZY9TxzSAPpHFAykWQldmCeKIogn93sZ8M0oJZT1OOin
U99C734RueRyf00oi0Oq09C4hmpaeOoZRiDrpYqyXWtkO/kf8bkMawL5c/EU5hcKbMqafXIHbgqu
XQ1BUC4TJyF1Xu/5r+eoORfFfxWJhD3XTWkVMzcPkcpOTXcItQNZjI9G4tbt98ZQewVv+AsXnfkH
/aTA08Qz4nCL1SOo+30B16yaPuv+6Ddq6P6i8hRj+E1f0KahA42J5RSHbRa7F2Gh94amPNEj9oeX
ZpfLsWddvo3gueZWckE+EXZ4dfCELu8xN1mQ4WzHymUMuJIMlfgtdzx4bx6fx8hnp67+o2dSO7fT
COeTb+Vu+Qu2TDgpm0pBT6WLG32a7j0502LJeATIAe7MEyCH8g4aTwb2wyfxeg3PLHZvOQN6jUzC
45epxUHT5TrWrs4lmygW0S5gZhWbqxowm0r3eNxpDspqrJJlGN/Kkk0VKbfnwkgp88br6fCdjJnv
UonZEKDPEP3rrOXI69YAFxMcPXxCKUEPNdJWBLJraXuT/TA3KouE4kTPFDMLO8i0ck9Oc7hVtXAA
aTFcFQi+pjwCA5chTgrXudgm+1JO/br8A8LnjWCEj1gIAsS4k22xRuknxWJgrJTc8JxOcY81lRyo
yWgbi6KA767YiHvm4rWMMWp7MLqvFe7QMzY2e2Yo9l4qMJDoSnSfS+4epTFLsj5maSugww+TtPQD
3gCZzZWY9l+WXYXtpB4PosTr0lbfr4FVSi97YBoVDmb0qpWwM6+x8ItXNRguhiUrKUdUyyNTmh8o
20GEFNhxWgtUPtgYHIpcnq80xzKZ2Tvbg95plb4ZOyd3dD9iGzVJCyzpZzNrlBP8Z4WMgAyzSh6f
4A59SMUmCmMpnEwxWARh9scp8fOGAw/wNU1Mik5H6bHOSKMbwcJVJk5g6BN8ef0rT9lpbcGWHjbK
V1SvNyNPZkReA5kl7taZvCiZ/XedLa7yXYjzV1HOnoi26GpNshZvrYqcUwS0DFnpBnKyuSOIZn7X
l7NlykoMkfwfaxFhWy6S6L42nP4uQINKPpomU+eUCMgu4Om/tlAQUHSq5aO5M5LLsG69K0qmp64m
94LUXIDC+WNfn6MNMhwmkUw3EA13uDkUaOLxweZTAOUOA98HAqfzDdaOmn5Q7wuuJ/dIjAnYa76P
hxzL8XGUvjFOrQjnAY8EThRB/p1MaFn/Zipz/8mv4xvVIhgHE9qFJ+hGefNj7hAjGEkLemYSUwY7
euOK7uWPo2n4Ere2d6lgEzftNyZ24FhAd0pSykczUSROg1ldsKXk8fyFPyqXOBUDovpVgroun8xZ
SDW9iJbVUlZ5Zd4mCFUS0Oe0MY8r3FWEu9WEQworXdAp1S9XTiiMo68MrS1qQMDOabJiVwkNDcCA
BwcR37v1CfCPyX8+vwN0lCIDPfgbo3tyNp2Xg27+TiSJv6GM3UFMhwbgCurlBlc0MHM6HaduqULW
m9Vd1GCW2H+GnIh/GzuSYLKP5BcaEubr8pncNHNuvMjw/SsMawaWKpa6PCrzq2a6q5lqWqrI3xZy
/kaTAZ4llurb/22qFFmDiVKw3brEhy7yNUeCpoRBKbIyWsdDsIFvQKVxK1Eglbpt8GWqejQ85sav
+NYgEW/INHXr9bA5HT6KUdkwkKqPy+MIrZpDWVarooZSsXwT7/RgiuO2ubksFPyCChnlDPNthIUn
oWWXeyNFoGbTvAJUFIIwrTqNhNJQQFK+oJXSRu0Wz1lQ8/25e0TQagM/BcaZheoYT8kKkQH7VaWy
xW/VlEhq/nWW/OzgREPw5YkiOvU+3hj5wt1aHJvHAyF1CpeMGRWwadzK/wwjNwhGJDMsr6hqjjyN
ae7EvMotm7wEwLuZiFOMYWOHllAhTIEjxlF3EL9xHiKcpK2ZaPxGO5dBe/Gc6IjA6IUHAnCa9pLY
6ScmA47wm5paT2iSVrfddKhSA9de3SymIN4KQ2zpZddFsnu8/nr1NykAlzQGok7nZhYclNQVzpvN
ArlfxP2RiqQ3HoU0lJajkuTjf/YQcClR4Ypgjwm5/EcZb+Aos19x2tVWI3XIkF5DUMXwaptGJ8XK
WKJxX/NTSwty3djlgPADMp1aWhAtvlifKb4AlurrPZP9e7AiLm37mnsE9Dl+GESMYPjHe3Ebq6eO
paFh7BxL3zItHPH8r/9je150pmttvLDuoR8sKV/9eAqeJK51NFYogprBekCRC6NUKAwJbHrF9pCZ
861eYszwfn7LDfbWTi5Bjnf8qVFJJwO5V8dpETAAGFft1iypRPknWU1GCYDtOKuRcVbtCA/Sq949
F4wSkftQmgdoSOAvRPtHxV/ypw0axrySe46n0Nb+9vfg+1Dh6dxHHmLcCdnHMynzsqMMk/t0j3yz
wO9UOfS1Wb1Xfg3XXsp68OeeK+1kSDSm2Sf5StYk5DLSsn2L2jbHIe6j73A4uDlDQkgC00pnpYe7
5HGFZ+I/oZ8xm3zF1rL2XLsJhxLgJMMa1PMWIj/BbvBTzDI81n6acA5r4OVoAosd5EBVE1PakJ3u
N8IVsnfjqqWGNGDCQAIpPcspcv8nZxQVqPjMF1ATaQReZdGiKNtgjKKkAs3lqoirzAxBwwJvMzow
J2cildM4uzdGNaoFPQfyAN/5eH8D1rTV19ZLZD/FwZaXfRVMoxGknq8QCK7lZvRgEoN7ytBoKEvq
kG9ZfWHrXMqOMy6jwA8bb5Mbe/4lnLuKVhAqXtVy7rogbf1GK7Q6FFH/D3gThRtXv119rDFXjpIV
oUZZYJB9UjhKEIlbjkmN6OITvdzptByUUW4ouycpiAkmyK565pNnlMdwjYUh0LfwVBDtdZpIygWW
SLMMo+05BOMims2gfsmcv4O8JlftZOFKUL/V8q1KlCgrm7nsediZ1SUt/PcO64yzzSZoDTRrvqyb
8omLxkaGD052dqa+38vqoPfHCeZ5nmluIF5eHvYW+llGwJshjx0wJYq3cTgcsmRUhiLv0p05v6L6
rj+V58BetAsj5rs284aubT3+5AClToubMM09LimGtrC/t3wfBSYwmShzRE4oNiA1GaRA5o3NnAM+
Vkp/sa1VLhs4tdYTCkGlkcGyVge1rsn/jhkHJ/KhkzUC1wAmFzD8y0FEvY2xZegHKvcFRCojr3KT
BXNoYTS6Eb+UTCsyWQXQpdjXySFNLRUifELl6pTD62uY5xqMnGkKukxrfQngu6CQLIGmCz3WaBRs
hKVS5tyCoE+OAg3IdNcQ/oqGzIfdslXghAODDoRFTf6LmSbubGFOl1Ht7Mamppe0lNqBmK3YDK06
hRTL5L7Yo7yAWBVR4ig59uqcRt7Cjvt9dRqlNZZI6EIvqMtCrj31QU98bd6fcrCDAA13fKbber1w
HgNO05WG5Xlj07Kr2VQ5FHxB9n7SkWc71K8xXUfSeYuIhvh52yP9mtygef+GUXC4I/OJikAjZfdB
xcqZBihA+8DN8Tnyf56B+xEV6U261Tb875gKH4TDE6Vj84U0IH6chfgyQAGMEee+mbO66CRLi16J
F5LPQtiFe0zJcpxq2U7KH3SQ4MF0/NyrM1bFP6i29cY/VwvE/Vi1OEj7Iyb2uDGe/rKQLqjEzVxi
sO8W4WHBEmSqNtGDDHlBFs/D5213AjS/mawpwbJiAXy/2Jx932Q+hs4UQCoLLJR2/URqFod8zDtb
dS4a9U5lo23G7Llej7AJvnhze6cIS9KRw09+lcsI2JoUlK4MN4RQM6WKbnlOFhsPBkSquTNa5Ex3
c0T+U5OpDxU8OnxO0iX77BVthd5U6aGPkxSlxJNCMw5vC3XfQqjD//YhS0YV9fI2jt4nwrpup3iC
m4KBApGMm5X2fQEkYsVv+4xmykCssBkCcB9ysD/mbzyy7uIWDhnGAklo37w7XOVHaqt7DVxEHwwi
7npuWBRJSaM6KLHvNkjFDhLdzPcWjzjSNr4x80bWLDcupTCszkg+/aNvOeRSluD7Zdx9bDcWpbAM
XI9LvvIzpgS4WMz/hb0sTkBoGGNiY2w5IYYBYaBe7p3NVkBkR0Blv19/z0ieqrxG/59pRnQgmwij
wfuHLjdELGmEk89juoDrXZ5l70sVq7duvDhO5AWNTq7xo5ha50+czPmz2Vf1ew1abQdEbzFvD3SH
4Baycgfx4Dg7ENJzfsoKdIllEZPdq1cp49I9Ar7hLs2pviThCeo/G0rcOEV4gSyRTS5+hKGnw6yt
+oENJv3V//HauG3gvEIsUokfwBhvNFon+GXDPHSLVnq48MK1DpkFe6hfeKGPgBIBWgtbfeBvmfiz
UFnwKrgMdh0cTEAcd06zYPAE6Ss0bcG3KTmduS1tFepdsaBaVnT8z9LGRoAXe7TJtIe3096hXEQd
aCcc56txs4Mau9bAkMEq3/0Q4LcQE06unSY6kQGs+owdT1OnmmI+6hJ9NMjs8RN5RH23J0DMoCIZ
uV/sqD5gTf9t/NBBjULl3ZKjgFVLBAF6awSY8SBYta5WtTPi8sb5GpbYgQJw4KLwcWNOsDilICl5
MVHDX+dp3ECM0uCZUqaSbc0Pmc0Nr86IT6fsBsJxn6ylo/Ec4rjWShFfmPGVg+OBMPyRwTJw2aq7
nuPG+En5Ki03khO1XXwr+tAH9IPApdM08/q91OxwNdbgAvUGtvontUo47uZT88npaUAAVmaTstgt
MkbvK6kXrsU9bcfPoETf9CPdLwZapZ6jhPN2ASyY31eRvHiKI33SRfBr3vM5ijZdmr6CUtxxfrTO
hfCSuMrNQ/tsreEIWrJtsK5Z7ZmJudiV86JWtRUg4CfoN+PeOZb3fdWZIbPCu566zEWsX/IzLmte
7v++cFMDZ76ZKbcRJ7umaRpijTZWOvRwY5IencPGQXdPf/qFrsp81413wnIRrXWwSzG2wWjXexzw
LYCJVR42wjAObIeOq+PSvwOrw5ui7EKTa6q/00dmkpJoSSdV+u0WfWHcDgbMPWk8FLKG9huCHpV9
ETcKqcJhqepKLnh70y+UI0zMBcTPtXO+emVVPb0GZQBpbhz9LoWHfi9JRUSr4XMXbmOUTNxJ7QyS
lpiZYlOJRkj1vEs12tD/F1S/6eEB54D0jIHCjUu0gs9j4qLMephs5Y+Fegl5JAVhIGPEHzsIkvOU
+Tst1afRmdSyL6BXpF2Rl3M3TLO16q02RzXokelcmu2RskmFkR8Tb51IFSQv+CsI3dykhsRlfQAm
/f/CKmmYKGQbUEbll5vW6Pf3Zw7IBGRfftfSLSQTAkAJDcOUmQPQr7n11xdFbJArM2o89zvkaix3
YO028pfcPk15ExC5CzEIk/ZoDfO1Bnr99YikM2EXRSyeuT8C+4pKehKd6v7BjsfIatLxtZBqSP3U
zoVjfbRePJQa4mGjjYI2BW/0VBM4DYjIh72AxNBz0ke2Qvs7cbMxWVHGPhJgMyj/Sob8kiFuYglI
9iEvkNX2IQLtSP68hKeGcHTFVIHkkGtVOAX5lp8P3IkB/gF8hgKtKw2uwuZ4Zwmxy3kkPfTJu9bt
xnS/I50LS2n2thDmlnfNgdrN7WyKrHzWG6VZZX8LuBKj945X8IW3qL2wk2FtQbYCrIKphXHOQSEr
BkEeGOELmAFsHB3S9K3N1VGn5tx62lgwCKfV5OE1JShozJE/5JeEcY5gWAQRFUsZR2UKBMTHOYen
kIK6EiECWulyT+/INb97mQw3A5zxM5ccujk+CW6Lk4CUJ/WmvBfCvHlYRYt9gFXiBrcdFpw+ZoZo
h0nsV4HuEgu8pmsFzdZo4x+or2ut+ftDMw6oU3LkO3hh91HvIWPy0N49gKQVyqTVKTpwUU0c+8JU
d9pgTIwz7kj32OMHj61P5dbaN0+peZdLVo0kfH4Xd+8taCYTpdjMWRwYCLlk1OhdKoddyzxYh+lC
8/Lq+4dUxqC4oQTmSbsCVv7I4TR+LJyBf/r1sebhNWejVM0FmFfUUGWXPusrg7aEW16aMVaFg/WW
mZyBMn2bovrB1jWJGt4f0ulugFltBoBNXuJzBiWz3cA+wWgoBTMvGWWdP0AfBrxL+Ql977nAJUyn
czDljc48qxUo5ypl8PuScOvbzvyw3yEqQQAOWiiap5yLSQTsELNfNHaNWm9tEhryeKCk93SfGUq9
4v4f5oBRksk0zXRX8ZT9gzu+tfl9L0cIQ8As3uJNp7lkHiAAEafxzlT9gQCGo9VChlZM6kSQ/hSX
VSU9CkGM53KO0GLG+m2NSIM3XNjD/YWfdCquSxWK7KlQUii09mgKeAWydWbC9QS6GZtOrgXcc27J
VwB7/dEwUgJdvnwGmLwY+iFo4lHE8y7u+sWa9UAebi8dyR+z7Nd8c+3n6/kNJ10g9OfXaWr6aNPu
o1v8EQab5ImVG8MvwlrWp+DGpNnlj3Bip24ReC6OZiQutHTrqAxpCbVvOpyc/n5i/gfoahShIQ5Z
lEWU0UIlto8QGyS5RSUIjp3pO92b7uMrdzY15yvsfkFV9U3xakWz3dOmVET4tct+rc2CrKqpgEb5
7c+D0LVlec3Uxj4ifPpHhmgzmRKd0kgU7cGu1aRP6LU/GdFCsVCYP7VYEAU/qThjFE+vb7yLPQIi
TbwXfEoMA7WZF6/MGXDS5sfdM15gVo61q3VDo/we7EZluF0dQn0gwptBJ+9uB1F0Hw5s/pU+YFow
mrNSHFj854klLPS8UcKnNdzRFj1JeDaL/0KYsa27vFcjAaKLFLp+AiiI9nmUUo+Q8dfKGZkygcDF
dt49h3h0qeo8thDy7dQ31+pW9QSX0qflAXetSoYM2XPUOO66ieN4QQnKVv9qu+F+zmv2vts3Tbe/
/pkZonmb1g700EqPFArAHA6+T1r8Pbl19uNX/LuemTkJAplHgY+H8iZ/YJaja9Mr1KUEKPRr08U3
8w5I8moao6YkRsCoG630LiUZfDR9wuvKJBdJlnpOcHsLFWCznhY5hnN0fXiSh3USVmlell+ljHDZ
Tjwbw7IDyrwYu3X2wdvT2erxbGrBCSLbP20wogM0BH0ZQz6yGkmEg3lVjBGkVo7sZ8bUXT3GZeLj
R6sR/Fkp3WpHodK6w6lpxa5h1RjY7Ix+hAvM7E3KT1F3Sbdj16joHNehfM9vXbkjjtTTOhF9PKw9
mXihuf4eGXlL2OD2yUk7fH9C+ZpYisA1zExFM/t7rbv3TvMNBGu2wnHw7hhZ8c6QkCGka81saiFf
Cifn6xmID6XY2XBs6TAxVh3t/IF0WUNY3X0Sb5LoIUlTMxYuVM6w2dUqYjxe+F5YZJ8MywJBw2Nj
WsuMq/UX5z+ulwmGba202zaR9wrqkL7JMegpTQJ/oKVrW7Ud6YQG2Q0GQCnewkDjRp2vVrB5D0s+
NkM3frLI3S37h6BA15HcjAqgmsiUPPbfxdye6gxjeUvGU3yW1zQ4Y4kVtd8m3BtU6RF2x+4uYEl+
apjRs/x1vkp6KTLMxalasmYVP3DnzYYe3DJ0pyaEuXs8vP7kuJ26Z2GiITdD01OntcDATbadD9cc
oJgneTiUwfOSZpTe1ZGougt15gEBmYywKp7An8Yz3fzWis5epth21IqS7qgpgfdXmBCbATzdWKmq
JumLofBmxHWMHbja1dd3YFqkDC6zazQ+KMHu++CsaPVaiq8Z7u8OOJFNxlnmlIQWnMamYebmTuY0
1XVjAusRh8l9NrMKKDZQX/CRUmshC3NZvMFmIwU2AkcTNTwOWW31U96E9aIyQTulDGxtKOEojDKf
6nj9pyn23I8CZs1HCtIQBkkBsJz41Oop2sYbaPuqZusk8xrbs43+0WOqGjVjoQlz43PU8gQ8Xunc
PReJDuwDmvBbpghyam7O43SKy9tzwapYQJy9htIE5+pFzhlzqJpPZ3nPijBzBS8LPvv73PiZmoCP
mwAOH7jY1lrOgKmOJAXGiwTc01S4zbGvPOoN08DFhiofNNLr556rQr67rKF+UcxnZW5h0499jQBr
5dbXe+/QtEQb5ura9WQ0LNga0MOBCn95qXVTCDTQx70ETYcnyxXXwhGjHryYHcUk3/zp6LqtsAfr
s7lsKNsy6i1N5mddSVSTdlHNfrpxYHTy7/bShg/yyitMN9Avr70Kg2Q93umfE9HjykYsQFfh5RCv
QliqekO4zJ/7sE9ZpJZsJ8UmC14GArCPPgBBO8QWjnrkuXrDBz73ZaDxwyN/jQfn2SLC/1ps7xP/
8Zqwpr+3cWTvpljdNwLjVZuL0xZNkX2W1ohwvbZQoVRqb2V6pAeTshXU/5dtfBjJVuApSAXnj875
8TToCrGKRtvgKkvz2el1Jktva6VSLViPvxINgR+pQry6fCuXVWU0hxcWbZB8hE8e+zkeeCeIHoOf
DDr/hgfyJQNMXjkDzWcaHyoVC9MY9G9K9czyqbj6a54dJHcP7bLzDUgLZVPKzPCTSHJAhyuPif9B
/Q9AEFCL7bYMB1cOjJMQe6uDI73btoVFJnKJRK6mu02esEADmkvRwDq3vUhG7DWcoU/cwYqJDTuF
4HrrvmTOcwJSKNYpT/jxWRd+NqiTQYZEpbGyRp/EgTbrNH3DdcJPQZdJKZ2QbmAqz1XGtzw+lUeG
+eRevKQctAqP+NW6ukeINXhj9PkvoY0ffhE5XdryHwEsIc2t08C18j99pKsmoOxmGX/q4ZDNc7c8
wygNySmtbrq1UbIIPuYlsR9mGVKAeedKv9weQC53gmYTezhiw9Vnts5lWsUj3HNf0Nr9e1t/SEpy
5YIV28+u4H59j2Xf4aHucWRpVkVao5AEIUDz0Lnib81fM6Cwb11tx8rsnFcKVGzLZwcoZg71rwYN
jYqLjFtEFpA55vrmuCuqAIxw6hlWSHaUCrbVPuEa3IM+C06qdKfC+MDorHv29y0QyfxjPuvSYUy2
yeVTtRbm5QuTd5znCM4uOWYLKI3oqe3hQEMefKndZ8K4oHDdAimE5YFMxD0KEhYVsf5sG2ITfjjT
retUqGrXuEj7r5BF+md1Ds8pjAZMVBP8kRXl+nhoUqIoq4I6TSYj0onVAnTa8rySV7bCTEwIIWLv
GUUpog+safvvjPJBuPcB5kcjww677zEGw5nYY/I30B12EDio8yRpD3wbaJUaIUmqXR6bzUBclqEo
m2NziysgE4CupmF83A/pvKaIQbhcMwEsqHA7FqdZ9387IwwUw9lYwevXTL43S4b7KkerGzVadP1y
GoQsSOKV4BA6i/FB0Py4Ug2HXo3ivo51mfZzCs+crdlw7Zu+nbPs/ES8DN+Ol3lLfpYn1ZbnMSkA
d9e2oA2I1jJR1Jcbd3f2Cbpyr/Oty8aEGi/d2owyP7MPeFGMoYYZ4/CbNeVg1P1iDYM+jNQ4OsX6
xWafFqSvF7y6aYxAhu0hwxNZg1Nm7DQET2B+cb/iwIvyQVVWn1u/qpPP0VtnW8PVHBwu2Gg8MUXo
B7tpqe5rz+LSdcnGlyslTUD6AAA9cjhGOSO3h1oD+DnPh5+SBd3XfDAgkxvtgU9b/atYU5s=
`protect end_protected

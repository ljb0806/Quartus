-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sOrmSo10I1O4q9/UFzvUaKjr/uqgU1nTwPJLR8ombVYYr/OPcvFjYs/4avtCugSsAw+vGNBfhmtI
bPuPlmuhJtaC7Cf2jq+Zl8qKOU3RojEn/CJHy0idFgZ/8nqENqaOLy6ck7+1pTMaEMDLTf6Sknqk
3qegBUK3o0SbV4rXhl9nx39ZUyFp/+itj5xjMGqqseKD3yBxvMxOLnJI10dqnbl/dP+89FYRtJY+
PYBtqWy2NCZ0P+GLyPLPPmsYClvAVx9NB/XpxEuU8QStv7gI42xat+FguswdRcORv911SV2BhD5l
10KQUyA/Kok6VsbhTgNag9KstErUuf+jXZRb8w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10752)
`protect data_block
Jh0GVz4SgtW8P359WlpvgDcn4rnqlx7GIunNylJiHS0aaDruykfM2t9GCxXJCmefxEMcSMp7l7UA
4xEzj9B4npCkvJpXoF9O3hg7CfaNxQhUno6AeZINUC5HrU1KyNztX2cWa2PLWL3ECb45WZMA/W6W
Pz+iL9210T6hTtltUOWuWAMdHlX0OgjKAcLyATXDWNiRzkmIZqTLvV5wlY21U48F/6g8WmMcFFi3
OGRBdSi7ozq4Ofa7OzmZ2hSwLkn0hsPiVa6rbQxuHnxs1Iv8X0NwLboEiSyPDUpRqL67VLnfWtpc
jRAmfDJ44ULGXnhCdlDFvvavP10N9eJLxL8H6xyphixrU9hVMOW+YS2DNm7B+6torq8dpHxXD2cb
tJTrOtWXN5dnzk80xAXPo1A1uRg0rQDcLzDelaNWwZu5OQpUU9Cu0ApxFmixedJ+A4NSiL0210Ar
8hBJ/I7v9aeOe9ZXj5FvEHdnw7258eM7Fz/+x/7NMn6sdbHvOL8ia2/4AQ0dpMPINzcQPRAlWKSf
yqgKCXrJsad51ePhWrWYrXlut5Lc+O91gs8ypcjq0QzH3WN60Fnei0HDvvzeCcoLEqD/uK7PjXTv
ykFfq9S3M9DG60m8HwIt57ts0aiDhhZVgnPJA9+K7Yv/Bc2hbLKxZXr5Bg29/00YyMIZA4pRatdO
C2EF9sw5BZeCrn3ky0XOhINGLWsjCcfsx7gRedOsw/hS/gnH98HB3FKh3JIvnhRTL8uV9SuZNU2z
RPt8bbTF9bqsS+TNy6J8FoHaM4JKSf5xM0uUwfaDFM+eS0li/yzzT0U4w0VaDjZczQYHcsoFn7GE
I2076QM/MbSQSX3NfRchibI0YxPcPi6aXrsWHQ7CUbsB+R4lgkFG91/EddtZNBwEXPSEuEbai03r
Js8QGUYTCmoOTN2W4wghlF/3/nUnzFxzSS9LRj3bniOcj6JbWnQ9oP82yUxd2Rf5nWXOpIa7++vP
xpL4OQ9iemJDpUCRfuhTZg52qO/veXfwgeZVkX5O2YzwlNP4ZRTdZStbWAMhMT1mHkZPFrjof9eH
rDjIz9qgbkc7LOAzh9IMVQKvAYmXGp4vq0xMv0Hx8RW21VdNnNQsoqHIibi1N6RJDPQFJ3JZOORj
HFkJ8lgKAdzO+i5GyyqHHmu3fCQ6Aj4aVGGRQxpvZ0FdC4gfk5IitO3euPM6XxoXezn2SGJ2hj4p
Wyi6p32C7gZ+eB3sAaoASvjQlT1ZhgOgsNTUI71vKk32nRb0l2wrKIDODldhwSFo9FMWQ9p4TfDZ
iaXaPtOhRuUyhvRd4XTicuXvN9NVgwjCO674H1bpSl1nwsi/i0C8Z7CL+zG7zSaNsWetpOcj+SIn
xpf+fb41HP0mEZY/FlY88IfDIe/HAo+rOGB0cQpqQm6Q/h/Um9YhbX8x/kOfvKVmXnoCdEN3gJe5
TDs+Zuv7N70DeGRIV5gJfW2cUIXn9XYv2kIGjFN7qLBOMP6tV3T3wEpzgbD0n4lMkkvXPk1ue9s7
IXjhrDVMOQBd0UpZU2iM5D35exEMvOybVihVhEPO11/703+mgW64F84cUksJKqyMLN3UVtAFQAl/
6gzE5u9gvoXaebzozhRrum4DQuKAXpntp7IJNYXpv+R/21CT/GPnMvd2VZ/8XBgBen7pgXeFb3sa
n5JmEIdKQkB6vY7QvQ/IJlnHiWkj8tqsITHXgQq5kAQrzaUzgSyeUr0kvorEWV7c7CirYE6p1a6m
Z8jlU1VOzWkKbY4WBS3+lo26FwEuwZjrR8FtlRM4Z7nTaoXgdh3PB9vcRK0zjayDUvpovQe9g8Na
kXYVlt2W2oJVR3qyS7Xj8GOYZWojR55VjEDFJ43xOQBtOalA62RezfTf1LMr6kYiWl+Jvft5qifF
JzVt/RKGzCAtHbNF74me9u+rxaRUQwIm2OPfXsDP4HiEHYXrJ3lgacE4kE+TN7+muygo9QZSZpn6
tNzU7/gOItJx/Hv1eUZkUz3f8kkCO+BHXoMUMHbqZ/W+KyIeyPiq+0q+qQrLzl2vGkr36ZVm5Jtc
T7/ThAsQona+nmZc7+A1YYk+BC3x11DKYMO6OY16UKX923JQ/eZP5fiwg5xUmjDZM+e9MaoveZBl
83vJVBGYLAcB/doBSpkIj3psU0qVjDi39UiYzQS3nhef5Gq2leHSLiJJWNXhA2Zg/S1UjOrulgJH
MLUjfZalY3xdSNHDGD70vKGFepvnn+Hs4tOK104M2sJZUOLr3kDXdVBnpb85Lx55eIyR4XNJwB6c
aBZI8v/Zs0VuwAaYu8Qzpy/bnWeywMcaNAIxmWJN2bHtkkeBPnlx0B+E4zUyU8N+Su+042KnlxCi
kpJZwiAhOUxfpVx8jivBsPiFMshXi4TeBiFz3BNLFgNw8UJPxTAttoV0UC5l5hHmu6MVjJUWlvGf
wUBMvgr6zd+yelBwn1zhjiE0SaHaDMTc+0oAyUBw9qRYe6JXxTQyvYQyxkBpanbLFyHuY6QOYU15
uujcml60siDU2tphlU9f4C9v6tsp69j2szJcZWGIqVjCg7q2ViQ5iA9mrsfI7Wlx1ST5XQ3lBV9w
zksX9YqddeZqdHW4+a8whO3miFhituoMNb01xJ7QxsvXO3OYSSo2sns7yZRL4yWKZutxNMQ/vyMV
cH++l5ByEDshvsiVlK2IHe27prRKEGxL2PimZkgD45b5zwkWO4sXBGNtvlLhfbxD/f6eBIP9V51c
7CM89XfZBIKfeUqldzQut5TZe1xmYYjnTYWoPPHvprxzARXkII67UKrf0x/7m0Fbl1S9J/hFS7cC
gl2zbnvi14jw+1NmpLfwIKBraAMRK+cwH8KD54ruz2zJjmSh3juWWvGPuoMP1HlpWz0nQOLjx+Pb
kyP1ZPTkUlifmbr+vXXBEnoVMm7irZhO7kfqssc/EFljfTw62g+so2l5HIwteSNhkQ7RxAKurFgc
u+zvqobht0sYznjQGSGPqvqnuT6nkofKxicTUBF7grGQDHGJbTwUDG1z79GeYynvtWppn5VBTiAg
C82iq+Y5nFzY7ywmUbXgerpFEEyhVTcNArND1Eqz8IOK+MsTB7mKxAW6yTjSyZf3q7EEfUtp7b0M
wUhIENklVPfhYZs4g8dMu/rz4HrnsbQtzr4AsitLSgMKUjjL2bxgAWaocI4Tgb5zr8OOGQuJidXp
LlFX8Vzpfx9WN1KrqIOBtfrM07lX1r0ts853wKIkugzoIuwJMcusByHCKyn0BroW++eY2JPkWrOS
Ea76L3NS+SMElHy36XSKHt8OojbSv61MK+719x8+KMZJj71qywJcuQvtfxMYhpon+tORfpQ1GoYM
mJTlqngsayIF9y0jOLil4Egw52tcZx/Ff8Ed1oCTC9NBy5peHpauxZJ6tHFJYVbIJboNwui9bx9l
mkJK+C6hB4mYhLRmoOwCsYlUI4XoiHm19tM8IquxBTAmtPnCwUF8Vj/nsjY7+69dg0/jfzGXnt/9
KSOJusPwaCFBojTgKlv2DfNNqO+AdYsuUUm5BV/k12iuPZQGLDKh/sagcDgs+lsdT5z7FwiyzpV/
Tslea1dpeamzc4lTvGcd46J8ZglW8glmzjGP8M+jvfTgyHIdM8yT7OlPnGn5T1egfvPrSJrXZyQ8
qGI5V+gtg7wnS6x2OUt3fDgSQurSGqnVMNIKnrBoaIRTm0eeYLixEqzmhWfXR5WvxfmR7Y1u+rR7
NWSW2liCtiUAPy1bHNopApLPnw28xQWCbLEn0OBHtcupRsU7w0j9tfWFfbonCXp8PZoxjePQOwX+
IAm19hx+U/5UE+cFl4kBEHp5KtkidLhPDuiapg4MIuBAu0/Zl7iF8kWmXanXRDdn97F/ZB6BNet9
2XeYi+R6mTYnM5q7+3nQYxyy5C98p3ydsAdeHJPLLgyMHVidfhIRk9QV2a5PZtv0mQ1OI6jeWUhz
UeXk4heXS1F2ASF0RaOcU/QqZkVsR6OOj+MZ80lBlgkd2e10AeOpiN0ki9quNZozZvNlYNmSSgXi
RUfvpdCmm4863+Y5vfH3jGtCM7z3Rj9xdH5H0RQFXZauvgLpo1toPMbF+AKOzNuykY9x9DuWG/sw
fPtiU8jXD9TyOG+hBfXCHfaKZOrnkewFcUWUXpc91QwUr/4vhRzt/6gIHct7587S24Mkr69kOnKw
ttM2hTYOE5u0Q5cNAWLcjd4MYOwYCC+sy0JDp2diVyxXP4m3S7R9HfiFhHNZazkt1QuE8DiY9E3s
z/AhRTep79FS4CyYc4NF51760RS+iCrkhHEI+hBspVfu+sUz8nj421p+IZaN+NnzDR/+XvWvVQrl
X75gjWObkLa5cSSu5B7UTpbEQXqvPf/E5vnpUUZOMo1wkxi3KvhUNGoUAna0htEacgNyshjgCUXI
CasETh0VSsdlKOyT0RTuwps70ow1L2lB/aelcTKF0H9vk/vGF/TPNxV+Rrkd1ckotoIpP5WsjmZm
q9dr4caA9G3T4ygGhVgM/nu5FjdRXc8cnukdL+jjZ18C1LTW4xxvAu7CojDvXXwW6ixM/LQPQWu7
ar8MrHdIEu9QMsIpdRbpApXQ0BgtryiiTZgpSdal56kBHoZEeo797hBH8pZzYT1xK97uiDePBYzZ
CYyJnznUKQQHVDgrhFAHYiSdFpwvgaGF5v56khrZ4FA6uu5gXH/dYEHoGbamhErOoDc5IgIXOryj
CLslR/nPW9wPxk5HhGx7GowyBDdUiQG5HnlICPIR1HlVi3CCG5y+zpG/ALO9p1XfSqx43vfTgsh3
a+FuIz/8xpkqWCxBfWhhFPazU8LrPbVtP97z657RTJMURCwC1+aKHFdkSP48zjjVwgK9tjf77oFz
4SNe9yDSzAx9eZQAVp4RHOTl4V1H8ynJ1o8TxCPXOMhOlmhGD8BVUJPxnivbwGzuZy8s6+tIpKYp
XiZ4vS1Dg/MXJp9j2+qj/aMM+ngmmYdWmTKOaVgUAtBnFmLnuP6NWfoz7g36DPUpya/8kqo0TaO8
iSDZ0i5Yf29OqNWQM9/xILToT/igkCJlEjBsGVv8FL6rGvrFByz+hTyGgmbxoypw9XVv1QTHF0rj
/iJqh0adfpEQWTKwQiIwRivc21TZ3/12rbTlqMEY1nDhhSKYhj1wYIWthQucce8V6VTYbw5oJYIa
gyT4FgHp1fUApvnY2DkdkqvoioKG+g0nLeu7pUGv0Fyiw1W4SbJe74tM40bnll+JN/A6EZx6q2ZG
5k65eGMhz3hjci2gR7k/IiIomLHMP/2OwqFLAdh/zhBZg2Fn7nhI4nBk77wZ1pXKCnYVX0eg2M2n
Ce8EMK90cXae8Hu3fqmDFvSTajv0ekFFGhragL/F+Tn4+g3MyiIxgNHUDCZtLdeG/kWIv/4T+xFI
o2mlkLwYK2//34TdCufmtywlL9PeHBwxR8CeWOW8M5flsL5aqliOLOQP8tl9+pWf/ujlx9w+CUJO
+9/V76d3RBi6aOHIdu32OTf2LNxaP04UK1Qf1+37Q0cXe7Ao5os6M8dCEWmBPgPAhcxGEONor/yF
FfF/sgb/VBKbNOy85C+r6mnMKZhoaAyzCbBuXLVlLqt6z1oJq5Jm+ewrFui8/4KQhQ8HgGx1LsMW
gl8zwWJ8lLEdj9iadJ9Lcsl49XN6NZuRtVnaW9xXDByGSOyE5nhrZl7l7b+6qiX1g5Z9bA61Q7kk
rHC+XmSX42WheNfU5oIQN9BHXGxLlyObmQ9/UlZ5apzZm8A7s4BJvGmoNHm0v+RMcEwFfCw0SnWL
jHBPxNPiYlGHdk2mRv1Xmq+wc4KbPh+O1uZOHv7gir4hs6VsgJw+GIkkEn7r2N1CjxQYNideHJ15
8B3GAi2UskbVODVTLNGF5QhJIBpLTA3ngSwNwymv9v9N606hXE0NM6aDM+qZLx4SE1NGij0gtg2S
dxI93oK7oLmSUr9BFx3D5uhDVxX5HYCo9mCZl+UppB9qjj0xnRjKG76/kYzqlfEooDhF5cEg5z8Q
fi5GbrxvNlWqcLNAxiJcA/QPbafSRYufp6gc71vzg9G5/3foAfZjIz8uP6kyoxoj+fUd/+EN7TNL
noU52tTspBEAQv26oDkFAdtbFcIcsTEy/CvXRIFsgkpwpB2GwhMlizDXg0u1s4A9odoSBvAslMA1
aKOdUTjZfiwE3LTYdcriE4LYhqLyCEcsn6KkCYzSphl+CEqoabn6q2VXo0KguL+kRABZ5HjLlfJP
QUH9D4OFNE/lwJZGYqcaqBP3vuBovtjXbWdlZzvqdlXlwsgHdaMJIS/3wSpurO9zHqcE9HYTvJYB
NQfyj6+0+7C7Wy4aCMN0jBMd+z9LCPuAxPOv7V/NGZ88BsA8y0raUNjWlevwhdc+tWJojuxdvgg2
ZkOl89EfI3+FhLgyUxXKh0SW16bhDnOJzCaQSRw2tgLhuKZN3q/uMVHssYvuOZxouLXdnQ7Ed4w7
PdJ1wBEa/LH438T7u7j5D5zbAeKHoxxevYcIKVN3kZYthDcKjQaHrtW1IW7qfgmXoLu+bLtRn5nz
7YyaF2U7MS3WaoGlmvfLmb2gQyUFw1Cii/H1TpshCK15LFjYTQ+BxLSTfzU5DRIjjHzW3PTjDZ/l
9KC7rR2RYRLu327Sb1u0y/0lF5S4yVXySGgC06UhEu8kJlCXyVr6fN9Idu2aJJCXwKyBvKiiUeuT
ENZC4XOoS9Ez6BNf4yO+CXX3xJvlU71M8TGWBKnGD5qVIBAWJ5B05CsRp46c9o3+iOgcRlgh0WXc
EcK/y853ze8/39nhYwGXjdSx7027UT6e5dYTyu8LjU/6qSIhuIz4NfaRDKuGO3YymnqB6cel9Ox5
COmdZKchTA2JXn8QoV3fpq0Pk9HZ+tvWpk+NZO0rwIgd+mBmECnfIFqN0AO7dp65fs7Mgo1OZRYG
Vyb1mC40h6aTCOTcnboCvyb/TIAB3sqvecok2oAKQlFKm+3ygLbGW6JkerU3SERMQYwt+reAOwb/
q65CYbwP+4y1+lwP1Jz9xIITu5si3D0FGXnM86Ghj8x9l6a6UqveRk91xIZs2P1t3qdS0a2IyEf3
+tOFQJqw0ghKjW2XEy4j71I7OXC+ykFWOelxU5OmaG6dFT/oiUEThCZlKjjKYy3o0Pb1kriJQEeV
InuU9haeKtPm3hsWcI8ptRHZ1l4yYwujjq78av5BbjNpet3+MZnAyWM2VtWe9Cc/BsnolW9rMkRy
UbZ3wXksY6dpO1ISCB3ee39x+QwCKCPj8AZ3adb7udDH6vT1srsUII3bSpNjr2/JBWTzOcckOGB0
SCB+nF/Mjq23u4RZ3vYew5EJ0NmVjZAwUEoQ2JzW63dCofJeWIgWbIujqalzzyMQi/Q5F8xh4nwg
Cp5hxE2NdU+4y8nK38NEcncZz+TODK4EodLkx+/SqSJ2LUVjd4cxiwS8oqlt51VKLdkQUYK4KMwt
TjHmFXgn8R6UzmHG6xniqs6tll6SDnqZmzQpvd9QJvbcyubmg/Hv09S8UTxFe/KGg4MTpzZTe8BI
/sM3AnssvlZdd5uNEWG4TMpkARq6ipi+sTwUazYFvkIMPoR5ET625W4uWQk49yVigUUnuOf24cfU
685whdsb3U3ZawIpiJkJW6gGhg0wSjurIBD2DyA5mDcqMN2dYv+tKh4yNT+Og8MWsDTkwuxakKeB
sGGqFIOAv2/X5BQXFCH2I2lEF+MHB2D8JyxlrQG/KpduT/3Va9pzj8kOQPA52o9efE4dfhp3DsF+
WZgOKLxrusx+Jmj37eByj0uKmhGQw6kiIDM+2sbHHipWJK+yhKHMxfkgnIqyZMbDNrLR5CSELFOt
7mOYpxqzxh33pS7/vkppIvnX2IuGPHbdTnx8HuKcl7qbVfZfmngrLwXiJN7gC0uXiBy4n4H8KQoy
0DOtJlfY5zzQq6iM1H/WEGAQmVN37F54Aog8jz0JlKGHnjWjMojw4Ez0RU/K7nMmPEH86IWziWFV
EUsPcxP6qtTPntulmlcMF4Kxew90/k2byrqJtc27XUtHKfWaDO4plyo3OdHuDVvLHjojnDndVutW
UvZJq6oE118H4QxN41bcO1M4HoxuyudrdoCg7n7KhIaW7IT9UGf3xkqwh5dEaFYp9FPb21jJb00o
TbBXM9vndBAr3VS/UeJIBtRTl+7UR8ZVDswJTJQeCPC73O1OiG7QkkI2L07M+XiGTiIl7Wmf1W1Z
L9brMZOr3aHT9hIYFF+L0Upr2/S2vOwSqpiMHx3oj0zMqqeX9F3xBibx0iI8ZVDcFXjfYgg5yzTu
WjaD+168J173bOfqYS7GrVk3k596HvIG0NQiOpHl0rLjwmo1mND62OtMvgyyQPLPmY4DXNiwL/Jw
iNuWCZ05ULKUl/SEn1QNOe8vVDx0KZ5goadL5aia73SZ8/ozVtbrU+9LJyHTju/7def+7qUzPWnI
ZKkvDMkslEo9nlEviMhOeUyLkheMC9GEMhEQK3rIlci+ltVQRYBSzyFtIYQn9wkBp1IjIn6Q+sIg
XMaadEUabsq/iJF6JJ4Z3FuyTMOe919An2ysFXKyJ9BQWP56lMuXQf4nI4SZTZREoZrsffKP0UDP
/1T5o9rAbAw2WjxXLSNfjA0DSDBGPyu067JrYUMaPWOMa8HoGmQcT3LLQ8oaH1NuvFzGFbabcXdv
riyp6QzLLGY/qD4AekVn1CB+KtNQy6QoH/f7dzIu1JELtpZZEygn+L1FsCnNthTClS4E8Lbm/0nq
vxGAtfFxuBAcUyq6tRfGmvd6J1/c4bNx3dLlRZXBne3kR9WOtb/LrCq7UfIJLY5TFnd1y5+cqRNW
iYE6e676qa2XVuKIyexKxO9KHwaEjSQXiOzCOsBZbs/zK7CxiH6hvi0UxMI27x/4oCINslRnujFz
Y0LsN4fqBwmH8awDWxxvUdRh2y5dJ/aUg1j2p3dV51O5u123e/usdoARbBRN1H/Dc/tDCbLgifQD
Z7SyFj8OqlLh38TZ95Og5evlT1/opp9BcI3aqqSP3dnIcGhpCF3rsLvz5qT3yf6ms69T0RUNL6sx
XsgolymZjOPU1RdZ9nhvBqV7tvbIRJVx09OlNd2wc8cLjyXurZq7w0jn0J1Zp5FVsJEa4UuzCHBm
uuYhcw1tyZXhGvY1nr+Wa5ua6g/erdOGTItqe/PU95P1okm4V9PBrJi1rhZYqpc5RWhSWKNu0RHj
1Y0CffsSfaKwS28jqb4Tx+CYw+XYvmKVpvufShxNsuYFRzTC1qv44Yn5+Ugn3hJBZw+6JYBiCDvd
LLoMmoPmpzEg7A4htvZTMun5rG1Mp8+Eajn/BHi11XN3R/uIlQ7JOUkT/2gnvXN5mypgssyzYzUN
3NLgSbXc0pmMSnaBSaP9enfCpJMCXx5LlNzhvNndc0tQctcv2DuMu6RdikZxqjVqLF40/S87IFQP
OsNE6rsUdPt8kOm3/DfW5KyOpvgbs8QYlxrqxlrjQGeBHDOJlwRFHLt6cXsQoEA7fF2FUYqIRhSy
YmeyowvCcIAjNkOy5+cyo1C6wtiVLRRRMQuwsmsedJhBWBvrndHaU7pSTHi80npsL8AHJ4WYAB19
H5YeeUfPlZiPIAUJBV3gb5sYIZcTpDIh9HuHfFdkXxGRx0AtZWCULXGNjzbhHNOPcC0ssjqGFqq/
JHsJ9XeXr8tTEuA25l1AT7wXUOsv9XBoWgL+eG/psMkqxOqj61VQZrB3tf47T0V1z68OezT0h6wG
I4Y7+GCGGZHjpMkECtWTDtg37Yrd7zYFVPR7ii5DquRYJhdIyISdrcowEjbjVkNfUbqWCk4JG6En
6YMNq0diaNQ10kwkIg+4Q3jXG0ZRD/eRhHmtPzqKCogHMiBXnkV0EWELjqc+t/TCHGZyaIiRkFO3
+EhzRi5ewVevZy4fSUroR/XT0m9LQdmF8kNgmtKo5qEZceZyGVGmAS2OCWhtQG+fFvjKRQiSA4dz
FOVOsb1MezsSQ9jFNJA13uWZUGfj3MuM5P/IMYjgVWFGVX/fM1u1um3J1tUzjCSkZ4stqCF+GyvJ
WiQQzcyMDFV53VXGdfVoYJuomdsQEUjOk10nxq1RxH1VEStyKX33nqAulVufykyl3Uo4KLJnGJJI
0P0WR3yau2qCHfdt6NpTBAMk4+L4f4kE3Q5XA/CxhRpSjgN1cpjZb7X2Ra+GdSJYTu7Hr+Ds1EvF
NQnjRI13+8I9kzPklFb3iO2eLrUzWXU6upKU1eDn9ehKJ9tINr8QJZYzSLulk7CvjiGOcv+b27aw
6lxxbCqWkSpqbZHPOZVfqmSWPwJ7ejqKnkGUSA7sqRzb9Qj/JXwY8x2yiUcfqufFK1xDbG7rh1/N
UMLIGEGuKrn5wDH+WRBpxAjcBu9XtY7JHcaBPUm/xTZEsid82rN0RHucFvBbptrSGKQqbXks8LMb
X/xRmf6yQt1TMCPgfAN4xVbLsk/VmY5O+BbiosTSxz5/WwYqMBnOeb1T9dtUo8drhDevMrf0sYD7
jKhtzoMcFtSK1uaXpoRiVklUsHBA7mYUnmxqw3kL1Cn5GXGyDLWI2CQvDBTZgLNb2amiNyqZ6qPe
6Gn0NMUxbIZi1fg0+iX9VDMakWA/aCnpYDOC/NnRn6POpadT0XFWBDYNajMClcM/qrdW1ZbjlURl
NXqtXRWuq2uS1JmBztonZy5uytPqs71uC65YmRC1iDF2gJS6v0/EFHiTscIWFQS7VEtL4aQ0xpxN
+taZYGPaKQEs8SFvaXCiKvOxfJA4/9hYyckRmafioAze0gCTQMYRj6yy9Q1J5srQV/rVLnfVRoBG
eyTRUyMJQ2exVUCy+iqhuynh8CQ3KdU9v5Dc2DkCYQiw2ELTVxILZgDFN1uPtE/PPONoy+W3cGms
8x3bzRovQ/+v9Uf//NXGHBLZ2HebKukkl+10/h/HczDxbWexgw0PmXiXiSYpAJ7K6G8nVW6ahDB0
6nhFKksRUVg5/d+E09AuNiMsKmHhBm0DyVp0acuxFtz7O9usftjwmlZqHzXQn4GhU41uWlAUZAes
3R1DMo10eM06p+gI0pq9APjM4PTN+NBVUNrqWs+uLF7zwBW42e6GPTraVi54pEomP/LiKt5Vl/C9
Iwwpx4pUmZ4u6Ibd60gbDTX/m4WtaDv9u4dKDggLLgECfQO5fuhrjp+bvMU/F0OQNr7PV5v62P2i
5KzyB82M1aVUqNpq+tAREKuUvl2nEzp13kLl1Po1A9momVPPizRQzf2rm7pISW0798p8Rmgge4Rc
o0TzgVCtHpGflSK5zQ8XnBCyLhLFAzvmpYcROMlNHfxqxRR+1MiGpDQCx+p0nS9Mdzxlyk3WLnmz
i0J1QSFkYtYK9/WLOvqunrAQnV8xQdu0Bs1juVJWcYKIZpUi6dseNySK8+h9g6e6mcMvcLjr9FgT
41vFlrAcnrzlpdjsDTDUZbBjUcK29xZJqmwoBASHISNbXF742fg91CAX2kMVrzCsJGVQiTlcSSJi
q1DUUuPhVFUCO9PsZxYrkPIPW3rkKGvlTKZNVeNqiv6fLZi2Rlfg+B/lFYEsPnXuH1Ek74jliDe0
CaYapHmCT56uMwh3eu6hmjj5rJQGV83TksxG7YQ7PHagevAa3HFlBRK2lB0GJHimEwTfUc9axhWZ
h4HZlnHI3H+oZvRNoJyMJoJv1T9FzoCyuPFSTJ+KJnAbK32MttEcHjSnwO0miWj8hXARpCrxd+VC
hu+jmCAHnlvSHiNEt1INXl7m2CUJkhF7eoLtiy/Su979uz5NR63Hf1/794JX7CHWSPV3AYYJvfbr
M/pjfTKMQ5K7zBTRoAMnV+i6YacUaS9jBRW29Aj7W7vPR/DCGSGN2DAMR6v2b0Vu/QFVVQf0sjsE
3K4S7OsIArOQ90xs6CHF1kr//udNHRxarnoTrOc1EieGIHzptMA+BKX+5vCetq0mk+QrpxP37V+r
Y7NQNCFwRLdgZruDRimRnfa8PE563C5sgAHJhdJF+II6Z2d96tWFkIESCl9nGkvGnflHQknFiXXY
J+dpaqEBGXeDxLYfeCiRNmiwebCDKSpD/UHRQx8o8ETC7GViGsQpXyvR85FTcIIXSNfufWsGCdmj
2I7ecr3RrVMAs1ds5Z5b5InDiDaZppPovC4snq5fczdUfeQSY4WgSVA8tO1d72HDruNe3AUm9Ymu
E2zPYyAw6qS6PbquLeAErj+G9REAuFAnXjyOFEwqZRanyZ+qCdQOUN1PIqGWCP9F//ftpoOxTxNb
JR+yZ15QJmYBTOjtpjUhhFAjJ4WCYFiAeaZUQ7cRTpoG98POKTYOEQG/BgkdmekhSbo32m0Wo6AF
6o3IChgBcSxT4qRNvD+eu9MR2mb7sZ4+Z+hm6DjskCXy88nJtSpB3FJujK/pSllY9NvKHXfgLhng
vBTgVAYVMUopcKagl/laCvBEWQ1702wEkDqbe29oUgMT4QOtTPFwbQRb3DKNi+03sqtopmfqh4An
/DnwxmNyCLFFzeqEdRGLs0556ThXLlyAyH0wSil0Q4nvvMxzIZViZTiY/Zes2kv3mt+fg2JeAEgZ
c8i/w626DmbSzJG6HA3OdJdk1dWp0X9w9VHZY2oUW4WBkpYxSENj7dm66Ozw4V5gAGK5uW1iE6lu
rJPIHh8CnAlnGu+ZJ6PahAkGnh19LixC/CUWBZ6WNL4kN+76WSnZqVzOTvMG6UGDMeHHpNAsTam5
iWybJeUXNkQQvU2P6g0t3+k+FqmEWNLDfm83lhxWfK8+sifjLHMBJPoaJ2PQYqLDdgNdauaDa+SG
t8dmCHVh5HYFSbxDQn3FLdS+MfUcPfjAM7BEPd7XoxPm9L8fmEALU9LHf4wf+DUJEWcF4c3zKlMM
W2fML0hZwAERdWEcL4v0uZKWPfl+W4iG6yocBvVgsqtUKMBcoTH33/VrD2fCu3+O6arHGPTZCNW3
1ZTd3MgLK9OjhOIRMWkTZ+vc6Dioz3i1Rc1oDH4LGXKAC5MGOAAaRbNktJWnmd1ZSiuo5OurRW2h
cM/dT+h0/zR0l70l3q5TGdmqX77whQnvUCQkZTVaRj5I61o+4pwNQ58EjtBYqfWnpYnPBaiFCtSK
jHyt6ZpDMu4UFZUR54OolSyi8cMyLT+nBfIyYKyBDaED5Pro1Wol/k8Mpsnq/93sij+Hdz3dT9I4
fGzhiQGkjZNq6yBrK1TtS9+G4oHVDCHPOctSW+MvpNp6EOF+xgSC7tkI/Odjzq8rBid/f2MuEFpO
nQNjW/4A+KhSXTfsydnp4fOXIkODsg3O7L2GSm8Ql8ZSp0HmVZYPbUGlOAKea2YiqPubS+upKvTa
FsiOktvYfYTogjQ6b1vOSY6c7yX66vb5W349q6orZl2fAeTb2Y3uecLG3KLdnNZRlSxZxR9BcKE2
9foW0aNRz9r7rxCQcgvUtliekQLhRNcwHqyA+DQF7BhM3scsv7Jn5huxaPwRmRxDjsB0OMAu+ttN
Pc2ury8Raeb1YcSyqWE7GrtT+rntbBKhK4ANvsSJpGptUD6w0kl7O9UhiJgBNvrkzf4zcFpB5XUQ
wTgdOJ8r4Nd9xbYKwe6ojvchyEUKLHJgX/YtB6c77Dcz567Jg+4TcrXkLV35tXHmymB42SoUt7zY
XGJHOyq1JhYODCrMrSB3B0i+Xj78DkcZnu64n2uPl6gS0BdBkTUuYuBjHnkQnrtKWoxo4qbMAgy7
38UlHqEjXsc3l8/r11iBp92VhbvPSGxeTqv0dQSs5tSVKoMnIc6xJnzlXkNaYEaMlBGzSZ7WBGoQ
v7rIFIXDNLtSBvW5naw4Ny9jPJ1hOh9usM7it4kRL6gvyrU67ckrQT0IHkTOMZ2Zc5IPTOWfOCre
vw56Kf9nG20+FxIewtgpSzrl2OftcrXp12Mzur4VZCVmZWrJvv7Q4sQ0okIsTKrPm7wTZMIZxvAC
+OVQl8WqPl41OWPPuNBjaCG9lBa+1pqHR6SRlcGWavVd28m12HlpSm4B1nR+QvykdjgOAkqF7IKk
Ckuvyck9cfyvz6JrF0FA2ZMd8NT9eCn7rHirLahkbNQms5dLo40qh74WylPeW6GFBM5FuHWsQnql
bN1mLs7PEB+Wpj7HiQ0xVb6IKS8qefQrUNriJWtbRya/E3BLi8XlSXQKoAXuVf3V0b/btuwfMy7D
Tphny++exYlfH9s5TFs+/Ay6ZCrDpNNnDdevTpm8X+ijVzEEiTzV28X+FfxOq3q3afy5ehEhQR6E
6e5QB6IwvRM5/+dDW9VFgMxqvxw7j7gYFQvjTZjJpwNXNvXYOvNuCEodqo+Yp1KqvyFTxhvau/r/
ELNuLjWaPa9DGbh0bLOfvXXX+u8cDZyTCsUzob7hdkeV+s0m
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VIu16zY8oZeIb3QmOC3HosqA6ozaQOeXhAmUtiIJjg18DqsM+9kyGrUIuNcoACh+s7alejqVnGDx
mDk2ZWo5waZ7gJu3XRMnVFGydwpzKoP34+JEKpdWGmabIjwnQtJBmInWEm29EPlIBCs4NNomyGop
AEpmGJsXkos1T5imyDJ5AVDPHmLsydMzGaHEU3poZszaNYGkjJogVZDLUdww3LA8K9c5m/IHjO3A
ICz84P3EizB8HsPNs4/GXfGQq3ZLO4kk2hRy0eb+S1i1rzXW8j7V9XMHjmw3m+UhJoCc5gGez5Gt
BPfKMH3eDD17AcQ7lk5uvF4FlEi4uPpRZwGKsw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51088)
`protect data_block
pY3of/yn3nYIputGDNbkG2GlYoFweicQCpUc84ydbVt+F0Z5zSKQEgpme/Ju2Eq79IujRtCe69b2
nsQ8PEPI1KBMDQG/NLVoas0Qf7j1y+wR2C/qRTpOiPJNFBkZGKtJ1JnIVJncqf6vWVSWYz3a9L1P
nBwQ1qiD8sCz3gAnCYPoPOmTMCLd8e1l2SMNPVZ4eKulJ8C/t5ibOCZwiYAasigMhpbpurgHxPsv
NuBFwTnc8ljNOxS/D+1M7vMIqvUp+xuRk0iYTAqmYXUCJNoRS7sW5OCiF/pr3UEgKMFofxIx/6su
SsuPmqcwiC08453kkWveLe2CleDayHA6RKtWgrGXUrqOCbXwvPt0BM0stQxyfdD44+yf+x0xf2xs
ArUlYY8tFUbEMmZVg4FLfYK1kuW/Ixv57v4cXhwyDR1da+jFTqBT2iWXQ/G7GzsnrLgIjmP/O3LJ
q2ZXlTTTh+Xcs/hMEfO58/KUQzKohtpfQm7dbn+dol0xAtSQA9TuY1/1Cb6iAsm+qJsCflzYWvx3
GMUvJmG5Gx6yuTDnfZ5K3io3GzS8Qhiqb9cig7yqVH0YxXPlMwq2z3sGE2z+nnFvzZ4gdxIFi1nS
1KKwjjlkyY5KDtmNpDEwDsuP9O3AeyoRHxC1CTEC6n45xXVikd4OD04BiO+FfKhbeH9yheOKWFHn
/kQf8uTf4NsnNJDtaOUd4qjbJBcJINhGDptYZ+HPgw9ZeEQ4ERQynaz70ghHkf+DfoZuI095Bqet
cfa4d6AbyaX9ZJqMVMExBT65qk1D+Z4EQwuwDZiqvZGE1kptIFxTw2eiCMz61Ue80YrciBtNe3cb
ZslgE99SrIkXnoFKJfGQV1OzWVh3XpHiL0mLEFEeA/RHyz62urrhpfVOURo+7ot/LDiQ8VzWxEAs
Z4CTLBYHGuu4rB6XhuY/zJzFqWmaenygMAnI+AYKtkxE+wZAVWWDaz1m49IN/9FYkzY6fHG/Y3a/
40Wy5gBI7Mmzp6zYFgZ01lu8NIGnc5+R5eT59Uhy7gxI/pL+wc1eG7y4hrUGiYZThdFWxuCtoe0V
JY+kC7Sbbo8e1cBL3DYSG54RERXaQyih90omAkWN2pbXMnw9056CoTSfdW71S/9a9JZV3xsMgUpY
rPR5LfZZxb2+W64hqKqXmxkHgwbI9z9ljbpMcCFUMuxwqYvtlBcCvN/W+rFrSZbBOCQKuKI+eqlQ
Krmc0MZOVXx9jOdJAeB4EFP1XVkzELT6J6M/ht3nHie5n7hPzDCTbB6pvcaxv4WhSiUbK+jPdVor
TrteahJNJEIDhiAMWeBt9X1y7DzpZjoh/AVyVhrBPvRJeSD/KkhBOq0egyMq+9R7ilVw1Ic0j50t
Rhl3SDKjhkQ15e7N9VyI/rygjuHjF8Rx1yZQ55VGPAOecfnUoyQBVMtf7BSgciZS7RwzF0eXm3Yo
bzcG3ZCkXYHTP+08CXynBfZbAcoT31PLYRLvUg2JK74hbr07Xw0fl28Wn1Zz0erJ//vvxTJ2nufK
0LGkvAOYynjc9spP01sab5GOnE992AgVnlJq5EBpsS/RNGa1gVoCKpN1997Lkb95b8dtKsXf0MRY
hWmJIQ09uoZcljK7K/HbiiTV79/hCYcYrk+2LUI/LShR3MU3pLuxbh5IBALQvptY+ZIT1Cj1AFHc
6a9VVsed4hSpNJJCK3iwR7L9jF47WJhMEXkee8ivTN28xdV1CxSUOasZ31SzhODT5Nxn4H6NDbWp
IBgxPwuZB+biFEcUuArun68nb0QBlFZaB2JWoyA6k8KKUbusQY/cToITlHY5OX3GERTqngLXed+L
GntZulTRgzce/0KgZ3f9RPs6dABzCXHlbP60SppVpDBpNvUGS81T4P1Zk/69zJoCkJgxiYavYSIA
955kM9oWUhKUIczl2imVg0hxCcZCzWaIieI5LAPsB1UG6MxI6a6zadUO1BwekbqktM+oXzJcLQwa
cEHtWVopEVRmSZliAbt17SiiTWrTQyL37BYNSKbCpOc/pzKppn3mpMaRgOqSjUcZRueBYnbyk1Vb
fPaU5tsezuaT8h5fxNOwT/BP27mpkvsPysJxtxKT0r7uJ354E9UfVADcD6vOAQ281/zSe0HGAzN5
k3VNcBcVrP+HyLrAmh/i1tbYFipnjAQR0gOfmkuWm1wnTB838xEsjxpDbZApWBi8If+WNlLKLDGD
GyB4xzkL3OhwmcyyrVPXUtik7zIPzINl56vVvFPrQa6x2Qb1WhENitsC0Mb/0nhTy2hn5h1ucLF4
Ul2nyzt8d0BOlDa03Cs67kLN+VLtaUJbH5vKWB1PhXa+S1bT5TJNGU0m/UOi2c6qh6U60ulBdZw3
Js8niSVcj1m9/xSpFyjTiIF+0JmlJw+ic6W9h689mIZnx9nTxNE/Eg0P/J5zIEae/Ta7se1p/4wS
seJ2xQTdT1LZ7YZAwAcmNXHck1gfw3t5E3gx2Pqb6JUCyg0ZOzND/eMildA0y+wSMXg04FEXrRpi
04+9WkgpcP78DKh48RR4dLxrwgj+gIaObmH4kSS+AjxnyukqElgyMNiO11gy/8Qmqp/XNuQok7Hv
eTboDuYhw/6LTmFRSnE/J9MmQG+oFvYIs6ZotE2YD6Ev12ET9n2pmRjv93rpsKyf4UK8+VCHqI/u
LxMYAwjjuaZK3de1bOrOuTnJ8nYmkxgJYiSaqnjqipju2BWZ+FuvTZ6o89jcManzYr20r+XZjLjR
1EndqyPJ3BZcl28wVr5mOzzlr4bRAKm6r5c6JkhM9trf5ozMxb6dI/h91bTrEe9wCsSqxqeLTkfd
6w7ukvo5y0nbeNCIf59OfxJdajdRaVRJPY28oLyUhECc26fb//Qp01Taqmxu5Sd9n+feKsjtMSsb
XwqA5uXrZNcMzzwCPoa+H27n6WxNwCqnAmq8rAUO1MpwhoPzEBoZ87wo2iSRmqt4PLzb46+vwjOp
/MiI7WoWr1ZsT5bVDrK8C2ZsWVs9XA7fS7OeGeN505XZ2CMwAc0y4zy5J8L+0D1ChPOnSmRe2lnB
8GTyjkwbZL9D0OiRm8Yz4wDw+zZFChJ7SfZAYH2YFDeDW94HGtAGYRsrKN7gDMNhKIkAWhLW8KZ+
TxTGd4A0WNgI/emLD58+b9k3y35Bc+TrJOFhLw049dgFr5KBXKs7vYZWj9V+K7HAC/UKi9EcVSD7
b9zu4ayZY9d9ZUT8FqZyZ+ATlKyH4XFywrxzgMA040TmiD6r2+3mYm9R+bKUths8yPxfpqbrkXmp
QqOTch9Vp2VfgL2gl24/Qh+1PDiu8iNKg3SE3u5VLFO9Dnnq3Mn4lxgs8XMtPCBdI4sL/zbpxQy4
llM5G/JBjlf2Vxqvxmf4Nsiw/d/vHqp6+skn8TYv+svzbx4WEnpctDoscvaENmoSLuhPDKeEIWQI
1kK7FpI4qYHrDbm+Xfhty65SZ4YsZMFUuUwZ68elXCfResrplDH+fq6Pf+FNc8soR3Am2E6+G45I
HGDS00BZIuIZaeHls4IOiDlehaa9R2voNv6WYziXVF8u6DurGE0VqZYoOBv9gzttRh4a4xaBPSYq
xs/QpWCqTdBIK9NGton/a1zJ71BFF3bqNCSL1MdyzLzEp5r3re3IpXLU4CWLUV307ZNbcdWR2PYG
GB353j51BsIllAKQ5elFEWDzJV3brFT0Y/4v//+dmS5PhInlNkQ6no8dtzw0THJ+cXY8f15uXXHH
HDxwntbsWaVHp5CFhgYZ31lBVH2wHfs4h9ZoLECrXlGS8A/cEj9SiXCFKQpHlQ9IKVVS7g/morjh
2szIonj6hA/RFbmsKg4yUGkbYZSnNLP9Dz1t8VVU9g0ijhRqfKzzXp3FyJ/LrNxd2k/GB8yKRiZq
c15cpeH5tqLIbwaK96i/bfWIamkfE/NIz+7+S216Pp3Nyf5Wq8gpx3NW0iDfyi9RWI5L0GOWOYIR
/qvhJo79HYwn37hgMccnTHN+EAjd7HBo94ECwmVdNKZaB2f0rxuib5FBFZP0t+T4nkWb8dXCF7KT
PssS46wmLPckdjlfmrcSEEVdv+WnEQz+O78JkKZ+yb8zchpP5kK/JAslCZZR7idEHeN7x2h/4zRm
/lxb1QafOoNnUeF557Jyc1vjdO+P5MY48WXY43XJDYETT8WaberbSzWCvKwRjsdGZ2f5ZMDphSol
NvuqwtBgIqCls+2OCxImEDMu0Aq7qSdspWAgUQYw8LjlvhDJ8MmODMbM20zCAZ6da6/VgGj57qpM
Xck4dfMAY29HjvIgW0OWCiGEvMndQ9ljBYwrtW+7TZz0d9BYdSQliBykyPFulYzxlyp7VJFivwRP
TWxy6Md3csOboBX50jYIzTmad49uCTSKwVdNswuYNxzj3ZBVWuJF44jA0hJ5wO24PSRpeIkjiFrA
SLGmYTBk4396bHO9yG2lBcEbu1AI43hpGSl5WuJc89PbYb/mxrgmKXspb80fUC1u2ENzzSZSUhNV
lxpZahd+HLhCdiSfsZrYLpjoHpNT4l5vR+ykLK5h/SCNbnZiFg/HvYJkkCFvBIBArZW74XdYfEaF
2bWtAKXLvfXXD8WwvWwu0o1xPpKG0OIN9HaujSe82q9TI7F6g0HEr74INVe0rbROn4TehJCP1/oX
lC7jkQ+yBcrtjASRdvYifiiNTjGTURaLMYY4B0bkKnGPSiFWiT+ndM6XDCa1iYF/vKXZsXyqsi4p
Ql6kpHzKTIQp4Je5nVujaoAi9SLsfMLbTHyC8a0rY85fk8AC6TuI4G+Y/CJgk/jmQxG/Tkxof9/T
m8WT1z27SRcbSwq0B1xkcWySApt2dcUvbX9G+O7m1erCRDAndWkITN5g/q0LULDMfvAlp5v5B3+N
MkWiz4B6t70vvtIqiwm26mgtzXi2xAU0XSef1013HJ8mnZOyQwEYawHfd0obTZwEnOPpJ8PzGnR2
2IzvE+JHF7b8a2n9YpEOqo2g11xbYBWVL1jBrr3XywYQRgEgAtADA0OiqikcLzupeEhY1EtUyYU4
OBl8XLuxQ6zY0Poc55xbJ48kqjqxM50gI/2XdSjd7ZLJGzqVVoWjzSmJsVdsB9TTSDU1+xMP8etV
lP2K9sluQ2Vh1W8tyX3QrwJl4rF22Ff8jHeowQJ6qOhpVWQK29Oys3tRGpMTiCTsyh7e3kAh/2Mf
zAhnpvmsy9j0KqjanCUzIfQOoVrg+tTAHiVmeCKwsZI0OmCtAIxEJhPCYLzbUKmJJbD6vrO7UPwQ
W0Pt7C4RGWGbU5dZnnYZ5zozC3fBsaGcrENNLbIa4CZPW3ykrPrNACJP5CUE3j9KJsOrUvIhM3eH
db5CIiqwITJrXuh3rsvglG93ojthMsjtIDnm2JgrdueeYacp9ryB6FnHC3qs3WggcjNiz4QrPy67
qOeTiSzpd++OE82XjipIHnlPF7ah+mRQCyZlV5aoqn/WSp9y2g+RqR/FCSC/sCejN35HUxOUMv0c
R55d1KM5Ri1jQYWxlEFUpad85zIvYhg02H8ZJSQuzG8BitQseVGM6sS/IGa1XBorN4SZoW4j42S8
DnRDAJ43Z/N3QEiPoMEBVCfOl8yKNsw7xmmKNrBbr9JKANV+j5WSh1axs3fTXNy4VE8qoa7sCFXq
sdyNw9WPo3zGBDdfb6Pz0T6RFh1pzaMBnTsuyE7fKbIKmiFQE0wR9fReW7Bz4K3dylrOJOSUpJ82
sC83MieFoqds089NTkS33BnIpDW7BmBHU9FVb4D9p4BFUhsqOMTODiTuGLOMl4nVWty5eZcdXmPM
NE05k7vfuwiRxj29OPtWjD4XWY2qRleDnlVXOcBO+4H0B3f3rEfa3DWUpDXDwXZAM5HGiKC1FEz1
twsiSMTWG2C8gmI3Y66lR1imh1yMXG07Mx0P5hJUfSdm3PINtoVc8Dnxw3oB7OTG8CxWZY9AgpUG
F7ia0XxbHilCxC8aIDlMsuDQK6l6fe1a2zaRFhL8h4VCho82TTNhhFDGjgtewKtmXbqCBp5UUeXR
Ps5njU3iearPvrr6TPRLjFqQJOQ+sJ0Tpus6me2m8UYFt8xPeqs/50mK4UNyNANmfVcGTENZ1WwQ
R5lmZCVdR36e8sWhVudCXoonBfZBBKOmdDorQlRVoAa36Cyrzd7dSdLkqOw+55fwm+4FvOuUhxq/
YtjCsr6HIL+6GyyBU7fZsZd1yPGXjKSn2TlSWfg1+7W+oSrETCgCIdWk4z8vZWnCX05p4T3PBLws
HiFELzB5QUBBOZkFZfw4Uv2/RCOyqK8oxgIo3egsVo0LeojD0nD5DMbZUmQQSVYWFJDaKibxmdDN
Ti/gCO2+Snwn6pFxJ31aKZT5n9QCi2dzY6FP25RK6VoOTnaoKvEQ+aennFw+hDRzkeQhMgccAvV+
dJ0CNncJf98oJox7i0fBrLt9WwW8GNLQ4kRvtmAbk3BIMitccS5JZxT6FYCXxvYIKR/gP2NkLqVZ
b6ir+63eVdJ8SVZZewg/TCjoZaUgFEiPlTJ9U9cyWMLmVHYbODitftQgxz+zwjdt2wgfhIGbHtCA
MDOj9eTSJ29pf2kLRjXzQ2cMK3/pi2QXO3LESfOvu+RYxgcTZUR9+TT2S4Y0pl5HykX0mCoG+AWX
plKXr9Zg+BWE/qs0RUxuo8eb7og4UmQ6fd9dwkCNJSSmnhKKxWzzWvPvGw7K0sZsjzkQbbI1FgBG
Vf7P1g7AS2O314qSialkJU1EwXs1KWqjmmGaBJ9OFNIEoQVtsK++7JivVhe2i1YYu50CJMgNwdBS
8pA2T/CiU7cDHS0meLsa7reSC9DjPgveGX+jErJRutdRYJs4BbEB8WEh6ni21v6gQAiQtrDVB2yQ
nWgNC4/9bumDMKfC4xsWQJGUOZOZvLCsW2SLxdvQLlhcsnEYTKQwz+n7pAtDjc1R8K53VzUP/H7l
rYr+rfAvzvcPXV5+ycP3FzM5CB2WPN/DzsEk2ms3NDoZYpkuylRKYi9JVk4nCoGCf59JcaHCzkkN
hPti6jszTg/3bXbHSrYTUgYCeLi0q/EqSEoV7s3THChM6iG3UOFm9o2W+02XcN2gjq3AkgdjUwzO
s+JaZa3+C7uBqRfOXmWbDoT9V08INt0LGTy/Js1nzWm1jfDCfy9qFPds9KTcDMbCHNSvYkboKMfD
8yXQBix9wIXZ+2VhTVarFXRH9bd8rsgIgvZr/a/5vEwWGj5ZGTDJSJHwo0ztdnb4t54r8m9YMXAC
hVA761K/tTndyReqHMAdl3XQVKxkbwFfqOUy+h1OuNLebcJIHZG91dHnkmAUzMuNs9beeZ0eGT04
xRnvw9y2/AQumohcRnMH2KEgC8nek8avdp4iZjRI84POY/anvv4FamD2NSVQpr7LjklTRBd3E8wk
jblLUa9QUdkciZWUTTEN2DGw+26j9e0kzF7Fknovn1xSDUbnlyD1XOWgjdbGHkWH/NLaBK5BJCtP
uiYrMnvqpXkIg5F5WL0BDJ/qUX02N1DDY7jNdyiw5uwNsD08IugOORoTJiSpt3gFV1v3QZbmzhbX
yCfdyVXix87XnGR9STNL9DYDakNcS1HHR0rklgkXUByuyt4C4g0aGivHod9/YEgy42CBP1uzbjWi
m2A+yWSwy4QMTO2TeNU+7Flibo8qdrSSuj571nbwMg2c+zT3PYhlMiA2Z8IrXhQN3iQyr9m+XXMb
7FmDOefMW57ITEmsHXgYTJ9mgeilK52ZzjCYI5BRx6GJzgq9PUrNPMooKvxHIln2gpV27MOGWAvk
KSLZeeE0Wzx0tRlmBMGM9PCUepwXQ5MCOx0pi+ORxGhO7Lxc9NGltXhTK10pCmv5w/zE+/c0rpBX
nVgHH+VT8vofM50f15PikfixuRhRebUtVqyJnBZc8HPPgYmWiXkayzVryAGbWasMqVPBQJdudknL
zf3mlQ3GxnxWvRHys97EAB6JKIE1l21twNHLqpriRSpLuieMxICLL7rWBxnP8KpbcC7aCoZEN3DZ
dW/76ZHjsGbsE0DXYehBISHM8saEhjFCgcS1hM9fmabTj2LDgsS95C+OEkiwUVUX0Q3PCUSg1D9v
oJt3SV/gWWzU0XHB9Zrj9w9uMXs2RUkv4iYhAs0pk36TEhRelOQ6xlAl58G66U45Acw8DebabNYR
VZ894VOi2ZstGS4+/KKmIXv9Kw0OtivRr2OPSvYnmOXdaQjG2UGlnU67Qzm/ayv99bDhvYpRX2/E
PTHyaLGo401J66mKj2AK68H0891eK5M/bhrKghahhJGK0xOvD2JsO+udh0CRPZ2ZTcriMrnNtdTV
/PbJ/071DHSYFuqoXR2alES17kFcjQKDVVFV9Vqf30091iRIxyqK0qU+pQIlFgpIQahaM8jcWYtc
QhKiSSNLbo+60TOox1SOHSvIQWFpi8eDLj5fLaaw6cWFoAObLLvnNTjuUkBCDlRzZc4L1tcuuTRZ
3Z8srUUPJeVH0xsOfnYpe4cF8Dk0rFd6UdjQD6JEGZkVcradwaCJQo40XHnygu0OBLLmEeM8M2W8
vJkehc1JWq9I+ufNv3HHQLt6OudMAsgtyOKk2uHsGy7zI3QsOqRwohzGalHmDYhcpcG8WE1EiB2a
+e+zEi7/PxQ9X/CoOH/jT+bpNYBOQvFDf6WwuKbwrD6BTumeFma+Nc7cx0OWxqqE4W4Lz2fl+uji
KC7AfViSPG49Sk8SHj3lAsmZnf45iYlLZvQ99B5iegBVNHBH6kdfViQsz9Tqa5cmsayn3KKLfgyT
Gqx9saIQc/iu/OofKMmn0tC5PKXTvkLflR42ZM3ia14dMHCDEBzFqIQ2lAywDgyL/wsKiXKWyDJ9
c31QZ8fpqlJ0J6OzmU7bol+nf1YNSxKp+nDIrE95U6Zex4rvMbX6wYtW+rEm6D2aLb/TnstWU1F4
17zWD83Cg/bGEENqKaA/MlG0KNoqEpJzdyOBNUYTY97wI2OTg8l5boo04b0QwJshAfRwcQx3dV2N
rwqkZsKyaDiJXP4hlqW7GmskQmhvPgbgwlz3g+XSB8BV4nKhEMbZxMegEBDS5KMBkB8TTZ4yJnsR
KOcdBwaCGg+WO3utfyFC8SLhlSwLHfV5nOrhJgWQybrPHW4CgEceymiuGIWRKg4kruhtp3+QLizs
07G5Jr+eK1iMZP2Od+m+2gUg1dZJ4btJRYNNTnh1n5WjrM9x6KCBtPdUG1CLG+aEBFV8ooC2wDwg
hoXUr4MBZWzlkVm8B5ijJgDCA/MY8KkxxmG6OmQk//YO4qHe/edF7KAG3OWNW4pLZISaXx7c2Tqd
4NzTd0e1ej48tL5Jhn3fdXl5TBpGYe8d19jy2poymak69nVg0eay9oWGPZ9vxppCJa2A3ZlWstcW
NZEmPoqC7YSoB+ftOrdMzgsvHtDgLp1pe5LHF7Hb9/hYY0523plNeaQeFCsUqi6pkDGMk1m1/43t
6vTCoyY6lRYoneevb5N0LDohWfmqxx55EWdOIEDvPAnM036IQPzGGhqm/EVGYiv2R+3n3l6D+Hyl
9rQSx1bBasuL/fmQmgzoJaaL99ut5Gu3QYN2Rcxhx2d+33iT9Ligf3H9vhZIzMHPmH0CWUe2UWqP
yB5fGXP0yzBZC7WHDyraiu96Yc6erk2JIajnuLq7qyrcIzUrDhBiyWbMCoXNFtjr1Ia4pkV//4wp
VN9UP3Zi81e0Ac8/XtREAQUh23HV71uZmzXHQrt+SKoueagNiRojcQT5Vl/LaVKgADBnMr42f8P4
zYwlO+E26qKh1hZdIA+3r7tbMCCOEFsuYEjDsGTYoNCuSfTHeTKbz41jrhMMzm8kjIwZRT4bih8w
qi6XVOVeGw3/mtYLAc/fn3TOQf4apfPbKI8Nj+gGOEHhkv6//Fnf6/c/I74pC1UeVs5CKqv+eULa
6VjXlwELKs/oaioHh/fqdN6oTfiIpvMgM9+1zvlLymg1N9jnhac4NE67DV0Ql3f2jpKvKAxJxvL4
i4Z9RV2FP7hzx26dmWnpYjDb45QLsWNhoaZOG304tpjMHseo5YewKwvmVj0+RoNQ529mVygsm8vy
82kDnMS2c0j9I4+DzVFzBDOMB51DhMs+Rf773Oj/bbJ9sTXwOaoIeWxfC2VgWXQpshM/QmVfiMqQ
oaxY+VHUQcDMfDLq5KECw9hWuXsnnF9Cj6U+N/dQEToS1Wuyi9unXLilpmp4Xq3sssUegMOZa9wS
E9l+B85KKUr6oLn4xvD3R05eLI88f3bzkF4iBMaSrLzSRoEFl2wLFoQrSMxtBfHNxBYeGkZR3YGA
A5pM+SA41YV8qWBHsqefBIyIrLvVZkuDCsAKWdKAWzeXBfpNXlkI7IBT5CpnQ5xZWg1LxJR3VDTK
gQkVklweMpYFVFFrgnSMjWo+tN2ieNth83Pbb4gJtHlv26G9M6SRMZKpzT1rGmFY5YoRf10WDe0Q
FrNDX6/2iANjf4oYsDgyRJyj75mtI+RiuAnbfaYU9aHvELpaPWiSLbxM0Mx6J24wm3qNnhFb6WSN
OMkZfuyxFpETtPE71vd7VblCQ0kzGkJFG5tPqnRdLql7MptsPUyWSUoVbID/BsyWsmFKDXXqhyT1
TE60M+yBtHxpOnajfdrSX1PDD5vkqEMV6MuWu/suNFCNGIQDZxYqzHDDT/y90C3ZUga/q1aATO8x
hjtIgNTCX27m6KxFcFCCCv6JpxOtVSt3T93aQkfHYy/d8CUROR85N1t971RDcpkMcPPLp6trrYh+
pfturhOd/6MMS0QS8IlOOkSjUKQnrdahV3VqGviqXG2X8qMZSJm79mC8La3u23xumUglaW/K9H2c
hGLZnb9Rg9g+a18tLPxn8V813gKsm5Pay2rvDUT4nANvop61NfloQvP12ccbmub/l1d/4zkmGJtA
St+DhG5H+Wn60asxjtyq6pDc5XifBX/+JKSR3MjSNZlWBHUvju/nqVw9LfsKISwWuWdMroakM0Jn
yCpDXjxZr13swsdjd7LvDkhJURv4i7RkxK5i6R8YrhmWzj5RkTWZAsUvc3K6/O7pDf2gxNpbbuGz
5JtLju3dpMlxqo4yydtFbE072NPIWzor3YrSZYw4uvzZT27JqSbKLFFlfZFEOqm5zYk0d3ZqCvC9
UAKGt+hepEiB4u1iJdOToWcMVlj4eGQNynL5tJlCVUBtFypAGbZjvf5T5bWF5Lb/uo0OQwQ6UXyu
G1BgFQF0Vv9CYJ8A7uvbJnccdJ/YDb2/GyFVxVHqtE664CHD7Zhf70UccvV3kssp8lCkfI+dbRg4
BydloJ8Lv/x59FcZUzELErA8DvrfRyc3gC73tK92DmcIJNgLMsOafLjm//9VUWgFrp0uIkznxvpm
zxgdSc9wEwloCgT0la877FEA+MdFlkJNIxoz2PwRdFKgDs/ze395gYncJZbHSv6VD0P0nKejQ/g3
9NEq+NdJ6cgqH1SiHoECZqhdHYh3pQVBjOShuZMkqxWcvaHArpxLuVukn9IprdljJIAZdQJvbJNW
zVwcXixUGZ+3x2L5FJ756pd+mfDKTBfZbrTxEVccFoE6UNPxs/KtoMNReW0AUSWUW0a5MLKFkG44
H9C2aRdxlMIo85pEy83bcLr/lrDCEKjBtMvb5FbNFinXlsfiKOgfMu5+IjgApiFuf0nemmv26BNi
nUWDfno10Be2qtnaVO4g7pltKjAHMp2pkeHWnSEgfN1i65Xk2F6psGbCdCND6mbveXgN/ut1wwXq
5Mfcy2fMwD7r4Q6WsQq72gYL8YINqZNFcUnx0gXZg9ckAT9r/xZ+OyPFIj9puv41d+rAH79sfax+
HbfIsu5E2+Y5AMzL+Jrlajk3YiaTV2guxswqAJezhyhDVkb2FC7gLVGWxe+GINAkPeHIdFr9+BOy
yo11seYXeIPDKkXgdQajRomGLKQy5weOOZ7z6W+u8SIE0l3UYFSfUFoA3sQQ0HV6FGEZwR8uuL40
8ufAy9OyRpu0CwX7mCIafT0iVNVp6HWdYK6Fdni9hEDOSApmw/2OJ9GaASul+qx0Dwzb/RvW+28f
FjKLaWNDO3BnP8V9+NYgl7LE5EWbhMrD9KzmZ81GZyZONJgQnkSLIyatklbKG2QL722cgxPXLLoJ
tyS4lTbeS9c7vDAySOJW1QfdC45Hm3lxctcrrTLzQihpIGjsCf/ZbET8L4WNYmI5E6lwl9hjDBOt
w6BWyiWkSTs+eYpZmb/sf+32rAoo330l1KzjOjo2lKcNQ0ZlibtrVuJ50j/EpLJ1IpUL6hMQtGUD
JUaOPv0S/s7q6wJCS3yOYGD8HJA4LaFmh41UuFkRJGxVOnA/ou4G7EmCcDbJZkpe/q/t0DopeaLZ
i0DHFitd/ammMTMmYSf+u+Arwa9ck7c8egrnEG7qPGHVP0lbmBc/iJ+rP4/PTdYqX3LtdFmdrnKk
iRbxsXxMt4NY2yfgh51aQoChPCOH5c6VE1eiMBiWdJbgJgm++qA/RR0Oy6QDoGcfKlVpFDv0FPjz
djrEkQPXTuuMvytXwiE27E8fLEIsYnbcRWSjc2qKbrBboX1GZvi+rAO11Qy4F6OklhmSVDl3aLv2
H3L81egA6k4AZPa3cBAosCtWClvIe6TDtP7D2msvTZdPsmTOl+DQtikTz0/dJs9ElUsJDHhyXa/a
EPmhG1U3L6h3wQ+SCXOsAo7pTzIy/4xgUSveE9ALA0ebPE2PJIhYcjCeHpvt0ZiivgUdWu4Sk/Ry
Qv2Us0x8PMnhNnqmhdMWvrOBKvEOsACM97sG7e2D7Psp6PXYG6EQ4HxWTRZTmRKohopL6kpahWmU
uwYCdAC3tHGZMVCkjgvpDt/zrvoVkY1vDZ3AmuUXkXztLXDSVmGkkAaGFmd5GqRfOfrBi9Wn4qVh
pstiGYZk9+u41Qdl6kJCOm2WeZD+v+/3sN3yXPAcrKyYm369gsLt0BskixL/y57u1aghbIPCd3Dc
TD6bVCCCYr8QrKVY2Q44xfljdl4R3NxNq1yS8U7wqUpWrFFmlhAG+Nn7ZEtTSdDtKrrzh3Qx0Bq9
/sk9SdjG3GAf5cUurFK8tDcsw0BISNFPIfX8ns2ZgHVnArEr2cnpg/ldGunfPmu5oKZ+dclfgMZ1
IRlZbA3ZeoK+HySXaKPijWFmUuhqs3k9HWhQxhmkrarMpufuTggqfAQVuVXfmbdstyCKNFsk7p3j
i28DzZCYev8Tg+ivtlAYdjtCuyCv2tBGXrmy9xtiyVD5Fc+Megk0IkowTEjHSotMgX2jDCgo8+t5
fke/IsL6cmDfMxL1Ug6M/bKlbg6QUir4EZiAc7sn8+r3cbtYEBcjfeArP4srhMWhStYM15s8yFbZ
aGN66zVGFingPIIYhBlIJJ1B9pSaK9C2gBHy9Do+SW0/2tnOaljD7Bu7zyj1Gjv8d9duQFg48sW4
eLkjSslmwQXepxtSWoSxIEit0qBrgLsMtgzyeppTOTCtU4hy31JyDIIf+tiSuH5m2LIv4s8ba8GZ
TWw0KKJLjZxNTWSn2HO7batQPvZcTOagUVqw8kkmO8wJ697gxzV7LPgXmhAM+EomEpTq2n7+p3mg
/S3z0oPTyepd1ntmegAZB31L3T/D43bmD5Pm7GSoW46PjStnSHTIzhPvxybHXigJdB/MmBb1kIrH
XDZ3lR3ZSs/dbwh7kVqujH09rdFxcwDM1cBCM2V/HXsExxA4FDy/wmofboluxyF8f+ybuLDktxVJ
UGnaiYXTefx2F/wEC/eo9UsbzShItEHxNxmbR7zZ203HmF53s8ylAZDAQzs9Wn55OFJpZ53cE+jz
Hj9g5YrbzKAA2Dog8jEE17DSN+oRc7eMMyUp736a+rwVj84gRCVYTCp/P6w7ceWY84WCoJ0h0y1P
JV9Hf7cdtigeGMFP/v5PrUCRgGnvcxqZOYMB579/O2D0eyvfKPnsZeHzV3uek6Ud+e0ytvEUJZ3A
naQbibaBHNb4YFxdUV3vDZJ+oElszLIhTJ6tupBhMVDkvUUPG/IZeDUxzw/WMsDcRRXyO9GShtQT
mASJxfipv3/rLa7/q1luKKsg65487dnv1XIszR1tg7u2T8o/9s4819WkDSF/HUchhil6FfqxLtUq
5RT3n3CGZmZAEz3PyMiWTk1kfx68iccJh4vz6YPv8pdOQ2noqpE8whtKyDYwt+mZHkoN+dtpswpV
DsAU1CGj6hPoBLrmpYNwnckgvoezIolpfKHjCqY2jzhPEymhbTFPH0TNhcIhq8JZphcsmL7ljOxz
3H3NPDfwqcKyRXM5KfArhq8BoBN9zj5clvyWduo+xTOs8hgdnMLRuMV6BduGjaDDQBCfZbl4ije6
3QDpzo8WtkKmT8oTuI3neMTU94rG6ZDg5R1I7kdbcrCn9TG9N1csArImeXdgP9hybJYPgwuVhO6G
yagSBNh7kvuLP2r1Xi6UzIN/UsQ38UoaP1Fcx7HmhhvdLoOfe4DGJj82GDSqscqSUyA1/gi7tBOv
6IPQwia0yoUgvnaOKGM0b9iL/0o8mmz7m+oBp3QGKtnaCeqAme6KllLi8+vGpeFDmbFhka2gFm9N
99ZjbgRsk22Jjo+OpZI2aroYe/vyXRC135gyNk+K8A7P4R/7uOn26zSlfS81U1LDS/rnUdpnQPR3
waNmuDsUzKMTk9SpFMoWvpM2G+h2o1K6TTSXg+5b4rmjiCVDrDdM+P1upZLElGzzZgY6dRoT7eI3
Rn2LAjWaTT1Z00TABNYT2dDi7xlpPZA3DnNiHyzbgk4czBbmd1aI1Wqzhtl/dxgEpVMDwt9WBIPz
rCxfF4hZPCLIHWhzybFmJJ4zQFCOUNsjV3dxgqQy8NKHHmv+kCaLEbEY6UBHKzfI474Cf3sofUjg
pLSZsG5kS1RD4SR8ICV7wLbTWep0TdyCAw9PrBBAziYP+kb8m2FbweCFWxvdCqi/La7DG2rywS51
EN6oJNrW3OTrNnPJ6vJnI1NfKTT2r9Y+rXgEtnN+31RKX9TP++gx4kHYNT2InrlzG7GE4blOtg07
0MqXMngMVfXQ+SgJ5hhoojgC5POSj5sPUuAMv+e5ZsMlNzzT5UvOV8FA9tUZglk9EN68PYK9Yko0
98cHRqgoU9uBb5mqWj4P9DxQAMj8eXcrKPIBOe/4q76oytr69h5P4w61/kOobERo1eWBsgxDfi13
aahcSbpZkpt29W+1Ym9JEbbJUgMvzBiN1yMUuN+kqCEzDVtgeyuVdMAhqFpXfbw+hLOZ5NrVLi30
wcpkV/6dMCEf1VsmY71B8Q02Su8rjGph4IQ8cjHZaGgsH6A6gd90Pyifa80CGyONLOW43hTAgFfe
PgPFKVNdROuGALjjzxXUTAi8eL7jmH7pj3Wok1bsWQs+1faU0iV391rReIF0npTXYiwkSmZmdakf
ZPQbb/kYecGkiiaYkpcZtmyF+iV6TWI0yfYFJMZWJEBCZ1sL0eMPYJVuiAT23r9APwsc+o+HK4Et
joYy0vERMHAS8hQFHYxxrOU5d2zSYTq7ycFuAoyhQ/IE+U9CmoDBKHcvIO69d+FqitfWXtwoKox0
TT/zW5bDEsmvocjwHrcDx6uv4BH3FReb1C1H2YR3oKuub3HktKde3SdlnDFXnKGqMdypuKnCsorZ
jahHbWOgMrycczBMbpGOdfA0nGmOUXr+9sUQGVMuIYWLLxdnGPG4ss2yHFdJefOf3Qom9UmThf9Y
udnZAMKYwyGoVnxtvOYNHD/yGmNsfpNqosrgPRRfVeOms4aOKKZjrumltWMHd7lRt/k0yycQPjL6
d0mF8ER99tMy/iKHwkTpEsv0x+9Tqh/pKDFOYZ7tT1CUGy6lkNWayLydHsm0s+3UIf01wnjSVegN
g8m7ofOBXf04O2lpA/zlFyzNET9sNiMFxO1a0XEKzwb5AB6IX7DB/8fllROF0XLKCuqB8X4QRm1o
zPiPyKiTwWt9OaAq3aoG6YuYFURpKjlswd2hK7A3nIuwGMnK+l7hdydZCGeEHHEWxrhjrm2Jwolj
DAzdDsb/nMSqPnf9hTT2vo9U8nmtWTSmhnR2VSbjWsgL9P3rHgI/+rtIFfdpcYOQOPr3KbircXQX
jRb3Dl+9rblUCvHV9kQx36uR6TAiK+y/jqCJVlINgGOAz7VrcEMYEpwd7km+ULa6FeGhsP8f1G51
vWVgQUFKa/UBsA9aGChpSFg/AJsfrXDg96SFY8DERC3LukSLLW1uwP6FwFogI2XpZnKcH7jpQTcy
ZeEvRF0b7CqpKoYZtbmq3kMnNpU6eoz7L3Q4Hi/QJvVTcCOv98uD1UgN01YwRd24TDsXBCNLeSWj
kuA6n4aN0ZqwH2+WtR7ho0jrd+bAMSPJ6n2bF6QmkpgPlNlPWhf4Mv6aaxW8CvvcV5fCoSxqjmlx
ACUaN6q63iCOCqjrN3DtJS+9CTdpBoQEsYRn1897hFr3Ebgv6dq4J213WdxetaiIqIdnPH6nxYXE
X3vrqDCa5KGbENe8xUt4wdsSjrxhOPNz4SUxIeW9XTYBX/T0VRsLdX0gurizZuLbMvwfwv4cDZSV
7PAPkCJ2EI7T1GAW8W6Z18RBjB/A5xbN9Np19SUs59r1YTvJSh3T1ahl3n2fpqftjPWzbhocZjOb
gSxkSsLACLONXiarw88PLX3klnVWcuNONcEaD1x7CGN6CNUToJRyfaotVmG/jWfzbROjrI86UR2J
I5AhF0iPUppr1kweeNHvpVgzOboJSYsYmoKlSBGQdPEQrWxb+Pzd1qiBjjsDn+LWYyNKjOqe+/IU
Jz4vS+2WpmC1FqtPwRN+82KGIYbTY2QRanpAH+X2mVuuJenlPqC1+BuBVp5G7bn1XNFoeIRepWqi
sRYWWaKVBR1VkcAoa6bx1qiXhcpAQtbqb+3GoqIlhyW2d86moDg5RsalxEi9V4KHTU2urhRb0fSQ
l2t/D+5HILlrGErruUNfdqIC1BcwFo0aCx8I9c0MBsyvxN8VVcIOaQLPlW9r/+BAJzdS6k0zBopW
P66Y2IARozz/yCJwQLIFtk2bBaNZtkhEECeeN6ljQI4VBeXfLBfgHNcbgV1CvC2ivyuM5Mkd7ae1
a2lOVUaHHPWCk/hTnabMwQHMgZpoabB7KLW1tVPV/5xNvdXEMmCOq2R5ZdkKeUeVI89XMV6ze+f7
L9D7HP/4+ADcT5pCJP3AKVDU2PAeNjUaBCea2ZmaVz2HrAALj424qBAMW31KsRUCLPiTDkBQ72e8
FXBuau5s1HdLHTnxwY4ax8T6Iw+/Cn6LDIySHx6hkm97HymgufIeoG9erm5R64fVQ+DOLHgNDPb0
+SqsRF/cJHnz8Q6mMV+aCJxmLuoRR9czNouo5JXAY36lUkvIjIj2/Z13kyo6WOz6EydEeBpioD6A
dFbwbpvH2r6b+hTLbpStSt9KFS+efQUZerF4wJC2rB73u09hjJO4jTMDbXhVZruHCFM4630/QjAH
BtQPXfzn6+8oQmF7gpyiiy1EnZFgvb1kekZOx55HqO+20c0tIFyh3Khql0IAQAvFPZ6agp/KxX5M
B5mVzCiFsJ+g5Hf5cf8VJ1OMLH61nD+0ZTBqKazfx+Xxi3A3nwlxf2pvxYhacFUdijws1JFypDqY
Etauo7mRK4hSsZwPf7ilIhe91+jrhskDo5mhK9946d4ZGNvtygRBaFMQiU97RX71KnZQYm6E2ZKl
r/pJlBFJBVKajFcqcJSdu5JE7KdMjUY/2ACjtEYkcoERmhuY4W1E/FnnDw7NukpGo546XOS6bnJz
kp8wwXnSEaMmUKVg/QwWKZ6I3arPKS0DzEHh+OaDc+9KJsxuuspLi913Bk8udx6Txz9GKv1U9dbD
02JvF4EcDEkxuJvqw8b7xq8XdXsWztuV6zuxR/fePLS655KS0UPcSayPD4L2HuRdp8B0Hsle9RDF
wM64Z7COfATWGJisdWBOYukIcqVfTCtlxQWZTbY8Bae35zoMPzu69f4TGEA3pC4xmLuUfDtjdUiy
JH4PUywVnH328gQ2e+QYZDr2XKrHMXz9Od+S813IQS4oQG2CnkIHuYDq8c5berEoVBm72YocJvig
BCRc34LuBjkZEmz65XvPskm9kHwUfyj8qhxYv2mgsvz5G96vCcYN3ojKf8yq8Jdnj8ylFV6ZxB11
V94Xm/tGoP5rSpn4s0KFLvEY1NGimzCLlDKe8EscuDm9JbGvhctTW9e4cKcUY/5qwyzS6LlNi3fG
p7U83NRqcuS10rt4cjoEYmTusgwxiw7yKrcPFhX0fc7dAsUH2M8tqAby7pbEuY7Ch14Vj4BohsCV
b7UGBIWw2YJ+6V28d+Q1wWLpL+54RIiBp3W938YR1BJGVhxAcR4qGgxzdawv6vqSSUTqwM5/D5l7
K3mEvz3hXdIIeHTXIoefwv5sw2BXcNIrwvNUt/ajoz9cYp1jsNVinjAmT4/sdthuMC0MDz/+GZkT
lzFIfmzAoSYTgnHPzM+P4ZcLIwHWHcjKsP4XDIgwmUzkyBRH9G2l+TQI/QdUUNasUAUEnbzqEtn2
Iqbb2OK0oyZIEs5ziDXuR/B6ThD/pZ40payUse/1GPkIjx5c54zFc4uaTCmyotvgwAxpCnxHxPjq
e6X8RqItiG89g4vlC6ASp0rxSAN/q0Tv1GMdWvVWxJX6joYr35ekUh0dZnjrRNalmyeNnwt1y7Hv
PME39cqaCw3Iur0x2CanG5OHYI5jQlIh4avj6/NBG17Xxf0+EqADNJjYsWPeDggXbjSMZJomlSRv
CWxU/vPqnyyCx9doa7Ua3xEklOPaoNA5siAFkF0nZdvQxvtIychGoJoAVDtfyj9NMgU+bDjNcFK1
SQMZGDeivOf6n1qScFGNQl4g2pgZMAEkMN+2y+6g7eKGgt5u3VR4HkrTxAJ4p662KwvQ+CLTXjGx
2+avOaBj5Ab4jM5wnlkyjXDkQdtNCA8Gw5BLzcHMou/7AdLTAWFij/aa7RwN6Ka1xscvo+Np7X96
rDKDhaJdoHz8kq2laIUN2nEa0SS23wmbMQ41J59INz1Na+aPGuRgBD/o0mToxnmCMD3oDDIlJJlo
a0CeMu8EmSf+jM0Z/l4aApGKBsAvf9LVHx6tC8WUiViaZzdrtC/orCv4UkP2B2Uwvc1Eo0qDKSwK
mBmTjOW2/fyFUcjOnNIInQRkseApSTBrBefB/q+v2a257pDYbVV4JPro+WKQJpzf5rBCK1ZtMSR2
O6tn54mNVZAcBDnu5SxRyph+QBoT5dUK3BE2T69PZocF5s8CHRUQAkDTpJlaYyCgDEuSO+4vVj2V
Qb9YW0D6SJ1lSHm30bySzI3CnO/XM47aYhDDIXBaAK+oyBD0+AR0n4EujFKmTP97ym4m77zrF4cb
jTaLEfWtIF/ZLyaI0ci5rAhPRiqvRpNh5tFjTIHuv9zbp8H/cmxab37neNr7S9Aek86QMUALatO9
gdLd/kvMbW0c39+6f1+a9NRRrdGxWRkRLu6I726l+dDw4bz+5iS9yjbSoFRyxNvoXT6Fk/tCV78L
yirEFlWLbEu0Wbfd9a1TaMvL9xFr8obsIFhMd0kfaJ2RPpDhO7x6RXjbRWNwqnybVAoxlZP725Dm
nWQs0VmhxLygZB+dQg+fnY3sz/T1ziwItkES9/z/RsVJ55vYqaSkU2+5VhF8HXJLkeedcg1xJZdD
c0Z39A13fW802Oc/fAhk417hGI5+vE472SZCSNTo4OCSY7lJobGU1K/leQ/BUh4LJvWykvOppHYs
t6jbZNhmv4eR4gL+nvWBtRHTtc8bv1ld7zazQUU49r7nCbrt+fj/kmkQVo4HJqtdL8TdRaCLpx5y
/Pzxpwwsz6IWwdcxx/Qrci5zLe/Uf5auKijFNkxcXZ5/Swp4USZekaBTVxTqu9Fxcj1lL+5ETi73
FWIt0cP/HmxTAq3fnC4pr3JEZN3H5Jb8JzuXs2rIteqHls+TD9t3vJjo8bQuFgeqOskDcz8Elvbx
n7fJfauvMgcMTrXvyHiF9Hjc6qoK+6U4FCpwbX58PyrabL9OGUy6dek4SSDq75tn8azUWiRaqO3n
PfabcoNu7W+do48DUoPxslEC9g7XGDW1ELiU5WZstV019TigTbmfR9FSy2s3jUb3qqODltVdrlxT
eLMqODweKp/rfY6ebdMv8RRUqzFA59dqdevAsDAZSysPIzGY9jakgXoFgWCF1Pl2zYI4DdmKKQGp
5hHaEAA188ITroKCeeiCIn/hsXm1/uNH7hey5hLXtlqxcY7RIdZUFrsYdU2y9D0u+buQ42oc7zti
1wBN117rXVOVQfxjV+VmU4RViooVH9tAvdi27sQZUnDK2N1fSSLIhxAe7hVAV+UXwIx/Xr7Q5xTv
Ij0x/z8f3LB1eagnDs/atNjwgprHJLv5acV3vwMQOE7Hd+ZkDBPKVSNuzhLiAzQdLj4LX4tGv8pz
svtbC0+SrpSbuvbCRjUqQonVE9EvCV8pnMmUCVxYzzjzr+SdGCjG/4z30AQEhQOxn0FQ/Mv/Mgfu
PDJqkK5GD50p+urOic079L2hP+zYo0ZCMfypgYwTHQUAJT3ALKhrCbCuyjTUaBbQREBWRgclo/qE
3pRKNRxMUuS3mqvkihclwdC4ux/+bEJyE1iLZgmgTtnUIJjPoCZx7SWdlbgDFxkufrWUKqNGGFQo
c5pcunKj4liZIvMGWmC0huEKpT5oadG1bIn8y7TA1ce8M41esSPjiykJGW7eacq5ZVvtC16PDZxG
R+qnpXF9bDk65kBpXZ7wo1wt1/UP/ninj4LjKj9sSfF+bodgOAl5wYStb1kL3QPo5lgPxRSxof7s
Bsu7v9/wvvnYqYARky5cJncu8yDA53xbYivNt6EZsVS6Qa9hWWBq77HxOm7TUV8jHexz+Vy0Dzog
XET+ufopq8If+Az52iLxC8fzUXmm8ZsTuEyahqez78FnNdpLoLaOFtIcwdMURwETST6Y414HEA03
JvdZuCXbhJ5muy8ZumCepA23tgLR/7jpVru0R5DDXT70iw0SdGT/rV8+unMEmdf2wjHrMtxClDr/
oe2ST0UOpay3kaUDYM1j9R1gTJqPinDcpcPkbcn+H8eBgZSZGGloCZF+JQ/pyVkz61MwY3oKHYpb
fW0OoyDrA3aKwNXHEI0sK/k4nob4TFyvNNLNLgZ7haS3Gj060rhCJP1E0n9SOrVskGEfjjuUOQCm
1arjts0hzBnC4gPxUYjvxACoeg0W3Qyd82JbyeEikNC00dRqve/r7sCWFG+8YTA+tccYxjY8EyCl
t8nV+BYuqiQa2y1TovzS8Y7tBavxVBcoxoQG3ysaV/tDrNxbpUe8yOceXwbRmfHSHyE+tQxRvbKF
8smHmNsEB2omk5N7Gjaa2Roe7aoB2RYcGOfPo3RJnBkqu5WkdeniRR6idW+ewBNkXnQWj5OXKhA2
AyrsemnpZjWtjIjW7xZ4C3HHhUCjcv9fixJlSM+mkEFLUT6sXjp22PYcJrZMT6DTyVHIomvfnuex
8QVpW6wC2saOMx3dr7vgGGurqI2AordqpfvwamkcfzhMfbrOiNy5bZjtyNZFeEl6Y68vjc5ZIazt
y7dv6ux5twW9cSRFVuGmPPmC3r2nHzZ8HNgDw3/M1ukCJ1Zbj8DQOyBZ32nOTbu6fW05d3m2AWLL
tRuNjbfQUdLdJYRGwHzsDhdKOHu1kxE0zNzdFxRcvr0MknU2b7qMbyX2sYMg+DArslpt5BIvZrwA
G0fWcgP1UC15ZQU+URZecCZ1LQlLXahotSZnoFcTut7dcrNYh5iTzOlkqjy9VaK1FmedHgMUVwob
3sQPqxQuuVgI2MM7clUku3Zusp/Ruqw66AMuwa7zNhB8UuxkCnyJuh77r3GjFi/lfwH4J/baWvdB
N0GRGpkv80jZR09pVcV3xTdRptFS8MrTGVTeoc6ivhDi8g9Uinz50MrgfmXw7ptdcVud3QXjBR0d
j9WniGN0o7WmnIj93QHHjGEFuHGljmWe74zPmd9xfdLojsk8magj/7WYngj/eqS8/ZqFKG3LHntk
tbJfNEasiUtaEwnKJ8cVM7bNAahZvuXHhekbqkJSPmcsoSmGTA1Shlhy/7naspm1XmZyxLhYGEw8
Z1eS4gc5d6bvc8KfC0TD8iw1KMXXjm9bOze0XL3HTkj4z0O8OV7fmDGZ83ZwvrDfPvf1kev4j0ft
qjHUvV4hS4cb0hTpSnMaJyKrbiLoNTHCxstpHIKCHCqnRbkyRBktHME+fHmapID8uv1Kiv8ERpD+
5cR8y2Ess4tZ+ZisbyJJMuYU/EYFJnb3MhHqyp9JePriCqVxclKTdsqm4U43yJg6VQozXGMz5zA2
NEg4iY/Rkq3byeSv2vcGdR32nhwNFKFtj5C5tgic4xBzRacRGPbKnd1+CN6Gt6nTJ43WsVUQBxCZ
PsWmyGAkUhvfKe7cvciu1j2oCaNTPUoRIra6/QkQ2a5AKS0nxNfKei0tazB/7WeUqboIftSomcSi
EeSPeCS82WFLjxczeP2BRrH5LNjIbkkHmQwN3dEHxnSKpNlCWvTur34ekne6qaK5xI911wrT7tw/
qTuG6zna1nHda9P3HYWo4flBN0BpPNkiRKzL+R+XaU42zohTeCJx7s0WisxhwOaGG9UBdZ+X9ocC
TSIN+ViYN1oVparQKkeR3ImdCjQGLOXh2Npe0bljIBa+3zlyVujPGvHDrOGsk+j9Hv5f8cO3IT+f
8CSHaXfwR4bpVov6A2C/taoHZRQnHVjqQ6rqetugJ73eqIpjkMra2rnMUSBDDp/p/TVQHh+Y4bht
IRIs1BUmJihMFM5EXJatIDnZ/d2A0S3/mQpwcQf99f7aXxINRwIb2d8REtQv9btYVnwyRC/N5Ecs
x7ujvJdgK7J6x95UVTkBL7MaFSqdgoxwjtf4G15KHXp5b6f8vigJYAcrGCYmhnM38/UL0u820p6d
YHda1R4W7mMZduBxl8aupbKmefix5ISmclMR148cgmvXa92x/Ss1Lvywv/TA+tVo5TEI51XrG9GR
op6oR7KzTJULVyBQpwuVWsYhrOqcQL/xQp/qOJMc8ULSigjZ0UgTYVDBd+wwRr+PqtMMHmlwv6f2
e1tCt7BSlyvgmB5SxmU/zq8YRgXpW280l+LHlPiizCIbPyknFH2WfyP3g//16ZG4W47ATNUtR79u
voj00vPZIpgjMBwBYabq2m5q1dCEJfrTJBTvrvVnNGeAzabEpYd2Znzrz8O0iLJ5gwgri3zD3DqZ
HGiFytoGfA1VKKUfZbN3z8o869dk6vGZ9XAUNXljwtJ2Ijkw8tltj2vnvywdtFc5Ap3P19r40FSr
xUwNQaCA9IRzgB+czmpeTkRUGEzWPlHdnVB5zX9QvzaJ2c2PbZosni4rH80BlvgJYQZ8ZG0skZIz
koziu1alG78OJ5WEuQZ5zDaVy0dJV8ccAgSsiCDEWxBO9I4403z28Fp9/wDEcxlQ4gs6FICFcciP
tvJV56bAh9s5WsV8jZde0vozr74yiYAp5qMaZIwENSTPRDkdoH+rtyvzibVxOu+XZd8KsJlq01mh
l4mnJtsx7Glp44bfxYY0ScoajVa371WWBAULJ077qDfwBT2Ydacr9qiw5PTob21GLMWtiqKYUYZA
qg6kkEOqs3WnhXAvqGRpCjvkNSW3G1zL6YwLkuXeTzRP5pZim7cilSDTdAOpZRti11D1FDQ2HvqV
YACBB+r7B71M3IJgeO3Adeh8D32x9MwFV7SBZOjvzwnqGVy5LrRs0P+zdgGZFEjbORaL2/l/MqkA
sQvkwMPwiRUrZGYDE0vUFJXViXPwloPtWBxXIWmh0DKJj2tM6TmC/SjLvPYqxO8uByYjOIrSYH71
xhZbRYi02z3GSkhcG1kQPZcDSt7gEVM5PheFJPm+yGEORjKPZM0znJa3vcEDnmchBLXkjhCgT0rj
gpgJrVetT8zpIlXiqs7xcBv0DYbrsOyqZZ7glRuRAD9lf8BXUImesufeNR+TNB1Qqik9Igd4p5H6
CCAbWV4jq1fyynRd3nv1WyaqTK63pT5ng4xbPstfKw6AIpT/GG8YujJFhoRC96KpcJVrGyguDi3h
n+oUMPSdna9wodTXpu/RNeuuI9JDyK4FPoj/flcEwCdeFpQ0egV3kuTzIruVYELq9o9eXIbCxPaC
9jAFq+G8jHXj1UVP4kA1HjnYG/sSMJAso3E1utwCFk3njbO7jsMhhglzfGJGzwPLRh8rPG3CqEuS
FBs732PG7WXqwCPj2Ex3+V2ZmJ1Bd76pBxCfLf3vYLwnLoBi7nLaERSodwqsc+10nPFlmmIA8sv3
XD1xarQ/80wOTKYxJcK25ohu0Lpdu0kN1vzfzPWHWHZpQob+lZOlrnBe4YDjjsbCjLXKRJHgBq6J
8FzwSEeTgeNw5KSE42UZ0I3E6yINRuJspBdbO5I5DSbzc8GKNgUdUQM3VOWll5tgM5x1bcQ++kJP
4nmGic9381EbR0/yV0ltwLTHHZ4mJv0PvlEoEokXjqGDH8z217CvVw6HGG1UVWvR+WsgWRjw7SCG
k5TW1SLVkbG8vAxiI0JFX4Cyn0QBojJg8LF4bqBqHmwz14+SoVKrTtzmTJ/iEM9BjOAe8J6LR9Os
MtbhKCSmcE7jN/2LDbK4EpxU3M2Kkc1iqJk9LJ4KneEw/uckO5IJ+nhYrLJyx/Qzq1W6gb78poeh
aABpeWtyg9vX+sywxJr2ZzA44FRql3OSN0Qs1vGvWho3hF8baeRN3uwosGYvVN6KhuOzkZqGrjJU
LgXR+oDiJoto9r8S5I/Qi60Z+ZP9b7Jtj2nQDrD8CAoyEWjnDZtHXwvW91YwvIUCB7Y4toBZARkT
38Ny/83EzXvQZsboq2yBLWVbKoZHbnyI6od6XrXV8n5oE8zhV2QaVerS8ISVyBXQDkNH1NEOe6kt
u/1s6iI+bpute/Y3atzopxEYpRdyRfvaqMFQW+f5XVkUyG7iruZGcNWda26MKUwJPHxLngU3dZq5
mJB0L3Hmx9pHNkyZxsinMC2qoMJ+SBwVv0K01rj01nvB4ne2Hy80mtYV6FJZOnaW4msP+PjP8/tI
KmT/8FT4Z5jNcjyMfGKxBqw7WDS3BZ8SX89vSl2LX7kB4QYnIktLqrUSKpNoln1BFglZKBXSFikO
tQC3Km4qDdkAFeDFCu0i0UztDRjCVgmXuwg2/XpAQUhT6qe5sLBqaqEweXI2aEC4QpFIRP+hLiyg
iR1OYP+7cSRksj7VJ5EgHE37K0jIxxKcgX6DKrvqRhi8sKD4jvya3iDDTSYmQcdkRa3orDugtn/h
vrhE3AAXtm+t1/cVOZ5PLnubBfq9PBn5DEJv1KwM8yI77o4qhBMSNbVqyu18w6fcUSvZ8FLfAEBi
RF1bjyreY0wRe/zHjKEZmupGDpP+cFvCNo36dqsL9Dc3jsEfploH9FX16ttatFk/Lyz7c7TmTrzs
67eLu/ULw+6M/VTRTqbrPife1dB44nbaPCS3hTCIfxJslutPH2v/Orub/QHp0+1bEHZuN3mn4SVo
A4ItAhLzijyLMBpegB5p5v3KVEIjFC6u4KY6dng/L9huwAiauLk8WXaqMCUWlxn8BubrRkRijfw8
xLGj1giuu3OFeMfuVljBioOU0++/KbZTwwDVQ6+ecQhSvZV7p3hrhdvWZRGVNdeLrsOxu8eh4Hwl
l2ClSbFqAwnLwFQ4KQSgD0LHUSHWL+SpD3dJW5pPwBY1gXxhn79dBv8dlyVWh67tMjb37vltugvj
JCOauDf0K5qZygPv86yY1/+Km9iW9u9cpOfGxcJEo+sVTGlDwRR3mzPTaC7yJs/QPAzBvBgjUx2p
JOO5lAbUD71+OnTmqmM51awf0mPT/2k3x7o88eL/fS4FDp6GUllKDa9sP4bJpGve8RfUnD76BueL
Nqytv66d8M0HN9M/gDfMb1sh7z4XOQDAneqeRwNZD7IjOUkdrkdJebcs/CLm4BN2F6cTI6CtwldT
usyTTCp4VUvKtREW7DVatNFj7ESnpZgjY0s6jfi+vqBHIhSBpUxyYyrNlNRWtWsaT4w3J4wOIGn7
2K52uRqf7N7sgH93pa8cToEuoMB4ja25/0nKKuM7Hxmk28RiD5txj+mjX9OT5NfrryfKdmt8Z5BD
BF4AkxSU97dKbkVx+mwo+c6guEqyq3wbrssRFuNVb0pQh64zF5Pn0xd25y1ZoAHpNQIkAUTy5Sy1
eHYu+V1I0glvWAOaLtxY+oD97ln6qgxjnJQNo7SXBOo9wnFaAl5KG00F9obYwFXg+fh+uc3uTi0Z
UiFZVJtVcshhZk9tQ5VyTj+v6YAVytD82qlf2AzED1yh1k9qqtxx3r/qFxZd5tfkl+uaRepyJ3iK
Eh1IpkPT8IsPiimCzHkumZGbgnupvblHCC5JBYMkI13Pfv41F1JNKwXxdwirMgJCvVyg/cJsnY2f
zyG8xTxDujmI5ZGdsAK5QPhRyNRnU0tKgxYx2wTnh/qMXJ0+qc0+VhHB5gBYJkiAnxAtLsoqroB0
aqmff0fZycb1k/hz01/y3KPXffuLw4chOzqA7Ut7v8mWUpLG29b9y6fioLc2HU+bnfJx/fwpTKnJ
VVWFLLL7gZYCnrHRwohnUqALvLvPJH+WobwsbfMnrralDij2ohzK9u0XQ2n42enT8b0JRTQNjbmo
wbHv1upxDd4gCVIPhxJtiNngZsjf2AdtzWmuZ5YJS2ZEEg+k0dS14mtrs5Cf4VLQhA9BWEmtd7/K
dgEfC8jwFL7o9dafj7hkxAiDI7B7ymddkkOvRqi0ojepT4QYRoDvAr3fL3Po2kuL9mkxUugGaN5u
GwvyOFOLhawa2mdej4XJbrN/hA5uwBKgBsGuy59U2tyqFGd4qzRCAhj9YJylpyLWaiD1Ln5h2hVk
VrX42T0AOPXdAm6kRyhTH9Q1EM9XxfX4hkavMFSiFWOtEGp075VpT+6C78J3LJeUEY1FJegodZKE
DYSjmyZv6CKcILyD6aonTNgvZH97KaqpQUeeZ9hlVys0Q+3qN+vEcmLVhU81x6HU4Jm4F0vgsZTV
u1mt8Zc2QomZR+ZRwmvAxj2Nw8PxDZqI3tYeyBOyf/FE1Qsy3xj5e5B0L9RQKZ1btB2hJUNAoFy3
HOIvBpgGxuRSPBmRBx0ish21+aKt+lEoOYhjlkNQ7ubZ+7JgOZfChP1k8XAcfKDjG0kZ9W9kR5/9
zUX2iCkbFtrrpFiwYjwiTGrtFxGoOtSIx7TJ/TyJM056zoG8FC3+K3HQ33X/guu5vqmsWCN9h3Az
Zd+z59nixhWhriBt6UJxt/yS+IAxidBvIZTwMD+8g/vrZyQDqAZUacsVxgoCEBuOOb6DU2sOGeTv
sv6rImXaTDLsjZOf7nm+DCMOuYDkoxZUnZ3BMsKYks0NXXBLjvfZY8D5Hw90iYgVACD4KnRaMCxk
/1pcKNChxezxXS8wdqDYVRhGju9zKT8FEuWLnsDYBR5Qp3OT57u1q4bsd1gjMcmsVaSIqPMzaVQ8
znPJKxbN/eTYfr8hoPWwm3i9ggmIVeFAqCZXnIyPe3Xg7NqDPGdqoLKOyuABL9SIJWEVtlBSnxxU
A295ighCgk59NvUmdaO3VEuJeBXS/q3QU6Gb1x+K0sa0AjifblrsLSnm3RChlTuriBjvLR/My5k6
MNw06GiWU5o+aLD5QUGxS82X3mP0YGI3xz3X7R4xJTqC3vpf6JIPLrwltYUW89XAc4OxJ+XfyLth
2nK/hcq6dG1lJEHxgpM/iNGh9S+rJYu9Vu6gddMYRXp8FowKaklcyAyludX0/meYBppCdvxI4AHQ
x33GgpfxUgsNU4vY7xOCshLrzLemoHpdPH/2rhjA5ZIQVxbXhgmHGzWrzv1vuehqfvZqjBYSoYVs
zEyNhC0lTAJppe/5gew47fE4L0LvHSr3v/bgOU2lsRQ1Cgj3nZ+GpLDkz0CBmNZ7IDH17Hv+Hc1B
RIQLt76HeC2B1NaaPLMMnBOKOa10TCfWdTTgRvAxaXRk7WtTseFta15l59mTIyMd+smtlYvAXlgq
jMlSwG69Z0LJemL/EOrST3Q2pS/+VkuX1uaIXcYqhfQqz95Tq08kmKxESNQUmZQQRiio5ukXK5F0
HX89xuqn7YkpQ6oJiUtTuZDO/wOlGvZcNXatCgAeavG+9rrC9hwoPMVK72bXIwRGgFh+kGrLLMpq
wffa0QpVxW+ftiSfuoR1W+94NIUeJGQlQpuew7dI7RfoRAz9xbfsLHdUcF6iH2BTt/jBTIq1D+P9
/eqt2kSK6/oVARjz/Ct0q67Lp7nG5juBgLlwbdq39clpmSWppF52jh7RUzjPhum6Q4c11gH0J0cG
ErnhdJMjWxB7t5tMwMDrBDSNb46FaT3wg9hKBNk9BHfHalLLIettqMEJZUDhSem34JMlLrKu9P+K
yPB+C+w5Nb0QlCUuxlhnNOGxAUEA28QLFcS3n/7wqgDG1fuhteTnUnU8QARn8MlGDFfcrXgVZLE7
T9hnxo6GwKsK+ub1p2kex/qoSA7R6EVZ4bzXvMsz8RE9gqi5JDIUPdeeKvN8nI98JXY+R1cKo8hB
45E4KQ9OLHtgNCpCqyWBoKh9Qlg0bmquOMvrMAVeCkVc2kzo9GRGoyDd9t1qKbaRsn9WBPdHarIP
EXe0lobASBvPLG/9mQEmLWweItyNTVUWpWvDZM7xaEXL7qsUmcLp0F5qwhO7To4Qk3AnJtdHMHlE
oexY9+wmEo8L9jtvr/OYdw87rJvsgVNIuwv9MkQi1t8tdELnbm7A1xOCQlM62wNzs4YY78WmtpFT
gwmv2LY69/qoZXadSGBp/sM007Fezs+P76Ivd5/MltrEf1jSzJSPuJSvxlAaRcqihhRY62tdx/qZ
JdrFTSTGS43zBfahnldyjRYD+MasPd7wgcM7qh8cvRyjkd2Oevjkwd2hhY80H6uoibt53n+az/4I
LhrIq6LjFc4NkDeodobQ6A7mMEz/0v/FEz2/yKZWspvWj81vmybRekWpFnmplh7KhiT4ERFws/Fp
qSe1vMHadbAt+zNxAd+Aq9UCtEG+Mrl2AbPwNJ3V2jx5wE97+DT8D/HACWoDN2wzAyySv5FmOV/x
wp92qcavvka52qFFnWx62jRgBJU7d07cgOMbQhKwWkhb3BMTJZ4h1hlDqFES28U2iIILVHpeMnH3
PKcd1SCgGxb6Fdn8EOd9nIlnBdNV1lrkEH+pAjlsSLZZhlyXTcE68fQXJICVB1Rz5DjVX7qU02lv
ExYWrHXKSP7LvTsgizI0/ucL+wgECgHYZtz6UmS+br1SZqgTkCUdJjBkzeVVNt5Z6yxqmRDgk4bN
Acj8/jZHKeaGvxLyHVJAzLt59Vo/kNvfhyrrChWxfGgmP7Ip0bEJbnFjJn0xSEeiFXQHuBmfYl+x
0lau7H06kNkkagkNRZxt+G26GmsV5k4GJ420r6nq/incHFPVnepMhD0sZEYoF0b69VxeJ0/U1y/C
yAl26A2k6Y+DWH4D/M4FAIlOkzFX2WQPNbNw68W7o7KOHXdzny313QW7QowA990P6JDMkJFHVY/h
suwiI8Ek8OPUw3byWe8irTS1LASxVkqF1f+mlmsRtV5tGDxQN7ovi4/M9nLea+F0L2yG2csU2Klk
GyyUQjcy1cjz4CMIpUaGLSRqtfE+B1rujXQcwxIxINCzHcI3mQrSjOVzN14owtpCZa5wZd5cgU2S
3qWqmyBiGqh4FdkkchMBVluplnNtApUKczOpt8R9Im++BAN91hNtKSGaPlURyMam4kFwKPm/Epyr
MRTRwjVN9ID5bbxf/ukTZKdWbsB5Z213tKVlipfQ7u8eRvG8tpdugoGCo3Bw6ePQLKtziCQb3vWA
D3FZB0tgLarRgLTVAdG93uEERzW1dYvOVUr7YLF++yxD0Mkos6nYHmAhzR4t/ZrSeM0GwO6dyFot
afjP2lqP0AI/Tbg8vgnhW5Ua2zZ0MUqK3wiKgDdCMQxeOpavVWCeA8/DYUjY144d4WppJg09cUYJ
NOvEDZTnw/nMxi241uDnrsAbC1Gn4GzX4TCCVTAaHo1aNzO4rugt/DZCsf+pgfRRw6ojX+Nu30y9
LBJACS/xS82fp8ayqvIgrh5O9lcYE9JcDEw0tSJdEu7WQTpDpolDAsKIsrk2oU6JsylAWpGRhCRm
4ffWV0y6ajP08xdYgWQq0bqpOglBEnrxD8iZffgAYfkkSK+Q26rLy4HR/oBk3vJ/7Y61Ls2ZL8gP
TK3/RRJ+MMl8KFb5vJHkCUxWF0JpI85JAoRjxjarNTCnxBEnQAqLwsOSj+oPNSiSk6LuNGjWkfYe
FsMqpohWUo5lqu6nmWUM4wfQVO2rnIsKi1nJcclVyfd/KMmFDKOELIKi3pjlMxEPkDRT7gIlyh86
W6V9XUbKH9LCvidBtS0kJKy2NIZk612R/a4Lj+bDnk1Q3gW4wTIEB9FETm2x1d8Egdyc7ELSCDvV
OBOePHnax4k++C3kTX511r3aXsdEsGjYoH7sGbFRMU1w0NdlWyOKkYvps2R2Ju2s3l7shj4685Yd
0s0d2I5T0C1mSqw2ShcN7fXQG05Y25+uTVhX22xNXB4myQmhoxn8uWw48ZvblqewLOBdB+l4MIfp
IFXpnBKIQr5HFiKrAvzCZcqa21oq4yIxoEccZiV9CF7y+d8i7LQBc18CHggEYsAopWGP5sC3WRJE
GCV+mSkc9OUBy82BbRYAfxXf3rGgj8WWVauIT/mZgkqCtbua+shEG8xzK6vJmiCnAexRrEXAhi38
Fh0OVEPeLl29ZdlUWwA6oNRZ0mz3CBYVOo8RWcQAYEM3Tr3kfNhb+mmLLycUBS9t6XvqiFl+583F
+YHirSmBR+lbxN8+IQ1E4IweUxLl4qy12rlGIEEQYHL/xUPwtnEBA6piVlCJ/Peuc4h611/94REq
6TWLi4brWdJG5KV7A3TNP93+sgZr1NFNBAECY+M9/HnjMTrvBzWPjL+GASYmAmhkUPW58AAoI7Gg
lUQ7qouRJsdgafDCEWvkgmW7JnQgcSFComWSDsNZPUxHe84WkwXmtXsDvvcbp1dqmT+apK1Xgwom
B4koUs/mcGpg/1y17lBZIRr242cS2K/WHvWP7k+9n9sEkKtUkFD0VQMh1y3KTQQoK3joR2bmeA+P
BXLLVa+ntNFkaBLlbBFotBeTuqSAoSkhGADgm7jyVHiQgmOQpX5PZkBCxK8wpeNA1yMzed5FST2O
TzUexVAGvVm3L3hmItidj4DxmMUdBwRoQcD7Wf55me1YLUDwLo2n0NhLw+F54R4QUCH4FadaRgI6
4a24Nu1R/Xy5STXo+xChtmgv/IrEOTzGtdAo2gteibjLag7vSqiQhfLNaJ7aytwE8aGcZTj/JT1O
DvN66h4evd6H3B0g/Y//ZyyMY6W00LU5QIz8XdYwfbqSIqYUzRaH38+egeWYIY7KI4U5keULfX/x
avjqnYUQvM8YQpZreXI7jbNnFnewU+bZ1P2/kIXiB+hNtyEoNexGjg95aZgdgYUNaPS/NcyOOZ0X
gvIPs/wfJR72D44oZlcE0uaTMdDcjboKiR/tuN7T3EOIAECIHUjMYn/MJj+kdzgJi7T6bXXYsmEw
JwkVhAtirQwRKv8jpF8GTnh8nJrpnohDtbfGkVo2B5I1JnpwKr14voCwKFEw3x7sBwKGH25vKoBA
IEelQQl+/ZDbePOq0ea83vXuq136qpgzgPzaTN4mJUlpNmW8+aB+blUWjpLoLfBesocL27pxz1Ow
CbWQtxCELi0cfxyOAj3csu2b3xogfw+ONmFKX6uTiJbFeMZGwRpX9Os9A//hb7hqubWc9Vl6eSYU
TO/hCVpZaBZZbnU7gtyvV/VVhlTAq7kboZ97lBu6s+Gm0y8Q8/TtB977LReThBFbLVNbSaxcG5rV
c4tq+fLbuuS2mZ4YuDH7sUDRCvZJYQ9f2Tl3GzpjloSf/0FMvDT6iVaAEGYS0ekEoNu5jbFXnSjY
tenVLWi91OZqqC1AU1iF0RWNvG7pBVB0IZE8XTXZsjMo5wdXsbdsqJkO5oTH0FDLKlzwvCxCaRpr
San+VJOhhgz6JA3a8FNrJiSx/ZM/jAxzEQi/S7aTitzAN/S/A6gxTMlU27ogEXQReIrhl1zkMw2n
FG6ElKWTfa/IPI1i33MUR5tV262H0O8zBZb6kH88kC2xUn4/XKyAeRPtjuL6G3d6sv6kPb/n5I41
U7SN/RnMZwMFBvXTbAPWGn6mWtwN8ALvosY0FuNz2wArH02FOnYQNYUlZlT3l7V3fjqtHQGTZldT
wWpr5pg6tA5qQQ00NvoDyuiWUebw3AQfYSQgl3rawo1H78T/n3Ggow/B1vbcONFVyV7402jOjm6U
cwYK40e334aFYjacAqbb/YZT7NJ6hFxzuUQqMo6aQq2VxYR/O+IfC89uP4au7Tc84U/S7Nf5vQkF
FjQBPETMnL9xNJheHNufBnYNSBwYTu+FYKHyee9ET4zyeSWgf5VXtgGTpk9hHFAChcsiwlzilI/z
C92208wQTtCnAMrj3RzZcjPvtYEQUp4dXdMsBBbLCt82gA6oEhG5DTbjNZbD2qbn+d5ZvID6ho02
IbaV/OBvQDWMiMHGfFXUq+3NohRkmEUxSqWKv07Qvj8ZSv1ery2GjFN5pvRcUim4dWyqTyXuLwvH
xYr3uH4KDnlnX8loADH4Cnab1yzmnOILE/IZm4ckK7W3zelRa6BEz4d1lM8nOPFOw4h52ck0Ckv9
KXb7n+iRelEEaVbWb6iccqZAFKRhUGnqJXs14kn5iVzL3xEHkaqcdY7dvg1BRTt0s6UDvoYXuWn6
3Bxpc8WNhLs8agFCcYr6lUSTuBZ8GNZRXAWAm6gr2V8D8r94CQ2II6FC2ENiGwnTZJ54iMEy2j3t
2xn25L3GwBDx6XJk+Y8Km1UiAy1r8YVfCtF53VNHwwKs3JR0hcO7jeTBueWuk5rPJowAyrh/YMGi
zZ2u/Q39hKNkMZDEsZvW8kw7Bp5fYVHfezHK6IVPFvNe7OEKQKX1t0SQDbYjhOZVj5lcoyFJf3vH
8d5IAJG81RLZcGd8zepfhEt/RjfISyXdHA40o8vv0dnnRe5WdTe76fnDZSdCO5G3fVQlD0MwcA3O
nmVZWhXqH064G+Pp5HsYQIOCZvyf3mEf/BXjfYqy2msfj4fGzQxeCQ8UKrL1BtnfYUvvXmj7ioTL
+O+PAUkNkG0fvCZndDTfw1qmH9u9VaVv42RTVmD/tdoAlp/J5TbfXmUm2TtMxTC8ZFc05vE4psc4
OuW+nxG6TywjUhwktrJXtaTABz2KPRWIWXmXuyjTmGYJkrflXY3+TAGJDmurinIC31z2olnG3xef
6UcywLSns4VKiF6fVBil8BYTDpZ8WYxI4HiRQ+cpyhhV9CxIH/oRS3bkqajHEKg7SKyZMmZhvYfI
8fwwI+jDv2eH+MYg8gerIph1lXVjaVkNg8j0PHl9qcr7oPAwU9Cs+FSaLqFGrjWvxkS2boBhdqHr
0hCM6hrgEDlBaCRHcLvB9C7LfRH+uFgtvNgR8gxMjWpq1PVhgaf2kdqAWrlZhkoovmdXWP2r/igC
WX38E1UznKtjxRXNOT+9rE2dKifmn4mpTdXqqpaE01oSsTGcLg5JXWhL2DoAUeypynrkYms3FMGr
9Z67EbMNa8HaDcC3nJH45M0T9kVpZ50gAcis4OQvhaHu0AtP2WwrE9HLIhODECDeAj86bzLQj+FH
4opOV+HeQzhJGWx3UzicpsHEgDZTX4Y7f2iT5F8vBl/d8vYZ0Km98B7fBooRjHmq5RfJ5FmNHrld
DzBLUEDWNuAMHpobJewe4cs1TrCT9GMRfxvCsC4QGW+0Cb8rlSfDOwtBxg3iHfNLN2X7pQNuq8MQ
1xqGfgeen/Pnt4IG4m2d6h2wclnjnvdJ0I4UtWXK2DuuQki9tqvHpT2iXt3sf8wwu9XCAV8kQiwe
0LuzqsUk+/m1RJMF3elTvp2rOa3gdRYwS2ByH2Tf0iWJMFh/XGXSHNfP04F1Z97UXSVYS2dYpJ5m
OGK03GQyRlqpw+K54lqbo13dj5ps+nBR2qpan3zGpPwHQRru7hP5/fDmqhCXFC0k3YI7OC9EFRXh
hlE0UfGMwcljGhfqTLN+1pxUt6EnqJVzlp8BnTgEWR84CtmzHdM4iPheofi4b+7o5n+cHspk8Uzz
t+COM1xV3xKvdXbCXFgTZu5w01Qc0Ukcgj/ieIR8wxlOVvtJ+ljgU+QAgAKsiY1Oc2GXoqgpeo7q
nZ6J66IsyKL/49rPRByve6r/K3MUz95qS5/qvcAXZyxMyzWsUTrnW+xn+zZjpEpz+ULusHk00pB5
GaPx5G3uaYhYbeEE42gGZvzizzp5FGGA7dQi5xpG4MzVPSwD3IkR8exy/UtRGRw5a4pMINkxKhg9
eaCJDzJ0gwko1nMrYejY3larS+kry3VDfofZbbeU0yWvTWUcluVGmEUEE7ejphZLhU6DhLKf8zCi
C0VW8m+JfC4tHXE6cBtJsZ2XJngCn3BESahFdSX2x+AY+rXq3x1xa0+3EEGgYgNmBQb8wg8TEmtQ
oKA4seWTX11SybX0eObZBL/DSv8WA23o0LV/h/fyDBsdnoZiGZkQ6mNKnP/2fAs4HEBwb2xnUeuz
GZ73nVfW3G5KE9J+ZBB0tUNeNxwjg025/h6IydGiYmz8ZaQlg3iQrwdkq/JzzkhvXizXav+uz8cP
q8uqMJs+BYRg/ILGpM3EzgxslDMhMcyF8RWDq6XZnaVghXYQEKIZroiX2mjkcbWDdUoKaVmZrYfJ
95qML6iaaS7vcPQA4qM+z8Xtnw0DybokriKJ/eYlsINAckKXylHX24N3o74afcjKxtLjPlGnkoco
cAapzfwaaDOHpnnKyTaj+GRy0/L3aurxRqEpOlwYAU/C3JDoh2L+6GuNcsI2m3P7+KJ/m4etZ3aK
Jfj2FVWQcpd0+PXz/O1eLPdXGRmYgzaxmNtjO/jS9nXl8475+90ytZEtK6rOTGe6MJZimva0NQfj
8UDmHNvK7xxIF54lCvwuI/MEYbu3ECZcPDABdLplrUEdknwXABPbh6YSnrcXKEiY55mshLpj4Koo
kefbdc7nYRL0BSB27k1qebVPlsZDMG+jGV41Xc3nK0sDNFN8rXAA0Z7G7ogisP6p/57JgWBSn5Ib
JHLLrbUNQjGruEEcsGPV8Q8G6MWtfmuXCzY2CvdHm/2biMH5YsSxyl3Exjvx8hH6h8oKPqvT0ddD
T0Xf8fd8/5/BIKt9E+gpBIqd955bkFg8VTS7yrb/g4IQWn4OwJBwd5QAFpc0ksnTeb4bN4kAFZiy
yXSX5rwmovo5z4tdJJpHr2S1473qz9oWlrYW1/5aG7zB8fnfv9zeQQevQWWw3AfoO1045KQ0h3ix
yUT1PVrJZecgBBrTJNIQGOZqdDrY9mwW47l9oWEYKY8F/EPdynmIPT1nZ/EpiWYK1Cqd6EPKpVgK
GeyxUC/eIODTBoKDkuoVoi35oMMSTkTl3Hr5GUdGLCLYS4MbbrrMi8G8Oc+3OkzAd2xXGp0BLoQl
GDyrrbfJFhiHwQIxgNYSNpc1rvgxrKU5/k/NyD28Cpajqf9Z0Uq1ukWGxN8EbBXqHlL+uSvOlTEL
sPQU6hnT0PCP24z8RwiY10Sc0mqeEmHcGgIUgPCULl6ZrZRissWjz0iAHgWpRi399R+fPkq9BYFg
UTHWFse4YztygnEqc/e9mJ3JVYURAVMqZ2fmbGIRNgOrdI4lilfX9EZ3jspPDMfTuk4XfU8CCwLy
TUln75w8T1sGtszU3Mr1KRaZC/nzUTt2ulv46o5M76SOVX1QLjjkRYrwsu8pzXI62ttBrPZjb9yk
ZH48PflZyQyovlGU26CBrXh8vePP9eN2FIHUuIw5Pkp4mbIXVhrOapGexN1jelUTwjXRy0D3X68s
IvejbT/sHd8scRDTPSAxDw4lt1we85SiWwh/s7SRYg9UM43kmeKWVFiOyv54cGGtSO0gKKFkrID5
493rKaoEnZA7hSlVweYEHMkCnd9twftJD1IIgLYZ6am5brrITti2896Pi2GTku8gLRttqzj80UZS
plhoP8XZd5xC9HD/UQAjKZSmEJ2RpOtvjlvOfJv3XUtrVXjujjFU0UJ3oWPYkFP+AGeKi1KCijgz
hezbp0JqAm4PwCAZJ2B9hHQe+8uKkT5Lex5E0loRkGZMbCgIuBieZRj3D9e1SaUELvYGY4K6UuH+
HoYKGEReK4buTSzDAyMBc+rYSaS37hJo/nvIL6iI9qepLVVw/wI+99/PoqDbzmgLVCA7JHhgy/+J
8BDfZ2A3QAFlWTWvfMRdfQytGHkCYYzgjC2XlfX6ipVfK7B84M+I3IbrRadseXL/qYScXGIe91ho
IBSltEu50YaphlaiUJ8ebjYHt8j8XDPhOPIeQj7+7mF/lIhS6+d2VuwTWVXpvxUKDesgkbyToWL8
CMrvg2wNnfP2wbaya8vgDaCm1LpuXpcgiKmO6i9LNHv2lchC1X4oW8wL9TvPxxIW04dxvAeIzDkI
AQHZhO+spdro0roswbf6lRKVB+peDgBqOi6hBXf0kYWLZKaDyTVk00ew9IjTgsalpu67tq5bkCF4
tcPD53PtNnNFWt5iIKBKdvo9aD3CLF9nQ9gt48zXhl9AhB1VzsxHS694Kwp6Y9hXOFZcja39o40J
jgB1QnjWYWUVbLYeQ8lZhIxRaaTeKRBbOSSHp2eGhQr0bqWvvN/t3ajF1F4sUEMY4kRpMgg/BM/O
1ER+MwnQgilgaEaJ/zAJG1D0hXW6TV5j6z30u5+0BdxmG/U+qWhcwQOmrhhgAJ9CKXz0m5d3DQMz
KP59psDUbV/jyMRZQdNiBMya+G9VtCATUwwAixQsxnmqYeaKHc0WkHPbUuGjj2uoeKeljBWPToBb
eMrqkztayUDTMcnWGCTsOspu6zEAJz0bz1HyepSG296PH0pb9wszBOrJ10nORtTJ2rjvh5jcYm2X
duYni3eAcdNzD6Gvym13xypoyrqSXJFuRy3f6biP5OMLDCDMK1HKRYjFPGuePp8Rw+2t1Hw2FfZa
Zy+aBKhVUG7HgyOe5TtEvy1YjVT81mpigjEYwMoJ/9QE5pR0zwkfUzvuYvyj5kK7ur+jb59dRyiZ
yKg7LHcS/4nvNWQMtue6LjquMefvVT5K9Umt5f2D2Kn9YTCz0EP64FqhHlYTuC8JUDRSpiEimx20
jQIUTUHUqX8ASB/UtejrOY9lvLanabGcbnJWvu/gB1rHvU/4fS9+gnjDr5M68/MNEFGap/FoWuaa
PEO2nLkOi2eI3Bnt/hUS4spvM4cJjSO3PRjqzRNmpY7mEpNaxtkWFf5XqskldyZ4mJahImVMfLR+
xJFAR1KDrgSpz4zZQOeLo19hFwHb+sKxMTwt6AtfwnX6leTbGInVLt6GNDei3txUdni6/tHw2YN3
jkv2jbc/SVsYjnYzOGXodDnc9i6kIfxRIdz0uyk5z+bELq87Ym3OqKITkLM5VsUIGEwKo/5JSy8i
IIRMiGkRXbm4xRz1Wi+H7GSzLQPhFpZG3KQMynnXZQR/z5qTqHvtSrgCTcimBg/SkvX0ivYz/NY3
bfqu9srH8tgULsKVvBmi34bLlGztnl5mBjyGT8+GeaAFA8lF7NMjeToaz2eBemDIv6VherQv7URV
eKi8yHDPj6swGNDGKu5hSq+GZLPZfAEaDe8qGukzjit6BDQCE3fR1IpHQf/JkG012wznzVbOBEpR
WZ0Bvvjd75j2OSHoc+yXH3ZBPBMR+NLlB8sS/i89RQX1F+IRDhFkeqGafzWpab7U8sX1rJYpZpyH
TFByvno4vVuD/uuV1GTXfShzueTBrNNIPW3jN1cpNCQKc+AK34xo+ZZUNhcuUlCCSsxdBnqZSJrA
PxhnmvfwspPXAvqDderHMpGSvzmMPVdF6vFYX5IzkZjIF+3VcGPZaKd7GeZLWjNHQ/+rhcPP3682
wr5/ScB6uxV1jErCBApD9dcjPL5yn5twB1ssm2R5y25RC+vY6Tt+cUPHSQYCPcuytLLD/gtkcQ//
nFt/Da14r0M+MOAvwMYk2yyvZnlFfY3aqi1w96cPoKbKMTfMSrat/EMVIg05XMRZgwWHlHuaVtmV
gFbi8eVASf5JklCNnj0pVXD6tDfz+Oo/HzGsYl0EDAqfXKwGjoh8wrDmi0+A3aSwk7FotkkLPQjr
m+amPDyl0kExS8J2lRpiXPyJMd6ThpmdSZynTpWLnfKGtUBff99k/2P+LkVvX1XUrWtx6QHMNfU0
K1ksn/e7xNeoaXG4KfNRiGPMxc1NLnN5kjTjwcsQXeii4vehRqBmynpobFxcP7FPOrrRbDY9brpF
Bc7ALuDVVelzklRNp2UkVQ+1M++3zdW0W0kg9NgUE04G+TTh1zAgYakutnzc15qefqnxLCgeAR5P
fOdnwGWyWVhXTa9G0cb1y81C4sfe+77xYTPrJ+KkYGq7y7vlrAtv03GGH61NxWtlLM11wObl0B+h
9ifwjab+M20BYE5zxXLDee70E6A4sFu0m/ZxkD7/fz/RoRZ6MIjq+caRspR+JOJIpigillodLeUZ
T+q0XrBdeDbPPPuRrBFDrZgapGUX2U+p1msFEpswT9ohTUkEpAQApRO1LwBwiYCs5x86oKS4vISx
BF1Rh6Ayq8xt+C1OkIZdb1FL+yXNdmFubJGM4BCZFx/VjQYdvnT9yXHgt46g5zUIJDiycEoK9lWM
cId9GMaddETAe/C/bLEDOBoaY4ms0uQdPeF0deZaUC4fU/efTiGqMHNkyNNWaDgftm53E2X5fhYu
FqUNwzALOyY/y7hEKEQQsDum8JxqIKjhjNvnQRYKTEKD2q6jlZlF25QfAY5D7MQLsDrrh7TTqbqL
JlbjnrwHPe/CvZ6Ryaq6w1L23oIjtwO9hH+DEqooJX3kDBEeCKtrHrxxmvRMm0Yt4SXWO1g9L3t8
jvE/8EEXr7wnbRHgJdrK/fX7MdX7M0nUDsFtfkXwj9aRfon8/c6R9H1affa0dgSmHOQVvN1WSscn
x4eHdtnqOO3EJi4+0iOyiee3MR1YTTtVbUTPcOoGiGfpmJT3dHlNBBHdElyeH4VO3BTZs4vqHyK0
fLobWT+CDamY/ZrC6yfRT79+uPutOwopZlXS9tTjgI+i+IQi42xeTV5VVMFLUJumxEdqVsZjwPNm
A7qgSnBkcw9CkH5dt8EyFhvSFRN1ngQZjRYCvjCdbfWZCeGQhdBoo4Y7d0PCmwS9vtSnCmwdz+KI
yLG5XJx5Eu1hJhrhxIU3snToZRNEe0tDccZh7A04R9IApB1mZH0xbinDUDPAvsRxPV7Z2KRLZhJU
oJkjrq39c9iCCEY21lgYVBKkbH1RGOfgepi4vLWIE2/6w8OgPqM/DWKhyQDvwMMZ68/7nigWR4Te
ZDS/HxEZtPWNYAToqa9Cml2EstTEL4MGIBbTxDaaB7Uzt52oc6lH70CIZbqabbpLxIDIC14YM1SQ
qjgT1bsNTq9D+1T/cwlkFX5bBtzTuQfEnX+Za3TstO4GLZlg8YrAcH0T+yw0c1oMxMnNIfbb+Yj8
fDFQo3l0spS0zsVlI0RCOA4GJXVBvsc0LmCr87d7jYJOXZFeRQpK19TePCCGAsTnx4eHhgdfY39W
l016T3g17SfLnowNRhT307fdpiH9ToPN8dYC8IlOEqvCWUo7a3KUWEFHuiywUp/HfRJiarcAhvQW
QIialjKKbkViHFILwzZ4giMpchK4kGgDkQpKC3r/lwP43s9rgxSc5i4JhH+fmfRLnXY3MExrYrtN
hRp1MOekEkjKwV/7QA+I2h0hCcWF/HO5+2BbEJXcFbOdRTtJBN+h+Znapi3pg9pTwRYOkcH2XBZr
wTLbmg8SrP0pITFxPXiKZ4dkWxVEURnPzOnMVssmVFbLsstXuhZptvPFSLpS5GW3jVZodTvIkaAp
5GHmku7dGhOzNpAMRYxWxtBw/q5AMV9HacaSlJBrm6y/a0J5vruq/BvBcmV25OCZx4N/8aWiqXre
WEIalmUbeJc810XSpN7A8OYB04/667FvgMhtCg9qcZvtuoDpIFdhgHLZWXqQ1t/rJBI2Fhcrd0+O
61r6Ij5wYrPRV/x1AIypEkQRBz4xH3/feba9LRqO2RKeQfCcyBEKfvPVsVF0KTL/jN2oHko44yRv
ay6sWbjPDI2xjJ1BhrYZO08nKb5inu5A+QjG2GNN5y1XrRCsPFyTp3UQomxvLoXTo5AkX36GbvqF
PEgrsDMZed9QQ9vMd4Mxl1H8bB6y8p+4Q7nk70EEH8pDGfT2h5W7cvQQTsIT3++VfxpmLaeEqZJl
x31cH8K3jPQtoYmsVeSoE0T4Anxu7WW47fnwDKRpZYzSfWiYaERWjDbLZTjddbhaftqaNTMjviXy
VS1lDHn/e2t0KQJ/a9RNGcFICnPLRj40Mw4gJS7Ti4jMJNDybGYu9vpr4voX3iRDBW4yAdwosdYm
ZsuW9bZ8SSYyeOrFEGUroErIdn8moyT/Gxr12oJIRdsgVEWBPCajK/tC8AmrmDiIMTG+6EVnLY5Z
KD/bUvuhnk1uz88wWcLR526I0vdexnV88vpeQbSQvlZx4IYDmUn54UzpV2JDH4ijWLoq86mtLs5v
a7+P6ruKbu5PNsblYz/u96R5u6PdKNNQhplFo11lF/pn8KR/V06Piy4vEMdKbw9AdRwyZ97fQKiy
Sq0NxsswI9nrqFqwIxreihn0bfobGBN9YAZapG/Bgryg24yxm0FX++7X6Naf2KQMLJM5Skgvl5eE
nKROw2f0IH8v2WtTbyXZr/BGClldbqdGKqO7kFe+6MgZ8/+GjvsBTff8MDKUduv3BiU3akHr5yXX
T/rpt+d69LSkEyOms8UJSW+FYJjFE2isGjtHaqQKgYDTEULjvfAm0IhVSEEbsKyplIuPRC/z/X4M
AG6jx5V1QOd0694lYgVB9Lq3AurKNOOgfjLtWOO720681LsVEw1HKL1lBsBn2euho4q2G5MFFJYw
BRzXj5o6+cOwoCqF2I1M7n7DuvZ91bhsYekMtUuNexU7DMG74iwYA46h9EQYUwSq3sctaJG1hxNo
qiq6Cv7E2SFUx4vd972q5e5SX3XcGnkvkpaS5rTsvJ7jjIiV9Z21EK+MYWo4+Pz2iQ4vqPHtlBwd
8Oji0LVZssNrpd225VUXPaMKLr5VhA4EuP1HFIseick3ltVLA08/aB8MzbHMUOMsCA8RUtol+bgw
j94M1fRxppCmieZHe8XK6fosXK6LIPnqSWINVH/XUsdBXjlNtCt7GKJzW14q3KLjNO2VQ849RbBt
kqILGTUh24uNOE/lKDJw9s1MiEfbJLk9arJSh4rZFEKcpIFL2eiaKWa2osSDuDtMsyEL4XPd5VLR
nlSrrA6qQ4gryqPt4IvzO4rUU7X/dwItACwtPyPA5gtkPg0nk9jZmmqYg45i8282dmpygefU0+MB
5e/ogSjHfmU9ugGUQCjDFRab2DK4QxLhSQoELdhH5BeqCIOifBxS1nzcckX//X45XX7RYktETzBo
jfPvb7wDNDc9V2EPQEGwEvWRnGGLDOX6ptaZ0SYuxyrnuuEh9a4ME5lNMMVBQ2SrqBzSHvXiw9yL
BNemmR2ll7QUVWtHUk8iDNxqvouk8BXaR3h9zJSCEI/VHF1/LY8D0s/LEJbIShbZDxmJobx9xZTC
XTvri/4YXXzfJHRjtX2TMXpdv+BfW0nMElnUf7F201/Nh+lwxH+WhRRuWDZthPHsSeIJRrah7R5S
aHPg0UMa8Js0DlaTps86XXbK9HJxo+cjXRymKVr/Rhcuc/zlUfwYuoNiFmpKvpGftcwqUiKxuNOM
VU94GGhtFWsadjPfdqDzdSw9ApmlHru2hPNz6n3BKGfU8wrgKeNKUoV/WgYtLz3GQvgGRLBTKwnm
l1BaU9gsYfnhO+14JMmI0os9/LkIBYGqiEGs89SLfGGB6KnVAZOEMxwEMbJjASL4EnEovW0tuu/U
l/l0H/LssAzD42r9ekHQHBBf+z5VqsE4DR+dfFPdo6rw3XT+AFMCDOjvKsY4tUx+x/jzFLTPFpff
NSdq6+V2SCOGlWLfmPBL+tJfiYJQAVC6QWb85388kAweBmwq5n8o5TQ9WvTgOcLAmIbxHvjgySRn
IEPV20EHavFEYNsmKX7mYSrGdNBKORN7YbPRpsnzSKQpBnM7SxoiXsEkwRl+6e2+SojyTgrFWv4/
XfYqXFATJZrM6cB1V0eYu/RN4Z4Da2wsckzHcCpl7QYIRHg9kzIZ42KRCqXJ2QFLYElqaH2QFetL
1WY8uu4qHycfgyFIpMouSOBS1Was+xbzbbrgvEEwYRo8qJa8DlfzN3S8nSON63pcA7PGbM4lElZB
txavPFl1lRkNz5X4M3ihG9ZyNHQOP8utMNM4DTop1qPG397uCQ9hxvvakp39hxWklViAZpqEPWyK
/o1aYVt0FY2RY2zk6L/OCNYnkAxJzAGRAsYsl8R69JSBGcUMaSHh1FYBOZwdjOjbu9U1K4A1v9MY
sq4n9zBi/0UcIX65Z1rOOcNpB05RfkGFHn+BBUFSefpz8OrWVihac2IUdTZywy2+VEpAdjsFOk1e
4mqrbrxy+UdjCsSN6hyQ6FIAKJVo9+JVwyyuOQs5RLwTvjaLI/jX+LiVQLtzG6f+XtGhiLBUrIbm
wVaMAcrqQIHUeab2opU3bNXbDfAARGekqap+7Ax/gre48fAmfatNYPFPyUnb4/3ZF9AT+WiJOsfh
fKGgKVf7tOid1XIIZk6bEf+kD5OvkMxsbJz1cFmywuUaIi9frhkwcuSBW27rlnk25l2xh0evObpc
/q393uUdCFACfGIFjN7pUXKWChseE0DY6/IIcuVA+2Qlh9h5IhjZqTzgLRplJGJVIWHAtjOTNjKP
DoxiK9uNXs8Konfi6VcfBOUuHLe26Io1N0PZ6J1o9BuKMxa3Wp4kFq9rtlh24kfurZ5sCXMywvc8
YZShyAZk1KEQIv7znGuMHqgvPfSZKaGHkKu4qYzhkd8wzsAYCq1vbuMMRbC5zRbAgBa6cNi/41uo
8fcGZnV63zG1Xd1TBkHeZMTcM8rhWMaeo3K9ZDj50/hJ39QZnTzXnIxMnWqR7zUSdNvTEiewJwTi
a8Cw6CV1R/woQUHKq46L7DzXl786FzKRMuoX/WtXovTynEEVpKv87W3AK4odibt9tmNUa6JeXubm
/4hFxJLybBrlqBJPqQRxIlw8eZHWQHUqy/AXDZ2Qpi0tjCRqJi29gPtR+83vw+TQJpB0bbbIUGmv
ys1fyeM27C/vGRpkDoMDhfo1Tl2PtH/zvunVpCZ/8oMqhmJ1bM06nt1prgImZsQuiMo+MmHZwrPo
5nXFMg3iRSwHwD/X0INENZqurETAhGgxyawGQKL7jmRk+00n2h+pYD5JvpOpb2mWtagtcpJ66Dku
tjbYmG/UKoHGQAkFwpneaR2XZMsKLsgzWuIH7IU8+29TlO6ovZPZlv+crDKAblT7Z4gLptT4Flwj
SB9qEBqgRBRVUDOOhVH5T19JAORen0Hm1ZCahPx7GCiGRVW2faJIRg4HCv1s1lcX301ALvyoE/6D
/pKn8YVRHLIEhU0UQmNUbIFWD1xI+Etr2veEtmJyR39hgQPizWHIyvHE/fuo7oSsF+kX0GCCuB75
wvSD45DqwSPRy4okPRtSMMcBp8JPkwltoESuICIRvQV4uwmfwoutM+pbkmwEOAiLULV0b8eYAUGV
ViLH3atLun5VavT0OZaSHRIGRC7MLFVJkoSFQMmka6nZrD7rb6soUNOPuqaKf/w+Eb+UkW2j0n2E
IvlNoB9ztjBPJS9i8Ps6YkDNIfN5g8pNhm3oOKKUL6P6HhXPeGYHW+w0BWp3xRkM5YHzBh0Ag4bR
8L6JBnJBN5+pbsjnh3GVRfpcu66qnJUIH2WxQJsMEPF7T0K+nmaFRp83ZnwzdXuTzzJFlj8ytST1
HBI0KSIEjIUAkeB6mNA68I7uboR6jzsArYqwCLquGZpqr8FyWbdmoye01NgUveg9+GKb53U/eCJs
z+FAUvNyxpZ1rniRI+kmODKTnjg/7EQABgBvdxHN2Y+P8x8EL9smyXkxbpDfFjXrJCDXsPYxGlRW
vSN/548YrpgBoiQmg7NbK969MPrMLkjkqSrl8KwbLBPtIieSc0FPpOeLDxGQC3a+bzoR9yGLMea4
iaxB5DaDPqbrZjT4A7SPuz8qapniXTwLjZVvQcs0EJtvD0NzIXj2xNV9JUusFJjApG9ughQNFrwU
eokVcP2o7PAKfqGkRyCbd2dZ8jQzM7bhGnMW/unLi5vTzki6vPqBz+gVe0BIj3LydKWxsZBRN0uk
mpo9k5NviHu3Pn4Yq63yKAeDppFp4c4tQbyoB2xd43B9b4nyb5h+btysKiiXjbV8hQKFqqkmriS+
Jco8E0ErmhxBalbEr8E/TF9EfjmZUOETV01syBkr1NHZC8lE2ip7y+h5rTgrvQtUp13h4x9Y+JcI
E5PoHqb4nMxqOCAOoZWkD1oA39JeVKIyuQeBl4Vqgvsk5QdFtVbnvulowht1dgzolJr4chWxTjEe
+zbAma29o6e9ODJXU97uo7k64dLHXVuHgyvP0cjBTadsEvAPN7ZTVhRfoHamLXIfdV+U0/h/Sj3T
v9VXE1wunkqgDjnORwQZzARuHQfM69tOKApw4P2N/wmaowh3KmVQo+LlMG4EUZlh4PrTPULNGdPS
QT2kKA/o/b4YcHqzUl28UxK+Mn4uqJpM99/6+P6hMWL9tMkdbaxfN06hAGK2U+vjmvAKh2A0b3Vz
aZR7pxdUaI9+YYECb8Uy6L4AEhWaU1zgDmQX60wCKyWmOSwqVYIhYbdZbqVCLYWq9HTYPLOmM09h
re+9CP+MkcZPqPiVgQ2BPh5NRVR62j5ax84w6KBIc9T7t7+ggvAj0Pk8W9Dccz8r3BYLqfvrKPSN
jfLUrDakPMhGKzxdQqtr2AOJs9zWaALa4B+NTAtoBBAjpnMNeDVK+wSGIMEaWG3nybmX+r3D6nh6
tLlEVbIbn7BVQRvfcx0DncDom+uLR86Mz+HrBHF76BEDCBH+N9KnLIWzapeogyqgdvvhd6hvHKl0
VK8CmH4FwTfi6amykfrkCeHJSJUXq/zUAa8Ast4DnpeAQWFn5k+dfrRSPyPNetS52P82bPXhM8M/
lbOrZjSXq4WzGIS/TZ67JfrwIhxp0T1b6IwgEzasAg8+amaUOhlfL+EmityI0BlxVvpexezwmSPX
CrWx0QvL4Gn3t09PZm6Pr2sgVHswUpHlsoAIA1qEgnxHZsoUYWoeisDDfBBmLmOmUuXMXDwXQEub
B1mESAV1ntewDAFXIK9ctZoWWPaK4OqeoYgqYy8SA+8klByFG1HXV8Id20rFnCvbh61guc0omXOz
guhXL2MRDQfVuZh1MUH7nuFA8J4o5DC4IA72OSU0Jsawd0LcnXmC74EGwCUVXiHMajlTxMLZQmMW
GnJPquIR/IyzJ7bKI3jnWU0bROUpHHZvHS2L1sfWeUd1cPK2RcP7FECGICqlylkeT/o/YbCQDXTv
mIWCqNTTzpoDW78sMe2Xkzz8HOrMAgHf3tkUjLe/4rfiJIXUIC+QaADM78vAOGNCAzJHtrgBtZpe
l7/1O9kUDt35irHaAKfCessQ3dvAt+Nuu6RjIJoPjhTN2MVGgthDu3cj9YoVmP9KsbgPm8RlCsqM
7JcVMfJrZc88OnAY3BYVjPVmX18NqjpoXmx8LwaLnqPjOnjQZWKoeeIziHdEcgLCdiBLtTzuyImd
DhusG5zXOohLOd1JdYX846gjHG6tA7087H91saRoMcnKD6xT8qhIFyRL4Y+bdx5qyKBZgmHWQT8S
4ee+cnp8wIQUz2GkWZT/y6qoEAKn/+4JMGv3YQEsVVxlqX8IqSq60WguTngBRzSHHWy9GxHONTHI
f8CoDikyjub7hy03vOGqX+Cs5a3LUDq6fSqb/ONp19jB50gsWRhSK6s60cPbquX10cZB5/8rxNjd
0IVO0TxO+ouV+Jy36nqAZWL6fsnDXxB0WZBbP+sK4Yd5XTKxcH3kyhF5HqwZByB9rjGpB4g7swQD
/DAmzjQrrtDYEoMjYfwDcwPZ5y32FeBIGI/BG3oWX1Bge/r6H/xqBjT6tVey/W8D46wcDHh9LJT7
yE/ZB8kC76iTwXw/6ivQWGjRVaOEnYV7zsgGgreCfVgCIhzfCi7BPpgrKPln/uAFH5BgqpS8H81x
U1FkFblQ8Quwrq7uhvyBMcHw172mk0XDju4eztaObS0vHowKID3TjIyTxELARXWyo04RocdrkPEz
LFHsVvRW5Zl1tQg60Pe1lcpvJliLh9APPZb9lLkMUWyOe3/c/pLn1GlxOU0OnCzXiSbhvJYVRzNH
Y3G/sKlp7dsrZqlWWre9HBoVtiYNy/qKP0+OvufYpD1FimVaYe6WzmGKQmoxcPpbdrBPUbTBCRsK
DqzFdweAjuxoLl1fy6GUhx+rK21SZnnlvVyWIqigWPSVp3e8Mwu0NlQ2opURtIH0MvelWIdN/gTz
iuHNeuCVwDHshJhqLmYU5TNCw6zlhi+Uu9TGZzNvHusuo/NnRq6bJWc/VEbQBFmCrSM5ow7CRH6U
y+oqgsmZcW3sucqbmnuQnKTwztZQ0x3LoD72LVEx1ZcM845E4GcGcZgi2D7uN4HUsd7yxgAjXjjV
+myv+oVwiEx9KvxNWSvziT1Cui1XwMJjMlDHDJ9nzlvzoxn6RtuTDWzoe9QJ68lzAvyT0itEIjtU
jMzWSptx9QHHheABSMlJPtr24rQ1q3lP4JGxfExgrBhIazQyKKEfYOPSnjM5DFH4mDOmY/qB/TLy
A3GxM6rpYg+en2PXr2mFSZ7cT6l10vlwHx/RuCTGHWpgQAHOkVfGExDUJxEEhSaK3NiHVEd9K7wT
0QiS7Z8tyxNdjJKeJ3QdIu0GuBCTs+OEAmaL214wzgCOzfeU3GLiQ6NNfrKVdwaTFSvn+yMiQgjQ
50Ftwos6BwxwO9W/MQGH4Vv0QZTOF/cYE4oquo9Vl8GccBQuXc0D6PjEr/apW5WNxCTC1X8KbQCG
BhjGUkpUr8H93o7OfufosrIdsp0RyyolLfrZToP3lxszCwy21vrvxo9XuBccqoe9pbWZ84fGDjet
zE0i0zaQGoddD25sM3fOGJmcC8fqyykeRo7YcZ5yyWnlImmE+O7w1+NZiSAKTOMfIi1Hi8K/WA84
77HuofKRQGkvg7KtWZJXtt3/4OSYI02KhSCAQlcYkijWDCW9KtqSg0NziiBxndFsIYnzUUsvZ/ys
QTt2sadGQh40II4g02Qna7muvovNOK8G2H8G/BP3A6GyzUnFQUiYVAS4oCXrqvFP46Mi6V6Nxk/i
JrQ4qVfwTUi1L0my6rIah4yM6BD5mHPXqekU9Ibtej1OCd9Nkak9NZo9NwSC+j1yvQHW+b7eudUa
oV0/1Vf3otdTVyV9zVjTwNPHA2RfFNSFCdL+LSwalH0mDSU6yRKQCm7mhjwWFanh9YQi4c0vtasB
/vOPnzvafpzzujjRAx6mRELLcexkTUxxpkdcyuSolCV0GP5My/2aoVAFageQf67iIp5yWgdI4E+m
mFcMxQxIwJZPmDjqXeUqRV+We374lgEXgodXPzfY6OUOI7TI7xNe8mKYGlhJoTvUhiXFv0b2NXCH
qH/mlhe3eTQ5CYmmWumaMXwUAdmgMKf0V6cq5UloFq2rrnYJYusJgg1/oWL5bYo4zCNUsQGuTuJm
rPCA+xjYKSHTDsUUYO4L3bIdbdkBaKDTdYjRtN4rOvgmLNy7GDbRP3cqd2f1p7SIeZx/2+dOuwSC
8gMLkwHriRTP+uJNLZH8LO8sOm5gAZAiQEGuv8GYStaI6dmGzrthOf1UTq5p6IRHJHCPOKkgOluo
kuYaRMm/rlj2dvhUEqDfCn6UN+jEL7JW7KHqQ22vEauOuOthVVA8CI74KJomuz0tk/+vAC74jqLn
mBfYcPx4F65YFXOPiJeSRUwVOf+kPp32NFBBwKk3yl9u0v+zAeA6nhBKlHZJrBdkiF1Ti/KHVOLL
BvVxKUq9JVxvlwLuVuhavbraDRTpCATbg3a0rPuareF+Y0rBWucqBjoyKZd8X7FHQx3nSypWg58E
rl/lRp33mHwIRtMGiYFJI1oaYQO2EyLl+w5+Lg3xZpjXpjEcTTKohGQJfB3z2+R5IrFLPBD6bM0s
YosD0GHuxmFbVMqBOdfMzjS/iHFlEHtmPt0xQ+c7ZbjjEj5WOZhx0+i070NLSa0WmQTKWv5HDOeO
wiHKyyQlSjRnxBPI2eaWZB5cSTQ0OURSWlLuC4KAZ2fVHwnvNLX6xO7QcVpzxTC1nO7v2MR88Kyn
s79/YZhKIfGpisAnitTPzYHEwvgrnxFfIlxrSH7un0JEoTjz6iZpJ6lTNtDkD3znnRSoaA0+aA3z
bPve8a/ceNgX4DXUgHYnasVnO9SqxsK525Oyyn5lWnrKM2k2e4Z7F+OG6JUDuNVSrh72JUOqRjOz
kBfRdD6MgXXHzBe5STgiOSNZNYwDQ9rRQqRqcg2vDRH2sLNyQojUhuPhiMF3XMZ3hQqDtyPFdQxm
vkfpE5gYoznSlgEbjhWOs4Id+cAlFKpXicmBUgUGaT6noUwDq9GtRbSlBdhlB75IuuNk/RKQdJ29
3HKuottOJDutFX09jbEdj2DnPmj26UV1BCeP7HfH0HDXyntEv1oCyDpcOXevWoAx+gzJjmDcbdlx
ecOaBResqzZiFD4A3rz8c9MiY06HWUnPMY/Gfxxe7ac4uIV9I/3UME7OeJAA2oJkLo8s7Sy+Kh95
NV/BvNRM0JovUzGaxbppblem9LxY/AMjHaXC/JJYh5nJBBfkoOLZyjYDnFyI3YbsRnA1fHA0KrX7
8qHrnysZRCC3tSpk7HkclFWKKk65E1TwD3NhAP3grZGBJSkZQeBcuw6Dezp4KHDXjEc+gIl1WwzD
ZHdEPAWL18XtnkFSjuupHj4m9UnTpysDL252xDNa6EFwwqf/uZ4Fd6hiMjNHAU10ZUG6vnvIvSvV
FHGp9ld+npJv9UZfwHbEV0fNVc7PgWfMSG+xzo3G7XNA6QGI5t2jDEY3BL/qs0HeVI+Q2/ce+CSu
o0W5s6aUG/LyCHsr2vdmUKFzahdLz4M6weCdFJTtNGZEjXDFnHCrKdGTIsUBgCsUO7GdkaQJYiN2
DhHKsamaIfRaZPh/sxGEeu8FTNMuOs/DJXQIyexB4h7VoqqoQZxHvqeOPCdF806XQRmFJapZdhd6
GKTMVKTAKj/p1182wzxMVt0VaOyjB0Tyd8Ht1giFwfY7N5xI4ecGnRhU+KKNR1XstqDXkL1qOtnB
xwJLPZpw/YrPVSM/jrL1Lhoun+K354MpLMqhcZmQQinhKoTiQZoKTpYlTURqmzj1rPx4NA5RN+Lt
yaWAp6T8dg01kP9sBFNI70BIN0KRDxWTmbat/6CETo9zKNVxxyqId71Ui6JinlDUMB2XNQdMv+QS
89DKNwqQkneC1qnROatJb/Ny+QOq+lLL/3q2HhXYPeQGiOVxb4hLOg9De6X5cW29Vyz2LP+SJB6g
6weR1+6qHuP6SiO7BR/y7pa6BSBeB3mChSAkip9fUfpFmQBqjgOOCyiexy2e8d6r0TRLKnqirL9N
Y52WHi7FlmN+C37eFriDiOQJf5LK/QLWMYEWSQgbyov4fFM+hAkF6STx9aBaJq20nv7qTbe4Q9Zo
4+AOY4sDRDOseE6pEHqO0t4Z4r/z5hTAJxv1EFw8Q8q6D9rYpbFbMTir6NzM8W48TsK5VdiNKavP
CSPNjD/F/NdjynnS9HVVTedeXXSAo7nSZvoL8b707TBSdJcRP7FkZDW8Hf8aP635jrFFQf58dz6I
C0tNLVAlI8WtREyQeY7xNVMqfP2gXSN7h4uJqJJrFehjhINCUssak4THBir8mAKv2C30Psq+LHbW
pwuwXnsmDhRlm+yyridkInvYfBsb2TgwvRq9s/oxS9yltLRN5D7t69/c1jILCv59kP166rSf6HlC
QNt6sqCeF/iNtBtjceBf8iRgyexYfHdu0gNKzP1qovuAXtdcRigKV0Gx2YAGPdJxui66a2TJwFvE
nlSrHMghusxtCVefETPD58Qu+j9wm/HCnVFYGgFNKJMasfaILaFJN0uQ4TS3GSaTyPACTJ4efSBu
trytzsPTwQq/98oLuB97q8BxI39i1Jpb4rCJhwIO11LSfB2kBJxf/IK3MsXWXW5pc9snWmMV8vl1
kkxcFyG1291fIUpXCz11YCTwEAqu80ww204nhcGMtvCu8eo+vbtliEA1Oy0ZKttp75U/n7bICSaq
4jdpGlP4L2LgCr991p/jHYYOs7Nh4xyD2rhMBGgpuCycBSb3zcWBXFejvn4pjtRfG/nV50qOTiF/
irwgXqxLZgapwWJz9hWAQi5lJ4f3J2Mgf5F9wn0Z/qbDODXtd/pOwcmsT+9Tye3vCk05Edqg+SFJ
vyeekcLZ2alfHAxDuh1Xr9siY/dd7MDnVyTWzwDoGWjWGOkINKVHLCunv2aeHbb1KmEuXn4wu7DF
IbdsGfPlcIpRa4/duqxYx/zP67vgPQqGjjOGDi5PAf6OAf6da+5AzQQPFywRmPvIsBzNDEFPYnRb
DB97CkJnVk3VOG1pjetmXMikJwZ7x6Z5MrDMWWwRGoFa5UtGU4kpr3sDNUVkQQc4tX7C1qu/JBWt
S+bRut16pvyYltOcp/cL4iYgucJ1jid8gdWec1hCVms93d2OuKVAbZDN00/vswTR//exEV6qkdAC
60ZzuTWHKmQORYB1nF2ico5aa1sSwvsN5HUO625DjE8PKHnBrpG3LIlQ4euN9m86xv6lUOg/rsg1
fofvm9xLCIcPjVuSNguhtNvM4UOueaZI9c7yI3ukhso5gMTXim21d3D387oU5+Esfu5qVPC8qfY6
2azguK9xFJeZQMfsnL0Q5h/Lei3lQgYHaXH7ZP2VZmSjgEDUpToXTrvlphC7mi9LQ4ZlRohh+sd2
3+3jgn6rYo6y6nzjNln0dkqYZZSOWF0voi5k06XvRq7752OJ6M+hNvIo06XzfFnWkCiGohUjpO4r
PtScOdHkfA6/VcqA+JDB4VYM97ygE+kCNEaTzuAt3Pb8NCtTVcaNQNEwFU2TSfUgHKWMJFZLmAqX
OcrsCVIlUKEnr2hIprp+6zDD5/RtWSSl0eTO2dad5Qor+ld1NczxiiDDWD0xdlyLeEyaBuxxX9ND
IfC9/o3GluRHp2ZOukqAW5u9RxV8ufgYJqrMuVDTw931WC0olNGrdGNLKJ6/8NbS4in6PCQIp7oE
ZkbBCrDLnaPle/lKZYt0pAshrEmirWjra/GKxLrmxyTHHZ3D+yXXJ1eofY3QoFbqStcMG2qMZpgv
/yi3ZYdE4jTZVroSY+OiqX6R+m3o9pznpdQGSknjJ0FE3W0fopPDJdazZePgaDXWdVM/R4VS5O4X
rJPfd+MofCSbjgLoEc1QglIdy5rbkQUWl0qXHHERy69r4cgE4ojRgzMzzw62kLokm5tVrcDWvsiT
K5NkMSBxj8ngAvhdTWqGZUcq+9jnlz1KBsbtGqKtC9TIDE3PlsCrDi5JOQusZJRNikSim9pjjLHM
fTBJeL9o+S2mODgTNc5ut7kC6zI08p+aY4eXHNVrSgbSW5IBxxBeUDU5E0d1nRCtsX0CVCNn9Zfw
CLZjxshbzbMTQTrIgqXndpRz53ZXxGxpC/PbChA1/z0C8t1tm4wf2M/p1E1ux0Ypq+YV7yEgVtcn
2tsTPX5HsQcDO6KpKnCoRRJONhS4sUA5HFa+Oyhz78f4qPSyrqlb3goa2R8ipX9XZiy/kl+iZzzm
1AESD6ap6vutEHNmGb0/XGwAUK/+mp/tq2MKWHGFH+3oQnZlkZLVk6wBpfg8rVWXKAg1ctVIbGJx
vDx6J+wmHghhZmdLgTmoj1WDLQhZwNGb8k5VoBzmEkk3tqqh+QFbeVJRSgRTwjpqoo2qsnpqNNiF
J2S67tRePrzCQXuqT7wV/nGs64qZlwfnKUyZheZd7fBqhVRwU5dJQ3uWpP6en0X4dfgNjzZK4MVf
sIR4uQqlQ2nhyM2X038X0anUlkli7PTlI9YUdhx/gGna1Vgvasr5A0HUWPn8RcbJmvld+A1Nnnmz
r8sVO1QV3dJCXqT9AbKWwBC9hfRdd/MxGdD2htk0lRXOpNdacbyX8XXzmiv2VVpe0fNos5rT3BS8
gxgNjew9i8v/C3ZjCmctI4PvfE+1Ty+D7/l/VHws2dC8MoApCjCCn2wcvEZZs/fIo/95Ye63OLK7
kXtZSpXHJSYi3JAdRyCSMDb7CONNb9t7gCdv+EBEUFciP8P9kbjfmRWNyCPhXqBWQhIn39+yA9QC
fK9TW1k2n+pdqg977QwKneDxrJgtSvxgRCQbPzcbGO0ElqyeVPcn/8qgICDCZAmAkzTigp4ThLuv
quys6eJfVq+fFUD9lOQ3qaYFTg7XJx/DQ7HB6pXgeqqKPKOkGWW5zse0rMZvIYHMI6hdtlfYAn29
kkA0y5hOZZ8eij5zxZXMkCksF5ES+WWoJL8jKQwv0qEotB4XzX+FuLOfcDZv/+mimQ7POamOZmCe
p7paTCUhNs7QSLCMTKDfE5qcGSbv0hbPzXJMSTlRvRAjSfcSI8M+5U7vWxGEZS0cDWZU6mxG8fRk
mJ/nSWkYGLiB98ovZoFBUIiOUHO0lrFCw93Kt3BK7I234c2z3Q7VqprazvV3x9SqMFMFzvLNksm/
Bi6xiu9kD9qz9Z/WQ1pjd7YGgFi74lVAShvQJznl3zR9MhxrwIm3J6yUsVwSjIT/CvVPHZWrbRVI
SyipDbANqYOrSVl+59HwwgQFNN6pP2nI1sDjfOSsYnT8pop9lxSR4vf2Sd5facVsybap6GYpnsXA
ZQQfqx6mAyYnfLDN4FLju43x3KHziCcFqWskJIvaQITz37/FEmlPVRFuI/kRzidhwtbtuksqh8bE
5q9FD80XXiUuBnYwXpJ/x6UmxIh0IIlXCD7xz0WosmvvGHDUvH5IU0O8rKdzZjMQzMY6rJWx9Ykg
Wjk342NmNEMC6F9IyTTEGcBRbr3/8CgjYSsYi49aF91Oik0GbzlBUtn43kbRRrGE5CK2mbqqq+qY
NSLeopGup5y3+IA9ZHu9VGkKi5hAtVIY6ZBRIwMUcsTxKma+xJVv2IF8Hnf7ckoOj2c2BLkos6ri
vffGS15GMpQPZgSF9eMoXUv2JiownIRe2rg+rDQUkugaCjQe2XJ4xNZ2P65GHcKLSU6+cTBNIH0V
T44CPrW7RAqzoZYXHgKPJnmJ3sXRKxgEh+MPBW+QEwxELxCYSMNpWh3+pDB5e04Yg9Kxtvkz71GA
/RU9DVY0eVTk3nvbVdNeJu4xbABOnNfz9BxtqMwD7HN642YJNuIrhO/kl/TN4FoNC5bfh1zloXwR
/uhs/IVyuo7ec6Oz6KJ/FuemYbc9oN52fUh/KkK6/VLgTvLBAUJR2Evit5cKYWucwXgU8Hwv4ll5
joHA8iWyDA/+wM8dhhHHNYA+2hnZwSS8tzURgRAQuPQ/ND7mkoFGltm4tPpYVGO6Zf1J/o8l5NXu
Ash/hiZaBR4iHLSovYNiFYRYn66beu0aU+THUaN2/bB3KPcQQ8QFUSyx9xPwQgmGMlQ2mW9XWUAJ
n+SLNDbSdid6R92qDHgaFwyCckAVhyfy6oPpvvTzmJiUHUUZANISy4p4XHX3W/R/0jrxVpd0AcDi
4kRpZsTKYIK9avys4T3Y+sMSkFjzj76P0p8wK1h3QjRWAJvLjZjhGvzIB7G/oGOcV0FZTLIQPFEy
kH5D0uu5lnPbpPDiC2hQUkCZU6xMb/Y3KH9/0jr0LzfIBwQSFnJSGnJaYzNOrgDtpbWBWbYXFVeC
JB6DTWJV5YoZz038QeI3jd5zDy4fknccId21+o6w2qmZp8uHxLAr/e0EPTnfhUpufZMgdIDMWKY/
mkKhK14BJ/rBgXqSlBvDBv4Z60vi03i7CB0ZMBx7Zgr/u9iem/af+kEwVW+VzX7yAh/46pMtqv38
8zEs5jyu15hvByODquZ6Sy0wXoyilVpL0qd1tpJLEPEZV/oLPmf+gARCvl1Hw9qIWLe5EA/92UFj
zZa37gizNw20DQS0rjkTgUOkZIAU3sugxmScZgCjINn3bTxYDTfhuBwOyzakduvRLTo/e0GN6hbp
cPaZS7ZnR0MJRAN1up/93npbvNFjO7ui2411X8+9qC3NBSQeo6adV1RVuafj1YoqBblfk4V7iAM8
QOy5cmfh6wMylvBfJ26Ur9t0xq6oerzqMblFAOD5zcOu06LalHipF6kFFtWgrHMeO1fz9ub7hD98
Miv+TlUq/IUpDi9EgcuC4ElvOm4vzQK1KaywGzHdmNQuRqzSxtKQfG9JUx58TFQb5hXgEngr/kEe
NacG42u4Vd0U81ESeXtVf89x1BYTe+lEzw16xWKrjpxSTbgjCOApkhfmTc0IDazW8Hpp/S/bX+r0
puYEjicBms1ylg2v0lvsyPgXqddL4zNhy7PZ1zlZvIPjMUdOshNE5Ipz7EEcQTjLvT+Up+K7Rq1t
FGAtk13VmBvs2JY36XSKTAQeeKCHfE2/OPcURxfs3gwLtQpGEASWQo7c5GqX6E18HzjQsOphWa66
YK437aEWYtY+E7OaQ5RSW0AHg4YU3X50AlhPg7D27k77GWXBH8LRGPOc0h3EfgE6i7OsIkKRk3S6
xESc2cDnE4ZeVEW8R3vTbBvN6HHWlC/DJivCO4b58PT9Qnly3ny/D52fJSNvEk/qdJQqI1Cz199A
pwl8WqjTpSQfjduGSJwsfiFYwDEBA38AaTb8lzUHDCf8lJhdpzswb+qTCBKut1k1LPv/z1A8BQ1x
7N3LWyyut9WXZEhPX6vRUuDcl6BN1TS4gm1Sks9lqWOiMVm0Z5GB78UutL0BzfjwqHMfH37G0x7f
ZqP4eCKfBby0YAY2xPupZuSd2bzhC3YAuy7NKyxW0mSylSEVAIaeKKPtikDGXaxdB7HxmxpRP7pE
sqw9EyeWV2LZSY2K3Op/IyCTffhWVylGiR8wjXA0m3UKvUbPPP65TqbTYtlxKPqD9wBZ7QVEWaP8
w66745n+pkyUQnuSQecdLlM1Pb20/IfEnJHXmk+1aBmPa1tBdDFKqpEWbrE/i14qPR8IQgxj+iXd
f3Vv5+XHYsch72Zr8v19+QKaw/xOaKv3X8QTguFjo5OyGW0Vpi1NEdMSPNK9Y9K/61HFBGavHvOu
M2Rfk835QumedZkc1xX4wFI1CqLE3z8r/j9Bj7BctRklfCFiL1j6l9hfDscFS3FWZ1C37UBnctMG
FMvB1jyIYIQUh6y0StK0d+qfUMtcE/QPWoMENwuZ0mufbxl8263xHloRAAS+2ga7nN1TWSwF51H5
qnO3SZhDGsuPF5T6FL+2yhMZzr3fqEOCirJAtfGFsrY7ljEeOn9Nc5f7YIBpth/ld5mq6fmkuEnX
BWGBUpWr+9MXUUIouumOV1OIhLnZis3XTjqpiyItiknVutlePlM2haRL/TnR+4k688sD7/B4STsh
QjU4wkz009L1a+fc/J7U/xCtHBFVyFuxLtpjBMMoQYy9Nw96Ryasf03aliBTrSsR4Mlo7g2gWEAL
wpcHEh4hC4RLu1wH52lMgeP1R7yA/eZoRZMnIoDZJQkI65KICyXtYZ+ZvJLuz5nW2OcfbvfnMWOw
pdRy9vGKI4A7JRpIFAuaRstb/mH3rdHria/WGLn7kW2pVChLY/zULPP9yTRf9o5trwjRaiXq+Vfk
Tx0c5nNv8tZrb5wOzX7gfmpfrxGn578AQ1Ux9ZmDah4Su3S4WqdT/aAaGoDbKnznJ051CkLifyot
j3Fx9YLIvvymHMX93fxrM0IAfK5Iy4a9jPvXFT3Zlsj8UnWyNETdaTgw7kajeQuJoCDfs4lRUcox
O+9C29yDIq1bgZiZkP0A/6IScreibPbVz8+QIiBpqfBpRs306Zppdt2/6EY7kQy/N9jquJUdYDWm
eJ9mwhpzkdeeTIhL27Hs5R+ZiuaAqaTTwy3WP3hjcOee/oNg7B/jYgRvoG5VASJLAIT270WQG90p
8cfDvVVhzinHCEgZcjJSn82AJEYtk/B+vRJKThDw8Hj7ZwXIMMCqObVBMPzHnfl4BH0zjHjJnXku
IzBUGf+3tDA7CR1p8tBmO2o4hj2g4unZzTS5i11fu95s5Sa8glVD4J9rOPCQlSF/nNDW/s205goh
FqVYZ/xyGakL8OhazT2Tx/DaYEWiA7ojIJh9qM+uLiVCi7RpC/gezcYatAU8T3CoWcfFwpZtfwT6
v/pdesQpCkhVrEN7/P/vnSxCw66k75u5iQTMUAgHRdzogX7qam50BFmSdLJ+AVwjZIFyp5teSPpP
YZL1vqflDbMDWQR9mRZyRA1uvhljOm3CmddIxitC5ld/cY96lgw3pECm/nHW6QbaPkM6qNUkKlGB
ahCla/ygppPPBM3vgDYGXDIduXKghS6Z67EhwQpuPjfFVrzSDzQuiEwHZZr7TJCAU+sSZVEnJRXZ
fCfjXIyQCv9ryj37dxn2QgAsjIlPCcNktMDFDBL9ujQKk1ipTehxkZEo6ifbZEcc7MhxNAJ08w+f
Kq8XqV5+DHlLSaIg7ae0yLYpaSKi+6HMXZrDs+LQiV/SsWeiVCrNzzIe2OVuY4wBjjbTd3rlbHU9
zQqrw4pm0iJioMl6vbDzFVG1/QysdNl7WMMQ30xuHRDCOtc8NO2CDDxxVJHSnGl+qE2uL1aXeWwd
uGUqs6P7sfPV8rFSQceVUVcTvogL0j7D1BEWSi90SBYlyE+oMRIZxDATZ3m9FkfXMtUi+AQkjEJZ
DSz+wXqcg+pfrO8Z6gi5nz+b/Hn4Us90HRqw+Db5cd0GRP0MpEJmNu/i3EU6pKMTVkjSYBm3VnXj
xebyT5U6nrPquQuYRSVuH248CEiRlkLctJ2qLGzNwRAigV7MtaZx6bl81wzkD4/SpK+7VdNmkfCk
/u9WL109NFbo3Fpek3sh1E8sul10w/JHiAVhX1VT9KUnb1uxFXhfjuQy4eMRcGydHI1JUzFVJSAh
mgIIVjdMCXVaNo5ms0FD97QZ59rtDRFI+gfPzcACidzpo70kmBGjslRWo5bvXWJgCED6Xx1HwLBH
9UVQfrwgH2P8KmeKWal4Y2RJWonZb4JGs+Xcl4CxdM/ehcYk6BsD4RvO67BMBMF7NdMhnL2Bzo3H
SzYCWo6nMZi9x9OBGM3ZRSMOxBEsHfOhrDUqlY4Qpg91KFXmfkm5q4202uqZUNQKcXQ991LGijX8
TEfylqSGPhhKQwtm/4CZAY+46flEcP95nDhDzsJNqv5NXqx0QOg1nEvICX0mqmsJcVyFewx7jG4H
Z/K5peaCqyzdly5RDJdhrxiyZrvHYoqbS5Ux8jbCIAtKUyhV70Ir7eEySwUJ1e49e1Vcw04/XY4v
I3lsuGbV/FatDU+Gh3kr/YtELO/Eoeb3lRxfrHehGEZbTI5eVglnU5LF/PcUiAmNVj18UM9UB2mk
BjD9OKyU61qRRSNPfjipPIA78XhfKtaFbwohJLN3BBU2yOu8GjXWVebIcCpMefADQMCnQnDTIVNq
uxuVmgXegYBNhyI0BCohBCzHKT5aeXb8kbWkeNLbfEGtdIN34Nc8D2GG5ximq5w4rNoLadVHDz8x
KLCnKizbmTKWrHVW+up/TQrx3LfBr6WC/ec+YuAZD97g8ab98O9KedOETUJmGdzsMrNnedZUlDkR
Sb0Q1euq1cYlUtoSwcAd+ojKa8yO0gDDnjwXJJrSV1TxLfU+ZGzXQfSuerue5CN7xnNnMrJZvVS9
20W2/4mSYHTUtiZdpyJxbboiu+UCmTldg2nesP2T0g+c3QofLBjUCpz4GM0KzRrw3BZxZntduzNv
5WKtzb0Fx2Y3sHwtcoeUYbFD8BTW4l6j6iOebk9qV4B3prUYnfy4m5c/+erU+k5d3KcxychFdbtX
GLJtQ8U5igrXy2CPt3dLUBTI/dMeUNQU9TJhtWJ0vthZQ8qSaC89fY8R8wfZrfBNr/f7fQ/TRUvb
ZpXMSXg42LP5YXQLLqDYBifaAEvtB+vrYXxYRp3E2olhaOElCZMXBopdHukuwIFQLsjVeTy/+alI
NVXwkvvldrk/Uz88EQWYH9Anac1Wtv+YKrVgfNfxQfPMr4YudHTnEMG2SDhJSOrxUMJzFtJmt7Sv
9vt/qHlnD2akarN1Ehux/ByVgdEl14APjlQ7CKEex1ajo9DyckQW0OOuIGbXFKoMR+JUqNNJsXAa
wyGYHrHLtCbQquGl9ylUxxXCm5VRA/Z7Sg8UM5OhlTn2KE5V4ShwfAPl1Mz/Q7rb0/UlXbcZAd1Q
0z39oajn41L4mnC1eHN0hEs24CZs1g4vua0eGZvxs61Nv0OLrwlvj0rY1iuRDm/YuZCxUn+ObRJa
B7tXgizkYMCOfmJJP6S7GLl0SfyXkQy87RueDQSmzX6xU5h/jN/Xcv93Xn29USb+hkLWPgkFrD6j
j43YSomsDrtjmAxG1NIwFxN6GHw0aVcEBzh7rvtVkxwTeoXNeKHWlOfCr42saiULpZq581swtwF+
b2COzpIsjSv5SU3X1X7zubdfrAItYOYQb0jPjhjJLJai6dvp0cDWc3myYgECwID15yxi0e+qIr1R
Ja9N9O077gmLxJEK+oIyX6djYxHxusG2yU+CpbiMstet0Fau5Xt9ZGRKdSDL4WOzC/VWSiKzIrEK
QmdUihmWKY0AEA1wRKFTPDrjzNyVWa4FloqM7Rhxu64YgPoZDoWhraU/Sa0ZqOigzRvwr26zQ8TP
lwJR9PLkJH75empM7WK/Z7w6bfD5CJOQBPssqMjuGwDY8o5YRAmahhSz+CmGcsgKrRMO1pBo3/5P
EbhrlAQF/uGyS2ei8qsBfIvo9MVogH6DTcVfYJ+Ob6lcsLlkLVvWqE3ItXVgXaZhjuBCLIxkX09M
QzGRRonQdKizcM/VUfA7Ew+ykxJaDHPA8lelt6aCzPmJizPgIQ2oQeNDceh8obgKGKTs7QmBAlSJ
iesIXRZkat77SeyOOvUWNYHPawGGkwKjFv0lpfYdf2v5hu9Fe7WUQ0uqfRCBj6QhqYS5p8OqyRwU
mbnaOM9PtyN+pPJRVNiAh0ZRnyXANgBQjjVLDeMYHCPLzELXlczsCrhAAnH8JEg0WOTqzht17Rr2
Fc7YL4d3pEh2ilVN+XQcqYgbz7v2QC2TjUzO+oBmUrHSQPpAo1BEAYedvd0YhYPiFyGvDJ1McDXO
3IoIxtPsmts2DQDHDBrz5ia56k1siJ3nujfp8AS5cKmofAMEostBwp63INCiJIL8nPYGhzB43f/Y
/pTFSUzpoyBDqjrYtQWuC/QqH5+qDJfrXGP6aZcw8M1EwcKy/vDp39UKes+5OWI04uLDm6NSUTy7
UJqJGKtpcRFSfrbMLM6ara2GuxkwkXOqYmSJ74wKmURab4wHMHXrxFaalGTRWsrMqsqDwZguFYYu
lQW4hL72BJNb2iKaVm0tEypCHNNdEkFgwvPA8JAGOHkPMLTLsXOiW3WY8GW63/2Zv7UwWIrK/eJP
5cQ64VwYsV9lr5rk/quk899esQQ+PTsgGKAbDMiWNtL+KQ5B2mm1RLIV6ex86nu+JeHfTyp8u8WN
r/Zx4n8jmN1iFp1923Ens8D7ecX6WagQID+u50qdepbVGH8Oh5/ZV1cgBsdT0OLq/mGB3La7GJFf
4dkzwthF74eLU83QqNIrwnWthB/W+T8PofejiDn4VqzHKq14XDqXOWDQG0QE1OxD+eXat1xvmXap
wZ1K++WCAmJ9rzMnUT5wHF7DAW8ctIZ4Nl+Gcf2EYrBUXpraxquhhtjigAIM7KN98BZG3D2Hgyo5
n3V887s2Znlv4oUUpLUZhpYcjbAJ9gS/sWZwRTv/lBMXyJn2Hl2Dcmk2pgvujVJEypnZ1eXEhDJP
oBOzsZuV1UGmnoqeCZVO187LGoUFm8bexCv7fyBTW4Io3M5Q019YuEbr2z/GJepkzjtkTlt7dxCs
Cv+0dgKf3uRX0VOGMeWajlpmoz3QMUSRsctnQK69mF7xOiGHr4a3tm0AC2ulGW+EggLqvCdKmeCJ
IsvgGBqNNvCHNaIXzC2bbEbsxRc7FcQzp1Hp6mJfF2e3Wqx2p1c4kXX+/Fi9NiI19oLubode1uns
VWHfG5MBRvFAsbMuyhvoTpoe9WugseCAcTAARsuaUKQcVsRLT4Dqv6OxZ7VgAfz8allMGoWcQ/88
Wkj8L0HGc/xJMF0LT7YnoINsyQQ0hfs9nsUIDpSig2Gv/0sEFhr34G7tpsCZVr/3ISMVlA8BM8gW
eZMAXkPDvx2XYWR76vovTR7zqUjuGEo7XjS4c3MJG/hedavbCgM0AVrtCR0L5ZfBpGyFP0KgZhfs
l1HfibQ6TWXxNGPSOZALhdfzjF4S+L2ephaJxnev0N5+uilOZY8JDQm8FrJ5ZacGfq9L0QSKdphI
NKoUQw5lt7jxYsfbkvmosvr0TNlCyMJluo0/LzM+2+46MFn0bp+d2gw8fJoxc0ysmg0SBRRKrkOS
j8T86icGjcaddb5aIjVFvBr3O1i/B8tcf4QkEHUp/sSPUeiyXt16tSAfIkFIcVbGI7BGo9isBS3e
JbKzawMouVI41AfCObuouNesUQMZD9uM34ND+85JI+GeJR/oK6Tuy3fyXXXz6UZdvvtUyLfRIQuC
svXNntaYCfuX9YnLxQnCP+GigPu+domkcEFEMWyqNJLta3U7V8l9hUQRMqmPWXCeJxSex3QPROOJ
99aG1Ybtgmy6BlPsnkAH7ONb3yw4hXL1TB14A8HZIZCYmsHoOdBISvDuNlF1HAFWB3DlMRP3TkEZ
uwqWXXCGIN+/I/MYeruQQOU16t/gWMzajFVsVjhRHHvGYC9gz65BgaH/hbomQq13qmML4MziA7jR
oDgb16t9M02KJecq42+Dd2z5OzqozOWtl8rmLbM63caXxxgxp79cVnevx83VfGpW73Re4SZKHF2j
l0yPLB+bQVmeTIHu7V7Hno2rXY1AnNJLtL1oo/RQl0yApwg/czecsf0S4WipeqggtdDuq6enW8c2
yY+Z02tjyDgsnGCH+hPzvO022LXCe09W+AIogSB6TATQZ2yNsHK+YA23VW35/QxHFnZG/dmwmKp/
++JuF2p5g/NmyW/d1j99QtDZV4eLBTRgFZhZcxZCAm9NPBCQ0d/dUu6/w9vmgjcQSP2m8L9bbQ6o
Ln5zfpNHXNT0hdZfEF/xtpXPOZo4U4Gy0NYaWnlOSBTNn1Ce77vilPaSMr9VLgvXj6NeivKkmTf4
pxz9f6B+EYuOutIg6RhjQDabEpCD0o5eWtgWdw+aAJQp4iR/UpkIWe3lO+xOLU55magb4r5flhdT
A8NYH2HRyg5P33vWbA+RwJ10exWLtpbp8AJ4QZX0QaZobKN2euxfHEnyx1STvZdPXUtVg+PnQTZY
GPuMQ/oxsux7+/ctDTDCHlei9hobliiS/OCp3cFHrzllkyhbBd/hq6YA+/SeTPQKTEZg6cGN+Qu2
kLpB5Px8RwaiZEJd8QUawnxZf4dPgfaY7com00XARbER2h5V8suFYy/QplWyDp23gQTbbIlRLhtG
HDHUD0HTi+jpBECoRhDiJuMsMe64d1OcN4Zqncpm0PpP130iNcyh9WirnNERab4C/9Pz7x7OLSq7
q+z2Bnu9zW3z4EoUibbsnxLjDsgti+leho2hMdgPdPtiWWzRsTR1XqskQ8Szpdk/IRCuXN9hEyqz
esp4KaYlPq+8R9LqE8PeD4tCGSMQ4qM7PjnkSmFxSZhfP7/l4s/0fO92KjPH5ttcrcw9RwVZYwOH
k0r7YngMnV5fANnj3/1LO+y3kqyrhV/rUcE3dF7SHaIyjs58NFHy55zZ4X3wB9Q8f5xAE9z8P+bw
j/Jb5tenVh/QP4mDlR+RoS4+u2V1Iw588IzsjL0kBuuYKx4IoVuyWHMzmNGyJPBZZiX+J5KT7uAz
vyO0HFrViCdYFppW8UEnEZiRXiM84SvX6e7YZoLwr00E1e9pUa4IDcYeCXa9rQ5p2WONPb8lfu/5
7YzXbjgwDfgthiMzPeQuo5dG+cq8Qoudx5mMF+FF17McHVKWJaVYck3wHZ9GS44C5hw3earmy2Tw
6gva3HFSLVwYaJ28+h9H0YjgVmwyzowDW+Ko01pJJ7xtJHKCtv2tWyRVgLx8Y0UNbKJTibu1+6Ji
q+zHEucOogCOIeOXQW5vzYfeCi/ABCd8xWQkLRxfXbCKzYYgwnIROYcsCY01SWlDH4MzDox91Ncn
cHf8TvL9MnpqnVdq6C0dcGBaIyst0m1J5x3GDwAs7KmSoHWb/sL2GGmiFaSz5bi2A97Uki9T1AAt
VvZme1ZGTilrWZ9J0G9iV7prvQ6pwt1WK90gALfugUWFD0bSDZkYUqzh4FKrCv4Rm2WQQHQRX+JB
77xJ60hxodC4OL/Fer0E47VqB+frjogFZyeYf5o6eU32/QC8oJgXfASRVBESRetFmyUBK1KScTW6
RD5VlOrWs9vi/1nVL8Uv6DHt94S7eAv3qqgEcuemd/h59+qg5sjLDVT4zA6ve7o6xF86st8VZCSb
HCEt5TEi9/YwnNkP5kAF6CDj0ZEdF+qPVY7WuLqa+p9RVDp0z+B2ebueWCP4JSMQGQty6OwlF+49
jyFMcdNbRm/3znENqYgyRF4dTk5XvZfnN7aZwDyKW/IRPkIapUXvMCqsBV8Urx9HcFtUs/dKBYJQ
REB9hRWjOjmIpQztLa2kwMRB384vfUZ0+7TXkxkheRLQxvHNiU97DsT3E9fubny2WgPNPsYOLWHG
bpoy5NHBng6GHhuWxbLCoSGhoHXQrvmtMDiG0MNFvdWrXL0I42dS6g/43nPwBQzhgf6IqM1/qpHq
dkZj5tovkEWWKYvXOo97smH54/0Aai/T0ScVqVBeaN02vMOvVktVvMRwD5dGrpOkNhfj3By5SKyW
Smj9EzS0t5dU6iYjCKSHxb8qqHg7t6OZ/HE9y3SOCA8ajYF54Dg9IG1kUAoTRuPRd50q5uxlduiO
r7XXSl9ovLH8mjukWavbsFfaav+2OQbN5a+YmCVCkdBffrcrpmZL/ctDIxtbM37PDc5PtPSoZ8w3
F0sZt/5COGdndWSDl1o+BeXX6Rsb64xegO9R4HrcbksifO1XwZ5LtSjK90G8T6hzQbPW4pzJgb+k
Pd0NssqvfuCXhdpvRkIJ8lsRo6rUcVMwxmO8eDKs3uJsvS3EMa0TemCVqK0sjkW07DDHX/mypSkX
kZ4unKcSq7dCjsFnGLO8xSmFcPmGmUn+bBywHUWfKgkfPYTfLwEGalZEhRj65znYtvGq3+QrfyiG
gemZu7ss9k0nQtCx3pVSkqWocGSFlLtbmdU5+P5yM0XeU82dRU3/PS/9PN45/tkT+fMLI2kWYrhF
4HHdY72A2rOraUX15BLdKviG9l++uao3ouvAShC/lKUNPMYRYjxMvidPXXNq8G+MxB7qIAE5mIic
DTDyObqTtBXg0va7LIl7aIZBsvCGEZxrp6q1PfMWrHqgYKdxoOZ3EdC9nj4aF1Eb7jgSqXPOjYPa
VU6sLzpty94XhzLEpS8F1qgQJWCy/Cl3qBQGe044hGacXpXrCSdK30MTu/ChttcyOgduezJdWhKD
bLxTSns9N5YOvLEp3IRQ8qjr2DOnxbfC/X6yk/TjYIGrCjJ9ghdRMp4G9KcvbKphl/g/rWlh3m6f
eYgNvSCthioeoMQypuwk4EzzjOYWbiAjuNQE0fJq2yMGKjnvHSUVNXo/sMWp8fidl06Y1OSLSmuG
6B+ePratqv6280Z9XgAqADz0aoaHLufuXZuXWc7Pn8S/gS/JVwHe59w9uvzIx20/WJun9a9nvyQi
760jeRi0RbIPQMiQYK6zfveY6QadFtlzkQcDrXcyixGCobpfVYXKsKMvGB6oV87gx5SKBN5nvb+x
eHW0UUW9au3o9079itWu+2K8G6/MsvTzSj2V3Dnl+yTLunwVPPxjSwyn5H3iaC4eNnwC35kdIyE2
YfcCIWgzT6+4p9Sb0Mnd8R1yPdM1LlShdvACPePako2yJ4JkHhYKHxcDKo5Bj3sEwNxk5OaaoYuQ
RcaT5DlJD/rgNET8/ly0u+dxScIGTquur0hlHrbL9QFroYzHILWoOi0GObRpnZD1kWFixBaRRvzG
nfyugOqLGRtf5Fea3Ai6W5/JIKxHY422HwweYfOxMICqoWfQ4pfdlcjHu+JJmE0xMwBecj+JTYY4
b17jcf0O8aWvxAb/qHIhs4230Tjl6AcHA6YkcD8NvVuizl+cHggeCe2FdADrLBW2t6Xh1S1X8ONM
BZKQQ9hVA4KnndCfCsp6EXPFFuOIk7zBJ0nOkek58PLGfNgMtTVwYiE0viLI63GIhWpha6msmC6H
/y8ZBETRb4ZVJagljNiQ1cSLsCf18h/OODrXwdnq2NgwtXMTqpwrwtiV+5LC4kVAIe9iXJVLRLPR
ETQnl2VIyiWmhWeJfXTlkzQ0chWgwABDE9hrp/QH6oT0uenGfxNWEwDlqFgepEseZZYTa7uIl+6x
ivhgw9Q9ZuDXdg1SUMWQMp25xkI1mxV3vqgDbAwtwVSFrO+S1Es9z1WeoSUrERI0lxBKvo7uK/nq
LitaYC1pYHPSJkVYz0Q5mGfSh5yV7BgTtPich2i0oKQwgjTwsneg3W1R6S3ruGOmQiUn3i3LJrtf
MQo0c2S3bP5lM+RNLNMHSxpWLn4CwafBHkNhooe7sFXMz2mlCuI7bCB5COsa5xgwGrtXOw64N+Q1
Ssme9ivzJG0DsLg0jG+nINqIGP7Um9RY/Reo9jczYkzQ1l7inVCfEY1FotVLmuBqtZr/7cQN952x
2IexFroPC8GiABo0D5qVEokYreA2H5DGLlcSSZRgamrvIWw3z4BGzi65k4Ug7feqKPnMbSfbut+4
Dik4S4U8pvn1ngxNus6Cc9BpNMF/Txkt4Cscpzd0O8Zc5jtR/Nz9SZLuKfYGP4ml4sgXbLPbSAPf
I6Zr4NDh82z6tWbyBTSA6+STt28Yb/sSy3SyujdyHlZJTk8PYdQBPJ92sANPGMkJVfUpGgNcN8H6
QH9CSCTC95UN2i8wJhE3Ssxm5zhhms/UhuUK7QxaF/TjzpeLGZHPpU1WmukduV4Hr54YkyMC9LnH
6qpPOY3L3HQGgI+rQQ19wVHRj6LWT3zRzzvKvglBF4Je1gz9K//JQDxi0EaohzCjeTInIoozrgMM
9gertSZl8ESSq2BJFavn53uiJghSI/4McANJK4vx5TKXrkcghRGr3lMOtRbaQ6VPPSAwoX0ReaJB
rMCAL0B5TBi8OzLsmoW9yWb1QbM8baPBmWxZJqp6J9zKzPXTAC2cr4BT5rjmJAKdnvw2wdFQcZ8Z
3uOSNBkaox9LOqs8R1Gk/9Kt+rzuXRRpBMO31GUEZmWgzOeOP4Do2LsDq8TqoIGpFJFqOMMXA3jc
5oId6HdPP08ZAjKhFj4VsXustORIg1rXTaqksJH0bBtklTU+QDsj4dzoU1DsMnuKjC+QfhtUYr93
rN0sQvFcpPtZMVZC18EU0QZq9hndn3bByj7SqraHovE3sIFCfzv7TXaabWNlkAEW/cMYKWw7d6Py
aZQFSLDPULcNS73Z2OHgAmlEFRbPhQcrNTvo6VEDQQsHwSlJjgGvMlxWx0fFcgeNkY4QvzjwK+Eg
YMv1U8ohiIJPZ4z9xYNB5A5wx4MiLFJ/RhF1vbMEklZ0szpo8opJjGzJJKzWS/tymbeFdfDPNoqD
+p+qLnEBRr4YzedprH233CWrI1Qvv4u7X5rTlklBiTczEPIBVQyYoSF4/F8W9GP5z7ApA2bsqe3d
ePM3HZhx1prjoHTdjqKct+97WlgoyasvxQ4QsRQddBX0OktURj3lBM+KxzI5Wxwa1V3PO9TEkFhb
nvasgjbsJX82cGmf8Aupp9cQDyjV5RciQ4ACaTcVcSDzNtabgc0ExCCtzvcTdG9HplWklqFBTLer
3B0ZYiapTGHOgrybXxriDUJ5iqcX2sYSNCJgTT/LHwv+eAKm37aONZQZfoM3v274VyS7PfC7zXYS
dFh9oX6SqmzPHLLYREdNBYLp8SknntLwzSofaHA7jpZBpirvPKmqHTbwoPqxMeZJzWPoBqDnuIer
YXoupJTum00EKgTXGZ7sfoANv1wt2JmuddBtbUHnj/xTTtffGWs/lEn3fqXSUxE1jimSWrJCk244
hxbtPJ1YcDMg6idHLu/vniz68i8mQJ5jM7FiPV0IqCHMhNIL9I3nrqFkNUBtCRQ8odGgIeiTzQ7z
39Khl2HNTzxIaYrIOjbbRN3bulPBOz1kP0KdPvhjFEWAt1tbrK7Da4ozkQW2L09/gnqpf+xAzgPa
6j9q1XlX/NJCceXBwMxP4chCktI1eeKd9QGApjpKksAgRG8wArzZ9JO7FpwfExkN/vdqlFFBqf4S
Mm3OMZ1nHJPKijAlucYgpdoj28QK3EsF3EaUF6FONQj+veNXx/UHEwUUxfLU4pR1+4sz1aVgN7FE
esdo+1gs/EVQss4Ut5T4XIhhDLzHFJthjCS0CH2u174vtYybmSx53PCdYP+ObMvZmM+mJTN/S6vN
OfoGN86BoDxdixhHUiaqaDJk6cDpBa7YiGj/91oVy6HoSApU+P2jrrcC8jHKpFMdpDRYnMV03M4v
MqNu3nOSzG9RTE1xmaohCwfJ3CVNvORA40pmCQEq8v1GZZox7sWa4+XcYwxstdYS+Y9Wpm/ChUaB
C4YmluLb+TBMyfpaGkKCH7tTo8VYMM3o7xw+FwvLt5do8PubsmsSXV4Yn0AbCoAjvtWHeIOqzLxL
wxvcsN+zGCP+bkiPFHjbRqnIxpxpC8MiavAZ9cNDR57UdEUMCCNVFbTqYDtwqIpT+wl6azHVH+WF
gzziyubM+zmFKm//gupu1hCOncRiSPkBMR/IXFam5k9Wo29/VS+0i3mWgxJ5cmc4FMcqzdr/Y3Kc
m5XxYZkp2MZdHCc/4ox0NPDO62wfV8fWmdJXDQD46O5kOuS9joWXfafJt9ya0AwOlsqIW7qj7/CW
sXQGz4gigrRrZWcKf0Q92J0dHGIJlNBrsfNmP1bfnOI88gMkIdRbakZydjNJx8AaUdCdCEmLvvRe
0A1TAU+tBHjKhmZLI7dZcraaw3Qcv7QxgTGPYBejfynr8+zkcXODPyCVEC+AovVcDbVDCN6zmkzm
gRxRPcCddFS/GjZnF3UQTCmV8PGV/V7+O1zF87GNvuJBPb/LExBrEK4YAI2lHn2sFMkM1TLmGB7d
F8Qck0rHtov3GZvVPQBJEGXSVZSX9gSTwS3dmaVUxi3R9fykmPlErHrcfyVdnhYoqeJulCM/sFxv
9TTDIrhh0wKfhk7lzfnOPqseZHRVr57s29mdggWrr1MHc1PYIO9SqQO5AWgGJdmievyoAKhoYhTB
BownULknyo/OA4hmj5cfB6eDcQdHCrBS4qcQFsDXbHfxvXeBoNVc1RrBPr61JbvfugXA7LANq8eS
UzKlNirwJeKtQZTUoYMIcEoQFK8nOGoh08T8tkOiBbfZZ4uXMec6XJYQLBs2rwI/h/DMyWoAD4kQ
NxCItSIDjt2lsMA74XuvzmrQbXSFKiJS8EpMWuKOPcQglTvAB50HyvNmVZooHA8IjMgEiseUfjfI
RBapPpboCkB0ytiC0odJgThrajwFCx1R5891SHFlxGoWC9MYtzZRNlXoXo1mC9gtBQ+HPHn+urCq
IdOoPN7o4+yjJpvE/6oijX58q9IJl1eCrk1fy0/Knb7uHJg+I4T3YNsNOkreMdWiUIuMHTfd4iqk
T2ej4Oi6PgdxdiMmtmoLEF6ZO2z8SoebKCKhjy+xeT9k4QzxIIY7EwD62vVuQsuOFrR/cfDcXa4I
XNoQAADNPD6J4Y+pOpzVkW0yyTDuhMiKF7Nc4AEfyrRvSTk9XVV70mRVYlA0QKzIvC0Pdk30L666
wObnjkufMJOrFdLHfZJPMM7zsdE7HY09J/gU42ug/PIhZtGORyxPuMF6hemgKPMOlmHLLHf85Do6
PqUaQxtdhSGIf3wCKSpALQ==
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�{�:�U$�>��lJQ�tO,<Dm��}۴�o[�7�Qꍸ��oӫ�.Z�Y��&e���Q|��r��!A���5#��]|��E��r��&8q^�Kw�[��G����ȓ�YS8HHv-��C��E���Hy~���1�P�v���F�al��$�C��]��T�T;Eo��&�0'���ǘ~�|�l)ϻ�L�� 8������:���{Y���&�����1w�b�I&w�U S�-�S ����觟B/@��je*b�r9��Ԓ��V���ssA�?3�3�IA��[刊k����w&��D��݅�$v3XX%���^�n�/jS~���r ��H����&����0��En;{�|!L��~q�k�.� ��� `Bp�;k��9 �O+@����K.��&�I]�]�P��+5�g��:W������\m0�;����vP���-nߪ3)�x��|j���m�����|�k�6��"��P�Km�37<�{;<	������:�&�S,��_�o���;�r������[	�>��V��T�+6t{��PĜ��!����8�k��OٿTfgHS5��D�jlw&j4�<����/�2(G06��S�I��_�9:�L�%���DF�'��'��Kx�c�{1;�UZ��i����E��/4�24ےSE�<�� +���qt�W*�^�M�>�F�Ŵ�T��)Yq�s�}I����J�1t�N�y�]��~��a��n�a�]���^�eK*�l9g�HD�Di�Ni�q3�2m�2VB��(�'?��������(�-�r�R&_�{��''���"_�ZH�]Fq���1خ@I/�,��_<�G��mSC�}`������0��&�/��pvr�N��������7��$AvJ��/u��U{��yxϧzU�t��"ɠ�J7R���Θ͓r��)�T��c���M/H�C���Y��BK����6@�w�z� Z��j�]��6A�|!���g]Xx����6D��M�NJ+u^��1%'6�9.~'����3�+�*�jT�ۊ��(tMS�?�"��0�NZ��~�ևz�Y`g�v�����͸ݮT_I$L���}�Ӻ�Wp���|���PQ8�E�v��"����������irOh1�����A�*1�l��dj-�ww�*}���&׭E�ΰ��������K�,]�󅿌ɮV���:�����0�@�(��p>��%�166�����H6-�c�xp���m�O<5oD/k�V�J�6^K��F�>f��[s��c��&K8f�Ѥ�ti���2W���Ej�{�pC�mag�<c��v���dRئ���|<��Ͽ՚���>�=��i����,��8���,�7����gA���,pΎ�����C��0)�9ZV̥-l�����LL�3t���T�7n��u�*Yv�}0��v����`��SXT(�|�>�O(mY��|�$�Ԕ?�$��p����u�:���k�U��6,���g�k��DOS���>��M�o$Ӑ*�f��$	�>��<��O�dn�o�,�ss��:0Ue���.8��b�����l�I�M�#��6�����������D9H-zr�W\r�SZ����g�S�RL��k^9�TK��^X]P�(����}�E�j�T�H��-89i1��KX	z��FD��ecZ��^h(A$�b�7h�6��?��pX�#��qL����>�P� C����z�^s3x�U�k��9�8_,S�f��'�пQ�n��wݞa|������(?E��������)o������h�K+�4��:i��5����E��)I�6^�3�#���^�{S%(���|^7��Ґ^_{���\Dx��z�?3/A��^5Wp(�!q����#������tLA�H�X��¼5�T��n|D%��N޷��1� %�&�Qj�7y������ח�q+�'ˁ;�q?h���h��\���p��@4����z��2;?V;H#<���h��F�?�l������:��N�y^ig�����P��M�e��<F�(K�:���t��\�%��_��\�|"O�\>9겈d�}��!�^�|
�8�{(}vm?2
��~����ZfD#ݺl{d�&h�m�T�@6�6�E�q�B�ύ}����s�q�?���!�����z�-P�lӇ+h�-�<o�/@��G�d�����z�H%�;�X�R���qZCK��^�/X}sF+>d��O_t7%7q~�Xi𭏦C�w�H��o7����%��e�Xof�k��D�kwUϫ��NU��o�8�Ό$V�0��,v�b�{�b�Y��T-	�fi���K�~C�I��EX�:���`�`�ep,��F���{I���N\��Le[J���n����H`W;v��Tԋ�q..��M�?m
e���8�ty�'E؛�<҅q�@׬Vٸ����5i��퇰�$T;J�pi��4yHx�om����w"�D��H���1)x���aT���`��sV��:`����{Lt��_c6(Gx젧� {V�_zd��D?ZT
�O�q�I�� .	mZ
&��&�g6SV/7b�)v0l�2f�Ӧ�e�ψX~�����*����U:��A/.���<�h�ΰ�7�aj��_(��׉ӕ��;��{�{�A�����h�['�7vP�.��g�� "7���g�hCi|:sc�g���n7�lQ](�Z]�zI�.�v*� �X=�K{��M���F˞16����>
�n����"PR���r����"���b:Ɉ�.b'm�0�C�o2i��v�u�TE��S���nuI����t�O����V�k�=*&e�/���Yi̇cy�,!&��5��#=v�A&�Q9��`��pKz�<�؝!�$����c�!��o�kPP��ep�N�A�mZ�	�EV�ȑ��jMi�ZO�䜖����w����
S��e���o�VZ]*�su��=�/Jܴ���D�	�Ȃ��v�_lD�[-M���7�����I%bߟ�Ĉ�_�����#: ��gzH�J�;.~xb�Aј���sH�煳���-�bGkO�C���<�W�d	Tr��Q8RE�z�
��Ã(�j����̓z��u�/8�~r'�bf	b'E`�sz����(tpDs饼�26�2��%sҰ|�j=�}A���"<��s�Ƅ0o�:?�ѹ���,�U���uG`�`e[4��@:T���t��7邢B�:�Äp�6����J��V�@!ד�@�O���HS׎'n�<,	e�K�$l�k��'��ΪYd�b�ko��!yu� zV�\;*�^��}��Q�7K�|Z�x�ۼhF&��`����"��uSw�J��6uv����D�2gf�R»��%�,Ɉ-όO?	�F*��0�"B�R�^���BN�:vC7����4Ȏr���ľ�N�(����B�?����Q��]N5h0=��`Aw�����J|mF�����_�K��F+Ӻ���[ƌ�9�QZ�����8�p�^l�y�c%{����FdU,��2�
\3�|�F��; �v\1G�2�I�i�Sk�ێ�x��vQ�4.[>�����5���`��ˏV��Vxr��o�� ʦ���<�6��*���SH��_Xൃ�:J�����R�pP��8����AU<G�Q�vD�cuһ�7{SX��O��UW����i��U��1�J�)0ɥ�4���+�3�� �W�*A� �S��_�=�i?���1m����,"�����c�
{h!%!�8P��{_���F�q��F�m��^���҅������5��b�x��qI�]j�����)�tvn���Ѻ"ԣ � j�/�]0��?wf��X��U!;�Ϣ0��+�o���y�
%g�]�F5��=)��[��A=�1�SƇ5G�e�9	���W�&e!�F3��a����gg�����s���c��]����3�k�mi�44�C^�(����ѯP<_�,� �� ��dq�ޗc�K�.�J�S>��<���u0���8���S$#֧_��Vp�I�]��Y�5�E��]�Mހ���-��@�-�u��Q�s�U`�>L��`h�A:P�(��Z.��,���:������T{���4�tse	6�	L4Zuu�_w����s��z51�rϣ���P��#}'��M���z>'֏�49T��� �a>���y�	i+�s�v�����崩YH��8+<^�L��:������b�/�*6����$���A�r��D´�CQ 	H��A�ϤWƆb0f8��S���#��h� W�i��K�,�Y�P�J� �a��Sh*UQ��0���țYp�t��HU�^�Ś<Kw#��l�Uݶ�ǒ������s���/a��n��}�G7��H�F&�}��㗳��" 衈��M��4	�ZX3�ך���d�[����pG�G�>>^{��/�A�7��3�h�{��;��U���N�&)>,H���v1���7��$|����_C�.���?
z���#XB&ߎkɴ���'��\̬J�|�������o�N�m�f��?�̗o�:.�V���
(�`����>�&jP�FUG}��K��z�tgHbJ,����R��QG�P�:�����-�n@�u(�.x�X��[`��x�B��X�t�;k���-����ܘ ���(\�7�8�4�c�;=]�$��i��Ģ^�}���!ɘ�pq�i�%�"�/�o4��[�$�K���h}m@eK�����[�1�
*Y���������B�t�B,Ҟ���I35�ܪ��V��oQ$x��Xd$���ov�=&j=�в�us��� O�
����bfXgsn��,nr�?�~�3�]����Q���Y%�9W8t�O:97 ��j�~�h���� c�n:�o�[,~�*?�N������͂�ʲ
0b���"�Y�?�hW(�̤\��d=��]�Rw�ylE�[We�_�4j%i��+�(�r<�c�K]5Y��X1¬���$�@�|I�]1��.N�C��b��It��>��xc���fǄ��/F����vK�,��W��*g� s�'a�j��� H':5��c��[����u���`�28��1�I��+OpE��y��րi�`k�nu4NHϱ.N�d� ��C� *M�R�lg%�?�N����M\`�|���A��:�}��A�<ku�;�ެP�u��&T��"R��*�~��4���w+
gJ��[��B��+0>���E"n�����C��-���XnEH=��I�+,S�?��<I0=��1k��'&�_rXI��^��"�[ ��Z*��#"�8^�|��j�X-��n"�VY�.�>:�ޞNk��%�]���M�w"������P,@2��P޶��r�g�#�����y��l��Ɯ��NC�Ӧ��S��	�Wc ;l���� �.p4!�ƛp8����% �&�a%2OeL����G%�[>ѳ�=|����i����V��w�/G3�QI?�9��$6�N��lӫB>���Ǽ�]e<��W���8��Sp�ظ��ڵ�{ck?m���i�aԞ��tTjԇYP��AK�Hce����5��M9��x�`4s��?X�4k6�Vy��N�"GT�3;>bEy
q|��I���⹬�3��B���	��1��E���	P����^�V�a�+ɜ'o��y�#��g�j����y>Q״�F���:�l���W!�ϊ���?��L�-��f���Xy��5��ؚh{`T<�G�v�?;�,lA`)��UV`�딌�t&�~�r�����"3Ȗ�{=���=��)�,�E�qo�r|�:�m^f�ʦi�H���=��d�ހ�w�}�*ɮD6T+M�7�5a����YL��<��������,����J�к��8s������3������[�B�e`�[�w�iå��?�+���+W��9�܃�`�C����G�X��jMN��O���O�>��x��3����z�վ,��
��Y�M�<\�B��%R�RmD�﷝꿣Z�������M��8Z�?7A'_�95PS>���<U��[];����m��9�t�A��"f	�����e�S�}dj� �.����J��F�|ֻ���QCևa��g��Jhb�Nwx��},ͫ�J�)��0�9�S6έq�\�� �`���3+�P�x;�Q���c������P�[�=&T{z�97^�SN��}�q�.X�g���n�!�awA���k�%�F�Y��,�
��~�F��흢Bx�� "g��=�Lx췣Y*ɓ�l8;WkS�
��9�#�WRp4�����w9{�N�K
���!�l������3�P|`�^N��E�y����"�ϼ^�DP]�Q��d$�X%�H�m�'n���y�b�G���՛1Yæ�P�%�&�-��lz��*��VG�::�,{�,+cC�<�m��ܻ"��- cc���et��T�\C�G�!�-�٣�p<���]ٱ�]q�7��d'x%~�-�����F9 �jXs���M�#�^��d��hPr(ek	�v�]�XM�w}̋�ۡh;V����Z5!+�<l�����{���=��'��M�:�H����|G�H�a�b��QE���o�-����m�U|�ع�N��ǲ�.s��5�L��vo����iM��������#���.A���ܭ	b�zT��Ou���f�ڟ�P��~���m�|Y��R��2>�5!�<�A�dJ�����Iv5�>nAՂ��/ �R[@SG�]�	Dg�r��Th&*�2���⍱�1J��φ��Y���O��Bu:����x&Uj���h����/��<�}�Z�ǻ�$�����Y��\�J9�'��\&{�g�>�Ώ�i����Zq0�|���I���|� �a���ga���}E�y��V	���@bE(녽*U��b��H�	����꼊{�\K)�J�X}�r���`34�QK��""t7P�f�T�@ve^�/�ǳ��E�����<��(08$�|����#0X�`j���J�xO�sT��К���j�vjH���1йח�(�����W�S�TME��������s�_ 0�Y��+
��1cF����Jo�Ҟ��_L��w�l���d�W�\�ߨ`a�5O�#��V�����{&�J ��V��������P��כު�'��P5��M������	�Ô� �O��K�����Y�K7~E������,�6�L� �9�>g@���ڤ���*hI$�)9�[ns�#˺vz�F��u�ΪQy8���d�؄v�����!^����a\b�W g���jB�.�{|}"��/37���P�a�����n�v����~��
�;�B��@�&�]�=ţAD>�E#A\)g(�o��ڃ�7`��g�|l�<�����ީ6�8��ʌ��j����`�67z�t���#Y���H��<.�q�w�G���p���p(�*�]�&F�NA��
��ƹSn4d��}e��.&�C41���9��d+?�;�ݹW���;�؟��>��_m��3�!��ZJT��[U�#���"�����W�b���QKu�.4jH���K����sЫ�" ;M/jp�t�[�x�{)��^�Ed��Y)��
��u�͠���ss:�/"dq�[Q�+��j���s�lի���~/{�b�6_]z�n���,�Ba��!,���+����"Y�3/%��A��?[��.���v;3��QU�:ź/�1����؛p��<�}�^���R�h�D��hIr�>�!0h��GD�<^D<�yS��s̹��7a�.�Ċ�8�ӋBRO|�dsy��l*�ߓM�+J�g�}ʀ���B��y�d�<��-���Z"X��NB�f�B9��ocpc� �2��;�r���2�n�oB1��|�B�+����~��D
�b�B7(��21c�Q�?�8��<i;����m�
�c �ݩ���v;�M�s�ߣ5|����l 0����C���vY��&���	�;=m)�B��M�%Co��JV����<���~'�^@�KH$�<]�k��a;�_��A6q��:!�
R(�
m�ek��)��j���=:*�Fh��J��l����ZLN�f�_X^[7=�*����m\셙ؚҿj)�͙v�/$Y���j����j���1��]�����dQa��JK�I�L�8�Y�J����Z�U���%ó�K_���=#��M��Q~N��ವ�ޠ[ٻ�>�cj抏�vxX�E�u��*��ʫ���?WH]t�L�_��7`�2ܘs�%*��:W���P���t4*��E�G0.Ȍn��&R��������]���Ɗy�i�ß"������_��Ʌ�6�a�1w����X`��E%;��U����9uHׄ���eխۦ�L���L�G���`)��86ŏr)�9��ȧ!���	�7�e��*�Fz����kI-�ݨ�mC~�"푁.b�$a��N��l�JI.L�9�C�^��|��_�!�s��6�������X�Ώ���4`�c?щNd���	�dy�p|��ର�����g��3s�S�2�����9�\pf�|\C������^i��8/�e�(��_���nﻪ���0�����E-��Sc�֦�1@nR/	����o6��`��;.��!uR=wb&�r���;M��s��[���{�p�<��ؘ*Vgcq�Y1���[n����%�HRS���	㝝T�?;��#�`;�I��4���z���SK�}�D�.�����?Ih����]*����&W�>�(�\y�8��S�N�)��ʎ���1 ��H�#oɣ�+74��
Dz�x;�X��G��[ޚ�).&�,�)5o)���e�<�o���L�Xlo�Z�q�~}{s�OvQ ����M��w�`��rB���T�h'�j�JK �@XR��< �W��D��0��}d� ���9z����o08j�N|(�6+w�}��%�)j���HJ[u�d�5E�Yʵp��G~&D��7�'�#Լ��:�l��K��\JQ/�Ja�3�������轠����u��y��K�i�+�T�.��|<Ϫ�����?��⏛T1}ta�H�������\!ƈ��%�_'ʄJs�g� oÆG��Uj8J�.���:����KQ3]׌�2��vp�r+�V���"o���ŕ�;�����]�>�ę����H��-�w�x�V��� E�2���Y�����Ov=�TGp���!�~��Fﰪ������3l��6��;�V�w\ �r�>X����tW0H<Z_��-���mi�.����
\�!oҁ4�vKY�n�B��=!�?G������n��:��P�4��Xo�vW�#�U���?Eš��:W���b�%�ձ�1�^6�Jm�i�,�
:����ǌ��8�� �"�!�F^]�~�#��!�4�T��j"���O$bw�L�`�e��u蹏��Ʉ�N#�6s�Dm� u�[	)ND�w9.�x����k�aVF����/�
T���O�%���͠�٧ 7�te�iQ��/\����>��&�ͪ�6ƫ��g�����A�I�pV��'�Q��=U�G��)�V��ʆW"��١�x<����_0A&%�zk.�웅�t�Pܡ=��:������O:������ O9߭�ym�5�Ɋ�q\Lފ����i�<t|�T�2h�ϔr� P_cܖsd&_��G�z�Z�Q����3��4����'nr�冉GƎ���<b��&�c�+Wu��V߇��]v��9�PdS&���u�=��z#F�.Pi�Z2��64�s�ٛ�9�O�_������'�sf�����j(�hr�d�/0��`����_s"�(B;��EF�����1�~�\Tѐ:�P�;��d�4�[���(��R��p�Ǟ�O.�qS�-CG��/-� ,m|�1M��>�N6"�vm�?��.��%�^"���v'k�㤨z��/�E��x�L+���/�􎆹p�IG�">�������Ww ��El8I:��o�֨�!;��f<#�S�Cˋ��e�٫Y�(M���ߪ�&g�D�p���9���aZ���O|74F�wQ�Sdz�¯���v�����/���ZX�+��V���+*u ��4��A�lϕ
{RZA�S�kAX�|�	O쳐�P��)��ÂOS�8Qc؉"�b�ܫH{Z���!4��l����P�k�&7��^�>|/J#[�(��[y뤦l�	ו���g쎞�&�m7���L=.����	�8�Kg�8�1e
9�E��$1@���lP},���Y�(�٧�������KG�[|u���e�7�K���`| ��f`[N�&f�#�5�� ׍�b���NZ�M%$���F\�s$h���V��.S�5���{��bR1͠d��x`��+����9Z��Or!�U��}��?R6-T�نM��cw,��#��~���f�l�߰fH[��`����=�l�Y��h L�"���|�O69��j��4���iД��£�WN�Q�v5|�����篢�\��y�r���BV��k	�B6M�&a$�^��6k�E�N��*�!��{$?g��p�-�0�j(��A�[R��0�ǽV0��/����x���g�0O�|��q <��tEWT� �N����MLlU��wi2u�p�̔���x{��PG�&	��l^3�Ѕ�%�s��)�D�l���ll�#���(
��ׄ,x}��Y���EK!�6J�?��*[��!��H>��&x	���K�9��ˈ#�cdj�)h�f"	 ����v�,
K��Sx"�Q�V��1�ٯf�1�Ub�)�fR|UP5���!�W)!�0E߳f�/*���T��2�Nk$�`P���!=˱�G ��R�&�"s1�oM=I-R8�='��.h涖�j����h�۵����/���+,��;�[�/ٕl�yX��n5�P��9*V<��nM�.\�_
PfQ�w$�s�iH��-$i?����Pm{�hF�g���]{���mW�Ň�� ΣI^`	����������=Hz� <�X\�����l�
�d�@��0:���¤�Q�c�+�{���%�m���	:ƷL�E&�ts�l���&	c�� �p�e�����t&fy�E d�xW��2��4f�9���d��-^l��/<ɭ;6z|f�m��NU��/����/T�eQ���T'`T�� �m����Q�-��Z�"����l�h(m~Vh�iM������Yz��O���hG�������aQ��DR�I�����$!�W�昆]n�1��N��������yP�KQ'���_jmop7!0� �tӉ�(����u��0��ޅ%�]���=�Q��r[������ FІ�F!o>6'(?��\4F�lz�<ɟ��A:�51X��|Q��?5�y��R-��^�}���u:��"����� R��ӿd�Я��煙F>Va�s�g�������Y�B�0as��X�����Eɯ�f	�g�6Oqq��	W(j�5�Lj�(�̾�7uC�'�m��'Ј���}�{~�k!5K��	����_�z�I��LK
Z�s�08y	�'���"�Ck�֥�������vH~(�?9#��0�ނ���`�ainf��4��"~(2�&-)�� �`���Z��լ�{�Qxl"��b���^��[������q���L5V(&�n���~T��MW��6���/9�Nv:#NV[�ذ=o� JU�9A���?%\b8��g�y}qh��}m�|�,j����lv_�6�i��aڮ�����C��4�qɎ���3�����P�5pK�0�2@�{T�][�F%ˌ�/�Hܗ*k&��$&lY�!�mh��a���%���0�}  �6q�;d� ��u���p�֗#��>�������������v���:8x@�U�}-�s��,��3�6ڟy��7N&�$@�D�?�$ŋ�fM$�_�>˖%�,�X�x�J�ע���R�!���G���N.o��T���/�����O~�	�G(�^�h	F��QL;���P�m�=�â���p �K�>��s.3[�۩��p5T	?�Q�G���d�ݽ8���0�{
����j��%ֿ8
F�}'w��o#��m��<��Vm��W��_�y2A�K�ה�}�V/�D}���_�zK
�6=��R�2��/@I�D�LI2�������woN�Z�-t�K�f�N���uZ��W�;T��]���.ũ%eBS�j�m�y:j�#ֽ�z�	��I�o�����ނ$#[��I\��х:d^�]oi0'cI�9��j��wU˹��O�i%�v6��70�np��Ғ�\*��U1��mg�ݴo%�g=Fe��RDt���]�7�
8q}C��P���b�Ƿ�j�:�	��tݲ�Y��hCo�����<�*��-�0q�Y�*Z'��=-�~�9�G
���+��\=��ƹL޴��fi.�P�,��&�_ �4K~3��sA�����AR�w+jwOK�Bbd�)�"��#�д�c+�4���;A��I���7�*�-��i�5��4�[g�S�됈!�e�����7w/1$����ƋH���PL������&�{��|W�Cm��Ō-��k(���ҩ�`�;�����,�<����0n|��CQ#�p
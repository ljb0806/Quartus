-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nUXqp8b6vkraQzbsTY9KcJpcJ/TKmog0PdbKYr06Jr4PH9cCY/g0h7T/vPd3OfV4Thta5kYYU6n3
IHwnM3sgHU/ib3T2z9ifTTkhBuAlEePTHRCw8+U1b/zgUUdMEPgqsIyjZcN6xf6uTIKnCGiCbS6Y
JME11jRlcMSQN6OlBnpa2sXSHoVToYsl/JM4ahM4EQPPibAHSYvf1K2wpWh9fVNMF0DysD2Se2pK
fo40AVmzGGIKIkUW8BQwBS4wq1RVSe8svxuRyBv0bVsCa3YTcVuaRn1M8rn5JmEV6S99h1VmQYbi
szzMcCkzd1FbiwsCr9HVboHDWVmj8n8YsxjnTQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26880)
`protect data_block
r0zhFamGqLIEnwtpSyo1K2UFotpK6q2oX+JYuhLoME8vCJimah5lCu24TRExSmNmVGF+dUaChKX0
mb3+MXQJgyOxZv+3/WQGFkAOyRojHFUYfjqFMFn4u0VOuOCnb4PZSGOodMAQmz3S2t8mtQPWRuGO
kI1xHTWtZAKo+iffAR5g7Td5G+cXMcczVoK+1kXrK4zzmyS53x4pDKa/VkrCCsVbTHNSd5rl73np
vPoQTs6No1gqCd42BDGZsB7KiOU1a+tU69/Ghz8jiQAp1Oz0BAGG7N2GfDPrp3mW97/XX+PF3Qhr
kxU+RSONORWP67+DvTL7fFt8xgaDjwWorse7PE3VNE1vd/KVrSGQtjzbchaKqTB7H9RZ2V8xCfGF
e4J8kmnvnKSa4wynsE7ZQiJw+69/fPLC75+Ixl/i5Q20BBr+f76p1CFmoVncxjxniEcyds0FLZI6
LYLCTZosM6tMJmCONs3m4jB7A9+IPBeg9a7N268sarbXMBsHk2LJyuz0A1r5d5HHQ76n16Voq5Mb
AQsXpfzDuKmkUw7CaH3tWbmBkKNoagQQqhFuZv92AyDCfM4EHebRzrwc5VETYt4WuRuB2wlVC4mZ
fSb3H/weCjhVlbJ1gVvFAVBOsJK8TnVLIFKIIW64BndWwqOyaU5plvwDQg82LKGydh5/aRbGdtXa
By4BPBZBorN+dRloS0ZQzf5//Zl5KoXa5uWk3sXzwbeVosoTsVom+M3FkemiR+UVRviQS5cldWuM
5OL0ChAqNmRD7osT3ez/+d0RNcAOu/Z40cDM0zHL7tM7lCoc/jHn1l3D7Dl3wK2rfrxdVfB27J4/
juaQpYpcTrb2Wwf9LUq++ZkWr0QPvqT8o8/GkLO4WHNVHn1G2safJYc2miHwMuU9JxV+ShG/xKnO
xfVcSHokZw666lwvU2ZHqbb6qn/S213KBgVtzxLqZyZjhz8EOoubUESzyeO1ICelkPsI+ffUt++B
OrdNupuiIQpTqukg7VPUbF76enuczC3usm+J867unToxSLCznR2i2ds6IRMlSBx5nGverpZgHS7V
YubmI+o61RmA+EOROa/JfhMOTRr1B7i3K+yjbWV9X1WkwAorTlYYFQ2v7KaSwp2yiAL0/8eEQE5w
WYKs37hrnwQnhCT5MUUpTWh+siyJTXKupcY14Tew+uw1me3Nb9yu/PlaOOr8vR2KNKvTXIBYNq98
a0q28UN/er51lgZK65kTZNAtgkDx2ps/LUu/gsUshS90mR1zKy6gtdK0qYzYJ3QQOS+xL07BefiR
vr15/ba6OHSx9aJ023UfKCB8YTaYOT/rtToldV/vAqENaOaaTyGBP4K0aqpdsT8qfBei936QHMlI
M/YxvuQvoOYJlbomrNMHw0OUYByYQfX7rAReJ4wqTOq4EYZgbQmyGsPb9Zv6N83ikwjvUe2nTepF
U+Chnqrw4tHFCpQ4sfr10SvJhbZolKw+R3OMEK9mNRszGacw79S9MIVZLGcK1yKGfxfCI8Pwp9oq
KnXbRNBeg7l9tKZ09UyP179hgN2OPzXP+fTw5sjkGiEs0Udhpmckbb2OGCH8CUXApqKYqoc9bCVP
UoskHNZDg3lRp8WhvAmcsNIchyT0cJqnSMWhHIwvLXQXCYTlOtD/PFAzpsUb34o69yp1DR2Joc9N
Z2OrGMd/Vi9JIIb9Opnrp/rNh5ZtvsJnjPuNyp9J72DUP+F+F4AYQ0drNm0igZHqzEMIjbGM1KUs
7mF0SloHhGfVOTHd+9qewdarlrgdWxNuYwvgJLFE4ucUk/IPHr+CwyXcBBcc6XNxGMSLqZvbhzvn
o8X/1rcxigbsoKtX6gxgBONzLGXDkabjeaSd164fKgfch2P6G3H6yvgUkzWyAEBm1Lah6LJIJkZw
vqmjwELqaW6J7k5r9kGEjTPeGrVYvgrsDEsL6wLjwAwgg6bB2BA/kT+6ZR3vCyrteWMIibJNLVjK
Z5AnCDXFapIn0HxRbAibm45nUri+0VB5730WtclMeRFCduGSbfi1vvdn+F2s30Qh8v0W3TlxuiqQ
WBTmOaoykGyxyZKH6MMrw172qTQyqVJId7tM958l0xeWNT/4wfA1aC5A0nVZN1FAEDFpDqkZMVsN
r7OoyS6Mt7nrVlEy77ugc8sYTHnOCGMpxUUFbbbi6Na3i+haqq0aD/urd6yWoYxT4ieFz9dTnyT5
NonKyDzglVx9yy3bknt10Rdu18O0180JT38jFkJ7tfhok98ybR2cnjvywHaUpZLkfh9ZFm7RY9ik
6ePKbMcC6kfWN2gMM1Wdt5mTtOWSQuR+QyuQoaiuXOk+CWVPzY//2yo8mN/CrQjaQEj9ccWADjeW
vPziHS0s+IHrU3dSkhdcou/Ewhg5foeT8xWRL7DmlmW+9edSnu2EPSZ8smLC3d6y1YQmyj2zdnnu
s1YMj5x/9Tn2yQSvmkUBbDIlP8DP2uYr8ds7y5f/xhYdJPj8AJFWfEshKhmBu6nhM+QGgovYBs4r
bBgOUMQ185aKh9+03Y50BkE7HJu7sisVxKgaMBmTV7TF6t0easO8hNugVd4OJYDxuHoyk9bGNm/u
8+nFg5wsAgF+KLrIbOFN5wOSQldG9j6j0lHEQ0RPDbZ+cR27xAO/8j7/O+ZQ7EnPT+Fon3D0lOVu
vqd3ZqzyhBO3Pkzq49pZweVdNwk6GQF0rpgQLFmzM9RC8+6MKIrLhnNKlHmvSDdKPf2UPbaifBqh
gqjoN8LKV7DhwGHP08sZ8mDCAumEJbc8cFqbSq4cng5HHzfkD6saVC9dk1vnaspElE1gOegACpIq
qRIIWE8g2o3RVm0QVztNpPSEYUrLvXW/aPDOfinoJtnDAeL++IhktsJMOTSBaOwdx8l55ma0a6Dd
8Vg8yhDpzPZraPJ4EZNZIXOITPIX1/eZWiws0snk2tEFfrfWQ4ZmV6KlVv/NOFzKeisRlxwejhEc
jopDJvVVF9tC7JRThYyA4e47vlB5L8rO+s5eXryBvsnlrft1XHJb8It7r0q1QcTK+ZPwdQ57mQIx
6BQh0hIWjdZzNycdibQ9X40u5al74mctRjZ6zJNDDh7pKloKz5FWDcj5HCDnYyAR9TDpwpRIaJe/
c+i0SWLIS6BCIY1BcnLkmzhsnMAKTQSDSiTDDIFi7vpCkE7lzV6JTMKGV7dITJaYaayVvAGI63ov
pefqWTgYKYlZ1UJY4CvTQESCqReTGRcKaVIFSfr4xzCu4lKLFbiNggyZ/2fd0QsiprLovNlSAPIn
WOdhj20H2WsH4MqcGsuTOVYgKtwE9Nc9rkyB7VGorQFpg7CsGeKJXiFncV+Lgl7AXJ25oeydPTp4
LJf8niMl3UqRh8mZG1sg87bVCG0BSc0jp8SInUkA9aBK6NxeLUrJeTP8TkUozr3l3d0cgNdjZBi8
f4aYRnT9QjJbOppQJpPagibPe7GGPYlvMAYMOa2k/mVJQCfsGLwCkga7AGbAA0AMr5qNvkkgXXVA
h27eQm3/oe2vjxjzjJk74CKNw3coSGJalcH0tCbbgJeiRzxnDQOIO++bQqNrGCBro0pRGzeWx9BM
QFLzj8ZFHHN3/A/YM+GrOhmDpZ+qZoQoOuC/cFP/0OtyNuOowJ5gzwF1iTExtuCL8JxZzPX/1GGt
40jPO3DWRzuEl4dv/KWb/paSdBFxG2kwgMLusEO32qNdQOPsLKd67MEXrLuSPm3qg9RBdp3hBklF
MoYTp08nUdqHzdL3e//8Y7vMy6JmtNqXe4/HtAU5iGoiHJMTQUvF/RV9r02LjAOxBjr+mLdWEdO9
RIn9+V6vhxbogAcJyjkefj6sdEUVFGL05iT7huc8A4nS+xf3hrrIKcW8Wk0lUg0SU71RK8RZlY+v
YEulqVm8AkUvU6LiHiodTjFNYEUUJyIn+hvuvg20p/umDlKbU8sZ/bjeh7dKsEOqXyJM1OY/QOiy
EdDBqB/jmlbKXkI6SHS4ZzkheMeSiNRLhmjvJqvtq4eNnHxvMtkEfsBTvDZkPZSLHLMX6I3IMHd/
X1bY2AVZ2V51oDwBHgZ75agRAQBj8NPneq9UXe1pQQjqFqUqf7grJM/GeRI7Wo09toGMdWMYecuc
dxaAh4DvaqOAJy6C8j4UlJEln7QqJ95DngNHC3f4nbY/ktGRLrV0LWGO23l8fLWqv8oo+Gzq/qWK
z24nP0SwcBfqh+zg6uD9ji1PjxyHDCHwwUPmOubCvVhRyqP8j5rRTrhHTtxOOQPoETBm2IqfMcj2
apsUkADY52KRkUAitKXqHvO46a05xJAxWa8mPmKapOvTCrufTlMoGFuVTUXkceFAcZmZpYA3wZbV
CunlFdRyoHpdRGc9aXvb0/e1rC7OKdDr+4kRpmnvlnj8AF4+UnvpD6/gXMAhWh7WoE19AvlN0hWZ
n1z+dNk+Q58ts8BndpPnxDsaDVIqjX8BQ5N5hpvmC3N4mUz2m8uRm6IpYgUOK/qzaZbeov8YHzSs
YL45b8NBRnDrCVCtZ6X9+ac4ksVxd6TsNTtM3dIoYQMyhJ/fVkR2RFf88huOULoQoA1T4TZkZjPt
l+OF3zGXCPzAFJ1QhDi1qRtC9PT4IhkphMdOeT/UDdwAEGs9l8/9eXusqrOKjZ5KrDrcOCTKfdrf
SlPvNI3fGSyTuibfKk1OfZvzvZc7xHi7doSipOZhxcQEya0HcZzEqFjxK6HnYfjw6Zj/UFCwR/cu
f7x9wOcObaWCXqIkjuFQJs8NbnXVPz1GCOzigWgnuZE+aDvrSCXRdhdgwnE6OvwMMzPXbNfOXmsQ
e2F0mFKd9loio13gC2uPnD73UX3g3qU/DCl//AQ8X3wTjo4UDXKnksC1H5wSNKGMR65tOUeFEefg
zZD0Tn/ESpcWqj61J4XgdGEUUkd9LxKvM5Zd2nePNDGTCs9jQcQXG8IdG1Jjz81SE41prgmhRfDD
nDlOeOUHHyGTXqbt8ym1jxl4VyWFXbeop11quqApF5m3O7Z7Fop+OQKSfhn32+J6NykfF4A24VwQ
M4uWkjuJ05AiARwxRQBtXQ3n5FyOYP0iKsjaXolDjxH77vrnlbeCG56FhtgtaxBv6/9/nWB/GYEV
bnYppd/ainTvsjTfWFCJRIqL8+9Q2CHmakZjyUcChqWC/t9S2s4L+sy+wSajZDRtx0ikUIceHSTK
lDw0vg4jMNNtlO9YQ1J0FVEkSps+3UFACHRkS08wFRYJH19nBhy047+sFsF3CYCRU9AEzbmGx2l8
BFvK9x+XAdWWfFwQiAMzHnw9uj/ht19+mmN6rghhGtCg+wM0047st5ldYlp/U8rEBa7zd/6dikY+
yW51dJb7qAEDz8XznvV9QJFMrw4vsKb/wPqyD9jeYtl9j9R+VLTWyFuWZO5FyxhyqLxuHb3OxfZq
z6L+uGBLsG5c9ssKFIIKeO1NM2zvpELYVWivOq9wuuAjeUao3sLvD2J3ahuEWjK9XtkduhgLhNKN
bp+17W/1N0Oic5YfDGrFNy+knF9bT3zFf3YgCoLw1uXTpMn+jYJmXFUiDrtXFtJqDbrKLeYxpqM5
9TX6ZDLsnpIraTx1J03eC6sodO881O8hjqoeqs0xJ0hlD4UEcuAEQ3Zjs2yHhPMiYxt2zZZf3jXV
xIXeUYc7Wb6W8D1vetpLMjQLlh0ZdXZt1x4X1PHOAWguCoN6RjRyZp30bKv59ArMerqSWyOt6u5Q
eKjWOCDRJKVm70RKsMwuB/nC4JCJLxrs0vKym9oZOi5ncEh04IEFbDkBWTHM7sgBHVMH2/WsC4u2
qUUbT1ybNo9IP64C+i/d+UCqyUVHdAlpKP1xJnC2sanLjGClN1UfA19OeZHjnLfpK9uiIV3rsr8+
YsQIjXVqBEQxq7+09+XAnSi1rNXfAaNElNkrW68GjrZIga4GsAHVlMR9pAD/21hU3+bWl5Y4Jqc0
K/ppwBgAk/Az12hHinb6oLm9XxC4PyxkT56yT8W++Pi8/0YawTHN6j8QpdGKIAvT4EtrcUGkglPB
yaB3ecleAuJ4yXxKyOMcSWNY8LHvKLyk6b76gQuCD/i3/pUuyWv+NrEe01KPlSD788rhvih403yK
+MIHkchR7ZsqluRy67fhgKJqp5Gb9t9bEOt0PtAMXtDiSjbNeHyRt1TbRoq1FNpJwnQjCbVMEmtS
CnG0hBKZnT7j6MiYTEz/8XbaE4IcBRKRpjV07H+lXfjPb468UXvQlRpIWMQA7GkTXmuS/dRuLHZu
kW6PbRVSkiLkeDOOslcuyY2GGIrKNW4u5l45AGg2LzXhjcKBIDpuLCiTYSjWX/5LAf8Pid7XGzkv
SmjMDggCEG/rHay++C8U0C0gW9tNf2zU0UrWCUwaUrfhgAzaLLBma/ldWR59hb+DwhQFI9qn6V1i
A5RaFIiuPu/X9irZjXUDyeHKvLeFWF35nIe8lVrfOhm7QMoUbnKZb4Lu5CgLhEavkDY/n7nczm8Y
LwflCCXQRcvgrRL1iJ2EnvwBiUPWdMU4l4tLzpTJtdo0gXxCQp0Dr3x2p2pBiSR5BY9KTfoJUOBn
ugmFysPt7vKZ9FR/jf42TQe+KR7NQ89StMRwhVcjVNdnWflrgjx4tdHHmRejq5fsg9PTkyaffxyX
2IW5O0bNZFdCH2JhcXf6jTvTEA4WAn2c5sA8eicJP4rSxYx3UByG4QfyMztBREpGMl1QnSn4A+PU
AXQi5wKlRc9uBddsCZXoAJJj0KIG15xVXNDBBOc+XsQE0GH8rD6s4EiZ/JiUczPLmyBQwI/8Bqrt
Sdb0plO1WWmKF5Johgo+KxVNsTX4jK3cz1zOMCN6ipwykyVn7vGDu2Pq9vwE3jwUVWZraGAweyoh
S9ma17hCK5nQtMMmwjEsWOlJPe0i3H5fGk6KVp7sv24wjMp/3M3oggoHGAqKgGxh4M6GrXKYVWPF
DmZYqZm6AjDFDzrvu24xotfFuMW2c+LHZ7Lm2TKmJ7WcolLErPtm8hGXzKBisC2fgvnJKH/Oh0/w
DHZH10fSxDk4oMZi/0dNPKFSYerqp3RtWsAlKLqejoS1H8mBU2yL3ig1C4hp1qPGsNBcMTkOM1Bz
PrrKZumGD4Mn/5bjaXZpjgoL6dKKEptdbxibeCA8xiCkOBjjBxrWiqQAqNKFqkiasjiDleBpLnTy
DTbQ4AbSSb9V5walryMRbL28oMYTFjcdLQN+2XQfyJRnJRXRhz3WRQF9sCs7ZxD7y7mgoyXBQtn4
WqhsGWnP2LQQsb+DhdRFpYzIbiUlSPevnSw/TMl1KMPi6zocIFhFDLmkxVcNURGFDqsgsMKc2RDa
bMM/av5+KoWEQZVHG9kwTUnlKXBABkhvDjNmjqjfAw1OZ2SZtv/eZfm/YPmUBTeqnT7k8lDgjEKu
/zA6IqSbmSjUr5YZaZtQxT1KU4n/MRW2cXmB8/tpwiNOFWlL4LNoHLCPUZK4z5WUG7bCJuz0gQFg
WPyCg2d6VpuUwOSao6OybdWM3BHD98R45XGeAMUAUPj1Bb7SXaeEPenqvPMs/8Itif6EIPB14n+l
kxMFAST9iHltbZHHT9rr2GBMdbxDdm+YSmIjnjGDaey9qx2mXLLqZKbs0XKyVQc2eEixq5nDfiC/
jvD8VANY2KZXVfLzWyj7w0OutYbH6QW8/T++fpK83rBYj/ncBNNUUk+M5Oy8mOWQ3WhgkZ1qt0Ai
5AJxjowcfdC6PYXyLaaPktcrtM8X6Ski5080+K8AALUxmQ+LeQ99QJAu3H3az6WRwanwIRDNctoI
NnhzqWK7sI9PgBndl0mMuqy6sPQzMjM/TByM2COUtN60Cavxa5FnRiyU0SMQzPS/2d+SQDVLs0ME
Epf5h99owVotpHW2AcwxtGepqqAyTzupeKI3szyANYqS6JQDWPWxBOGWFM0oF+5M8m5c/pcdx8ZP
3wLPdRzvkpxZbb63yt9NZO0T0YnTnWCbj7mbVIbd3KZlqxnFpeaLfqXdR248mkkcTGFoOf1G5fpF
AsDmcT8Xs2wVg9T+NTw4h3Lv5ErmgyHE+H9yXiMhymBI9UFWqi6q4uDBrP08FBdOGzjuICbAp+/v
8MblBY6/aLGRQlfsR7u8xmfAjJGOEzdfhp88wMqm9ZVWPlUZUeSyJj1nllL/jDX4TDwPAyWFBI5J
+7BxoN0bmERKm4hrj4rOGKlKYgz8MVNkRnkWx8jnoYj5S8nR0Ll1V9uhOCCCoDTWZLkifFaiinWJ
TDE3MTyrHN9rgrj4ykxBw22ikTanf8QbIzewB/C8HYTapkbcx4gUWH7Mtbb/cj1ED9WQpk9WhQeZ
5FYpsRk7QY8XKRIQZttBsboRkGt5K+dnGDB2JT3KXyga9EKOdlJrBdZuomMR7AgrV7v6URIdGhlH
tAyHM0rv9DfYJMydedBIc2QE2ti7qgT6jPkNOf9u955EN/zC/C8zAXqPARkkZ+DZNAgRh10k/Inh
nyq3NoEihFqG54CqWscWODAbe3q9JcwJ/bWfDYLxeufNo0MDP0jl1nQHoT5yYPVTd5Y9eBJ+dXtj
ZK2CP14qY1rWgLuz3un8VCqI6Bq3aAFmzgYOUYkf4XaAEX1BUn2elAFLa0x3n2sAgDvW3/3fRTxG
vyjrpU3GVtu1RHYIdpG6BNNKCZ51uMkpLsoz6GDMWp1U2et9CraJpc6ml1RgiXvGell0IEc6upLZ
tA6xsu2FFx/gtGeTz+2OnUZ1pS3EJbxz1eVQ70BDUowBKu+1aSv/Sabj3RwgBLOvO7n2NbdkQKKk
ng4jprNkZK0VFI2JolfxK18D2NAxqPmOy1CtOLxm4CCcxmwpchR6jrtkwwrlPM763gmZ+91tX3IX
aE4zNrpwFIH4VbPF7BrhfqzE5zcEFA/C03BehwIfmg9gDegaJFQZQv2cfpkSaWXDyA0T9nuxabDL
HJh4be4+Qo7YEpSE8JnhjM3J5W1zRh2YPSsMxtEh6yvaffD8ldbS15ogo+gNSgWixX4SwtU3AA01
44d3Kf/TDopJGPPbFVbknEMhlka+/qTaaUHCBfJwZNv5tW7VPRmwB1G0d442b2fLtJoNtiELT197
/9kAbcJRca4ZZoRZZTmDTanMwP4NXemafIZZxYwFw/oSnNXXkLVkDOcKzp5NLvtmjZI4mdj8h6Rw
Abo1BhiXg2zNkWJ7oiYJ8D/8gQGDKgwn8ST9pDlw3RTBQ+cj4zG2LgWx6mLLJrCk4RrPsdGD4k5l
37hK+B0RwjI78PNs9aixW10Xvd4YdrJu/GBxqto8XPGt/P/OrN/hVAwrCr42KHQpdNgw1pi7de4B
CCJhb/aXuoY8fKczCtlTd0nhU/7/pMz+khpPPhbGc7eNXcqLJRlfwwJABhroFF9mKoqqJfmqnaY4
ihG+5jgrtobR4++bqshZxa0WF8H0eqqLySKuiDz2ZyGiIlpr+6/8u897I5yPzmi7wh9Xb63/AuX+
Ooy5XK4suLDSreED2oLkhQjg7GeNBIhEhi5KcsmsOSQgtoJaIkRNwOw7qO3CBY9ICcFhnpqv0qMs
UOH3muVLu57/GaLIHXlg4x0hIArtU99nCncroEZzhuz6GCsUa+DDCBG4vosZle5nFSHBzw5HTbAI
My4XXQgG9afQ/sPHTu8MXbFs8MCJ1OnBFnSf0cpjLnHUV8iAi9sRchl7pzJj+GpvEC8wo0prX/hQ
c3zMqL3Hr3VSWan2aKVsYvCi6S9bzgTl8/n6MpOdDzFzrFtoCXRkclyl+LfAPgwmXcnlcbnq5osG
+tUlfSmlgcYcYf/cjhpTpJzVuXlVqIqU0C/XPriA4FVoMHvp/RW6+Ls4/kR4bEL1plx/npTfd3sC
V/rRrNyRRenvEqguUapQDS8prwiYLO3RmxY/gNlTwf8LnB7Ytv3ZA1nUO4PhwmqlpjjubX6OCfPU
8VsLvoqywiE1iWHlQhEHdOQybZfvTAd2KJ/Q9Pa1PAv0zEfVpYHlw4icA+fh92xZWik+nX3EaK2+
wsZtUENIpQ1H5gRCtKN21WP/dvCk6UCSFcLkYln1FGGJihSW5dBcsvLR4d1sdSobrCSPmqC/S5D3
cedfVUHqSG9DBExCI0WkT1SnVXbCvwy3As0Dn3l+RT+X6x61x+B6Kh13Xp940/4ID/JCffVltqIg
JQWOiEWBs5/FyptAEufqBrJlR+MrV9q0EvfLlGmV10j7v7dsI4KxbDCWuh0DTee6p4ZFS0slaBaH
sn5zEV5beB6Pjq7XewXwv4isjfpQXRjypqdwfcoFOPqupstT2TXEqme9EQOdazvDu+zS/oDWRKgt
go+g11Bc9kRxGXpEBYlsAyF7DwoBXS0O5tG+KIjmoAtbaedbcCkEStVnN4sNwVm01tMB2AU2vm5i
meis4fQO/FN3cI6TDCireJmBRVs2GyPZJVDXJPD+2qvndRfxjw70SFPsuWe2rxuNp7DXb22FW9pU
8hzypuJPdr8m6rmeBD9i8e//UP9hslHAwOl0WvIQzFyLfs72+yDWZTqt22R5xyavO73BDfboOH/0
9WQmHIbjlY6hC6hKWqb8DCaF1W5tm5wa5LzVwUXkbhLaBaspSPB4+MhsT5zK4N+Ps+jGAQlbSwbn
9Li48jTG7zMQBBui2VfeiwDNtPXFtwEfOkUg7W9kqZT4ZP+sLcMF1l77D3BmczE/rzNbjaiLg2ro
Z8ceXHxqoWBxaHUj+MK1P5dZRsfFHtVbtpW8nDin7hpzU2+nQtd2nHrWhuvIc6bnLNy1ILdAYuFN
aHgaP08dlE92ZCw90Z4apMi1gfHONMNulriO6z3hWzGwBwE1Asfy72jCYEphLY6y25uzpc1BoDNs
1wiOjtBT0PcONEbh4GpQ0bgT2Oi+GTVq9ylYf4zHFkEdVcfOgKV2R/4Fp5gwjrubQZMKYxplmzdn
USQghDEIvzEV+Pk/GY7ennqzwOpxnW8j+9uE2KpXHCSglDVlxNOtzkkU1ygMBMJzzH9F/NP3fe3p
X1nTLygbkbPEmgJL1k9hI1H2aLu5IxRokJX/Uf8DQf9mmC6GYxVV+ktSkCPHM/Gl/NwnH2fRqDoG
QG9iPqZAop27fNFgaGdIQJaNzMg2H8sXO6bzJ13pXp4tHtB0mU3/LZ0qwMvwp9J+CexBYIk0/n2n
iS2e9MwK8oiLrheBN2Ez+twfEEV/rgxjwVImHq40kPSEv1AE1Ei+GMzJvLxhy3/QpJvgjau+kHT4
J/Z9197E6ztU/PcCnyXPTSYfPBmF4dY2FpuFZ39MYxoegqfbxsrdR4wO90ekPHtelahQV9kYTtuz
oYjWXob8Vg82kUCxmQ2vKBfA9IU6p2GTHj422FrkbO1qQVYfUA60tn/MTB8t0QqW/tiHItKU7E8S
nJwSWiarvPHPOJwJjldYTts1eLAVblI9A2mB1J2Sudqp460NxWSfKiuQ4gPKZLzdl/7g54Cf3SCc
zN8OOAyJlsU1Srz57WpCO5J5Ytk1BJjt7vbXvqzigP9nv5sudveoEwWaBii0Si3ECEbU2mBrcTMF
+lL2MO5N39HOaq5mlkW+GK1ElVfAFCEq1iSxpZM0yQJE6xoCrV99usoTK/xiuTPFxpySWO00lYjn
WQKcGHZn6J+1yJjvFUlPrX5AqsWHyJDP10h3pEI/IhYUpjn7AG48MdO7uRmUq0G/1Skcux1LWkNQ
ebrbpRFD91b07uSxJ/FrRAp8ptwE0AKbOeZ8u18RoSoCM7+FghQnRt/CWXrzqjJfkNTxsiE89pu3
PaCDUsOAbsbUqJbS9PqaQcTczaEqCl0iRHXgFdnMLeXQyfPtQn/OhidcTal08eet5GfP+rOZ+4FO
AIolua8FnvuRRPtCgMky6jYIjPEmezntFdZY51LzkMxTriW2MLGOB0X/5zkD/Y0bN3G1sKZ3I2MD
HH/XIuSVKtKdCI5Imfo+0pVvP2xosyQfgOeAHDTcmHupsmOBpaHbmIn9cX5sGwhgYBm9bNc9ZwCZ
VsWsZJu2lt9hZT9q2DlgpxS62KorNEVmt2ox7o69XRbItWa2+5BikuqW6YRDCKtb5sPTuyr4ebRw
AMVY4FBbB0n/mPNX0pvvoJO+8UylhkKhoXYia/r75xt774jRDYIy+3kKJLCodZVd6QrJru2tQAUO
9SG+Rw7DjbVW8F5gK0kgx/qHJ5b9Od58Eab0rDMN910LQqva1+t92WgIKp1oSoGfVuAFTTdn8oFv
HEUOZGzlsbhH+GbshZM4ai00mPX7mSc+JDQXaAAvhOdga7vGnW/7+JBAeoEp318sC4A9ghJfyO+Y
fslwb5O5WP+W/JLulHYTIVRTW0tXsyJQAAO0EDfVjljfJQavs3OPlRN20KKITolLh4RYJ6TLcFGW
0v+5o7KkTxHHbyiLdeRwdWEQrkacVPwtweK8pZ4ovk9RFUPVybjBtc7V9TNnWWlKnwr4oo7XbBuH
9vkXeAjON6Kbz74PCGq7axjGYvlP6e7FQqRBq9jFQ7HWEmDNtYHFJ8QSx2S2drZV3OzwG/NsH8oZ
hdR/XVjtdr328NvCblWdgwsZ93o+WqtSjmv6JfhB+7DdeSYe6WCX7QDZ6qGmOWtQ61JXdrncnJtA
dSnaAfZOfu7jDPkE8v7R99ex3F4Ntu6klF6QLC0oJDuNhuh65IeEVZdNvrorZhZ0t3sjctVyjCnc
IB+gB7SgJgDeGb0Ogu5Vd0XVNPkQNHwB48O/UNyyYhp3lls1QMIzEW6nnnLVeJwovIVHig7PXyuh
LeEzkBoUHVtl6zMpc81yEbRvLHLAwNk/PKJzwD3xXZbDdoRGaupfGOC9GhwZNb4a1g5gXhemnMYP
2/AZddK/tZeSEWZI9IcCALcdUSpicVswmRY+5ful65jUKsbd7dK+vh8SPyYOL3tEHvGU6ciLTvdV
YtZk9pdFiNpQ+k8/s8LjWoTnVkoeIZsgT0sWm0AujvRHaaoDHwNpdN41yWGkSc2mJQOpuAL4FNOT
5rcervbwTauOxhjqIlktJBHUeTExr85wjnIYuix8IJAxQ4xypF3yMwatgf7tZiDYTSskSdT2Dy5v
OnLZ9Wwd+FdU488jFA4GRYMuNlS6iMBiNG3Fr7XFab/OUWm80Bk8CLofp0c3dKuM1OZ5KeJPrSN9
KjgAs80zoljLJASk/1RyGBOqV+QjkTnXPu+PJbXABnBMcMHkqcyvjThtdb5MbJ0VuP1Voie7QXXL
9Tv4Lt95Gva8nutgKjMooFn67TDUhfrWhTBohDu8HVwYhqE6iqowRcbD69mNqPi+jOGhntjc7RoI
eQeWmtuh0XDLJ8sfJa4nhWKOh/5H7CdXnZ87DhOZ0dDJY4AV/dXScKdj6wQ9N7N54qNxh+f+yf1N
5iOydEQXI48KoI6H6vUgaaDT9Zz+wio5cK+VINuJcwduCqzB6m7PMb/WVeXFuRK+zDNfMMSMxoBC
7aJwvNbhm6rp7iD2hyNdveJ704iCj+oNv8/nXE6PjbhReLbcFnDaPRSX0wm3GUu3mmktkdSkKODd
DaBo9aocAj6evpldK/5fuj9R9fnz7HjvtM7GwQqYZiXIWlHr2s8gjaq8cwZzp0kwWbp5BQY7R0k9
paNCJVeEyZxTiofgP0O5FWkAM6BkghsZtsKwixRaJDZadnUUxCVj5l/PxQrGiW7tKKqiXK28qJEN
yEShUzMqeZpY9SG3OSYdvG/sqlV2UI3xo2bDPv9qLEjH39cPP+GN7XIQGje4X67vQcYfNdQFEqFu
oA5qkX5xLkK80mH9z3/90dXA7t9T/9AdjInUIj9+jAX8pgycu4RTqgkCloJpcrPkGcv/0k3o0zXz
bwtC4Q7JFRKsSC9dl/zgFxOcr0Qk/9ujZbHtYnIC+8d0dpqhB5whKG0PMbvsM8aFim6q+0vTyTq3
FH/bA7JpyRcaEWJ9x7ZeKo0pLn+gyIEtAjxYXIT/Rv5slV6ZwNwx3o0jeRRtRJ9gGCwbJQCqAKtT
GHm1ggTEFrhFuV9aGWUFgtDrdx2mvVPeSUzkNy6iW2nAK0LWaXTY1EZqocnL4p5pwe+thFTBEoWA
F4L85EXRPMdxsuGL+G1TgsP/uBuDwrsL/hACI+X0Soo1iESan3eqJ55REIZ6z8k6i2QaLsN1gE24
lTO7LYCOmHeAnWPCBDrWSbKuhGvkE4RZhpRDQ7jIsgfKDuHJyCo7BFaDR7SO96cwr4uzfUCUNXSf
bScxhLI6TiP5WncTX/QuTIHjGG9fEIMglHrbAIB4gjZ38MH6fs7Zn7f6kWr/nFP9i4x+lD23rety
qd/VNOcI26CHOErRQmu4OgpgxR6kpXIo5ODxBISMJCa4DOex7Suz5BKsYa+efFFD6Q8J6AlgI6Ie
2Mr4zkHPNh1+7Wf4LCkecP9xD1GGIMcgId9+bX6A5Kww6o4lqQKfhcyu/X4zOnikIneTukbM5Iv7
gyNrRMQOSL6Dcxyv6TcIhyNQXAHI8p1QsoY/8X6+WksgO6NuITjCuoAiI0nVuKed9yKy+RztnG31
DLalZuuTidr2zied4GTTHF8FV/ArAt1AvFiAhVFRl5Qm0ESa+nC/4fgroQb91sRizKTiQP1q2+JK
LwffwVTdpVfsn0aasvTbH+pVouIcmIk0OcPjNGpTCiwX9hNOdNL+FSZGJvoCPEOYR3CwDBH9Yhw9
p1+GQpaRUKIu23y+3/7XcbvsQoN7vpE0uWTMq/KrL/MxUpb8bNc0w7RQVAz7J2qcXeaUPIb3eYfe
sWD/5vIrsx98UqHROQmzWSWYYluoWytbB3+CwXjrv30oJ/lqXxE3rqwQUFAdVcUSXEVW9wRoC0Ub
3Wm3bwaby1JJaw0ZdY6U+QXMd08H0sXBdJsCV397ffhGyRwaYIYocR0y50d/29h0eHJWL06JPL0b
KAIIquS9jpCyWEdzxxHjxk1Abc+mUqyzwXxgDIV/RyDH9EWN/HYE3loZaJ4z5TNP55qTCqYdadIb
yVCyOu6lB8dTDSpme7ymRE+ULcQsFXNwl8ayqLOdspJb+GQJ38cT0uRqpG+ps6pH84fX9VFXLzN+
W9Wwa/KYmJxZr6yMPD3VUKRnL6QB5wergpx8FGPSDSeW6e+cxGKZl1e4cRMrV4EyJmu9qpOsdE3a
O4YN6I9T9jCvXnjoLvJfWfsYh9skXxUWqNtw4/eNeOTnbJ/rdQZwAev98jGzED8XGHsKJQDPf1Hf
AdXq7WQZkZ+SI5pcstLRjOXsQRMQtKNnVccaSw0+eurX6UyFTlTXMh+VS39drQIzJrnAJPznRpzq
nHXRDBtOYi804L/1vA+sryHB+ZFXzSezpf3eDqgg2QB37qq24Z7+ZBVKVdw5Z06PRQIbaqnP7Hqk
QR0US9O8eXZsVKKKnAjOIMbRgAAHv8AMx263B0Ahi/E6IxaZq5+IVO8OaayPP1/zdcm9FEqv/xIU
83ABp+VQqFRnauWgXts1soUxL0BmHRQgiU+BIhcJYWTy6kcUna7V9R/u1rouyCfXG3KBKePI6Jg1
hX2kjCApAfApdUnkmiVQcRBCAyMAslkkO/GVNcLGzZmZ6/jFiE2icq9y9Mo//HuK7vT572Rmtfuf
ebudy2uQsP1FVytO31cgtrBxmp7DiOabLEmf+UyQnVNJNdSymhdkplvU3/suCnio7BIiZzTn0yy2
B2RdmDNF2PONGrEpJBPFWckauW4Bo9mhFCoonBrzC600MydSQFIshbX8qqJKfLSmRmwRGyiHDMjk
WuXIPF6fX0/LPP3Gl6qLGzUmuB/NP8Swm1PejXpTVmlXzsL54ghs/b9VU39DmIQonUtQwJIVkx+s
YkGPJ8XsmKjmc7Jr2YZ5GwxmTU/CMxli9LJ9+arkxGOmoMj2TCaMRGcUpyZPFxoaNgsefV9h1oYC
++UtJ3yhUnpKh1AfZTe3Ta6Cxp/vmieIV2Y14SWrpQs3ZQdJatk9eO+0Us71yMhhghlc7TIWRwRZ
crY95azhHPNpECdGd4ZEicIcRF59Wl1Z4m2xPEiyPg8e/iJsCghcD9Z+Cg7TEb7zzo7BK30cBL+a
ZNsfu7WPtiO4J5hXs1Ac12Rqqxgl5n6net2Gz8GG2wm4n0xY0B9zYzFrHWLg3B30AjX8MCdWqXvt
C7NwCs0x4lbu5WJtfB99vkRgBqvJJXjtanBKPa19gI+lo7ZWmHMLBEUpQTEYNSByICw5Z6u3Zlq6
w0nMuIci2o+IpmQ7OvxnUi0mBtGrSzVXMQaYoeuucZJdzHAoWpYAqQAMv0MpuE1iKbusez5vw4lb
DBOLhH7OH0QqoV3R4BHy2t/GO3vmmxv9ZlyJuEDSns7cx68wJlMcniLcH+Ed0rnVQvk4TBQVCxsT
oYVGXlOcr4nJVZC6E+xzIYWWB/gOHjy8iDisDlIRImfdj+lcl+VBStcWiYLfSwajGeMEHQdUA4F7
pESppZ0N2ldLcENiMyw9b/4XwZkV0HFZE6D/dmVEk7jgYeRy0a7fVXBjFzU483i7gOeUooaYSKby
v8TGtu0wGvXKlhk3SrMW88IXFjtjx6noJeWILQwE9fL6sfmMBwzVdrmFBKelZn0Lc4vJriSBTwx4
x7XQ/62dpy9ogZrLxzLw4dm5S2ze0zYFenK8mO8/0m8cKwjIwMpFjcybswuN+QrPaosVylAWbKQj
ZBlGI9bHEXWFv9qosFK3WxSUB8/vwyIMQirjQaISM36xO0VE9aDpduzaxsmbOS8iNgSV7FkqNvxB
cOojWwRZKRsE7/3F+Fl1g/8wmytcZVFxB8fPurP6nMimEgpEVXRrmfxG/FxyJZzqzwFzMYCJEn+b
JDDEKEybvNEYvcBkMKxF+jM9RCYDgeMJcCZ+4OfsCuFp9cU3Djhk0DkkiIaBEojsxDrqAcBPAjPR
FsOMWBn4pYETuSw7MDjuK1gaYVHjCMpP32m2qV7Cr0MbERr+4jF9DNSbzIJQSaKdJAcPYaereg8+
3MTQbqwuZaTPPjIyasgtjvxtwJtL6qdBzq9rQjVXIJwTUqlh8rCHIiUOgPWWHfIS1mWMVYGfnusD
IdG6lz9TZ5I+8JS7FPSll6snPrmdqoDD0urOuUDGWW/jNvsIdJNpXxbnQ9RygNdMtw/6owb99yBF
5tx1ACrSlatMps6CWpQwsPoyGsmYTOs98VAwB5G9AC17030Cj25zW4CR3vXjtUzL0kcV9ZCKmmqQ
0uj7XFPgISdFb1Zg+/PI+3Znro1k7dIN8fwuD4dejxXFOuZMJblSYaP8cyfzMbB7Yu8IS3y3Q1C1
P27lcQoTfXReawliSI+ltJwmKPQdwRdPT5ATkjnsf8YP0CjWhM8qaQ97S/+AQyZzxfkumQio5HBH
1+E3o2rJgBhm+uazvk8i+JFVvrUpb00w8YpX3qZyNm30umSf5fDcD0lz1gL7+cSLAMR4yR43RDL8
QZ78ISQfeMknbV9DU621Gr6AKvvStZ5YdYvIIK6XWBZ5inJ5ss8cXQ7rOvD9ADTdw44HnRFcU0V4
HEaGZUPA9TyrjDbLsxDVYoYaIqwr6W4BCTNgYsstoi0cOFmCCvfSOkZtwIDlTKZ+lBf7ggJDJ1Xg
gi5H+wIQds5gQZxkZB/jdk6D7BXgdrqcUJsSE5slGiAOPw3IW6NcCfN7OBk7kPngHXkF/4kR1XiK
iHc91Ea/qW4+pZFWzEDBXhj7P2aJntIo1G2bdFXVbVImd7rW68UDGRw3pTenfrvDZW7obdz/yI49
svIelYW/o1/KRTfCsNOBMYIBMj9gmacHsf+Dp3mzhUAuzSMbF98yHezkPr5ugCqnTmAhJfCgLgwv
KjIWJVd2MHTun81t8SfJLrcdg3vgSY5NytYS8PDlWjG9fD/ti4QQ1bQmFoCWxmJRx0S8NAZmu8TZ
6BFvfWFf4alzMiAUWVG9ab8nHloJnCn88d3OxRPssA6Er2U2wUSFZujnrPbeOI7MlTLwl719awO4
K3sWmhYWK6CNwRLc98C3CeWesbs+QfzAs9dggYBcLiX5yca6IAYfZUFgIfgJEaX+vB5Q5XKr7OqZ
ScfWL/ZkZsDH7Jmg4iUCjBh6us3o7fpWP43jyToVbu09IZ1W7vzhXY5ftgTy8rzTpNN6XOzAMqG9
/c+HG+hBzHCADu/MARy7q/9nlI5nVLHZGYcBIaCd+YTuJ1df40pIRFCxHDLEqiOdJtkUK6UQnrZw
3SDktX+zv26RGWBIXCsdlyM2QHXXOltp+ySrLfTnqfgTXUOGuqog3mUmdabaYEZHSkUuop7BYvvc
k1ez0Eh6y6eUXKMNOdTwBRlgbsoXM/9kVOHlHRGVgjQYg6czEJXAQMXFVx7vnNjut8J/O+oBE9zd
l65BMZUv25KkpcWCpyjsg15gvAWXGfUwiFishs7dYzQExHJtnwyJ5oUZcKtMjhRs9giFa/2I5W5F
IGK0HqFuvR1F14k1OaaeFLYyHpSTG0zClDTiPOIFGO86Rt2DBkxAKyDzGo9PND2d4AENVuNYb0a+
K3EjR9Le4wTcE2iUo/Z5d7v7D+viMhqvXbhNzIzCKujAvcgfNsEbQ9OWfuWff2+PsYso22pSWm3b
dhrsuMREnxsikk3aoRyky234SqtNZ24lR6Xbk2oJ7aXdVW/U6AARNc/Z11IyKTIuDwj+srVzic1j
jP62d1Mnjcy+uGlbvkpW2nDSFGcYw5AT5AMGmUkC4x751H1CryMbuh4VTz+NxmWe3crN0O5ZXxaB
GpIrY90S1PqKdxI7YhDd01r/CBX8Sb8z2+nXeTKq7gc0XrhwL4O5EJ3pILF9nYvxBJegd30GLgaE
wfaWux0H8CvtMJEIlPeCzvNLcpDI/ZW429t5PzCdpitV8UVMLm1Z6rG2ESEDSuHPn1jdtVgN+RzT
xWGNxzS8ja92bwKNKTZ9ys6ASDoyvuuB/lRGIyyF/tH0K+NkQ3f1OGSJ2GBiR43AVXVIVC+UiNLO
MeN0SRTr7Fbjqd7Z2FuM6sh813EMXLLl3/QW3Jtcg/oovP5h7iR1HMHXh5N52GZq7jw51JCBff4x
OuKeqosDUZizz8ByCygzyGJW9jYxC3TymkVoeHzzibvT98od3g5Hl5sbZCNlhuqgMYeyEBnr6oB/
+f7XbZHoawbxRZdbLyUOtsIUinPiAMADueCMj/6rlvqaCx9KVxTeKiSihUpjRvOHsaovB35THnXe
g8ocVpTj3pPWqQOHRRWXtorC9ZD3kNCL6FnyakJgvOQ24TyKDM5Cd0XaAvkU1jYpKEVzPjCQg2JS
fVkJiZ5pD2KhUX9I5e1tWWuR4UFNB5if3OF0cY73TORiOMaLxCvOQLEuxXE65kMlrF8TFt4Hmp93
vW/icCN2RXD7rQU0Wt+p9+olPoflCPQbrXTPNGOsk0ajpcvHjcahfCQDkQeQ49rGONIenvP8zRtv
VUz+7vuPbALoU6ly5tkAOxuJ4v4iLoI3nODqtY1fTwLaaf0ECS6GHuGyIZhn83cWhahoRqRN5ZWL
tMPnBukuQlFONSoa1MaQwdu1wB0u/oj39SigWJDJGsgGdurJJFag4j8YqzhUkZVvkrikV7LzxJ2r
InIfpzVRIah3Xj24EXDMu9lbxty9AfvJB/8J/4XwvUbbY6Bm/JmyyxLXKb8dJNTbXWrAV6rgOHAu
mRRUp8mdSD/qQ78NrFy4zxpC+lIJvEYqS8bVyiCyI9glW0dtDT1uGJ4AUAlxqUzVhLmCOrdIP02c
EDip4f1RI0paooYOK95RGY73DiFEWobN18STLW1H6nsxmOZCt4uRqujVK9/rBcQYixeLoR9Xrk8o
HKVexp9a1vL5c8H2F5SwD5wWPJHAqnmF/FXwFE676QQ4DaAAx7lJUkc/kA0HUhWHr45AMU0nVQSV
3yiDAtqBxtCEZ43Vp3qFmHl1lDSJo3vj3Ek3W0xkSzS1rpqNSZ0s0mEWmdNgLON1yZdAm7dSWyE1
mD4TzTkyG8Ten/eBXd2GoaZ6hiF/yYOZopwWBi+lLd7Gaf508S2tV7pr0/PA2oPJzrbkOBshDxnQ
mja1gsOvKP0ZyW0sMCmE1Avt5KwvksV2kxdmQ+d+MEaKJ4smDIAMAgBkiw7k+P0WxPterX4k2VsL
8FHG7fZRhT0b+/Io0CevayIvqSn0yIggup26apjKFRpRPMzACAwb2A5n9pHXU7zG0MuZfOqf3Ym0
+JdwxL79hembCy8AyLy2w2II7N5eg30ti2yoD1+zDYFVan/L/LBHYFlXYFX/t2fAyjezDoGBnzrG
KFUYRXB11H7jkfXkjNH3YLX7N88OfWOyNvJ/SEsdRQX8Ft3VC+A7H6zBmbfgVKg65885jJiF2ott
RQgp+HVUWTW1NRkdLe1gsluM99IhQ408flww6ZtJI1C9Ub9J/eNKmSL/yG9T4+P1RGz6FhKS1+1K
cHizRhpoSgiMJ+niNyMjdckYKyrcDXKhkRpmaZjqTm4YJHLKIWa1ICQH5RAdIogvmPsjvnMa3CqP
HICQ4ZnJuv6DSzd3nCDLH2ozCDJIOjASwbliT6MhTwXDUtcg1qBtgTi6LUxJjkKuK/oZDt7LM/8N
/C4eIY3MOXlAlmWyf4NseWdkwzBKlpPTVg0hCHF5V+k/5x3FB7A58ZLlPzIexRKulFeM5+872VXH
PSC3ooLHqVohnlP2UzOuHPiluSB0Sf5i3NrhEZdn7SG0AL8XBtM0RETI0ISbK3y3F5SFfwA7RVvd
6VmCemy3PB+iJyRvJ4Akg5WryUEZesKngC7yV4hdzoJdeR7oXgxcVlM8i2itzafUY8NPDWYoqqD2
Jh45eZwVB8XOcwKVuJM1lEVrxeLwRj7ZXylrKqzYt1sImlqgIDKaYvuSanr+5cKUwbL5F6l1kfyJ
aJgndn4XzjwY/0YqntvmMkuBNHUIjXd5HMVXH29gfpXVwiUpSLyLZ7zu/GzEpr4UVObLRc9f+u7/
bINLmQMstrEQirqV28NytJZ7zwRlLgnaHQKpcvTpfyrb0Zr34gPw0jIJZCEL5LWP/6wqXb+koi0b
XJTTGBOpb81poc+72qvZfgrAXt3sH6AvL0oU4BF9JE1m8gBneUXHEN+DcnJMlpgdCeS7RC7LXdnN
d1cqgWpQf6XXRsoM7gxl2Bl0ve/D8DrP+qSwv2c5Kw00qHa50SP3QtMURFiNP2eAo1tZggy/VWtR
BvK2eD0euZki23p27EP+U3Q3b1J9QstXZ5DqDP/MhgpnbXYVux8DA5JQ2GcZYw5sm63foj6uj/9q
dB1zPMeSqyAZQROI0o0DBrdRvAVGWh7vYwqXpyCeNFCu1HQhBJrVVNBFJTW43T8yWGRM5x4QDjwv
y8eNKs3fMwf++IxEwEuetRCoagvpyZ3SmlKTzHx9E2zJlCaToOGDGZzFvqMn4TnUvuCge15KCHTM
94XrYTGvM9ZjFBS1968poetxs16FKpfPaup7Nd2d91uEuKQrJRN8KWxkf3M/PdCPlPnYDQligT3U
OVHrtrspO3uEwmzHVU+n1SJw+nsSFr/oPRXAOWiXmIGoOam7IWJzBuImk2IVczH4CLLUVWVaVyEG
8GhzP0A/MmgXlODyUdZWdK/FmxXM91JgEOUMldU2ItqDDa8X4P8e3XlTlnivppTpHsj8ZOLyPyRE
kNioJEhMfz1kkqP6Oa6J4SIP3Qfa6pC36qNTAuxOBesPq4DFqzS/v+jG5gPVSY4p8exmor+XbQQL
9HsKaZnq821/hBc27UATMoETQvPJpsawUjz1btJ7xDYZbkKwHPMt5y+6HIM7FDsLm8J8I7CavQb0
YHg0eQrVYebSOE+hKNwQ+mkGZsM9VvB9+/6ixek/WBueZSd/dFZrKEXqeCNZxM6alccCXYqwymOd
g9jsSfSMF0t9E0cnVjqeQbnPb3CK0zYAlFoNNXhyn1ljVm782YQkM2NCfP6lJRqNmux+imtkOIL2
9HhZAyZhkJgofMYYAzjmkoSolKz7BjXEQznkaX/G7GmgHMvhdPwbYVdCBfNw3Zs2au8lpd7V+Rzo
sN7U7Vh7fZ/lI0VfhL3pWoijc0LJM/NkO7moZU+dZCslim0v5eLN3IBo5Lkem1jrlMqBxNl2qXVt
gMeKiN7IQ1fbwAB7AJgqpAcTE3sNCWQEb83MEKUXk2TlnuVi6+NlRpTZA8Wb29hh5wiRQQhzyFnu
WaL1K1fJOeS2sEzZ62eASV2Qf4yBGVY2heufMrZV2LMELtSeF2iTP42LnyfEAvNA0RgMmlKrOBPv
NUgNfwaKtFzx8kgVus8OVix8XoUSVTJxtck04YGVCRyuP7PpauZmYAIy7lOYf5zMwgXUVLDOQmay
WVTfJ8PhrPozxpHMb7qacZ6WqqiQuzz8u6sSOwOtdSqJ2MouhkFZvqhXeav1dqBQgQhOxtWpPUn1
i6jl0I7thwNCSSmAUE+N6kHW/0XRoMEsco41Dmou4AHGiUjOO4KH+Lmng4La7zIFDNyD4rhTPDSM
mSXIiQvtvyjfBdVjbwYUBs5xjDqjDFMT7WV0pwvTKdBy5TwzxATnKo+EeBK8sJhm6KM/zP/ANzxA
oF+1zcJjvonL+Xahwp6ge6nDRLrcn2FGQz8urANiy5Fk/Qe8UQpseiimpD1X+Mi1bEdZGLosqlEz
SHxIMYx1oZT016Ad8L0htHHk/OJOoN4xyUoUayf9qISsOGWMyekZkowUUbkA7MM26NVM8l6UWwBl
EKbryUY8n/pttSUuLamcsV8U/pve0ILDepQwoeRgaR81KKmim3cOnjkvQARh9RYNX3/PLXwT4w01
CkSC/uIv9cfdgG9U/KSsQvifa/tuWzeYkTOrxBFJRuKfvEoR6qrxHZlFyhiUwlsAr/nM6WZp1YKL
Yc1cQINJTdH3U1TPYZHUG+t+Xi3tZQ5k9lhahADIBZ/QHidgJqGI9YryiSpjZ8TNHOvLPrsYVim7
kCtlvJWAMWy92ggXhQJ4KMHzmHnwfXy3uFARfw9ii6WEk6Z4AyKp4rUosOklZmyaN804yDoqLAfu
tVgnnTYCLG+wa2I8XvvODbc1azJKGQ29q0/8KSgOVVZ3j0pCIa+Y0+jtC9ZJP2mJyUCAx7702+r0
L6EF/eYfqR+OyMp2oP3gYUsUNfxiHot+TXh5lQpInPaIl5H+Vj71VwZKw7RVGDbEn9f9TlFIYOqU
vzDO93vBKlXCyvVRdQQkeE6of05RwIHIyrD28rSxxkD4tTpt1sXbUZ60iXO0bvIFB7/hvHVWzp0l
BYyM1Jh+IlzLnM0FuaBfyJsyt0g+xwzUT6tNokXrIgpJ9WBn2E7PPWr0G38et0a4CAvseD/8Mvdf
PpkgKzIWY5ybHDLXBt3yIF9fU6whEQpF08c9pUWAegv4m5qUdRVzX44T9d1BvI05AwzRIFlkMxHf
SJdCMvzHLL/1Qs3myGrONJPSfjB/RjC+jCYmB2buoUtLZ3j6lZaFkW/yQJz2evHVIk8nUVQGH4Em
I6ktHhi5bLKdBiBRd6CrY6bfUEinkWqZVC9U+JPQmuX/37SU2AaDi8/onX7U7Ok8wq8b1wo1kAWD
W1DJnMLoldNrWMD/yUiqlTpBHcqUktMI/XNX7jHTjr+C30atSsy1uYdAtJtqAdVKE9w64DsudcQN
8h9IQ5Y9nkcx63Y+xwd3DrHyL+3+eKzpSL64PCx0QoVy0DPIoYLwvCfvAvjLDdOaiNDP7wjMmnE6
GeJbECzrk46fo5/YXCgpdTnw9Xy1QvqXhju4MwdI1V6UmJWEw/nI4uACWhzLNz4cui0WA36tCmcK
PDqjR8lzefoaIqvGMbRzaBxL0OzjHC2BTjMUW4Z7qrBWZ/JaRm5Qqhju6mP/jHdE11YA4fyM7GJn
6aJWWHYenp5wPRpydh+p8BR00zGlMpdz7MJLJnauSa4hsei2SSPVS/bIHPmW1Pvw4McUXhjCfKQx
PX0wN354PY85koJeGDKjkfRMQZ9ZRmKtIy0IgpqlK1ezBVpXZ1uteaJ1fbPbo3FhE8MDKVnPzqwP
MjdGrnImQ6MmLsbIUDGS02WBxzGgXmMkgQCjVKI90D5Dx+lmby2AO2nXRgbJnc6q++wRgNawNbHW
zAr93irPrG112FPnof16Kt8gl3FAF3ZLPBX9bTHCkIqIS2FcDjX1CQ7Zn/YPM6KpHewUOrLCoAKW
tNg0qKagAcwGLsBIuKeghl7jOIU9KM/ND74F15d+gWP1VoeIKIKJsdmVpUr8XSKegDkLbU+dsaVz
e3uQz1XzX3a+rtxXBPUD4dSLTL7+EO2c1nahQTCItDuCj2zdaZuyZ0/iER8ep1rl2USuNXCQ7h4S
ZoJBjc/WRZXEWE8rR9glKKO0aAGVrsCIw0WYiIsN8ZVp4zBPefZIhU9Z03jYxPiEKjYapFk3D9Ks
P9/uob9m/zstZ9RokXt5++St176sPAvDK1W/6eBe/CsDbvfhW0/B4qpun5MqUeKhmjft2oR62Rxz
Bp7gCs+57FFFXYf5+ZOh4OzQPR8z4jpj95mamNahF8jiRYmb3X5CdifycpsDeLu2o6HLseBQt7CA
rwbMQuPi06SpXLSjhJQ7HVFce6iROdk7eUDBBCLyhJwWMTou3vR47egC9IUT2PXQjKWl1TF43o4p
Usrhij1o0O0Z4acd0qRtgVhF9CA037xsYdmMTtWPlDV2Gsi/3Y0cOoTncTUgXecg/Aewi+dpo1ly
s+SKHAbOMms/MgwMsFTQrZbaYHAqCxUQY7mUal3allfjt00X8FKHuDM966YAeeLViYoUCFCBBJNQ
kKbGbHZNY1RAcaHKV6asXG++ruvjy2WxO9QjQ/Vxg/HPXwlqSWox7U/fSk2t4vH2c5kGF0gTCMEh
KLmCbfJB7Yq8AGr5Lj6C/10OXyqenh44ufKg9ut+LcCusgzJtGSr0N+LJdmfVP9hyM5p5cg2AK+g
jTVSnDvw1qdEQocpR7J13kcMBPRKSm+JphZXZQcJmRJtOwbfeDmiH5ZGvBVK0Rk24TZY8/1gCotR
GP/nI11q9yLms2ybkLljljI5UnTpkacKF7CuU5rTRYK7JfYtGnAnzbnp4Qwbv67GlUaT4sReim9B
IzXJLZDBBr0K5ztcRNgQrPmoo3NDYaYyI4Lw7KTWicX6ao3n0Taj8uhCvHhGppS0o/ZPvMp6BIs6
VY3ks5hlPtWJqY0+QH9gglJGZJpKjAUzCqOkdjNfBI8y4/Awjn+UEOwToXLSn4FdenKb7HDYnlow
aMHgKSoooivtW5iVhtJuW/5RhuUFKtoP/SOdEo9qxsOGLojhZ54Bc4x1pFDHFiS9DfsRAnKauZ73
AVoLdxeyihd8T/w1bBjsDalf+qQD++eIWBa8fYli08BPj5foMwUfrjZ6cTS4HOu7B77GckPj0KpK
zdNjTuiaPDE5COorzlUNkO1d8IOmaQ+wTt4RN7TswwbwRn6munWyPaTE8RkPiA4veOAJXWQlOOD6
iT/LXTYSCR56x9Tjm/itmenSTLVtw3UU+dqB16BFIYd5BdSuOtF30/7RkMtXg+oniCYC+JjaqDVO
tCe1RUb8Y3NluEBXDNC1UUE9pbiXLxMfnSD0xYzL7U3WIR5sdloCh0upZhtaeGfwTw+8TsHGorUq
vGXTBMK/n9XPJR3BAAcu83T31+evthiO7QV3xFnBnDS1MIeFclYXqozkg0u4yfj+d4kQEAAmG1SL
F8PXmQ2P9PqJF+pYUFjnJqwmauk1pdP7KB/sEoNTsDCyF1ESYAr9kU/oLZIsedhg+jSG28Q/DSqK
LltyGDigozcCqdAg8XH903cVgFj5sv0PIoZVMmb5E265FnaKFyIXeW5pIkfjPbGZFc0MCEWlNo8b
1CgT5D7TyS8lmPA0Lca2ZzJjtA1/IEGKT1bhxtayeKpOMtn74AkMDGc7NNLt8VuUJsZcVgSVCjUx
S1w6kcSGQgt9fYEL9mGvdo6wW1dBr7syklBLKVWi08JJ6hYiGp3g8un0ICpqQdPMox1pWD1Ims2c
PCbOos5i/utMWTNE5w5SjdpuzO/SBggs8PRrL0IV5nlgE9yZ314iibqyu85lDn/8bvx6+GoBCVaW
fUKahc+jgJ5wq6KYVSkveaif1tTyuAbfF7pmQ1vxyUJc1a//vrNAw90tzgUQnvFjuTLfZhO41TJW
scmB4qvud2W2/CB0ATbHzLb2IUbmC3GD46e+2UViWqafbeqrHkmiBfToFhyVr5aPtnm7w7K8dBy3
qBmFAo0kxRADY734yqEzuVf86+XbThyhFS3ryo0YPRLWs/jFAjj5GMnM75JLkaeKGSljArU1j7wP
3gFU1dGfr7N6dVG96eScgxFUuiManSDqwterCby4pAZpK8J6RlR7rxQeVt0wdyubJYBI5yanB8Oe
aeMA9rkHhVCT96lxDkfK8T8j5qKcB961TIjnsnBQhzpVT7do+TgofLzUEXKhNNVQlW//xENe1TP/
HlhG/4rgmIpSaW0bQFBgRTK/6uizHohF3IfTsr5e3TEp91T4egWa7K/lTxVKuc8nDqLQmIGtu8Qg
G9EDD2hveORrOMLlawBqlCM3dtlXhyKlIXJYkkBdamNg8onUbscN9AsGiBKCTZQ540xq2gPGq1UX
H1Dc28cziBJygCmIXM0Fr055RZlMlgVGo7gCQY2mloCsUFcbhA9PHAvbkPJLY0fQZfmQj4ueI6j/
vaWCZhVIZi9CIT9xqdrYuWfPJclHzt5CbqLDPAgsxF28Mw31x+W5FBZTTisYYQoiFEEYcuoby6s2
fo/8Y/ZNHUBshGkDKv6HHepVI2+KwJ8BCsViJhEmSaPAQmTw+VFLG2Uvrr92NsYyMiaaXSgyYWiu
N8MpQd/LhbOhNy80/ParHlPpc+lybuUUHJ6Q+OZcNSzxMmCaNCFNLkQfJSUtIEXsKYdsZa3D6IbX
FByQxb7fEPu4EOrHvKV6hqxKozrJChhBgi6E89odLu8wYWGr7dUUSUO7ltaXRxdXLBDgnydMxVu6
uBoLxHnEhiE8AIk4rz1saKzYb7WOyir+iwRty6htqNVz+8uz+HOWdhHKCcONIZlprAqWzqbKiGK3
tLDkK0hqcrus75QquxfmzxJLNk3lYxuiKxel7bEj9vR1lomk/R4FSXXJzKqo+yGrY8VYJ3ZSHzcD
n63QBxyw/JkjerafefzxLmXMO4KhWIyw3fqZf46aR4Z5XKHrYdfAwn7XeyeoIqufQjO4QeXXhw3N
2fhvcstA303xKv4FTbyX3R4aPkPRXwPvnVIb7TpmOt79qTh5quWetpMVfNS8T3yM//cQ8Nk0C0rP
hDQyhQmxFE3SpzFGhbjZrgNDkD2Xu4A6otSuJ8ouQLAjyDEwdQxG464Nz1iIB20wI01Fii4pcsMo
1/s79k+Ad0+x+c0hqaE5kZrWO401SnYu9S+KBUlec5ghk22g26fxRyCO471d/SUGVzS8WlS0qi30
0a+y3xSwA6r97uwm8hXtCXQJyb0fI5lUbqtbQ55wYUkle/mY+wNQRQiwgXJPr/2cfKoPzwOH8ML7
nDhlLAVwqgdAPo/CnqTl7x6K1Lrx5ViJWjMbqLK9ggH8BPkqqj5QVq/7nJj79+9w0yHEOTmWka55
GQeF6Wnwp+JTpEPzIVaoygFdnXAOIJdtRESMJQ/ola8w6hmzshRdLacstmfPZsH84UHuRClvMewy
j3A9uKrQln5yoAc6Twk8CZGTMLuE7q/e2TUUyJ8mDVNzqdlIJVStWHfezExioPsPIEW7SgoBcWgm
MaD8ckYZiblpmoUATvNkZQVydPQeQzMP1OZv/CMe0MOValFk99ZnjLpGb7cDfnx1HE7nSLbr3P2E
ieC+HCw1VVFcadestTbbUj6OyT0M8CKrh8yhse71y2UFiVLDUAQoHSsxDSUq3Bgc3PNAcq6wsf7B
Lnjw6GxTYG4pD9Jx8mOd5mWbJ6ma1r/xI6x9Vh2SQZs3vVXglVUPWXFt+HIMOQPFzjyoVW7JuY44
r7G2hYHyoxKjgzxDgdvhkQCaV8FkF5BUQ/dtNow4hjM3O9yuM8fBolkvH37Cw0ccc2aJ+TtKJ1DO
YR/b0D6lHO+/fsV8eyC17hYb++T+mEJOhZTSvnaqx0ZYHNmlDkgzjOFcnfxhSrLO2VlyyBedX1nb
ncG+o//grCJv5rP7bISbkEFJicrnzo2Hp/nJXGCuSm+jz3RxjkLLqPO/XschJD82L48G91yUhctd
dddODEyKcjYQLPuh3IHHeRsmLFkkumuATg7BLTnhmzoxxiD++Jp+nsw71JhkiFK6uB60Z3UfIKj5
4cc1y/V8oLnO7wsquPUPCqZGQhuJSCwdSed/Zfbb8zLoBjnY+B2dfq29HC5WHAI7r8asmXvGhXgZ
6N0MlD7wwEAWgA7SRKPtVMKZwyjvPCce9Fr6LoVS4AVUAnZkTlXof74A/a2zSL4OC9EfozFAmtrc
Eb2b4kmbObAraX7EAr0DwBHYMBpq2p3FQAxnC1uvdnI4560a8fG9eSAH/ahd1Htas5KQdR5TaBIZ
6p5cDJspu3VlVvzFeqQeq/nS/IHTEgId92bGNggGQlrwNs4zUUHZWFGg4Y1nt0Qw4RIRMGJz3LzD
cGuMXSJP5kVAQKcsCOG8fT6TcXkO87I7fwwHUC0YSUxJq0zosmR6AkD7hYbO9Ozz0YVmPv2DWjxH
taraWGMaR4MTYh9dNZw3vJvFDBcw3zL/R26wc1omvlWLkF1DlC0TRTC17K8LV8YNr8Zlr1X1BXuV
5OtmAucNnAEmcGFu8E+M7/wX6aq2kWPetIxCbHkFhkPgijCYAE+vL66G+v7oqEA0TT143y/oRBzm
qX8Lr5jF+rnRztPXzD/lTNBTXU5V93QDkj9mLq7v7UwkD5wl9fb+pcXOGurL3DgfLOrY4iCLZT5g
Zegz6wMomtRJC3M6aZqrmjA14XH1SntNN2mrBuTDQRf2IIgZ72pwQGxllce1DQRB39IDRaXiyWjM
Zaafn+Ifnk5MNonmoXWqVA9HeBD1KkJmKkH8ZEygBIDDCIL7N1REpSfJpX1HCKrzrmU7/djVSgJH
3voUCIcbtul6YcXtnNdV+uRTcAezKwJ0T2asdxjSfLY63+CUxqaimEJKRM+TwIOXiOSeUA2EC8Fr
Fb960XrouC8PRjgvoHUdEqSx/2F6eOqdaMjAG48tnHdrzPq9i7b0Ho72fX4QNwpAHMteTmDNlKaL
FXslg53HynevygV/Gu/RSgzmRzHndIZ2oyZY3avPqRrP/H9mZy6L1KFSmrxV2o/w+J7TYY2fZQRh
vnZdL9mHb4kMsZNRypsKq8PCu2hiRcvZGQEdlznnFwQz6owiX/uBY7syeqfZZP6BmQSHc1SZkfh2
r1U5fsaVLm8IANvC287bk6lO0TrdaPeM536TJypkMTV0qgMHA72harJucdF5L82iM0yiP3giF7ar
FK9LVGq7wV5jtJ0VZ9KVv1ShHTN31Mf4IW1zna2feLZ3vnpGKIQc4z3+ZyAJ3LVKGSvivG+fFzuA
YM2ZI3yrQPO882zVfpXgCgNL5i1Xvv3xmxA8/Wp8wmXu1E3bCjlefyUtDQwPYh9hyDLtpNaWE71z
6qbN/iJktbY6CRk+di1auYCbTFlrSgh99OOMLsqPAqPQtF01nIUyN3nBflkjTXfbcnMmHEpmKRGS
t5GJRsi4FFjmEy/l9qB3mFA+bgjlV7GkWMjeEYjv+HQRZZuKbgJEdFNMBIepohAbmmY5ZB3Ng4FG
2jnDu3uqVr4JqjJoH+mH2pyUGUS44uQl4+bhwBEszC2zJJa6NSoQmJs1UEAS52A4QW4mj/BSsMqq
eVR5YZuu5GrIsfK8uItiFL/VqWUP4imhCvb9P+CPFVamw/Axw5bzX66DDzPU6Xeb0cy2dD+kzudW
5REaAg571OnbgEaLqOj0hexK0mZHrplVmx6yJombsOw/ilCNUL+a3EA3/eAZGnKdz+LuhdyKAOGA
L2rpn0L879Xtemd8K7z518oDYtWm/gv/LllqXHXgApbioR3ptYU4GfQkOPLD60xmkUB/0G7Bydpz
/ZqjCKXj0maUz05X7Hj4+n68RoU5NAkwmAVUg5ki94XDwdooaT7Nn7KJV6ih5eDwtPOAJR/Mbxa1
sD0Pv+fAx2wHpxSOt0lsKNIsr4i6bbgqja9avYXCEHsgii0fSbVviXSLwwWKZNC/uPuZeeWL+j/4
/p7M/LxlhTVecpTE4u08u0Egx8tiVTTKFglMCM0+un8ZAu8Udcjikf5JwF0Yb4Sf+fWxH+stIjL8
TQicBazUZHiSBGZH2MFYidHb6x8YbBRdHuFPh/JOidP2Pk6HXQeK3ukCpV9nsL0U4ONt00jnCSUJ
060bXLuJbJrmfAAbswVGav4Xk2Bkm2qtYzBlMKYPpWTtZc2lH+AlbFCrQMtVDvEFSeL2By8JGCBo
g/vSRBDc0c4Kz19OqXVFQ8TFf17K8koP3sTeWgAuQ7hTc5KtSxHafrGLM24RKQMxQes/OYEoZcJM
G8RktAs0H+D2eBvqgwChSofkTu0fNhOT21b6uwrZx4N61fmev5bTBal3CnyrpYid8HoX9fchjooG
9bdB/NbJSi8y8JfFOt0HBIUcuFvZBmHbc227ieFF8no028R+1d0Ktu/R7aJT/VQxOhFJh7cM4341
oIrj49HJ6zyhIAis2E4tYCttfyeZw7VnOK8YnAI9MzYKL2MjAPvyb8z9jXOG3V+lSMyy98LVxigY
mMZTEhx//oDQV16TenOjlj24d15F2bwr3y5rnDesI/KjJXRR1zYDj3E6Md0/GKjIPx0ZGcLPokfm
NmBUf7skLWhVbkctNEyi2FepoKKG3xhBddqMGLBoHRhVurgBW89gqDt/91YLTRn7elRUvuXfz28Y
yL7JEzWNVY+/LRBlGgyIS0cz3Zmna9J1bNi1icr+l8RmTNT6/+c4sFKG0pHvZInFBL3yl5qthWEL
S8RiMwIgW7CWhh0y5C1RvK4bSixKuXy6jq+KlljYwDcZwyBE0pGd7sMIoiVBMyOOTquarhqcX+AO
lgickuZn9iyDK1DXuL0/lC6ILwRUjg3vyzJbQSQQhqUf8tF8Q/D3+tR1WlRVTtLv6rYgVrSSabXz
58Iv9TH80GzFeQL0y50pewKVShX4F8/5ltN7fM4/FydXiALtF81mSHC0JtKvlMkWYEByzBfHJfep
l3vpbPNndJcpIOAH74MktoqcOVcs6MuPedk5BR4ecQPLc11TPiBuJ6U8cKBDr1pEm3k4wByZ+4NQ
dXyZ5nFR10o7jKgEt78er9dlcgIdjA0jmMA2ysnLaa/Jurtm3JNeF70QxFnVokcQ+OF1xOMWn9Bt
D0xDHlkHNZGAY4lgrT8xTkuwr9Z/0HtzSPQACNikgn6Ji1Pnr5NDdJcwXzI0PP0xw1kcBXDcu5zt
tGgI45O5o3fDJ8LE2Q+khaS9ioJech4AblB7J1qdWM97+rg/ISMihNY7/4Kxf2QR7R9d++vjsgLT
gP4hePl+RBZy1OAR8lRAAAbuM/APQd2W/rAjNXT87Qekl3bk5QPBGuCgaGX2XCh4+JU4JL4DKYPN
n/cp+eb1hV0OK8m2EwtJtM7Mp7h7rvUlAhATunAHklY+LaxIKp8Zt1XykKccXNiDS0abLfx4BRdl
MVOuFGxVsUnfBEQNAjKucJ9iA5c/wN5iv+WaGngWe4kLQX+b7m/dPJEC6iR5pjUu34E03CgTTxnb
QbfpDSFtkYJaZYHM70lcPV6SgK+Zth+bkg+R2XL8p0IMM3HRH6PkGjjach51CTtLj3ClxnuEPrgy
Nlc1Orc66BwdY89FI4+DKxjQDFtysvQMCTi/qqQKVmLeOHo/Yqapox3gfLhflzWO82IwdG2+fKLF
wk25wGyeToxNXCeGNQHnyEVaZZ+cL6gLa/jSf3yyqb81dbX2wsZfyEuifWUiZSKM9y4IeHxArmbU
+KsZGO+CZmLwdmLXHxzAg69X4T+dikfQ2zwy3RfjJ+oT1H9IZyGNUD1k1/Q6Blhrc0d2nwilCN6A
i399G78rdbXB1WfQTFdYf36t0Y+lHaH15yqriT3ZI7Nn1Ygv7InSH3HJKr/x2613/vnfYNe/QLXZ
W2yARTNfD3ZB3IBHCygBLLnd8wmpALNg/z49BCQDebRqyft2snE9WIwhJjEn1hqrRbUlMX6G7fEI
EmEx11RRcSSUeOXpZA4n9Mk3uz3mJmqb46YV04uduLNXen/3WF8Go7zVv6On6teFfzVZCUEuFq1S
/pJsfJtwp4GIGd6rglDqY5XoVKPUjvUhy1VFXAf2OV+RbPNLFvJUKHggs0D0KoGnynLcjca55zR2
Ft5n26MkQUNiAzia0nY3Mk7kHT5T1NBrGdvHfuJTmGk1cAi8Qm5jlXrwd40Tz6RGpxBLC3x1zKi0
GoQsI6kFFwtN4jiw2Do3Qtr6co4KbzzPzUSuY3VzmfKx2JKVkW/LLWAWl4J+O8Zrhgn2mBmhWLxe
YNqLrlPccqoNQab4BmMWUKojL6KMD6Ji8aoDxzyCNrT+Nupl4HI1uEXmfOhFH6dSogeJoCUuu9cQ
DjoCTJZNRaoYzbSVSvUKmxQQBTfJ6mH7EAPVxe4BN2YpxP81OMgNk6nNBaefMKQs3e9tlbuNfmgC
bttLEMUC8rPt5wpjpXZdJp9Sln/RTDKVlkYU6vY7GkGvFBEGvSqvMiAMxizbt0Gd7q1wm+Tc+9qi
duexPesMV6K59nI9Y9SG7w1WnIIox/SPc2D/QmzcSsm6vpZq+jrICm/HMlwFZk7X2jWq6Gq8TPk2
vVipsVnP6WG3N/mLSoLlHvydEbjnFNVxsO+innMiCVWNKHfLbPJIAhX934aZ1jgby45G4lSNrwqH
k+pAtmECjCOxqKB83kmnJjFYwsjogiOvGezgT1I27QHcZrUOAAttNJpZW3kp+vOessLtI16ItSei
4JHpQRv8tTizbpLjANSilLZ8gYgN9wptxEdl1f1yx3jciGwHcF1+sogxnFTUGrEdK4Z9FGVjxjiK
Y7lFFjjrsL47bkuA7Yu0TNDKn5HNS9Qt/2tQLxbVgVO5Vr/0zutvwfvbvOGHRySvtnoAsby5oxdZ
3Df/nXDf4T9UujsGb/cWhZeDFbrMZtCv8Iih+P+2QxWgMqLnwtNSNq1FMMw552exehcP2XuDW/Wo
fGcfxfjQEt5Yn4ngXzMe6/FjRWNh5M3LJ69mtubJPP+DaG42OaFU66UXUVRPvUZ5I42M80R+9vJ/
iaj4tli/RyOqBjslx2NBOZOHyR3s0WIKWW97D6Am0/MV4AszZJg7ogxTThQKr/9xsRtzRahlXrrw
YmKmU+SsNN4lwW0x+sl+UwBKSATFbxL8jmnmL7IBZ46VHCj+kxXcPc/03tjjKuwGplCnS20MvC28
9uwL2EBwbocL4THmZ21ZS10Rt8Ru5nq4riMPb97tAw55iMcgByF7s+vey9QSpU41qAEnSw7ULh9b
mizRb9I4wTUVYjjznH/DydcbplFHixl0gr17r9H62GfcHGyyOPKS9UzzYd7vYaiZoaog1RukCbuX
2PHU60Kpse7CZRk7BCNHA5i4KBLcGNkn/w9oT2nrMa6fFwx0PavA4PT72s469CiqolkFNA+FwM7F
HfA69OjT1VpNv5il/qfpF3UK6oWr2gMVFvw5vXwGfXPA5CBPmI4H/tjG36bzNPzZUdy2sQ7jJlES
voHAO/8ZPYPsNdeVbfcyQh6T2oV9a9meN9lgn7I1EHf0S7UVKZRTEj91foJMCS6MPuphKscDWhsL
Zbq5eEz+TM+MnlMZqmmKDR1/tgiy6KiD4/obOUrBtvQpQhhuDb4eEIbBqlCw0k1DeNGJY3cGJepH
XMjmEBW2YcuyvlP3Rpf6iydjdaOsZEM03g8Vg6yGDTJxjuphdxyVYbo2m3iyd35yCANlj+1VQ3ZG
rsHWbuQp616//3EeA0vZe5jSAkbVFC5Ks80XGkh1biuXclKN+VkPHw/TE6AGuW+A8z+Q7poPqtj9
pW3oE9l7PQcEdlpxM2g3gf730NkCTsh7CfFgVoM+8IvJSR4DC/8Rp+8yZoCRwFYhOC2YCXTGgp8U
cKetxXx950WmY8faFca/gb0xKhUrac1ls6jRDVCM8aRdmA6cvNsVOYLTGyGdKVHiCeM7sZUVICBJ
u4kQVEjC+a56s0ZcsgZdEFIa0bxJqwbOZ74pzKcxPFhj+kAmI/fQ5OHGxrZSW2sz8U70PCHoYta1
aQbvCTsV4NU1c0Ahe+8Yc44V7O+isG8e2LUJ3DoK9vHGQkMeV10imJDiXT1GyPCEpCnLnRkaL5bR
AOtALTNRRHbrMeoGLQuE2WWHzjOMS3ppRRrVHySRv8K2NsDlf0jvtNGr55ZxM3qFDTFyuo/pB9sl
2opEAX/XMdK8z4euexqmtgaJDWKoitc6CxVCoN0b+etkrLgxuw/OI/JvAOZXT3sO61nZk7kuiePW
N1OWanPDj28r2wSKkn55IDGFKkguUHFhGDH0rThG4A9WEGL3KFsKCJ+U5qgD0A9VbndTXlbspQFA
n17542f511CHv3tZV9JJ0ZpwL1zD35C9Mwf4vKb5lT8pPd9xeR6GQ63t2eGjMWUKFmtrQeFZzUzk
2ZgtUkYxDgZsUY/VRVIE1Dx2u/u4SA6l5t8ciZmBQ2HZZaMBHovk6HUCFPju5XySZZtHRso/UqOV
XqV50yKv9Sw8T1wJ5Dh82r4cY+2lo16k40t2k+vQI0YaIUCjbiYylATMOq33zHEEY9swzS9Ef5tM
rctdvkDxHWvZRsINCzmNk7SEkv/c1Wlck6ivDGsDw7go3uvBALV14J1yhqgwlHamqFgmve8/iW3U
NcN8GKwo8odI4PIriBjB2LiMQ3UU3RQcV/O4FiKHGnl9QUytMwPQPypthesCgNth+0e4GGdSo/Ug
uHyltMhbs4nyfUTrcnIadVOiM1r7gm0yx99CBWRomq22xJuvmQGKIfQnO94M7L1hEpryuGiXqaj0
A0XlEZSSCOLCfW7JYugDM5WY/J68aW5hcTDTWTunH2sd5radtQvRSha0hFdcPs/E5oV+YQHGQaAn
S2QEzv4zgaxsVYp97u/pMZP0s+nMcLM7NO7+Ecb7arqOtOpIiCQw43pqiqXg98ptBJbjwej5XwA8
OFNcBe+8GcB/BOyZt0cGHgTisbzqzEFQG+3rblun4JjtzmdI48BPeQrqKZu91CLatT5LryljtdKH
JtWkbO+2UcCBJLCm+OGC1TJIQN9wDCfvzIFhjqMrqgVlqmKzXnZXzUJ2wSQ+89wDziUMRpi1Z5Np
AEgICbcnPR6xSOi8sPJ/IuA8m+I2wAmVyk1TrXIDx1QZ7xIBOI1DRizEdzCemBiod1lTMxXga9rU
N1JVPhkierVuQWYwChsUR0zgjibI1zuFLU/4ApPvnvKwHkk024707LGYVORxZJtyaxuaONndoePX
ATHodrI0fTJBAz2qknrMmxXfiXev3EbvaxKQMJ9CQazeKRHCdxGyIF4Hui9tO1LhWg76gJk0bvsB
5Bm/pWfjvI2Ah8XFJRG3K0u8kxBN8GONV442rT1nG/Q5vj51DH2lQfd5pKG13ncj9gLrXZVBsogj
uDTW6KRkoUaupDrW3ki+rm40D8JQ3ODv1MaaL70pefbJtr4cq4KcBIdHHLB2NwRreEnkyExPtLmY
7FmExlp3rkGtUllrXlfx734H25aVlFuRpU4VkwThwsk8nw6XtkmYvPpsOb+YRJ1eI7bqIfkqyFiZ
ZNJJC0/KmXOjhMl0vtgs7BLwkYiJk4fJFCQT74NkeGSJymUNz8Gdlz4agijZIqBQRkcawr+1Z8O1
7p2CdMCLtxBXSWXmtdmOy7dLuDYtV9o89Np2pXe+7VAz5DhJ1N7ChvG01Sufm5uZD68E/An7jd3s
ErsSHgaLZrD5/SQdnwiJuhNcfpy8pFaXiyNuBlmF+hmvf0MkcT0ZeceoKWXTmKhUtV4UzToqBn71
wLf2zqL8oAUZPPqsako4H9a9Po0brdRcSyAKTlpOgXgz
`protect end_protected

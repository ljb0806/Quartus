��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��YN��C({r��E��v�ɣݯ��бM8���^M�Փ�K�9�aK���O���F�����".{s���8&�\|[����i���_�Ish�FX��L���:��Ȋ2)���G�i���=x�`�l�~X�O,�ڟ��;P�|�)7��0M�݄�6�X���!s���x��zrq/�i�Я9�TX�ؒ���C.��Z�{:���Q��-h݇ğ�c�iR��7�� (�ll�'�)��C���&i
�e
%��~K�$r{dv��Mu��X&�,>q9~��~W6;��ޢ�#�`����G����z���W�{�/��{��H�,�D\��i]�=����v2"��:�-�|�����Y��I<�B��W5���U��i�zR���K��d.�NDZ9Q��}b#�
�
\rc
c�΃2!�A�o܆�`7�P���t,�$(3�*ZL$ñ韚k��hd��vj4u�VW����Gڦ�̰,�d��,�b�H)[�P�Q�I����Z]�Y�)�=>LtP�iQ��Ҳ�V}͞��b<��՚���c��mF�p��Y�J�t*�����9��,�rX��5�����K�q5��z�ͦ��	��~������k�&uP
���*$vL�݇��:�<��w	�ߚ�	�j���R��5�+�[hH���)�=bI���-����-�4�{i�G��y����ڞ :�y����Kpc���X�gz���}F�qK�"2�/�'p�*�;��M^�D�}Ҹ���#�@dd����Ӌ��Q�{�^��Y~eXw+��
ݶI�l���<km���/��W�1��=	Eiw�t�ʴ�<��u��A�}S�c�@��.���w��I� ��H����� ���W�!C��:�w�?j���f	[�����
�T���ZX���Ҟ������|Ql�a�woWM�Y�������դz��-�~����V����0
�쩦�#BlwE�k��5�'��!8����=r�ʐ�sZ�
�5�����7s����VrI:xB
�����8]���I������=A
�gEKV|(�/�㕏�
,�4�t��*����=�lWsQ���
������4�"+KoJF"�
�i��3�-��'3�}��� \* �ذ�O�~¥ %�\�s��U�NI<[�[,9j����;*�\Y� R;�q�GYt���j�=�!�e�{���+�ay��	
O�{;�Z V �a� �F�_�����PE�Vs���Mb�=��2{Up����%�ѹVᵸtN� ����S�#��.�۾K�a��K��cN�Py��a����.t���e��c2[3�1����4�a5��܏��zP��p��N��eK�Ǧ�\ �n�k���d����0�}�:+�is,Go�)_PI1#��6�*<5B�=U(<�s�l�հ��?}�ԏ����po�d>s�r��P����^Nbl���??�ij"�ȏ V�����/�p.�#�Qx��@>c"#}$��C��s�����	�����5L��}�5̱�����	��$�u�Ey�F1
/:=9�B-���0�:Df��LO�!p��Y��y��ze��o��엓�cbqŏ���叀$�bY/�ʠ�B��"Q�����GqA����?0y�G���"�-�8�����V�f�\�Ih�1��G�ʲ�U5����#M��<�K���iALJ�4���g8�M��L� �,��Mi45�v���e;:s�o�D����V�Y��LS�3}�����cp��`	��*��qY�����g//���tO%�;?��|[�l�epX��J�����(3_�jaPT�ֻ��p�kI(�<ı��[t�Q�������5@��?��`������Z�#ױ����6�$b&�D�E��%ȑѶI�.�ӓ�YT�#��&��Ȩ1��ƐU_���c`�(��y=��m�Bqg����ĒMӈ5
�*x�ox�<Ɖ%�� ���*��@��S�.�G��7�*���v�8�dI3�?~`����Y�)�>?�UV7-����R��`�p0�X��S�]�#��f[|��ڎkTj�m���[��26���;�2bj��jI=R�9�����F��u�`�?��\/��󯢶�W�n�8b�� ��6N��ir ��5O�S���y˱����?�F	��բ!�k7O��կ	[��x���E �RiO�bwvD�A�S����>��ȕK�f�J66���=�H�� ��@gfP �*����Ù+��o��G�
�W0��7[ã�rR���U��jy������8O����5z��(vE�&g��g�(�ٛ�2�3�{��
�X����Z��0�`[��=�J���m[��U<l��g������wP�v0��Z�R�+�v�L"��m��'�i���~z��(��8�>ci~rl(_��bI/�=�������N��8��q��FLOO�e�QR:����9׼`��{ �4%��e�3�O<N������&X��[.�/g"�=���Ƽ�����x��\���NS�"`����M�kp��X�KbD�C;�Q�Cl�3�~R_^,�.A�l����2�*hՕDJ-�X���L����5�)	p��9�}vI�y�͑�����6�F3���L�����74Nk+V@����.��9�D6J��w���w	Y��]����h��VIT�vc���aD/���:&G�O/}D��9%�U^�Ŗ%���?�p}��2�����A#��ovTB�_C*���;&b��n~�,%p_u�˟܎ &̗��'<M�J��X2��$�J��$�y�i�\�ct�Q�������1���ݚ���;:M�zxSǘ]������ӘQ/�q����u��qRY�5��'`���l��|��u�|=B�lս�P��X�~Q���
����S^c<��:��sN�28�'ZNzR��?ɯ������O����z��z��=����|��H���b��Z1�>Պ�!Z��p*>^�멽R	bL���	�0^���B�t���,��s��ר�R��M�ߋ�Jb��i����W
p��k&'�v����\������A�O��S=1�ֻ�;65�!���8���N��_N�� ���N?����RI�U+B�Z���r���lq�ogr�a<�oT�b�,I�Z�uFw�ɴ�ő����m�8σԻ�����s�UfP���Y���h�F-%߶]1w�f$�{b_8��=�"�Ԙ��#P':%�צ5�Fa*�E8����K�%w��n���tE���\arh�7�Q�B��l�@[Uz�w�rC�OPĳ�}C}'�ӊ�/Y�����A�7� Vޑx,�A�!�ҷ�3ϝMT��[*��4`V�l���rJ;�(��}S��˙��HzRG���w���)V��1�L����Y���7Z���[���P(r���.A�{��g�F���C!5|�h�:�.M����u�Y��%��Ʈ�.hÙA�*�m���Oj�,��n����?{�+OR������J�f�,�$�5&1�����"��� ��x�$ʄ�Ov�� �-�-�R�;����YP�0�JR�ɮ`fq���R���P�Fz������Д���v�]۷%�4�c��}�����8�+X�H���Aap���G+�	.�D<��~lM�:A/t7[H�p����֗pG�*,��q��o�"�.7Y�:�ngH �Wj)���?�S�Z?ν ��#�!e������4�%������G�0��+F�鱓���'˂����xя�v�V�C3�V�)G� �B<2�7$�[�����-�=<�<�dU��kqf�i4� �1�P4|=��9�Ϭ�ޠLc��Z�yƢ `�;���!Q��I�C8]�]篼9�}��;�-8KP�^o�8�
�N��e~����y�gJ�PD&qU����7����CC��v�(r/G�HH��~��� }N �60�:Q��U��3�C�A7��Zn�<״�����z�TH8E&���T�P�t:X~t� ��!�����}��X|�b8��0��Rڴ�(�~Qx�����#Sz#�u2�;��a�]e
����.$_�U��;��Q>�rKE��� �{�x�������2��>�VNEE��P�TQ.���#�\�t5�t�dd@?�i9��3���`��-�iGt�
��2�x�{����|�71)��S�-f�]6x��e�xJ�oh6�v���Z��옣w�R��A�fk��#�d�F�,�����(`\��r²`�뺦�4��h�D�E��#;�-w��������>��֊�ܫ��۹)�Le8O�r�O`������C�s�^^~VO�d?`f�)R���Qv1w�����K6];�seJ7DO��T!�����L$��8d@5�	���V�!�aL��#/h��kP���x!�,yj�8�'w8)t���}e�	���Pn-�eJn����Z�-�V �Z�/�!�a������5%>��e�9l!2r��F�1��$���ă�sh�m��GΙ�o.Au@(Pd?@�������a�2�x�������s}C��pnC��~N�bNe;� _$��o�����Ne��̌R��$"Q�z�i��h:C�)^sJ��*ź#x���$X��M��K�2�bd�k�;1+_H=��/��P�0���y�+)Y��Z�U���UK� \�J�«ə~)\fl���Ka��&�> �X��C�D��K�*@c�*�f���Tk�����n�Sh��\���;}y�S�8䤁���R��&ܷ�O�-+{��r�(Fm	K�/_�D?_��*�l4�n�+�֌�������S�e[j�g�S.�H1,K~�u�;],�Mҫ%�)9�Z�EjY�g�׾�x� V�i��5ަ Z���C0Ӓ�d���+� bU2�8�n�u@��?���5$M/��9��1������w���6�a-��Nk�,��_��m���ﾃL��]�|�i��Oq�kf@_BQv��ǁJ36�(E���� ;!L�?�����a��$���#6�����*~�Ǖ��?#�Y���{\{��[��ʁ����w��vx��H8Y�+*Y�@$Ќ���	�ɟPЋ��&�H�G'���\���y��\�M)��!x��E��: ��V�_q���b杊aN�;ؤS��wO7_�(bu����I��T+�X}�Q�}��0b�4��/�U�kǟ0�3y�p�Eނ��	Z\h��>/����ʹ���&o��	՞��z�Y%����!M�$��^��I�?�Ã�,,��n9\�{+O��^X�M��U9�5&�!���B�P7�H`�P�nd>wx���J�O �e�G���Otݟ-0�k�%P��97��9��HV ���F��d��6��k�����I0518)�~�,)|�NcsT!��8�����<�рc�nV�L�J D%��;�R�ʱS�����<���%|��o ��|�ʨϖ�@�����W�S�_o6iϗ�L��+�XC��nF��3��+ݦS>�7}ڨ3�B��9�l��\�&zG_����{M�9g?�,��Q�Wm�+�Ԥ����1�������܎:t�G_�q��V0EI]6�u(6��EX��o[� x��R��:���T��IT���V�ஈ��]���=���IE@ٍ[�
h@� ��4 CS�����(�z�>���As��i`�!�%��;g>�[զ��PY��fbBB�vٵ�=Q�����ь���i�/հX��������� tjt�4�J������}�:�I��>�!��ps�v�&F�g�4q�m �:Q�ȱ �����-��@������{ �"��$o� �מ0�b�]�uC/.�f[����
L������Æ�`2`�M�4�������+���ه�6�H�9ګb�
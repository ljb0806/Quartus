-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OJz/ADc90FC7Xi+vCbt7qjMyVIS+5JZedtcqAZsAWxoyn7xDAxMn5r4VEzw3Fx8PqApEK8RcH7Rp
EZkLSiTuMt9x1rWGDdNjLuaSd0jrTi9Vv/7+lW6R7DCIVCwnz90/AAl7WTKrTeBwpkdxFDuSZsmF
BPcpBoZToVWPuHpumdZvVErvfyA4rnse60w9MVYCbW6fntwgewPPP1OSeXcxgymWC+8CY6ORIf9G
m0jxEi2iaBit3FUW/a8g8bJwQsXpnQ3wf5LrpyzGFB1dAaHT5T+x3ygFTFyypEGF3nO39x54WvAg
XR00zuCiYnjevEj0al05RHuMmIpbgJWSss88+w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
wLh3BaCLAiaaHZheHM/+56HZYvNfhOUzgCKgkQTGwb4NgI4KrtYlqsbyUV/JOH2Vu/ojMu5sjuUg
LA0jmBwgud4taoWqA4vgAjEi8SZb4dRgwqb5L0R/P84fM5lgXQMmt/QcDPEiyFVdq9OzJzTLnQuK
b0L53KVNW3uX3qhdKRTFStQGhnvTb/UgKET8IEXyoX3clAdZAvsVm4KqlVEKcFFdYzGNy9N8TDoF
VYbkZkWDB5Or20AVKcK70iAU+bM9b6BEBy8okaxyEJeI1tllOIYxnJpephTLN/2I87KWBfxDLokZ
OlEojFO2VI6gr/3Tq6nJCJyKKV0GI6kiKyXx1XWzyugDH3tMfOpzBpi/kJXlqGyJTa8BunASF1QU
JA3MCV3JrWRTXJ9BmDb5yV0cTTAYqGo6qrUZ/eD4HANecq4NOr9EDoXHZnsKxCmmIVCNLm4migP7
sFtZ4c7NgeyOHmdYay1m21kopf3RbNLMv8sw0zs5fPrbsHb/Hitj3v21L9jfx4KvUqglcht5+l6s
tCNLhpiRrDMwvCe2LaVd4PPD8A4zIXcuIeKH/IYEl59jJVK5lucylAao/g2DUFkuWAMJH3aywzNo
rv0pgT09/Ha1zOiYZlluC0JiC7vlG75ifjxtY7uhcawIjXsFA2t4rP/cwckWbWUa6M73W6IYjbip
KZZGMSahSmx4hEEtwoekNUuaV8jIlHwRSPXi9siyusSGGfoa1sj5EDSZ/ieZEOwNaL4bAtCQKiQE
MXsD2nyHIl2v0h37zUtaX6RzHuHMKVlmssuVQwIzQ/a6gNdZ3oCUwPcMjcv/YglvCiXKh5uDOXEx
QUZEEtSnYxrhnyEZqhWYiDwsUQCxUifH/A2vfPWGWZhELI4UlF0ibUHEy6ac/i7aGXelG+PaDVGY
kyPyAKemYXS8054p0KgP6yzVNz2jYU87/eeU38+8igFW3BNl7m9G1apymvc0e8UfmIBPVH7b/nlH
H8I58xmn1sdIsyjKb+YGZ4BoShJEaCiUC5EnmVHUx7GC0LEOk+OOckuCyNpa0QwY1S/afum760ER
gtsCBG8r9wbOqucpiBeAH3VOW0UiBxj4F1KRIY1ZIwDjX1vxMOWRRO86KnNRusRFJSvTIGVSc0bM
HGkR44wku2HhMXHhZhNdBHl3QW3zM1C642uYNrSORU6KJt0NaYVx9S3b8tF3480mz3h8j1txLsy7
RrN84dRv23En39vINKWg0DV7GUo16eG/vS0EtT4jLflFn9BR/AcYdbm4dP0D+4scNK24cZ/qbVne
RKsdB767vD4RmMhBMoitvxR1ck2TyjG9fbktqx9m5Od6/CTV8aUuqsRAyjcr8rlPIT9ftbT2rwrB
tqpR3UBIwmi72ZPi35BynA7haNHGLBzOMNzJPQU78lG0gn7pabvDDWcN3oOt4k8x18NqEI3aA1QN
rm8MN8Dpn4U/eO2u7VsVN5wCCL5vnzyi1J1WBivibO1at6ppP/KFVSxKev+gVkXppr/aB5Dar/1P
1PTVshVWVXWmop3sSeNK3InamoerklCIHF3lk4Vm3MrzYX/+51EXe8iqDhBEBLACDm7y7+Bd/SG0
D4HeHG/14fUFOkOalj+Pe9oIhDgUy+7EanYYjgJ+sqfwZsle344jXD6+FV89XhdNBJalo5SNutRZ
eaTIGdZKoFL9zdVJ8MIydzpICCn3livr86f1pPb6tgoBhFdvMgjSFP0mDCfgjAt0fy3LC7XeVTC3
MBgD1AwAuuNXBhOflGrJ7DsIcHFT2uTCQ5sTG9jm9oJXR350YwVk+9dhyaIH/LQ3poW6xa4trNFD
Of/BIBr7jE3mh03e6tgUJFZCCisqAs/EQIarRZ6ziHEIKb+Un4JeB1B8u2OIw2O6CikBBRg+J2P0
xAhHHvYZ9ymEv5poW46G8bjMTB631L/d4VM+DTbgdURE6KDkUkR0L3aSnHKw+ggX2G9Kusqr4ju6
dWRjiZ5LWUo3F5ykj7/bHcvoVP+/Hg/7XJRsAfmlpnweBjrYFsZy02mIrKaHP2FX/2Zd1bejcCw6
0XFmDf/2a1zcm6B3+/DXZ/SnqYO3ELN/zdTrT7jcjmJLJCgj70iPrDbMnPTKfjZVWl9gxsZ6WzUP
Lad4wMl9xYDGe5L2zOt/Ei0Hyzd/mdiHpzVEbKNIsfJR+FP5KANZ+6XPhu1XcaM9cN79A/SzBSLC
j/fuFPJfQdxX5XlxwIemlEzBl2xKNXQiUI9EUyiy8LMgC8WLjt5eiUiH2BfbjNRbDGpyUnrkubgh
27InM35BzVUO2PZ0TJXK3LbJpAmGRkckGXrphdcPIyhE9CTzNQxhHl9NpON/tUI86/rq2SheRRAX
+L2CkthuhDKKLf/63H4YDRIN47NQqQe5Rfzh39KR/QfiTLhw7lMOc+tSLX4sGhHYlqRzXpkDDH28
yiuiOKCBfQKHGnCtIXnfHKZH5o8gi/0IbB5d1QHRc3D9QgZDJxRKPl1hXHTtYmmFfLVRXbm3F05u
sRlWAsJoykoL5h6m6XQbexd6e5SifVlrix2KGgCoCajqhhYnIDYJR3n/zC05/K4Uh1o623kNohY+
2BYJY4uFQmqPXM3CDRnGhiTmNZOrr94vE/HEMo9I6y3OMKfwHikrmkgXi26ief/UXjgThLRwZZ7u
B97FpMobPh0klfoleWRV7tjNJLrfzgUERp5mx6tOoj5mpK3mnXHDuMkcft7e9a/KqGmTSGKkj744
oPjqraFVp+DOumv+XJh2n9tBha5MWmc11L/+rWiuUVp1XENKxcCYKSg4Fn3qZ2WJxQHJ6OMi4DCY
5Gt7uqZg93oGIj1TkVVehNykaJ9XZO4hBX32TpA7mcfhpk7vGPQwZLwlagGryigxMwp15zAaqzU0
GcyRzigx0WkFe7W8HuJuFyLKuGD7+MkFm+0Ra5wxat017rE9xpe3XgaEigSdh8CYTfMfbw4i/KzV
vtqEXhX8cxxIWqZ3/IQ4h2LiHpJGBn3CCfCtlp+ENK8aJ2Iifbxp+bOFHowtqGsX9tuOSnaYcx+m
iG61DngpxuB+h/JXmbEprojzMhejCihB8nPAxQjf29okPcad1VzeYHXvait8k9k5Mq1rqomsEBrW
i/YQcY8NfT7pPwgDIMUoYi5Ch/Mb19ARi/GZUBVIBV/0ftabwEL1TDb9lw7UTL7HJWWnmLHE87fz
k6YACzf+3riDCerS1HexDHqI2N8jbSiXZRQ/tlF1Y1+9fNfSFPrp+eF0vhNAivpXJscpIuPntzI/
ZoCK8EDxFTujL0bbHaBoiDmDGYnEnsY3+ZhenXeC9qupRBiyUuyKdpYCbD0CM9ZJUzMhkIwr6HDu
XbViCeB7KNpB3wfJdn5r7v3LOr+et7l6F09eR+Zfcr+0GcTiZ49YKJONz6vf3IKfhuEAyytza/eR
TPyFVTCxFqh0Ecw2sWBgWAR9H6u6Eozbu3TwzXxdZRrbr3WKXTP26csVdH/mKPJv12YuUL1W+tAT
qJDm8oOSfTqyWAMHP5qZNKI62U2e4TR1MBB7yytk9lRTWJjSIzS3Fr5pScSKLlubo/Vw9oXAc3ST
x6nDiq9HZ5mkfcYoiRS2d2k+G9vBsXkE9TMp3jLnPEG1BsbA3v57oOCO90YfaNpbibOgrZRDZN9T
lqpBiH5pOw+CNwiM+ev7lOIbA9+2qJeaDQJ1qzhj2LT5uZH0xosCNkjCsGD+zgvpu1Pw0Ir/x+We
n6yyEklTTwh8cls1ny3yYZEz3XExjS67dqUgNayIqRJgvnuqTwJaU4lBVQFIlPLYrKHy50qp3Tew
s7uc7d+WnnUCCYzuzIN5aWvmEOD0n+4fAXqcR2L8nVjjUsW4QhTopwogjSwO5GbE0TKA113GMrPk
oviwUARgf2NLHzuqKzZYXi7gdJN+yOQx1T3jFmUHdoZPCMdIyIotBXzbpOrBUaANnUsIds5wJ/JV
0Xc9pdlqmKgExmhiRxg/1KwnS5EBTSr8O1dnzIKVVIXigtntOy/8tZOGSXNc21PcUOJ1d4EpXiCu
A9Xb3KhpPRdGnPZs71IdkLFEwUSzxoITCk+0a5MFt62CLCAHHcQ8MNNFOnMEbUWuq4GJZpp6i0dH
cKr5E73OBIjGtmzyZJv1ZN1OtLS2cgYn1XYKJErrllAs6wCZm6JWL2fL0OtGSZBFrEWhG427rZLJ
Gbm6jEhRqGDoxgyPqF+DCkb99tVh7HGsqib5dzsL1mbPIdKRjMFlCxsC/k8gJMHUuRi3UOOh4Tub
r3fjMGZmTEzoL/uorLfT/IaT3kgMCQ3fV0ATewqfgACq0GYEK4H4kIf7hngqMLcz2BkcOIOc4Ybc
jwugEyYod4v4vr1/1rcFNhjMT04HYOtIkf+CBobREeK3iFNo/OrRaf8VkbphEd5o3xigUp8CaVca
DZKbrEKmj3SiwgjhEP03LdY7IwneuZaxHjVv5yHYEkpgj3biJKl7FBcOonarEmIKjJEM/z/R8QWK
EXCGKT7rV2cD0Vjat3+08BL3UUfz2Mz3SORFk0/OjjS0dpABpR5FsiUEoq7GsMdJ5q0i9SlwuNdg
BGfNw+zd9JOT15dzczW5bQm3wbtDOmO24B/mC1ZdBEObuyxIMQ9EwON7bZDZpCDVwQ17BTPZ5aOj
Zyn9dx+6pUKKlw6Vwk6ax3pHfOvaK6uI3faTVA8L+5KANpAdTjEN6p725BFBB8oncOvY9GVpPW9X
uI36p+Hmkdt/EwQuzkqDB0odYtFLKon+ojN4yitl3rTE0OnYZCfsff0GzuiNMmQNmaw+fhdHUHxH
EnTRyPtC7zE1dknF+uYOljQb/bbLpcHficVQeaf5GYNZT7bSkogMR/ofueig2cTplAMzTmKLu8QI
T4NtUy3jjwEGUvx4889dZBSEOaJf7l34UskYCylPkTGKjCD5hyg6LoLLsH8BfPhBUy0linqtKxKn
LZw8YyGIopTi+CbBV2S3yecMRx/00OnTwI5vNSMtnSs6SZhaoiKFKlXA2F8FqwXa4tPFNFPhKHZz
01lsJwHpgEk41vbakfMd0OmRGENbAUyRNl1K0YpnYAhY/0GkA2Csbe2vDhwu3cy/JPOHQOaWZEFK
uTCAdGbjxzO2dQe5bOgCKYqqkyL7km4/MnU5bJD1Xok1cGeMO9Y0n54VvdAdk+DvLE6cWkGmSMeX
OEZD68AOmavlsjIdO7kIR6RTUZFq4vliDnDBc1Tg7uDrNr0Da1Uv0/SK4NWKDlq9AknhjdXh5fvp
36ISMfbUqTphUOJ1mHhZsP1Km9NKNCnm5Qazf3iQygETFdLKnCHU+SzEH3cDityLv5ZcarsP0T2+
GKenV7g1dQAFBD8oTLiozbxCBrSCkKdyGYz2HI8WPYc9uz4G/P9VCkeggsdm06wOUkeZSEthcijU
vxOxImxVktqbOpbU3mHSoLdVqoQEI5eB2SH9XjpW0Ts5jEYxN0Cv2PpyCvjR+P6+ET0g/yQa1YEf
nt0nRL3AxDr+/LKY51QRJVZ33bB0ZWIBvPMX5Bu8hoTC8XgWFscpjo+BgxLA3KCGQ27wLqdRJFDb
4nSKmJEkEJFB3Lh0VkOSatQd63+3J1wK1yQ4lAzZhAZT1t4zC8PTUwmFE+TMxrPOZESk+TTokx0K
QCM9R0meiBBgx4NH8NVWscY6q6Pvd0mTMfwBChfOJY7jJ0YCAUEVSb6epsBK1pbCZAUFm06mCHwx
nyvkkAG4JiLn11KpQ42mUp4J1gBBXX9da/OZg8J5oL3QlT0ylYeaMnpEIGUfZu8j7SEkXMMEDzzX
76ZwKpz+y3c6xngJrzCmiKTSHKTkkIgVpxRX5O4AOE/RkKDU/+jRXuLP4iS/msFBNxGDfO+zslfE
wXBHRxgIXBAEtXYDtBFbRqUFHahF9WTFplvyT2AhY1yao3LgigNt8I77OcxqyUw75X0GVtD/asGB
oOXvKJRCQxGuGwUS9gReXN/J5cUqFeCDJBan/eZTPfWwmg1x/HnyuMEvRjbuGAKljNzAytfvMhwS
W0vJ+HvXwPAV3cPaY0HT+XcckvkhenWszFXAwKV3WPNdJuBiuTL6YeqXLyGJ087RMxulkaIKlK1P
cQX2vTWmo8NFZJ9jecUnbT8kIpZzE9km3VhoLItj8t483DXAF+XuikMxw/U7nYngrvR8gCvZE8gF
jrcGUR7AqGGmNSwuurFxl3nqMI/KoSE3aj2nBygYmzE46UHbl4uczbHy5vFbuB0UzXiPF6glXg==
`protect end_protected

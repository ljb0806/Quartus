-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HJPWQ0B2xGv3LUgHo1eGYQaQX7RPb/oneQfpyuiAd5IIgmyb2+VTV7ciRuYrXiMYFNf33LE0Dpyj
e0ttR9NuLdHYxLb128H2XxcLZ7qlyYsHnGxY7ovcm87DeLYWd6NysoLPIn8rYnWyyDdQlMGLb9zZ
jZS1Xgn7ZtTQVN7oJ0vdPJDvp0ZepF7YyBQ19KJB0F/pwpvnG32hJ8ait5ZVC3NNpea0wTfPHBqM
IGSUUNVhkVQB8Tpv4V+L7MvTwIe0TO7Y5ZkcYIdhOIYPPCiUsEWJeSosxAFYcGdafHfsoga345uL
I9XxQgg0sryhPCCYFb49ckUQUfInDPM9UVc7Iw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37584)
`protect data_block
/+djeQ3NsrYynMeoXBI0Igta616SpKmGIJ+09/NGZWfF5k27LJuabaPedDwXZF3WrV2AHWx7BeIU
ZqvvBL+i56hs1hqPAGiaQe53aX+Q7Pl1iDJhSvhpexH29MmzgLvuLl0xj50eQDsxW0RspZFciYjQ
iUpirO5WwmhauPB5jaDBFLDHLI1Ya2+uGyfmGtBmH/XVwvJs3sIgduk+vj/R8SShCEWWQOWutkSg
Honh76CWxzaMiHTY+/D8CvSPqX/eNhQ2JFBEIYM0/IQnRTpS628dgoEM4GYBlsYjoupgLeBMxsIL
Fr12zU4/hjrR9aNkO8gVEaFEh/DYdVhPvmrbs/fn+svcWV6jQ2YehUrH/R1xKRtpv+wjbr0KzdmA
aRj717wKFmsPhfRCfrbIO4hKL41QqDgfazD0CM4GYn7bMWqcvCZWmteNWSAXu8YCqedWiHUBb3pS
BwBwy3WA/HgkeD8sYTVL6mmaUrizvmxTIRwpZV3zmtbE6QOauCtIh9T+L3rBcvxtr8XY9TL6lEbe
8IiGatTHaGsp1GPj0jdzA0ZffpNMijPwsoBW6i0kYi4J1Vh1n7u0TJR1JkTEYI6eUiXK2nPBIsgI
cQmgI7zrx5J2LPCqwt7QeWJ++w2/mC0fQO631VHrD5Yz7Ykpz9aa+7xoT4XCiKLAxEBFq/Ci0Cta
oFi9fBZcI8gOoutVxjTMQ//OydMwxlMf5HpmeGVY2c9n3Tf3/OUjv7lZ+fh2d5P/QxSanqjP01kj
vvFxF3ATzhd/evcXo/EuIHJ6f7ST5kYZwOcsTcnoRZUudvycpAL4cxrIJjRUW4JnrdQe6Wqv5FWd
r/JahRMHziS6nraoYFya+NljVUIO0JWmlsqQrAVt0x2W46DcR7E2SfvlnOk0KBkz+Weo+/37xTfM
vg2NCpQPx6BUGE8nnhNSIZjU48CGVwphrjNAAU5oZIQotGUwhUeQIfZBh2H5OQZCdERcGAmdCOB0
MP+Jb4TTmNaPRKxAcopdO1m9a5L1rIlfsAFOmii1bW8UBsrkGk8X7GE8sr2TA1mfsmmN7JZK9X6o
VQdBcsoBXF9AB+kl5oEK7okWDi6BveU4SooBpElZ9FIij2qtYGTyjfChbvA8rNX1MwKAjpGWEJ5K
dZugSxNekeXB4JVewiXr4y9DOL6/E+U4rV+iB5y+cMItcT8cty8RCSYj88nKphEVcSdiyiGR8sp6
16hRgTyV9zxNNZk3ELna0Nak6PBcd+6puJ4twn/pGuyAokvf7k/AB8hllb71tp7gPicbeawPRnrY
O92rmoEWJjsBT/91Ag19o0/gzy6g5jUXKu/YfIgtUwhbsikDgQAWn4lcC6R7HCw6qCBYEiUa1Oli
a5n7+YuS/PscGN7WyLDuRE+k3KbTKZlhMCEU/RNXogW0KNcb46oEu9eHo1hRrIXF/TPBsluUfmtS
zWy7xmjDcS/S4k6zKh3msoU1X6hYEThF6KXAchvu+RqCLjEphvXLFIepreQvUL5y17BF557RJRIh
RqM5Q0/I0zbVHrMe67PRlX5jMhNSXiB538k2QjJdFrr8H1/AKI5F9BpDEoOkGtIOUOD0zIhFwsJj
lLUxR23kumSU2BHPI0HrRbMOL+Zw5gu5RqvyK0Vi7/2TKEVraiqUDKLkzO3aNhq0B/fuf0CgjBvw
jn4cxmUG9EYF4MXYRVi6LXhUbHvQONz6BIC8wQYVhLmG9TT7KdhVPXOGh+0fVHQ6RTUPjRXurrcI
igCpoyfXEFVBOglt2Jl2NUYddewS2iE7KkTEJzuwkZdIo/Bxrat2k23fOcY+7qPdXdpNufamoeKn
vLouIaPae4BtNT4Xoa2tI2DSAJQ5UA7KbyKQ/Mi9J5qQf9DRZBN/62wbEnZCM7mlMA3GOAh5q8p0
sTg9R7l6sqS8Ax2h8f8tBpC96ovdq4k6OG/VibZDmt+3pkgXeVL0Wpp+9/jsT0OukzwDtmm63Jb3
IY0HR1+gpGRkiu/xHHE7tIn0NQLNW467sjinRHHRXhG9Iiw1FIyNB0I9NOiUgSUFRg9HbRmAlq20
wyS0umLxmaTxte6vzj63Z5k5/5nSiupRwUR/hQI1IOKmxvdOK98HrFk6wubeC8mPLTYQHlTbbieu
pW7MNpyGYSk5in3wc2Q4Ff8J6W1P/NSh2s/7JQZDvYoykdI8EhPXMMX2c6UqNwlsvh2l48TmWqMN
qcLoSikoWl9AwjsbBqjrdtZinLXklW3lTKYVr0/jHYBuSYtiSUoUClWQPzcPBe9fN3cljibKFJPO
gmQc3DbDWkXcrizitLW4MwQUwY1/dNbZvgU4Q/wTUN0hTyhWg4DXUI8W0k8F1TqJAcsOnK2D+BWz
bhzllZN9Gr0JU4qbNQd8HHr5and8jb9acJ/N0nYoso7bcXit7X1m5qwFNlLIR6tzdTm6YyvIC2iz
HKW88bKZq/ylF+q4HcRHu4qGQ/gR0k8SeL3QdzljSRmBzfPY7su279BwfedI0lGRwcaofr06WcqQ
d6GWejGxqJDOIbTYIFZsGmOh1bdUVaeHci1/w3jzoPY5nDpUrkrN7gSwcgWJkLGWPVw8rakor1Z5
li6VeScaXEPznwFmrYdYBISft2GufcrmT2jiHIlIA8l+CMdee41+NY7IfXB0rafHApsASkpBQW2L
hEMLeJC/UnHKMYDStdxr8o4uJ1GAd+NDozU9f8lk+tMxLYwd+aXB7wH3E1ATcJ2+m6ZLh4m/q7Eq
4txu0gL/v6h7DZO6XHYTfPFMokQYQsK5f9JxXoQfk6kjsa9C588XdO0WPq9se+d5j+Rq5CMjUzg/
mNNwRP5rc/0ech5CJS1fGQhNMzWxmx3zt7h4oAP/B3BcpPSAyw4WtYZUpuMyLOwvVZBjZSdR9RAd
xrrAY4PNZD20ppV7IJqTV4IFTC0N/BhfiQ7RlJK50bNsa8EAPocTX/6b+rccBaPh2D20UN97sMKS
gHj0c4w7+DGBZRWOw9+kwi2Lo6UCIadrMU4vk631qXXBl2u1mH23aNq5punjsOk4lgjmVldwe1Iw
VImqRpki29nCT2ZXD/S/+81HODfmK0u8SdVSlOtA4S1X54jbSL94EpFbrMcYLR4m6DGVTXwB0rX9
5gx+S985EKA/iklaebBje7ufAC3opyRwhlxStBO5ZlfyF2l6LgqepDsR3b87/4JR5KcWGiJNgc1T
DDp/W3ANsIGQZA+S8eqSjUnWWCJBCA+dsB1z8J8rmcG/nvmxxvvd9WCdsr2s2/mmgxvdjxaO87oF
T93wvO4GRheAZpPVYYsj/EDD4J3Sg7qMpUXzUh6EzMnS1Jy6rXHdlKIb30cRveY7mcocp1cJSht+
CoyXChhudEvEkbBLeaditgAEv92e8KFKzKSbDwkKtk2YKI766QSEeNF8GSDktBNSqnakbBRf1xku
z8l/Kg3BajeXYdB+r2omhamJhOVGnGtdPDuHJzDzOu6GZvF81JTAmiWql3wXEr/AqNAk+DUFWe6g
0NSsK3fyJeTwesyxPNZW2qU4/pF6D8WvYdOQPx8oiYnyUGd/tPpuDESRzE+sm9fmFpsPUHYJw+Ya
pBJUOAronra77Ej24MGC9x7ylItZ9HsS2s2dbfaoM/KddaSXAS+wTZlx2HD2mqvdr3L7zTGziyo+
G6SJ1A1Ef7CwH8mY/oVrYmpFA6yGijX2KQw3xFFb1tuNnx0EWngw/7djBLiMxkUqUn4CDWrizK+L
1rPiVYI9a2skX7QJFXfF4oQnD7kR6h2ycfvAHAXncvpLbyAHcnQ+mgrMUpdzFjNJThoqVtiqR+0M
ZCYlGorbUQ693/moFSTVGdYqSmv25mc/o2dWcSDQlJXJd7l3S3CMRu5cd/fTsCjE2ia8X4Aceis7
FZyAmTOjPwWle0olnREovzEH+8zzAGmePkQVb/7bEDxe3WgD+OBX7utF/bcNk6zIUKDzrA/OFbpY
cSwgoR4ALax0zflP9zXzAuwxgrLdxrMqcxWJ94P9pCH7VvMrOawMGdMC95CtUgWPI5Zga688KKO8
XC75w/ujrRpaPbfrqz2kpZlTReeuBRhMe5MJ4z6sJGufV4ffsMjGPdfWC2WLu+dIHLvEgdCTr0sh
nLiKTPOvaD0JUJOB2DKn5ikAjcUOKu4StPGINt6Ga2hb6d9s1cs5BeNpAXtd5B2Z9tTygStxk7x/
Cr4r9bocLa81COa/K6L6b7AnYnORPIUn+JkOUPlBlJWSiuDApsmtRJ758/aCQzLM8V6j/vZ9G3Bh
GbMj5h/IXKJaNHddM0+J7hz61Jy1IW9wtK/WX6bLlI+4X60kY+2jYefZvFeC9igZmEC4CQlYUjIn
HVQDqVOAaDR3MtKZczKWlk4ovEMDVM37CmpHiXEnrN5WKrYAZfVf0vWxCt/eC/MGDM14+Syt5GhU
HM/84r3vx/CwwXWDrcXfPKwSgdMTwYdvB/Qm6Mf387yNIYLFRg4iqk4bnqNfHZOtyF5cNw+RVwlv
zlI7gsBI87I7bmVBkwbGfCOhVoPK1cbNwL0BUy80Im5luqiMfJN71lyoDhyenQGUs9JcE+ACqauo
obIrrrTTl98nTkmRFjW7jJW+hV1I0Ag8St65cuSX4C7GsvsvtDnTgC9KYuQSOjmSmLHiUqrp60Qk
zGp8yxzKUiQVHKA62NnaKPu3vCE+SROSpFpdIOfke5A+Iemf99Eb9Npq6KfTopoNkk+wQsUMw3i0
sFW6WSvogZ2gVdDbI4zZIpysuolemfvF+F5qHUzfo3AfOwC1m2cgYIFFaDdq1qXQb8JZj22jlJQH
5yWb5smDMsoNu/4QttXOng1FGUK5epNEWoSX+Qk5HiZBh+QcH2iJDxhUof0NysVYrsU4A767xUU/
wq8VOwD5BEy123PBoVjdIR3sGK1lPTSz9CcCX31idmD4PZRfETTU6Ec8LOvIijw/jwF44DQqVxbR
y1rCLezRCa1NJEF6s8cD7zHuDB5E2WDx9bTBkxPb7MmOHI/3F5DFfGo3bk7fidaAnruRl6rNvjsg
vnlVdH7m9dTzhgPCHitAxFIP57UXiZKF66Q3hc4cIHktaxU1Gs6D2vsOVNBnSgiTDycGFywEU/PW
7k92ibtmZ4MH4lrxgDjssnCqK88ylxCci1uu/1STOYX7fz/AQS1QnxmrBkLNvDTuhFJSaQC29g1a
60EJvFtZ0pawKJzv0FCpZsVnU8eBfipLrWBOUTdXc3nu8BgHVtxLCDtnzUbGnj512k7qCaFTcGdk
WW1K/Q9doYiz6nGEC/z4W7DggeVOnNs0MTOL48G1sk0PceFbI9y21cshObB/qAxqJk6ZP4996oTq
DRoVwbewe0FS4ch01GLUQSWUagYEePEE6y7eaFDRl2pJtrxaWLfkEaI0w4Cr/7iRO79FnfmkUUPy
sHmqRBGx+4eM8UJgIwK3h0moGoNELenRzU0ACnQrzBdfGmqK04TtJzUwC3cl24Qi0VmGI547pZdr
qMMWPeZHdNeg6RWKmrhc4Dax4CmvOEtuu+VKwwZcYKWKYtLrSuK/8Xz5bzZG9KKw1YAU9+e+LWQq
OTyxbNWot3UB/lW+NNLx4V5SWnPyiO2bW174xXy1ArbABjQ7rjukJj3DPkXwam/6EhEqrrIoR+S3
Q+J45KXn5YuJjYpOkzHKW/jUOekbZwuwQn4iqx7vbUIZC6bcYQy0vQO3HLq+8u1u1NonkBhLiA42
I8O2LsF4AKd1P8iP3+CGVmwO9uUFCXL11RvWEQ1pzQON3LpKCMq1+fbmrRitTjNx0aQmk4qVVR5J
UMj2m2qN53l5FiSHnmvPPrukKh7vxcMkGBLnIyLV1DdTD3OoSfXP7cljZbOwilmS9CreigjLy2Qr
Bp6Nf7TGhfYC0yd11budkxsg5oN48K48DjkKC+I6/xcLZuKe5bMRVGl28pFAK1nezSqSrgVqg9gT
NXkY5jv8i9mBkN5X517WcLkVEAwkuJIYZkeLNpoDvH7P0oa8korckJEt+Ls2ZdWrRWRAs2ZKp5Yd
d9DEl2HddbUoJMDHZjAQjDDpA5QGVYBMfqwt8NahFXAQZ5TcyQUCGfdZkCmuKB221JexGSwnt67t
5+X6TYaQKX0KMMkOsvbrH4H49kXB3N6SQmHFQclYcnBHCFhRzvBQRcFmcZoJS4yVhAEEwxh2Znx6
3ddSIJqp62FpttHT997lBty0B6WFZM82Orjfv7MH1na0s1rnBfgZGpldcH4ka9KrnyyCunE6GK5e
PiMK7JcpH7Pe++DWxx6kgSWGjmgo3dT/Gp6yWAyezbx5WphU2SCGwwN6aIJT+yi2j/npGO6ossoD
ZEkNt1BzOa+Kd7kc8693+PoUVH6bDEqemo+h9Q/TJSG22v6BjTQQGUiwbUjzHhY+S3jmTW5HhyG9
HRWQAb5TqLbrkEIeTYyPIxgSGpQHnU88OaJQex0YDWFFqGQWSEhGkiWF7XowiYtwkgSNrZWUlAJO
u2Pe+9oEX5pR2/0JxQ203SpZr644EjE7IoFc55D444FwFNOpM4q09G5Sq0wwgTR5Zb0tOX1R9bBd
WAL2tuRozXxbQbeOd531seZNkD0eASYnU4JKbc8I1rIGrcDV5FE0ys0G2hIk/VsJqT7lvzbeUZMT
gLnD5Rftb3gz3HlukTHzHdr7qPaP2/f9NdcFM8qq5H/Kg1CNGqKUCYdSggm/H3ZnZHspiHIcSQJR
LxSeQZ/7Y/QzsKhilgZLIqtDV/NvE4bLJM27uVT6nW+VohfYudHLF4cn1UX+S2bkGCRjUJqjJAQ3
tAZN3ADPA6yeEmCUPsqC72Jziwx3rO+vJ25NmInQSKpScKWU1mc8Ki+y2e90JGXtJckSX1/2zbiw
+WgiSrULn64ST+lZxW391WOMm8QATCAEwM5ZD8vqWd54bDgzIyw4IowMTIrboKtzzaFxTumsVl5o
cOJPddHK+YQy4LlfFbIJiOI/E64eyZyyODOwbMqA1MgJdey5um+0ubEOncdklzZUjIjDgXSMcOce
FARmrhfznHzSpTQEywzeO/LLZlAoqVGO1NonN7MoupT/BEzaxvK3AOre163jxp29Wz832VFBlYto
7CUKjvXnWqPsKUTSmvEZr2EQHNupGbVrd3Hs7KoaDpw8YjrcGsvtP3JSQPNgm5az9/d56jQvo2yR
B0sZ3+XjYf9hA/qshwbcIY2eB4hnp/HMj+Bq9RIpQeKuYkLj8gGoI8IA6Zqv/yYHefrqmGFz54wl
udhGioWvT0uVuSmxYvPiwhMGoreF/WYAoELRwO0u7GHlI8bmQpxWspy69BsDd/7V16zNarstZkFW
mihERg+aTZNvtDendrR1sPz8sbY0gwPVOpTgBprAoggvObDXwAUeyfCna8UE4Z8kh5yuNsjmgGTi
+nbxyxab4lJ/btPoG79Q8Cz7CL7j5KL2r/ChiiCL9WfEOUQFYYfi0FEodz3+ufF8vR+jHWuG32VV
NpoOk48zT5Tk27F77TEYhBkaBgUCN01h/eksEWXMzL8HS/5rVHIW2mFTMxAjqixxKSlWT6TcgfCt
rVOHZTaazPVPcpEsuqL9yHqpdRDMT5jEYCvPo8CvQRBA1EidTkI09HGBbWI+U/P1QcsiIyIrzlfU
5VQtluOJ1StpkIqv0YcFOg13Ru5rNXTKflyPvuvJCfhKvNKfl8sX4Jx0DuJxcTl9dmyO7sqJFVJp
991VBL8bJle1dLetAHnCoHBbIvxG/NYWbwHaJ2Ja65IfiIlQT0Fecyqk0rdk/v84exAjO9ivEa80
GxyAbCv1Laq4BB3bo9TH71zF5Uzb+LwvIA2Xh49pJ3opetNg/fVgt2UHG5Y191iKi9d+39z3sk6G
rdhq/pxXBtAb/d3a5ebG/ifHUH01WyNdp8Q8xqtZJlnHfDRO701z/8IRft9HQwlaIMzcGOCFwjYp
sEgjofs6C6IHinzSkaNDDoZLqyAfhT0ufhuwD9nqUi3Y8A13jJduxY481EsnOK6526tq5ahY1gxq
G3Tfd4/QpdWV1e/CtUEtXMMi96v8+sc7aH9iqRo43GFrhP7pELqxUPZQYXLdkVXsikNI8lt44cQV
aPeXrWHNTyao8cb/5XzA5gHRqV/c6asmhpcQ5fx0FKHefwF0JPQzv2Brnwf04QVsHMSiwW9urQeq
tJxCCvR+gUptk+XL4cq1UARh04MEUi2lNHi9yWeeiYkJjWK/kM6DtJ1WNud+eSwRqCJ2gbgZHl3q
4cN0YSYOl1QqgqzKWvaNNnwytcOgRmW5qt+sSLZzr92+DGsOqnxtIWCOmWvMBaZlpApXqwuXAV/D
L4sKuA3zPz8j8XyIdy57NElwkGhNs9YR3FkooNGw4j235k+84dJz08RebPcRk0TZASHSz4M/tZNM
9Qp/iO4dwoiR2P7YwN0bi1OxchtmZMMUIB990UjpQe6E+hsb0q8AV21oBk2qlpDAQzskALRXXYk4
Ofol0KGSJoRenYUW2T/FGo4Y6hr7utb9GKsw0ODAo3ChkcAd7ldsqT0WAW8pIET11K0lxuZONbyd
0snZyr1VNaFxOxOhN5RDA4q70och4XGZORzTih4ONiAZvZg7hsY+LwxGKr8UJOMLaYwblOn80Tx9
oYwld76sZUeHVNLlp57k+9/73WYB5wxLKvmmaN/6DRBsoPyKPKrF24N1PGSy5KDc8gGBwGVvOp/A
PKuuwUlf02WOtJRseRG08s9SG46ogdbj6nxt2C8G6EO69Bv11tpTvQ60mndcaoy749nqlMJ/RDWn
GUm1jWZ0xGAUwbN4rY8xKrNH1Hu/Pnbeap/LfH+5zax0/KOnk12Mv/hPNVlLu5YG0KIvCVU+wqd0
o8GtDxbQIZQHD7CdlMdGVk2GWyWRYROyiEz2x4FqPOHozBdjOXLw8/MQhB3QWPl/SJqHar8Lb0L8
luX/XoEuQXn6erEq566fgXf19jsZvU+MsiFd5/+NmUJleZ83ZzhSqXGmqLlUSD/FR7sVGVLNqBzL
GFNJlAgTfpUlg91hswRfDUi5y92cy01qHXUqWCK8HeJ2GQfbsEkVOBTLJ30j0J/DE9q7FXdrvYUC
T9osfWve8Po5wbQkweRFpJIkYpo2TYm9RRvv0ir5C/7CBwwwGCuiGTt3dvtiSUutKNld8RJHtJ81
5poG14uqOTWODCGuBj7/v5ldMRXTbCc7xGmD+sT+Xb3m90CDeL/CExBctRnHFfvfypchLUOmjDue
I1tPAEQBdYxwSM1LA+UMyKri7IdbRpgNCOXrVIfbey/f2/k6Y8j6LsaxFfBwddFGe2HqAMBCHfVl
DNHbzIPa7miESacoynzNUOY9lRhu6gzFIlTZVe0yNeZ4q/6IKg36uj9UbY779cObhIHj3XyRUZ32
+f87eLNK/eg9rCLo3uHzXt4KOZbLQI2nyaSayUOkc5014QmNyL05I63HR9K9CVI5NpF95p+8PjTG
VjiAuw6H5VfnK52jr35zUPiHilWexyj2WAFk9FtjeKeNeeJtLXh75Q8uib3LZJHoab+YPNAJjqDc
KhF7Cm1PCEccJJa27mpwFDNYQlgbicSdzr30kC8VDsn1jLn0cgg5YEYaYiQBroltybfhan6odTEf
rpf9oAzAYhVbm0UYfDcFm3saoihmF0aeebAAYlaEnarYMnJiV+dMQJm5VGyiBWEjvmDp3TnWTyQU
IwdTgqFUklRL8tbSqrTs/T2RFICmZrEF2J3cDL3NNd2vOA06ZPRLDGb0uzI8HZT3Ehg/TQUzpjdI
ySH9p5U4h+0T9QYYbmHHoGaCLC5C5JX8GNCEIBA42Lrb3FANc+w5cz3ruqy72xyUjO5dqD5cOtAQ
qvygmFkjBmPJ56cFUQiJnmOa4/0nFB3lX41/YZ+0t9bcJHiBgwOQ4MsjNowW1nWZAcm+lJKV66fH
7lPHkAxj9uS50yaZvmPZ1dM+UnIHj7CADzH+WCPtPZ955lwbFb25uMoafX05sDX1zVkkkDgm00dP
5vu0nutA93nFITdPNYp42sjrMslI7/rK0EXFr9GCRA9G7EnvnJjNDM9OGnMsfX2L/LhsGsRhry35
U2SV7IgEF6a5eAGW7aaCZe84og3bV2etnrJOodyw93qLdSEeKo8g48VtM+0+ucTw7MduCuqvMTzU
uHIUIpuH/z/2G6RG9v8Fol+rRLsXR21ia/0FxZ+ysJ3G4mVm2HHwkyhCmSkSh6XawTMt7yrEw+4L
RagwhcWRhVZzLN2gARUnHR4qm/Nl+ZOuGprY5ycF/M1LHzOe2mhcVYKZAMp5gufp/s3nDh8n1dKG
uEJOvFkjU/txgz69qhkE42+F+sWf+oLIDJNiZtIPIQv6s+sqt4uiX2lTHOJOxITVQ/2VmoGLeChE
V/TbB0qaEJtzY49doz0S4JwpsIluWwSxkOwA94ZeaF4Cm/f9sG7tiBEEmPiHQZRvY2qhskxg5IyE
9Axrs2K9Bnxk2gf2POar46PPG4xyOcHWnxI7w31f5HHmU34DjkgrLdePCWnoec3Hqk9mZcksfTBl
4q2fYoyp22HEMzSZw1dInTW3hlitDLxYr/bwbvoyweRQT5HZPGQRokHKpkpRfwINsY8CuwQUt0bL
CJ1ClNMatSL+i0cUPccgp39NSLBs9rLuI2jtRtHBnEduoVzadt+bL1tYGva1GrOnkqO7sqE0bl2a
VbfSQTgOMnQzdxzEKP0CNGn4y3z73H24RRjkaZU8LbfRntt3O4yTf+tYSDoaUh+zrd9l0y7xP530
rrAKp0i/UyUpbyNZyzP+S+5XZQuV08Y6nvdzpcI7WsPOiQ84TJeV9aSKd9XybUGHkHfEcbAnDMNH
tIh1xj9X9Y7pa456dn67RFIyzzdYtGFIyiC7Ahpe5qUdjKsC/uE4RGwYF+7LmBg3+dbfn1U1EKs3
vUxb2dyBOOcyTxcL/332k8msD1cOWmZESdpqWCtS+TjTJdr8p7TZqS47zRKMvHS54alNj4x8fotR
CC1MjzxdecQLXGdK/yRg44cLZbkWCIz4UU14vmScblsOqNZVyhuA5lj/5JHtUI+b0ZLzO0m9uzLf
aQiIT2VgxaGWvC9Z5sH8gZusp7QAu4rs2/3Zs9Ref/VNMYZC5AWaiv3okbhrxPaNQvkiIP0qYXdU
aoKVmHdmsENBXIIuGfeF1zbxbs1pHhALOMeIeGVEedyiLbYCG/iR36A3BD8imoxjWPsmafrtWldD
mTFPKQMnITFxUHFopueEWDrmFGsgYj8DRPNG7L9gTmnncViQ4st5qBKjhctuH2BqXxU4oz23Y9/s
KUv4OvFSF5B2tViEs1TbYwaP3MvC3L1+6TfuHVbND28lYVih+krpPAYl/iryjqAYkCEKB6mP1kYy
JV5LyHPUWXhtpxDOg5lkLeGDSIi8WBudxvdKS+L0aZVCCKG4zObZfvWhIbrv4mqDUgmuMees7a5d
/2rHnyrkNmL78jJ3tWiri2OflyOd5RiKTzeW9muZsowvQQqKzg5dJuwb4R+zEQq8NejTtMJriX3l
Z6fsN3ue+Ez5bVDjaxtArWmUk1mit03SZklfPUY5dYr71KpAVelrUrbStJjewlfJhed0KCVptKl0
goiV7dzXz/SnwPNb7/nPi3Gg2e2wueEnf2lBy/qdBzC/hfZmFGn9/9oPgBbITcHSil5YnOQolCfA
IrnzNdSJI0FjT7kXcQb0GQdgmCToklrNrMqEla/tJgK3lLoRSANtyR/E0eMJNt72OjmQ44xB3IB4
ScYoeUAU9znQ5kAnpGZXkiWqFj/DP5W+IWTjrO4f462IlZgZxfreFBbpmmo+SP4doa/qpllOUm6R
GH/lAqMsimgetJOw2PmlzYiS2D0ukfzefW1WTAtKBcnKg17N+ntO4BDGXLMdeQpMorwDg4Ir0HH2
9N84cDVw9dd72PjJ8dwsorrIyBv2illkj+/ZkRJm8nll+pnkPkUV43KGt84ScP8Gej1lBgKSXOzk
sHLWpKAuWWHXNKvFsMnBxkmO8VmzMwT06fLKR0AtukayCMk12+Nb9nd7T+BbmsYMeybbCLpXV3L4
fx3qBYAJs0gr/hh9YSAXu3PgbPbUKiMtWAN+dwLXuOlWZBhdEsXnRrAE7ZKftfEo8b+sKn9q5d6o
IVkvF+v4clnS1z8K1WVkQB3ylt0oTvN96r7y1ACU+XDr9xIje8BuYGY8z26+V4BooKcceCeYY6Fp
WwmQ7p2dAGS3DkNZkogCFVY10NmIB+i3eZkM9zE2c9j5UlySpmPVcfT/RiNL+JqTjs/tabLsNweo
uEgobXQDqHg+rmMF4kcbcUoYZ4dfnALdqHbijr82oKuigdpQTMOiwNygiXzJjW1mkCJ04XlP7wSs
Gfwi3G1x4PU3BWqMshquCfhulRJTCOiP+v2Et3tx4rSaqHhqVTu4EgNk5UC7gpSOALhac/OYFIqC
VZ6KvjYQh8OaJRKB+q6dg5quYGL2aqW4KIlStJBIFdLR3AQ9dCA24wH/hEIh6DbzmdNPeHGpRhYX
nem9Z/9sfIg14dVh1z59yFpGn5TqGIDkWGueGQ5rDJsztXrKQjdzsXqPEYRMf7ZVmuqHbWknAxXQ
GS4i72dZ4mgrlVpN9yTWbHhpmROurprDrba6JMbqVBY7gkpsI4HHHx8iYGC1VctjhMAdz0Cm2irN
v7ymwgLiqCETb6wNvEQ/NOL/8WmaMrh9xwIlMjXq+ZEhUc39OudU37aRpb2SJhiS2+9ydEF3PLvg
EDWSipoD/OAbKKDTlg6UTx61jPdLl5wEpaSaWO2tRKcfShZCLH19JDX+dR+goz0DmfQLVHVaI3nj
AVpQTglcW7JdbdjgLR7QrCNLVYLDzReEWM2axlI8a/oBX+5HMl1ZoJRVmvAHdVAliRy3/k+5pbU7
OtMQj3sYzRmikr7qFaCDMDgBQbX1C4tsIWR9OGhHuPbNEQNkfTR+Vw3ZdtZtmg2bSH0TF14RRvuz
Bjc6Sx9U0mo/DymKDGTXVROp2MKVpLWaMUhuME9/v4Iz6DMvbIofDFuG0wLrYr46xJpdUFZzqIK/
6MQ0XwzL/EIONyKEucOrOjvoZWtH9mw9ZAUA2zEoJpgmYOsUPQdefel9QFth3UewtRUWF/F3VWAr
vbR+Bx7RSfjlDYwG+2Y2LE3JNmIn3aY3CpGtafRwv+V3PfM0iLrWW7Tk6EJrjq4PvJVx0lACxOmd
DPvE1jWY5IoN/lXzZ7FVz/1FAV8cEOIUqdb41SXhSJXP7UNZYWXeRxpiGlzV5su4+RkF9MCajn9X
6nxmHbJHNJ1ETuaNrphqu0yADYKauzVfJMfB4eIy0YZ7nnIewLV6LyfxJei/4SXl0rlUkyu+h+kY
NFYGrNoM4RXaiFls1al5TLjEeP8YONRWA3wxOGSaJphHCnOO05Y64ixdbTGM1tugQJaXQtTn9ivg
uJ2W6NZvyU/Dg2FSduVJnEF2OEbPNF2ZV0CiS/dtZbgB89Z/0AH16JIbpYsVhKQpO9hvvJnUc2ap
aVmb7zYeFk0KcOLqpDsLb2rQUiE+xC6YcwBnnnmdWHuWVqqC38ZyKQW5dDPVM0HGX/WuflMo+A2r
NYLk3NXVJb6EQJMQSawO3NpT1I27Tigjq67PPMgkGTYfT2HBfUjCKWeVUn4hDS/j6COF6wKvQuG5
3+LtwwnCVo0clKk3VjHt+EPXnKHaA2t73E+XPgtMxALLzpBfmu5imsuwctHIl4vpMB9sYUsDaVkX
HdRGeO2dq4h2vDyICAa0oGuKY/TbC/qXTwJSZHqnqs5EkCCwg7nJRApnj4PjRZnuLy2fPwmI/eqg
SAsPczwGImsWortUYPYJLKY1pjEJf/HHbPu0WD8XD6dmP1Pre37eBFQR3EgXXD968nV+fU9iTCvu
jMIIL5L7bMTt0KQDqja7zDO47MDRgUo9DB3ZLAdNwY0fjJHbznavz2NGBcFQxW15ceTDuSRwRF6b
YTqlIixHJpPUb8mzMRvtRzZqTSlQzhSalZ6sL+UEvnROuWdafya6bnweKR+JjfI8rz01CztSGFdz
Ls27ruSvJ7SE7+FCHDkQCELwtFWAXPpwhTRveeiyrPkkKGLEmc5vSH9Bnkx8LAgw5f7fIDIHNWM9
tB1P8naAiOpHnIGMfZ+p9Py5XiXCKS7Anle48RP3r9YO3/yhkgfJE6zB1N9w+gZrWmbyZ8XW8ozk
vOWmWyzPHemvSp0g3FCFS8R71S7NtqYeJ+xelrKLcQDchx7TxTG+/ceisbAMmdnEgAIGD2WNmkC2
pcRXmBHQcjXduff3M2vNZhQXULCBiF2Su9Zt6AOjyw+wi83rW7hyTVf63q0cej2dfQbi5fii8xXp
JNJz3Qezuy6UExd7Q+DfPDmvbSxuoYpRNRy6qo7f2310jcbSdmw382Xwh67eAPto32SCnT1ZNFtq
VNCxnOs79rON2rqt4G43ZHSKmQ2Yd8U/hv4UKpnzvYV3WM21d6Vrk8PAJP6ZZIC5rq5NznNluGua
8SwagkihaacHiTX/4rd6Iq2zeAv+j5hkMPdJCBYgZAg0lg5TOvjo0pRx54GSl3YeGpoHRap9dkAL
xEaCGVo2rV1NrtOwOv5u3cWnhp1jH4KO1kOP6fYYLNsHhWLymHvqKjpeD6dkFeswQTs9ei4ebCaR
53L3OssxA9a4pXM5p8vjH95Nk0PN8h5G0RhJ9LCws6tEeGoBG0SFud55L8M0WjXgL9hunGCn7TE/
auIkg26KoBjlmV2Cj5cY2yNYiVQs1NFQ+rYPifSopLF0l+A9er5NQ1Wrfbpe675tMPu/X6hfP2A5
Of+hMzUQ8JbgtHhk2sOmJj5pHLwanQ5Fvs0FwF4VnH1beCL9sz/tcMbm3V6DlqTVj69XNG/gbnbv
alktm3WNbxoMwCraBdM9262e695qBHst1yKEeRn+OuMeKlY4tOUu2SKdryv3pmWPXEQVrBmtAq0M
uyFr7AhPgpMrRYTWw/klscvnm3gCxOVslpN2fwEzhgr5loFPq/ZzAno5Vk+p0tPvWAcMevonfJsw
MUa4jL2U2/joXRFMaQa78a/DsiTMu67Rd8kohUYehgkusTt370t35bndCIYhCEhbW6HlhWuXjCjG
vM9NY2yLvMqGztczCTgZhx74iD+MK/VJMCDihED/LLzpMswzDao/Dv2n8aGQNeO4fZiuuzi7DTRG
LeBml1Jiajy7vRW/WYjnlADAiaeXEmy9IlUCGy2504S7LM0Z5vfK/n6ETiepwP65jTwAvDGATwF5
0qjC1UsKCteZoMpy8toxgCLUW4GrJnl77pQQGDStYXmyMpMM+o+BClg+9NS7/UMjHi0/BsubRVRv
c/M2NZbXCHowfjVFpukVyk5VWVKliONM7N4VofDGqmoOTu9rMai05FxM+VcEa7qTI2WII6n3DRxc
Z4gqMT4URSALLc8WlP3ZnpN9izhbO02whm+gVpvGnL48hpce06bsBze7vFt1BeJCC4QGcaTxCP/A
TU8SQmT4kN1+QjV2INueLGj7GkE0+Dy26oiFba1KgKBSYpKjFebosMqxGMoIX17EtPv99UjXgVXK
UMWcYkzJt3E7xgfk8s/0nmYiAKb8SbI3uiJeG/574l7ZrfclszaAu+5LKD8sX5RmVWecUOgYr3Ws
FeIMj4FfLWrFz0VAIBH1BNJBFn3OLkWpD1rxy0hN9lZl0eUpCRKCxZ+uEvKfKOqRPtNlNJNhzoeH
TkE04gL/gU1h/3LlbluJwCpnFKFNQDyMQXE1ul66uhcqjA/niz/6GYDPbuQZlb+E/QCtXpV05vTQ
o7WYg9wvMLsrzCkZs/Qv9V8URkQsPs9SMoomVMJhKTpFgxVfyC+bTZO7pf345ZNbRaQyQ9O+fby2
pe+7dly8HirzRtUtsFmAns+rGpkL2ViVs7hn5n2KiSRengbwaN2uYoyDrkoqC1b6xdduz2vLTdeB
H/M8+1T2IoQSGdH+XcVnYIL11hpmlLks6TjTjUEVlLc/lw8VlhV0tFGu9trA8eX5uOjISzbl2fWk
SetPL1lUMk3BRVjvO7Jw0IlLGEg4Je2R6DQbtFta6Azn2XwIwnULPh1KxoR6M46nr8bgKwN/W5xp
XUfr2bf52xFnqltilEgb+TaYYTkXXJcWRaseB9Ga5Lw+re7ZSd8ADsaSnmJS/6EjYHzOEDyedZM+
jMeJNA4Hn/feCHOIHWZIdjYeENd0f6qDmLxL1XpEsWHMg1crxxZ2NT64QIF810VoiSn3k2P0PJk3
rmeg7XWRR+WT1LENsdidK3/q7rE1uwrQ5mNbMxbvRHD4RKM5+BwMMVfRMa3wQB+2ayOjvbD8taJz
0SqqwDLDmuygfBJqqay42q4pAYrHvsNGdw6P8XE49e6TikFgos9FSH4Avr0Y+s3hKey1k1iemHyo
kW5iHYs7bNeN7eJJQe68OFL9o9TLTjdgo2N4ESmUaKlhUwdmRPfo7/JlEYOWFaWla4oKx3/0JGnL
8+WrszQFYmdB4nxdY1aVwyJ425Fe9WmhzXQxJaxE4U/RZEl3ggFfPFoKCz9p01o8U9FaWt9cl4PA
lsRcTC2Xal1v2/xnJRgxxVeUxtST6aDBbrOI6GY/7avIdImniB6KP0R8Cncgj7W4s0d2iumrw6Kd
VBrbYF/8UNwTrd3S+T7f/znfPV9O0vEVCPyyXU9W372lfs9O+FEB9u96nKoMo5Na8bu6bzNyno5w
Jw/oZaRyt4y8fG1cG88WgF7WZHtVfRxJUWdPASGs3AED+F6LOyNQYmu2UbNvH7Q3FZGSb+zxcSd+
q/igwn19CFdi66lA00HYqxir3sKFW+s8Bw9VlHJzaXfVKUZeAHj/6ht1LUAzWK7rJ2VQMSmw7XFo
AKJ9WRgKDFF/AxcU/sp/EojDpd5l9Xf+1cg3oRZavJgM/t+smTtfi63ST6lnaxQEwbsWTSCAcrlP
93+A5Gr0sVFWMwge3bIMMpff8kqPDr/hZL8GtETBKRMM/EOG+izKqgVVIPlIaYQPQnsJ83pnxh9U
VM7ybz9z8Vj4gPI9iEy8Dl7M07cdREjW+dZS+KVdBPlzGW4HeGIxKwihz9wfQPnoyyubTsStL7Aq
+02tU7KaYPF7H+aijRdyu0FQWL2QElUhpv8X9m+eOV8ONcpeZG/3p1C+ET//KswYGoQBO61albTz
PMtF/oZFIlMC8lYIT5h65bFI8Wu+Y7amzwk3BSgWU02+t5Qow8MPAjJwGMXuq90LclEmD+SeQpg3
oaHTPtIVYF6/2RtVKX71bxaniHBz5CVnDUNovkvbgDdPHzoJPhqr8h5/61p5uzgA5vHx92S2TCab
7HFMcsXHfNFjvmUPcL3uh1r5/I/qoWQ4+Z+fn8fTTIWAUQ56ZCHwkVDVTHPucyQOcJRcpoyT0sll
IC8wrJ4xwxT22jWP4GZA2GBTOIsgyRCF+5crLWN3dQVXTL58HfiITrr8mt3WSAmXRS89T1rh9O5d
oyBRDO16b41NERG2FSiwWd/w78UMdd5ZavrXtKCnbuZRlyPQVla8CTgGFnzO3LioRp1K0uScztp/
tbicApxdEOrBU1ZN0pwjE2AfbBwPiCTwqOpI2FiGF8xYKcniTRe+ADyGu2J6n6KWrxlCtSbfRqOo
AX0J4zEtH6juHavC9ZlL2UGiECIemnKaN6wjDKV6E2OsoDK3LCvZr5MyX/qzxkEtGtSXlaJ07QT0
3fMgGnDwK/ZijhLRiS8TwYamJ5nQ16Y2d0pXlhSmwUYXYtOfRiUV1qIu9z/coj5kWqWUpuiAKV3n
z2l17kfKLjuyCE+l7eHTqNHvZ638tePupTzBRQpLTWNgmdch9OsUcMtfMxruzjh73A7dyDlBBeK/
Ph1NMfACo1EJz4uvKVN/GbopR6e+/NCPz5Q8z9IhC7leOLYYLHT2qXh58aZ9exyUnzRAZVlA5/93
Q2FY+nCCXmqx+mU33tGTxtY92LMKSFe67v6RyTEiKD2l6ikNSWmO4MN+1ta9yJ/EtlsU65IlIhRo
cNf4W5OCVBZbejFYd7TcGCk2E6Tn7KR+uYGg6/P6J4bcSD8sTShGhuW3XziQWpWYrq06a0aT1H8x
DE/5xiRmU7bH21AyYacjM7e14kXQ0RlTYeZLpN4DeBooezg4pzWB5qhLsb8QdWhnEn/ipV1ayr/l
5mTcfbbo6KtjNmRumjzpfOudvsicHSGSZ8UiPtwxZ1Mu64eCh2YYvUDpreVG89oIPTr/XHULIuJi
cImN6Q878jhquaT2Eg9jDZ/3lfefTwkWo+DPbxbFPjYRsmUbkY04MqEPkKMmDpoJOaug0yvHuIT6
Y1g6xGGnz3GKCoEfSMaor7NpU9+wLfLy9XK/pPEbvuZVfEx47nX5JQJZ1OPf3Da1nyRhmnL0IBcZ
y80rKqILQ35i/GfDfQJz7ti6XTXS6Gqf/H7QZSzbI4FxNnFTaRNNpnHsWMtF3LuyhkBPCaT37IUA
EPqmhbXX6F8BPJhqzYluiHpWnfRnguzad/hO8KXD9hjrIU+vepsCfGAb3aem2j01dhvx/t35kTjc
JYBkQDFFvbOo5f4AJVvp2smSGq/oB43diVUQUjM1fwwotd1EUAaeTTKjwjPEe9EANVubxfQjLGws
amYYdLicPDqpyAyllJ+SdNnLldTAPgTy8B08AxWN/EVBhNNZWQYR2qiPgcowJxSb+X4ISyQm4G0N
gjXo4gIqjHswf7EsqdFSxnZtXLOaz88t0RJmaNBOKrvi74pyAQXfAz6kyFfUh5WUTv6x82fpppmW
yZeZGLmwoLMBDJarKiM8B+O8urOnDMB2WAdn5s3kj4KKfEh7ZSAyYlynfVp7u7NgXhV+fsYQvTfD
dls2ay7CEIxHbIC/37FOncvWV22E6pRTh6qx9OuPiQYu1yDoeB+qrqjujvpiTjjpuwHA2umI4mXs
wnMQx5zfFUqxohh28sx3BBeTW15T+mmUD2YiMjF4rZG7bskwsh0DoT4vXqwNU+moomZcdOGX7SyB
tuOOrLUwRbwKvJB3+oV6YMWkefvCgiENB/ei6sUXWbcqOVMXNVvovceNFjVePMsyl/uB2iTilSkE
E0G9G0+sGPiEy2XxJCVQcf4ZpTxE9UDx5Vym8VJe61XQo6iSVGO4KKMFrZwyUwnJsHZ+KC3DShfM
7W4YI8EK4dyduS7tpyhStSquLbBKiGvmo25mgViM4+Xvh6WwzrnM6wtjOnvwehMNEUXrUU6clcUi
HqO6yXc4xzZJvegctXFi9euehl/WrYvlG/jHn82Xcmt8EC85dTunaUx52PMKYyPU6lek8oE7+wSv
Zq4CUyMTEwLE967NjKpzibMVInw9hmrq7FtokAQQsB0/W5QQR8w5zOQcvCxb/x+/33lf+1SyQtRk
r3UbxFFMk6O20BboC5rVFRAmtXNg6FPJJSZIv+Xj9UpmZMhWonAS6eiHwTfDF+hcLdlwJjhSfw6T
BKrv2Xx6HucZYvIis17lub/8qlJMpUWjmIsZIQDgkLDPuoCVxKfJcOtxEHVR7I4P5bcs3Y04S2WD
WAd0LXqMjpJFdTJ4uN0TkChUDgX00ulpKf5dAkLJ5uJYiiZ31ZpzHV2xC6PH8Otl3X82wOuxBVBK
Nhf9aSYqvMAv+XvfbihqJJwMxvXjm1ysl3dB9CfBGJUrYRhlNXCj8qozLQeEofRy/t4Bnw0J8ZD0
k7z6i8TIINQeaesL9MPxyNA2JoCUoYMG3ANavjkHg++UOrUBwPTSlvwIlxtOgw/RylJRej4haA5+
YEIYwC+WQgQQPHye9aVEUKcznj2e6njeTbT2f5zcurHjwL1aW9q8fvuNjVC8LRjDcWrYpt1P+Jhu
ptWQVyLbCIjZVxKI5xenXfBzE8OjCYPw6AGMSc4oDlkVm7j/Coo1YZKWjm1LIP7nVXLbgM6jsuSm
ceb8Rx1BFTOFiQvPnuWzGAsR8ONebSIBA3zBW/nGNXuEXuEoZOLl3HGxtyzV3lFIufJcXjFk27Yb
2h4Tnd4dSHV8lMERDQEnMUTmtwiS5kNuc0O9+vLS1c6iY2DIj+owJ6LYLe1QqtBPtPG1a38zVfEp
lVoNasiFHm5J1zlDz0W8I6krHUH9gAGX7z0TTGeA3Yx4RZmyTYhC9f7IsNawTutu97gN/Z3CExf3
3oMDfKniNvrdGdEGiOjdS92rH8FIepQ56Cjoo6+5yFT9gwEU0PwyyMnoAINIFMHFTAc0E4ckm7VR
3bbZAz2QXnUzvedZTEZfCJFFfqDqq5D+HQGp6YN/2XEGmyprIE/nwP6OESTfg+kut3s9QFSA7+sU
1JuiVs4hJa3X7uBpDGe8HPbNF4CR/y+nFTwzYbNjESUxVdtKoMFpJXEpaHKmMrSUjg+TNgy/vmPt
JQZGh1RumoYb+rJzroG0xW7rnjGUuczTn48uM7zLUAg8B9qfKvUJ3sQNFXzLUsGWXJLvHU0O0KY/
OHZRNn1AueiE7lhqo4UHdBpZoLMLWf7OJC6PysDpPUJjshP4G83h1iE2psJQdB5k/YBLiWLa7Rwy
PxwvrB/kcyOg0iJD1Cl9KRZYM56vbuxzOPgvJUCH3WAcrRY88X+EL98wOO42yRbOVY0QGIih9Q3Y
ejafLnvnUTmQ9G8kY4COJlemtk4sKKOr2GL1HR78MbMz4SMIQHgzpdS37NKIjH8TOl2LvCZvF/+g
7P34M46pAOngftDEyOrX1g3v5loQmVAWc3OG6Bw/9Dfv3soyBEf4lwTSMcrZjLSUkLN++D52+eMZ
Hv+VC2Twe1tXSKoLzZ0svBDk1pjlxCi/Ea3xjKxCwgJ5vyyoeLhBPCRHTVAtbhuMLGHLMyIVt3T3
QAbPidyItWVT6u+h2GoHBjLpMy/W79mSgMIUnQj5XJawNG2UzwkhrH7xMPE6s/jQMQhvCIhdXU65
69ngY19x9S2goyPQouAZo5OmvY8EsnBiBuFEd/iVflBl1Jh5PJz76Mbev9ObR/CwwtuVZ5i0SgxL
+9ZHuvUekynxQCH+fyZzEu89ZiGPj6BFZuOyknttUI2IRVn+wpQwI3DkHlvvCSlLOBGzIN6Ia3Rt
Yy8icUPeaFLwzRzscw4qewjdbrz2JnCKsoAWdWAcx68UZcSJSuEHb5CNNKLG4/U5wIwWTxU2Q4WZ
XfsXjV4ZydiyNgMWTZnkMYM4dkyMj+5RWQonhGCNRDJAf/cB204tPexbyGgr7XDgN9GSiUs6thX7
JYfqZKGswldRX0iPjbNmvOjRA0sx923IFRAKKuO8V37usErtR1jiDBHwgcLyBnr+98D3ql0F/AZZ
fcwnDGTfrX8S62XT6WoRz/4deZHqzjoNHBGu+FLDi0iR/7tAi8wwnuIUNkO0g7sE140wQNplGVDZ
cnLJXAgbLPTnvc+ggR+RZuvi/0lIzmUWrL4D2vEX+BlX0qM/m88oXlLoHQSKT+yT25Sz0XEQHC7n
MWS6O/boUxRyjqEb+mSc0xU8hZaXWO3HFiKk6fsKVXTPdrdXI+eWz7azmEta596CO2RYNaNrOyZM
B+9OvEr4EKbTCx14zBwAn58GQti03VrhYGygAOnIKegv5DpQiINdZmHaU8RMskFkus6UYCU67HMu
hfO23RML0B1tyTR+cMclgrpvM+e7vL+2ZRZ1iAANYV+Mi1Ce0khBEW/aRMvfgem5j5puIjWjMftL
ddchv+vOpA57dKdVhuCMZgz3Wh2Qxqa/VDTmHSBTtYOusdRMXYlN90UoWeWquIbGiAwKRKfAjDLu
E+fRwYzGD1abW/G7KIkT+MZW9W46EuYHOLA9R+A9x51ascSPybRyj3YPC/zkGqCU+TtGAzzyxvMY
4vlebSadCCn9+CBQ5EruNv8BFTNVXiANzoYDd9JppZtSp0aplYzRo7LCVjddiYztq6Xgc5P2foHe
CbWp1R+2Jsq5s2oBtWkVWP0or4zFR7Ns2MtTzQ4Z+sqHjkrLCHsjrs4NWtJkzJKMoqQFggETYBia
G62PZ3sc9To/413YUzcNXpCGENoP1W3Qb1PDYIEc338Uxvlp4V52mAGEwOzxokRi6UGIBToCSoWM
pctgjb+H2R48se/FsC8T+5cI7SNEiJ6HaZIGNgQjEtHYszvWeUZWt3tL3xRGGrR1W4XdGr+i/Axv
Y8+cwQqeBnoc2MFrVHpH/PLg114XaZKcEJJFiATfsnc6K4p8LFrkNywLFjpa7iYl1oJma/L2kVA/
DjdX7FavEs36AuBY+3/HbDEATT6UuBb7I6MnhGiR+2XM9MIwvXrwwqPFLESewacuxJLXAn2xsysD
F1kBqsKztbW05wJg8wH54Z1qlVtkFUmXGzu0pjH8tGfMaiWiQwhe9Hfz5G2HBuxJ/IM8rTvVYjWm
/3Il22gSWDKbd71JDRs5egPqBU815NLu8lJoXGWmd2Yto/w5YOd5Kiz5TEKhYD49dWDlpDJa1IXm
p00GamtnYb9QaEaW9HDA94jNEK2vZ8NjVvwTNjhSYieUPvvnBeGxf4hDVDfC/2/sUzPDU60/I8qV
LPpIcgV+R9OpGvHyAhG6rsCp90SovGXD4XH1VNpl4hcRaKDs2QDtOH7BUZ+N2ad86xgAEoEYa3p6
4lSNeleRt5/cJapXu+Br34uKleie8q3EaIbNg7yPeTsrm45949e25Ej+uD9PP1wI/duZ9ogiC61y
Tv9/tIFyRaO0X9g+mO8kEAz7jmsTUp8fnFLExxArljRo5zOmPfGkq+87t/gOQ29rDeKVg49BK5xQ
eC0WEkHwKaN1Aa/x3STyOzJ+FsA5snziu8q+unpOxF8QlW2skIJH/vg75C+8VI1NngghvBDiFrZD
xk1uf9V+hEiMU1elRmcBKgP1vVgy+51kPsHT5KNERWLFcegeUOkqev5R14yagtENKRt/jJEi0x1G
nS9MjldOS43NReVfCCWEXjt5Mem8zC3PPUXmuGk09fh1Hsb1fzegHBmiOi9+UKOUICHW87hYcrio
eojBd/eFxcS2fZCwcml7xmidIoC4SuYNRm56Sdd2DMBsZLMphreKWIMB2M/VqLhk/IKw++X6VAmp
6kp+bjSMPhi5z8JwfrJto+8VPmzk3ygWvfZH22shTHebxYjfFC6e/4KhfhzC1RQC+mhcH0O7fOTX
A/MqunHL5xl3V2NxXM0kZLvjiDYMtIrQAjxhs2IUVO6wMcsW9kgmIfqkCHpTk4JMNyH+CuedoFq/
hHtzOSD+P/fc69iUfr1OKD938cqso7xKFJABY3HkUs6aMjlPqHD2HDWpTRRpUo/EJ79+y97jea2/
pNLRluUtYkm2AGvLslLLo1J15vn7aUVptv+nt041OMg4B+yOCobqT53XvSIrgNwujHWQmfCN9zm3
SPIdPWTejnWLY+HZfjm7ct9ANjMC6bERScw1jSFpm9uQbXJDYrVdYvrR6Kt1fqS34V6X6CmOYfxn
qBlwQxQsXyWvN+7exbq32nzYHDh6e7iHcIWtJUo+JrvSeOhs7+sMJfv0IzImepDzcpSau00TaS2C
+GVmf+9iCU7anXp4057PAqQpiSNNEY329kU4eGTUHhl7w0q0UXVPECV8x2j3OH5azPJARqLUWhtE
zMkvhUFu64OVkWY+UQHjORe6b4DXVfcKDVBdxGL2i9HTi2uWQJvnacrBvRBNtVjm8uqbCDtQXtmo
BnHr/EmPn26KlFZWxzcBj74Y+A6Qle38OLz+2Mh8ijnjWuR+V7p0vtmp79v315heiPkbPPAcRejY
XIKDEf9w/8Zk4QSh+h0hRlCVkOerzT8+GObGNBoDPnXPpe4BhI/rUjYQpGJTO94m97dvAzz2OV8c
CGEed1c3Kbldv3pTlk9Yn08bh0xPytMhPudkZI3jTIUcUNfxJYB2gn4cswzcJehKQfmQCtF+BW9f
dLincDriVfe0bpqfJhMBFCkKYQEj0ihf3mBhqNmaOAbi+iHkd50Kq8cpcuSyr3nQ6ERjUS4kpXBR
3LA+vwDRttqzIHmg6+TFJX2MCLDlIuPrRLKM38NsvrObsKRIOQFMPNTH304UmjOJMob9hbO1UgpM
F+/dtFqGEqnUSm17GLJer9jAbNsgy7uUQYYK7KutV00lbg/GrZ3h4R9h18enxhNCBe/Isud5IK31
tyaf4KX7f3YAtwIkJbRLMDiVUBbHmWd0GJzN0saQ9AJzRIaFMH+1M6M3ev9KmO06iVoPirxqvXxj
uCe1HxZ9Fu2SE0ylmoms0G/uY5BGT9Wrw7ynDjoZSKl5Q+zl9aHBzRVG6IOJFgc2aWWyshq3EM1/
1tR67p/nd7Xfn8s+ec1F7JKrqSkNicFccExsKd438y2F1ObQEMs+aOn5Z5Rnj0sXT5U/8nQLaZQ3
+eNjLwLEf0AMuE20KznjwI/2IlsNvfZh2jVLB57T3QYq0zpi+qOlXaR5q9Lg9tx64dU0SlK6+Lid
5771EjJShk3tF3DsouREN2BCUP386GFDvBQvHM+5dyos1T3WeE9GL02Tdo/JguVxfRNe7/XUMX54
hTfTcMpxCiWu37klG7c8s6lxt/aM8p+K3TN2F45Ammrf5OsFHkA4LhePrCRUuTiYKrEP9qRuf955
0AeAUvMkgjfWFnQAv7YAGIM/bxGKzuK6wLMimAgZY1ZqTaJP6gl4v9kuShO9GkV6MfqU70E25lkH
2J9ZvyrgOujy1StXTeiI1d4Q89w/0vfLadcEA0FtRtBPenSL9LBYMT3B8i+i8BKXeFXM/tQkDmBc
A46UB5Ozmv+mePjIp6PXOxKEvqq+A23S3+168jUFWmuD3v8BxFSXT9yQwynfO5EPwQTBeO1r/PXR
svYJBOamDjxQrBd3iMlFYG3YAr4rVrTDMq2AT162HbwRFJbS8R7kdX343K8oxIPxOrP9wiMXpP2D
WXYSxmFcpm6yOEheFkMQrtlzHC/as4CB+mxyan1wGd9HMJ19AS7Ob9WCf6rI+Sj1gjtcNckipOWa
cyS+An6MJd4rppLcZui8EhqyjNIglWRbYBKPYm9ii81IryLA/AE78HfZgVl/G+rupBikwTCbB+Cp
kzVFso90aFLxGyTtHw5JRbg9zPMivUrwI8sfHIuC6ROFsUF32fr/Ve+YBPx3mXxR0f04W8G9IuSW
2h5/K6yDCdIXsYirlVDBeaRlqYee4PUz6zDDGxCuCl9OE+JshYLMCU7NX1sjV0dba+7VQxFomCAI
p19rFPjmSRwYVnPWvo7SH5eQP9K/dJIpCR+p+UL1r1e+IMTlp14pbyhF5WR8fz2pbeGmWyHDgICd
Li9CrcrACFgq2yMrHwoc2MKLLdngTxxoDuDaRtikBxKO2AYazNDJSMv+87Sf+xD1hqBONPf9fQyV
qOQup59pvS1hmCWsdw9N4P6tAl9zMgYvlz8dqJQmpexoE99kyg04JYQ86zqicwuzXaGiVhsH26Wu
WsJLNgZlxH/fj8r6Emz2rI5/nDMCMevKhAFBix6XrJqDWZBC7tf/Et3V8+vTCtvEBeascZdpWJ3D
OOjNVRW9rzmQTpecLSQzWVHaJ97m0nVEZMB6uJMwOFjoAuopqgd//9/j4vMvMlQZOPm1NR+X4qQQ
HJxMFeeHLjuFBPQMZj3rQPFfuVubeIKZgeU3OcL11H5rzKVSXHstvZyNwYfrZnR0L3e25U60feTE
a/Da0L2UHtCYPp3RjoXgx68ewr2l3korsN8tHq+X0w23SL+4oarjnPXP/qYVLTbhalwel92dSr5X
/lQLkjZXEGDfe0gPZq77Ne4BQ4PAaGGueLHT30vbwSQmUgpkWmgpaN+UQDzHwSXClahhzMmBF4mG
ve1kBd4yEKbRMmj9VQpCeD0yX7xHTaNOhX8j/8glcYNi6Wr4MvDQmPzxxISQJ4d1F+O8AmIziMAd
R5KPhvP6yMadkLRF0uutCzDseGeRMXa1hCPJ/P2DY4FdqKdH3noQeUSfxlP5AL7JogeUXYXgm2Ko
vIgDAmHW6QirnmA/sShqJPKgJXqAsYgWpvfuxSETSKEl2El5Tb+PTLZjwcpld2J4VPb0ozhZ4ON2
tXK66qAK9w4AFvrIE6Kc4koflVpDMWILatsDR9/Cw8IqyTHYNHpMSm6MOn4+J2e9rMBzHtdwtNJd
vetrUMuAEtJcrrQLSvkofJq0ls7MUkw4xrPnTafHd06l9tFAA2+AJFqUUbpKUaUaWhu9dWRABpRa
XGD6Est/3qZaGckJxp2R61QGO1YOeIEd17OZdhkOMX6tWtkdVl80O5TnQfTtm8E9k7eLdY5rxksl
vpuyP684Bw25jcE5CNYMTrlylvQmawAXzh7FCsFdRVrYCOd6CXF8uHbgwwjQZzBpu3ZqZzdupuU1
ywwClRfSbgo733hXeBCnBVesPZfuF6SepeYYFUv8u8Ve6nlnlUGy2x5KJuLNT3omTAqhBYLafYrF
AyVrSveN1yeHonbm4q1k0A4neHnDtEUAS3VlK2YWxNW+z1q8nNYi9+s1c9yKQlGr+ts/JxCcOx5x
GdlAYjGUusaeGrtq31sn7RM64kBzfCRTgrMcsD06iouUc4XFHMpSIY3MrGmbD8Mu9mus66pVawZl
4Bgp2jKu5DEg1VZIceLzFMjePVeJFp2RwuNWllNwYJkzKn9NWRQXKG3mrQcNQpkMjLE54ijlq9oC
cI7d9gZlZlB9ahTa5wChb+jSNF3cA6Emzg00/Snou1rbUxhUwOI56qsx6u6o6kBX49uysvhIVITv
lwf1ANNQGfVaE7VvAB0lBaPPLsRILoTJCkiXS1Gi2Ekbr6sM1ABdxqu0YcSlVbOPd54sELVhFn8M
uKYqU2Qear3muXMX94J7azbLITSU2BWQ8V97tL73ytoAi+1AD2QOvmRExY2UGlmOZ2X2bS8xGCho
5k/f6cBUvjC1AOhpzqQ8Wfca+HcXQwftAksQibETvKFZcl232cokjQiJtF4AGWJpgKD2MU4+JlwE
YyMrlB4gUfECiH0W4KZCZs+nMEuJ0jMs4aCnFSIctBz+/3/zJI0oaIxMJuV553ibaK5kSR771iVL
JeU2Kh+FQYes3QH7sB/wCreiYhxuX1INyL9VhPpiwH9BrCgamKoAIWTZQLxp+GvXItd8c8sedysa
621M8hhfn6U8CVnuolnVwgRJjuBJU2VwFZ4qqAPki9qWR2MZ/hhJuOWXkyBrGRBnAsdRCh9ic0Xu
qooaxyliVOYheytvq7fuKp0yA/q+SdRIsDcix9otPZU/Rj+MjFkmCVNCSQz/u/o57byUQP1ZBp3U
7jcHwqsKKoirqkol5zTqIwQbMMsImibvvuBkfU/FnnU2N9ZSyQDkirdcQvG46k3gsw4WG6Vy6guw
OF/ClhHfRVh6HMfAO32ITXmAE1NnOZkwRHno70NHWMGA90V/MGGpq3p4iQskgH7za6amvggr3xq+
ii+p8kHyYhWWHupZchbBnV+PN+0Ptq42Xg8ITvzU3xkqpu9eTv7K5CqVUf/CJNvB5K5+nDjj6eVI
ckXOmqWgDvf+yLRMLuUi0VNWtbyoZ8p9KvWBihCq8H4T8TWggtJN9XacehsPKsBE35xhJdp5VPbx
UYAP/rcjXAdANACRE1u5a2+9McqqKDaOo/9JeN8A8gq39mDLXN77V8NRFccvmXJVMoragJefYfjD
B2ps7PsbXwBfIE0OD9gxEMPwYNoC/82U32HiN1vo0xxNea6BylvOZbKYQihZen3e+RI0IuPGWqhH
aQi78rf36W8bXKHUWx6218rDQhNFHg/LW/tXcOQwll4bTGKViGusbSmkxCPO61X+6wnyS723lesu
Pa8qlrTzMbALW64CaoNt2txIF5xic8Cfq/DuavvnPFlIdEZZs3JirBQ+KKQ8oCtCaPR3vqJTL62h
3m9nfi2mzV54uuvBsqWrGj2204xTmTEgFyOBumZ308mEia5BmdUZv6rXIDxJxSkA9zofdgiyP3/0
cILVVBbzmT7uk3/khdUr2sO8wd2Ac3u0PNVM60FtCU9EO3QCfMN4mIlWHX0qaviBtXuUvz2Za4kV
QT1+DWvIYRMLk4MOu5ApMki2edIjf6UsXInuFNv6ZNWlZSuf1midCtjd9qwFWiOocFohkM7l/k9Q
kRVXET8mBi48uaCL7AnW+jvN8wTh2X+b+jEQGWFVTyY1Pd7YPpzFEn8F5kVF9AtIUd4TWTcLh2EO
DVrQvDaAyT0XxwrHh9dHCWet01yk+DWjIqPmWorbvgwGAanp2iSUhWeC+CJ+aBXrMrzTnGILV8tJ
4HGOqUe/UlQB/R+Vt1eRpz2JEOkmAj40r65x7dDfwKaCjW/GmeE0xesPhg7y1tMH2FOO8NPAuA6U
/pE9nvF7ES9LI5xDzINsguvTO5IsgZLNzBLdXHwV1qzdQHLzQBEKMu253RNESOiDqQxDl+dz3yrI
KfRkgcSJKeTdnspvTZF5JoEeLWGPOkvKKEY3eU/cQ/slgIIuUqE5k+bVb+mUbeTpgfDSQuqws4Lc
NThnAog81qLpRGqb6EFWXP6utawzX9+34enqhmDX/xJnRtzlIG0sWTQtk0xwjBKMk7lMqCU6+ohV
bWFvUtCGve9le6i3VmsYI1xkvBOt+J/aTen8fAm5qIO/ue6r5AB8md1ziRSFutOa99jgzS0ZKk0f
flBlQMJSEHLaX/99i520r/CEtiJZrcSk+bbGlZBeyP7xUZuxX4VE9wcvcY6IGjuokcWXpeqUea6N
xZ0kIhmrqfVvM8FEc4wGpS97IloNmoCVlagG5N2ldpLihyCotFS9JZB+ude9+Kid2RDVkdTv4S/e
CWI/rkUcGfB/cgJRJZR9O87nPNO1JbcBR9urc9ffd/EUUw+JiFPOjFxjESvLshdnCQS6W/bJGGNS
QOSzIuu5VyIVtouAiut+dGh5sE9DOnY4tyPydIFgLqU5WHwMYS2RlAGBGcFIfTI75OIy3DpuaEp0
Acpy8GrZq3yGv4QSOWXpzc09UHb+ptt3Z7rooTUK+0kiWpkyeMLEzWAnFuTsZAfOekaVSSHCjTqu
DPQdEmJQt2diveDNCBWOjSJuLFOPCG/fXLfHDh1zX7W9UgdMw3espDNttfxelsq77RmOPmxMPt3t
jO3KcbRHc92W2S5cUzM7ObRryeikkS5tYM3AOTpnz/57qRAOcJPSoMpKg0D5j1+cLm+1nFyFB+l6
W6qa3kWOqLXofuL0eL0lU/anqwXc/XpaUQdyPACUSvmSYKML+ZlBeHtAHx6WPzMBdvEQSXEmWHE5
ofPDTORQ23zNm1wj20Jw3QCcvQHGXsONw3tOxA5zV/8xEvAzZveF8I/HnRzZgZ0QEYccfEGxPvTg
ygQdyR0+fDQ/PSkzxDCIW4+qxalEKgSOM5wbL3U4dr7MxOTfWPmPwThc6xYc0pxYc2whNShop/VC
2q3oCoPPb9y1dWd2vUriv32LU4QIOQYSBrdA+Ck7ni0xXARiaZY7mhzVB+TJ5TXFLtni3YePf0VU
PSus2DxCMY2sMDZ2AhIIW4ahpMUfjaTX4iua/ceBtNNImGQpQlcLXg0ojS1Baf+b86/ssI7S5+Eo
/CZeJgwDg6K77AGWPNA755SkfDDCW6dOQ1vyIdM/GONLhMdFHCworq/J1PpsHkqMRsJkhz16MV9N
rDrPsLCZI7VGL4yDgjz4qasZjoGGWQsmGckgUcviuXN58MmSrlGZ39z2OB5fQtNAZU24Vwe7hPKp
dTMMRELeFj2VZjdVTNeiJY3efQuINRdAnM5fEtrNcpYOPlwoYtZ4+MCnsM7BAxxZq4sA63bzHvSM
LYC0OIwxKPJpR9y4HytkjoWXNYjA68bkIbA/vxfvg42gjqHoO9FNmQ+zd1wHr1bTAbTgGF/bp7+/
ConFEoF75NApBVO/GRrloFCTr296P5gqXLkvntxYf/tXv5rfNX3PwdCN+tWZuOsqH1+zNWZFPn5L
CTQV4cssTmXOS+8RD7cFkOgChH9DlnYhr7mMg7tpMzLP46KCYW3J/YJ6q4MsnMAJTsZ3rGMuRDLz
bLJuqypWDVRxNapv7GOuA7Lt4F7FvL1PkG7vsy+rbLpXDotrG1zjjUBjR46mxWEt+Tr5NdSeb5s/
+nnxmn7El2Q4s0ceWSJIMk34UlkJaU+tZ9n5j6vx00S4LkEnTnHCGWD1LBJnRQ4JD4F6HJMu6KIo
d1BwsrVLRQMq+IZcAZlxzpEum9SiPznbEYkYUebx8bDTKDI58tOhXaIEm91MA2Af4RxPMMXApqFN
N80abCfg7QrK8WtBGqA8kpJfBMpKMzRN2DMdaoAOVaNBCOB2vTpUKkfYJGkyoOmgguwnCPvlcgJw
w5/JTijtvlhTO3bP7vfcd1cKk4wk2LwZKI0a446h4muI8AbL51k/AqmjVdISXx2EjA3BJaVu8Kgo
C3/u3NZP77TAqiScovTyGZuM7PRqjTsvRdkgVEDqC6HW0Q/ISPjIztbZUKNSZ25VrG64aN49EesJ
0WiNcmvASADH8DCt0OfSuRa3jxX/6+1pccUaplbafST6MyUAaZQkuJXq/J4vfo+e4p98ZT5lVWEA
vMn7rcXCImoeogEyLrOTJgjAr9Veu7UtDJg0U8Hf1TRiu+ZTHSMNeHUltxjJSI/AEQWWotQUCaWU
Brilt0B9lq5CiJpvhcJXthuWK9thLzSeXkGxR+XfmcpSxQuflpT6uXNeiPMaedcICfngHiC++hPN
+qEr231tEWKUyVM+7AYCRgt0Xez2v/0fl4YJopW5jPzPYgkt4fIiRj0L4aus78jmq40DTvBLmiJY
h7Ry+s5Jc/vWWVSeSYgwr0WBOZbcYAylRgDnYURbvkqP4JHqlrqNFbaHM7wsHMzjSuKLVNk1WWh+
pG0AWeFtHtsfhqYIl0aHcczkwKMmzurwpmBf/JyyVIviCLUw5aqZfccTntY3mlsQ+phXnKUZ6M8y
O8VMU5SynmFCSB6DitDzpXXIb4fcU1ukCs1K9dmEXUnwMrHrV+sc5KrEEitQgjb9K/2A0JpcGRhJ
c+Cmal6OxQ0Ph2Qtd9PwbHehu6JBwKH3s6DRQII077M7DlIJr3BN4BiVv6a+ReOK4jViw99NstoL
3UTGSWFiIkK7cX55ovqoiiGeesx9epF0nnva4yYB4GPQ+k/yL2Bb+HcB72Gc+CufvlfyqsHn18mj
Q1YGTXEX4iEnthM+nIGZ1p7rcWz0sn9+KgomevE+IOevmJhNHoyLFR/6iF/NPcP4drbKP7T0Qb7e
5aymX67+/lEgh+tW5YrjhynT/U8BiT9PSihMsfdO4P0kk1pjiZEj53cO9Lj/k6w63SUcyf2KMOui
2BiwOZhp5WAxuRT088WXL9kZ86lIjZbtY930awUphiuaioEWXM99jqY6PI5XfviWDwLN+Hi12TVt
VmGUZtjTXRnWDxnSiVD5+kHEffW4EirqJ3T3CcP4iJ3qQ0GzfojyWtdmOWi1APsE1Mi3Z+DRRct3
esKiEgNLnHSlplndpYtiMuU+uQBcLqQ7sgFzWahoxvxH06+4Zvx/j4Ou1P7oTips1Hojd061lE/H
9BVS6AFTq3d71X1m7n4S6U0ayfdjjrMxvFfGYOAWLSjukiuaUgPL83hVK2AAA5NCwPASRMZ3tO3w
cyXTgKvzdgOHFgjtTcv9jE2s+7FZzOWDIXhJrofbCg3EOi8ykR4eGlunpl+EHjCA5FnMWN/fmJGw
WqCXpI306YXPTVrdSpUaIZM89k8OppNMG84hSSNyZw6brtGEaCteKp8H/DGFwhezF4XZRmAaLWUB
0U7v42G46WZGuvpO4RHustSykEn8silazrzGmpz6XyTM7d4NH4MLVSMIJMBtXGnUpLMTqeJnCuLz
0ndy9o+G/S9dhh7ilbPvO65a+Se7TKhc/bfQBiZgoXUM8R6j+5siYwGARxwAIIp9COx17Se79tOd
YOHQHZ+z036+1Mmr3IrfNii/f+fSFFLJq8nncYVQbgOCx8hIGUWsoxUwsCh8Dba8zV8AR46MS+PV
xUrS3uhyIYUZ6dmD93jYZt6KIaIqY7tdvEj/3psvIubLJh3w5QejY1ZvPW3d+Z3wG1dpKSVVIadX
0tzEV5ldTOOaOQqxuWb+D9vsek69jdgB2wW1DyVnje5eyO4+Ej9unLYtZbQkuznyTI6l9jP48Y7R
DbOlW42qyMXU57x5XU0mEpvpl8FF+31r0q0eHU39of/ADS9Su2Umqiofv/eF5dtQjdAjDGs1VBh6
DR8bAZbks/ybuwYC34Jizg6eKFvNjM2vNbiKw8ebJYmTgxe1D7C6522nGhPKiPMRoGhGxUFWv/q7
pIMXS2Co4MZ5C0w9FIZWjKaRcRabgClZ2n5Di4nKTkCbjujy6DRZViuWACagBjNy1qudYolO6VE1
He0EdwdeAc7sqJAyXhK8UPebw9nF26UoqXHy7erDrOp0PFXC8KWno+ACfWmssZbNAwBR2f1TinCF
6U7IqczbejynfUWqk2tFc0CDhhQ5CYNcB6nfv+3zqU29vMixVKKoP/iouZ3D2k/CC8pyrBlO16i8
TTZEB9z7bh7rNUMcOZb47Imprnf8EpUSxaZMPTelUvQDWPYQq/V7BcoSWyXvXSoVMlI1QqPCnAF5
Fu/XxmSLVWbmSGi+tsEG/vRtKs5d+KwEBydA72SjEaBc+CO5jBbc74BIqNB7AfBD/LYNQk4MbjaX
IRF7U9GOBiuTWeT0ZP/1v4nVhkTKVl8PhjpljwTyUbYCTWDemPiRUpS/1+W8UQAqB+RVyvFC/bNg
If0qNuTUO1GA+c/ay+0A4Df4LaV/ZJZTMyN8fosZXwqYP/fnJJ7+Mq2IXkCsPWljg8KnEnfhia3u
+qYRgY2hhdeUmzoX0PfYx7cnDtuKtGAAZnAz0t7YAON5sr6xNLxmepMb2e0ZCaqKKMsN+2wYKmQr
OrUjPP01a410b8B+co8w/3Ofm4Tod/VXOOT2O+flrisjOBAfjFTCQY77pc3Ei0A0PV67KCzQBk4f
F3QaVsxwuYh8jdu/QEKF2F5N2uiPFUo7RbQrCfnr5GhWrUU6MUaDYUmsCwskp9jn5kNm1IUS2YlV
zpMVdSTTkJJ4weOs834l/N3A9AyOD+l/hYv1EWeHGszwSJN0UdV+FxumeGmjP523yVvaPMJ4AJ0I
uugBuiPRjxljJe6hOxFSOENHsbWc9MiJSGtj5rUlkfvdn3NerHho5AXDsEJNRO+adGnOomkj1Hcx
uqtSPgQ1OY34ZSIvaGnJ3Kc1tLpUljd6oCZdCtxfhw3+JXgLNNfG3JlkCC0my2qncwyvQXShOLu7
geqc79jvfcVmkb2twhzdA2Z4aSjjXPWHzkm5Ds1H1Gc4lPfH4PAnGnXfSXhtkeG8CdUVFY306F2L
lgbqTQ1V7/lJqZKL0/i0EPGhXtfY48JCXNmapStwCkZIINxGk7bRfz/WuOxsgv1XQC9mVMZU5hBV
1qjzwXcqqDz1z9nPj3oSu32FCy9Rtb1LmDURWk7xoUPnDBLeFmmiBXGDiELXMR4AquEY/y8/gn7H
J6bXZ4m6Wu2T4wO8gvVhqaPmczHMF0uYNaQiVtUVhcet7qHYW+JkrVn8/5JFeDUU5tIiFkGy0Vgf
pskXJq7WXtMB7QpFO4J/vBMrpyd438yrWoFEiAkLaUkKquv4fYQN4iCCIc7IP7Uv04VxlNPijwro
8eNEuOTuh/KEbgJeH/wO5Xc9TSX+i1rJI8dLSJV/k3zzGTkp4RIcVyLx3STkFZpdScruuUqsK364
V90U3hg8m4rhmk1a2rh6VqwI3NLEzzeyArsvBQM3oLpFzw9Q2wVq2pMSJterE04aA2D3oppESHRc
B4F1TmWkmoHSYrDWyvTjCbqV3aOqoXfCFTJZSxGJYwMOMvb7xUlbA6PPoALc/d7ay4lLL8lWbCFk
vglX4Q8Q3hGAXE4c16ZiFavT0AlJSykHyiP5HafAoRvIhfE9q+3AqfB31jlw0Kjk55QKUtvVJhgd
ERixVYZRIN7b2T4BVmZA+7s5brI8BYi03nHBD9HMyZk8hJgfWCeldMfAZ6aEubS6qbHo/xvE/cAt
Oc0iKs45XggFbcCk+lSpIMJXU9aYvkLEM5AawwmJGabtwWv8Qq9NdUo6XQzIqEkDD/Y7eFxNHhw+
8jMJua1DXLIwmhvirhyaI1BjQvOlHYQWUZtb05pJz5DYrsaSQnwXdcC3PINNw7rMklqbiS1Kwfhc
wcxkaBXxNXpoQtOhthlCWPtjG8kjq7rs+w+dmZQSQoQMcSTowKGzLvp1ysRfkUly4ZZLSghr6lDg
oTvZTkNdonwGvPNmHbG+QL9YgwcN7aa9jxENr+crYHwLRh9M3K9GQKAZ/gZGfIdJHD8Kreq+ry3h
p3Z2FVhOPXQih6Nrr935vHA/Jmev/rnmRHCaifx5w9Mg4ol/RUC3KY3UKzzuvw1xXK6ioyhLRBp+
ccw0y96fOey+cl/AZxuBhxOgCZotXWGOt2Z/24Dp18582XX8xFH6r/FmzAWB97Shp4u9+anZjB20
NGWqqCSK6Sho4t9foWrn5QIJXcwG6OjK7gvHagFXZKX3mXQvGaNYTE+67+fB9rq5bwaoT9Pd9J88
wHZgUD/yBW9kAkQsXGfHlC5voY5ZjrbFidMW9WfxfTj6N8gMd86fn0GDds6Yie73LbHH2dQdHoEb
KIB0KURWsmsXOQYag+XTRgcZJtSxNNemZjDN0JuWYSvfyutDqRTSLTUevcBLEY0oHWAwiarlFGvB
O9Oc8h5tdCQ1WyPUaiOoEe50v8+LPV3RiMvPa++QtJRGLpjVIPA0pyXSqcDTmY7hicWWcGSPyic8
M3niTcB+RJd9+PjQSi0NopFEJIgO1e9aP6lxXzaINzBJRbIo6/2Ds4zgXiv6O22DkO2myJsDujBV
lrauO4y+j9MhNuoxhJl3NmM0T70sLsWCpZ1UKUHoJVMAJIzbxmXzp10RjiqzDoNYGA6x0Z4HeYWd
RBRyqKVSr3m0tv9iXakfxtiM9/ba5u3g8cVhogZqaR+/33fn8tzvXq/0mLsxuvHd/Ymkbjo9EgBy
rCNVdfdb3/V6T1l6zJuRHhIc5yC9OCnAqwNegC/OWhIkPguZ5HA4thiVGXAKShmRtmKfk5Ww0rgp
HEu1SlrhK2kZpibvSqevx+CzveIMp4CL4ibFWV13VJCxs2DpkJ+toi5tBUVWVpMyL1qhGWgnKWiM
wNaQ0OE1bcbK2a87mRFz+lZvCtBn5fEU6qafoGq1VnyzOy9SZj10YiDVoBjj8ItmEYSSGDaXGFM+
/+joKsdlZEn3/X9LVD4FF/HNQBfzHt34/jjfpC3rTaJj876tVITZ+mQfeOPxfCq1YPB+39hcHCZQ
+a7lMs58bQ89CxPIaSuVroiVbrxhrUW0tHh6Dsi6oxnIR9LPAgj9C6kY9ChgjRUrx6kSTbOXfIph
vH/HCUJB9QVzLedu1djz3GdmcOk1zWXGCAhHACZMY1YKOjlGE5sTGWwUVM2b9mPziyrWU6xFQggG
o1/W1sWw2cZTwXt24AiYOA7A8s8WP+4oARo4UKFzHNJNN8HM7qmW26WHPFJLUdGmesSU6Ndze57T
ywsi9avR8nb2RkP4gB4pSU54mFCRA/mmbrXFxZBsj+g0rYBD/23jNCsk8Gv83Z+rwGHws2t/CGIb
a/v/Q5IWUbhsMd7hexZottoYRQZm5djI4mwwSx0j4S7T8UmOuvu3yIcxWb7rNPWwcggDwdPVbHvB
shic2aPt80d1Bb465bG4SGkRxyZ845X46Ypc8KO2cmtLhW65v7/nJKDlH9f9Zj344yFGq/LErcbB
wXUHK27ya7kKp1z3wIhMyUXREzL7CWY3fLHwicxqhqB6pYHKpIPti1SHEVjQA8EzVmr29hbUd6Pm
zIROGIMTyoi7bdPcRoNKoY6T3pRL4SZ3uXTBEe8RRFRjD32SnE57nWhWHWsW01qcRmm+i0V4uaMZ
Mboz4CrpliRfThGXAHfCC3ID5ElHK22Cm17C+swr3EVq+JB8Uwy7eSRIZCZ5ySDC587LsqYLggTt
luUAZ9et8gMaD66HkUumJJZCDrU8jZhH3F6gvyAzOz0XzAmdaadmjFzveq1Pa0vs46/BuemMNfbo
dSUf2SX2DvqU02PbxXQ5AhvJiD05HAJ4XXgjPQ7AnRXYyCIHG5xdoH7H2XjqntDUI4dqRQ2OhQ2V
8pxD7vFYc0sg/wpizDillR4sAPnLlcK1hAa/PaLRWh9LERg9X8aFgX0LdCfPrWBD/lZGOWtb+n7K
VAFnMqdy5EZqANMyvTU00UsiBDvmiM9pP01GxDPEohT8JK5VMBes1ErnzG93N8jvf/GHHl8ziwxm
MI2EtBB0oJodruwCHZhnV4t5kiKwwbxcl0JGXAvObXTCaTA23W30P7lUFqR0X00Z8V11qvjhMaIe
Y7Nl/QWEabd7Gbb33/gq8lP8/RZkXSgfxALJq60lAwo61k09OsAd4H7K2ZEqIJxIRFOzEsi4Cj2C
MilYhNw8qdoawebSJXkCtzsw1iCjo758Ee+xGJSrWtvQaRt39AaRCOOlwiPYMLiCuVg++P0DJE1a
fXTpGAM7ZQc18FFYozjK3xYBTB6dEmOKPiVToe7F0FJMsL9gT11b2Sq/1NMkmIGXTJ+JZ5DhS7yd
Z+B1bmDDvLRlYZMUpLeyHDWWxFnbu6sR4E3femWCY4UxlbQsRy8dEiPEXy/FoeQtDpZjs070Gml3
25lgnJzRFdUH6gVpqsdyNkjik7LJ9HbkwcQW4NVLE+fmAxLcSPAPj22L2qIWg0dI+8kauDgdDIZW
uVc6A81gcf8B5Kbfi56KT5pql1iy9QOi7v1DW1U2RN33ZQRnIxwTlJN+s73SgeJAU+guNQ9PWaF7
AbSLrW+Aq6tN3+osPmiyNVyNywnzK6kA5k8pAvxF9z7AOfoAFj+dblqf5utzE+A1+wXNmLi28El3
7XGnqwOGyDGrrTpWBmjAd3gGTexrDsnZRWI08bvMM4BR9Af+ENxCc2btqN3S0QbQ3v9fkTL9ll7L
dZ7cPV97awgpj1n6ZSfuQMvct074sIu0kYlfYmI5VNep9NNgsRgIUg0dM/ya0yvKcqCCHVrTkR2Q
ubiebw3c+4Iz9bQlRICxHNdW0hoekqXn+WUJ6W5WpvvnH/+vS/PBJOG2QiEaoj50eRhiaidqTBMO
zbxd2CK1o7Z8yLBXtjTR64fMFTbET8Nqf1UGcY1mKKX1Tb6enqYVNHecmyF9y0PyXR5xdcDSo3Ya
nDyI69tIIXjbWrZPhTrW2woAPmATMwbEnv6B/dwUkZrgBl1m0wKZBIUrqYPNi8cg0eb3IN7i2t69
LodDxggsDGMylMt9r+C3sBiYG90/jDPTiKsELsEGHC4E9x9skmEdvu++9AZK9p/W28bNUfy02Nx+
ggy8YcIMw5kFRvrAZNKb8gRiuvTISK07b1nlOUpwYOZbzHDq8fV/cSINTDvG4Ym2qKqqwTYgpeOT
DUlb5a9G2qGYvK4MhiY88XO0ijDXc5UGRBfeQ2RUbVAr/G6U5kkakqzrfHAmfqLtYDoUx4s8VbVx
QIW6tLygRhLd9pT6uy9149qJpEo6eQ+NCij6FCRd+W9wBNhtVpGehNxdRifUk2RDL/v1l0IasYzT
ZxhZin7yPUog94KG2edLy29aex0soZoE+mfSai9/ych3bCqK+MMt8pR75z2kgmn0EMVpnXqNe2Ji
3SxL24A0apZhOEWpUHRLiClRKxmCYzlJ1eqJhQvN+7mhdv/SpkRxEKPc/e/3sRs1mKtvnI6BEUi0
3cqNO7RvhEz760DL/c4WOj/9/S/mZhzG4QdYG+d6kLv3yOUIUv+QG35S0Y/ybdMkh1StocbHPOV4
PJjpXw/YI6mKeDLOmws0HMOIwxpnUbKO4G5vp1eoO2YgSx8jIGig8mZK935guYYB/BDKie/7g8Ye
TtYO94ydShXobXw4bkPSxOYAPPJuXJRbLRCugkOo1rh33+93tDRVicrZz2WMIMTWI6hdgVylwCTU
Ymd0ZMq4Ihnrqhv6YyHqForVipJVrRDD0jGeIM9cPDjdd14jFTcprde9BbfRfRb9qvU92iR61y3L
Lq1MLv9V17Sl9ApeFdWvXQmIxoRK9jTKZ7fMzRLwDw643YvedYBhv5iV1NwfOh0aE1crcfjAwQIp
uEDbr4AdkZ6KdAZH328KV5f3V3PorSWb4/2No2ZQA9YuAJ8ClOeamM7LwIiWG2Gw9pQWGP9zfUBR
gUnBmeTp+YnZG2sQSfDkY5OyRJI3w0M9rf+XXGrF04EDqTkYhsmgHW84x6ony7yum0YetSoDWcDk
39aJnhl/SIwUV+sr54E/O1vr9KBzn4LjJ6wEVqoPck1tQMVJJtLOS9uDUcsshiqKYBOGmEFAV8Ev
rdcQVH5UDsabX78aj1UVzRiYkInoukVq4xAKg/FN247XgY6sPI+LBlJiAGm+MMu0mVlRyuiH4hVy
ep1XWlvzR9H1cjIl/c3O1xs9S/R4vGTAQdRLt0pwwoWc8ZmMWhDvNhEpP+pfmDlnBH/uK5UGJHtN
K1PvcY64XwuQX8kOaI4CkHhDJDlXEi8NREoZyjEh/elW42+rpOcHuRySCZa28Gr3mgSlKFGECRZK
XBHQz+w1bDhI6nLyuCnRiAyORPYNeRlD6f/TD5ntIkXBgAOjLqtwtpdbRUmmEkdS/K67FVbed/xT
dzYEDUdLHAtEfPyxsbUi/fv9p/+KbVc6JX/1DLRJrHfYMfqi8lov8F1ovJOjVBHnBe2O76epBBvc
X67fIMb3rvFoK0am2YsdaPxHCKnJoLRIuqoG+J1t4iopNNn+v8wlR/D86B4tqbbSl2haDmfJ6QpV
DOeP3BtNhRS3yBTAIGPQXqJ3reh81POVehgPhxCYJjg7E5Vy4EMCzqF8ZMvBJ0XXn8WclIf0QPY7
/My6Se3eWY61Kz4QZBuuIht7xliwh+5u12/0bKEu6Xg0GJ3Oz/zy9ghvh/eU+eN2uz1FWkKYxFvW
qFa0sbxP3gDLHixLyb2S4VdKujGkDkOnFfIvYg/MPruGAoag/7wwhoow4KVNNbJFy0avEXmCAmFF
uukPADfebdeXwGv5rvPn3RRWDSFo7xGwcK9TBa6rCKYBLsjw2erihLwNFJkF/tBAaXscnoADWQQq
xPLVuMxFk4ss1v0mv7TJ2viLbdA12ecghlPDKJLLWQkAO1Cz2wpSETDn22n+3ZOf4M8wGoaBgyMz
CjSWgktH62AfbhJ6QGX5DKATUBJ7MMm5vXNlqvHNYihmO+2gdQ5mMzfDBvDWNCVVET25hvFOsiTO
NBRqqwnuNm1lKsR8EKBndeNNxwaqZeCOC0oTk6szfRpHkeB1HsmCp5s/7ijK7AAq03BhLHwCIIHA
TvPWXleC/r2vb2MmNE/K1aob8/+ofZq15rv1ex+c6HurTXyXf5Pusi5i+sVYHZDQmslVIDFyvo3L
0Hc4aEqXBmLajFEBf56Z+eHZ/iGrYkuBD5GaXiQhuTR2UfHN0jjeR5Z5u6D2R+E/If9bFB8uQPVk
XBQlrWu4XWAjs9AWQEBRnll+vmyObbQz6V5nS36lIlQ6eQR2K4Dhdii7nS5MH3pWfoOzjTcuz5nN
qyjX1PV2RIVNQk3yPuvWRNDf5Fud44CPtSNn7zmh5nQF2byKKRohoG/QNHVOxJRbk4q0gSBAy7cK
aqs5rB4K9bdjMR8w06mL4XKK7c6+/XQezWnCygthSkwQznkuuqsR4ksUL9YUWkrn3JL/hqGFopS7
ZEnD8JITxMwNIHX1zKny5Vyg4PjqoKBPKYoTkUC+Lf2VvYKciT49YOulHptbtHneb05XDja26ATu
9wB41s0vP2ib+guMrQZAp5uZWOw669NTaQr6U7qRVus31L6SN+frhwRmPaBjpDNVS52d3PC1VIne
eWmm9c8bxp+WozQiIM/zk5K6Xhqwd86t3OcHb9+zZXP8MEYofM9Rte2jl4kMeOj67AvcciJneiHj
yRDpkLYavOIlx+hpCbR6oLTkBqvMEWWPUinT6qmrXTF+Mgj/87WWnIiG9yzby2213yLKVJCoHmMS
PkAhQ5qSbE/qqFw6GcoHLeRlodthIQitPGhIfeZm/wTVQPjee2Rm9+5gsnzNvCkTBUoIFpi2/iIi
h4DUuaFkn8LuEkuR/EfLHLIQNxMJZMwhzHdxHwmvHhB/nPQ0jYLW6Xz2/05lFVQTXglZbLOfWKDP
suTw2ZsvWVLyVigtXPP254QO1by775sVadfAe9W42ShhGDJ48u1hH8fEezuV0fae2xxOZdfs5Gpb
pmuyJ2aIeMNPoHcrFU4k591YGT6KrjPfzGh4ajHDSmVg2pkyOMdlkhJa1OupJzWx2v8FOReDICMK
UUk1FF1bPPtP8Bym6LYix7pF26UkS+Oee7BF5MrkTTLuzhVPPiodjJeh12r+1hqvm3/sAbF0wx+x
Y4Luon4Wfzt6b2zazkEik57wOxAfrcCLqVjV47U475vZhBruMoxEzK7BllhyR5ZQha1paqVU7wD8
bXuchcDwgx3C0s9anjRarsheD2thxAn+BFCm6exVLYYDXEC2xXihWrSdFkVgOCMBaKrrDDlTCN91
iasMdPQ0LrEPulSzutAPfSF03MBqnN4OU/MfBTJWqup4Q74XKUrEjh550WEf+5AQRMkN2Vz55z2o
kXMHPVBNLtS5QHL8bTCjwdVZDOPLY7TiqZAO7oLjgHlt8xNmRwYaat+7yE3VbYfb467Jf1KEXKgU
aOf941e9WGhw9cP9ll0JOFNUMATTgltb/Udbfq5ujisyYp+BzG9jKIR53ERjfyILedE1ZXKS2KFK
z3UdKaqjm5+hHMDHqtSZnYxTkbCvv0G0ClvvmJejG3UyrV0Ecz1LWWjTAwZMuK5v2P7EoMW7Jyrg
wWiMjK8Zqxomd9pdqMW+oWMp/Mx5S0OOiFSFGfJPNlbsQLtt4ULm6EyuFulmNcxged+vEHROZoV/
Rw/XazboYwV0fJtQh4B4FeDZNriUkZYGW//m/9iI13/mJO9BAPQJ8pdzBQwqSowI6KRnGlngvX0T
ZiVpeBf/7fEsAGsGvmmN4HqGfu5F12rwPKbcpPOBldQyIf/wYrgXk812ATw1UWVLYtbzLx2/ZNSQ
UX77I1iWsXV7ihEJR5QQaH3e48vTJkT91wR/hKSydTz+C2Hb3nrvGTlmFhujfkbKk8LT0feI379x
ryKdltK7n9QkERXpBjt4VVCiti7lR5B/iKPQc+JxWjQVYNOzv3VB05rJn4kKtRuIu6KftEkffiFP
bDHNx/YvAcWiZb8A7tWFzrTBoPPrQisUi9RlAs86MQ9cEhC48N8A3pb20KdRUEp0efFt6lAE0PEW
Nqk91edYuGH3qajrAqT+t4XJ0cMq8eVxDtJzkBu+nEPGUJ3Xo8HEfhUjeOiLFWE3t74UbL+Kj+0R
1MyJFDyaj4CW2ZBkrO3YJfbFr3eSx0rJAZiGzLt5UPz4iJgAuz/h+wxBw0Y3XuaPpuua08WYaHVH
0METikPvc0onLjvb2qgifAebwcflz6ehN3DwLkTjpI1Hie67svesq0Ki5PfHadO53BGFsHwhQTNr
jy8DVYVkWZIjUzJvAo1vPPDqUJffqX5t9zbn6QDCUZf+nEVdA/pgRC5QkgmefyiM61pAaqVZU117
viV73Prsov1J6slRkfYzcNTOra1IJlmRB3vT59qjRuqluWXTxuPjg0zwqi9gNCvp6VnVRXr/lLgJ
VypT5FnLz03FJNWq14LCwBY3g79Ri/K0BePcixJf2t/qWDr1/1/yw/Yzw9+95xjYMhfIk2XAyZWs
awMzRB+ZrTfe58aBEJg9OCPhJTVjTNTciKbE/6g7itBGPhW6lC3nLH1UO5HcPiqwy/LHKw27XC9D
dmjq0WH/atsjfcULHO+n4owoexqw0L8JoampszVj7AqNusndL1FEo8a7eMZ1+SaZuRO5HcFxOh/F
nhgbspsyBp6AgOggrFDNGvitxgeiiqpx7aqLaJ2R4OKWAhvmuPZ2USmbOsZljE70TgDlvr6oE279
A1cn5/2D45AF7TR5Od5bJzpr2+FJGCvLYPlG2wqUw9DbxjS3dFz6g8bHHxTgG66hkH3YUqjRvQD4
BZNDRzLbGZ4xV9zR+mpHz2yQlBErum4zeLBDfuqhcWdP9TTF8qDAZCS+E+caDWDbr6gcHRqibNUt
uoMzWkpYE0I+IAiJ5YkE9kgDaZx3/k47YzAJfeF47osGsBWXWU51PSC2mlEi7s8XMyQB88S9OcT9
DlLk748LbXZhAuz6hwy5PvK7mgMiEqmSPtpwicNVddtt2wbPca8IR4gUHIH5azYSlD9cs2JAbUAA
1w2wY2/BP5751auQ1yv/xPkhV1PlxS2MH6VvaaOPqF8nGx79xaQNa+99uEjhAsZvaZFbPEWaYaPX
1InbxkJ1AWvOUaVlxohgno+gvvYcaSGokNi5Dr0P46KYoSAXev8Cyu/vlhEWR1qcemNvVVIMJsW0
sFpXjw9slrJ+TGKquNb9xf5kyzd4EezFzMFW0iWlAOUd2tWvIEj9eOUjTf/GTQSOaDEkuWGHmqac
ov3YZUnfCuPv000QPDKAgb1BtvewR+nG8VuiuVEzLN0DdepuYxN6Njnm+Zt41v3yhIO3S7NlZ59o
7s4WWYi5eID3tI+kQCMx1a0dD83H979BXCTJgT/4ihJp76BssDu3sUMD8XASMmDN6PjWnK5S/FBf
5lSWLhS0h/o/DDtIqy6s+TqPruOG+dTgKP38SRdSP39LDi+H9LUnJU9P39ejpyv4Xe33DyF7rUjH
BOvpN+fXioklwz89zWMlJJr4xSb/XFJRgwkLS00KZYujiGwLzcr2OsGrURQvt1nwEpyYXl/DD+TL
/gixXaUzRBW2VDLOxr3EqhN9GfLy0oo7t3mpDxcxeuOqpZgcZYC9VMqu0EWwUreVb8EXCeAd/NhK
v3+tQXiN4xzinLP9Nc3S0tw5i3Hg4iPSHIjcnpUULH6OpLFTGletlyeL5jL87Hif1v+ggRPgwFeG
eM2gJ752o1JUyNq9FpHou+i3bgV34CkZPuu00uXrMvyFe3D1P5RJxlG71ilGZC637hGg5mByQCIM
JBtPiIUzqEfq3A1iTJF/45amcCBiY0EIBu/TFd6QpVGW3afXKitxKZ4r5XD4YHir72X33ymqUau7
XCu+oC7UpvcWVglYTey2+d64vEmyqvFzdLJmuv0iR2S3QKFKIWIxNyCwg9qGSZQBVolcwQXX2lbm
5YYhA/DtNXgSzbV3MLdUR26gNDZh2ZuTDJz3T1G97JQ8mEslAG/Ec6TonvbSgZjjLTx94twreyxC
eIx284ycIAN93pCXeedz/x7G3/g+PhQfA9NOaP2HDJfm3Dlm7dJrS7x+ACUYbf12yPYBMS/8aRkN
NpNwG6L+HUJIazmgQ9+qO8ZLz/HKkKZCfPaFugBqr/YJy6J4wVkG/kknlrpHA+6I2AbCxfdbGhnk
dFlDD4iAtST2vX+QoRoLkaw5MBfC4tYG/SgUDjkwIxRV0XdG7ZXKk4NKmPN37kgImyoCZ0rWwxIX
WCXuZYhsLIPW7VjOFxJsPZCybz6nmA+roU5fHNQwyt8aUXhniiBBbRB9/Bg6TQ/jRiQtT0x3M+KE
+lGTfJz+H88X3UcV4/G08MAoo37E8USqJ3rZII1D8559aoAZYjg3EPBQFdp+qX/cvUaojtUhi5Ka
dtjLpLz/vw7dLDSZFNG9kAWUoyuybN4UJ3S370YpCl+rL2DyLTEOzPYbI9CI31xzo53QMjpiGqIG
n+9o43r8MgpeL+puuryUJLYcbLOJS3ojqf05KGaYAmZF/rwOnHZRfOBA2P8uNnXFDdrWh51k6oAN
Z1FNrqyRIuOy9ddWGLFLAA5RFU45WtGmHOLVoekOEwOBXzIgwkIEsSRtUEjLSN0zr8U2X1nbQcdl
VIiujxH4RxO4qjzSgn1esxr3/Sp1h83EoFeRnls9loz1WZ9fNxlDn5fW8xL/p/hX9RLkws2EbkTG
VJUqFmxD//xZf1NLKIeL9GL/+DvueBULiZANKPhAgY/Inovwejj229vlnoRkPMneTWHgtbL+Jt/u
/mP5jARytpfRE2N33KmGueCnqDM4rRKHVhBkwWQjfnt1wALKQQrFYUeaVHBs8QPvWl/Wa/s9Ea9b
6HlU6tAqVGAhNf3qgii/vU/YZDdnZ5g7TZiaeBwrIxUbf0jtFvVv3hyCB3uS2qc6tqHkh0iuwC+u
qvyUCGZhhyU8DUSv7hU3E4dHjZefKNxo2ozYDSPugKsZ82Tr0r5XyAgBrgp+li0aELVizD8VON97
81GgmlHnQzqd04EGNuOqvEfXb4kyTtlymghxBuz+4fb8eKkRnBrkBIwkSpXgr/GbZggE0RF2wx94
GpygWZt518knKhb4odSjPCr8dxqsdkT+EAt2O5fBZz/lLyiDOatMFKZoX4vqz6pe1fCTiM11PRUn
ipz1eGEzrvZcmO9LpuQQO1iIaj6iC1OCZQvCk8W7B/pNGiDzJU89MGxBbNd+Wh7wd5xK+vnKm3xA
5F48/KeyjS80TdGu3VWTqaVYmYX3amhMcX7MqEUFkuN/ePLO/PrCInYZAi0InJf7yvH4vCM2Y4Cm
7soJo396kNGAY0oHjEFoVASPLRCq2frIcRfO2Z3da0/Fv6LQll9DAje4NSxb7wR7CWcxOS7N79Dx
jFDTEN5BNhjdlmLYzr1SkNkigSehNrLoyEy2x2oUfzvqJiFHRaZ5JRBVN1LYyxTfASayydfgV3+I
qXGmNEri/7pHbP5roEP7YTx0sb+wYr7IdTp7NlvbnXNzqlTLZBRO4jlIU7BSNo3Ah4YzIqeG0nQT
X5+AeDoWMwqlUpgZ2pDl5gcXgDLVRdK/qyTYCQ5sxhdaMK1LwpttarOKEtpQXwwWlwsHkFFSVtDW
TY1tIiNVnXQwiI7tYvP8Ox2rd/ulaOrWHObsbx6rMDemOcbCnyQ3et7e6pViKuJtPqvtN+poulK1
Qu0zG/1Izd+Jc52zvabb/dVZmlZ44rPXFHSISPQx0oy3opz9P1sFf4yNEdQldf0voQaUqFvqkU/9
g1imgX2aX3pchZ5at6Rr1eQ7fvVJxF2oqIJ+9f/7jcw12D15rS/DKMO1haW1+ZuP2N8sB5k2ddAK
ldyDgbFeGjzEQ/OHTvak8qs1trp8V8bBj1Mg9enP/Js4tkKikctmzerMSPulCVbGS0VN6f/bg80e
oKLP6NyeaejxvczJDHaK9HVCYhJl0cDZinXKxm6jBHmR1O4CTOjoxuADLnjG7ZrKcqo24XIQcEG+
p2mWcCYjuXqtIFLlKLCfWZy687+jT8lFtZynJexLfBuo9TQjoR4/PtmV07D9dUT+tNY3vCQ8lLDn
7ENB9unGkOyDfN46cEP7zaMkULN47Dfs5LGAfAInIOA2Opt4RLnKcQAq+9owIEO+IEViO/aNbiJu
uNvBvV4m/KrYsW5IKI6UFegjRgbHSBUvDtZ8nNpQLQAXnCdknH+ppDDuxYtaT1+awiMIowwvCZvn
+957r/4GgeEqkZAu89Fns/Fx1SX6x3fmISR+foiT6GY61WNsd8mh5tVInSuVYyDsh+CfNMokTL8j
+Txfqnhe2Hr1iv6EFUQ8LO71vIfwX2C5ZIOOj0N633AgNBKUCqwiZ+EqECzKc4aIHlL4BqmwdpDS
Y8goe8KTmHP13GZYqfpb+UgHJDLht+J0f/9HjE29Sj2O42xSehyJCCFhR++u78977bqDuu7pWm0C
gNexEtbu7JHUudfJ5Lwavb+O6eZfNv2fJiv/OiTNAMua7R5SoMnWLnInUe8nym9hCozYXL3peUdw
ZR07UR4qwwWVHTWxCyO/eAce1GMaMjYjjjmrbK9AURYiZ4wQbxCZK/sgijyU4r1HGyzsGorFY1ja
1zVIEHmQxa9ucoqELptNKTXVONRdLKA+GGcm1d3n4o+xXzlS4iPOCl/BuG2nNsEF9hDDaOUcc2wl
o2Q57isIZhyUAUtOpf+5uK6QqsGX59MXZzqnizqqnDR4qV4hRfoNaNtRKdeQfLZnmJFLjPN+GZ5j
GrP6Tak6uq/+sk0q5j6/5o454TwUUzN8mTnrhMuHoLBGtJeVjAVZWtAbzVXvhdT1IeJrd+SO8X4Q
IEBD1rBeu7fiNlPQ6L2IZpXgii8YW89/TbzGkpe/m3BzHLlJVjGAp9QDG7nTBJzq20saIEICKVW3
S9hJBXnpstRNxEI1S0xvVT7aVfVeln+N1L74mOp0w7cUH/SNta2bSVCqMZ8H9ZQ9TsSG2irfyNGp
velrxRFTAfbCNfDyil7L0aBcoaXjujIkRep85He2PypsGHq1p/BCqol2anX/lSb1pqM4NNCKiseP
Yk84nd198LQ65WYbOZNr6ZPYTsMuXfQuvEfVj22g8IP2QpnT8wcLoysLTstGep2wRpsC1vlAdxwX
RQbKMmSNSFv0Yzfh0jsVrWtpLv+vEPyml5NvM2Ga0KcpmUQX0NhaLlX9NXVxlsXYOdGzyKBChfxJ
YfSkj9x+tcGaC1bbrDzCVAOqdkblOIJEDD8TQfz2QPecffN0yQhk4X8/z4fXzCsGvJ1iAXhD4/XZ
0LsE+3pcpyRgt6DOkNZ+nbLZv1JHWWHPVBSNSrZdx7h0Oniuur0bKKcxofrs2KD7sW4WynGipzqq
nFss+pyU7jq6uH2qPg3uQgz9cUU8ohL8oDMEiyb0wA8nKqrpIVeDr/F21XHs2D8vI9dl7pO5xlwx
b8pIjTLYDbbDfjCq4RDOILmS4654s4P9TGuMjJVK4Qmlbts9ncAM2/6r9WDLHoD93pMd+fzBvOAc
wRaxiUZsJnTH+opV35ZY8pXX4g3288CwwoVnKqzEX9y9zLm/GV15glJZPMJ2dDFbnyTEQ5nY7M/b
Mk+6M2dphQ1f8wnAoYqkn6qE7uDDNL1rIxPjTFSuMUj+ARHTw+mU0An3yP3n04oQdPgN3X0Me3nm
m3oudbRdmHpBxOOjjngr3V8zPh3w9+r/XleV7lMH7C4EIp/r/aWwlmv4xVUTvFlbiJOyv28/LAVa
C+JkdVC4atj5URwcmRKBETh4ehhDHoUoRmVKeZSJD4g7VTzsKpKDdamBNERJUBU6WUi1P1/cGCXK
b1pgnCul6VF9hSIXexx+9YOmaBVzKztarLVMVBVyW8v1ueDDEn54m8BD014ZRAsxD1Dy1RNuL1Sc
vr2hUf7ozyRW55e2PfUAmg/1Tvqwtbt7ijloSttHVtHoNQ4FIqJzYdIORpKCZSTs+g89c2amGzy/
77PN/mO7JGaOREX+D/yytnADfqp68fFmYfMmxQ0Ic3y4JOhQM9ENYAL6Qwd0RTPh1hV4KmfvZVOI
ecifBNDvVlN8HiAv2aaIE2Wq0nE/omKBnJykKBdIWm2S8fqZlXa8wbk6c5csmpsh85ytpBp3duFN
zCB/UPyoNWCNGldCq/ih3/N8ojFrabSVtz84ipvndsFi6MYiS3mSDsY+0tK+UFLtME0milXlek7R
wofTmp6zK3oa4QfChHec2ubpgYr96sAvVkknOIuAI9m5Qfr1jZ2sdz6AEGzYauO0dIV0w6ue8U3B
8quJAPYkHUzC3hpX2JTUB8y85FbJHIJYea6AfhiGrkSw680rMGtBqtKg8GiP8rgpmn5VkFVhxoqI
gc6YmqCHGkPc6i0VEGsiURAS4sISoEZfYwK8tMq2hQVfpaHZN0W2B76YMSTTja9ZiYwmSBKAUU9h
ADYOJ7xWBYuXnCW5O6I/UOvdrWI2pqgV4YgW/12fgrNBG8m664WDrVXt7UXCVIhOTlrAaDK0Njny
AYZfmZHNDR7y3Zub5sXWvOuYzikeBASnVj/7ehdRCGS0gBXsWDf/OvgIOA6x++iFIpOkAuJMt8rR
04hlMRN1vKut3P0vM469R6TgP0XwywFhYLI47aUOTbG/TCmYbbuMwmWQpMLyoJslEcfpxbP0gRYH
3XwLeajwNqZewOYSNLsoRgFDhneejzBrQdhOJmdSmJtwzQ+YQZVVBbjF0qNahEjKRfvmTCL5rkv8
8bD1SeoVL4FyZ2o62f2yCuflweaVAZQaBpwc2T5eAkr21owdRQnFbQs/agAWxtfZ5sYoItv5fw66
TKGuqDpkEdo/d6NLyXxHxibG7/rV9+Eawo975PriKqotPgeJ6mofGveL2gWBqaxmP/uSDqlO7MDo
eVy3lzZ8n5FJNlUTfOzlPQSlBd6G4nkOCw5OTZ4iKI/agx1ZoL8wIq4AVMvAEvExoz1DdIKI42Gi
ODGN+iOVRwxaw6FtkH6KhqsrhZzzoeFDJHSIkbJuNysz5WT9y46+ye00LIjJWMge+asLJXEF1Hla
buYOUDdXHkGaxfEQLadcrbunPtsD3OIc+pSf3MZowdKGnCFQ/575W+hN7md9a0ZyKdxI7sVfjm//
pEbmOj4vo96hW62iCLfButlbxyutT2Zb3rszpuoXh8BLepnuVN9dNPBKS2t8a1U4lBcOeHnm9HNf
6uVCJw60bjVs8OZ8xxhYT22G49TwbIfoT3Qy9pDhPzJ73fT7c2/YoW40mcxso3qdoI2Ec9tbJVFV
v25cEnOeFdGQedy7iSN3IqUsYGflRckbdX2tKFRD1zjSn3l1YJVquq2fr64VSxM3rNMaOKaScTIb
4K6Rn/cs57kxJUDe+P1jJF7XjHK9G1GUTqpU/b+RTMOIGaI2YIoY3AvX52kPF6Bni6QFqfzBQqm1
KZIjI1zvTUlg2woAN1DCqutcyx7taeKh3NJ9aawohMfksHbSj05OSRFhXQkGrxsK8FRh2g5B6HQk
wbxDP1/8tClPskv31A+6IUCwG2iiFV7+Nu/zxjd3nwG+BxEn2nBHw8EnXah7mlBZE08Q7/6PupD2
CSNfaApWb0DhK7LuJGI+X6uRCMQp5MRuHPiTIEialQqZxYOY9er3Iu7xfO+CFKaQiXUSs611mEtR
2I7HtccRYwFlkXT284X+lu5FyPKDmfoVI0q3SksnOVRh4sJJDhiO70xPkCaO0dY1FK9wfVOFcndv
pXYvyMw8JwnZqZX3Byb0RBy5GetAbSQn+d1gc2xJlxb0EqZFuZstG0EXgh+FXevaNTf7xdGzyvbu
3UHVFcetJmLim2pCf4TXa8cFjLGT0R+N/OgxrzhqT0C65yxSV8GQr123jG0baufcP0dkEnS/+uZp
W92UBJAdAXLl6Gpiz4JYLxhKvzypcfVLKvEHdUoWu8R5nuXJnwx+KXyCuvpLFxQjG5n6Q9/dU/78
WhyOEeOSFRV09Zy1yRZO+fNyXert9N1tmIoZrc/9QgjtLEcP+KDzxcz0GPOhnjFwllPB7jG82qHE
z4axQ5VHRHVH3cteo5LKCES/QhjTUIDbD5h/4dQxgwgud32XpTpAkE//KzQvqBirsVtGw/VG5nVt
uZ1QlqwnbhUqSGUpcgBB5I0Aq8S9rOuqEv3p62a+3d+IdedZsgPSdZTwjqBK4R8K60wp6/prKmHC
2U5mUZihOUbX2EjDQ0BGKT+IB67UjfVuuUYipwP5tvn26iYx87ClbFRgvs+DCY8pUH3JAslN+Q0D
Pt5LoEAdArnC0g5Bt30Fgjoxq7drcaruKJoc5U/2eh5ul53CI9OjZit1K4cYYFVnVZnXDDSh6FWp
jPIyX3CquYmYrFbIH0UGG1MQSAUxWxTjYK9F8SKrC0sMu7TFg+i7rUV4SPqzJZJRQplxZoPnk1bG
mWM+uwMTcWgPwR7viKVSo3WIyXuGhvodSXSH8tPBefeuQWREVrGbEBH+EkZ8HMBZM/cyvjumCH+R
en3AmFNx8uy8OxEwtT6tggZVivgL+YQd2M7Wn0DElNVqQtSHl7CV2OrvjIcGwAqy/8S2LK2Xqt+b
1HoVClTEYb7A6VV27XrAnKNldh29898ip9NjUvGR6hFfw2hoLG7iWHZ7jVEnnDgBqsET8QDZTd+b
+vcPX0sCBgDdqYA/GslEiLdLBmzkwBgg3NVQpBVIiV8TdrMUanjKfp0eoUY+rMJHH1ohZgtqV9lx
ON7hQaCQG0HBQz5eh1NT+3cWtmHxDcqacCfgWv/hTYVrXaBViAoGqzu42rohwZ9MJ6gSNjBxhr7z
XuxPFzsqPswAp/yNA5rkhz8pxZy23RWyVoaIPRNEg2QG1BafCVPpjtXZuSj8dBrUdfBd+C/Od+UH
zrHQW3lfsjtRVsC0IKUQmSmQVTb1+vQIiRxVcDlLQPn4/euPuy6iYVg9Hk2rjaF6v4vSsMumjTzK
mH+0fx5v+TdII26usQ6Z5HWJXLMN
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y�BE��Cp*��2�==��Ȳ����z5�Ώ���rJ��`wt��y�m'�vH��j-������>�9�*��>YQ�҉�1� �pLs��[u�4Sʱ�eFWa���VM$�J����#+�.F�ۙ܃:�t�`����i*�m�+
z�ު�Zt�EN��Đ&�n#F|Cp�$�}��eˌ��
V?G�5���+�C%��^y_T=O*��[��iF����X_�"y[������ �Z}����uH�����d�_V�Rv��]��T�t'�>48������L��(�<�OG,o;/�ț��.ʁ�&, ���]&��M�>�7UO2�Z�R4W`�_���]wT��(�j���䒪:B�C\�Z���:�T���2��Ϛ���^�A���z�*�ȇ�i=��/�︳kS	�����٣/*�P�4a��`�v�~n6��嶽P�D���]���'� ,*#d��Wl_����)c�*0��|y{����Z=$�_�K�H��i����뻚S�� �C�_�/H�Ir�.\X!ّ:M�������.�����Pf��*#�;Fҩ�>��%i��]�7��ΈT@�x�ܹ�Ƌ��C����e�� Z�\���f뒠�������n��ĭJ.�mwBA"�����������om :����(7�z�4�[�P�MSt��ɬ8S�>�:���i���}`g-�������u��VDס��_'���\X��&�/t�2�9�6YYyst!��Hڗ�jB� �m�Ӏ�/�����Gx��v�/�E��)�(���]���\W�>٠d�o9�غzRT���5�*�E��r�]�'���a��l�YoǪ���	k�[G<��Z�-<U[ ?I"��wY����<�w#���!�9Lc�V*���o��ޓ�M��s��!�n�{O⥝�������w=B2�;XJ��:B��FM��U(WA�Z�6Yī��I|<LI��������ݭ'(���fJ/�LQ����ll>o���Ht�q.���x�������Cx ig&�iB�Tp�,��'��Z�Xީ�4�.����lj��0]���u'��q�hG��xm�.�ͼ��Y�ǖ���d�=;�v�%�H�&CG@�%0w盏�8�6�AM���"���l5��V�T��~�u"��~AGwߤY�ux�������N�;�ˀ�%���<w�<z~�?�I��N����Ux�K�x�x��Ln�S��jR�O#Ti�||S�a��k�T�x�N#���E�@��@[�.A���F�|ź������F�����!
X�(��&|���E%>�j`#{�����xӒ���`�T���p"�|b]aG����6z�%[��s������ҿi�8�o{B�SnDmEF���4�W���a	Q��L3r׹�7u[;/ģ/Y%L����Ѧ��&I?� 6.vOXR=u�8�Lp�6�0E���nv�-�*����	�������6�Wp,��J$�5�Q{�Bu����)�LR�H��v{w�Z���N���x)�%����$���3i������`:L��/~�����Hr�2�D~�넰�	�Y�?�-Y�fŧT���ٳ�:V��7�ґI�$a=��@�{���*9����S6������
R#��Ό�F4��pU��� ��7�fF9���q����m�9������B/�^i�(��R���t��!tJ"��I�ɧ�������S�i��#q�F	�ȱ�N�ՒT~#X1�(���4K4U�eAQ��c�{Ԃ�>Q�������� 4�4*K��17���_I-�d��-e��EGM��ai��/'�\X!��V��^ʠ���G	�)ᯢ*�hh�g{�L:���⶛gg;�`�z-�2I�=)V�H��n{o}'ÿ�8)�W���ݧAs��Rq��+�S%�)4��҉��$׮�L�H��ny3(���B4<˓H+�r@�\v�=�X���J���~��T��.�|_�cr�	7��<�:���(��K����_�Mմ�n���M�i�A����$�8�V��r��f�q#\���
� �����&�)�	��J ˦Ցt�Ez)�h~��7=7Bb�J��r�?W��&�P���rL@��B��>V)�{O���L�%Gx�=i�L��|c����Q��s,ء=�+�6xV��[Upc.(���}���#�kV�s��[��O���<[�k$���&����1�Ց" J��6d^�zG�¾�����4Ko��5�Zi0��]������滐t^�=��TD��hoD�#��/�瀡ݤOme�%�{s	���6g�G���H�`�(.1�JA�y7�m.̘����qޓ��Uɉ�����(V���5e�}���N�ݧy���s]?Ѳ�#-R�OV#���O�e�(�)B������!�1�%���6����2\����IPU�Ν���i����	�c}���	�Ķޞ���_� �F�N�T8�}{+(���$���&oh��յ����4�P���:�� ��a*Ø���n#/ʻ9i
@7xAth51Գ��k.�eϷ� Ч�Ջm�J���$��#J�_��N��ٞ`ek���Rb9�����,�nnb;�Q`�;��Z�zԩV�ܤm|y���}c�!����E e^33�����!t�����_ 
�+��T?S�oeL��(���D��X�JAح��y�-	����V�ei
N�� Ks��9k]�ve�7��[%lY���f;e�UKQfJ}ڮX�^��nB1�,z��#���uU�Ó�W�1�;�3kkG��1��v�_i=�/\Sh)���D���Ka��!@��p��:
�@4b�^q}�����z��!/��W��gU�fi�3a��_������K5#�
��z�;�N�d�)5,y�<�S�ִ|���2ܹ}�XS_���*�o�1�7Q���?ƻ�a`���f4.=�C��0��^ۮ��9p�������$����D�;����wx����Z���#��`!*��#��^�^2��\(HsI���ܨ�P��|��i��p��V^����/�WSD�3}l�h��$%�X��@~�'��d�۽ �G�W�YR��zw�6�p��V��
��x]���}�
�����#�)
@��_$����V�Չ���Pn��+�?`�,�rm��r�8�XoV�2bh��G�Z/o9��Dtw��	�7���H�d,8E�%���5e|�]����yB>Tp�7O
c" ��J����o9��CV4;իpV�cF�+te��_~�j'n�)�rR���F�}�DD�o����P�g��#��9�L>!��`
8�\53�����s���.6���ɟ�(�u'�!J��r��w�ώz���@�LP����:��1�;��K��urZ/�8����?~Ot�Ԋ�D��В��M������7��3����`3��ӮS��1ց�|�Ƿ�b�2ŀ��&5�[fs�[)�8���W��L�/
��3&�B4Zd�ԛ�l��D��4ʼ����c5�D��H<`K���	u�!_lp(O�.D�kr����� ��Ǚ\�  �P�"ó��F�wY�����z'�'*���u
z�%4+�G��gt;f�M�y	�ݺ&��+��'	)�\���b��]�<tLxn�d]k6�pplţ��,yMj��y[0 �WG���z�!���S���Ns�KЌμŀ����A�g���31a��6>M�wj�����?�`(�L����1��6�I-�j9�����xy�����M�/�|�&�ۧ�5�D��>H��w�uW<��w �ԕw��(��#'��8���-�)���o+��%�y�Ϧ,��t�.w�s��;0V�@���q�d��$�@��9�wo��cs�tƮ�7�s�e�zi(g��-�[tZt�Z\���������X��l�<¬kh���)����G2���_�f1N	g]¬�9����kk�C�S�C�Z�n��h������̪;_�6���(���T_�$h80^J���"�`��tE;���8.%�f���Pݪ���S1�S�����Q��tZ�A�aBtU�6>��e=hu<.`���(- r�S�VDr��+l8������W�O�+�=Bh�8��j���)x�O�� s�a,��+���|х���p������g)�@h��3E��o
�q����S����A!D�Y Y��fGj@ų/\:bEi�&�_̓S���D�eG�R�}�'&TgSy%P���e4uP�ÿNL���6q��GI7N=� �:�q]Gr�TQ������!ڱ^�.E��rQ4�͇��q�����P<�_	���u���2=ʺ�/ũT��p}�`&����1�A��`^@ׇR������/��Y�Hc����פ~}������dx�G��$ɴFH�.tכ�V���5<H"`���c�Q=�r�;�i�=r]
�R���-`r�/ҙz�ɷV�i����~M^��D�&�mnc����*X�wj�3��V�[��+��*�Ư��� _�a�5��f5�*>����/��S0�iRsc����m��)4�g���L���,���ng��H���7��(����,�֞���W������J��9f��h9o�E�\�����n5G�$޷�X�A#��L��c��_3F���skz��^2����3����-:N���@����������ƶx�,�/a�����W���U*MŎ�RH�y �P)5�Դo���=�h���oDn~���R4-1�N��6C���")b�	�Y׈|��8�?Y/�
ra���0P�l��<z�&��
��M�ԅ�t�����X\[9�/ �k�-����p���I�����d��$N~z��B5"������BrN᤾�����ض�-���(�V;s���<�d��n��g1=��Q����F�N]��Ԥk��j�3�4Gb�W����s�C�ثqK�ct�SA8\�X�6<��	�-zS��@3��'P�Y�Wb�;���\�k���?�
��"�Up�?���3�|64������}�{n}O�����r�@�OeD��G��CF�űK��|�+��,����`(��?� xi��b��+��y*����q��|c��hT�9q���>Ե3#�|��8A�暚c_~��)E��(���t���/9��;0�tUo1gI�]f��.Ђu�/QȽ9�K����vͲ�Dd�	��y���tdv$ѐ�D�u�8�k��Q��(a�}4�[�?⣺���U�Nr�&I�nJ����[�Q:%�q�`@�;y�?S��cU��=���=�e�p���� ��?d�y�e�Fغ��F��ڣ+�Y=S����L��g������:��E��ݛ��Z�ό��&2צM�7�9���u^F����B�AX�8ß7$%�ː�<:ϴ3A������f��.
N�Kڙ�M���E�K�}�ce@��Eq�𻐒�\�ɓt�� �-({�e���qKk�D~t0E̶�.��M�*+�=�5�4@������ ���-_�k[,�Q1"��Z۔ţ�����D���<z����l���܎7��4�B�����ꁋ�p�#���Y�)۪�~> ���(�d;5��,(@�����oU1#�R�}ՏK����0����-���GLv�K��8󁂢1(������mpb<�dt���oBX�3���P��Y�\@�D�"�J|D������#���<+�h�xvvø�j�����[�%L6�w�{ͷ8T?N�ß�NR��#�o��]lz�&�ܣ�EL��j��n<]�yH��+�߲���&�r�N��h�n��/a�����CDze��t�pQ��6�t�)$�ē%g.v)���(��Һ���@T��F��-p��E�,!���
 �)f4���x(�ӣ������i�.��d�#JӚ�6���1	 ��0�67�:@�#)����'~
�I���W�T��̨�n���n����Y/�K:�*�<�Y����KPs�?oFƧ�u����kcT�.���u������p��6_##kgF'R3GF��!_r��*F]�dP����-���|���w!�nr�߇PL �S�������^`�"��#B�)�T��J��/p;S8=D����"j�Dg�l��vH<A+T X�Efƾ���5D4:!XC��t�����Bႉ��E���lC9*�d�y��~��ꇏK�*',8��W`����=��0�I�w]	��Ӆ�;/r��87��YaQ��N�v8�_Vs3=��1��	�YԺTr���j��|ʶ[I���Ҟ���u�kAM�"�uȸ�%��OA�l�za��T����~�-�ŸM_��i �8l'"8� Rm���Pf����L����m�F�BL�ݓ孝-������t/\��EihiÆ�X�#������L��K����Pe�����i�lɍ
���y��+��%�9�r|%e��/sd��1�s�;���k�>>��j�jR~i��%��+�ri먮�_���{��i0BE���W!���M@�~��	�ol�ؚ��!)'AO��3ÍsX�	� q�y�����G���"�5����P�ӻ��(��_�˝�bcW��
�T�/\�B��UdGl�t.�fV��J?�z&�[HE#{�S�.���T�'�G�Aj�.�_s=��
V����T�ॵ�X9yE��ߠ�I���7`����uR�uWS����ï����.������?5�=�'���@5@C�	�$q�����s�r��}|e(s�8�����B,�� ����
�l�qc�㝏�#�E,�&��cL�!ٟ���fA� �OaP>���o���΁1u=�_S2��tpGf��::۹���]�R1�.�{2��!u C ��MTZ�g�E�F����i��[�2ui	3v�P���D%�����P��&ҕ��Q&Q�_����uC/��� ��@�H������o��招�-��uR���� V�΄O��;�#�T�Z,no�j�����n�{����ҸF��N~�*8氓�U��1�c2.��h�4%���}g��N~�^0�5xd@d˿�{,�IK�D�1~̞Ա����sTTaS��D��w����h*�[�W�����`lMT��S������YA�#+��	�y��H�XLK��ɾݻT����ĵ�n��WW�daԿW�ǐ�c`�i༹��[2�">sO[5�N�V!RTK���]���rq����W��K#vm�ʢ�hϏ���U	�II���>�3���A8ӛ��5#\oK�=�hN���\��@)��.e�~E4�X7�e����c�Z��G���Z-�M1l�S��l;�>>qC<O�>	�>�R�:YzM����_c{�锻�q���(a���8�}z�>*̀�wQ��?+zl���N/v>|󨁒05V! �J�r��¡bFR��W�q1�}09���J��,�ʿ<M~�+�$��b�*����)�$�/�o�^:��.�x>�������}�#��
a��݃��$�@b�	0���8ܱ~�	F��sѹ�����z�}�����L��5EEKW�s�˘����~�)4��|�>�,�
�+��� =R�� '���@ݽ���7��NY��ݢ��r'w������L�(�_O�8s��&)�U���7U��<�a�Sʸ���^��GJ$Ř����S�1o��h0ᠪ�9^��P����6�uX�@�޴���U�l�e�6K�������p�H0�΢k��gjs�"��p�is�{ba�b
�j�[�&���-�<'{����Yo����U'�4��*g�sR3�=��(F(�ޤ<�=��%>8�i+y$Y�%�}MNu�j��G�^dvʭ���2g>zIGO�}�A���ϝL���Z�Ǜ�.��| �6i��Nf4:��T��\x�ж��?'�Efm���e3��������/u�Aom�Ι⌼�-�A�)2�3�g�&Kn[����QTznX��kQ���QX���+)���=ZA��%����K��A�!��e��j����q�I4���6\�9�R�M��Rm��Tӫ����
0�>�jʍ��k@V��Z/��>0�o��6�x,Ti�\d��N7�sMd>ڈc����Y� #�c�x˛�R4;r�n"�y�|}�?��rE�@��b�g����	
�v@��{�EsF�j��я�k/V��Rp(AO`���䦵��u�SŌ�S��V7�v�~���J��}G�}�٧W�}��ġ�����&��CJx��_�O�0~��km�,I�=�أ!d�&�Q���[7s@���:�
��K���we�9$Em�/p��)[��[8�:^�Xo���K0�#|M��bAE��jcd���v[�TJ�AG�� �G���D�����`��PUl����g|N�M���2�Y�߰N&?�yԅ��AqA-�u9��NB���77~�.W ���F/����=U�H� P_(���S^8J�V�#cz���ia,SJ�+�H��S�����Q��������E��,���q��$ m�<�;\׃)#w�	�oR�"�������	��Ђ��8��8S	��j*v.��AlQ��^���Q�~���r��.�g����(���,[�\�����J�|Y��>�zh����ܑ����9�(�|����tiXn�^�w�J��n>䑐n5��<Gr��l���d��(�R�>������Z�ܕ!P�|,7������B�]���֩�D]�0iӝ��D<�H  va"�rQP���5���"�$�Ԓ��S�Adݪ���L��x���P+����.�b�BܚT ���Q���nD�� i&k�]L���6lb~%lpmj�g�M���Jh�Ƌ�i9;Z�҆��s
WnU ���ӴZC8[LY�I*Q��EWv�N 	q��t*���k������.�\iT\0&�M�^�Ҕ���-���P_<�� �T;������s<Ѭשg�3���0��)�S*]SVJ�n ��=ф�Z��ȟF���P�������᨜��|��#.q�đo��r�K�K��n�H�%F�����pu��4��(]գ�=:���k�(�cJ�e����'����b�q~�x�`#i�䩍Z�M�['��8��%G�8ב[�NF�d�S�p@P%'�P���g*β/��3�i,�gŮ��>�6�Џ��;}-���8>���ԟhD0��U߷�՚
y��:N� �խ��S����CX��-Z^��6D[��K���ٶ��:#1Z�8e�)X��ym�U�mH�o�W�W�]��)����i�*|�(3��N����o	��?�d�gdՈ�,��;F�s%��-��G�>;z��_<jEy�%�{,��&�:�Y���O��"�h%�O_��G �n������8k����)�h�hs�NVG��>"������T{�D�y5������Ѕ�{�EM�O��^�~磣1�>u����XY-|�Ɩ�~f��M��Z�fr��GڍR��r�lF9�E���Z����LN@1�Z� G�U;f/�菶]��'HvЙok�S�y�mkB����NX�f��������7K�!���#Cx�V�Fe$��Nj�5�Ǭ����#�iĭ+�ķ�p�O�|���p��@���M�k�X"��������5�U�-����q�҅b��#�:���A:P��V&��p:�ۣ�_����f
o@��݈C,o���P����g�&� M�x���gIL��a�b�u���;Ҡ�3^8vb&����5�;HUivx��cZb�݁,zO����ؕ�����(ů4��a��G�@��I����26��%)�@��5�&F)b��F�/̍qe�)��)z���w���\5>�1ۂ�"��o�}iH����I1�o6��HG�&�;n���G�.�� �����x���=�e|�h� Wb��'�;��e��Ԝ[��D����q����d}f}O�����%%Es���v�H�����C�*���E�\� BB�@�5!K@7�\�8Nx�ܚf��h��U��%�>�	���Z�H���M/�Μ8`2n��||0�4M_و����7kM�N,E��-�5SAT4/_��.��8��4[e��Q�����_�̓f�H��.u`���Dͽ�H5u����c$T{���
r	&���B����g�	��Vl7�)�b��տj��Z�c��b���L~�r}�@��GG��P���-�X?��&��Qɟk�"_Xt�~W�����*���
v�.s���S�6y���D��BzA��Y�5\	n6H��Gʷ��|h�nm#&��qߩ��AD�ߜ�-�o�k�|�#V�nY�ڙj�iH���s�N��t�%��	^ǌ��1��x����D�"S�j!�ukHa!:l�doKs�w_�� ��k��:�y�Uz��z©2�B<�"j!������	@�͞/(WBSkș[|�H�ҷ|F�!�Yo�8��O�vY�����t��M�ތ�T�5e%� �^g<��S/ףiE���LkѦ�KX�����>�_�M��D�Zml��iރsw4��t����{�˒K�j�ȝ,���:l�ͯ����o�M��?E*L�ǜ*��֘�"oHL=�ɳ�����8�M�p��2�,��M���!3�:Us=_��l%Me�3�����|�:Y�%�*�d�)sl��}i����:���
��Q�u�3���O�S�t��{�h�{����L1�~)bZx�SG�GIe�"28P{���[AX�z����.�y���G��x������ar�+�I<��!/i��W���8"�+&�fdȮ�f�5:�/b��T�-E��&�>9�|�3Ȟ��Rf�gy�Qv�5v��4�2����91�9v���8��'��g���)Oɣ�0��]�2�`��O�u��\����;H�L4�K�[���7E�T�\<�5��Y��^`Q��GX�ċb��8�kSL�QrY����\^�T��e�R%���L��b9@�� u,���9��u�yU��]f����]W�Ң����K,H�c`��p;�1g�=pm��p��E!E��cby]��<?�6��r_)\�<~B�����u�|1��D���˭�Ȓ�n�bw��q�B*���\?pZv�+��FSj!��֣7��F�-��B[9ܱ6S���j2��V^h�P��*�6���NЏ�/���̻�f��z^�� r
�7P�1��
hS�mf�c�{����$��W�^W�����Y<j���.�>Vl�0o�8]��:���cY�e�D�܉��ou;��1S���B,�T'�k�>��DU]���7�8��>�j|�������Vc�!��c�}r�p����(�L���ˀBVΗ�����w	/Hsu�Ћ���'��ax<�=m=�<�4en� ���l
$k Q*GDz`�(���=���$�U'��	RX	���R;�J�\ٶ�e�z�Lvq���
�r��X�v|t�����{�ޱYw}���dyt�/����ۼ�ڣ�:8��W-e{���)�O)��.��[���;���<��E,���]?������w����rH�������@��M��0,��N�,��Ni��Ĝ���1GBJ��ƪ9�5��K��x��f�o��5�Y��]����
g��?���\>��a�ɬ��}6W���:WeI��� ���I�*l�E�q�(J����C��X�5�72��`���2�ޜ���}����1�-�^�L���V*TӫΛ����\�$��Di�P"�����4ܠZ��c�͎�����;����s�^Z¹P�#����g{!p���i����&A)���;B[�t����"	�Sa�����wn�吖j��˾m"$��Ԗ�� yeT�  �s7(��:����d�*���ً6��ʼV�w���(
Z��ce{ko�q�m��Ӿ_ω~��$���U	Vz��&��!WAAV�; }���)�	g��q�K'+��TCB�}��8{`�6���ʏ�͕�6;����Q���M �Q����u�OAw�&�j�4*�۞uh�l:;v���H�U���zDW�������f�/L��\�a�=f ���kZ��3��P�f^˃f	����9i���[|���`D�#�B��۷�ZM�bۜ�d���R�]<��@j��7D�Vg�V볘��Oئ[��f��6� ����<�ȃc&�5T�Z��-�Q<2,�� I��S��#�&���E��r������c�;fE��������V������P�,w'��:#�*A�
��4
�S~p���@�%�Z~��������>X�1���0�ۿ�����x�&�c7�iHd�{[��t�w~���Q�N���ɍؙ'��n�AIÚ	�l�K]W��K�A��ţ�#��9ER���h�x�+v��2��3bE��dE�%MT�j~;�&��ONrf����i�tDe�O$����r�OG�Wa�+a.P�0M���p1>�)��)��}`�`%�L��K�1w7%���3Hes]�|c��@�"�{���˨r���!|�H<�4ߓ򴩋��D�"H�y5"Oyp֝���g��Ґ����}�AW�r�A�Ɂ�-�(�s����\�?h-���N�ˬV 揿A�NU�x(�;&i�[�����؜�c3<�n@�]��Y&���Z�CW����$*sd���̷5����E���!�- �L��t�xֻU�p��453��-w���7����7������$�-��D��	$�s��x�?wo|a�P9cH��!���0���.��	Ҽ4v)�s�G�� �F3�*����!bX�=k������a����ķ�T-OX�ݾ%X4���oqkܿC�V���?*��?���H^��	WHv��y.jU��8�g3j}d�֨n;`��!�1y�Q>�������������U���wt�p�2As�(J����'����X�5��j؜䠨�ϒE��f
��xmb����F��<�#��9pڏ��|�Fe��<3}=�(r%t�>y�j���+��BW�����~�S�5�e�.��tю���l0��ʝ�b�S��H�c[*��Um&������3�GZ1�kU|c���đ���n��@nnr[�����0�P��#'��p;��2gЮ�D��V�;�%�{+h$(�.C��M�B���Af���G��GQˮ3�|�M֘�Đ��[_�ȁַM[�Mf"c���g6��.�:���0J��:�릔����M�e�K,d�t��Bi�;��V�DVA"��`XW��7v5q�}���$��L76�=�4 ��� Y���u���r�a�d7i%Q>>W���=�֪зd��d�H�爁�}��lt��즽.���s[�TGhx{>��!�cA����l�h�l8�Ϛ��dc�4�����!�X�2[�;��u>so�J �6<�F�X�l�K�|V� ���%	�\�;0-�SV��6Qe�P�Vk#/���s2'&�V��Ķ/�e�VGP%H[EpY�:�AK�V�9������/����Q*������4�-���)����������g�N��V�s�� ��X@%>�б�>ךbG��N��x���@�2u�(��Z��e� �y	#��ݑ
��z)q[��ո����+�>����v[�a�iy��<T??A�-��Y.������43�JT
ّy�����B�p�ZI������ƹ�z^�~�t~>#���MJ?��p@>�><nf��mEb|�`hrs�(��X�Hq+�,Bs���S�h�S0�A��1�6���v�s+�I�|�_�_.��M��Gd��{j�y��6Ȥ ���S��L���}�<;�r�B�oᥘ�mH<e�z�|��=긍�����'.G��a��9��di]c��e��\-�Mga~�g�܂?���ӌQ���6�%��(��-��Cd�l�b�Vbڙ��'Z��&��)ia%O
�lY7��Z����H�9B�wh�&�@�8���&�Rvm$&Z%�P>߬z3cE�#]�m8����ZtSy�R���x]Q�L�O�K�̻�V�������ɏ `�#����PqG+�}���.�`�'���wy���"Ba�7x
ښ�E�P�j�w+iӛ���X��_6}��a�9���[�5��#�w���W��@FڋB�@i��OHL<�-�R���vX���b�2�ȾNڝЯakm12�ٵ]��;���7�5�h��dX�s.߷�C��$r�A�+���ID�4��6�{��*�������ڐ���.E���9���QJ�z���C)t6��,�e����.�#7�81��Y��+g4�l9��.J^粺�#�7�k}?����C�w��8#��o�g�2K�:��!7�H��f!֟cPNZn�췪g46k�43��<�R�!�`����PI$�ۤ���jf8���P�8��&�U�h���lMBc~䎜��GkӖv?��/P���7T��:���e^b��Ե&CN�n.t��d!hHޞ����v������I��K��Z
��Xr�v�Wn��h"���K�L���7�|2�#]��:Ʃe�>�#�ԲY֮ۊ���ȃb7�UgL��Q��g�)�d"eN�#�Q6��C����%��ao��F���˒�]�m���7c��X&TG�K���yG���ڂ�a�A��f>��T����K�>���-���A����@��-�+���$�ө�KI<i�%YѺ���Jrky�A/[�B���	����cl�]>��~LG�%e��Tc�Fd���\Ѭ��G�ü�E,�K��lꔿ��]�;]]g7,��4l���[��8�l�$1ok�lʢ���^�D|8�z���H(�M��f��@��h�i�"6h��[|3f�v\��jn�=�[���?
p|�_�Q�|�]�Mir}У����� ���| RE*ݐ>����������5�X�L��ף�����~;���8ZK[��2����������H8��HN��HۆW��%�;��� غ#�� #���l��c���g4�ٲd%�[B�+����v���8R`7�<�V��&]�ȋ���ޚ��+�}g5�#��CF����w�HU�IM�.�u�o��2�t��y�jm���_g�ʼ�Hw	�C�;6�.�[�[ڲ�(wȡ!��8�d���N�0��a�by�e\���yM*f�����kH`sL]�U�k�C�7��L	��O�)8qt���t��i��������2�jѹ���Zi������9-1���@�;J�b��n�����tI�L"�
v����ژ�H�X*Z� /����G{i�
7�h	5=�z������j̱۽,��ܠ�%~'��$Y�N2©��,r=ϲ��R;�4m&&��5^��#��m�ȧ!@.�����Qa˃ ��
��^����K�"e���Π>���M�,On�v���<��[Mw{v+�'`܄p��(�
���k�`ᙤ�hQtA�j'МS�!��˄�%%�xX��K;�ࢄ�D�xZ�F�	�,z)B�
ߖڿ�v�ֱ�k~�E�DQ]LClԒxf�嗀'���e�����R�qj�`��&o4H�ǯ+?) HIQ���v��
�?Ҝ ���`U-<����϶��s�4Qir��'>�䃂sZ�n���Z�/�C���iL��
��:6���j�W��c]�(~�J�m;�e�&?�*��@���r�h��hK�K7|��I��@�ږ�� E�)����L0)b���S�K���ci�X�%#��@B��v^��݁�6>�5	����^�\�l���s�@�u��7�+�V��%�z���u��&.d<���ʫڎ3��#��)���ho*�q��ĩ��Rz/��2��l ��56�VB�[P����韇[eT��f�82���
��h��ؤ�A�������a$	�����*��e�� ��wS���N7����֢� ).E���K��Ɲz}(�hS.���0&�n��_���)N-����Z1_���9O_�����]3T�^���	�n@���f����м �W��y3ygz��q���T�k{�ǭW&v�8�Y��LhWY�0����4|���e(9��7Dx�mMv� e�LUL��8�lZŨ\�K�K3��&T	�)��Y��n$(\�|!Y�5��Gl^�5����ƽ�{;S �'״R~iY;c���q"���`\)7[z+�0�R��#�;T�{0 �-���2JVgz	Y���Z�$�ι#)�70Hy��k��˖�,|��G�ۘR�����L�I��Mz=�8�5s�t�DC�Nɍ<2�A~��X���*����:���Xt���1�u؛�K6�Rp�5�%��c��$B���`���շܩ��E�k���A��mW��^e��zr���o��DX�_������P}�n4sN�2����j,Y�9_M���:�aߥ�	�g"����PC>�h[�E��]B�|6C�[��UDF!5�_b������0&����.��� �ģ��/�2C7�wm���%�l	$	����f3��sC�+��.��&]�I�Fχ{��  ��8�X��yo�dH������9TH�n-S�تT���f�YP��H~��U�&��r�!B f1�x�1�0��^T�p�nܦW�~~�s���~Zr�ף]�,�iuI#r�#�f��ց|T�qNg����q��R����A���<�,�T���GN�A)F�O/���;�(�^a�!!���l�u����P��
:���_T��ra:4�6�����l���fh�g9m� h��=��Q��
���:���.3���Y}�vTKa�%�v;@�%~�t| �v'�l�l^�f�C�1���u)tm�b��I��ֶ(Q�D��QS�Y�4����aF���[�T�W��x�i��4�k�n[��_�S��W�"��mӈ�zz��1�'kǑ��L���s&��Ap/(�eA���e��(ǯ�ͫ^��N��ۘTz�"��Um�=�O��3ܔ�e�fF�WwG>���JS)���o��4��ѽ:�/I>דP��F�}u�;6
6�L���ͲW4�/g/�i�Z��2I�U��~�	���+qD���ζ hl.�̸ʍ�Y<�-�;=�����@g�faZ�˿��(k3
(��R�m��"~*^Z!ѯN
���0���p���q��5�$�<�>��]��V�Vo�U�mH�ƌ+�k9!��M�y�Y��K����8&�Yߦ)�;0����4ˍ?�ڈ���^���U��kTP��Z!;���-�;W����\��Ӈ���8��V`�1�)v�m@yX�� @�x�a�,�1�%]���𪡏���G�乡U�#I+����y	�%ǜJQ�ԫrG.}6NP䔡�[�9[�(<(��ME�miK��iJh�s6<��3¸#n%���kQ�*]���EQQE�#2����A��y��'��HG�K�=߽3K��#��G�eo�Z^�v�偊�)��L�5�7�UF�/
��������3� S�j�^�i M�����
�����8���^ŢU�d�6J�^n>w��!?��=j���ȶ�=NU*5����;��~�ݎzς�m�a�;�iȾ)F2�`�
w��'��Ӑ�k���,��\ ��<JYŶɏ?��>Y5!A�r��xq���F����x��X����x�6��6�#.'�%�%��ȭ��U�uWwL�M�)s)�+$:�����	�D^�����e��b�L�C]ߚ62��@j\J�^Ʋ{<���Z�Yԧ�tc����n��#���/tT��9;��q�BMz��Z0�\)��ɲ@�-/�b�1�� �5�HN�ܿ���������P�<6��)�ͣ�Jn���UP�l�n������8���oةr�=Ka�Ua��H���ʎ$;g�����Q�x��!dG�G{��|������#Un>7���-/�[��������۔Q�N�������k��W�c�F>��N��?v����h������t �9-Mt���v~�2�N<)<�����.uH��!��\h�<��Ժ-�{]�.�x���B<+]��+��o��)A�������¨w�4s�w����BJ+J|����7�Pޛ�'�}.r+R||v4%� h	MPnp�9ʶ@)@���Ϥ�H]�H�N�m��9��MP?�}�f��[��i���?�#��hצ�˪5���L��[�rK_B��CrnZ[�*��P�.e�!��Z[o�z�B�O�/��\6��(�y<����#K)Kq�������H��X���ǵ��hl�a
���54�z���<w�s�����(�Ȝ�3%�X_��ў�V�5O��qpr�����T"!t��#�Yݗ��'|GA�
�o�+ 潶/)G =�G�W�G�vSӎi����#f�
��J��s4�()b��`��5�w(��?ݧ�|b� .ȅ۝S�P��_����31лɂ��V��|G��3"�td��,U��>.�["|��Imz`�d(�V�������� �Ȏ2�5�5CK߃���c8d�w!&P �쭑�����\#6!y{�����c�`[$�L�`_`���y��"��>�'�\�g��sp'��O$�a��6����L0�vZ����pl]�	"D/A��bd���]K�&��bm�T�˯2|z,��p���Y<����4Xb/W��˅����Kl�).�]NT&�� ɪ��ϥ�̴��}Ҷ���ՠd�Ԑ�=��	e��4�h���ȷ�	a=��rj���p��f�P�.*�!zOHS��gJsZBjY�����ǞZ���5��0�w�� ۡH>�~�+q�_/3���qz��/��>Ć�<!Mrë1Ke1!j/p�؀�D���a��,5S�R�Y�?��AD�hò� ��j|���5�i�zI;�R[��9R���OQ�$�Kc� � �*H�i��4�y ���`q%��o�g�]�!4��GHH{h��ms�c9]��?�F��jsK��?��u��/�ӝ������`��M����QP����@�)�m�e�!t{��u���ѿ��M���ih�я�n����K��,�bŷt�!��Qef�e�4���ų-I��]����v� �⨆��v��W��ׇ�͡�R��r�.O��Y�J)�JQ^����f4��s��`������Y����E��t�����n�cPy�Q�j�����HfL=��{1�o��eQ[��J�:z���Iu��}ﲍ}�%>!G����x�Mg�^a�8���b�/�V��㮁����+t{X\Ӱ+��^3�_�VӺ�o�����-xB	����!���Բȃ��yFGM��IHw!��L�KwX�hɉ.�	p����X�>�}t�5L�T!���{"``��Nf�}f�c�����A�O���J�DyJ�I��P�m����%�Iru��o�.i��˗tԖ�I�D2F���@#���V�G���Z����/	����80A]���$�'p��sS%��4Q.��[O���E���es�N�������*m�TNr���������HI��������µ��\�񛮧R�
+�M3h3�nY�Q��2�iO�����i�;�{�ˢ�B��e��Yc��:#�$�م��vOɅU����7/��,cR _	����3T��25N�ߣ�~��x{���nZ��$�)#�.\!�y�uWTxvS��2L�P�[;NSb�#��B\��)P� ��g]������_�I5q���1D��3c�:�\,�N��N�ZL�al��(���ך}`7��fOX�Ŷɘ:����dw�BY�Z�6��b�*@v�O�xJ�c���ª�X���4FH�l��@���<$+s���ਲ਼�|Z��z�/;)$��9��te-#�=�V<�W�顙�d1��T�:|g4N�r�%��3��#�K�.��z����=�
e���\`�p��FU��+��U��n�X�1��5��MVG��Z�6X]Ե/Й��cB�Ԗ�8���F_h��_�4e�l��c	���d�H@�����`@:�����{��P��p)J��s���O0��Ȥ�D��a$1.�FV]R�A֜��R|m�O��NTT�n��F�%Ǆh�2�A��5����/;�s�@&<�6�h��0��S�;l�^6���Z��$ �9�>v��9�!t�����Q�_[ �7�\��x屗�e$Y����f��3�G���짣Z@+��)���M��)_�o;i%\�~i�iR�t��k��bҪ<�íQ�0)�54���MY��7-p�zKC���Zׄ�s��e��Ѵ�bA�[M��
g�{�!���䈍9�XE���`#�E�I� /|��������nl�j������=��`1u���~��󛉬"����*m>�b�g��`���ޘ�J��,ͥΘ2��ê=%I�Ҕ��i�rΰxi�Ԁ
�:�m�������%.z.�r�»m.	5͈�ܞ,�A�/��Lv�H��J�
�9�=�6�kˀ
����\S��"�V�=5V}m�^��N1� �Ԑ�d��F=��\��#�h�5�C������ZXT"��d�U���^�
��97C�L$�9�z��3����n�o���ÎnI�YT�*^6whA
Y�H��,Lu<�lZ�C`u%A�qo���â�Y�^���R�$����b�&�nmh2����ݟ7�~-��[��C�i��[�7<>�>�I��l�BwE/��66=,z2�E0����^�䟍�
�YPk�28=���[6ak��f�ب-J�2h�X��to\ ��ˆ���N������*7���;��10/���p$�$�<�7�1'��*}U:��W��y�e��O�Tq2	5��8�GY3�.��x�D.���܈	���uѫP��D�������'��>͒��}�&�6�?h.��fN#����Ջ���,(�$#s\�I��6���9�Կ��RUq��ؼ~�*��!���v���Eu��?;�0X�O'���]Hn�҅(���V,ft]���"��Z�s<�-����JS��b�Ǯ�1�c"B-�+�I�lf'b�Nw��n��U������a�(�w�N��Ҭ����S�yY-/�A@�IX�� t��̓��Uۛ��?4���޳nQ?Z�pr>Z~+5j��*��6��|�d_$d�Ɔ$���G�HC�H7�Pis�#&�C���� ⭈��b��ȑ��)�Q;���/뮬��&�q���0HZT�E,^C9\���r�Y~��>sJ�kX@�	P�O�)�̀:z��
7"q�jK^PB�wP ����KХ�̍�XՓUT�I��I'�WeR�M 'q��W�
����;m�n�9�9�P~�p}��xG ����*�Luw�<V��Ȏ<��t���|�)��B6���9���/F�:3P���2Vw�`��~�/f��t�_o��yc(������3s��>�|t�EDw��iU�������Е��2����iy���n���"�v��$� �K.	.�X7oͲ3�����f
T��ғ�G�j�U.�eOs7�iX���EUSR)_�R;�Һi�8��O'J˛�cRGQ9`��eG%ᷘE%\N�.(���l��� �8�,MQ5�����&�`ʈ�6�Đ��򶝇�x���X�'�͑ӎ�g�)��0k��p|$����N��R��V�K�~��vC������(�@�m��=JNYu���L�Ͱ�U�w�Z�`�Y:��V�/�Q2��5u��(�m|����]ȁ/�Q���/��J�zj2�"��b����j�N��'p�S�W��-�*>��������bg����D�m8��"��I�y567` d�Gj�eRNb!l:�Ģh��\>�h�UCG��HL#YMF���C�%�O��n�
vBpi"���s`w��B6�
�/Eqo_tbXM�H��?�2m7Iq$��������� ��p�A������6��+�̢,LA�ܪ�ǮCm���i��V+�O�����,P+x,��a4s�A����W7JC ��������mj�ld�Z�<%�l�';Ƹ��}�'m�9	��;��ܙʾ��������I����h*PJ:��|�u4Xm��\�ut��[>$x=�0)��@���*�B�(��s��A�G)���[�T�f�%�"�һ9���%+8/�)��*H\�>��-�rX�MF{�� �q�\���_��W��a������a�,y����,:?�=̤��=��OlL�~�$ODW�����Ĩ^�˷����Y��m�s=�rɹ��D&|*@�CZ������?��m�@�K�C�c��(�d{�ʺFi��eI�"�`� �뼯;��G�����#���ۤ�9�C��v�n.�k��c����wF�@� +��Y�j
�^�ґ����_M�����%�{+�Sy�µ$���մ_,6[aU�bWU/F��fe�F��3�7_�^(�	�,�Z�0A���)I��ۧhX�u��dU�ͅĿ�z�����7��(���B'Q1�}9���u���b|֬m2�ޡ-b��â�&o;���f��\ ��z<7�2�����Ӯ2�$��ی}mO�q"�!n�G��)C�Oyy���P�H��n��V���b.��k��WEs׺Pg�1��e�����)�yKE��ER�j��~�P�s���ª������Br�G�5ELP�%����vƭ'���~kc�f���]T4�5q�D�Z�r>�vTw��	*1�b�*���հ� ��{��H�"S�sH��*��0ʩt�1ӓBUl�{�̒D�*�'Wk�)7���)�B��)��ŭ���W;m� ��S�^?��28��[�8DSm�b=�,�Q����4�b� ��h��٭S3٤��ɠt�^�h�
�� �y\<������^u�Q��R}�b^�z�O;�O�g��.��\��S�n�.�k�#�&����9x����np��̎��&�»��mm�/��t"G)䇷_{��P��		�<?���� p7aM�%�;'����D��R�AK�Tk�ٱ1\1�,�[���4���0�p$0�4�NA��;l�u���H��ؿ��������*X|�֚��Ԫj/0Ȩ�����3�瑫v���������q���+�R���r��,��h��t�0�]�j�!`Yg*��9�0�mϺ�XF���ᏻ�q�!��8�@�w��4�ZC��������#�r�@�/��a^cZ�!�Ae'������j�/��'p5vWOJ���Q;��͚���-���Ք�+x*0�eŪxU�%<ě�?��$Huv(���ofG��o�;��/�Ul+�Nx��[rA����󗌑az�6��1L���ɾ~�?��ց<8=�,%I�e@�zj�F�tn�q~��Ц% �8�m�e=�K������ns��Oy��/�g��f��K�g~�/�2�9.iTIWI逻v��*�A�0�Ihyȍ$m �?K��*N>qq��M�P��y7th@|�2�������
7�����VV�O�����#4�m]I8D��=�����m��JI���
� �u���7�����^�� �T���蝦�y�eР���H�y��n��]%i��0kP+ �L�u� �xtH��H�,[�ftW&fKf]��&�`Yg�����X����3�r��5#xc��(��l�O��r����.�3[���y��C��hy��>�h��+�Ԟi�9�z�7�z��j��«?��:�}�~�ŒӞ�+��z�|k�]�i.�L����.5� eқ�1Qסd@Ⲅ�δG��NlKkG1�=���A�݋ђ��i�|�����,ߒE� ���H�����+�6:mH���������O;氣{�75W��IN������FN>�$�x�p4S��G��N�ͦ*6��x�֫�j�=�i���v���W��G�/�����s�Vn��(���X(4�[.��L�@���E��2�tá�=�:j��߽U��g�C#	D�U�SW :�w&L3d����0�1�S��@�s�(�nw�C�W���Č��W�v���Ś��'kh�_�׆���1���I�G�c
 6o��{0�+AXu�4�D��;c�K�B��jr�r���*�V�VX�pM{d�ؼ`[3��������f�R^�2�^�	�o
��4�i���:��ØW�_ۉх^����!�,���N$��Z�F���>�~
���O)�jw#M����X��s�i=ڢGi߽���#�p�X!�)�����V0+p���*I���^ƀ��8����l�6�����^*[
�ф��BB�� �C؟��/n!�2�y�\��Ë���]ܔ�и���Kp��ꙅ���(2�H�2���	%0��y��/-[����щ�-�4���w��&�y�����k��;�U��3g�����<�������|�N(����ޠȏ���|Mv#DZ�p���$�wzZ2�pPɵ����:�5��1;�I�pj"
\�v�<�����2�^�#X����$͍ �����H������Wb�=�06�tM���#�-�,;ɣ��}b�::�_���ҧ}%\qz}�VD�������uJq���Cl���9�'`�����Dk��=�V�s��oɫ�rt�31+�u|Cq�F�\�@!-�hG�	h=��C� ؅&g؇�DjV6��`d�g�w�t腎�QZ��;C?�0����䳋"�{��GQr^����Nn�vW��lx*��R���Rd� Q�q��{1PPnbp�f�#�B^T0���T��Պ��^e�G(I��0�I�+N6xr�O��;�FQ��ȴ;UY2RY�6;z���:���j*����d������		$iu֌�ݠX�Id>Qp:{�����[z @7�����s�� �+0|�������
Y�3��o��W2iU��	�iۂ��ND�����G��z�B��(;�8v%�(6l6QӫLG{.���%E{�]����k��l��KQ����$.Z��ll����-�I5����+5�'�<�ڰ��׊UqIOHQAޭ�-��&��(O�.?YU���ʵ���N�@J�?v�BTAڥX�Q�K�� �4S��c#�;��;�F�>ٯ/k➣�d��>t)]� �������Z}���2�̿�qa3T�nB~�%�=# L�wr�n��toM��|l�����̫Y����fݗP���6Q�-(�#���9,�_���Ď���-T��x~���XS������Bt��=�� y�O���T���.f: �}H2�b�b %��-j�&3��.MeU�ѽ/"�gx
�* Դq6}½:��;���R���pr�� O���VQ��L���Op���k<�3�+c��;tڵ�t��g�~�`6�nMna�,� �G�C.�b��-m#);�2˔Ҏ��S��L�>k�G'��۪GP�I*�l.+�-Q��d� R%B�I9��r�;�*�C��h�����f��w���(�@���/�el�O���5���ob�e
��G>�J�1����` ��،�q=��A��9��!���,���y�NUlW��V��X������pn�~`�i�yFya
�-�?��J�EnO�������WIȎ��$D��A%(�&�{Q< 9��O�;�L�W٢�1h��^������7��\9}�1�3C���ęG�)�p�օlAj3��r��� ����n�5X<�v��ܛ;�C��Tzˉ�!-g�Đ�8?��d�Bw�%�u~�h�����5UEMG�:�o�&?J�m�{�,�fw�箸Ҵ��3f����C5����4�8�*��%���<kC�i*��;R��!�8U�Ad��k���̲��R���t��ެ�$�m?�I>>ُ�Қ!�q�zJ�#g�:q ��k+�a�+�(���Yt7� z���(���o�z7�5;�u��i3��F��;�=3��?�.���U[)�E�un��M!gm�������>I%l��͘M�ٔ(޳ˑS�EG{3�*�c)���Ͻ��nD�'�X���F�J V��8���z�B�u��ʖqCP�� '����2��
G%�#�����8�
�*�C��U0l�{'\d�DܴƩ�yZmxN�ˍQ�-�LF[q�n4�L6�3�K���A�x�̧�f$3sN�Ƒ��-�؁�p�C/�QX�E[vSSD�u��O�&!�GWoӓׅ��	dcPC)�SF?u=S��'N��(<8s�g���c�%�o�y�R�'r#��93�/&ʐB+��~w�;��6���ץ�Uʫ�ܢ�8���6Q҄�JB�8f��1Ĝ\��N�Dm��? r�S�gi�Z�w#6�-&T�q
�:݈�#�'j l8"�-* k)iU���H���ha�J�=�aR����Xxy��L�\ZAr�5y��Q���*�*B��X풆�f)��8�.�Ϸ*�?�mɈY�B�͒��1x�=���4��$��i�i�а���Ҁ�y�U�rȦ!�Z`����m�B�����6���<��A#�k��ќ-��V��O/��!�����U�9��b������]�ZN���#$���9�D8C@�u�~��S��m1͔�d��|j�q��u̪W\�p��7~`�G��,��hWK��lQ(��Ȼ����/ϓeɘ;�{�'��Ct�z�9y�$f���0*��87��T{�������KQ�BYю7�ez��sTB��gb����H�ezSaCR�_iRAp�aId��\W���l �@
{�R� 2/�t$EL��ti�Ά_�*#x�UF,������(wU(ۺ�$|T4r���L�/ai��:�}�c34,��au�Զ�7��U�_H��LG��& �B ��m�>	��킘���,�����&�
�)��������N]�[�{[�P-�F7���lu��( >�i�˶Ck��IO��2y["T}j����$]�D�D|o�i�pg��1�,&a�=7�����!= ��v|�t�_�[����(�1h�{a�d�7��|�թ���H�����K��7.��e�M��,��kQwY�g[a��[(<r�Xm"��BDI	C5ݒ�{�z��?Ʈ6AI,ɇԒ��9,���1���]"���n�:wO>��b���/^e|�d(`�2�nԮ�yJ�pe�r��;a�� |N�u
���W���s��u���C���<���%�!�!��u�=�lb��)|��ֱ�Ϗdg�C1M��..�֐s%�L����v���ao�^���#`3"��^��;.Ens��Riӑ���hm'��w޲�;ek!F�+�K@�Jy�����,bƏva�͘j��d����1CM�������5C�R��l�K0]��`g��&�S����i�&�W`]�:�S���e���bl��5�c!���m��(��Y(� ��@?��NzvQ�?W4\�l�;�A)��j�Ȼ�8����V���o���E�;p���;����Qz������y�}Of���<�fæ��ה��	�_q���HG�d��Q��5���LL~�����½������f�䶫BQ�$A㩙'$8C�J�U�U���!u��I�l�-.�%�h{���7V�ƽ��m���%7����6{��M��%^�ފ��t lW�b���Cʔ��闒~:#��L)�S�%�b���6B�͈A��-0]�@�P�\�f}n��a(�9���3h���r�L~Q�K;�f��u��/�{��Qr�]Bϯ}�;e|�bo�_Wڏ��De����s'j��#����=;��p&���% ��C�~��n
7���@����Mr�SE�K�.ws�4��Ҝ4MTdt��q&�/�碒,�s�9���6�-�wc3�=�;^K�O�_����,�.�Lj��M/چ<�ߠ'�6poc���(^�\���_׳:���(P�I��O��ck� ��_뀍��KWT;�hO̧�H���
� gў;�m�\�|�,2P�T$((T�;�[�pG����G�z�B���3#}L����P��C��oq��~a|��s�H��q�6�%~�$�\�{m�c=
P|�K����}H��T�@#�s����5�,k>�5:G
���M����b����u���N_����Ί$��嘑���b�e�q�������e$!1]SՖ:���!\Xk|�E�#���IFu&�j�?2(�6�H��0Z��
S�|n�V*��7H�מ_����4-�<�m��-uVȮَ�W�J<�I�.��Ӧ�ʁ������N{��ݽc랔I�,:�V(0./M#ؿ:��ח0Xt�:R�j�_[ɩί��[�?�B�4l�A�-�䩬	%8��9����g������Q0Õ`�)^�![��u�v���/:f�����XVh�FQ�i�75���F�0 J�Ҙ5 �B`�J�H�k���MA�=���z-@#*�'�rV��/m!��w�Vۺq�	��@"�d. �ѺĞ���{w,>͖�1�T�`/0��(�c�f2��}��W������v܅-��=�6��8U��+���/]��d�:ï�m���[͸O�|��g�LF��"�/�q�@L���2`�Ms�o5/V�꼡��ʩ߷�f��8iyYB��9AdN�U�W�t�����믝!��,���֕l����ɩ�=j�l e��Ӣ��d&6�B�:��*����tۨasOn������K�'��Z6YkƟe�bah�u�����G�#���jF6DVR�l]
�����\l����`��THV9���l�[�ѸoH�ב\}��9&'#k�_�=a=~��7Ռթז�΄��ȼ��2��p8u�$P^��녾 K4��o�a%�P0�e���w�Q�H���^i?C��T@u1X��GIl�����4�(ICҚ���4�X����:�<�ז>�����-
����g��dMa�$2:��.��΁�WC<��j��7=bGh�'�A��K �Jp�zN��@yI���!�9\U�@����L��N� ���H?/�,u/�HC��fl`s�H##����X8�yA20�em1�-��HN�\�Sҏ����=�<x�Oet�}�����ݴ��Α�?A6��Yε�/0�E7��*;�y
|�c�7��<��V�}U��蒾L�'�g���C�V%�b'9' K�j��B�2���-~�(���t��o[��6��_o�im
5�2㲷h�jm5n�gc�����tl�S9m(���?ytY�
�pQ	���r����|$Q�*�(����DG�J�AgA����� 3l`#čr�AF8�D1���c�"�h�4e���pt�AO��C�J�fB�H����Qe��߫Z����K���o��{ڋ�{��๨��t����7x w��J8r*/UXa��!����[y�Dy�8⽚
D��s����J�[,�4��ݱ�y"�74=v�Ŗ�ފ�l��A��uG6���[}�]e5�2�'�R�VH{��"�Rv����^��մ��~9C�^�2�e
K4���{��`�����i��)��XO""��X�u�h�s2���Ҝ�RE�%N檮��" �}���䃾�Q�'�ٰ��dV�uI��D��� |�u����mĜ)D�>�
(�������*<Q>Ak5�,�(�`gyWK�}Z�l��hꃚf_�}����{uK]�v>��:��PWk�;�i��y6벇��'Hz����fz���
��Ju�o���LN�h�y
�Âl�mM:��/.-bu?)�&�YH�����T�)�`���V����z$�3XƴVV�ի�)�!�Io<�!+r� j�>�����.��SтԲ\#��9��;
#�i�y�?��mG�6�j�-�6(S����^:��D�5`q������a2|R��X+�봯`�J]!'tR�ͤ�~�E'S&�QY_�Rf����] �O�e��h#C�>� E�z�L�'rwޜO�(�u}��c $6�(��,�_����L6�!�?p>.O���5�<�.�X,�6L}U�k_���Z	w��f��P����DiϨ�c�Ĉ�ǖI[��s�*�Q=�ĥ�?A� wE՗3oV��2��U�⊍'=�(�U��� nl���[�T���{�
����GG���S�j�発t
��M+��������*X� @�K@73�Z��u�|���vu-�o-�u��X7�ba��.�C���&�}7Ƭ�w�Ѧ NQ���}�Z:����R�0�y���KЅ飂CU��?��)�9�ʗZ �����r��U���uW�x(��O�L���yۘ&bx�e	���I-���MWgL�
����n��V��0�B�8��h�ww�$�(kmjd�������ޮ$��|�҇?F!?;�!�G˵��^b�h�7'�OE�_Y�0�:�����to��CC�k��۩e��@�gԵ]�K1�������C�0���4Oo1��ٗшș�I����_��r���N9��Q�
��+:��;�F��sd �����Y,f'�~�Q�_��tL*�Co�\);?�D]לO� �Gk��AT3�'u�_vE��/��򢠜���rUK�-���/��hP��+�ǰ�*@���m���p?6!��dW��O�����"��� B�� A�$S�E�H�-n4�b�}�QױJ����⣮���w�2�]�j���{T2�(w����'�cr�v�hk�%�*\U���óށ�*� [�*ѓ��c���0�����YP`�{�:��p��4��`R�����$��
Ý�_5Wn����h=�J��!%��E�j�gI}vK��>G*�ٵ0�j�>t�go-�8&#�}O$��qG��4H�D���k���gN����3?5��_Г�ZEB��W�DU�X���֫عs�ө���2, �m�}jȼ0�)ͭ�F�Ӽ�}�Mƺ���CD�[�x��(����}
CZw��=�3rF�V��Y+=s���]�C"�hm�h��QQ"�j���,���3[ 0_u7�Tȳ��D_�ɪZ?�z���~���;�_�#��	�,����Y)�H4vuy(�Ҋ��F�|Ta� �C�4�g�z�<"<G�I�n�yhQlt��P��/$v��é�/��{*�wM7�*�V1����/vJFj�����"3bИɤG��}Ţ]��	�%��G)�(�G�9�����W%�F�kX�i�S2��OD��P?���5�gB�}��SӉ��J��d�
��W�J��
p�9��f����˸��89D�Y��q�HM���$l!�k/r�_���GF�l>��+����j`2X�,�i�q����$P��UO�m�so�x�R�٦�Rj\3�3RlAg�����
�J�SF�K^Ifsu�Ikc�XO�-��Bq ]�{��)N�.N�#j���[M�sM������Y�C�Zj ��6�g���ޥ�Ny2WT*�oa���Sǈ CsRN��j���I��{�FR�����m(����\���"õ�5�s|���Q	����Z�s����	[靍���?SM���9�ɼ�����^�����Y\k�D��t��Kx=��%)�`���՞� b�����^�A�x��R����8���.��13BW�tYm<-����Npk�����*ڴ�^A�G�ޒ�5��Kwa��"tj��N\j�&��T�g�XG����5�?!�\!�������6���)t2x�
2-������	�;1}c���V\��S��#�$�N��l�!���Cb�nA�t��*E�7G��B���o?Hh�;�tV�!���BSVf<��Q���Z��O�O�Њ<�����?�� A��K[������#�%�^�[�l���w "�� �&�k!��ȁ/������<Ș6�r�g����)��$�B�v�%Pd��mљG������G
��g�X��o�v!��㚠��T�V�����3�4ѽq�Q�`�����;_��N��M�
َ?��4Tc�,3��w�}ۻ����<T)���><��d�PW4f��+4�(L���B��\���ǎӈ��˻	�e��z��;,<��9Yjq�������W�J6*�<N5�����*S6`M�`�7%�U�MI��w5�P��K6/Ps$0wI)%Ȕ�Hju<����&�.�h�aK��,,Z�e;N�+�Ț�.�Nϖ� ��,i��j��b)Q,�	�C�d�����������v
��_5�C��S����"#��/��o��j_M��|��D�֒��̙|�n0��̈́�����jLq�4&��X��qB3��јm�TLR�z��׹N�b�2���-���n��K�lo��������D>���dK���P���cU"4\���GV�n���h�����Pe�%�g�-O˘,p�C0Z��y����D�l������o����<=2��6w��r�;9;�L��	A��F U���[s�)�Dm0���ItX�?�cW��Lu^�(���W:�:S8'f�%� (a�Yl�
Yɡ��p�aa�2�����Wu�kGô<�7�0���&+�ĩ1�%�/M�V�^�ӯ8'�$���"X��$�t��'<���?	j����$vL�8wǅ�?����2��)�M�[�P.	�fc���,����E����ܾ
�}J���*�{��0LW�ϡU�����w�sb&L@@�Y���5E_��$ӮP½,F���(��&�*�L�W�fB�'��o�1�/�hw��/ڌ���3��|B��~:�}�Z%���	��v�Zzԕ9�]��W�A�����ty-$b1 �?���Ǘ�-<���*-Sr=B~��*�h�!%:��IY{�r`v��؂l�69b-���;�+�Ơ;x�a�C.�� �3�[����/p���"��K%IQ������`����"{������
���.�t?�@�ǫb���G�b����O�}��=1W�=l�z��*2th����p���X��!��R��8�g�_=n�ub(�M���ƿ}$��Ψ�z�jR%|R����
	՚"���^V ]�}W��%�jz�N�_��������G��=�J}�p���I�V��m��Ue���t/��y6qa�7'<>��IY<�l[.�4�Qu�?��Ŷ<�}էw�%ס��R	׺&�&G%kk����b�j�>�_P�d,��.5lI�8M�;�Jq��� ���|-��7�Hv��9,����qS��ErS`߈�k����қ���<����[�BIA�gR�<��Ik2�^����	�6/��>]��.w�纥�i'����5��0$b3 
Aѳi�%�$ek7����NrdCd�����!�s����4<����Ja�a6C��p��A�֐���Y ���ۅ�Twm�d�EX$�|�x�;��m��8�� 2T[r���<a)PmP ��0�řE���$����(���ђ��0�lҍdf㴊xv��f�~=G��d���2��I�K�מ�	�;"+�'���B�pjb�8�&�+t.�w`p'�v��|�O�+<
c����MCIU���rcA��'{��E1�\�ǽ�J?~���r�LdV�"�n$�����W�R�ұ��1��4����>��Ս�)��W�#ccI��`D,�Ng�`U!��>y�T.� ���ዲ<E�9�Oiv��^�!�'��P47{h"��a0��i�}��P�D���&��u�2kן֣�-#����a�����=qw\�4�%0���,WoW95�ܢ�b8r� إ̌�b�Uj`��Y�u$�����#������R��8%laB̃������։�+Q�8�ھ�l�������oIqfB};�"M�h�tUd���8 ��U�_vJ�X��^��G�l���nC�d�����
 4�>2�X*����W`^?0� V�������@�Y��.X�x�L�E^��p��jtoo ��VdX��%����l�����fy~G�z��G���ދ"�ܥ0�Zwm��ڪ�5��_;3i���8�M~&��aa>�mᅉ����fŭT�1JV{��s~�݌�j��D��<$� �Jy�O��f�8!�7�yhh�:�|\���Z��0Xk6�ʸ8O�
b�6�KO�\
�����КK�#����q�j(;Ӂd�"U�K��6�!K�P�z��c&$��Tg:ܑ��gh��*��l����F�)9X&Cx�Y���}�=�6�K�~�a�^�Y����^��ӞM�����ZrG#���A���۔/�Lj��ӨNV�C���"r�D}�~�<�8n�p67�07��=k'�?�w.�P�� �e_P��ܢT^�M'����+^M� ���,�Ş�)�2_:�g׹���L�+�^υ�b���F��pΉ'LF]P/e`��4�]�IT�y�L���@qi R|&3Ye�E���I�J�BE�1�y<���QLGsc�N��*̱�q��K*�'����eW�=�����(&P~i�dp�QRP}�Rx�� �L"�ӄ��m�z�[S^�5/)��b� D��e4����4f�Y���&�gln�B�>���՗�)�OKb��Av�(������vK"WP�1,P�Su1Y[6���w|Ī�nj��_��Z���q'�h�%+<iO{{��-�)��;���H�9Mwv�v�;_�1~2p�K��$9}R;|`�^@C���������pX�iyq��hS�Vb�^'<t7�J�*��p�}�y�uq�����t	�d�Y�9��"8�VV��W��^}Gň����"���)L-R[�n�ayI�)n"��Ć{!j�D�,r����V}�V�uSl���s�
��@����IUlr?Ms�����S����u_/ʎT���ͧ�S�E�1���Zl`��$D�en��⍫j\�0?��Z-`=;�Ns$����Z����I����,y>M���Uq�}��P��5���b:����tF�>	��&�L�N�R|�D�j�]�f��{��,�M~y�4LKѐ������y��d�@ty<JH��@#���?�HV[�O�g<���w"�Q�ې��|���QQGǲ�Jr1��Ҹv�@�I���w�����e�0u+�����v����	~Ӣf{��5�ۤ���6�~�%(�v��D����TA�<�D~6�z�ωC��ZX����ۗ,53�5r�D��/�F�n�tq2љn�`ݼ�bM�Cv�L�&?��=c���Pnf�I�Yy�Y_-$j�f�=�A�����f�&�ӷ)	�a���BD
Q|��ـ�QJu*�8:.Nt`����-\@'�({�ov�FΡ?���ܩ�� �D��	g#�l��ۛ
��,|4�l�7y�M	�d+�,�\8�y�ʵ�_(�f2~�' �=�ްg���"����	�� ;CdH�7�X2���=�`EV6WY
2*��l�g�X���Տ�0�g�̑&�����Qv<Z[�-�d���lv�P���L���Ag���^(�6�ڂ�Q4P�aWƚ?r��%��M�"ԏCOegL��p��Ȓ?�Y2��.N�>� m||�d�K���2���4S�*i�X�P�e��a�r�I��Y�%� X��qS�5թU��^��_K�ma8�3 Yn�to�����;�x~��X=,tly�b��Ҵ�)�Ȁ�m�!(q.���ֶ-=����r�Ǎ1��f�>��U?��1G���.���Qd9l.ѷ^	��o=��M��8�-�%a�}�yX�"�gź}԰D����W(S�g��D�̯�5�����W� �&�:XL�%��g�i�r��G0۽m=Sd����~D9�)B������:�<��0l��Z���7�rv4�AfWa�O�W^����tTF�ӵiN"0
�����~Z���e2�W*��8\`:&��A���i(���«�Ez������"Y� �g��o3xK��.(��Ʋ���U��Y��,��:�)�N'���b!�Gj"] ��e�[��yY�B��L���2N�p6�b���К´�rz��(Nin�?���sCt#��Ӭ�B�C�\0�P��#$D?�|�"��"ҢzԘ���
�P�[��.c�D`Vj���** �!y�#���+��|nt⯐�M���gXZ4�s��~�?^Q�*bu�\~uLD|יI�m �,�L	��gD!U45qޚ1���ڂq 0/;������ ��f�"6@��A�Ƚ�c]��*��U��ˤ�k�3��T!�8+4et���H=Aw=��ɸ�b���`�%��P�량��o�[�=�ot,����^l�!�K�~�A�>(�3��=�k�T�3TWq�]>��U��T��ϡi�N�0����T�~D�E�W���_����^IWj�3���] 7)36XERNl��`�x'gZb�ߥ2�zt���g�!����ZB�r���Ζ\)�!s	4�v���<����m�f�%��$7�մ���$�^q?��hM�cY�R���;O\���Q=8'��	��NI�p�S��8L�X�'��z�ͺČ��3�1Z%���#æ���i���x!$��9�*��$���$�M�񑫝��p%�{�[��OE��GݕR���Q�4v���~�2���fv�7[��y�فH-�Z`(��������ن��P��\߫)~���vu	�,��8+{v]2�<��Xо�mB��Q���ՇwL��4[	�]�E�m�ʇx!ɚ>Ly�y1w���m?�����
v�<+��~�:���_�'/˛��cz>��_iZl۵㟟t��Y����hʑ��nǧ�k�~�wjW�L��?rL�#���֠z��lE�������\P�fA�xIy{[��9?^uK�~������d���}́��U�z:�x�>[�~���2��7���_�-�q��b�5��?v�����i�JG�mq�ۄ��r�����Npgs��+a瘢�seG_{���?�l۟�9���2���]�Q<������n�Kx���1&� s��x��n*�G[7?��PJ@�(%Mj�7�_цG3KZ��/ah
7:���w\�:IĦF�7\:_���I�S��Tm��ڗd^S�����	?,i�&������<���$>��e���2�@K,I�62��#��Ϣ/�KL��U��˹w�,��y��ںd��j����<���"3GA	�
�Ǿ�>s�����@jjGB���P/Q�1��>Wv|Դ�D�*�L�n��ĉz[�	�@��E{�����8�������~W0&�U!ԦtF���q0�/�$�8o^d�?ς�W��we�PӰL;��'^}��y�뇀���-i�d�0m���̑J©����!\�S��_�S/�B��s�j��h��A�����-}F��Q���ZHG'oD�3��q[����߆�E�����l�!{?C��
i��v!�7��8�	)�v�k5r���c\�\R!�Z�0a����8S�A�����2}ܒ��e��񰇲�-i�Q�e@���Gt�n������X׬sגJ���T98z����9M��7}�2@-��i�|�$K�R]��M�y��b���?n�o���]�!T�Su8N(�u�OR\&��,�0d0��Ph��&H�^Ṋ�awlDRr�[0�_���=���V�؂�e�S����<ѫ�nf�y�g���KP�2/b�B��A6dL4�g��F�>)z�M
Ɉ����yE��茛7�V5�X�$b���ֲ�����>�gzBU�Kvq �4��T��՚d��d�U��Pqx2�ndxAq��e_!�#�����g!	0����Z�)�����\q��/��z�)!� �ú�T�bV%�cұ�J�1��0T�,|�WpZ�<+aZ���7�����f��v�n�˕� ��Oj+y���zI�|lc�����a6�_ �y���tF���ǿ~��P2�H�3�~+�s�Kp���X��-���
q���g�y�0�9���(	X�З�p=�c��U�8I�ڏT5*	����1m���!6<�aZ�O�2@l�� ��;�p��Q��7}�������s�5�r�@���yK�����
	�Eܖ�8�:������X�$�V86���]=� �Y������
5H.��Y��J=
EY�L].�	��G����������A���t����f�i$�`T罺 5ƴ |�Ssq�M���~L���.>��z�D��]�|�-p����җ���g݅w�}�ZB���qOA!΅��3���j��:����_o�����Q��o�o��Wf�&@c�`UƢ�m��uM�ʖFs՚WX��ĂԚ���:�]@����96��3�|���c��o���;�TZ�����A�bb�f��e��^e����#UH����z�d���1e�������K:�2&�˅���*��ʚW��s\���F���h?=g���ҙ��8�����O7Y����P����>�G�J����-���o��w/c�9FhŲ*�ď� �8\%�ɻ�����0�k=����p=��,���l<m"�(�A���{�{<��;[��){n������c�s�nD>�d��� @�J�;��@�ˁuN����@��*E#�*;z2r0��+��ґ)�Z/�2o�k���E<�����ovfX�b/�L�`..̥���1E��!F���W�TJ���pm]��!&�A7vl���=}x%��>��o�������)�Ke%]ΐ&J$p ����z�"��~Qt� �Ϋ�<I�5�SχNE�捤}L���?����������ƨ�X�������=��挜f���k����)9SAK�}�d�� ��Q���D�L|�ͣ�5��5�n�!�?̭G��;��on��W��c*�:J��<�L5�D�K�kC���7]�5���py_9;z�\�	Χ�^0�7�'٣64�ڑ�7����>�M
����ҩ�<�Z�s���'��I�tO��9m}5���ע�Ȱ��x��"}�?�8e���xAA���hsU~�8u�d]��(P> �pDH��]�ҡ>\;!�e���&8�;��F	ھf���P��o�B���`ď��<�W��~M|i�<�#���;�������$�y��}�� @�'�m�&Z����^`��s�}������y�ڕ<q�j�6�/�)I6MO�]*}}Hߓk�$ē&���(�;�;D~��.X?v\��cG�#��(�;��f�ɀ���*-��9;�Վ���qT���0��n���翺\���#�
��Rg��8��X�&��l���p�Ů�&G�K7���	�J�y�1Ǫ��h�:"�j�g5���ճ���jo(E��׎��'����^��K�����"òQ'U�t�B�h�y�
w#K%̦!#N9��eS���~c��8@,uR�Xp��]����f�ț�%�@*|��MO&�����<�d◌2�~�c�T�{�T!�C鮔]�v�p�@��m����a2º�0g,N��Z���on�o����a�d**���3[i��*2�����4ӿ��z���^`�7��<��� ����(a�7N����6ͭ�B֊����)W	Y�u�&	P�������e���=&���i�I��̭U��N�Eu�vtJ�`�b����!���b�'����I��i�xM?�Gj2��K����0à��'�	߮t8�sk=6x���= ��~8)1�~��ec����@���dH����� Uo�q�.�P��a�7)��y��t�yE�р�Dn:� e��i7����xj�$z�E�����B�#����G�����b��_.��"�;��.=/(��^"��-��M�	q{,��0H�@�pܙ�0Y	GHtv$���>����$�]ɩ���Ci[+��J�{8�;[?�-..%)��['N�H�����8N�����"����/����Zu�:�]��C�څ�	6�>EO{��/S�Z���r�~���̚��y*W��
ܱ_6�`�Vp�0���T�c-{��;�β��`�/s9��D�Y(� $�>��W�;A��ܦ�p�[H�H��:�����a6}�NE��*��y �����q�=7���ܦ���$\%Wl����������}��pmmy+��(�����7>�!�iʭSt�z������7N,jC-�X��V��"�?���C_��fɦM�m`�|�"{J]7I8Qg3V@=�$�M���Ϟ&T����3��[.�j	�r�b"y��|�������3�����}4��=*�`j�l���",���۶&F[9~1���9�Z�7���+��Z+d�_B��:k"�柢�r*-9����iE�t^2)����,�D��6Y|�4ھ�I�X�f(�[W GE�K�7K썩��a�c$��WؒƉ��@��i�܆��&ܲ�}�O�
<����A�Glij�T��yq薖!���|�L~݌��]��A��N=lִ*&�3��xl� 
�(�ˣ�N#l��a�>D��f�[C=T� kP��26��M2s[C
��cٴ�\�,ZYP�vоϱA�w��MDU�����i��=.z�-�ן30��z� y�{����mμ�����0L�o�Z��6y!���2*;��^�˽�9~�~�P��>+�uf�a���/�$�9߃�ҁ�0�Γ&d ,eNˁ˗��n�~�2�9O�h�=N��B��3ɕ5���=��ymj�̀�H��K�:j ��X\����3����A�����I~����w���s�>�����2r����=X�L�{�Z���v\���"��;~r6o��8�=�n$6���T�i��u3������L��2>��{�8�2��?����[�'+
0�ь%��n�ʧ������y�yc�kT� צ�k�32-8�
�YuQ4̓ "��%*WiJ-�Xy�!��eď�k��ҳ��I�����ĵ)�uf1H{�?�9s��\zӬ?��9y���K����sHޜ�`�8Q��iX���E�SJ�[^�	�f�6�m�m@o,A�W)��-�x���s#���ӕ�p:�0u�!nM�0�Ҫ��3�辱�~���j��q�4)���TO/+����B�����+��V�D�ƝS�ո�2-�T��o�$���8K���d�?
�v-[�8������m�Ҝ<ƕJ�6��.��	���sݯ,�[�[�H�"������4=��7g/�pO}z�����`nT��4B0a=vn^З���b�$#���oWi{�ھ�!���[�����_���놭E�Mn������9!�S��Yqfc[F��M�u���Y��xB3f�g?A	e�/�9��ܢ$~���)��D�iU� �vz �n��H���q ���yR}�t��9)-�:�S,�_DNV�$3���s���� �XK���;�ar`eD���	?+�,�%׳s�%�ٗ�D��i��uZƁe�B"|�#���P�2-�$q���%�A*&�����kW�?_��7#�?�ms�mU9�ߖo4.O-�U�Z +>�@���^�k\?��14>%	~�����BK�
(�<����5�lt(�ب��ޚ'M����)p})(?�h����sowP
脳�.������!�^��!r���ܜjxX�-C�w8o>�!��Yǒκ�R�v�5&v@��x�W4F/��T&6&?\ >���h+�l,��IO�	�ժ+67�zaM�ޗ/�
F��26�J�OG��$�!�{.�k"w�Q��sB �����?�����k�BL`CW��0��! ^�y�����������ayd<,U+8"���l��-_�}ys};�ټ\����a
��h+�4h97��7F���zmՖe�z����X�Z_�O�}�y��zl��s-7c_�8Q�x��Z�?�(+����PLzXCU����p�P$c�R%��nAm�EoO:�D�LK�x��U7����C�ȿ"���W���EYN&w�n��T�]�0��o�&�p���������_�p��8��Tm`Q� W&�����i���ɟ�k�ݯ�#��F��jx�Wa�A>�\�����<L&�=Q�ʵ����Q�u3�͛M�����C
@��uKn�{��������"�\)�n�28��$�YV����/�<e�B���B.{��������X=��]�ny�Ol6�أTI����P����ޗ�v��&��߸Xͼ��A�r*�j��d]��qg_��4g���h�fe�EV@�M$����ަ5Q%������]k���=�TKS�rgbMa���Q������$����wyr@�J���Q�76Ȕ<�iML'M06,�q��<j�^=}����'͌nm�Ј�J�߉�Q+/��䁳��_Ii�ra� �1N����R�@l��I�D�� X�� ���Bxd�r�r���5*>=�Vk��h�+ُ���GSȣ�g]�;��M�������ro���oᒬ�',�[���lr;���.�v��5 �L�*"��q�͜�W��sq�/>�*���� n��R ���N����5G%��B��(Z��V�k�c"�w�f�
m|���;�g�Qz���kSVga(�<�ڰ ���	4���*�J�'p�mԨm���A�����U^�a���kl��̒.�A�ט�k��L|>#F����Ɯ\yn���|ۭm�H�4.7 �D���	����R�ڷHO޷6/���:����`���d�����7���%^%a�^�Өt���� ]TN��/�[yr�syS"���|�߁"n���2O�5k��{��{NE�)�
�ʎgv���kCc"��}1�����ݗ"��n�pR���=�E�,�
��fP3�"ז��2w~/����J�כ�.��R6����v�f)�c�7Hd7���F�v����s��C��6����~UF<���8�+�:��M�]�ӈ0�y����d�����J�T�͎H�!��:�æ���G�4��)	����Ĺ���TwA�����U<�?y�%����$&��LPg�(���*����@�|�����a�cǉ�/��DLeHn��̣����m���W&�轫=֢�K�J�8�̀,0l��~6=}\e:��Ǔ�8����W�
���m�6b?.�c.f(��� ��kĵvI!F늖{+�Jo} ���@���>���^���چ-,�x�ߎ����̫غ�͓��P��&��՚,��7������g�mV)?��'�M"^�z�g�.%�΃;�6ȧ.�hV��z:��O�6���ͻś��_���=Q�"	s���_��� 9�@�1���}�m\"3	�`n�e�~�_�f��I�uC�2A�:Ć(3l�i3e`�QA��K����'��?z;i�o�K�'�֗�v�I�+�ͤN�א^��w�JP�6�b�W�yi��e�D�.�X��c�w�A#v%�*¨�>9�d���O޴��`6��3fB
�����rl��[��W=����j�n�����w;DtE��p�.�V�����!`@��{�(�"���*��䎐\oJ[�)��y�TK8��L�(ū�z~;�B��zE�*0AU�xz��dD�Z�3�A�R�m��ʚ�������s�B[�������6,̜ɍBR�P���_�[EO�KfL� >;*7!焽?�e�*����!x��PWN����5)Δrq5�O���mHK0�G.��R��~,��G������������P�;AP��p��R����X�5���X�Au�O�^�O�D�7<Y���ChE��6�3�����딯E�Ç�g�^�zW���ڒ+%S\@�
z4�d|a\���un����0m?���!I\�>J� ����L�/���ɿp�.�m��Y_B1~�Z>�g&;�Y��Jsz_��.��_F����A�<�嚓C����%�����҂�r��p��8�emi��.��?c�t������b9oN_��@�W�7Pݕ�'���0�.Wu"���tUb��	��kZj,�T���o�!ID�C��t�F��xvQ���
e�Y}R|9�|$�N{9jF~B����I�.��|@/}�Q�E3��ft��ȁŘ3W�L|���6��G7r�f�Z����4�+��ܻ\'�)�o�ߑ�|�Pt� �BW����X���dW�@��M�M���M�2�^H�K_3:)y|C�ҟ�l���SN�����p��1N�=����S{'��ݛ��K9���w�®�&$tY;V�{|�����F���82B�&o�KA(bc�s��
��	1����h0��}$pKÉ�jU��U�(<i4�'HT�I|��!P���d�+��'�./t��ɍ�_L�6{�E+E�Q8V����P��|����$�h2�8$X�Z�=t�-; ��]t�B`�p�	�j*�}ko���]��)������V�����Y�[�U��վ�0Z�=���Q"���}TIE'����������BEW
��M?@ ��>k�y�b�L���j]�#�Ҫ�KoW$p���QͿ��s���#� .���"\��m���D�R@��J�U�:��)m��������R5U���~q�y����{z/~�/���F���n#4sB�zӬ�\��3����1f9y�2��X���"�W�{�_�;f�;6L��맳k&K5\u"B���c�l�!�Ikթ���A*k�V��NyW9�����)-m�����'b%<�B這#��M5���Ĺ�P�Kӝ�u����:*�#����{V5b^<ѹ������z"*t����Q�ႭD?<x6܆>\��O�&�/�y5�hU��j�A<m�-q�W_�D��t[���"�X���ǩׂpic{�E��d[�u�n�l6Ȋ/�q8R����D_����쵍j���A�Z����~�G�soz��F ��.y���}{�zT3!?;ѯuu��K!p�Φt���?4A�N��|zUSo�IL�������4�������]d�;�k7��Z� p��&�:�� x�^"@��=��D��r��i<s�뛿q"�j�~�`U�[�	V}-3����a|�%f/����������J7S�ݻ6gw���>����5��Gh����x[�dlV�(2mo�OߪxtD�8k}z���]�D�xRy��3���U�m3v�D�������e ����F�ѡ�����A��V��Vz�]���_���&�j9� {,�N^�ŀE� �,�Ƃ)8twاWk�1���MҦ^�j�����sqY�~6b`��Sw,|�k��\W�3�DdJy:��.���оRV ��B� �p9v���ȹ�XR�g��'M��x��9��Zh���9��(�k���7h2<�4�چ� �J6Ƒ�2�j��vȸ�1n�c�1���>_9����	.�wiq����lT%L�SKIz��[��3;�$����yh��J0��k"7KƄ=��duBpԬO(/4=�5�Uy�����:d�QN"��8JM>V*�f~����(�A:�Se��K7���ihZ���d@�Aw,E?ӗ��Χ��u�bYkŪ坽Yh�,��e���o�4]`��hOE�T�.Wi����#}���,y�u�����`���h3�����)�6�y�Z�rw����5O����6VU�-�KM���<��'�B�J-��Y��9I��3G�(eNW�Z�5�
LK}a2�V|	�$�_�9y�!,{(, �n��zF\s��ⴲ�V&)	��v��V��� bHN��4J�����5�����c1>^�wWufw��46�~svӽ�����ʳh#>�xHת����h ���7�C�G[0N�{>*��5Z!�A	�A�i
=d���F�<���p+�����Y��J�?Õ��?J3�`z�?%�Y�����,���I뻞ea��iܸa�r�A@~��#j���d��!ZC��8I��Ѹ�} >�?��Ak���` eqAI��"�[��4�,Z��>�J}�$�P�Ct��"ӳPݠ*�6��H&3��-$�)�Q#�ٞ��S�<]n^��1���Ş�^���T]���B���Ӆ�m׎�f��t0��jJ��ߤ�N/��K���8Et�1�`P�ܵ�D6V�Y�?���Z#�q��������&������y�����B���8fAr�����$@n���Di����[�XN޺��"�SỊ�5=�{�q+k#�C�<��N��������D�ؘW}g��5�p�~d�ZE����)�����~��
���\������'�W�ٞ! �OZ�� (4�F��SW'�MRy'���&K�R �SH�uG�\ܘ��^�Ӕ��b3��r)�G�7]0 q�Je��Q���E�D(��G�\��|���E��i�~У@�yW�	l,7�	i�q	�A� =�Xdn�u6���d�΁������n�:V,0F}�[x*+L��
/�\��R%'��^��(���R�Z=z !�8M0u��M��Si	�I�8٣��z�y϶�ؕ�y�uӱ���5�Ml	��Ϙ/�����|��-$:�?+��-����
Ƭ\��=�g�=Jq���)�eP�l�D�Ď�KO�������BK,_E#����*� MZ�&^1-�I(R�f�ME��9%Z(:����H��Zvd�N�ј���������d�PX��458^��_򵕗�4�Γ�C�"�f���� Ô��z-�Q���Q�����{�Zy�퉔f�+�[�*�${�K��%B}���>���>6[������2,��,�����v����<�[�����r}����%ڛz+��J�ɨ�R��-&"ˆ`M�he��#�4\���bАR����dZH�����P��P_�|Kv]]f��P��;��H���P�T[d@�����7��EMU�o)�Yr�"�e�\��u9 i�TT%ʓ=�J7���C|�|�"}���zA�%�%d3�#F�t)F�L߈"ڢ��H���k�R�w�^v�p�-f�����׽�뢳y�i�pmj�ƏfYR����j�h+R���EM��a�w 	�Q�0�C���>V^��y�3�t��lb8Q��v@���ڧm3$�NXC��?�T]�E�˶W�sU�{�0~m�[�P�D�J�O~s8��0�pQ�*�V����ȋ�x�a�����Yև��l�P��� ���}�46�E��P��;3�!���ʠ�W�ܢx��#�p��&����>�G�pN��(�%��f?k���?>5����<\��Ȣ�xA,9X�ާ����RU���h-�3�u5�r�)p����,?��8�Z�S��[��ݡ�q�E�BZʪ}S8�j�T�a,AA�M?H[>q0���x2^��IMI��I���Fn�b\�� a�J�}n�~hW(Ff�g�_�l�8� �T�s�js�<Q�)�;���XZoR�F?�'��4JF�0���xgGX��>�j��1��4��K������h�t�X����y���/R8��;�n3��d�
{э
p�E�<d)��=y-�u��tK�e�U[4"
�l.�0CF-y�_>�i4���N�ȯ��ߝ<W���,L�LKތTl�)�5N�c:�a �͉�>�
�-�A=q�(L�f�$U���˄�k�f�����6�$;ɨ��0˗�������>G�xP ��&W�0�tkp����{��C�
p�1ѰYKӓ'���e�å����I9X��"ĺ�3�IzV�w�t�c�� 
4�~-� h�U���Z�(��`���x� ]|���˷K'���;�.#�||ĸ6@|�]hJ��+�g^/�S��F�R%4}(��P�F:��ܮ���E$����f�k�mA9��1a�N`�$�����V;�^[���K�b�����p^�x����z,�e0#�f��UR�	.��}�r��V�^�,��g;�J���t��uI�Z�������2]��	{4Twe���+�+2_^sz ���H�ImU��.7iG�z�c������ �'_��י3 ���b����9�`5[���^*�ᶕ��(fgmX�؄�MR6�q��k�Dr�%q�o����b)י����?M<2H7F�Q�޾B'Utv$�D��G���O$̅��8J���G`6>�'�)�$~ά\+@c`%��xUl�x
OL�7!>��0tA�wf
bl�c�7�|5|��S9oZ�D�HQw+:��"������0�e��&p�0��$ƫ���h�i?��,�1<���.��X&bA�����{����u;�7a������P��Goe0��I�����Z��r`uƹ����v��\���x/#?�o��!?��������E���$�@P9�)�By{+dh/|t�1�Fo�9
9�szh�[��<�ge��SF�yI�l�c>����q�U=0��u֒���#��:�@�bSs�X�}Ǥ���<Ǵv�дX0�jɶ=Y����mHE�x��);?5ns���=ze��O�(�:q��G���*B2��O�3V <����/5w�f=n��ڕ�wR{��guG��;V�D0��)5�6��$5���Q��fH�8w�.;��(��Y���C$���Ή+���yS�4oz����#`�
���U��h��]����խ�/ ���Eҿ S��_��omv��Z������⑴���f,��^��&�@rsэ<-r�]�-P��?v���)��Gق�f��-'�p�aj�Iuc�j"V[�k�ƹ���a)ry�������"�/߉к��GCM�$���V��4
�vW	H<3������m��	+��55�d��y����0��4`Jw�U�*R�\����d8�=Nk>����Ĥ�0��c�:�,<$3o�pƍ�^�k�b^�H�<�S�
�m���J��ۃ%���Z����s����Ŝ9���7�����;�kOD�ThMzT0(R�f<�@P"�,��݉>���05�H�>1	�{��3�"o�(�� �?f�� iJA�Fާ�.�c��Z��gm�j�s�H����_���a�,�-
�	r�L�9Qb:�!s�h^���n�wdʘ��Am����r&Os�U]��a�'�ug�6�􏦃s���;eBb 4h~<g��z����O�Tfa��A�#�eƤ���EG�`?^�lu$J��y���>;b�B�}����ìo@���ڌE�4�1d�]�i=�g��34/tp=��=�nL���>��������lc��Ѳ<1M�f�Y��}��!���#T�ơr9�G&/YPpzM_}��ؑ�H�J�����J��i(`G�4V�Y#��.^�9yéVp���䏯ηG	y��b)W1��3��*��$O;'�r\e ���"te�<�J�^S:���6^�ī�pqQ��*�����Dl0l�{u��v���s�#�Y��I�ٗ:Inr�����l%��O_�;���8V���X�Cd�k�+�j:�+�@2�h���h\0Ђ�v�9��\[�fH��R�2���6��H��_y�`�ŗ�BZ9o�oT�4�}|��	3��C�<����$>�Q�/S�
��|�_�H1���9�g��������v��ڗ�9�fR|)=sB͓ ��ƿX�a�ܹ�m�pMYaĸ)~��>�:���H�q�$~V/lb����E�"��6�̂f���D�Oqs�+E��!��Û��Ws�wey q�bID��EJ
��R'5�\q�2}i����=ge �B?A/��s
"x�'�C�4��o˞-��r:��o(~KY�0���$k�����I����e�����$�oC�F=��-�<��l%��|�{z���v�r׏�2�"��Y�������z��#XS�� y�
�����;nɰ�dM����� n���Ik9�ⲙ��q)Հ:H��8e޽d�i�h�У��N��N�EAp�O�@R�Rz�uP��Pu%6*:��&����t�lv�ڿ�z����c��վޏ&�V)m3ߗD�*�74����Du�a��dAs�c���'t8�p2��L.a�mHG�(�*3Hc��{�YiYl"����"��?��(�d,��2/�#t���?=��L��pA�,�|)J=UIEO��$}��a�؏�"��!+�f��wO�&�ŝO-8�i���w��D|�+��ѳ=�����N���e��?R.��(JD(O���ߣA�����I'����5�~K%��S��������-��g��[�D�j��{�7�b���Oz�"񲼗��ո4]�1̞�K�7�.}�ὗ�c���~c䣨f���[w��P>��b��m��^���8�M}�it��)�s��J��Dl��{_8�;腁[��)�!_�pv7��5p���R^����ڠ��(�ԮB�R�x�`C����lE
ڤ@��ȫ��pw����[���㔗��ڼ
��a��_���93&ID����ƾh4r�RH��=��%Nr]��b�Eg��o���:����F�߅J��Տ��Uh���u-�t�2�kG�މ�b�Pu�8�Dդ'0�b�Y��'��^�<��:Ģ��G�ky�C0;��hb��ah�mlw�{�������OX�p8au�_�t��c��S_�	D�z��e����!fւ�ʘ�_s��i(H�&&N�����1f�JhS��9O
��X�ɎA��(͂���Ws��q�;$����H@Ȥ�7���!W����ĆW�L�|�wm}ɥ�������'���9,�<�������S MOQr�������VO���؉1C�Q0B��
t���t�߂E�v��q�fL�P���;x���Ru�#��OR�q}:���*"��*-l��i�8�u+��F|6j�pU+�/�� _Q��GFE�u3��ڗ��$��\9-�V�f�ޱY��{�����JQ��W�0/�N�-�u>�:B�Ι�s���3c37;�l��!��W�nD���ZnY�z@Km)$&1V����_F�~�YI
�^/�C�nu`8��[�8��j�
q��V�?7ư�iHz�r�B�����Cz�w7T<���dL�A�1i��r���U����R�i9�A�b��U���F��� �B^ſa�{c[+d|�$�-Ӯ5-7�˴�d?�:,�FB�t(b��6g��53�ҰeO�rQ�i��4K��f�����
����q�Xa�>�u)g�$���</<�1-~ ��L�	�q@{��A|j0&N��	~��b��T�Ǡ6��l���X����ҕ}��A(j��#!��l|����X�ߌ�@(�D4x0'�P��f���D�O��F�I����'z>�yo��L�t%���=+6�M��@QD��p&m^p�����=�7#�E��7Y�m�X�^���[:%Dd�)A�QM���-	0�������pz}��b\9Ѝo�fz�M
�O�o���;)ȑYsx9u Dj�6��0���I`������ȱ�91�L�mm�o"��Yn�W���X����[��P�����ӡ���E�̘�y�@�J��P�#�ޥ�� �W����N�A0����,���qm6pբt˻�t��K��<l|�ܱj-/k�_n��)��~jQ$l�KHm��ʿ�[� d���9�T	�	l3���?b2s�Tr��-�*!��g���G��	�TCG3�+��
�/3[�r��,���~�Y��:K�5�;u���{[
���ݵ{����B����đ�m��z�3Ѕ�pк����6s�t�ŹU�c�/������s�j@�
�<�:�����ܔgR9��I�7H��y��4����9�#��H\����}�P�_�׏�S5��E.ꪷ9���AVC������1��oO�JR�B�������\��WF�:��8�#d1�|:�� )Ƙ>���}M��� G�L��t8nh�I	Wu�k��cc(����n����Hw�����H�[�7_�Y0y=���sO�Ij�E�2(�끎Pյ�}�N+lgl�ޣ��%Kp��P���t����t
���\�"�)�3J�+��������,�X�ٷs�@� nSxGpaO���J��E��u<]_⢰P�!�-�o��f������l�q���w⥃?Q��D���@��tV*�K�bЪ�Ԥ�Lܨxھ�B�<��T1�f����J-�0;�AΑAx̭M9>��h��������Y��R��]YB����ۉ���+�f��g�/�0��S� #�[��	��z0���n��L�,�S������ϩ���_..��]ϟCt�x��a��ǀ���|�Y8ϖ�9A*Ҟf���B���n�Й�\7��� ��xX���w�Z�`o�)��͇p�)A%	�r45��l^}#$����U��ta��W�;~aO�,���6ފ_ڕ�#2gq��`s��C�A$�H�J�V]uTp;��V|n6a���kL5�s.�[�"gp	��X��i����a'>�KEb bl�&��p�n��HA��$u��Lj���L�N/Bp��ŕ��|[R�r S��W�����:]>\�:�
>_�@�O�T����^�8cH���D���$y �� U��T�%8���0�4��x ғ�7a�f�ۧ@.�Qyk�b�Ξr�F�V�w�w̞�y ���O##� �X�F�S�"�J6��ީg��r���l:KOR��%��W9z�nȝ�/���)�GuO������j5���~Ai�k"�S��R����l����B�-_j8T���d��׬B���ľ�0"�%�!�5R>��h����[HI+BZ�u�?P/���Pi.�̓�H�%_e����jÔ�I쪍!�U�����zvDԧ�������U�G�jq0��lu���zc��'ƥ�f���*]zʮ�����.HA� �����TM ��D���V�+?�!���E1Q���˶~~��t�K����BW�g?�e!�[(f�a����E�$fn+�v�z��ց�8vF�A�y�'�Ox�hF;�<��)�4ai*:����G�yC6��}s��̿�2,ӠX/� E�ԻNs9��E�3�sY�ٹ|�[�M�s�3��hD��6�;��Z��b<%VG+���������B���U��M٢��K�>�C����}9<�Q@�B�8����Ls?"ajcC\`��u!G��gytwn�#3�m�F�kրW瑮��ӆ�����/#orH�mAi�����~�,��O��(�,��&��g��(�J��+����}J������Nn�$��s�LX�dA�#�[��_G~��I�����#aC���_=���!��zD>���8֮��e��T��\�D�!�H�Yv&��$��(Buϗ�Ůp ���P<����o>߯�w�-=7��9d��^e9��p6�`o/�-��|��ihZ��y�gr�{����@4�]�y��κq�8�ۅ_R&?T���X���&�s$(�^gDx ��-��=gv������'N|�RQ���¤��ޣ�{9f�H�Zn(*��'1��BM@	M���ƌ�ױi�C�����8%�&�[K���e	�����͉�+��k��Ր�{"Ɗ6�ԅ�M�abN�p-]����:Ƙ�\;�!�۴LY"�7�]S$Pp�a:$��0$In�	�:���3*ItЌ���#����]�틀	���vUa��8�=�9���=�Ng��-��S�X���,��wX��6 �*Z��_N��.D�y�h�t�V
�S"ק���;M��"t��w���:�}&fR9�j���ě�gQl9h{�ڟ�I�Ш�B#�{ /x�9���96��3����� [� R�E�2f�<����&.�Q�)����q��;�߲>z���62��E�%���}ze3��2�H���|���A<'m����CK���.��� ���B�ۣ���$��^�޺:R�q5���i<_C+j�<��,;Ho	kc�z�(B�P����FI^O��}%$���3-�+�#�'������?�X��!<
?�"�gb����G�P�i�N�B���9�dh�Zk%�f��A��+K�L�����+#����M�d�V#:��3r3�v8�1�GA����ф+�)�.�U�-i��)�'.�a�X8j���m�<��H9��w��ۦK�;Rk�Ç ��`��Cڝs"�	�,�G�B@'Z��k�ra�o $���e0��Va�օk�\S-���I��4�o�H�S2�9�)������ jZ�l��H�sy��qΎ
�9�H8:u��6�o}�����ͦ𠦷�[ޛ^*�"�r�2.�l�?W:����@\L��y�D�֓�Ol�ݭ���hh셌0I C�Ϧ'{6V�a��I��(��|݆��E�6Y7���L�Ϧ�U�>
�	"̬�1��_]�����#���i�=gxuC�%%1�WaM�&���BG����\�L퐟��}:���%q���S����&\V!RzL�>��R��ś�"���Ne�}�~�B>�Z���� ����Q~򲂐ETԕ���=5��W�����D��T̼�\Q�w�6��ʈ��}�4�E�	U-(�;VF���2��+�͸����MI���w��Gr�P��C҆k6�H!7�ⷙ�Oa����S�9�5���~m1{��g{He5�wcVԱ���b�⒦������czP��f�Ia7��Ի��#��MI�¹�.��+UB]�.�f�Qh@���0(9��H��(�E:�)��3r��Y��:��=̽J�	�V�ОR�9��a	O	���x�8~+/���������	���i���۪q)�Q@P�a��ȓ���P��c+݋��}�8[�xi����}���cŏ���IE���w/��R������:�Mw�h�o��X��W�N��s�[�M�%��*�4�� $:��_HĞ��X�@Z.i��V�v�pN�t��;j$cqڊ�O; ��N���+s7D���G(�{��Q\������F�Fo��o�O4ڷd"|���>+�4f�ᧃ=�|y�(>,
C/��I)e��I������B���=o��N�*%Hs��G~�����O�{��g�F�	�w�ob�J�-��'<�8E���G^_g�R���ʠ�M=�%�]��h�ډGw�=�걌>Դ���JU�XBp���'��� 3~�f��|*=\�h۞kK���9N�v���W�r����������i!��PKQ�3���MSs�2���C��nӗ�kV��*�2ƍ�>�L1�o�v����N�P��@WA��䧧�0V�������	6G˅�CW%�6����_��K��ϊ�`��aoSp���J��Cƴ9L)�uİx�q��M��������NJ��rX�p����"��#�����V�K[Y_X������\[�:��2�M�˙Gt]r�̂��'�#�zTR�4.�7JC4�J�C+�sZ.��p�E��!N\(3U�4��nݢ"�P�d'+�u8�Y�f0X!��J�~��<�Ůo.JQ@cgpi�z|��lSa(�{�l�@��!�<�Á
��Uɓ9Ը��3����R���C���}0eIY��d�j�ZU'P�0�o��h�g;˲��}��ǣ}i���Д1������OhT��=(L��k(��XP}t�6���OV �g�x�+3E��7*X,<YT���J���}�t��zW��r�� ���.&��y�)GF<��Dq��n����"��Z����9bz��T_~�QWc�� �c��0z�03ȱ�6ze�Z��]����.L�l=S3�bl��ر�8�k��!
��d5��^�劔ğh�Z`������&�)��� 3�-L�0�[���@F��W}Z��,�8Qh�$�$�z�[+�����H1�]���fT��D����i1�){��d^������Q�?��9���ʱE�3WaU[~���a1^Ԁ�2��ʬtwX��b�b4\:;b�ɂ��aa�%��	
��g�8u �A�O�}V�b(|礀�>�Z���#�������ܤ��Z���8)p<��s��b�Y_ ����T�3�,#v�:�}�*Ѹ��"��d"��\�~�(�O)46���;���:��Ym�b�(������L�J:2�v�z�#�pE[��\�8"G|��z�[������kȗ�L�.������EH����j̓�wH͑��rrb�����.��V�eG�z�C똰_��G O�s�����Vn��%��ky������R2�}�q��9)}�8rl�R_�uBOf�,������Vː?n���=q��l�w�	i�h�ir�pH���$p���<�@ۘ����e�m�7�PAb�y�*tY�hX{X{���un]�O���0UX�x�5�3Q_{�11m����e��Җ�d,�7�cΐ���u.�$��a<��n���0����V"8b�2w���|0�&2��b�òv�k/��jk��.Y���}29_$Jڲ�Z��H����j�]3#5�� t��8}����x����- <"�
����z�ɔ����oJ�׏�v�Ⱦa"�t��M�n@N������,�<ɢ'��3F:u�����]�ýje'���qv�1��t�V2ϙ�p8�?����D�/��0��8����f�(�!��oE@���eh*����l��I��,���m��XBi���N��InyĖ��c5{幵����� <���H~��B�m�[c��9.i�a����k�
��J������!:���CjF��m���u���Lķ��v~?BAj�K���Z�ҳ�˴��z_��Av|,�6b�e��GnfUE*iHR?)S�%����?>���Pm�n���{G>rM�#y�!����������5ۚ|6��)�9R����0ƨ�I���fp��.v�V{�T)�8@cɞ��
��X�'0�����W��W���(^'ÊЮ��?�~޾��r�<#i��!�;�+�0�*m�|�z�)[<_f��0p-E�����0���V��o����/�6��w�K�G�jZN���,�7�T^�HЈ��?���
�4�5���}#�Qk^�;��Ze�|���LAS�~�\�EAQk���!IQ�(qW���Sy�5I��; ���mU�[�R�{�-�\�*V���..���
ǕX�1���g,wNRC�t�g�7��Q2?MPX$Q�t���[���ҭd��.C�^-���h��zy#����{�;�I������h�ӱ���k	�k�R��[�U�P^A�m��?`b-���+�� T��(��ś�UZ	���o��n��O�Q�ǕR� ���>q�l�¾��DJ�-;���b*���W��,�g�GN F���h%	4��~:��/=
���J�X�S�/xo�R5H4����>,�JҜ�@��7S�$X�0�W3���]�J��ɟ7����m}��T$r7=Tg�%�b��&]^��w7��Au&tء��w����<vR%Jm�S�J9>%1;:}��E���v��;��Kg`�B(���y8�$c�?\B91���:��B��
�!'�*q�-`���?����x#QaQ,4�:�0�ȷ�,�Q|��Ÿ����[�e2�[�I�NhSf��<la��f���q��n<ciu��{�)��0�܅�s]��wF�6��>I��sֲ��Hbh�QE�<k�Ű۵���綞!!��+��&:�]�j��Z�Ω����Vw�H���wxu���Os�Ozם��<�B'U�p	v)�g�:�`��qS?����"=�h9p��+0��2;/G�^�B�Y�"!]��`�|z�'#-����:3�Ǖ�����|�ע^��؀��S�}��Ja��,7��0jYa�M]��ܟe����`��[��=e]\�����0+�zioȄ��ҁ�Ƙ3x�$v��=��4����n��� ��������((�P�-}�-�꟬#
w������L���m[�R^��թve��9�mrº*�w�W�b׳��aL��>�"s���m�Mu�m�NF)�^-���<��>�p�	�w![#Q�?_�Hu[؍P��ˉ�[�%b��a�NrkJ�]���p8�\K,���A��.���v�u �����zQ��֦q�hz[����e�#s�	���gʢBl�ʹ��q�e��d�+�[-�p��[���z}�dP�i�jW���e�j7�.U oVzuF��/�7;O�ꔯc��\`0�hs���^�B�� F�Av����|���`Q�t�z��Of�ܵ��~�H09z	; �?L"��\� Ǧ����J2Q�6+gmy�vZ���! ��_�m�Y�A�K6h~C������aԉ���ʘ�0q3������ʸ�,Ds��O����}`֠9f
�lj`��v�b��X��^���c���u��Fs��ݶ� �H����rȐ�g����.�[�AZ{g{%Ld,#�j���b����װ�3����Wd��~��������n	�̗8O�,�
�I�����9�a����d+!�^OG���5Y�c��C�  ���c��#��õ�(� }�U�����������x����@��������f�vu'�82#��f��vǚ� �p��<�����9����?�ɧ'����]�`��"�t��*�L�<:���e%%�� |�>�	��#;l6x��^����mA<���}��/"k��vԺ�!�ڼ;}H���K�^/���P����|���>>�~h?xo�߼\b0���'W����
��C֏د�x�eU��#�����@��w�u����@=�Ԫk��]o4�E�e1[�z�����r��L�IU�"��f��S̹�E�R�YE�[Iogk����ұWȦ!.l|ԧ���DR.��iaV0��|�̨vX4�Kc�Vg����m�S��T�{9w|�l����Ԍ}GAe��(��m% ��X���&����[��/V��!f3�oODt�\y�+��3�=�\ve��5,��{v�������n8L��,R�� 1o�L�}7@���8:��sD����2���j��.�O>Z�F \��Y�][���H�3��! �pu�mbulB��@�`���!#A>B��>Fd�7��ރ~�P�u��p*�{��b��y��������Q�0���fM4qSM�ɾ+h�U�L��(�O�/�EJ���(�!��.��������O"�ì *�Oo#"���=;m�hݰ+�h��������Ԣ�I
{+�U�#���ke|`�(mi|��se��F�\����%�$��:�^�!+�$��>�.�u�70k �F�DR	�]�(��&V~Z;�%��$�58�v�o$0�0��m��*�v ki"&��"�9$�LBz���8-��BA����@��cߋ(��oyUؑ�#1�Ȼi��! E;�����q�k���W��1(�(���a�ϑi�*�
�W?�<K�w����Osw��/�頤~��.�B�Z6#4S�Nѧ,b�q�K7��G:DVݫ`�}o*�#h��2aJe���K��
(+���Q��׫u鹇�D�)��#٣���5Ӱ>^�kmk$M}�]K+�c��It!va܀ؑ};�5LU���6i�#n+�n���c��4^y���������piW'�f��\r:�foE��;h�T��aG��V�H�;�s�0O��Y��h�~��}������q������J���S�_4�{D]��ܧ��]��y/>�[8J�����X�&AZXd�Y�>1� �G�?7�6�z�uJ�A���8D�R۳���4���Y���}\���s��(�-�37*�-CN�ʍ�F�,�C����!(i/��R��|�-o�c`���Ɣ�_R�>$q��3�D*B��3�XܞGvBS�IX%�ӮQ�h��~�.9X���I�s�8�z�.��-�����J������e�j�g1�1|�γ8����I9�ҭ�s�Hp��J��v�h����a�^G��a�6�G�m`:� ���R�&y�N� �K�*ت<Nj��Ѥ�$�O)���C��	)��vqS������ K�ɵJ8���v��@@(@拱��N\�q�ei��bx�p-QQ~�"����=-9dmU���֠��iG�VhD����&qަ����
��B@FC�o�s����6�U�j�9�e�ri�34n�+ Kq�[N���b�CӊiǀZ٢n��ZӬ��SK��!�<�#�+E���0Oc7�ߟ>"B�̎�A��l��o���W�!d�yQ�����th{� ���}y8"�8�M[���U~�L����]2��#*�۽�j/#P���ʡ|d.����.=NW��Y"������B�n�ק�٪{. T�-��@��	y���9ּ�n��ޜ�$����C�j��x~�2�b���f0�����B�xe��� %���B.`�5�t�z��Ty�2L,���g��aݍ*������
u�֓T�w̴
fA�^5���]G�k�F٬���ܘJ����9�!��돳%��-�m�t;ǲ�,��8 �' �(�M|���;XusbC�J�s<��W������.�'�QI�����~���ޤ�_k��5�,"��Rl3�⹆5o�ǜ�� �Tȓm&�W&3Q��լ�K�Bj�yP���� �\�`�
%��c(�F��b��q����"���AD#ٯT@p����ěrG��^!}[�4,o�,��+,�O't��8	$ F��O�p1;��a2r��d�wg��!�47Za��e_M���MяMj~󃻋ȏ*�ʬ�^`E@T� X��o����
l_�c�C��5��XBe����o�~Ԃo-=>��6v�B�X�=t�8(�3
$�}cXF獪1�D�-8�W�;L�	�����H��.:G�_�Y�r]17b�`�;֚7uU�c[�Y�����V��mwq�!2[Zc9��o�ka�4E[��=5m��#�B<䛮�>��A��h��9���jX�k��D�����஀ѱV�;�1q!9�X)��&.��8��u�
B�a)g������"�ZK�2S��u���^���R��RŤN��@JҔj�)7�!��7o�d�3>��[%
c��,v�D`����ɝ�N1<S0N����%���n���Z��_�=�)��	�KY�D3u�;/��~?���
k���!��/#ym�3���Vyl�5>��gz��	�y�9�''�w�e��v��y��Ӏ��`B��(8���K3��B|"sr)I3i3�x����E�5�q��:4~�B��\��@+�)BA_s���Q��?_���k�}'���	B��v��f(���O8�@����3���+���Ն	��+��ǡ!R|�[�Pd�L��*�QX�ܰ�K+�&0a3��-"���y\�j����k�����M�`�����A�$�c����ء��&��#U��j�B���e��R��/[:�Xb�¸1�>F� uh��� )���!>�_�բ��r�*�[~�E�`���)[@���(b����g<�Vk�����򙔉���y򏆅'Th�ߛ��F�v�:-y�ĠA�̉�>g�3��c[Q��?�<�4A]7�b�[���~���V��	�=~�o��5�ix���?�&Dڎ��(�5=�_�����/��<(�vl�O���1�R:�&�0�G�Gq���

��3q��;�|��7�E�}�BmҍI�XĶ���-��.6����O�TM�:8��0������K�&;P��*G�ow�D��v����X �#������}K-WsSzR�4��1,+nb��3�/����̰'?��]�#�����?'��T��?��c�(��T����
p��ޮ]�W�"�0Q���c�,�N2�3�$��e1����7L�.�T��~]�$:U������]R�y��͇�i��w�o�� (��)w�~nFjx������6ee{;Lږ���3�k���K	�9�rXtG!�k���K��gc��S�)����z_8�:"��/�7-װڧx�S3e�W{�V��;���=�h�(�)�*��@���ks4,��~���̃f������=7r7 ����E�#Ə���=�z����c�yI�ě���֊�la�Ԡf�ū��L�K		�D��32{�L�J����h	:��s��CHȏ�j?,J�����1���c���r��#�[b�5���e�x
��u��\��%w$Qx�d Jz��}X�-�.��0'�o "L�O��˺��y���4z�E�9'y�H�1WB����؍�
C$>�t�|f���پ���^�jE�6��ĲJyI�\��q7>w)�\���7���2�����������w�l��a��I ��ى��#�0w�18�#(A�V�w���0�����&_�`�H��Ø\�yDr�Y��e٤á�)�Җgk"��;�k- ���*|�������Y,�|�����w�?��$^���g6(e�)+{�U��3�v�絨�
�eoz�
����I��
%�#>���P;iMr�u�:F���I�%���j�.Wϋ��;���Bg6�yl�BwC���t�[�*�n<M���)dmq_�.Up��u�n���Opȍ�2';�tk|@t�$*�̔cJ䬞�x��U���6[��Sk�6$�O��a$�c3��9� o5Jp ���{	c�0�����LX�P��F��AN!�@4�,8�Z�!��X��n}��T:����7V;���pF��6X#7kX�ʳ�;8d�l��Z!��y���!U���Rފo���9�vC!���|�t'pQ%�A�>Q]S����yO0EһT�L��P̏Pe�m��' y}��r/G��B���.�&'9'̗��1|�1���)��_�
�Z@sU�[��~����*��̡���v<	��}zlsSU?|�}t޽�w�uՐ�ip=Nd���w���u-V����FG@��$�!�2�A����}0�-L�N���v<
m@�h�)�㍣�lZm� ��qe�byQ0����[��:����kN��hV?Ǟ��H��<*vu�w�R����g{*_�P�n�2�8��Nr1^Q��M[;N��Cr���*m�gw�й���q��97OoJ�ۃ�];t�s���̾��w/�+/��c�8k��g8<�"�4.��6K���Gh�ؕ���4�oySF�a��[����@���\"�'�(�¯��\�=o0_<��р:��/����!���C(|;	3���Џou!Cs]5�@ ���ĺ̓��~�Y�����cY��	GwE&�!5,o�����HPwmw�}�)��Ţ���.f��G!���M��s�C�騨�_;.7�E�;_δ2�k!&=}�m�y�6Z{��l�v��VxZ9g`#
��\�rC�J�(����ݵ�&�k����fc�A��?-�M�<�z��*�'[:Öm����\f�����T����/������/�J�{I�?�����c�}|������%�}�44�Ɂ8�p�ˁ�ZL�H���P	��ک��a �Jͣ�%����g�x��19��$��k^�j�=�\��98!���J�IK�G�Sf�e��r�"��q������a���Ӭ�U���2L6��R��3n��"�:�߭�`�%2�ћ��,�0���0V/�7�~��#e�=v�����O��T|b�I���N!t���q�	y���5+�P�(Y��V> �)&��??x3���D�K-x��#��QJ�À�C��جV:]G�Wzם	�:j�2���&`�ti3������V8�@��*$�H(�Ϟ�c%\�חI����jS~H�-qU��W��8D�R;�7�uP�Z��7�g�_��_���m���×�R;�5�7G�@p+�_����1ohv�!x��4q�n�*�8�r�,"t-n����Aƅ�5��.�����o�1�C�;ho�ʊi��h)��[]�,����40�"X'�5��:wR�kTϽ<E5�^�m���יk�z����

h<=��!d�|����wd���DR�+mE#�*�!091+�h ��ɳ�8"��۾��T	+�>�h!)��E�s����`,\+��A�_
�j�k��� ���3��Syw��+e�����P12��?��X�,��	 ��V�1x�>N3�uYu�$��ij�);^7���7��=���r*�&ƪ���@8&]l�+�:�r��
3 Y�S�.�_������2��5!�U�BmJ�t>/"6z��|�RP�����A��(�q�#�r���tbI��ݛ\����ǂ0�g�b3͏N��G'U5���!�~r���A��m���cKM$�H��#�g!�Ū(�N��7 2'�e��5
R�jC5[��އ^�u���[R�����+[������9�W�mz`_������ S7\m����a�zW@�Zm�)�F)A�"T���~���8~1τO�x��F?�io�#K���g��]��=f��E$V��7a g��A}Q}h�G��c�R��c�� �4�������^5�N��H��G�l
k���V#�烒y�ʥ"��-�K YA�.^\�<��o���\z-�.�Ң���^�q0�
-ytH��\�x#|7�4<9a$������W��/Z�߮Lv�
��CU$��|cgh���:Ň����[g\�fG���ޖݬ��yߐ��bG�Xq��`d�/����f�o
�HX72���˅��-?C�Q���rH�����%Jv��4���S�$*����)�`H�F�Lh�1r����t+(����F0W��0)�W�:�Y��P�F�%*gt�����;j2[:�_�����GQt���$<�U�t|v@�G�s�_�z�bH姇�f���?f�����ŔR#�<j�Ie{km��Ç���24������y���7�6�g
�g6V)���3�=6�#��Ʒ �'��#9� ]��P��J����3Nz�œ�r4yF����?����L�����zɎ��(���L���Ҵ�Ύ�J	�/v��m�X�vn�v �
$��÷��6/��pX�Y��c�_ۯ��Nkt.n��k�<ɻZ�qJ"/�>O?/�dQ�������]H�Ȣ������3�j�0<1�g�7�(ܷē!�ڎ��h7�<$;��I����VKAF
�Yf5�Y~�ء�I'�ثQ���	 4��.��Ƈ�
�~X*>	`D)�*�/}�X/�r�X~���k=���2v����~���x�K��zJi����p���e�;�p�KP%��,��/�qL .^<H��]��Q����
���ƙ��[�54]���b'�H��#�ݡ��p�%\U�,4|���~*R�R,ڑ�̑��9`�痑��ٿчB�܌Ţ)^l%
J۹u!����N��ۉzX�d*���$���^�y8���"�o��H;��Gr&��1��fp�����N��*Z�=5�4�����=�{EF�Ɨ4Y+�\z��4��!t��Itɬo�(���U��w�@h])u����MČ.A�TYql��dI6O@�V�2�7�d�`�$��XHaU��!DYU5]��]>��|��z��:y`q��<(�K^h#1��r3��~A~����W�,�>5	:DdH��5�9H��0��K)Z�j�!G��>��$ϖ?tq��&ʒ"�U����י(DN�ׇ-�*�o��^�^��p������ė�V�}{E���N\�\��#��t��l�	���8K����u��Kײ1�7ߚM{�ɧ��3�f�'�8V�H��>"6���ʳ��GDs�XξP~�ꢅ#���
�`#l���.�0\Gm5�w����h��;)@H0��wz����y�9d^�;$�E�"G�H�pPǢ��;����J<u	F��j�/xl
��7�u
O��'F[�%�/�yaϺ��^�P�k]Ũ��+v)�V!Π���R�����8ԩ ��D�y�:XQ����Wѻ��?�c�ϫ��f�+�<���ϷH�3�����2G�
��<���sp�ƴU�y#Ҿ�3LyHwG�*fZ��M�v�2*	Kp��:���?1½Zt���*ɢ+WPd����J�nQ�
)�L��,*��ip�WXh��]�tK�\��p'�:����r�2y��
*�\yp��<��%V���̎:��mtQ.�얳�rَ\n��j|�%�+B�΃��%��0��s���e��_�H��B�Z�v?y����ᅓ|赤�f��p��u�N���N�S���3�/s�X�v�]F�_�1��/k�<�� �Q��M��2
�	�e�����W�6���_#�X�tj~�����.�n{��J�Ai�9H,?�z��nI(�;��k��L7'<��#)��I	��<&�j�e�(���h|ko<�i����A�=����Y��<4с;��ֈ�xM�IѢ�v�v6t�	Nȟl����F���P���.t=��w� S�7�2ޮ��	E�mmԓ��Z�}K�=Dوk������J�f-Ŏo-,+��j�#54��L�݃�~+'n��#�n��(�`�
p��.�~�
�yyǫ���5�*��
W�e^.�7�uVLJ#K�
,IvA�*ӎ��U�Q�ի�b�Z'�A��<�ދ���}��_�M���7 
����,�2���Om���T��ۙj��i��4Y��gE�\=����ʀ�V��\.pG�_p��S�%A4���Q�n'�s�[�/��8,�S\UM�
-�����ZxJxki+�#��t�u�re11�=d���)�[Ƈ�K���6W��~H����EK ���UH,�ˇ��f���WK��u�WP�	�i<�$p�˸ @ޞ/�Jڂ~��n����>��"�`$��|цݍ��@��寚�?��X��Yd�+cr��=��
2�j@�.k�l�0��4���)c_��=�
�!�*�УTa�c`���&���^�ofG$~�È"��_���X$�'���G�U�G-#;���%Ԡ��b����=����2���/�8�e���Ϲ��Ĉ��6P�a�I%j�Ǳ�n�е=�#Ǳ�*(����$q������$����=��HÇsV�:��mt���GJX�'�5��=�enSO�It�"�8?�P��HL�ى��f�9�����a>#&W�2p�=�KqMIAtˋS��GBH��xZ��w�U,��Ԓ���y��T�]�g�)���P(�M��$�'�u9=��Ғ�N�1;ɶ�����=��Ǆk��Ed��;��!~��φ�`��V)�#�i �ܓ��n}�#n�k�闉%�����4�kB��X�H@�%�qqE���߮l+�?�Y���O�6��XZ�{�t��@��M��x��:j��c��]>��W��5�D1\0�K�Y���蝍4�.�ՂQ׷7�t��ǖ[@=.*�G�|^��s������yx�%.��Y����2׶(|��a��S&!����E�����u�[HJBrR
��B��k0�7��=_�ݜ�.(��;��Q�� �:�wOW �J��<��V��S�W ֶRƐ �c�:ix�:�J9��]�7�V��}cj�����6�l�o�&V�}�E�v0��=>��as�N���!�MG���Bx���9.��L�S�I�_�/��@o�r��Cܟa����<9\Q'����2��������C�ˑ���1C���.u�`hw��H�o�X��@z�Kp�<��$�ޮr��m"F���/��|�06F<�S/����g�8��T,�����bo:r���v��F+9�w�m���MJ��+���|e�U��N����`H ��Q�l���W��p'��e���O��})�/�7���ɝ5�kY��/K�Fr�K�Ne�I�_}V�p�Y0w$�]?;�+�Z"N
�P]	����2]���>���XA$�-��nmJ�����:�K��?����n�����`\.d�� 8���f�%�椽Kr��[Ί�,�VD�9�.�:ݗ(��~O'�24j�U��S/WwgjE��LJ�(P=o�~�ܬ=`�R	��1*�f�2x�\�^T��oC0X�Ɯ���������"~{��yX�H�~���N��Ց�b��tTO�#A�՜(I��5��t���'��55N�T���������-��%����*�g�A��=�3�6Z�Q�m]'����⍵yHW�B�ޖpF�a�#��� ����t&��qPѷ��c��3�I_�LF�Ď���$�_e��Ʋ�(�dǘ{'e�ސs����Eߎ���0 9����i(mc(|>��+kbe���R�G5u���l��|���X���+�(Pw�]i��-P3WI!3�j�՝PQ����Yu,R�X>�3�1pϓ"�wO�o���m��K�p>�0Y��hKk�^v^����ј��N��t`cs�?��yҬUa�I�c��r��T��U���!�S�۝g�5'J���6B����JRs?�i��ʞ���}d����-���3��;Yv��~���߁I"���ޔ'>Oގ|%�ib�H�h�)��Ե������pk�G5�ݽ��˵A����m,��U��ZG�\_��@�4ɨ��O�~�}6c�~6D�]kū���I�b
ۆp��j)+dI��������]f�$�xE���X֌��qT2?�.9�51�_��m;�d���-�_
l��}�����A:*V[)�s���t;�t��8�G��M����	(��;���!#7�9c֛܋�"R��3N9�Ub'��6�_��%e����R]���h��5�A���#��D�V�
l����>�V4���ӡ`�����Ī�Z��nw<�Ep����$�,2b�x�y� 	��kv�� ������Pݰ4@2q��Ul#�5�ؠ��O=Ђ�O')���'�����x���'�$�(rndl�ӗ�*92�+h��3�"a
�7�ɖ��@.fL�«R=�x]~���p�8�����l
�W�Px�s���^�|�J.��s��x�'If��&Lt��� V94�_�D�h4�z��z�.��X�i����P;�7��4'���'1	�Aw�Ui-&Ao�ZT��a�R�ئ&���\�],2gfw�X�	ʺo_�G��jR����r.��P�q�F���[�*'#� ʰ�u�ÙĄS����' 7�����ܬ�q5�z��@�T����)@�c5 �҈�cVEK��;�C=}��P����t��1$C`���-I����U��]�$w�Q���+d�'n����7P���Y)��h��B5�GCϻ�i���OY7+C�.E�6��3mC�v�=ff���x��� m1h�)�&ͺ� �Ab�"´�{WE������(lY�����ʲ:Q+��8e ;9~�|Ŝ�p*4�'{�3�Il]�P&:NdypN��K[Fǡ}i��fZ�: �BِɆ��Aڽ�K�����T~�=�;���Z�TC�޿�C���/��	���N{Ǩ:���v>�Te�BH<�{�`&2p�������44��j�r�9����\�S��p�lEb�'�SR	&����f���C$�)Y1�u��;�+�N/sf=J탰!�?o&rd|� ����u��Xm\N!����;0bi��{,��[�t�S��S��у�T	$�M���v�f���H� �B.Q#D*q�ث����T�P(�Y}>�u� �@kw�pcx��d��N,r�B�F����Ȁd︩��9d�Pfl�e1$:��#���5P�$���g���������^i�I�p��dX
W�tNʉ9΋ת?�z�}x@�u�/'3Rs��lA���R��W�O���Z9GeG���;�p@�Ex��@����~q^�!U�O�\t�+��@P�^*���ԖwW#��5y�\�H�Ǖ�I9�ϞR���+�=�ܶȊjE����I�ݰD/z�����U��s��3����e�?�T���UJȦP9��I]�˹�{b{XG$��R��@y��S��F������ɔU9��VHM`�؝	ʬTq�yh�5�E{�.�Sf��`�SbrO��s�(��,2uN28�~A����ft��p�m(�"+ꀲ���	LfW�#�\��e&x5\W�3]c���H	/����Y2����H��v���|�|�R�A��b�%�P�~��j[�9WSv斂�8��j6 ���~�����.�<Y=d���Q�/�t{F���70�S����M��T��Wn�7\�X�!;�S�˸��{���j#�f/3��|�t#�E�Py;��R)����bw�䡤��o� qV*;j�=.Jm�/7oL�h@:�����H3����,���?BM�~�@�=�F��O�8 j\�~�i_��A�IE%$a/��� /�t������,�-�2�~�����Z���|$x��I�tj^>����?#��*ꙛ��+��0P�M��FC��R���_���� 5C��ɗb5Vg�ro�2"	����\�)T|${q���y��3�߁�t�����qf]�4��
+*����ű@��c"���M6҆���J�ED�}5PxpϷ�~����$�)�n����~#�#���r%�Z:��H0|�J(#}֢�Rx'���z���P6q�|�jC�֏���Q�h��>��ί%"t*a�r�<�Agx��Ǡ�B"0YZ~�:�<e��n�����g�3����b��_8��V�|Fw��d|��4PL�7m�:���E2�Q�UI���*��]m�l��#���A�����wtY+���g��^��4�[p�,�F��\:B��?)�!��V�ލu�m���ᔃ��#�s����%ÛC��97�o��wn��%����ڥËI�:�n���)&���~���G隬�/���r���@۸������Qfѽ`�j�P��)-4/VO��e�P���X�z<�܁�&7(�oi&���b�u�)�YR�L��!�n�hQR6����v	<��6��<C�Wz����#�Qk�*p� �z9V�.�+/M�� �Q�����~{��j�F��5���EP��(����r��A)7�M�{+sF��E]6 At��[.ƚ6r���='�ep��_���P�Е�[�&��9��ܲ�kTx�D˴���;6{�GV`?gF��%�<�bΔ���H`����pn��rY#	s�L��S?Y=%/B�5Re��e:�V�#����OwӜ�篔��0�.��Wтh�.Q�v�r�.�b�H�S����c�\��m��vٹ���α��]#z'�F�*vq2���x�m\��(:�[4�Tq�i���5D!8��h��xb�D5�)g�J��n�槀�m��u��|��al�59\�?��L��@Y�����+~���|6�v�vB%��:�n�	�6K�����b�eq�����ô�GR��%��e��l���י�e>5�WYB����^Yv�zS:*�k���x*��Du��4�<�b�7v�7����j'���d�һ�}Nk��tx��g�΢�,�d'��v��<�%�"�y^��uJ'�ڂ�������Q̟M��.�A���ü�V�5M��7ʞ�����&�4@�F�H�hc�=f�����X��%��m#Aii��M�	N?-n�;6��i�˯��?(�>+�p��|�]���
]�D�����~!t٢�����H��BLlՌ�Cdi	��@=���t6����pw�"�AgE�qM�)T6�gU��K@޴�)Ra���ϝe���?���;�0U��0��9ǈ�P	1���Ԝ

h�ئ�ሕ+��Zܑ�3����B�U���FQ%*Z?�@I,��q}� 9�Dɫ<�����㝿�g�SwhSTm+�T	�U>�7\�ԡ��H:�h�Er�銓ht�E� ��,�-F���&��1&��V	��>2��	���L�	�O����x��l���]�tÛ��||$�K�x��j�wd醥�#*��l���ʖ�
�Z\���b�L��@��g&9C>�)��*��5�Ǩ�����IjO�5����D��ߍ��	�EuJ�(����W��R����,l,�頭j�MZ�E�4�1�X�#EݞD[4��%�FE���8|jV���@o=�+��$1a�E�r��s0�Y��&&��7Eg"]����4��I��L��>q�?�v�ԥ�K���m�ݓR���Y
ƄD�r�4-��~<Aqӯ����9��c�����Uͼ�٫܎=~*�\;��E����}�iM-U/�a�YƤ��!泈鈣�
a@L8e��D��V�Ȟ���j��z��3������WL��Qo�`��T}:��8��i�E Cg�2�׹���^��M��<�e�8���K���p ⮥��]cꜢp췐�C4�U�ֺ_�4&�GȔ�?U�ɟ�x+�Nr��2��㛆Kff��|��*��>����d�<o�_�),�N=�T��qI�Zك���t(d���Ku�cp�ȡ�I��%u�������<L]�
�H�O�`�����&�7��N3	�x$��@h8BD����6�9s�l1���\��^���$���b_���m�z�I	��P}b%�Ks��tr<+�0��A�זO�pH%؅0����@�5x����T��F��%KtZ�kc�l�+~o�6A�e]SE06��l���`��n����^�ݮJ�OM�6oz���\�\p�k�iK�Wy�Q�����\�C���^^SC�$J�=;�U�"��FǍX�E���P��x�����.��wlU�5̞7O_� ��ݡ��˫S����NQ�B,�����wR>�*e�M�ד�Y�
z�q�)qEg�l`�8i�	����l���Ĩ��-I�"��}��/�'A��-���7{.w�3�S"�'r���� � 3]��=���.��&��Z�fȌ��m����X'p��w�}�/�H�L4�ALr25��7~}�X�u	۽�b��C���yw���ܳ�7������`�x��%B��������nZU�E�49�����ef�nB�G�n���Wݎc�����$�mk<��ߠpΦ&������o4� �H��=� mYXE�����Uh8o2X��R���: `�b�$UQBz?�+S@�x�� �ԿZC�:�B���"�`�%]��-rK���1��c��.䏶?AM� ��;��֞n&>�yM&��U%��� �$8�r�͈��Zo���Ouzv���)� ���f�o��Ho��đu�ɜ��<�t�;��e|15�pG���]�
cGJs�`s�2.��v`�̜D�=��L�tl�|�,^/�ȭ�ۄ^}�H����%lf�'eq��z�L�!����v����N�|~�a`^tz�D��v�iJ���P�raBʛ�i�0�@�`����_c�"��R��)�k�}c%^D���]�3�&�c|�������ݺw��6�CiA�$�SQs2f{���I�[0Rl�QF}��,#��K��`Ro]K���y�F�A����o/��Qϟ V����F-�s����8�X-��Ƅ��'t�=H���gŽ=�����bN5p[�kJ�{��q�a1����O���4p!h�̙�sI��$�T�%�����@{��0i��go�݇5�u�)�&0�=�q
�1��
(��CךsI�9��mK�Q9.f,�7pY2���C+�67�1�6rW$�����{���M�3i�\b�e(�Fy�J�2�_T�"퓶["^"��!a�#X}����*#�-&��.�0��w �Km��VӚkߋ92r�*dR,s�|�"�×�P��.kˋE2=�nD�3T��&~L����P.H�|���34��l�v�4_h�I�)pUjtE�=DT<�*R��*�cEU{M(���Q^BvB��|��	r�z ��殁=M�kh?Y�u�3��� C����vr�&߾u�`~0�E_U�l[����*��@�Ɍ�	��&*����G���i~._J�M��2UИ_�8IQd �Ԅ�G�]��
��ttoݓD7<���s3����W��UO|�M�4�`����Q�G�׋b
Sp���>���&��\���^*�Ֆ��T�>��!�]OeJ����;ƐZU�5�V�Q���m����U��p���$��A�N�
��,Ey��ݣ-�BM���
s"����U��.���^�T,אbG��[��j�8逛��q��y��i�w�e�ߺ:��
'��"n`�������b���h뽖�ZN݂����tR�7S]�������c+/|V�|�ݬs�}[{���0V?Xxw6	��N&LAd�v�s�h�_�<��7��~?R_'��>�K���g�c(Ά��%3�{\�`MN%��2��{>;��Qۢ��f[�J�<�X�3r�|S�p���pS�o����:�,/W�2{&{�ﵲ�l��}���h��uA�'���HX����g��a<J'�Kg>[��oّ��{d�L���ɿ���S�lK�&��5^N�_S�a]��$�$�ބ�ϓDfL�=��Z�{R��!������ޢY�2)�N^��z�<,b�t��6O)��RY�U@���6)�Kk6�3������x�YlS�M���s�xcu�
0+똽"Ly�i�ݗ�{�UE�*������u�f�$߄�	q��s�p
�����Hj�֠�����'҇���cF�qX��D�Ӊ�2ǃ-o�)�}N)���7��������J��W��!!��ͽ��@&�!vB��i}�k7I�
,�����p��:; ��?RP!�ib���5�=�di��:�Z�r��0[h�A��8��:���V�+5ؐU����F��\xo-�4��l�0 ��p�fŋo�$��kq{���K�ad���Β���D]$F�a��4�ZL�T�Wm�38�1+6�d��(&F6��?�0>vTQ9�n�Or���p���:����~�r*�oq��R�R2��p��ݔ?Y�۸9_ ^eq�T	�k[�9�IBp"�M����)��g7�zF��G��~�:�����n: ����:P�tX�9+u��P;_��m���_�O�lk���;��VJp6����Rh���	f��~a�<�gԐ;�ќ9_.��?��z�p��9Lo.�~������L��)I�<�s�O��>:�8/̇h=g5�1���T����x��)ݓ;[ʣpj�@����U[�Z�'�ю�y�����л���8���lGX�}����z�o p?���bLg���Oٺ5C����j�"��W<�3y�;�m�fD�;FB*
1�W2vy��Uo�Yz���-�+�V�|�4K#ja,	^��d� ���rĘn�^�d�2�GdJ�N{�;DyļCI3ں�ܟ�u��	�e�<���Lc�S#�tcxJ�Qg�y)N �O��j0�zeq��PnVǛ-�H��q/���Nκ����6�P���|n	��B���+~��
���t�@ZHt����[������0�(���jx�;��̕І���!�R��d��I��u�7k�-��O��@�A2�k�~��#(�i�P�ŤVQ��8�[y��� �s���M�эc�I7��K��RA��a\�~��d�R� �Vs�1hs��G��C�K 1F�Έ7�a&)ʸ����F�P����|i%�Te�}�(�_p�=�b�����}6����l/��q< s���ƾr� Y�y���!c�8%�#��c��C��d8�O����^����9�
�Y����-�9�*7��<�DH������df���'�e�n��$�?�R��9*s�K��8w�簍��bU�F�m{ؼ�C�(Aw���8�V��Z��s��d���V����%!%S;���?�I�Ψ �|� �`ѬI/�O�q,��Q�p�\�$?��x/Dԣ$��uPY0N�xt)�ԕ8��e�8O�g����=��B}������U��/�"3XؤhHJ='���0��n�4� �N��+,�Į..a��,����i�XD���������g��7��6O��H��r�
��|g��ȄIY���G��1=�P�OX�)��gݭ6\,\�X$�>\`J���f}��Z���T����X�i3'�Pb� ����g�Wq��ƭ�c��;�����p�
�qlH�+��K6�~*�}�iX��xuuAA�"k��r�υ��=?�zz������b����!�ƃi�G	�ᾎEB+��~¥�X��������qb�j<dݖP� ���U f͢�ɫ)~�6�ע��<5�|21gE�l�M>��߭����?[.��-0��'����pg���p������O�86DA� �*?�
�=V=�/��ʮ��.:<�_;	��������?��5c{G�6�¡�Ϙ!��$]���O=:.4<*ʞ#�%J*��ԅ%������Z;�S��z����4��Y�.ӄn�\��I�g�]%e�$���)�&b��*�Ky��X~~8h̽3i�x.o��9�40c��<�A�@�Q##KN�'�F#;�1X�/\O�-�D� z�̗Q�m3ҝ`�����|:[��AW#�2C��dص���|���}_�/هN�����C��[�D�����Ộ��v;�`����*�]v�R.eXKb�m�;N���[��i�u�4�@9cHg��|�1z�I�z$G���y���-�[�W�t�@p��(,<�z pkAh�͋t5L"�/�����V5��b����X��}�b�#��D��Ü\�}���@ɕ*b��_��?X�ȯ
M�*9��Us7��;:C���K�v�~U��Q����0(4��<�8򺎇��-�k�_N�X�l��x����i��J���O0[�v��p���Ee�f|Җ�vi�q�?�8��ID�=~R��@�l����7��ٛfG��_�'c?5�M|������E;����,���I�Y7ױL�x�(^m&s�!�l��KP�
��Ҝ
� ��V��!�E-�j�˷i�JЬz�~�!9�x��*�����Y"��1��0�u*�w.�1� ��i���`��o�HV_]�(��13���s(�dF�9T�L�������k ��u�@qX��^_%���%s,6���#b��f�K�H>T��+9��}df��n�f���+"6tn��������؁�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�P�)Bs|m�dWc5j�C`�wJ��
�A��Z��Q�X"{E� *�Q��T{x#�*���w2 ��;�3qF��[?��s$T3h<p�B�SilEpxF�
gi�� 1҈8u��@�a[h$J�Y�ѿ.E)T'⇏�N��O	&��$��G5]z �q0�Cj1���e��U.!�S�US��G���� �ӊvl�%oXCL�c9l��6�	/Ĥ��#���A�~���%��M�O}��x�c�Q_ު}Y����Ie���/fѴ�~���B� Ke�n�P��/�Y�^\"c���L��vI� G4��eG�O��4@듛+WNo����9Nމ.�4t��0���� ���P=�fa��ATDA�e+u�Ҡ�Bةj��Ik�Z���P�b֎�Fk+*��K��\������'xa����W�O_0�W�Adz��k�z�q8f�ʖ��tz�t���Qd�C��	~X���(@�a��z�L�kE�n[�P�\�9����K'5�g`�8(�B���
F�F��|��)r�ד��2[�����%&al,���0�*%�d5��Z����Hk?M�q
�3Aҟ��Uf���>G^��Cg�S���9�ݳD4G^E�9ݠb-J�uU���hD����B�Rt��C>���g���~.롄C�'&ov$�WN�⪂1��1�4h���~�t�L�i���~�Qv�?��U����+e�I,�U��m����7�{�Mf��!ˢ�(v!ɤ�m�Ѡ.J�j�0�)�=9jr{�\�֟��m���A7�ԛb �A��� �Tw��w4�����:r]��U`��KH�	��ʅx�_���z��o�2�$Seo�t�����ƛ�fl�r����n����/����<�˂0��Z\+K�vhxc�P͟K�4!C�ʄ���A�&����V&�N�����G|VN�<���XyEM%'S��%���+��(V@*|�KߗI�T@̓�f��ڵ�b��V0�@���"�u���dP�3��˫"��d��g�&����=Y�*lJ$6��[��Siu ��BRT��e�����/D�q5�����e�+ے`.l�K�����)L�R��\�.D�$�$�Ag6C�����k�D��R -��G1� p0���1��;1w'=lr�Z�x"C�c(�����Wga�����a������ �W��dB��,��@��ހj+�hp���4X[N@Z�a��H?
yX�D�d��}˓}�o١�ߖ.���w�k�o�S�!jޙ�WT�<�ؿhR:���m�h���nL����P���XG�>Ai�z�|s�E������V-��!���|�0�ٌ��։��-�9M�{�\L{䞦�b3^��*/�F�A�8�Z���vK���m������X~Ljko�WvALφ��Dm�ݐ<��8Ōrw�@���:�Ý7��'%��í�O��1S_���z�N? ���@��z%�&�)�����_���8���*�7�څ�\.��*��Q�mI�q*K?)4�T}�`d�E��Me��˨�������E�.��ooRe��pHK��c�`���_V�n$X���?td�޷WJ��o
�ǁ�����M�:=<����h��L�U�w�q�U��+9@���f(��|QN;t���!�]�a��`�Y��弁� b���n�B���@*�Q��[F<��\�]? ��>r�M���l�x����N�3dJ��Y��vS�s�#Rп8o@�x�+�r�A�4���F���<��6'��T코p��cH�����7]��V�'����.�� a"�͜�@�Z]�W/��w��o�[��9&���-��u�}���жNѢ8�i9�R����h���!�B��r�ߤ�$Q�Rs@g��?�������%��NțШ�dj���;@�5=���w�k���OX\���`�A8OpH����W^X�8;tڬLy�SN��T������N&3��w��*#�RE�]V�q=��i�
1p�K+zZ\+��j�@n�l�j	�	���ί���F�J/�F��W�9X���_M#���������� 1�u��&�&Þ*s�6�L���9!�y��fI}��Gq���=fL�T���r��0���ԏ��s���#
v'9�oI�P/H����Y%��J%��Ն^s���l�aNT{VW�شb�:���r��^�!��Q�P��Ԉ\�t�܃���Т��^�0`��r��]6W�z���C3���4�Rla�ڬ�`T���O�}�d�'a������
��̿�F�Ax��7���)��C���o�ZO�w���阞5�%C��)���	�M��bW4q���T�?�ߧ	~�.ߨ������.�`�kX;I�9�a�V:���r���QH�{�{Ģ�Tn]}'��6�����c�L<����"� ��IQuO�4�;��i�R`��s�LHf�����BF��"������ϗ��ݫ�w˜�ݹ��0�|T6�W�g�+菜ly4� �{��R��՛� ���n/|$ء̃�Vxt�{�V�y~m{��������d��l`&�e�k?P?\�U�M�$�*M��%ٳ9E2��O<80����ˆ��Rva�>���|1�G�Dk��ф%��.1SAy`�罼͊9Cf�Ӛ�*�otQ��.=���P���nX�c���\��"_����W��hH��3Y�G���ɽ�Q��ן >0gAI|R	�i��Duz)a�����|$��W��hxT����h��f����IS��?<�+i�C"�B����W	��*���X�U�)��;�l�z�ׄ�%V�dOB��>�F�����L
sNa�S$xQX�x�ue?�C�V�nhu,m�Z�����i e���;�i(��k+�Jj ��Yn�=,R��3˾�bT��r��.�JёW�B�8�A���
z�Ý���Gw�������o���C+9K���]-.�&�+�AgЮ�%�7��]��3������m�ף�C�u   ����?�#��^�.p[PY(���b�(kiϞg>�
��yF`S�0՘���@�W&���6S�Q�����D����X�u�@EY�۸��Χ�kB�T��bf��>��CبUñ�muh�"`�E��W��:G�����[����&�e�c��t��X�F���?X��}��Pަ�?������rr���ZhX>2,���^-�� ��|��/>L�%�Y�ʨSU�$K����(3C�NI�W�U�
��H�W�R������q5�u;�]}1�uՂP�wa��	vq.�!e�vz�F*�q�Ze�؀�~�%���\�EccU����Cg�*�ܛ�ܫ�@{w��s~N�)A`%�Z��}t"e} 3��<?f�G[�
�=D��<��"=�"�wr��:�Y&8�%�8�oL���TBQ/m�,��'P�	Ip�f�{,����	��N`��,���K���)n�X��ď�!�m�b���m��R��Pp���K�o�IU�<Zcγf�\�,|�[a$�����c0���  2��P�՚�Ϭ�����Ɠ����Ty�]��#!�L�=��.��|�MFی����d��X��ߛ���C<�)0� [uf��tlh"O��(o�սj�J��l)�&U� 4xÉX��+��3ʥ����C)h4�a���ы�����	�V�[�@�U�6e�������Tb���s���so"��p[���L�
&oM�v�]�j2�PċMh��qZA;��<�v���b:�u���e��9'qt����y~k`��uw��l�YO�R�=ֆk���=�H�D�Ǵ8w�\��rF��R��-�^>��߯�Y�p�	�b<F�%@������4R���wcIk�,�k$fNNz��:�n�5*�H9D]�]J�=��A�,��@��#�ӯ�=4��w_��90H������kk�4Op�����7��>���燜��ۈ�*�?�H������ٮῄR3�Q��<�.!ix�����65�`�=�� ��+�H�[I���G�K{$�g*�S�����˰̹]���4	v[�M�t����O�k�k,Hj	Ͼm]��	|h
I&Y�l�<)0�?��H���&��pE�*LK��Lp�9�Ģ�'��D$K2������oW�O��pp�	)z�����mf��A�d�R��;�Z>�dm!c!� ]�/�Ea�+FI �X]v-Oj���g4�e�����<FX<3��Ѕ�S�)<�mk�\jB.�!��ΥX�<٧
�1��1N�B�� �}�L����^j�@k�q.���"��x�֨Nn>�Λ�/�7=�"��I q_<���N�%��%�-�f ���ޘ�q�/$�|��r#��a
E�E4����(��}-O�������׺t��<h��Ȅ�X)Z%6�<��_�.��P�S�M�!���s?���wC!OP,�>�=2�n�^���HI�{��[�|�Niv��)q��Ŕ]��$�B�w;^��VI�顪���O��<�Qē2<���N�p�����r�.����K�����VH���ص��D�.P,�Ǯ���3xsm���	�9�\�rc�!w�*�i'�(7�K:�T��8��ѿn��Ci*��cL��jG��ƀo9F�h&^7	n�s�GY;�E<��^�����Oe�;2��,�7��7�U����Pu��mw+�,��Hk T��5�vǗ� �h�����D^���GƢ��������$�OLc�Eoy��C_*(5�A���> �s���W�[�S�%1j���%s�N�f-��ʝs�������� ���M��g���>�M���j�\�(�Pѩ�w�۠�M�;r!�m��i��7�!г,�,�7��wڂ؂l _���c�W�P����jΰf׭V�]V�v�����!5ۤk}|�r*�L�V��ܱ�o��M�M#%&~d�����'I���t6qR���T���4Т���ݻ�����ϭz�zz���Y�v*��Tש�]�Q�����Ce�k)�P��KH���� �X��!���)w�8ɿ���������m��>'�+�_k�S��<\db��
����Ky[�(e�K\mqt�(̯��d�=�X$lG
�_���o"�,%Q{�?lg9��(ॊ������pu�6u���$�t��ͪ>rX2�on�X�7���hp��C���}ή�y���U*B��h����ZI�J��)���޼}@L�6+*L��؎�{+-�O��q��_qk�sȎ��TXm5Y_6~n�����`�c}��/7_����}g��Q����5=���V��L
N}ݺxa�݃��Y��_Ҡ����Ssf1���~��j�3��4� �,�Qiۂ���y��Mfɹω)?!!�=J-PF{�,̬��c���;��2Eh�-�M�S�[^�fn�,����P��"��L�V^�Q�=<m�~����y��n�V�K��^t�FbTj�=Iho�n���0�SP�úW���7Yʜ�}�HP}�^�x�s�Wn_^apY���+9�O���c蹫=�g�$��<ST`��
�.�A'z��)d�����*�����b������)�f?��c��N�JŔ��v��HZ��;�<�R������*�����Ir��1d[A2�4�IO��$���5�<32�K ��	׼���{��h�+v��H>�|�Nؽ���O�t{��x̣��6�`�Ь���j$��Q_�+P�X���ٜ�>�-���g�����ҹ���J� Ь��f��b��V�l�R|8��nh�L<6��n �_��y�A`�n���WB���_�&Nˬ�����Ҡ*]�k�Ǡ�EWA!#� $���~6I�1j��y9`Q�y�f�='� }���a�I��^��AE$�4�ꔓ�b'����c`�IؗfQ�:cGut�������*�.�14�S�K�M���@Tv��w*�7�a}�~�\�k�+G�l}؎���+hB�_Q�	�b�5��=�d��o��']]��)Z�M���x1�uu�@���<�c}bwu2�	
8S��
���?X��`	4���s�g�;�C#�&8_{[uo����e�T	-�=�G����Y��Z���_�/Mb"�����"6  �,Xo�����re4GY���s}�fk _jT_|C^Dn�ځ. ���2��*����e�t���T,��SMz���]1�j��f���Ij��w�m4-�gew�����P:���������Ro���%�d�b���m��p�C+yjZ�03dC��#��-GyV�_����H��-CB�3�#��*%�}J���A_\
봹�=3tkV��k�qb..���fz�س�Ҁ�'��n�7�K��F-76L]��/Q|n�!��%�6� ��8����h�=d�����1bd�>�Q�*����R?��<oX�v.�/F�[�P)Tj�O�g���4n�dG��4�%�M4j��A5��8}B���+����
�ʫ�����i�{�q�r�ys��ׯ7z�}(,�2�Կ���G� �"Y�Og.�n\F�������0�>�����[!�G��P���dF�~ �d�y|�)�=�ٱI��՚TU7�hI�,�bpXY5n�"	�ĵ,�Z�p���7uB��:���^r�Y�\\�N�`�<;��{����Ifɪ<���] {:Yl9O��W��d�Gqoq�4 8���D�w^E)V�Ҍ~��oi+>SY�~lA=��A۠��#�!2��b0Z�_���S����T�~fCn|溥�iwO�e�j�9�w�k�A~��:�XQ�ӕ�$��+Y}(+ϧ���Zy�o̨l�)��'������`zn��6{�5���}5Ҥ�����w+
���u�{�&X%j�<�v>���$����v����b��E�em��eé�婞5��G]��+�GV?�ub�N��������h7�I���@�T�0������N$c]���$!s��B��j�M~?�lG~���k&mN������	��]�9u�y'�i�Nœ`����aω�vb�7��&�B���`x	�qS�sC��VqI��q�"0#��f�VoO+��978��Y�����_�����C���0�QF^G�l��`e=�Nb�O��6�9H�,��@���
�I3�nOp�}��
P�Ǖ�r�`�ë�_7HM��^	"����M��4�-4��M��:������H�'�C��a��f���F����(�U���z��"j6�_�nq*�i,�g2x\Γc�h�i$c��E���o#<TӶ�8�f0	������z��=�YZ�y�gb �r�.�01;����%gfH�b�=ck;F���9UED�=M>�QsTef�<Gj���V�hW�P��_�zo��q4(GR��]X�F���d�p�9�m�r�؄t# �����g6�Y��Q�F��ʰ���0 h��]��+zIB���1av�+�u��h���J���c]<���F%�n� ڑ�΁	 	X4����q��j�b�p��<���}��ݽo�Gƴ��3 �����[Y��'�s�t y{��з�v}@5B�bg6R�P��汯&y���wI�`�CzN���v��[_@H�O����a�����A�Kx��k���οCz
kd�Y&K� Y�Ч�Cf��DTwN�F��g-�Ζ$�<!��v�iX7�2��ڍ���?�p��>�Q�;(�{�Ǩ�BbY�yVo�Q��6�d^p!���/:g�Na1�O�|�q��E�JV_i�J��*d<'�Lg�ݖk��b
C�~�$���$�%)K��p��h��?lJ(�4,ieMg��ˎ�%#X���A�U�7'M��r�n
2�ׅ�o�e���VQ�ۉ�jFrf���F�EL���u�"	���U��Sk���l�z敹�Ag�ܱ�.�`�8��?��	�c�Qm@s?@���XX�';����Е�I��n/|J����ڽ����;�}���-�f2����H�siR_�z׼����9_��j3�g��Z��S6��e���*N��p���c`����H,�-�K�@�d/!Dgl|�' :�7��,N&�n�[���
�~�5�ܠݢ@���0�)�dLuI��b0��2�ݕ���{oL��F����>�\�[����lDU�w�Ư����!�2)��`��9� �x��6j���r#��h$󸋋���}��:�>���qQƱ�~�L�X���{���L�W��raNk���&�=~k�_G�z'��G��v���%��v��U$�(]���C�<���| �.�?���$�e�b�j�Y�h����SP
Q�K�&=D���%�{_
�7ʄ��Hor:�]V���)Fvk�z�	��R���/����܊3��uR�Gǟm��H�i
�tq�%�џ�����9v���5����ɗ�՝�[־�0泒 P���b�]Ӌڂ覟���yR���&y�x�*����R�bv@�@&��ǪS 3I�L�s{�C�c�[�!�U�㈇orBcԌ_?�^��V��61��D�?�p�ʜ>�qO(4�=��j3�u�:��d�0*���>����]�+;�ݺ��,���V!Z����hh߲�l�h���d���%�{y����k��(/\ǡD�R�$�D������KWIy�7���66�6#��~m���Zqc]he�6h��,/5{E���oz:��&\ض59�FU�sj�@����3D�=-t�GT����f�EOd �Jj2cF��p� [�hz�ϗ6eݘc�.���D�����=vŠ�mQ�,�J˅}=֍X�j���j��A�u��R9�G�I�-�� >C�:� �'P�Ɣ��_��9���+�t�}�M.�![����j4��\���+�3�����jq�׿;�����!��2�[CTP�����KTG?bef�܀���p�(�P�v�h6)��-���^~��F��pR�t�K�3ȃ�.���o��K��r6�UjX֛S�ѕ�	��1;a�r��0!�ŵ��m3$�����غ����$��� ԛ�Ӹ�����<ɷ�L�c��!�yk��Y���C_��e����/�>�Ӣ`C�g�Ʃ-���#���Y*����G�ESOw|$���Fgwu{�ZI+ǙV��4g��i��ֻ�_�/`5�U���i*kWe����~���7�7~!67$5�~~;����v�}6�{����IŴ�!+<6('��}��#(%R#,�y�=�)�9Ͼ��߰��m���������U3g=�8���M/�!)������U'Su8�=�)������'�5�Ջ]G9������H?'���?�o�-��sƪ�|Q��P�+ɴK3h�)�W�yL3^�4�#SCSA�p���XdqE�q��m��v�V��3�G���u@E�Z�LX��R�T�Z�0�¡C�8Ȕƶ�����Q��
��uǧ�!�Đ�#8<�V�Kr���Ջ*AcبB ����	�ٜ���h�p�@�>�Qk��FE�U|(R����L�wec9GlMi����A��kb�q�Phy��_<��qH�Buyi�`���j����ߘ��w* �M��W[J?��9p�c�V�?_�{�I˧m��1�+8���ʌ�Ho���,,��I!x��`f���qc�H(�js�"�&��RєlP.qǚS*3��	(H��[�YD�ʾ~�,�DzP9��?e�����/���>�~N���]���gωL�N4���س��zk�����?X�uH�yJϐ��V�1�7P�ܡl��L�ျ�{1�qE%�_xc.�q?Bu�Dбy�S\H7�Tx���<�f%���^xO�w-V���M���|�h�x��=��:���ԁ��
������S�	?M�/j[s"˱�G*�O��R����{�ý�&Ocyv�7�o�6�`�J�<���E��\��2�KB�����h�I���0;�)b1U}���]JE�,���������h�aG�j��R���11��W�.O�+R_I,J�(��m}�(����{�V��Lf]QH7 ��FKM��Ղ��m
)�͠����SF<J����B�3I�pN�G&��-��W ��FP��h�;��P����=I�U��2�"n�k���Y��1�zdqG��8�R���Z���eX)�^��z(_z���`�6�H��E�vѨ|�.����#��cm��\�h� Tz��`�;X��oS�C}"=sz6��>y�,gk��Y���w='�6�kۊ��Y�=w�-W~ܠ�����9�t�Q��R^�X^)��[��c]~��5����·�>!QK���H�AbB����E$�M�Dh�BH
�H��Oa7���S����RK���v`���y�`��z���0w�S�l���#'i`�9;�N��3���`� z'L
�� ��M�Hk�?�f@�H�"
��`+�a�V��=�./��&A����\�M��dBpWp[H,[	.�MT�W��IH�OB^�y�iZ�1l'4�\���*�M%�>���� @|�9�9��w�{xѳ�BD�q0�y���³�X�%>F# �z�{��V�P� ����~�Br�v3/�L҆�xJ�GO�E�1��d""�'� �N���W�� ��z��~G�����ݹ���kN��C��ui�����9���5\z���p�D�1�r�Ӣ&�t�t����S�͓����r� M2ݟ!!Ϸ;� J��;�#w_���Q���z����
Oi{����:���Ϯ�������n_�a�iCM#CX��' ڶ�!<�*]I�t,0{�N˪��M^��@�P8\�](�D��c��DRؓ�����@X2A��P�zii/���Yh]NZ:6Y��wF�n��\K�I@��b=Իf��n�Ђ�ș�U�K��\�n�l�Jf�a�8��gn=���X�Q�w_8G*j��7�������4���
l(��н�Z���d.�%�!�a�f��y�%���sBl���ވ̈�*�$�����~rh0�����k4��Z���%I��=߄��o{�C�B����ٖw3�7�Ml��s/N-�L��-lҪ�e^X)���I����5�3��T�[k��lϡ�9J�K 6�����9����$T
���������|���5�s�B����pZ}�3^�zk�UN��\��6�pk塚W��cdM��-F'}J 5��4$����֏�-3��l]��\@@�ˡHX��0�߶�ŷ��s�bj<�0�is�����J�T7]NL�{-w��������{<�*��+�̊qu�Y����R��8j��[<k���wz��R��f�m� #a/�'F=N�7�)�̑ڭ�HxŇsw�����<^�6�N��<I/.p�� JPT�}�H����t�>b����ls��L?�PL�֯Tc�f�G�=�� _��d�
dR,�Q�Ow�S�x�,�O�e�z�Q�\K\#�� �P1�@���X�!�X$����*�b!�$�׵Z>�F�r�CwF���D���~ᝦ9�p5�j��F$a�3�&Im�Z�'��i㠖�4p#e�!��ց��᯳��t�����b@��˝@��gߙ�
�������&��a�m#��ߵM�'��7=�Wr�ﲰfE��t��<6�)xM=��ӽi����L��=�,J��@� �H9L{��ԇ��٢�����J���;֥є4��gq[�=�N��C	Y��&Vs�nəkt^�\�O�`�R$�&�)UH�g2��u�m��J�B��js}IF��%�Li��X�%E�p�m������i�v�
��e$��Ŵ�y0KUu�~�-��#�<7�U�����n�b�[�@r��_���j�:�����3�A��B%�p�\�?ה�7�6�%�<�{q����p�U���8¢�L(Oo��	.4����#Nq���jĿz�������aRL%�%m��/V{�!"+9a����^1��ڕ鮴��f5��\���Q�����%�Y�����z�z���u�32���|mڅx�>���l2�ӥM���j�)F3�pvO�u{6����r��'?u�
kfp���\"@���G�	�~����/z�3�H7�r�S�+��c��(�(�J����O8��T�~C�Γ?��^��6{}��⶘��!�2b70v�*ϕBR�_,���2�Ixs�;�p�<��q������Zb�r��+�����V���_[���0�IN p�7�#|�>a ��5sڞ-/9�4f�����hT�6Ѝ�S0H����X',Jxac�Y�����\�a�8s�F�HZ����k��U�AX�.[��0��1�Q��Oo�_3�Ӧ6��X���4������H���RJ�T �Q�gA#�6����1�g���'���~>>�Q�fP4�lŝ�t�t���{����*�m3��:T�y�Š�OY�dՠ!�n/��Rs���3�CB/� �
�w�Ֆ���5��/������O�.e���i7u��[�;(TG�X�pi��wi�>���`����/5��n�*ԫ�:y���� Us����.8ӯ�-3����P1:4�������� ���;��0�O�Z�ى�����z��k<d�P�#��7|(]ؿ�;��G�D�j�a�4���`�}-�B2$�(�;�&�1_��!�d�\xI�iVIBў7�ݡк�	ew�A\s���@
�v�LE���H9}�����:�f�w��Y��B��T�#fm��m��8�C��bVz^Sl�O+kͨ��ZAtRk��; ��	�[o5o��U{ʃ*/*����1�iΘ�}�@��j��x�\r��n�N3Td���So���ǀ��\����#�v7�xk�Z���κZ�r��4.�Fx(Դ�4�w��qX3�I�Dn�*�l�v"º}��{��;��P*�oz�B����x�׶�z�����aK]�Db�ҕ���kKe$6f<��7�/p�\�w�w�9P%��7��H��(�E�k�j�^��6�хJ�=��'���^�=����M���]$A�l���c]�AH�|��Y��
�<�+��{�oދx G�8�X-�N���=���ŭ����tҳ�S�rX ��!~8=���e-p���q��b���~��&'���Thk6L�,���������h��l�����	��a��ߎb�Hb;�EQ���';�(��v $�06J���m�J�UP�Z	G1Q��m��q�&S1j?��}1�W��$k0	ʲ�d��o�]�?Q�w?Y���U � L�
4wJ�_>��G2x���$��&A�3�GH��M��(��	n����E�Txb���:���D�xT9��������m�6�w(`�"�"���w�a��2c����[�ha�����;/�P������gNN^%��V�J���&�X��Z����l(ܯ�譭���4zF���T�=E$*Ռw�ճ|��J��d�0L����lX}#{b���iLq�k.��X�W�����9�|7�����!9�ݨ���Gz��c�i^U���Rxl5�P�,юM�V-]�KU���#��^�Qi��3S#=���bek���D��U@9�D1/$�k�,@���q��{�-�ܻF��[�8�:J*Jw�se��H������0�E_��vZ�~6&���& s�{`zM�藘�йM*�Iz�h{N�I]	 !	,n�.ʎNq�)ოy7|g'.��{Ր{>-�e�?�ɡ����(F~��xǥW|�Ƿ2��uz(�W?����$��.��͢0��kQ�$�����������UL�F�>w�=�m�(m��;���W���y�.Q�ٵ.nQ��_��*,Ի��/�#�g��P�Z4l���k�Ƥ[��r������"i��_V;0b�6@�$+�m�ʇ1iI�M�lJH9C��q��4p�-�̡Sz�!o
J�F�i�XQYk־�6 ���)X���^ڧ�:`xX�s�<��<��ob�|+����m�j���B?w1�L@�������0q>eo��JӤ�[*�az"w���#��~}s=[�n�4�6� H?x��|��0
s�p�ݼ>��%,X�IX�H��X@6�[6l�Z@�	�!��4��M��f)��]�霘!�J���S:���K���g�많i��e%��馹iIF��#�Im�����:�t���&X�;�#��U�by�+IO�_�j1������:�r`yL3��[tx�]�iSqU�e�-@]�c?5[s�Xuʛ�+H�����ae����o�7���%���$3��t���<JD����@�] Lխ���eB�\�/�P�:�J����3�AU�R0`h�:�%���-����b����v�MS	^�qb�n%��M�|���\�W��g��`@i���R�_ $T��v�����P���_g؇��E��Ms����-���M*�%��D�aWkPj��K��:?,	���C�B�����T>�Ө��\��u�}�$�x�N��&n:�%ղ���ZS*xc�O#x�������"���c3�|N���+�+M�0a�
��iD~��`���r��r(՗��*��q����a�#�K�آ��q��m��xǹ�0��_o�?�m,�v[��"_8��s���mR+2wx32տ&���)��۟>v8L%�8��`(�&��xJWr��(���fW$ޠwxs`!�2�����0-�ޠm�r*n�E��O<��˝����%l�:*\Xxg��f���z56���K\V��[��u���u
/}#��Z8 0:U||�`cV�dMٴ/�v��������=����t�`�U�@]�OL�b��So����#�Ȝ��$�1�*᜚0X��
|x�/}'�Q�
W��Po���|�pG��[�K'�a���ݣ~z�^21���/P��ԗm�
�S��Z���q颪�:
M�����G��V��i��*���-Td�
.���?�}�%5��]�F�����d���"t$p��������rqv��N�ep�)�H�"<i[��5"b}_D5`J��f=�<�F��~-k��}�F�t�.��f��4���l+��a�>�2���'0��zݗ����	bI�p�,+6��������B�?�_o��a����9N�ǃ��"�R~u"]"��2���n`���� ���]B�\��7��x�x@��N��RlL!Yȝ�w��ٚ�@t���ñ�~#���.Ū|��Uy|��=�	���"u�relU�~4��#�y��4,og�֋�<w/� ������R���,���I,���6���T[vA鶡,�_�e7���<�8�ף�Ȑ���L��9��|ܖ�M(��1a8�Lt���p)EބO>�MM����=�T�KGG/_.i��S�����-��*ӂ��0F�>~�S��Z���0g�3Ǿ,�S�뮱��ʅ*��5d�g?y�*v�4*���d.s�d�70M	��/�|W.�F�D�o���~|�0�YČ89�f���:2;Qi ���O���>��ϩR\��l&f������(+1%0�e�O[�k���hs�Eo	��.U��b�*��ʀ32u�GY$i�?��ɟ/Ɯ���E�$4��*H�5ש��j�f�w{2�Y�g�PKӾ��8������U_x���4iw˩7���z�)�������ML���gDz�#�5�{Eڝ���x�9q[y�?�Cq��RV��)._�j�Nۧ�i�/i�֯��G��������!�ў w\?3�l�~2k��1^��8���0dS���K����`NW+��}6�t�v������Rsh��f)8HN-��[@u��[
�ù�]hE��LHrwl�e:FD�aVx]k��kԟ(��wuj�s����.��R�U�l�����xc�^ؙ%3=2Y26��.���t ���X���o�
�!w�#���DL���)-�ڝ즨��i�.C�z\�s�No?<z�V�Bh8��w��Q	 ���~��͗M$��_��6T����[bA���?��8�rˉ����2�O�V(H�%z����7As"3�[�u���o����{��,0��H�8 ]��g�͠I��A��h� 3�\��^�+9��w�a)��Έ�: �q��|�o�rIpD�(��2�$0RX���nf��XF�uA9GD*k�v�s0�A�w��m�Uק5�D�1A�rCGڽ�b�-L��9|�4�(a�g��jQ4� ����9ԳTZ <r��?n*Z��xSL}P;8N,���Mۂe�<������<��e|����,�4�NI8lIU����h�T�R���=�W�=�쭝;�����P|"�h���f��1_� ���ʼF��ˈ��(@��t.ٕ�=ŸQ�8,�`������t�Xr=ē�ۂ�f�b+���m�D����8�ז�`�[Y6�.�#`RHA1;��7�ٱN�nz��l��H\���j|R�dR��y?0���ɿw�D�R3��+Lh�l�n�{
�چ$8f�ǚ[UO۱d�
�b�Ѹ�ae��A����រ	���������S�� ���4!!M֭����/�R?q�|�0Y�c�&�܄x���y�V����uy��-�����_�1�l@,�<K�}}�j���yJ��f�B7�;��dS���Z�ÒPA]�׾Ʒw1U�3��^��>Y1wɤ��@��	E�"C{�o�@���@����H�iGj�יSE����������J#P&�@L��<�:��U,��b�#��Pxt'G��i"�$�J�m	g����9�2q���%��\]�B^��Ŧ`��3�e��á�s*KT��k3{���g�3��Α��L���-�?&�`��mJ"���4I�%���1+���צ��m��lܠ���tx��]�3�S|˱�4,䇗�k8�RJ�R� ��o\���f� ;X��ٮp+Yu�,�v�U�"J)�%�®��Y�U˅��1���ؓ5[�=���7�����50*3�r�r\�D5�Aӳ�@�F��Ŵ��+o��Aԯ���Lq�:�.|�@\�_$���is��O}�^��Rlz7�L�����"��&��%�M���3��f��%\�K}�$�kxGT����n�T@y|��p���ȅ�����M�}�x�{a�T�ǎd� H7�j�>�?�������m�V��0�E~�x-��p���V`��H� dц��m�Qx[TC�a����חêE[�R�:P���Ǵ��:��ՙ���c`(�&�s�म���� ���w�5�,?�I!�[��t� �ehD
8����zm��`AF��-#,��j<�O͟���}6�)H��:�Tvb�� 9��Ї\�F��#����>L7@"�5���ǹ��9q��JT�G��MU�l��'B>F����L��@�NVkZ�Aj/�َ�x��O^��������Y�F���bS�ҵvDiTr^%��l��ŌTNE8ru�,���*yͨ9�b�iK��J��r�_���&��P�?��oG^Ŷ���R�@�Fv���6e׵@"픾;��x0OSP*�1_��G����v���كu�c���y�\��OO.8��x6�P~��|���j��5�#��	�o&�$�6uډ����w"/�=��k/�Z�=�G6��K��ޜ�g���'���<s{�K��.��/Tˤ;h�c�ʈ�-4} I45��?���A���MU+D�<zӆ8+&^���%=F 5y
�#����`
Ȟr�w� -2���S����m� ?� ٬H��C��3O�e�޻#�ޞ�U5����R�����it]{��W�'KiZ(,�
n���=67�/�*�T�BM�W5�r��1>do~C>�8���<힤"�n���(;9M%�@���q�Pu�jMEȊZ@rTDY�5o��B\�4�]�*Ղ`�D���޷E]�A�D�54P�✩�!��Ad+��s�����_�.�@L���o�I4�"�*�\3=�uXJøh�3oU�H+gK�X�.�Q�����@3u���*�w4x��o��-P����lŊ��8ϯ6�J�Ir�=�gUys<+L)٣:9푃~�'8�G��}z�!�.�����`�Ǥ����,���
�ƕC��0z�dO��g
�I㨀�O��1̽�)�+'�˻���l3?���ac�+�We�G��W�f{3]�ĕa����d\;��6���ȏQ��o�D�|K����B�?��*ou�#��و�$z�\'��pK��P$�,n���%�k ��8�8�9Gz���(�����SH�I�<G�.á���W�fΆwb`��X�/#���0��!�OTC���~���	f9����sS{o�,Y.���O�G�����b.���'z��݄j���<��惒�����>�����
��M�5�~�,�'Sc�h�}U7F򖰛��б.�+O�yB�X�
[@��@ϣL��-ZG�z��<��\Rh��x�QT9�N�����Kc�ES.+c{A.�՗2бB|'�#��N#粱��$I�[�]H�K櫖�3d��v��� �XZ�9�@����zw�D�tX7��[�����C܂���%�tW��)O����ɖ��8<��yG��Й��.B�s�������Ǯuو�ĵ"�#�N��~��F
%V �%�D��ڔw[H��f!W�Ty�V\m��"ҟ�� �%?o�~z���B��>�u����U!}��ત���/���mԾ^҄��p���������֞�y5Ǫ�wG����$]A^������� �#
z�"д�ǫ��,�4�<}�*�����S��I��H[���|�c��_ǫ��D��`6�w�>�7R�Ty�rb�o���~���� ����'g�3���\;-""��-& n!�|#��m�bj�P���z��0[WϨ����?�}WI{G���9���pQ������ _#�������sk�n?����¿�Z�=Y�+#�*�4�������8�Z{t2�u���8�V�uf3}�<t���is�`�����@W>��rr�pb��`��ܧYM���_;s��0��	K�N᠉_����#(��eIq�&�ƃPp��-s��0�@?�8$�.���"O@s{y����q���Z�����X�~���\������ �oD�M�N�<C�O9\v]X��8
0�MHQ&R���� �,���p:W�/��䘨JnY;3qe[�7a\��c�:
c§'���>�
�w&m����s*O��2zܴ:e@�@��e;�|�B��S�t�+�x��]aX����U��J����$]n��o�"21�;�@^�8�%S^-��fȮ%*�&r�KzcW�5Y�i��޹4�Z�{~g;�\sf�}0g��
Η�Z7��|�5����պ׮oֲ
:���~݈�R��<�j�[F���߇�䁒;���Ē�s�u��3�~鋙��5I<��֋�!��Xo��
c���H��fWV�M�0~��Ar�.����&(�qVq,�)�s|�)�LXĳ^�?�o2�B(J)ϳ$���8�(�����D�
:�1l�������X��ǿ�����hj��ŭ�*{`��`�)N/{k~_hVp�v�OX%[�4b?�)��K�|WNW3������{�[��"Æ�z9����
�3��;��sg���`���~�Z���$�H$<��=�n�	�X��;J��
�����_����Q�])o������v� �J��A�i_sVa��TJ��D|i|b�������a����I�܎m��xE�Uی���,#�γ��')?Y�_���s�D�T?`�W�ģ���s!o�$����%Bk
t?Q���
IR��x@��Ə-�Ѿn!��۹�RFL�Y�>s8n��t��2��o>���}-vA&�����4�)�4����7k��Rk�?~�U�H9ۘN��\�#s�v�?�-�@L��C��� �@��4�"�av w��п����Xy/?n�	bx��U�*��:�T��0�r��~����%A�����\�4��&���
э
��K��v������<x�2Σ��ė�,uN��e����Kv����\����6pvz˂�m����z�����H#�p���yj�N��U(�D�^8<2�����<֙w���~_�b�A@��-J��6����Sl�\|�{�����?)i��)���^+���s��� v&��"���Y�pcY�'�\FR�8��|#��4jn���!�\�
)��5���~R��7��B��9����̙�3f�w�O�a�M	JR�L��&s��W�x��E�&�+�6~�D�	���>1�`�1�GS{nl��	z��T�b��b���t�\��=w\��'4:a�7����I1��ȸx�,�eh�h�+�{�A���z��k�{�p2�P��̟S\^�/U�:Ȭ�yyi7�@��D_-D�0X5K�̘�wYT��PU��(BF�x��-����4n�T�� �����/�73�#�Uo|0�E�{�x��ֿV���Y��c�Ͱ��m��+,�I�T�#)/�6��пU�:�J(6\B�M��y��d-����ac�X�v���A/܋�4%��r9[��u��D���8Nw�WB���c��FI�,��'|D�gx�`���bb�M�B�-�p��*�\��9I��?V���(�W�6��~�XE�/�7��������4�%^�	�8�=)VDՉ��nꗃ�����+�� �3�}NU�O�8�#a%�=��l����N������:��Ж��Y?��Q�[�B���CN�'��7+�V�c �lL�L�=P:���T�<�Q�[�[��[�d&9��=��
��B�ְ`k^L�6Wf!@�w�6a���m��Z0}E��e)'x���%��A�>�Y�F}�ן�5Ap��I��Qh����$�*�`�;�dg'�P�Оuru+o2�?7�^��lK]T�9���~�z3�I��G�^�{��"d�t�a� �!���k��2څ����s�r�A�M9�΋��r��$�s�
���9��Fv��ua���,em��qI� >,oc��7����EЛw�u_ߥ`�U=��_�C��,	}���z��U�
�]����7�3D0�Mw��@t�IfF_�t��a�A�(�,�|��͡�SP�ܗĩ3o� A����6DRD|wBj���¨`g1�q�l'���i�T��Bf�ԬaxCHz"�2E#�Ky��t岾mn��5���e&�?U:�s����%8cԠ�]5����l�c����գ�C.9�}7��&��ə�V�ZӃ)8vGo*����a���k�N���8y��DN�����yH�]��\-� ���]���u�gϵ��L�`[��z/� � \Q�P��&�Sc��S�R�`�@q����R�RĒ����x	��Rc�,`[�O$8��#p�w��09�ߪ�j�A|��|�-[̪EAQ�Ğ����}Bj�ikx�1>���`e`�f�B��u�,I��W�O|b���+����~��#�f|e�1�Z�9rY!���<�~��|N��d)ն����H�W��,q�{����n���3�b�Wu��*��OR�SN��m�o�*��	��J22p��)K�#�G ������Af&�-r_:�t�ܖ���:�� �4�\��$F����}/ɂ�[|��n9j�GИ�ᚻ������Z��:,fH��b]v��6����3�]'c�I�t֠2b���f�ӹ��=�2������%*d���cf��m0�PP�C%�3JK��2F���r|Tؗ��P�:�Pp�%}�TBR']ac�j���-5�h���DL{�&y*���VG(���;�KTW��C5l�u��6ڽ����R�]0:�>r���/��<���Ҳ�'��=����z��͓�YV�%WU���%�$b���@��M�j��t�k�W���+�3��k2B}ZM�w�^��K

��;pT��9��#�{�0��5��z��ĥ��6���i?���Pm�~]]<�XA�li��]�v�c��O[�F�}�N7�u��i؉5��#j���T^\��������}��S	.�<��w�t1S\�$�0�zb������j��_�H�������n��;痖�8Um�����jk���
�c7~���/����]�\��[(����\P� ��p�����*X.�� ��~L88���5Y�əΦ�i���
�ς�Ѹ~X"-v���%H���\���y�
I����X���t�\j����@�2^����[$('+��v��u%�+�6h/^D;�M����Y�H�̫���c�]�^j`���Ro��U,�؋}���kc�a� ����)�é��岛8D�zk����{���#�߆��YȎ��*:x�ܘV�u^2����{�'�\�U�i��N<Э���m�;�3�~J�ԌCN���e�"��
��M��At$�8ҵ�[�xS�Y�b���CJKr.`�Y�g'g�?�����eY�����~&��|�� �~���� ^������1����k�eಌ3]��v�asM�p��T�x�%U[\4>�����j��P$s�J#��M�ϭ]�X]��0P��.X�bv{�=ס��T��,.�t�V�E'�R~m���v1:�`�
�����Mh�*8}���N��D���2��kf�� @ľ�K[�y�������x���`{�@�T#����%���o��o�*G�!I��5鉮A����`q�>��)�L?�L��,��[���6�5�9�Uf~х؞�/�[�W�-|nJ��k~����K�8��f��JA���)p�����Q��;@���o�E_�Q�=|p�l�~���If4$鉃�^[���s�����[��]��(��h����[-�(��s=�y �:��g#���eLq�� �N峈5��[9��tn�ُK���`��J?:?q�{�T���нV�/�O8W���$<߅<#�ܬ����9r :z\�MM��tH�
(e�8��hg��P)�a^����G@�ۑ|�^j�U]S���Gz���R��T��H��ȡ����R8.FK��h�v�u%J*~�t� l�Η�S�yw���ekwWl�nk��(�@/���y�R,��\�b�I�=��ߢ�'���na-i����&9iU��V+��0r��
F"����D.� ]��;�h�Uyu0C^��Z7様p>��մo��G��~!�E�����o[V�[`i_��ht���~��W7e���c0<��t�e�y���j�k��ߴ�H�Xv�SW{�X�T�;���s�翼0s}􆓏�]�����Q�߹�歏�]���fSuʉ+����Yu�2d���f¶c�>.�g��oT`���x=rf�:a'��|8(v�HC��1�i��!����^��������S���%�B�md����s^``��b����	��j�ǻ���/.�Uy?���$?u���KeHWv��ڙ�<�N�&�#k<Ll��b�fʕ�/Eu��N�s��SNB#=���W�R��~���je���0_�	���PgM��J������}�����[�� �vƀ�ձ׳��Z�)�Z6�۾���3����K���"2���
��&wަ>M�l��ש�Y��U������B�kP�d�{E}r
���
<�����:"�^�G�B�Q��t����.oZ������^Rh�q�컉ƭG6�ȇ��cP��ُ���:��-!޶�,�|�w�60Z�|[��J;�C�N���r�"����1kv�����^�6r=�(2��B�O�>2j4/����c�/6�M���y��� ��N�Je���(E�5ˋ��k�m�c����e&� ����!�T�1�i�=���c?x$D�݉yp���NU�m-!&}���Qt���d�hn�]z5�gZ͜�9�mD�+�( l:n�������{�!*R���=�+ܝ�˛�RK���uBDtB�t�;v���$=B��J6���Ғ"��ta��~}�z���K���t举E�H�GNLt��*R:9i����`�g|�h�%jNWʯ3�7h��A��בߟ!~�V�p���!���=�D0���%��m	/i�������n�/8�͔1���Ye����N�ms	 *�1#������}o�{���
���ΰ�(p{��7����X۴6YE ����U��'ۃϣH	Юh�Xy�n�����ਐ�|[P�۳x1�ط���}հ�����OԒW@���O>����7��d�ӫ��{�ģ6��Q�*���-	��T�Z��ҁi�"��9E<=�ÚZOb�3/*�����r2�����:�?��x锵g�jlC�E�~�G�I��Ep�rM݉����>�W�AW�)K��$!�U�e���!x	����7'��-��XS)��%�v9�� �>����"1y&`���;n��*��Idi�|��0�"�
;>���׀��1�N�d��#��pl�g�߿�>�{_|+P���~�`Dт�*�Ǥ?�2v�^l����	+�џ�.sq�dG�w�M�AT�ݗ��gMM�Y���%ʢMkmĜ]��؃.�2F�]��z68WE��V�����F�y.����ֵ��]���j~X�����F�\l�r���{��K�"+�w����Z��H��P���S�?��p��!*��Ի���4�M�#vD��&�d���`2���H���U�,HE�T�Y�he���3\CSZ��&�$��%m����*Q}�m�P��a2�FS��{J��+9�v�tv����)f,$����� ���w�(\r3|ih�(J >�" _b8���U����������<똜Ƭ�8Qm��ٵ�<��c�+A���1���(&sQ_���٪�s@~-o�� �+h	���?c5:��	�lp�-N�u^e�F-';eY�I$�j̻�n(Uח���9ZiU��-f􃐊��<;�<�����8�0�;�����8�W+�03)�+�2���)���&��(�	�1nq�l�X�<Q�7cl���Ox�pbrB�+p�u�+��n��Pɖ#(�j�����>�+Ȣ�{u���2��@l.3�%LK�B[]~�C��H������r�vk�\^Ad.S��<�'��������c����E�D���EfK4�|�v�P!E���Y��.�]Ţ�[��G��c#��8�/������*����!q�VM�B� d:��u�nr8���e���"�C+7�����T*��O�6`��j0�7@���At�"�=.��n��at޳��u�K4>�X��2G�L�%�X!M��\9��&�����>ߘ����EƩ��uՔ��j�.��"���NH�f%d� ��y����}]�.��(�Q��v��gl����^ߛ��|ހ��v�����2V��r�gm���X
�\����p�|
�b�l0ҳ*+c�	v kPh��q�(�8,��$;_`��3�]�-$^������s�ռƩ�̗|
 ��9{A�OHm�)4�ޑQ�w��9�N�h�pnRk��t���I2X���=lߥ�(!XtU+�t�B�ҵ����WP�q�h��@5�\
P������J?������G�*,������:8*Jw����b�V�K��^�/��iw�t����"����V�����6��~��ſ��L4YfUz�%ʾݰF�Y���J�\ )Z��H�P��R�`����2?���`2�@P�8�43���XT	Z�|U}�AՒ���v��o-�>����l�|y�"��f�ԋd�� g`�^��43�(��� �$4�W(Z5�IV_�p�}�+��'��5lA�'BK�c5a�\�e�ȧ���r�
 �"�JH7G�K�=���EZ~�@(e���;���Mܺ҅�Q������qݥ�r��w��T< 1�ѐ��D˯�Q�����SOg�R@����~)���"S�hmR}�B^��B�-)��Z�Q�"�4�2����%t�������������=���Q~j����d{�@�'�8�ߐ�N�*��[7F�iLs.��c�7n����J���n��"������)0������4�`.C��B@�;�����,��O_��j���5������ܻ���uXB>Ja:��$�D�8�i�7�1d���3����w���Ѵ �z:���P�az��!���[CP����7c}kw������滽��0�qmB�՛������M:��qF�3�{��PM����gL�d�4���������i�CO`��gw��Y�=dh�Ä&��]���П2�}���ysr�hα�8�^��`%�����eY��N������]�/��c�x���7D�n��. ��7d3���_R��,@��L# Xӽ�D=��%�G �V�G<�Ǹh�t�����G8��PHOy^�N}�7k �0i;3xs\3�}q! ��Swg�ٵ>TC%>�*�%=�������z.e���Z�R���R5*x|�QIJԚ_���8�|���&M/�e�-��0Oa� �Y�MW'i��y�V�W#�F�P�����<c���h��7�)+�W�W�ݫ�M��P!`�ʒ׈�b�tq�m6�'�Ē���d����ʖ��+�8���q�)1�纚�8���I�9����*�Dn鉤J�٫�,hĜ+�k�
ۃbme�6Z��7�Wr�܌���}}c���4H�ܡ�#L��ޑ4"\�|�J _���P��)L����rH:��H�-pDJ�!ٷ���	����hV
Y�{L(����%��Ks�*
*���:JjETf�S&,J��(T�|�a4yԵ2���Z^��j�I)�2K+;��í���f�����A[k^�vgc�%J[=�"�xy��bK{}�2��g�>���j�����N.>,z�G?���|S�N`?���q�"����jr	��"?�?����^�a��vw.�<l�_>/{Q����0yc(��=�tE�h�q���:��}��@���)<���$^�m&�����R�m1�%L���p�� ���ɡ���k�nOP�0��Q�~Q�ǖ6M�e��+��jZ_B�Ry��4T�P�_�	"���T��h�e����<df��<�Kݪ�Q�5O��ӥlF���%�����?,{�h:��FC����7�yq��Q6�O�cѓ�"���f���`�Hޱn�ݏ���jXb Mߟ(�gx�V��eᮙ$�d�*-��?�e�IA�_N@\�@�5���to�|� ����1�=wDEDf}x0��c�%[ ����K9��jڵ�;㗗�6T=̓�O�B�W@o��ٌ}����A?�H�a�C4�y�Z���Ź4����]��+��DHɯ.��>���b��rA�
�Rc`���mrxlA�����B� �MK=�}҈�g`&>:{6��|�'�q#��~a�:��r��C�-&	�4R�J�5v!��1���FG-u�L��)�
����T�G����$}bt��kZjB�g���3�-�7k�]jiN��/JKap�tEI�M�T.)bi��g_:�׭�lY��9�1P�N�Q�)�^z���1�8�����D;�q��Ė���ܖ�z��~�o�'�qbC-y��:���uu��O��IMB�pP�(��u���=�}�ob���ݱAJ��b��� ���2B���u��,օ �'���Bc���k������ڦ���������1��H�
�'�d�[8��f��,��To\dH^�7����ef����z�b����T�ӣETFP�!�~���Q���{��-�9x�sڷ�2.hRA'����Y�8~����WBv@P	�Edj�X��������E�[��nE�R�Ӎ�k-gܷ:f&P ͚W׎^]���*<��@H�(B�@'qY��]i s�*�.�\x��L�H�wO�Q.�V�\�3,���/�rX�RW�ܒΫٱ���~�~����棨}1�b�ZJ��~_�ܡ�t :�#hHK��fH���1l\��0�-�����H�r^#��
�S'����x��1��t�e�Geh�o�[�.��U�A�B#)�����#Z��T�߿A����j�
=���x�h�ך���9p�+���x9��7i�<���jݿm���5����A�YVג�?C\ﷃ�tM��v�*�L��H
O35����.5J�*�-i,p�,��5����+�6�� �̣�w?es����G�09��3�7�ܖ�鸊��Â��p9�7؊E��ȩV-B�ˈo��Y�Q�Th�.�?�xCOyI}P��!��м�+J%�ת��!��H`J�6��hR��Of�Ο����7]����e�sIW�e�v2���pI2�M�Š��@:{�o�1�?��X�=[�v]������<�i��2��/o�Q*C���@���� o���pyM��x�+�uD^*�N�[��MF��Ů��yz|K-,�ݏtQ��^�H��;m�bUS��wce�:�����<WB�-1�D-<�%'�o�
���0����������d��Ar6Ou_��0y`}�&w�/�5�p���"������䧲����
�$��J���"wn�J��d��T�-ܞ�����ư̈́u)6Q���~X��y����2u��ؖź>���ڠ`ȗ������>c��+p��`��� sc���$�yE��Ϣ{�)����y������C�W�ϲ���H��>i��ȧ����da)�D׊�I\%7�F��K�@����|%,S!`5!ݠ�K~��f��\�֩���W�Zy7B-7l"���s,kŶ�ګ�5�_���^H��R��b8o����c#I�����I�ׇ��B�S� ��R����1���Z3��N7���.~���1i���,��q2O���a��̎BdHL�)kRl__�L���gg�����X�x�"��@U}����C������-fw+�r�e.�	UI+γ�S��I��E2at�G�Ġ��'��/_fF�h[�����p̋4,�0#�;�R�Đ��z[��N2��q �Y�lĦRYn��f�
��W7���/
��/14�.9dst�����k]��8�7�����+���������H��e���6��C�NU�BÏU�6��\A���)�m� �}�X�m��R����©��{̼�dt+����r����]�`a�F�W�����W,v��L���	����Z4�S=��9n�z�Iʔ��>���њ�}j���?���J�D��E$�Tn�zn@���X|EHM�ƒS)xTm�Z4�W���0��\$�8�#��Y����9�	;��Qx�B��W�����V@E��}!�9�z�΄��o�`׏�"b��N�ce�>b�gp��!����v�n��%��/�~�[���vx���+��M���K�M`8�3�a������kf���(!�e"��@�������H*�]-K��y����ЉCx�����c|��S+#z+#t��<<?�,�fl�dd��zP�ō���{�'���}O��q�~�Ԉ�B5"�®n�ʾ�'���D���B˓���㞈��V�A��<�]�
�)D�4�".Y�Ѧ- �(��̦7kFS��#L��[ �Ak��Sl����<'�a}x�I�R�+M.ᨘ:"�hO���1]�'��0Տ�Gٚ��J#�ë���~��N]�M��Kޑ�6����p�Z�o_K͈�� <U`��L� 9��$frB v���8��n�Kg��%ŪNL�Us5�x���-�l��<��!�	C4�-���
�'��M3p���T�ų=^�T�.r�X{�#�I�ĉŮS�ی�6�m�B)�[ݼܻHN�3�Dr��ID������?�zBP�]&�h���i��S!)p��)QQ��i���do����4��&Us*���a��{����OBIR�7;�&1��ї 0\�?��*[��X���5)6�A�����]��u�	?m����&�G�R8@Wd��Ͳ�g�T���+9'�b���ȇ;d>�����g�7��1�Z7{Ij�M�b�BSe�p9%����2B�7�{�+�4�m��r�Fj
�H��l6�@}g�e���?xґ|�&�o<�?��p��Ļ���@|��<8�'G�s! 	���8�U���ܸ؏�d�ub5���P���+��e�떸��p�fD#����R�}׎�R[��B��ƶK��hP�ƌ�\;��d��>q�k��S8$�Lz�+�k�8���6dȁ9)�-�#{[GRL8Uy
�q�oS^�JK�Ǫ�T��8)�hC��� J{�J��_=�R����^N�oד�2�U�3�qt��wE	F��]��$�D3Ǖ�OEF.�ҋ*T����A��)g���+�����|D�����j��tw�渆g��"`�Z�� �+���d˯�;aq{j�����h�����)��(�0ih�~�� ���M�vck�;��R��e�#�;�R"�G����_�3 ���I�fR��z�q���!�遦��tw�2����48�$�nE?�	���=�Q�7<1v�P�%�#�%�S{�y ~m_��~@}�������b�[h6�"����}H,B�o��'g�@���,�Td�L�S6+�j�����f��u$ܤ�w�0���@S}�6Wn;�b�	��d�Q:w\�,t�5o��.�p�9�I�O��5l*]Um����^��J�4xV�%iz8[�l��j�Q��{��O��Q�����n���c�ݎ\��옮9z�X�@0{����?JU~f�'�w�� �&	6�h�d���H�	�1m���QOD��dϊ,�:����9N[\�u_��@Ykz�]���L�,�`��Q��h�7)�����ߩ�@؉f�o�ޟt|��ǁ�Ts1.(�Ϗ�o����=�w��1 X��ݼ/��4p�\3��.��i�Ob)�:#3 �2z��[eo�aE���*���X��;��ß
�F�V/zw�;�.aq�_�`O]�|�1hq��<���*Y��o� ���� a�S�����g��Ƥ=%f����N����}9"�� G"E1��4���
a�\"��f��9��A�(\��� �P�<���R��U�k��B�p�|�z�(��-V����:��*_�����̤�����BB�ϻ��IC�мP�.�#K*���B��ŠOe=�+o��"��f�,c�)O[	e�R������������
�0/KK]��{,�E�<V�w�S��nj�П1
qpX�� ����a�!N��>��B��C
+D�Rb��{��p��'��ID?���ș�y~�C9�t���F ~^���FM��ꤟ��o�pb��&�
���G{�&؇���ρ��)�+�dPr!&��e酦�c�<��?Q��W�0�5�l^�Obs+�vʌ��e���k�s"X��
�$0�8��]2�wu�-Bd��	��e#�b	ze4��r�@�#/۝(�S����j�\���}���s��hd�G,���m��m��8�=m���B"nx����'��z�����M#_ DP�h7������S�����#\���٭W��nq�s�ъ]����2�+� <-M8e��o&B{� ƒ�6��g�ru��Eչ_z���r÷/�����������y�d�cc/<���џ1�t�h����a3.\at�WV�e�
6f)���}��J���.}���96��ڜdU�I��ڗ��!7` ���{~��no'~�	 ��kV1��4��~&Q�O��h��!�j��5����ER�
a>�P0:��X���o�3�����<nD��ȇ7ۂA��M�������M�*Z��r�6lS�W���ţ $��r8=);��2�VJ��L=��Z�:�Yy�R��
�����!�f;k�d���G�D^�6c,����\�f�MV�W�Q�7��M5��`��j>`��ZL웜�̝(�z�|��L�J�p �n~
�q��℆>����Q�j]�\����X!F�!���J=Z�dC���:���fv��Y����I}�K�sw%�������.L<�w.-!��<{������ �M�$�ۈ,��#^֙���Ol;
�c4��ņ�;;���:�"@ڴ=��z�N/HVI=Oی�Yyٽe����e��7��*Y����?�?"�Kp���OcNB���=���A��Q!f���\S�)R�$���Q�6��A�}��U��Yܻ�1` ��|��k�	{�-I�y�a��Trew� c�g���!R�AI��0���얩�����FvKV:���������K���	v	:=u�/�]�����β	Xo�Bg��Ʋ�%��6������M&q���<"��3��d��g1�Z����%Y�%z|�O1�֜��`����yF>7c���oa��e\���DY��u��#��4�-�����k_3}N�.eR*)�1�r�O ;�LB's#MT�塏<R����bL��Y�@����P�`8}v��}荇���^'y�Qa����9:\��4�v��m�4�]D���\-r�f�YOK���A�r }���Y��+)"������/���q��HP�?�H����f"J��2H���o����M�[�|����&!�Iޢ�i�z*�Q#q��9�|�*)������h��	}���.������L\)�j��S�`�I�+�?Y�%�Rn�:��/�]*`0��&�j�;�|ɱ��J�p�q�G�y�a�Ӧ� �\��U��5cM�S
�}uf���j�8�E/5����M1mI����w<zP֨`.�Fl����C�1��������s#K����3�5� �c�u�o�"&1���Rp�}$����Y��@�F�|7�/8�:f��%�b�M�G6��gP`��Y}��8P*lf��q�m�>�%� ��!�Q��%*��;�ag9�kL����Vq�'��r^���T���8�L`��^b��.�Y�]����ݱ��G��L����z�>[r!R }yq�7��4�_w���Y�;�>�1�	�OӇ0�iZ�r	����=p��@#}Q���u����,P ����RH;�G�I�F�(��#�L�u���I�v��w4r �;�8
�E��6�Z�R�3
�J���TO	L�?%/EX�D}�$\w������`FT�*X���O��"»�x׸�r��"�K=L����̦��m��v�Щ�^L����{$y�bϘf��Y@���N�x��г�>8�{q�I=s�Yˏ�@�á�O-�($>Il�7ӝ����,�����E�e��Z�dH�-qS;7��3H�X�?J卥�Io2� O:P��H$趮��1Uz�L#6gf���{�=R%_(�����c]�w�/�.��I�々�,��/R���h���Y%�o�S��4|A�T�����^�#t�㐧�^�>`r�J0��;J[�t�"HN8a_sI�ᕎÐ^6~�&��~�.����1i��R��i�8��2'�ͣ+�����ʙ��������An�[�։F�҇��6c���V�d�K��(oO5�ϧ�iL �=:{�u�tأD<���x�� oP;p�|>-Vv���:+"��{��%Y�J�:>J+��2��a�ӱ�\�m����}��:,�sv��{�m�h-�k��ᰉӢy�:��G��,r-�_Hw�?7����φ����A�ް}&�
�K��q{�^�*X���;��C��pT�sU�����U3^�����ϼ;c�?�U(N˙ױ.+c�W걫��ߥF�g_�{̛et�q���X�fT���f|( �|�7��d�?�&W}a���ë��ڝS�b8�+�l���C�/֚{��ss�U�Ò�A?��oޘ�B�����d?Y|�er80-�D4��H3����6�	;+8�nQ������d�YP��g�i�A�ο�~���7���g��6$�A*��!qe'��pA}�j&F�4�>�osq������m�	pQ����W��yqG�@wYqx��@��-�W	V��kǽ3�h�8��9.� b=��gꖓ��&��7�D$��1�`}{CN�P䮿d��nK hd�t�yx2�cT�#��V<��<��a�i���
UM̟�'F:«�ak�<�����07��YT$"��*hD�1`l�����0���I�"��,�1�m2Q4ek}��ݥ�8ϸl�Q�mҥmk�d	��}�[$�IG��3���`:��_y2Π���ysc��D�3��ʸM�d��1q>�˒�6!=q#�DĹ����I�
J��U� �L?�#I��8u	�XM���F��p(�u�`L7���h�ɥF.�&�$j��
�ƴȘ�mVH�R_���n%%������hK1$��Wm.^�~���A ni����	nAG>U������L����:�~M�>)��u�#4,&_�*�a2,ᘦk� ]����������~�擻M�
md��#���L�$lԄs�]�Q#jq䶦Sq+:s��C��	ߓ�(3��,��\"��U��;|ߍ.��um��,����z���~k�NM���B�P�R���k�u��P��ƷP2���5�ܺa_��xT.��Nds��?ன<ŧn���0�d�xQ���5_V�@ІȎ��a��>Nu���W�bP�CR���+àm4\�����Eu}����u8'&�w�?�vsQߕ���۝���� �ն a@J[-)�����K���o*������l�����ƶ�t�$�!�q�=�=*'�gT-�a
�0o�޳B�4�}~���7@�򰓊,p�1��GJװ'�RJ�S�r\����p�� {[�h���=���d�'�l��� �1J�h���0�}P�dGYr�R�`����7��)�5�z(�!�:&P0���C��O�������1Go�A�Ǖ���1���(a�R���#`4��7��7�q��wn�V3�%�>�r���}��W%"�(�C9qgqNn0�x����g(C[�87',~�P_S��)r�ŭ���P���=��u�{a��|Y�u=.K	5;�؛��חz5qs�aG�*��iy�f93��nW��H��DX��+TT�>�ϨX�d�����Y�O�Eo^nX��[�:���m�B�nK�o� _vk��jI�v@/I4X$C�{^�ѮS�<�����u˚xĝ'
cya�(Q�yp�9�C��J�uU��!�yad&�c�k�C���g�td��+�q��R���]��w%��]�P��!�����`�3.���.�H����7=j�A9@m�֐����8w��i�   �	�A>M�&��~c'��㯴��T�9�|w<��ь6M:�e��)��#�;2O�m�����N���fœ�r�����5��v�i�6���_�b�s�*r+x�?����I�򧨻$��M>�]̓�;�i���s�ҫ�g�wJ��lG�$m�ٓ,/��&4��8aâ`��(��F"_�F3�a�	���!xB�
�1硾`7u��'����8�/�<gc��C��6f��P,�k0��8]^2����G]�����#s���XD�G�wfٍ^!e�y�!"<�4r{;���Aݙ�C�^���Cq>=.�|����cu�K��<�@��1��ag7����f$�Uv��>��y�2,��E���V�?.�zO[�����v�y�s�4v�o+�ar���b����v��B�����X5h~�~���?���u՗:�-)�O,��Ꞹ��3��1�rc��H������ޮbg/l�8}�2��8S`���?#����#o���Ū$`���֦�y�A����Uq��F�l,[�D��4�1�$rl��pS���k���#^JpED\W�P@������E��CnrѤ�\��i�\- �H��V�^:$&7?ę�at �����Q��v�W�&�V�.���(^�S�Io���ܑW���'i���(+v���n���[>�tΐ�/�� }����V�mt2��t��?ߋ?�
H�cآ"����w�#d1PM�bz\J$Z�F���6(F����t�Tr�Sq�o,��hsST��66�`��@��N���HG�/���0d����t�_kn�B����D��I�8����4ԡr����ٓ�
=�!7��N�k`%9/�������7N	������#@��_EԤ�н����ρ㒅���q�RĻD��`s���!�/H��g�3���������YFܨ�T6�k�a�Ԓ�<�P��Н��,yC�$a�t�����-1e�dƺ#�"�@�)D+���5@�~���u��.>����)c��=��6���F��]/���~ Np;�8,��f!4QUз�*II�8�?�$��3!�F̠��dъ��+���B�c����y�|�Q��%�r����u?9��n��RE��7v�98D�}�1��N`�{G�S���`�R��1����4��0\�I�q���]<ۥ��=U��j$��D6���*��$�@����MW<^9�\�FT���7�<�)H���HP�V
�Za!��l.޾cm����4p��腇p�A��Y�lL���Pp�ǩ	1N�y�nu��M�,������	�$��	��i3 �5���ZE��?�*(d�)�MO�%_·]���+�j%���7��>���~ȾTo��M/jx������֣�C�1��W�YV�Bd|l�砏k�q��� ӓOC�8W���.��)���σ]��J����ڍ�@��~�v�>Ѓ-�����D�Vx���i�|	JO�\��C����w��� ��򛟱;��H߮�:Ǳ��~�H�=���֞}��0wBS�t�ͦ�2dm�*'�>Xc����q,��8�7��A�,����m=�����1I"�޸�H«4/�����*��qO�1�tWV���=��J:T6��	��E�J�[��R�D�����J(�*@4�Zu0ћţq�P\�QUC��@� ݟ���q�䫻����^]�8����.�ĩ�y��Y���8�R�t����N�1�ί~�G��b����0�͗�{\���_{���^���x��p-I�����d�Y������o2��U9rZ�R�ݺ�P�^��?gA�b��ր2mS��bkz5L�r��R�������vTxK �E�6�<����vU�`i���gL=�?|<�Y7�^d{l��|�\d�~/�:H�
�2���$�V�$�
Oh%O��	eQPo�GJ+q@��6��q4)�Ѱ�ʣ���,sr��)&S)㫐�ّ��E)�Y8�[�Տ���Ùe^�<��Ő��<���H[~d�~E�P/H����1%V�=u(Ҥ�,� >�Gv��Ѩ�re��3Q:#�)�nN����"���������`�?U�����w݇p�9XtV>��}<c�1 �&�	�N��2*�@�����P
�DWP�����5�ji<*9�ϡ���^��;�#{����i=C�V�z�5$�C����պ�
�/��-���@I�VA�a�m�I@���������u7�"�;��<���B�f!�>���A�+�0 �Hw�̆�l�wTi�gZC]�E]j���3��}#��ߤ8��[;���2'?�N�(�:�Fl�j�#o(�z�Q]l��r�)�����zf[�L�[a���\�	g�d� � ��]��_�h��z��/�^9�֭����aK�с٪mчp�$�?�>���G{�@�**�m�dl	Ӡ�ʢ�:�� ����cG��FIu��U[t�|v��.�T���N���)���n ��e�����"���f�1�6f�i�\nZ�`���*Kc;�H�ml�D��l9�����S�t�FTL�g|ڱ&a>��_V��|��X��_Y�Ç��ޘ��F��اr~R�a:6R��A����V�Cy��9��,Q�P��5uv����Hd�nU2/�B ��k!i�!��Э�vN���7����y���F�Q�P����%6ň��>�j��|U�?�tk��s��YLV�g]�s��R3z4���6��5|��P�Wk3��/�ޛ�3m���'gf�!ꁷ�<$��nY���C�12���p����Hy��?(J��p^姒g$����!�b<	�~��v���5�N����H.����GN�T 3I�ce��V����w���٬
�[�� !	�c��v�VK:�P��|V��`&������lE�;�1(�+��yCP�&��atD������-�9 �Y8�iೲ��C�'�g�e�/����=�&���oA���{��ӧ�@��+��ԗH�SOo��泘��m��Y��E��wM�un�u��Ұⓖ�B�;�S8rk�^��,tc��:�Y��Emj&b�ma)=�VT���b~t�"�t E�1� U򸤈X�n1� ���?��;���-_K*QM�a|����@�
��Nt���L�>��wk:ys��i�[Q�#�G�۔R��m��:��s.`��a
���������r�������j#(޶�-c�n���Ƞ�������nу��� ��i��rƞe�;9���#?l���"Vcߠ�#`���P%���}�\BJ���8f3	�'��σ������B�-��ļ���NXSշ���h���0MP���R;�ۖ��U������"z�}hΌ�T4���ڇ�^�������I�~������?l����f�͜�F	R�vb�~�Ev_/l�W��8<�.�K�ࢱUZ{�#!�Ǆū&�Xgէu)p��۫�
����Hh�7TxQP���=9����Y�T+��%�47&����Joɪ=2N�B�Rl�5�y:V#3>�N�qx��]��e9���d��$˾���Sز��8d�"���A�^M�v:D���j��n�`�Yt����Nc��2��(�zv)p1�t�������|ڱ5�\�q��� s.�_'͍������	[גs�tհ��X4��`\GӲ=�]�̠X� 0�#���qL�*��n��L?*������k��x�nph��~�)̟(��9t�d�G�v��hBaeS��]�~%�^	��x)o��r��K*=v����7Q
�~��{�NQ�$@@�y �ޙ��e;P1Pd�̄�
��51��i@�G�S}9*~���������5��k͆q�%�|GV�Ef�H�̢'+*���c����`��̴}u<%�|q\����:Ȁeti}�3;Ψ�o����"~0����`��hq{a��u3m� �T�C�U��O�\Х�	V={d�����{�u�: ���6�݊�9m<#�=<��i�����V�9��L��&jJ+�؋P�A�>���̗1�T�"��Dk��l��}�Y;��w�9놢9��?~ T�2��JY�zD�c�-��n���budO-����=�䶇��@{�U�F���Q�O4D�]�� �:)�����D �gS�?"#k~��$�S����&�����KՕs/�Fx�������!���S�o+���7�"��`�K���<�ȟ�:M@��M�9�j�����q�p�*��q{�\�(��j�P���_)���%\��@�� ��s��2��eQJa��7�XZ�R�R`i<�)����/-�½g�P׮PG~=���_�=�����B��\ݳ�*���k���4�qr�T�6<�:�|+Y
e��6��Rc�>@�@���vbk�s 6�6��3���%�ʎ���cN�qM5�-'�F����v��ܥ1�dQ��	�(�H�֍8�1�C;�ⳇ�h}�g-�W/x�>;�'�����hV�v(oZ��`��p|���ҍ\��s�2��#��gr��x�תl��z�qw�p�Є��p��;�9%ނ�,��!u����7�jEz�&�
�m�7��z���%���/�co)�4����y��uտ҉� ��|G�.֔6�Y��M�v�*�JW�\��9a�-���MQ4����>Q+�Ű��C�}<_ͳ��>��RɃ�[���6��`��G��`DQ���C�/#g�\P���KƵ���8ԝB`� �;	��n�E��S�/W�Y̵�����M����w�-�;�7�f�K�B�F'p�6��|����{�r���\��j�{󅤨�އ`3�oz�y�V�~������z�9ذ)E��}��rj�_�Lq�-�v��Evo	� �y��n�B�9,�̃Rz��ڏ�FG���OO:�=8>�Ҿ x���~��P���=��_+Q�;O6N�>���L2����:������J�=�l�I�$&��S������Ba�ᆀ��<��ZN��uC��pJUh;+�^{��qw�|�]�;P���z�I�� ��(�1�t�����y ��.��b������I���ي.�� ?���S3�Qi4V o�t���d&릉��?UQn���U+���K^v�����R���pt�LI���Xn�ʡg�� �f��Y��Np��^�\�<�K4� �{��������9rƓ!�~�i��[��I��}�l�� �0P���\��$�j���e�'�N^�"��+��U��C� e�@�A��>����Cly��>�E���F���x"�w�9��=�Du�0�p� h�f��W�бN֜�>&��Q�
)r���g m�1��-$}XRj]�>H'���t���4�hr�I7��±bsBz�S4*�twr!t�,�z?O��ۥ�Ok��<�5��lۄ�n�20�n�*$�[��齪X�#e�t7�Z�y�a��a�K�_��\�ۏekN��+�oǠ�����IL�����a�
�؊�[EF%J���ò�9
5�4+~7�[�0����a<0���[0�{p�lh�����مu��V�U"@�c��g$?g(i�Ġ��Ww�>����K>Z@&Y���Y�R����F��>Q�L�E�8_����`5�*F�~�vDU�,D!g�ì��*�
� ��"���D�Z&FV����F �>J��f�����A��1o���2Q�d[Bp�ADY�n�bS���q�Lܠ�������%/6�C�$�6��כ[^$�Kd.ah���Vt��������м�%�b�0�>IC�,5X	9{��ZB��s�L�R��B����}�G�l��&��Z�3��N�Cɷ!_�u�@�����&c����w���8���c��p���W�*Cc��B8F�u>"˘��h�+��f���~tI������`<��S	�4w"���t�~Y�ΰ�����nE'0B�|Ŏ���L�ć�m&�6�h�7�4�Ϫ��mBԉ^��4��JO�25Q�����(����}E�!-O7�]}h��b>���]�_֩�341�qײ \��EA�Y0-����HZ�����"l��\� _��n�P�,�;#��Y�bY��Խ�&��Uj����>���{Jt��^��SJfv���'M,Y�m�-��.�-�j+;)�2X�!��O�F���w+�E�VM�Y6
rd�G� c`��7��l[���|3�Գ	9��h�/2&>�x�����!wQqF�ʬ��ǜ?Ӧ��g�b�@�vH��g>��E��Ya`��RS��c�x7ُ��ymH˷�Ȼ��.�� x�b��0��	Z��L�����!�w#|������C?n�++)��0���e2�@�o%�މQ� r~��z�h�/{
����x�쭁U�b���w$��J>ˑf�zE�@����{-��1��@�ce��Z�s�d[to����3�&�ĝ7��#Pu��F�h)�BY޻6dO��:O�E��;�0n�9�94�L�=�p��onN����wM�1b�:c���!A�7�.�D@*)�j�؞�g�R�p)s�.��5��/��u�=.�Y:\�C�iv�90�����u�Y��'��4���Q�(�gėKC3[�����J����X���Bޯ��a�n>e�2:��sq��+L`?*��r���z��௑�?��1�n��2g㰛�q2:(2�\�� �K��C��D�.��]�M�� �8�B5]��DS�0.���Ά�|f|�3A׌�/��h������"*Dɯ��K���4���[�9�17��"��|�������]��
�'2�pU�p�"�S-���a�cnCeͨ�2X��n�n��u@�2s ��e���&� Y�g\�V���ɯ{4Zj��
h�u�+y��od]JD0�Ij�
)�Qn��<B�����c���*ts9q�+1���ٶ�_[>T|H��Ϫ��=���C8F��<�5���aj2Ā$[-�?��_6��~3�o�Ŝ!���#�F���l&��П��4��P�)V��/�	�'�����O�E>h���}a���"UGb$O!�+rJi'��~m��T�V�SJgR/��L����%��c�7��K�A�����$�M7�7*/�Żp�yՊcfF�T;�G�-<��	�H�>Pd�I�<K-'�(��'/cM��ݖ6���Z; ٹ�q�VW�>M�uU�cϮ%׌ɛ�_��3Ek��?�뼅r���+ˮcaЧ2Rȹ�z,�c*�$<��Qc9�o�O��rd@R_vi�͈U�~�u޺])�1ˆgÞ�2{t��0z���i�I�ݙ�:V]ҫX�N���(�M�|�0�xlcҜ47�+H8U��	)��p���-�~m�!���9C�^`Z�5+sg���r`t���6�Ü���������%�6��Nn��ma!����*Y\��l2&ف���h��-O���C~����eT2{��t�l)Y��~/��!��p�p8.\��|h|��U)k�->�E��xx�����YM�_���L�D�fVa沷��bR�-/����&G@Z"��F�hhQcu�`��6ЪY{�3*ul%�E}Slֵt�60Q��a�<�[
Ϧ�W&	!��s*�ojL�TzeS�f��@����Tw���Kcsҷ��p��B����}�ҝ��Z���Ϙ��g4�f�`�%:	��� ��Nc�'�?ɶ>,�Tj.�����[x/�@�\�j;|?����R'�A����2x"Z0�S�g���i�s��I����UQğ���!�tXwK�c:Jj(�8���sNU��@�v�'ضꍖ�����1�J�� D�a�7�R^^�^����i]�29�p�C��\Ci�Y��~��(3�Q�K���#���Ƚ%|��Bt����mgȋ���E��a'�w�!WY�i�������c�����̔Z��}j��� K����z�P�{�N��}=�SY�J�"7���U䳱�4�Ŏ���hM�O�Tw_����j1MZ�W|[��'x�^�{g���Y�5�[�b:�3qȬ#�d �/��}��r����R�%8U��~7B������UNX�;�|�w:�|�w�ە9�����<(֭}���c!���$2�^�ŷ��p�S�f�鎯SY��Ua��i���P�TI>��%LJȟ"���$Ҳ���A�[�u���z�U�p#��a=(��}*���z���]��S������|�R�=U���a�`����_g�?��Ҙ���[i�	�K�c��b� w�\p]���Ga��4y�SNp$�O���V��n� ��%�HlW<燰M���6�$P�����e��e~��IpEr�����ï_�ѹ�9����[�ƚp�ԍ��H/'M�nq�@0���1>�{$����
ypm_F�_&2�B���Im����0ci�֎x�FX�[Ջ��:R�j�^�	�^I,2
���F�۔���Fw� �ΐ�� �n��K�$)�[��Z�/̈́[Yn���ާ�����E�W �i�N pц{�;�T�n#�S]>��)�jpJfJ��J��	.��v[N��x.��ȯ�������HwS��1ۃ�G'�,)%z�ո��(��
��%`0&
zGL��f��يܰC���V}huY�c�3�FĠ�gb�"3E-#[�C��r)�%v�)Sڵ�[HA�a5�/�dC�\�V�'�\��+�܅�j�㵧̬�A�@��0O��}o����"��Ui4���c�C�B��Y��� �k��~o����SP�	|u+�<WzҾ��V�g���<��u�j�Y����Kȩ�ј#�T&�7�DA*�h�^��U��xWg1��["�bj��~]�A*�j��$37��Y�[��0|�Gvc�z��W&z�Vdu�ȼ��R
+���~��L}�A�6�i��~�o3Ի�*�]"O���� ��Zh9�6��;ߤ���_S�sV&H$���:�[��g͜����ds�R�$[¾�+�3|��3��~ l�I����C���Ժ����`�b��z(����^�VW,"�U	d��Ca@@� x�E�;M�={��.Y۫�O����݌O2g�l��ص�a^�O���	��ʒ�9��^��0���v�V�\���<���Ҡ���̩���e�t��;�-�)V����o%E[H:�#6;�|���&5G4~^��[L k��3�I�C6�B@�֦MS�i��� -|������#� �	�7�H��ڟ=`�!� -l�L]����� ����O�s?yw��1�&���d�;�3�f8��}�k0&����f�$l��-�&$uaEf�����@� zY�"T���1��d���S�M9va��K���I>��`8'#A��w=���	C���}�¾�q�kL�9X��bӹ���il�P8���_�W�<o&?#�{���l������^�!���P��e Z�����G�ga�v�:�N�tM|//��)�YN==��NF����t�<��Е ����d?�@�Z�oC�o������<��L�����Ro�~�4�A��*���܅*xMu#nM�|H�1�HN&��B\��s���OJ��&]�e�K�\S$N���������{�T��B)�q�F��1�u�k�MQ�0�\'Pz;�����
���"��{:Q4���2��"����_Ζ����4RW�o��#�.2jF�R3�.ˮ�Y�B�����
��_H�:o����ܱ�N`��&�Ԩ��v�R�Zw`����Ls״���I��D{���XB��Lă\�@�)Ç�C�`�@|�}��R��_>+�ǁ�쨻���NIWҽ�,�|l��L@�A����$o�!H�L��똭��t5^�M�sf2�Q9�H�	�˱���M�p��n���3*���%8�d�$�vģ�����J�F``�ʞ�GqUD��O��Gü�~�{�-i��y�4�uW��D6��7�W�鑘�h��&LL,�/�Ġ@�'�\�XZ���fw�AH�����ƛ����ۆƓ}3+���iҠ�s��� ��z!�O��j&f��g]�w:r_ghH˧̆���6i�4���͓��B��>�L�#��w�����t,�U�~b��@UF�S�O����&lK(<6l����ݐ°�����"��tآ�@e����3�qw��q�d;��ɢ!�j�6)`Qԡc�#��Ib�,H� c����#0b��2�#�l�U��݊�}���/��C��c,9>�;L4+:(=��5��񀐴��!�)�*�H9���=vc�4~s��e�V�[d�#�v��!_�ޱQHDP>�w�{��=�הkO�J�}����_I��#	����՝N�c�>m^�$ɕ!
�����I���̎Ƨ��<��`x��y5R=�FM��\O��
w=���%��Qf~�2�!fM�{ꨡ�n뾖'3R��m�JоO4�#ńhl�IC�m���������@'��K�� �ӯn�b�a��Y������&��>9�@N-5�GN<�A=>>�d�d�2(yL�}]o��j`q��td�z��?�@�'�x�[�]?7,@m�jYU?5�ԡ��u���6�~%KBX<�c!] �T!��/�$jQⲖZ@n�����}طI�vM�/4n����s^�D�B�(UC�?��]2�|�v��N�m�1��YR���[,���^E��xoOҶ�=�G�(��!O�l��`qX?/'�*�,誱���V�Jy�Cb�4tRb#��~úp��5�4�fA�1g��t��[��-]�����<�d�H�	-U�Y�7P�nf�#�u���T�����_���|6�p+�x5O]��o��>�J�6��/�Q���֤d��NY�����i�z��Xk�e6*�d��"��g{r�_)�*�W{�-��e[S��!:�lX�F[�5Sw��}��8<�"|�0�6��m�(��)e�6���aCO�s��f&m�/g�H�E����ݒ"_"+���)Y�Ҕ���L�@=��U��FJ�k�H�����`�y ���Ȑ0�Cw0�Lj�� ]R��Ї�똑���gz�$B２���{�6F*{x��0��WXe+�"�}�ҳb��[�ű߀7o�ֿ�}ɜX�۩p�#���di�c�_�O��|���u��;�ŧva�EEk���:�1���狟�7D����`<��'k���Q�RP�^�<�r��/�0X�"��HR���U� �RL�h��L�hO�#�wT틁�Ni��]���s���� 3O���]:EDN���ǁ�.9��v����]+�q���Խ�|:���������)�dbF���a��f����e�%�͚���8��P��uU�Abk�X�<�d��j�K���W�6�ٓk۪���p�t
�$�w q��+U�S�T���T�7a�-�RLnh �cyP�3��"0�2'�+&��)Y[:���}������<�ܕ��u���/'N������deͭ�',�JҸ�߆OY	2eϊ���[�G�@��X+r�)7�ec�&�J�=2CƓ=�h�~�Z����e'��!�xw�][�tZ���Pq)t��X�ru��r�ġ����A�yo���2U9ĺR=E��q�.��\�����18{�'�l�ۄ�Zl=���@�.?fZ�#E D:'d�P|ةQ�+S�AP0+�ݭ� i�'�n�]�h��{� ��T�8�{F��:�g��{`i]�N0S�(�j��S
�'��P��.�c��9i�QJ"�A{�xo4������s�`$����l-�'�}���c��5"�ڸ��z���R{~����vH[�I�T�3D؎Ȕ��!��	�?�����&���o��p�&M筪��;�U���4�h��c���夣�A�`
#%���[Bȸ�_��?6R\���6D���xL�vGM�&�j��޽��ҟ�Y��!�7�1.��f�nt�t-D|ɩ�v�
z��!�K�>�m�h^Ǡ�iEOc�0ޓ�F�T�.���`���#���`�d�|I6`s��)Z��N�ɻ[�<�Q)�����K7�Ǭ7��ֱ�m.X�<�٣%2Ó
����8� �0H����j=��Dt� �Λ���/rG���&_�GHd<-���H�8��<{�֚�.)v�r�f?��[�%��Τ�3������{�.�=4	j}��TDL�d�}t"k�c*�@��F;�W��#eǬrT�����s��Rh�L<)�W4���>3~�S��4����L{��� .ЩO���4��-ȣ,L|�c��e�}�Lm���Rt�. ��.5���bIf����:�G3�$�<�ڎ}�4[�H�럐鍶Kc�^��^�l������̛��9�d������A"0��;��A��gGst�ߨQx�^���YO�#b���ի�<���v�'Vdˁ(��s������c>lzM2�%;�*,�	���c�'�t��g)��@��(ѽ��E��S6����)�x%B.A^�Nk�6?��sԀ�����X����/^�<9"�a��`k=��d}'3$G�^'��ۆϹ���������l�_,�'ř>�~�_��7�'�>�E�����lbęV�U�FX-d�P~`�(��L!VDɑ)�[��#G�<�fOb!ߦ[����KI�z�=�z�D�Z$�3x�R���L�,:��F�k��k7y@F����Jͯ�G*aS�&&��(���HG�C�:�"�GƵ2]yZ�-wp ٟ�xu�	;�u����``0�EW.��6�j��#ҋ����%�dC�P�>��PM��ggb0n�d���vW87ڀ���/.�w~�S6�6.���K-N�A�\�O�v�(�*s��xQ��ez��⊰R`>��N\}k]���K�!�{N�%�R2^���B^�����_�QS����$�pzg3��Ϻm�6�o���Z�ú| 7�c��g���%|4=�W��E%rw׷�|��{�M��N���!�gg)�q`�b��	�S��ŉl'��1�!7{F�\6m3uZ�pA�pV�b61�f�(��t����XwuTRC���F�[|�'�����0σ�E%n��ރT�I�Q��O�NP��5��)����u	�j��Z^C���"+�˂�l��Y%�w��Q0� H���0�$��S�o!>�����R]w|�|�'-�z\⵭����&!��`�'N�!o�dKz����K���Wbwa}Y�Û
���%vf0k���o�Nk1uJ�¤�ܓ�� �G�
(��d�"�PG9���^�H��\Q=�`��X���y�#'sK5����^�����a�{_G@�gv�|.O#�	�CdVR(�Ϫ�iM#R"9�y:$oE�h�g���;���N�T<�U���~ܘ ���7��i�~�{S~)2�*A��(R$yb���{P�BB��Eu������g.�@8q�{�����k�K�bl��v�����A><hc@��w�b��b k@��"0nF����^�$�ت��VGܫ[A�d�`�Ww�8xx���**vS��tn�c�2+��fq �z�Mł^n3��2�Wp<4��qӆz��L
}����؉j奼vաa����s]:]�殊��OmC02�Q����.�_�!w�:������R���Z��O������9��,C�y�s�?U��QW��.���W�_,?ުI�M���]�.����`]S0x<4_ϸ�΄�Pn��r��s��w瑊��-Hғ�{9��,"��s�3݁�CT� Ygnu�ԡRr�6զF�N!(�����z,���4�wb	�b^z�n�\�7��\���381�o��5:n��\��53�7}X�%��h1,V��j��B�4��4��}{��G�%Sd�R� �`���ħ}��D��QB��e 0�BSHK�����;2�����k�_�>�`��d�O\�ƥo{��y@��p�=MP���WV�ß��W�>�u_;΀�k-��}�W�d����Y|���M�}*�8�i�}��h��U{���q,�J)��d�A"n��N]�>�[�
58��Bv�u\�h ���[��_��-ǆOfCb'��3&�(�����O���ѝ!Ϛq�/ő=�#��u%�s<o֮� �@�q)tH ���f��~F��[7#��f�_�
��z�J䰢�����4I
�9q,�J�i��`t���\�O��Ƭ\a ${�B�,�1�f[WŸ��)�:��E:sX�`�m�V�2?�C��C��I/�۪I��H���@��R���=L{LZk	�Jl�K��g%@��d��M�$���6ћ<W@�y�{����}Qv�jyɌ�Z<6�7N)���Ys0��dH=�N�E�
C_
2�$�w�_�ޭ��D7}Ģ�%�T�G��ثH��4ʵTk�Gr��ĝ�HC��A�_s�>([zy�>k�ŝ^�ն��w)K� �u�Bظ=�#ȏf@�)D�	�dx�n��?C�k�ܸ[$v��v��⒊5�н7o�8�#5�L�R�m9���9�j�P��S$���VM��=8	7T�,/ZX����ɓ�c�#�[�ƞ���e�MZoMi�?�|�3D�P�mQ���7�8�~���}�p��%+��#�m�  ��D�f�aɥ�Q�|�=����	1���M}�T%�)ۧv	�_^���<�1�l�0W���";����P�S��',1#��f����|���y�V�*�?�HFuJmI�i'皭��m��3�l��-+�0�"h�F/o��[X���b|�t\�&�>o$�V�tG�r�ug���Z����F��8%�A�Q��N�8Y��]n'���ǚ�����Y�1�$�5�"��-��n�%}����Г�*� +BP^4Oe�U�j�iH&����V0�zy��Ē#%3�,�5V�h����7��o�<8˲ç`,�ţI������¦�5�~�P
���=�m�=�p� ��'>�;��N��)�jY���i9�������Ȇ�����B�	���0�[�{�#\��Z�񣆴�A$Q�4֋���D��N%��:O�L�Th��μ:PP� "A[��?����G`:�N^��>-�sE�����pB0T����+�ݹ�癥J�ܩ����6^�(� ��0�ꚼ�#�����=�YDG90�K��D��]77�kظr�~5 ~�;�KJ�t�N�"E����@�#u��Y�{�E��0%��48�_��q�T��!�����m_���|k�X�j
o��>����ٵp�0��:-$��(׬�=G#��)����HM/O�8:���af� ��uy� ����؟=J� 3���m�Tw���M{I݆-�1< �;��=-�����=��I��s<]�k��(�B������.k(�z޻���= 7y�M����C���:�-�"�A6���Ϋ����Z�H�%4�!�R�ʜ�x_I|z�@H>����w�`��ޱALy�{G�M�eŲWofr7�q�>�ˉJӇ0�b��=+���mͻ��r:�ݬ��R�C���m��{�A�B�?������}�s<���Ε��b����1ܼ�bt�}���MF�vGnN�<J�������ל*�-z������1{��k�/G,��b���|+��J���F՝�|J��\�&�m[�AW�����l�?��DJ�铻��@�Dy) ����P�������[;���S��.j��]��l��q{���W�������۟�t��R�'��("����@'AD��* 7�G��\u��~���
ՙ͵�&ٛ!�	�n;��Ѐwo�ɤa0��b:P�!�;@������O�>*���,��[-�dۚ>��h�{vz�f7$��6k��tB����W�?��:�b���@��Rq�`��W��==��"�`��!b�U�ҥ�KBnힷm����o�Y��Y� a��Pȼ�
��-"n��8�`^p�<���x$�ZT�R�dd��
�$������-��ŃD�kiv�.-�z���g�&O�X��W��Y�ӧtD��^4i�Eq��������*M`����u5�	�3l��1��4�������p}���Ѱ�ݐ�n�E5W �ݧ��`�DY�H�DMsK�m9	ӂد��(���D1�Y%�Na��b�fZ}?���`GӺޥs`yj��$��_9P�\y��G�������}�"P~���b�|g*�-3E�(K9���25. f���&�`�M���&�~ЏI䜈��撃#,���[��=[��ঢ�����ΖH����}�Z��!39H{sa�jEfsp��K�V�NH��cU��W��l��6�B���1�;"��V�8&��z�XZ� ��o��RPtWÒ����,�|�����<Ȱ��)+��礿I� Q���c���p��&l�-ԦV� dj)I�
�����[үC7��oQMu��FD��g�JP"���^I*��q�ϣ��UE�x�pph��/�J�������Z&n�jm-2B�%b�?�I�z���b��K��i�Gx����-��{���ޡ�@�T�y�� W�%��"�Zg��zN:�]�e�ҡ�	��Fp
��s^ߚ��ƒ��)�>�=��cMmv`N�?	�޲�2k�=�v��?O�V4��\)�֞Y��k��3�\�`�F�3G�	��E��)l�Zԛ�6�\���qٖn�P)�1�+��uqd����0���J�H�A����BOģ�?��R�Z�k���תrNY�+ �OʛI����Ԛ�OA��񕗸�����Nwjp���ZD*�$G9*/����yhSޫ{V���u��Q�o{M�ܡ:���=�aM��GXٸ�m�D� �Y-E�e��q,<B��A�����+��%��Xz��L(ĥ��&�,�!
�\��"���Lǳ���3�՟|�]+���B�*���{y�l΋�ǕW��C���=c��n{�G������,��OK{]]�\�G�!�T}^���n��f�Aq�2#☓]�BMD��{��sk4��F����(�L��xB�<���u"�H�k^�AbO��C�x��"���)7>��4q���E��/�c����X�/��c3��T+�:��w��cÖ�1�;M8<���3s13�C�*�yn!���,]�&K�����z�����Y��(M' f��Ĕ!^���qJ�-��Ѻ K�kw_=�7[z(�}e��Q�q+�v�j\��W��w��
�6�AB�[��4W����ǐ�2��e)˓4���߅�5?&Z|ŷ�=�\M�`��.}q]�����ٚ�J+�ډǤ���3��^�0`�<��\-�#�*u���4>;�i�4 �����£��]/O%O�}�{�6=a�-J���-{^h1�z�-�����BG�gV�[�ό�n�w�X����f!0�Քώ])B�?SGߧ%|@$�ކ~K�ڻSP�xl�=��{��V)���U��N�3_V��[��"��p��@�����X�:gl(F�=�ˋ��M�?
��H�wd���a�(�J�۞ܽJ���Ӂ�#����JA ����|���O�
�_د�xُ��"d���� �h�V����be�lT�h�ler`,�z����Rnn��q#,�|�Ȋ�� `��v_�|��(l��Z����������y)G+��Z�Ѫ���R]���5�O�T�#�~@t�a����;?-��W�{c}��7���B�GuM8	J\�3q体���D�r���D�T�,����,o]=&Hй���ꊶBT`vK�:?�(`
����qN}�N��'�>>t!>f>����n�F�/�+qeK`�C��? $�=��d��$+��69yL�SB�.XwA>!�裮��ɷ�/���<�H�s��ԭ�� y�|<c�s��T�p��%�a�p0{�u�nuV��N0e����풨)X�q�I����o��t��[i��6'��f��'���f)�<wLr����~��fUN�o�d��ńG��yF(i�BUS5l= �L±=|;_lm�	�Z��/����{���E�hb�`����2[�:��U�[��(�Q�ZY���J�J�)���#ZM	FĲ�]@C��WJ��#�@������Dͭ�:���U��'��9��Љ��}"w:���V��~��3&���.�����vr&#���T�!;W��#)~G�Q.�U�m@=5��ͣ�o-5#��B��_�J��s�/R�Q9��Y����f>3}�z�?�Y<��*����&$M, �-zgo�`Q�bL\Z��i�������O)�� �$��ݕ��BJ��@	% �fH�Եh+�T�۴������*eT>���[*��z���qu�w���Il��ёFVw2�i����d���C)����X>��J��9�eq��Gֺ��g=w��"��JN����èv�B7�Y�sQ(�#�����^�@"^S+��2&�����]���V_R��(��
�{�1�?�$��|9���p����3/"��Z؆�ʩ0]j�����zc�4�'~����<��e�xK�G�i��u!�~y�抉�t� $'��t����Q'&c~�=��C� X���
U!�Yws��,g�5��+�2a5/�e���KCp�0�(�V��?�Mh~3�y#Q6�Pa&o�V� �
)���и�	+�o<�8�4����Y�1Y�_r��rK�FVH�{�UV+A@��Rw-i�gJ�G�q5�p
�{bs(�j��E�(F�ף��ީ�_"	��'�t@Y�ى��t�x��m�e��f��Muq�B�wv[J����SV��P(�i��sѢ�E:���?Cv�������0�<�@t�
�߬�0�<R���6D\* �Ĥ��NP��g^��G�K��yөI�(�X�
o�$k�8{��CT�V;ˈS���;�a��V��&x�)Bn�k�̑���	���Z�ű�λ�lK���>.p�6���In�)��j�kǅq�_SJ+ݤ�����?�/([	cI;��i��]Cn�i�&_��!/�k#�Ez��Ӗ�	�P�cj�u�bT�vD;�˓ܠ��#�l�H��S�����y���iZV�T�ƕV�	n1˔�DDMe��Rŷ���P��r�B��әv�C���bw��׾sSuw��&�@��`�*��n��WI4�쵄;k��Χ۵�k��˃ �1��`���4F����u��~,X9�D2N;������#�
E'�������P��Uʆ:Sc�
سj��z�\�׳�;���t�c[`:���@�&�9�&�q�bA��?0{���w�cM1����YW'�g��~q�_ý��F6~A@���'6w�۶�Y����t����2�ho�������
\�0c�@�A�3��Os��5WLژ�Lk��Ǫ����)]�BXZn��? ����R�$�мk����q"�����1h5���Q�3��S���a�e5�O�іS01uY�\����9�R�zi��|@ʹ�nR2�e)�`�2��S�~h�9��Ȃ��ð�����|��1�*��C�Ӫ~�]���&�����\�Σ����+�%L�Ch��^`ceM�`�G�9W�����6\��Q�3����(K����V27�O����]��򹈺?8A����pf��#�L1e=5"d8|B����W��%[�V����e�����[�Q<�le��)CKf���
5�k��3�����\a���;��2.t�}j�̕ȔCl��
s�TC��U޺!1��p�h���:��|;JJX���q��/�\��U\���(+�׆=� M�Tj��Fb��4����u��Ubg�' h�Cp85��d&U�/�?f<ZkJ���VjP�S�r��_�B�����b죞���V��b&�~���K��y��L��]ऑ��e�[h;��j�tqྈBcPz��$L��ފA�L��Ⱥ3�[��Vi>�D�uDd�<�&J�����@~���3��
`� ��p^8MJ٠R��Eb�G؞�5�T�g{��)aB�K&�}X�8�����/4�K?sK ��)#)*��۵���3@�x���C��~q�O8I������#�g���޿����پ/���x�]H�v�jA��C�m�����~��&��� Ȟy�"*u
�?E�~��HC
�x?l�M}+���`c���yl����,�8�|+TN�	��*����>�n_$�:��6��}�F�R�a�-�����Ȁ-P�,Q&>0�ٲ&��R/��Գ�o�d�
]Y����Idn��؉~w6̰�|�]�h������?E���La���o��!Ǳ���\��jQzxِ�a�k����m+�h3'��J7/��H%���+����F� �Q�Yb�����Z�*���~���v.��&�8�٬�׬�[�9��M)Mٶ���t�sm��/����{H��''#Y���%��ٝ�b��P��Wd9�JȎ�>�mg���e�f;X���0�˃�%��G�N։�l0$-� ��_�c ��0�2QG�u�a��Y$�zJq��|ad ����"Z�����āoI����`�Dg0Ǘ��JDNR�����ڨ��$��t���Gi�\�-��H5@2\W�0�� �ʈI�P��ۖ]n��i���1������~�$�a^��~�����㏶���$s�)y7𪴛��#��8v�:I@!H	�|�����.���~%xd*��3�j�cO�ZU&�׼���-Q�z�5����ͪKa+�2��S��:Y|�~�?T-�b�Q�+�R����k ,Z>�+���N/���u�{�lF/�ju����B���j-�2yN�T����G�X�{�-N/��Tb����߽��Q|`�p�.8=
`@�/�f {]��"�8�����d���}<>�ďH�I�\'HF�t��D�Χ�.8�׋-�_>Zp��q�:�7<��{!n� �8(IN���@�����,̳Aץ`�>��s@�1Vv�δ�ɓP�(�	��̷��^�27�㒑�Mȟ�Q�wzc��4��=����O���F�ћ���*�l���9(�� �#�����~��I��*b8;�_���ĥ,Ϙ��|kA��t��� >������bw/�?����8֎m�>2Jц�b��T["GK�
TjP��9��] ˞"~*���+d�KUݭRs�!\�mAؖ�	�����?2�7
[Ӂv�-��ha8��E9y�1)ӷ8��ehU=-;q�S��|#����;��`NiS�8E/uR�x�*�5 �e���\�h^����5�z2�1]���p�A"�)�y�n�|�Y��?Z�4�%�J�`�B�h��- �"XL�D۸�C*1o���:5��2]؍��4�m���{^�[��T�4J�SX*`z0N�ɡ��XӴ��r�h�;P�8�E�˖D/Gr_�_bZ����Ͼ��e���ůN��}��Z�^�4
��R�_���i����R���c�i����f�F�5X[{�)#z�f�LS�(�מ(�
&9x���#A���sdJ��%�Î0�KΎ�#��lU+xә�[1������J�W���7��D7X: 
��N���)[�@ � ��ѡ|Pt��<e�	�eX���	"�	�ܢ��E3����x�^ �&P��3?�83JEͦ>��5䯹,�E^��#yf������}]��.G4�|�����g�׵����7��q���o�?�������<�M�'�|	�!�M"<CR"]�+n��)���\ශW�K�,2�X0�i���H�D�l
E$Ƹ�2���$�1�à�k��S6�G!.A�5�D��4��V�/����ɳ�a�~?�|;g���Sa���0��$4+"K�u5��p��%?���%�挭C��1�܏X�dx��$'��0����������h���A�z����Ma|g����u�^�5?�����)���h1�C��xFҮ��.�$�5���~��"b���՘�3+y[izSm^R��)#�Q�>�.�&h���D��Pt����o�S�P%Xٍ,��'A�b|�y��t�{~�;��%+\o1d���p(k�ƥ��V�?\��Z����=��x[��&�)�bא�����7�����c�J&?YZ�iKt�vR��]���Q��ri����+����"�Юa(��2�X��9��XOB@1]��l��#����Ѓ߻_?�4s�Vˀ��M�A��_�\@�@S���V	y����۞,i���<2c`W�6��ԁ�S$>WHT����9,#�5ν�s"Q%�L�^�'4q�@P@Qe�T�Ry�U@60�(rg�E�,��������Q
��X5	@����Q�����漊V8��`k��&1%)�cI��й
�E� (ot�+eKg�̼�x��͇Zeb�E���d�6�)]a�-A�N=��1b�n���ɭ���ǰ̧!�W���ܑ=�:Q���c�]e	��v}*�n�bw�����b�gZ\D�
4T�׿$s������R�E@^����1�>y�����Զ��x�̉��pZ?��q��4�	(�B�4X�������}0t&����To��|U�:��}���6�l���&w�5��̠���'�ڥ����[�D�a9�M1R�&��	�&�)�<���eV�~6�N*.2�#3!{���yp�w^���2NT)喠k�U1_��K�@W�x|ı��-�aO��`������������'e��Uq����}b@-R��-K���/���'��0�����O�3�Z�(պ5�ڽ�i���V&� I�XÊ3�Wښ�.d��|n8��1�uƓ~|W�|e>�3�V�T�����V�'5��m�1�t���Z���w����+��g����Z�7��ʨd�����8�3bL�mo<4���!*%�����䫳fb�f��|��+ wbw�O
�����9(QfJ9X+� Ƒb�q|-��Ic	���Tw����υ�{m]WMR(��J�AݿQ	���
N���ڈ�������z�>���0�3���g	B]!�͆��=*�\��D	mpq���P,<�Վz�o{�\9���#�*��w�?ӯdh�^/�ճ_����X��Ḁ!J���*��uzNQD��l���t����'v{>���N�������w5��L�ʪܓ�j)|�����)�� ȼ[��)�XC��{A���E���݆�≰����b�$Vw Ӣ���0�-dnf_����I���s�z?��;�5�pk�9��[_2I�|对�,�����4��S~�;��<�Q�J�"��u��?���������u�X�+�"��!y�Hq`��0v@%�Z;o���{��v %D��ʃEk�[!��Y�@�
����u;5W t\Q�X\�F"�Eࡪ9���:E�ps���g��(�{��b�r�������\Duy������[w�F��A�|���:���޿��IAd��t�8C` ��U
Ȃ6N)�N1W>�~�V����"����6`E�<���決�N{
"x����T�hm`ˉY0�y����[����������t7��LT)ao;.5�~dq*u�k!��J5E	�(��p�.U�"�d�f���D��֤_U�,N����O�_So_��&�vR �g�]<�	S��$a�<\�y����/�G��[k���(�vw���v�.-�G�e�.�BUʤ���/�G}g��5��a��H$������B��Б������ffӷ�z�q�b��>�(d�.��ْ�8�d��fz�'B��_|'�z˝r����o+���R��wU�J�W( 
��U�˔*y��hLmO������U��~e}c���U�o�z_��3��]�Pjt�ɵ��/ʶ�����9�8�yi�i�uǩ��R��4�M��q����?k_sr	{ ��/�v��j���0���yBU�4P����.<��ε�ݥ/J+f̥���qd[؜�2���fi�]��vx�"%� ��!(�sg���J�ƀv�,��20}‗��r�rASR>�74h�F���U'h�A�d� ^��L�HSȏۆ�i^��K��|�Вϻ���f��vx	�v�+T��͔�e�+լ��5�Co�Q>��2�k��u�]�T�.��(`�'Li�򡭉�e���괃��a�Cf.�&8iΐ~8�/���T5�'hZ�Cc�^��֞� c�}X���MŰ�����AK��]����;v�f����P��5���������/�qr���|j� �/�����m��)���4��%	Dt���M�kVc1���*�W�{!/�]��)i�\c�Z�܂�Xp~�e����˂ �P��2��GB��Bؙс{.��[L�Y�eMlBz��R�/,^�S�e���{Nv��+zE?��}"�ű�L8�о�w$
�!]�h�c�GB�Y��J��D`s:�/���S����N�,J]=C�8�]o�0���O����� �C�#�k��R�q^3mdO8Y2�=�ɧ��5�B�\J/y�^�/�u���)�5�'���_��o#�i��p�N�1w�J�B������d�e���)��L��.XP�V~���,$m�EbB�J^�J)z�]ΑX{�����h\.���2
�����e��N�O���04P6�������g�=>�fC�Ux�l_�j�vx��O/���f��h�$�I1F\��a��|JR˰�!zɀƤ��sW&hǅQ��E2����yL����r�e)[|��Ϸ9E�'��Lz�5�F\ˋ�.J�м����Y��M`R�b��(E�~<U'L,��ڕ+ޫ<����}M�YH�/�S���F4MM9w�����,s86��w���7ɤ��d;�y?i��ڭk~z�?��P5)'_���6v������� V̀�e�����>����bg�h>�-�E��@;�{�ؐ! 5Th�g���%q�B�9+G����N���7
�т�1���n�t�#����dO�5�R�^�7W��cå���KИ����k�^|[�g��U�Byƻg13Á{�2�5׏K�5o,�/)Y�#W'��SG`���.�&�SXa��o�s[w�k�fw�k*�6{���(J�4(�oH� ��(���`��bk��x�J�Z���2���'����D�<ԫZ���ե(kt��"�ƴZ �E� ת�ǥg��X"�>�ƽ�ǅrO����$o�mE���8J�,,a���Y,�l^�4$��%^��c��#[�$�Z<	�d����Jw�8�q�S�~����o��Ǟ1�B7_��b��i������9/.��a������i��:^ �#���/�DN#�{G2�jE��Ŗ ���f��Rc8�5T?��ĳ��M�O�xf98�	���3�?U'Y7rҿg�z�Ypo�?�������jL��6--�	�n�R ��T<�b���H�`Y[]���z��7r@T����\t�����[�%$0)�����c��iW�:&�E��ӧ$X(��g�9����o�/Zk$$K��6_��}@u9(S#%�R�hr���<�����F�6��0���$e*I�@H�*�eѸ�Y��ۭ2�����`F̞����x�x=hlK����U���ki��z��-yje�;~0��bja�J7�ơ�ᶽ���ѫ��[}�APQ:���|�Z����`ϝ>DV4��#!����X�~v��EʴG�(��}Q�Xvn��8mU�p�y��~�7`	y�9�H�L�e����Sy*�e3����.�@�ȐW4K�$TОI"��$!�(�c��M�����d�d�M����aK\ں�:�!���"��J@3�W+�4˓�' ��G���pW�,��؆%|���>��3�me�Q��߃GV��e5
JG�e�>_v��\����C���e*|�v�<'�ؤ���x��WY��Xٰ�~�ǧ��� ����c\�S�߇7���Ҏ`J�3�s��D������ՆT�s��tж�O'���N�${>�����e�@�������u�ܧuO<�Ꮍ�@˞A����w���l�����E�?�S��:�<"n��ˬ�&!)!����?�H�%ڬ��%���6�Fk�,JIv���3bL�ET��%��D?Y/���܈4���Nf7>-������&��Tcy7u��)ý��$�+Q|ҩV��S�v�;�%�1F����*��Jl���Ti���ۨ�o�ynHv]+�|�1i+�CD�R��>H"�u6�>�T7j�'��o���5%���2�JHl���zd7���6�ˑ��N]�D/�k1�E'AK���+ߣ.�V�w)���)U�@l�m���Q��@u@WW���UI�}�̬q�>��d��nj)�)�����_�5cWUr� ���.��9xmđ�g�@�C# ����s���C�`�|�/#g��ܑT2�y?W�����l�%M�O���+Z�̚�n�����@V�xW��'٢���}7.Q�}�'��NG�u^����,�pLڑ��ev���d|
�y 0��%3ɯ��-�p�<�A�aT�	E�a�,$���裂B��d���Y�\�}Y{�w�kLL�0�3�GӶ�?+>m��S׃Hj1C,�A0yB�`܌ސ 8{$�]zrUQ����n�3����>W[�a��
bǷ��=�n	����L��x~-1�v���]_2q�O{�=��7H����qa�ՙ����樾Hh�n9"����3x�.���cP��c���W����j�;���6	�c>$�tk���˞]�#��
��T��R>�8;10�W���RaR$�l��ײ��Խ���lOi��F6X��X
���������F����Ȇ��W�l';�*�S�zg��@N�����B�2\��ʳ�$�$F�\�	fuك��U�^�dv�}BrU@s�������p�F��&P��p�#.ɾX�.�v<ο��>��s�R�KU$�Y�5,L	������U$�{��^��S��1I����vݥ��D�:�G� �%/�2F����
�����9'��y~��'�
�+8}P�C3�r|�=���_���z����$�����s���� �8ata�rqD�I���0��M"�!M���ʌ�D|����p%_�hV�ۖ����#<tz6��}�L��|�*�mO�7������e=,�۞B��5�AQ�Ri/���s�!�`�sx�?y4cĖ͋�mزz�X��扥����?�7���h@X�S;E��`��s��in=���.e�\g7���W���~o9�UYP9�`�o����5+�,�����®F,����]�s�n[_�3�ٺ,�q]o O�)_�`��yn�C�qʖ�B U��&a���MN��Er��;����{�\(�'���q�f�<:/+jb�.��AΝ������y�sǀw�`���.p���H �%����@em��P�>���d`s�1 ��U�7�^�F�f�
�3�j�(a�Υ����dø��U�̱J�I�w�����f>J���t�g�L@��ω6'n�06i3��#�nP��3?��V�#xa�S',n�e��EM��ũJ2N�x���?����&�G��0��LH��ԗzw~��I�;'-+��]nc�8�Я]O7���u	��!l�^mLও�=���br�Р~��:�����z��,��p��t�p�Fx���dÌ`X+�����&F�v��D�`~j�V��?���ˤ|�r����]m5�O����r@��i6����١2��w]2���1����#�ʐ�D��иD�B�d�P=���<2=���a��ٻA�XP�h�"I�u ���bv�0H��懵:/tR��^�zN^r��y ���&xyΝ�S(8��x9O˾��V|P�q��O~m���M�-Ko�\�ꉼ�DtU�X��X��p#����I2
�SL�ϵjU�O��PV�/sHi�=)6?4�V ��	�@BG�);���X��p:g�{�� [�R���ː�a>�&�=�xX�����d�B� �F���{Xt��I�h�anL Q�V�*4��ػY\�.�����!�۽0��r;���~L��vj�2UQ��莅��$���F<T�? *���7r�'�6�T��M}'9+v��b^�ˈQ$�Ce�\fb���������J�1��ȎⰙg�Nr�I�T��
��O��b�nJ��TF24˩�?��@?-� @��H�@9O6���G0��r�V�sU�]���\1
(>=�R]��u�����ZN���'w�#�ba?V"�ې���^��Uq���T�A�5`j\�(Qe�^'K�o�Eo횝Y���}kZvzˆ��=�Wm��(n��aP��S�p�P��T��YP"Y��ۤ����� 5�2�	N�YQy���` �>��!?��7W7��Đ=6��E�o�a �EG�{X�����PTҼ��Ss�V)�B�ⵯ�"8wv�5�j)��L}�4	����p�<���j�i�YC�#�d��LA�WT��� m4؜�#�b��,��� �P:W���=M���ڸ���0=�>�m*�p��]׾�߰�0�@Fmǥ�&n�|�û�r���t��?��6Bn�����&�'�R[�B/�v��;[��/BW ���$�D�~���Cx����9�����5h2�cq��kl�@�+$iY���x�h��Ix2?b�`)�B�"��-P��/t�m�N���&|]c�1��<6�	Y<Ш|)
��	�GJy|����ԛ�qL�a{Ay�GF����g|:-s0��P��g�;��l��QV�q�$_�r4.�q^8��?F�V��x�%�Uz{��8_J�w�o\����9*~Ɍ7�u��Ϣ+/Zlw��G7�[�EQ-�um�Wb�d(@���2&��．Emq��p���~��3�{�4�=��9Zs%.������M� \��_$�����0�w���Z]�*��s �-õV����t���ooyL2t5� gr��Y�$������x��eJ7��ݢl���ls�^JQ��z�>bñ��8�y�؛��j�&�-h��C��#:����/	OY�G�8TD��'�-��NiW(ݾ׀���"��Q}0�4�*w�_h��e��nW��Q�#Z���Pq3���_�g�V��V�0�k"�Ifp�jO�WXǋ�лG���a�����*���7�N�M��R�8����R�Vf\���W8�pzq��y��I7>�C[�Y�V��T�����2I�c���by�?�}~:?V4�#�ۯ�o�4]EC��oS����yF�;cv�9R�Wx��"Z3|sl6�7�W�zK|Ƿ�E���?;�0A�
y>�����I��*����W�h���~ZE�;�����j�4����5t#�)Ғ���i�:���"��n�g�y��̝	��1����q:x3��^���0H�l�K+�zڭ�,�Qx����'��YS�Ra\�*,��z�����p<����j	�\��r!��t.kp\��:�`s�t�VO��#��2�y��Xu�<����B�⇈��S�N��:��
�X�:������ʼ�n
��gG}�-�PwbA��Bt�OT�9����<|�q)����Q�m^���� ��+#ZAhP�*<[:J|W����jQ�'��6U���i�oA��>�t��yg�n�s8M� ��D� �ug�"F9C�w���SI�5�_rv���D6`�%1�f����F%�(e ��Ld��GTK��%x�7�Ew��ߨ(�F���5��}��V=��2�j㰜��
w���P?+XI�)F|Br���
��k�9���xcsi�G���*�F�e�	���A�K����*�:�׎�p��Q)���,���[3��u��o�LF��E?zV�-%C1ty7J�+�R��ᇘ�2�I���ʗ�˫"�����N��#T�E ��İ�:p���Gn��(+�C?�=�W�Y�P�P�OL�0�i��:�vI�
�Pa���?�j׽Ұc�g̫?����ӘA�٘���㬨J�
O����'���kGs�@az�z�6/Kr��DЗ�0o��)[1]0xƛTۻ����n�b�yW'�?�-�͖߄�'��xXTʝ9�b5����o���>�M,���5)���/b�{�rJh6zP�}>2j+c�`��ג\1FH͝���~�����N��j�����T2��5 ��sC���0'_��� �l��J������I�pXdf6Uj>�T��Q�&Wf���Z�V�G4� ��ym��DɯrO�1�Q���a/2|n�q�����/�m�<��?��/��Vx
G�5+,z�^��\AS��!�$�Z�}�B.�`�ͤAF���G��ȢM���
���É�D)����E���l"Bu���u:h)F2�l�E�u�'��I�sXJ3�q6Se�&t^OY썾/I����g����..u<+���~sQ���;v�$�io`����,l�������%��|	�C�
;���G�$蟑��s&�5��Ϛ8���p�;�ONԊt� ���5�1�l� ���C�Y�Ҧ�#�����i�t���0�i0^��ae�Q5�_�Z�Zqo�N+�-0zU�ɯ����,��2 s�_{���o�f^�~~٬9j���A������Z�)�����1�S���DN��F����EȮ�^�:�yPh���uQTmMt�'�ئ���'�&y�4�/N�$w�]~�/<#g-�=+��TF�]��w0��V�k�I��ks�Y�d٩�F=j��4����c�f|]���iq�O7�yf�#����P|GOlMP�hfY�G"P�brt�ɪi��0���j��a���D�&�حD`�����ԞeF,�g�<D�Y�f��r
�g齅3��I�NT����w��YZZ&�CUvm������Ħ:��b�W���ek,*�.��eO�k�IP޳Dڿ1�f�'h~o���=��*lV�i����cUj�RP~πf����}�W��а^1:�dvKLE|:�h
��D�`�U�1�g->�;�vtk�sx���2b�?�/�A�FE��/@�l6��O'�q�{��7D�
[�܊{x���҄9�S�x���e����ttÈ��?�J�k`XV�����j� �	ȋDz��%�l�W�4]�d�_�,��)�A���<��5ds {��8D���Q�D���=W�!�� Չz%���NO��C�iHdM��[~��W��Am�6��Cb��Q<��Ǒ�Q_��C���i�x����(>��S��=�8���o�?�;�zb>� q!���"�W�D"P F����_���-���"lv%��wT͵X��I�ߖ���ە��]���q���D0�΁EQ�Yi�J ���X�a�zƹ��,�����j깂K(W�j�jw���_�\A@�e����ګ�ni˟�n���?�IJg����8�XC����#��A�l���27����Rf���_P]&�t.%�x}�CϤ���d#e�������-5#Ù�����D>p]��
:��~�� h��҇g�Se���G�B|6��ϲ�q��EW�D�	MP�Ţ�7!;����¥FbDȠķ��v�;���6dXx��e�X6�[N$��l�P�NCj}oyM��L3aA�����*�?p,j����&�sk������m��������I�� JW5���La����Kz1���&7Ŵ�����lt������&�k-bu�T� =
�+*��A� 5 Z�PRxF���vTZ�L/����@�
����R��a8 ��C"��P���-+��[p�w2�O\��û�n�SÉ�+�e3��<��1Sj�l̶�����%�1�������s$�d�=��Ýa�����w��T�����Y�/S�^p�XTgȵ�ǜ8��5Ε�4T��۳-�T�����XU?��s�t�m�!V�L��#�:��鐂��<= !{^��\0a�-�G�Wq�UL�"�U��6����o���<�X�ǧ+C�F�+�bi��g���q�k�-�chK�ۤa�}���&Eں������= +5��&��a��G.G��)(Ó�vg������ty�$f����V�߄Iy�!�Y/5�.�+]lԘ��=�pv,��p� r
�/e�i��G!C�0��x�ᕲ���W�0Ǻ��	�c�<���������x�8����ڱ�\��.�pg���/�:���؁�a���4��c�n�����qn�H�5�-����Bg/E�Su�~���JT/"��b:�-!Fl�AkFbz�8!�&m4P�������龹N�%W��H�2X��r��P�}HP���P]/%K:�5M�,�N���6��θ���l����V�������b�r�|#D���W�A'S��8���|�^����������nd�	�(MM�W�4�*���Z[fd��&9��	�H���6�+8�����ԉ%�[�>]�@�׌�Ʌ]�$G��5<*��D�p����.P�w�}�x5a���7���x${oE,��!��Ծ}�.��#��o7�QdC����*���֌��k\�T/:��ܸ�W��5��굝���^yF��z�����	l.^�r�3͢��cȪ��"�u�;��>�I$��t��d}�� �U޲i�O���"�M��n%_�0����pO�g���k�Y��7S/5��8)�� ěw�P�0���a��Sw�>�� ω��*�1Z����!����UX`��^|ɀ���ٶ 3[(-(����3��wc}4s}�tj� =���������KOP}����`� �w�-���I�� I�
`A��H��ZM�,+i�1�P"��QRi���,��)B~��E��Wt�ֲJ�|�M�^F�����E��p�\X�ZS`��%����x�S�ʿY����j�/��i���G����M��Anb:��o=�
�&�6 ��iAv	���<�{��*�v��K;�u�x�;�	�J���	Bg{��$Q�]�j�0�)�w�y?�����	����.���D�$�j�ƀG���?��{i	�H
�
��ͪ7uVא�^J�O��s������d�Ȧ}D[+$9��ҴCk��8��	�ߚ��aƚ�$�_�����Ƚ3R<������+Θj�p5ٜӓ�WPZ�m$��h^0D��U	�fW�q9َ����)��x�#�c�r�4p�dpn��N�A2�3|bU��+9	/�����>o��M
P��Ŋ��y@��oPdR����j����:�)��ǵ3)~gq�D�Ȩ<�3�^$��T�]dE���6��!*t�/^��G_���E���y�Ȗ��x�;���R�Q7YV�8��*K�+a��Q������Yd�g��>���g1��]N�\�4&�[�rm��ZE�xF���	���a��T��͏�Z�vx85�Ǫ瑜w�g���G$�f6k�pC� (���`���WQ����s�{71�ݥ~��KZ�o�Y�w�[P���˃٘�g'u� J�P�pbϾE��Ќ�,8Т6���mI���Yn6C�$��k�#iP�E�*<c���p0��icF���f��:�Z��#�"�5���`�ݪd�����1���D�qwYv|7��9;�x[�R�q��T�is:�4�Ň8Jі]�-���#E�r�d�oW�`n���4 �Y�I�Ml�C����nm������s�N.�?m�n >h���*�q�_Cl_��s���\�V�����K0��%`l�������-��g�]=y��-Ǽ�utx n����;�AD��\3��vX4TS�|y/�����0�S��Y�MZ�$�#�v���d���iY�����d�K����\ԩM%o�ן�K�v��A��=������{Wᄘ��`��{���g0�Wr�o8�o^�d��@�ŽaK���w���N�頻�j�����|�[��Y��k����Ei�j����j>*�Fh���]���;�m4Z���%�+��g~g�X�c{�=k4-���Ϭ}D���:X�3G�X�HH��܇�h1��c"(� ����L��!��c	��@��Ø�7�6��%����%	4>y ́Cِ�W��m �E���w������kg�½.���ې\��Iy-�。�[����~����D�eQ(_��x�͇���U�W\����4����W�L�eKT
�f��G�=��\t{f�)�O�"-Aa�mF��UE 9\N]�v���:���k�Z�nͽwH�1����c�睎l�f	�F 8��嫒�t�(��� ���Xe@ k�*�˻*N��'�
u1sD.U�s��c[p����/�?]pJ%�E��z�ј,���eZN��(.
�~�f�fV��Px�L�3���� ��	:����0��"�O)�/�L��9���c{Ƅ'��l�Q�% ��}�}*�����RW��V�'�2SAa�����-�1��Җ�	�G:���\F`���]�r:�v���m�A���n�u]��_�ڨs�m����~���gqd*coS'���o:���02:�7A6���&�Ch�d�GO_�hAW6��t�
�Rz�w�j�3S���72t�כ/���b��&-��e��8��$�?��G�H$�
��������UM�p����/�fP�1W�<n�i(�u\��\_7��H��>7p|"DB��m첢Ci�3�N1���4��~c��p2|��U��fbL����
;?�龌.���DG��Ɇ���DyKFZ�j�k��5�������,eW�"����v�RY'(L�֏Q�'��
�U���[�(U��]=$ַ�V�aJA5q�n+�����4E��\	%�"C"�dHاN���uk��b�e�ϋ[V��S��4r��D$����Dj�,Q��1˙W�����3z��4�<!�1�2���$�m'�8�OZ�ˈ�g8r�C��&B�I��kMAܑob۠;ׂ��J�{����_�w��e}b
b"i�
���{����s��[gF�@<+��������U1Tܓ�Y>�Y��3ȃ~�[�,(���
���~�>|"O��Ŧ������`2��r܈��c�5��Y3��je�^+�ՈR�E4L��,|�s��{TwEGȦ��P��{%���&��3Pi�
��ԠB�{!������p?З�l�R������ɵ;1����t�5/p�J��K����
�������_�Bd/>�K���+��Ʉ��b�ӑ������8�P�C6ǰ���D�s�2AE@���B��bjtp��ƍ:b[F���Lp��&c��}�R�T/z.&=���d�q7�����/-����-$�ZQ@oi��
F�5�Y��\(+y�2�o��
�_H:��' ��5���q��É�Z�w��W@p.��x���^Re�@�~��	��
6A�?�2O�{�V
MC�%��)�iO&��d�y_���TMw5���38�4�턃º���0vo'8����Wg��K�+��uRQK�Вਊ����j��#�
�Iō�����-M���s���H���C���t��5/�e�O"]RG�A/�^�"iꈇ�C�)̊���<06�m��5:�[N5ޫ�b?C�T�p�J���d�Q��L�@�db'� 9;�,�h�
�*�/�G���Дp�~
b=��>��eJA��ﲬ���� �_��6*�/�T����3��.T�3~LK�%<V6��_}�Fy���R�{,	@�ij`o���cľ8�z!^�1�|z���%>qkE�h.^�����PF��p����٪ &���qjm��TWt� �=����-K�
q^d�ư��Ƽ��x���I�c�5�|���m��'\�$TǑ&xG��`rV�U�H���F�Wi#��k�c�k�w��Р�V����;�Ǳ`� ��Y��u�:ʿ+��(S�H��h3(�G2��a��XJɓ�k0�4�9��-]� '��70 +أD7�5@t=����K��t���e�߹i�r�IB^& $=>޲��p���"�.pؖ�ȧFWW�%�;�;ji�6d�<��/L���Rv/���5��{"�?`1_>�'G,JV8[�|�����sPr�-[�Xb�ȵ����U��S�z��0m�ʶ��������ߪ�&�P�s�-��\��ܫ�{jఒ�ڬ�>�ԙ��� XW�U�W1._QK[|/�˰��}p��I4�Y�ͦ�5�0zJ[o���Sάu����gid�+��UK���L���X�^1����j�nX�X������|��k�ٻ�/��M0�p{��|���2'E����M���� q�^ÏPO���S̋`�k��H��'�e�aق��ӖFbJ)oS�����ٮA�B9�+�G{��4H�{���l�h1oe�%ye(|P�0'�9���jT����I���D��І�(�Yv~-9p�*����q�
}t��x:{a)Wr��*��&������&�}�ViH�;B�It)�N��U�>������|%2�p�᩶͜=�D�B�z��)��OH�5�@".O���D`��B'�?���0���Ys)<�5"��	�]�:���Cnp�Q��v�_���u�)]����q�����0R5��S5+��B�n;���3���Ct髟���<�si��a��f,��}�Dȍ�x1+�)��"b�����ص:@us���v���',��-1\f���}u�s�2s���_P�#½�tg	$ϫ�Bw2��Hձ�QZ�!�y<��K��C@W������i��6�X�$������La؁��f���ڶ��*Y��`�zW��+`�|��)��:�%�� ��צ�����ygk��p�݉on|e�C�iqʯ�׆�����֌2;�qc�eZ��&�{�J�l�bLns���|q�_�K���L�G�+�K5�[��Z�D��߯�p���o_��X���|;ԑ����J�n��>s]=�R�L�Ub�K�e������3�^�sT��C��&{=ǎr�_�!�I�K\%:���t�*B�JUA���m�(�{�lB�dF�:��Ǆ!y�sWK��a�B R"T���SX��%W/�ݮ�OW��,\Jكg{�0D�K�@o^���M���s�j_���5$�G�&M�4h�M�\�Hj�.+{E��;^X�^h��	
��2�Y���M�l�m�,{��吱Z������,/Uo�7
	#u���0�G�J¼&�]�r��+����M��l��h$ �P��,���:TiP�'Lu���x�O�J�(����s)�T8��(��|��7]��P��xl�{$�9g�e9�@>o#s�4)	�����dd&[�-}96�N��r�F�
�i나�z7V¼���<I�`H<笍rG�_�گg�֦;��r�QC=�}��1B�}��GՋ�GM��m{� ��.�;1t�p� ����Ӆj��v���j^�! ���L3*��sZ�>v�ƃ�e����������磳�ZP��^"HZ�����ǆ�v��6�l6�Ć}0�� �l�i=�u��_{>��6���T�Z�F%���:����U0��|*��1^�R��J���"���;)����%�̣sE��d�G��k��UZ:$s�����$�9��͍*H��Κ�ǩ�5�lS����⬵F,��}�o��-DrI�sPn��+/᭮�Y
݄�P�?�-��~� /�Q�G���t�ҋ0?���a�"��r2�BkJu��0��`B츬��6o��P9�4\hM�3ӷ++�b}c*�r(��l7c���J���͓���*f{��ϧ�μJǥ=6��Ҽ:����A��5�@7�{/=�[��,�O�#v����#bi��������!1�TU�*�KÚEh�ॠ��È��-�}ɗ槆o�s��<�؞�[�$�8 ��W�8�Z�d_�j2�F�*}�\"�C�=���T.��@����G+UQHMEoW�\ҡ6H��wwعh�h�����m��Q��1E�י��OV^��
��d-�
����O�وd�ÜYK��Ng~k��Z5f���+�;ܗ�ţ�fh��S'�A�ʙu�5��fu���*�s���^��&�s:����ƍ����6�:+̙{-b��I{iw�t|�O|J��ו)|�NQ�T�!��Cly�KAHV��9ҸUU��� I�ZF'�yę2�v��ؚ�V7T�-ؔ�#�F��,Sv��2b��	�O0R$�F����/M�#܂���fJ�v7:>���cц��A�ep��η�`���}hn��Ɗ�\'qq��-���"��_��}� �.���Y����&�t����C	^&�w��O���	z� ����O��Ύ���X`ԎD� �kB?4���������Hcl�Q8ty^�����5x�Ǳ�;wkU�ĳ\8���V�pɪG����,/���eS9J��a×v$�U�μl
�ʑ�3,vɨ'p6�˗�u4���%�u%��_��/(���E���Qއ'g�
�AEU�*��N�r�鷚���wB�,)H��CG��};-�|��0gB�.�����ݵ���WWt����GgH�+���Ā'���7�V�E~|h�f���{C=���1�
�KX��K>͒�ٌHb^4
Y��G ��#���0?^��S�#-�����Q��eF�0�C!��Q�l�!Q�����t�v��~�	���t.�)i����z�ڞڗ[1��!j�|���)<�ߧe�~w�utl�t�t�/��	#j�Q	K:��i^�0x/��/��#X8��I�K����{&��d���Df.�x,��IIM8�/""�@p��#f��i�\����,�z�<�d�"A��c�������W�9^_�]�P���;����rhs����,=��z��D�vC��1�=3J�c����A�N�m��f�#�̒:h�,R�FՍ�0%t���~i��q�.B�����7�ޤ�.6�s�i��W�W���������`c�}���8_e)|��+���*�m�����B �0)�|��WhX�`�U�ʆ-���V�l�
��,m��="ƺ�4m�T�R;�9�_e@�/,�ҝ��C�2j�.ܤg��>�ɒ0:��)�O���1�8�A2g��T��n�j�Yω/x���ƁHB��Q�ߪ�bVYKBp�Kwz�Y��M�P�#	k���a��q�7w�M8�:�:�B�ם�]�09� J�h񼦔l�Ԯ��E�U�wcYޓP� 9�!�꩙k���m�����:	|�~:q���"�}����a�R�Eh�?��%��}����0��ϾET�+�"��r�f�y"�du�Y8����Ų =��@�e�<��=�臘�&�R���bgq<�4?���Z�B��N�
��y9H靝�kM����F*���Y"�ܗ��	@�>�Rl[�g���^;�v��/U=�s��U�Y"��, �P�z$��o@	Zs�fg�<Ū�t���Y
�ᘕ���߲�J���'Y���0�*fB��o����l>0��,�=4�z������-��p�/u�8RVQn�A2u��
l�k��=C�y.�8rnp��0аx��c��Q����������G�9���2[íߡ�Ǖ������C���p���[,�A?�4���ف��S�Sݢ�Jn�z&,����I�6� ��|� �����%��͈��ݵ�,����O�����:D�� �I�������[x�ƹW 2T�S�%�����,��"Cm�C�"ŪF[���SfptG��x�9�+�j�S��/�u�p15f���5|)��t5���΀������@@WI�\��А�LN�_,@#4M 8�(o�@~�W��"�۠m�rTL��^�8:���r�a/����Mn0�Kk�m��P��G��:�э�ee�⺾b6����t�aꒉ�,K	�O���j��w��J`O�J~�}�t��B#)@����`pB`�@�I�3��\ �������z���a�㜈�����������9kL�j`����F^�zk����K6%���aI�]��A����r�R�q��ý_���ڼ
@{7�����\�R��.�3"��7f�Q��.�IEK�Eױ}�<{&;m�բz��'5V��D�`��� M�j+�$�
]�6��i�r��w��K3�s͈�� fԪQ��W����`�zS����W��i f" O?������ZO�u�y��1�8���Z���QO��<�t�%d�2'r�o�6������q��4�q�(t ����2 g���mD��Txz6VI��x�s��bm۷�^O�c7���@���C@�p�Qh$�	���a�+�ꄗ�g��Rց�+��O�
]�EҊS��ix8��S�`G��muu&{ �YR{��ͺВt���6�+fP!A���R�M#���������?Y V�m�޸���rD�+S�l���R�p�*��h���;y`��wI~��ІT����R�Ѱ#���d"��e���H:�C^�����#�w�&�?�ol/T�!>�z:�X�Af:JN
��V_���y_jk���;�����N*�$� Wz&qt�g�za܀?���LA�?��(��=��(ۤ,�I(:�N
��җX���҇���}���Xz��Z+�{�>#�����H��M��t1 ��T�F��E�E��J/e��'BF�펰�R�e�X/K��ơ�s��rOf�9{4�٤�P������5,��R�K'֭�tR�����GM�!b�L�5$�%Ə%�`��"}tr�n����)aS�������v��޲V]�8'�z@5��u��A�kT+���ݖ�Ԉ�b?\�P�\�]�7��SO�T�G����V�g%m<��e26�j��/껀���Pw�ćXWP�ҍ.0��E�5 �-Dcm��!��&ϣPrY���"p޸��;O>d��0zs�tv���k�����^�k�[H����\^v��E��$��b'��7۫m4�+#�N�5�5�>��R�j�>h �� E�בdL��#�n6�`��D��\�b4�X����%�n��T&x���"����J�w��f��gu�Iga1�����\��!�İ��r�9=/t�����X ��fJ�'���y=�)m���@�����7���Ԕ�ڌ^�Bu����:qDF��f�`:`\�p"����Q3ۋMH�4�۸�Y���x��9O|6|N�� �hfqa`�w�쒪J��1�%��/Jx�w$n���Vp���nQ���t��}z|]vM�q}�z�U�����R���GM��<��rs4A3k~7����ߑ���+N��)b��Z�\���<�N���������!Q
�S�$���]�lqv*��uv���ڍ̼r>5�2G�����#�M�m���^Z�~�}nh���)�4��R��z�.��6�5��*ۤ�=S���O�H&�5�g&:��k:��J�����`�V�ݕ���u��0͠�
�sVZ��sU
�J4_^U���p��2�������3�����<	p���3M�^6);��;q>����
��Z����(%6��`=����ģ�ֶ �[� C`�����/��X������$5�!9�]��2�~��-!y,��Q)��/���sH�}�������@HlXh�/�+��Z3���_<��B�OA��{$���8��&Bh����څ�"zc��n�ә��׻�Ҭf�lf	'�^��0_��z{���a&�&
�)�,��X�	��[v��y�T���J�&��-ۘR�7R|�^���*����Z|�T�3vr��4&t�iC��C;�E�H �$�f5�0R)��F
9?%qĊ��p\(9����}{���^�U|26i�X���zZ�=9R��W�>k�X��-�� ?'��j�����=���`�t���>�0M�<�������Si��4T�T��b �Z�|�0�I��h5Y
�&�z�#�tóA@���z����S�|���a�.0Z>�K��b@�y2T�#�<rV���3ތ ��mi��&S��ҧ+��|����}sx�{u(���^�\W05�&aʚk��őu�ˏ�?���Jʱ�����6���XIY��OS.��=�绁�`�Yr�����ʸ�2�Ot�O�n.�3��2�B
E�E4�1�7�&+�o4�cNQ9Üɼ�Pe��(�-rC��]�)��
	 �DϸϘ�@���ܹ��p,9��rnv?5�3J��Fl�� �}ɖ��@J�s1;�b�܌�|�?��(�]�����)DiO�2�TEĨ�q��>C���0�$��t5�q��X\xZ+D2-|����,�L� W�$"#'��0�g�tuRgK#�Q�6^�ka̒���r$��F""�R�^����t+��`d@�?�J�Oo ƪ۟���F��������`�VWܟ-�l9s�xn�bu|>b�PDb!�#6�1���r�j#�� "hY��4͛��>p���N��abPb �"C땡��k�ݩ�Z��� ����I؟�E���r�'�u�{��l���@;	A� ���c�^��tɫNT���e�t�B�Bt��+h=ǒ}z�8:>'��O����2NUV�/�����:~!�1�
ZT�]4/���L:��b���Ð��0�m��%Q����|���Â��T���	C6�ؗ,�,�qO		�P._U��mB�ZWd�Ԯ�#z�X�0�I�5�o���x��4Գ��Y u����y�20�����yI�P�Q9�#�6�19����pk���e��Q@����������"(`?T��S��Mdq]
���x���[��5g���<��}Hw�^M�WqF�_~X:  -�|g�,^�K?�32L�W�R��ME^@��p�u�t�N������ǅ��T��K�!�ɂ��h������:�egR�����b�&��=eI�.��X����3��O,F�-�[��m���Z�����k�6�UeD�jhoz;V��c����i�u��Ǧ:I�	&3�;��&���o�M�/$�6���ё��j�QX�J�J4k�BG�O��Rg�s7h���r�����Qꅮ��s�&�%��@cAS���Np�D���~�S�y�
�j{�g���j�5;}L���j�0�ytQKN�OU&�]�-Ol�;�\J�wLٺ+3 0�2�� ��>y��13�˴@z�uȠ
9�FK L��Vf�O�kiQ����"���Q�u����5Xܙ�IC�$H�p��01p�Qy�ݺ�mO�ghi��s͂g��q�Ȳחw��Y�K8������W��b��9xw\��&.����:�l?���V�w���(�mӜ2��w��?�?������ �Dli4��E����!���Um��m(\TT��=\SY�:C��:�f��b��u����f�Y��Y2��U�x̝.��<ËX$��͉��N��!(�ķ�Q�?�'����I� {��`Dd�qivVg���G�Wvo��S��,�;M'Zn�P�b�����Fi;�u��\���W���92�m�f�!���%ð���߰�1s*�����4O/�#��0�7뿙�C�5
Ҥ��+��U�ƁE���U.�O��yj�?X휀��GxeN��k4�\	�ؼ!ASM�l�f~U�9�*���űa?f%D����- �������J�E�s�H־�b(ϠlQc�$�G�;��.kԋ�܂��h��꣯�
"iFR�  �0!�B~L���m �;���p���ǡ0RL%qOX��~r0�m^�[��l��쟓E����8�f9m)��rZ<c��[���l:DLf����=����jL��[7��	��kdh�6���J#�����oq��0�Le)/�	�9�ݱ�����A�(�/`���A���o��
�H���O	c���͵���#֜�{Ձ(�r�/b�f������|���@�JK�J蘝��w;Gq ��&z��:^�e�!&YW�~c/���<TCMn_2�z���G?�Q�_�~kF�����!�t�*y�yR�+���i`��a���^�1��t%'P{��l��Ϙ�ϋS%��/�+����F�V�"ؽu��I_�O�v\�F#�a9��.�(9�L)5<�$�O�X�*�[t��i�6#.-AB��qI�z��]�|	7���q���L�����~�P�Zu�#�;�ɱ+ץn�#����`��H� ;^*�˧?�'�z�D�d�� �ض
F5[�����/˪�v��(�J�#8'��_/���Ao3����ٗ���L�����m�(�(g=��$�
��עuL$�D qM�"@`��*m㖃WT�+�{��d��.�d�E�/�����(��X��)C1;ϞQ�wT)V�(hk!u���]���R�k7 ��C-b�s"K$h}%Z�Zآ�k2H>�י�jd�s�_�ZI8�W>%<� ����6���Ŕ<�^�`�0��Qo�Sڹҳ�Ye#N�tD!�g�)f+�R|Hv[�ޢ���-��I�2,�5���h���|��~�.�9ѿ/����uK.��6�r^7r�v�ϸ�(FK��l"��l���$Y����Orf�)��Dj�i�^J�!�(�`�*u[�y�@e5�. oh��e��H0�n�������4<m�27"s�r��5���2W�Z�k�S����^^�j��ֹ�zE T������b�-s�:I�4��.ȶ
j�@���H�g��SV��|�¦�F_q���>LD���~{��Qv/�&F��L�$Pli���H�gq
�����tv�i�ΰ�j�N#��s���}�]�?.��>�kMl6��L��T����V��C�G�W6=W���T&51�6�+�,o֔�������&܄v�3��G��y����	� �79�E<@�#z�Q����`�6Ә��Gn���Z�k��/`m6f�6*^�*
)9����w:e�q�&e:�؁��kπQ��G|�@JF�W%���ʖ�l�WP)x�M?��i�ܽ �����x㪆Ƈ�u��腑�:�����\y���Z�ӿ��ya��ɡ�|H�<�&0�1	g�z�0�k�mVȐ!ݥY�'��Co�W��J�B��L {�>w��_m��Z�YH��^ ź��>���YԂ}¬ �����>��~(�(Kt`��^ۿ�>��O<V����l7�,��]+ M���q��0�n���`Y�ӥ(�(0SR�QL6H��H�c���g$��s���q���ɤ3� �b�md�S�}�%C9 s����mJ,wV�8KT,�7'h3(V�.6� #rP-*�=F҃8�M,��
�ڑ�o[E�!}�,¦D�x#e��$��NIԫ��!5!����MÕk����v�:���p4<��d�2���2 U]�^�;;X׋����#~�h��&e��%H囝�U�s{�F�={l�DVI�73�a=`-��������1<�����F��������B�t�;t��B nUK�^�An����Q���x���I��A=�`�$��q���x^�>�ݠ)��(����ބ��C����g ��f�;q�S���ߙ�v��=���KC�iCd_B��i~9�u}�84�!lrX�Mq�Y?�A�K>��kXm0r��xy��p����P�D�J߱�EՔ�m��ƣ��| c)ޛa�������J"��u^[��o��l�f�u�v��+�dE��|�a$��ꒄ�{�Z��/׀j+$j""��1][�^_�,�G�8�,���q��h�r0��/�0��D*�
�@3�2�G�ɍp�\�� #�h���KK�g��_�^���]�jus�8�Xl]���zKw�������|���i�p�uj��b�j��I��Bʌ���*K̹��
լ85�������.��A6��<Bg[���$a��5d�Q�l^:�/J��V��=W��F�|@�)g��6����X#�����Ⱈύ��T��(V?�0�������������;?b����C�d��u����B��GT��n��� fb�j���<�ƣ�������eWX
ua|�]"��w�u�h���q�
?��H�(@H� ���k��auh��6�^]��L�po5Yl��Z=b�y �}����q}�հ�q�0��SB1����HU�����3������cq���XS����ie9DL����]]��M���ЧxH�m&"[f��pnB��F���Th?�|O���E�ۓ�No����xn���s������[��R�٪ڔ u����++"�<c\;J��~&����fA�$f:�f�-O�EB���P����۷t�T�e���`ɞ]n��Rg��Q.����R��#��"}���׏��R��ݕ��Ӥ�ַ��2�"o����,����W���8w�Rj@R���AxU(����U}���9Lq���z�G��@6 �${��j�
��;���p�r�>?^n����f�1H]������(���!�_���sN�ʑ
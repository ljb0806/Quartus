-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kTwoRWo2CC1iKoVwUivKh/GDIiLXJE3sg1TD7ElSJalBAi4Cg1LeD8tcA6yfN8kH4yzeuE+/4Tiz
mdmXqv5hyCR0RZ3kKJVDb0hSsU0GQhfUPzPC230I7zonewm1eRk2fFkkcGhRMTdkmMDxu58VK/wt
WsYrjHmdMkL104QqW4b0co1V6Cqptn2t6rzYfNqo8TKUAI73WpX4SG/71N52HkYBuWEe7jM5ddKy
UAUi/OmCpxenQGj96CMCL49FiPkilaCijsgMvETvo+9iZfMnM5dhPdKksNPeh3G/8xDhxRbhzLmU
KdwotYwsfbUUAH9PQ11zkrckENA9cjzGNNFIOQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6208)
`protect data_block
tYL2X/ehFof5hkyJvhriXrvekS2weBUzVynOe7nejrrptt0ozbQdXE9Kx0j08pEJHGnwIfLAWGXQ
2w3dbqik6W3qILwFG+KqNLdLPGqOvO5akTHdI8jXITPZS3KFjnf21UnFkEC7y+q5M3L5fWWxfVQ4
j2Y6ZTiUgBxW0Ir9eMRqiLDFkoGP9o72srpbUNL9RkX9EIbwSW7MRvzQxgUuUf40t7jnTDSzV/HU
KyiwN7Pfi2brRkSmUEj08O5yD469H4YEVNORBRm1OgHGoxW+k+6G8tDI/hL7hZag1/KZUOtKZSGk
/s9pCncbovmxlgk3lNxywE2CelJDLiSiK4pX3QZWhRM5qp5VkR9vo+KmDBrE7GOOJ1Or26RuOdCt
pIrRTFRhQDUSqQSKH+KHVhRu87fLM7tGOmE1zODgC5UXpKr0WwBKoI5HENosIr+chlSVo2v2Xq0c
Z81jCGOFqTnEqFneIPiJwj5Zdd+1weYyf3vOT2EiqzLge91tejrbwjHdNN59ffT8n8XN+x/JqrUH
EVSNjH224ZF6T4A7dGmwCR9UclNVBA7IZE3nK6/Tf+ZRG9bTFJ8PZTn6gCHPICHlHv4wUSU6PTYD
rtw0QtxlWCGAqOsPXonbpe4bQDDFlfk+0N4/IdIFbnNf6vKy+jQ5RL015iZ1ARsQrEYnn+BuWvyc
db32VbDkOOQFqtjA3i6m7g/Zj5Oe5mBxyhYH3bYPXXrwBYsMyNhBtiynU3rF+HmIX0a+DHssJ+GY
Y1V0TX0vsCkVCZIzE9PxyOmI7Y56NgFD4lPJs6J2JVBDihoyBKTpao/SIeIK7ERYfjQIIljR+VkE
5gjeziZPYxHTETDORd5h3nWT3l+e7nSLWSmA4H+f6STu+I+Thz+21JCFV1N/R1/YHcHGu1z6ngVM
u12XEDZnNiKcASNEHvg4phMXCrPGUgq0OwLXko/Cm3jqurDvcTJzTlB0VhgUOMeH9KhQjbO+w28j
RlBw38i0IWWcJViQp0VvxNjRH9bWo6XXbcC8xyEqpkm5vaOOtK+DyniY3PUJJT/caYOqsdBFSChY
umsauS8HLioLVH466/9faZ1v36EfUOck/OnzLKU+iWsx74HCjPUlKW4dZj6l0WU9FSV0dmeTBHFS
kSUAYD7cWS7YrlEwMdqDcF8TKGgb0VjMlt+echS4oKa10ZswrWXaJPfxXZfyeKNVvT+DwEScIO7p
QOnej5Nlv9sogBamcAaNH/waZ9jBmyX532JtCfuOItES9ZZ031q2YLrwdl0Nz7XcQZqaFer+Rnsu
q/qPFYjq1+mGZlpaY4hesCcbwUCiwjPz4Siy3LcOmlrXSW1L73ei+0d7xkT3mLjsX/YEOsBP8hJs
z/G6BKvx0K0ou70m4IgfBvbk3g+jvsAU3lU3bbItCFlTJpn7nn4/tq2yT+CXEcx8R/L6sMACeY0z
wyBInLG7K2Mv97aLs321dhv4J0HU/zudWW4lPqkgkMkiAb8ZZBCaZWNyqBrNSl+QWqtDb4y2JFKM
jUPNYilanAnxnuVvvNbWEokcfWwFkbNiq77U8i2C3IKv7gXbQVvA1oU8g4cAFI/+5MXMSJqGddr4
b7Kf139rEj9CclPmcKIVlL91YIc/prMsuBw9fbdkr2KEL0HyaNB/Jo+j+W/gcudFGfKEpPcqQWde
Mr9MMmFEDWdckF0hWfPFvFTm22P4JJEShgtH0K5xeQXOfKQeXGomL/ZY6zwRQaELV6QPWEAusPmX
P5RJq4yEQWXlvaAWFHSKdDfJmlIrsQ2H/oKOxzkMhBZCRXWTftrH+eYyJjWJ+ZmEIVZhdEe7sw1H
HE2dCeCJ9I3fxg+wpP5twJRqFTFhfZWVUg09kKwP/oM60KlFBmTFlckdJcE3INtxd0YnMtReVt2I
jJw4OmOjIZvKvq78wtrCW/Eg88vi7Q7YuH/dG0YwsgWAu7Ndm9rwBNoCQEWpjtjrg745D0E34g6n
2EEka3Yw8wD5gO4kb4q1CwnfQCbk+wxN/nZ7R7LmHEw7VwO+/fNAzXmcxWOmIMLqKR0G8HAey1jU
gxX7KvXcEw4SPgjhRbeWv1T5edPGNYVRiy3suBjXLv8NwTBcv9DCveTMTyYtjb3BBt3cbzmWi6wE
pS/Jyk3KfbU/payknLS7Qw5R1eJ5M2E947FxwQGOAaz+w+E4gdQEbRs20VfZ48j12tEoRwRXrh1N
Pl4PpcIcbq4736QjsqoFekdKxlpabyndAZYPVgUIH2EcWgG2fDqKzWB3jFshw0QpjTr4JchFBpBG
KyZKWYsmejuNJwvLG4a05RjQMoLHbqUUUJQbF9PvJRniO83yQF20x6ZnW8EIiydVtHZjZ//5SrQW
MnnIMF3Fk3fs/AIZuf7WT3pYTvRIB5XH3LPzISvlEquoH0Fgie5vOcB34EsRy8Bon5pzLbyDQWyM
UZFFXxh3qT38MUKsBblNexMmZ7K0DAQ9JQMo0MhOGM5UVNZIT0T2vfXs8aRlTBSGFy4o8KpHoMzT
yU9jWOsZBRJrs7rJhrTUHHTp/jWMLziYdfnUDSZHA9MpzrMYtvl6ZLTYhG85E48r+CVSTiN1B+Cj
qJcdSX4jn1JIlRsq++aI7ukXDgQ+/h7X8/5XS2CQGT/P/cpluTXGnmqCpa3+yV6dsxny03VPBa51
UEvnSsrV27RWaNEo7wy3VyIwnuFAmzqVvkl2zIl49ldSiirLb3X2nDHkg6rzOSSqYNcb3uV1+a3T
I4HkiEnmF4njsZDXmyvZYo9ueHEidigfk0JZXLyZPFUQNyFv1hJxSH9kCLZmr2EaBEV3L7HpzFoc
cbfDveum1CbF0pLCFleNJK6T91aCYHNnnmc7Q1eC7kFnmJRolJoeNuXAgWz2dZlAcE/oesA8xZLL
wCiMcXnu8JfZD7ooGhNeWC+Gy8Zd9NRmTmmMr6M+VAKeWv74WBh+rps2vCHo9hQNXZ0wayOj351J
Bp0DZl4Y/2XoG4XZif4gatBFUBPKvZhK1ATlJ8OvtYwDN1QeA/Gahzgkaxk60x3ltfa2gpJdgGnN
BKazy5OHMg9Q5Hg+z5aj5NqyjMgiXH0uRPARpjFnalmEkWVmlkijXPrAsTzoIv/+EFu22qPgSDuS
oXGva8lTEbj8hQ6ItboGuaGf1Tc+w4HqxSdag1nkQ/xHK94SFBcjoV/q/aOfFMB6chST9uVGtJP9
eHA4hjteBggN0PpOt8f3dSpJeiIMqNDNDuYQk++RW4LgVdi+sEZrPx0rjwSDOzCYkxB3wbC153VB
TSdMyWWsELrYS+SFfFARRxFv+8241zuRn5HN6ytJrMRmqYreRUeIiUw/MwsmWLAYhjAiinBpO5YB
9xekB7E/9NVK8PFsmargGS7kBWxkKUAhFcQYxE8E/1xYpF8rEKDur98Xk81TkXUMjmMFy/ndLQsq
4XCMhi/pe1RYhTvQvsgjXg1JBaf7JeW4lCdLD6Oo25RrvRFTBOmp3V1LaxxqnGC/XAgobaX72QQU
LY6SQ9tI/rwjzdNEEMhTKWxT2E2uoiEi36016wW1TsptXhSFHKP9Gxewmwq6dhgW+rhePHc0vuTE
becY2gsF70xja2RXP7hZuKrtODHI5L/UGpOl8OESuwyVv3C/kxGk8odwXi0gF9IoxYqVxr78kl5W
HwDq5C9+9ykrbhp3gxMRxVSLFzk9Wsm/kqCiQXc6+9t1Sxteac4Uw7/xA1rEf88ldfT3hjHLD+Ml
i9h4ycr+BGKBDBB5LYMooQTbqle3AYokoCwfoRjki5jI60d3EP4Mh8EUXS2BbOC7K3KZNBbpVTXJ
R87CnTcDNMwtoiiF7k55JIV/tS5rOdJnK9HEgXTe/8WQHMOfqoSB8wBo2pWx4lHeei5kZU7jyzPB
Ug3o2Lk0Dm+4D2C2tF0tft9m2W/LvCX6oZASM5jjg3xyYYHhxgTSwpOCyKBVfKkWS9x3+2L6UkoD
BjsMQ5Nmkiswa5t4IIlVMT+8ij40eVAivNFjEIpZ3T9p4CgFB0AecmiLS6QgmqOm2vXl47p3Z2JT
wmzc0eTHhKIuxh4S95ra8ZD3UKsn00lGVqnR0RMsZVyZcip11iL06NSUCgl6J5aFofaJMJ1OUE5X
ubEUcN/L7qBhrIiP86iVOAbq/PrXL0dWy5BjJ9mc7iTkXccdEEBZBH8+eRyaJ0ONoVhdLIQrFNea
V79GyCcovbj1rpyRi6fIjsg+5sV+Ow3bt1L/mvaJrkIxIXFDvDjyCUkhSY0t4Udany+zpvp6VZrL
4HjmbMZtnUkGGzurPPZCjSfJHexqMbLAkPyPcnIKqwZkaxdVMJy+sZ3jCVoHFN8+ngVe1nLjtQ8J
w1CJGF3O8Lrwv6ryGNd5HYA2NX3JdjIoeia6loWXOxGvH+FsTv+aHqzgomIjH4ZDfYlmYmjuAJwP
hwxK4WRLVMQrX5X73NIlqigQa/5sRnys7ff87+uPOmX3fFqdn7S/T7uHKZssffBexHUxPalCGBCn
pIQBZiyuqsJi4lhK72qjYGYGFGexfIAWyI6Tb+Rj/LCcg6GUZAzW1U00IV4Q7SAvMgMi7Pt4qt2u
cMcYCZo3unj6e7EGrPqkHqmiFFXHwYESkm52DgeKSpNlURaKBKo9JMzyRdmyKaS9Qc3ELI0MwUI5
gfBQ6LxqZovZtb0nk/RiN3LGfQ6QkcGwkhwT+LUY8O1C/W3ngHdWstif4o2L9K0H3006xqi6CebW
RecgW/3O6O9ZVIab3aZLRTJ4OOYHTn5R4FO+aslkmWF0PDe3HJcX2Im0N8K2H2soR3QLaPUahKek
YzKNJxUBXWrVRR+CB5xVS5vhOKCbw4WIafgOy9hGip9LKlQKziyaE/kXAv65YwCSdl5qFcClyh5i
uFr+aI/NTUUN0fZK/RimI3K8Q+qxijsI9hF4KRG2rg4gHiyxiE3smSagh5wUMyF6/wkIusZsGR5n
klEtLqF0kg8mxLRxxnnOIThDW1uDcTDuG2Bt6A1FnoZ0vX83zssTbH4JmJtPlOtWNZXmKXkOT9ls
oqsHKk/xeNvIyUHZF3FpNd85Ud0KCo/BieZsSfPbq6BmrojG6e4fuMLvmHyloCFMSYJiJotJHgFY
hjQ5SJctIg6045EPpw4nc82H3NcKS+5QOiVZFs0+Xu1WVnm/TSiUK/q4b52ewhK6jeYit4CdLcyJ
/iy28Gz8OOhXrmWGKhsYgvlmTQLkb0VsHlU9LDZHsrOelMsF6wPs/z2G/tyi4lfs9hVWI0JlRJYC
hEI92QnnRPgVHmS4bGwbmjpPObcKPhNBTMXOWkJu4OIadKfxuRk9hlKt0oIjWjiU8rWR+GUCutfM
H7knM4ArGnpWpmEM7/izRYqZimzfjroeSYgmEiLjiMs6FoB4hpZgYLOUXSkDkHCXewZF7rrAUfbG
+8K++USOYecNxRNSb6vM6LbemwVeBfve2ntlZmIW27SyE9JophYQ2yNp0qhkrePpwW08Af01n30g
KKxYLS2FjcCFLEm+W93q4Bne8EXyEpb++er2FAkPsaMy+BHyr0ubHQJRmuZTY9QlzB5fOPPbF7E/
Cj8q73FFJCvkN5r5Y7/IuCpwtbJST1wGyo1grISVSJ7RjAVV+bsb4Zl7aQLDBU/7l5Vr/SQbOZBW
rCbrctTUGFCwHoQns3tT1SzTWewGM5Mc9drIM24+PTJi2xmpxojhOwXVLlMfPYRMFt2feoXOFfJR
rbj8wu/KeE6PDLhH8RlnhlmcBxIr1FECR2vIvEkD/zTchBla99UZnLDZPZId9/i0WfWOw4tj8eva
mm7LKDtrjHTvnPWSaeqJUy7DBZAvL/GHq23VcApOdmi72hytpcBWJ2EGVVb9BZAbc0I4Q/lBtjvO
vOyfBNA/gv+pLxIhY6F7vH5oPrUZKrqNQgY32aGl+mvxHVEJWcmgdNkZn9RUm63rT7yG1ksB4kOD
LRldi+WU2K+tMe55VmLDLoMFTISRa2yMRzmDHJZkem5RVW8pt5QzJQhpivyaTOvYj7lI3qpV1df1
2nHjF3lPY05C0HjpG23hcbuhHjr5WlD5PgXHFoTFstmxlnI3ltJ3niIn6sDcSsEEFggGKXCu567F
/TVD1/iGQ8/C9Ktu2GLOcgkqsrjXARs/7ew3F5v3UB6pEf1cFT/Rh7tOk9jLYQFYQodD4ZKVDSS8
Bu+7q3a5VAaBCvr/cyGC4SbFpEt8GkLIW2oknBmdBxO5pFCIhGGHSjbI0V8td+yIbuXkLOXrldnR
k+GKI8Uuak7ObfCJNOyasJXStAsmTov5wpmMCDZiq0i4TXQa5qyTCZ41aBMvUKIdRztoO0DxxHYd
R8zSbv+jQUy5u0+yKwvUVdvj+KdDsK3gv6eew3hQz9Drhge2Dpin3dRNTbulMuJTVZ7RV6iJhUdk
t/uPl6QWbCQT3AiOy0ZGRZQJRxwEPrIVzCEzsQJRB9VJww81MEY//Kmb8Nxj9L7N+4XFXPELAYp7
igsI/v34g9LdmJlMeAvkk/6xz/dL1nNunXMMslZA0ywvADa6vNQ2XFqQbOIQtdhZHA1RDYH3KSss
LWCRf2LCVqUVkS3R6dLkxQaoLn5URfbpww9z7y21VBOcKa8B1Cx/5/eXA3ID8CBrAjalinSLwe5W
3mQqngvlSITUdwliJKkZtGCIPu61cLAm+MzCXSVJCZY3MAiCGW5xGMzYhNNEoJUY733TvhxCVaLz
hQ+ctYD/s1Xv9UR/mZCEOfeIQip0M2wXH942EDyDyTeIvyF/u/6OjhXi3QuziyCURstdAizr9JuB
deAgI4YxLWXMYKBj/1xaD3AJuGZYn4j24hi9V3XMVYXkMHrT5XcQ4XyS01ZpQTkK30ogP2IGjTVh
N3puUEEy6m5aT7u7gzJcGxt6twWdDZ5qh3PH88Mu65D+vUwuKBl/87Dp/oL40xUifzfMlFylkgxA
36ShJ43ZAlbbhukGjy83yaEEFgrww0TcoYIsjgl7JYvOZh0FgVtai0QMUq9Liavvn+n8y9kU9xzt
m3JS/fihaSbG9q1gDnMNt3frB2ty2Rc3k+I8dIC8CtVLPPzLQHUMDYryuUWzVj2DUr44jvusLBuX
uk8pfM0T9CD9ugj4lZ8VBkMhrH7xSFDCG6bZt0zBqdFMi4hUW5lvVuypiCFSA7bPOMnsDh8MoSQn
qIIUu3GBx9H12UBNersDv539eEr65E5Lv1Aw7cRVaDu+E1WgAUnNwjwXmOh5bo9txm/iECHmjbtO
uiaetoWGoQEvZt/usErSTUF7Ak+gV1/OXmxVF3UB1z6N3CUbXxG71AE/7S+WtBqCOI7n2Cc/880r
fJjgQ3guhipj+uHsF0tdgd2RpgKoXWhkPJyt29JFDCd+g/D7C2zotEyYJu24TAsrWLWH1YmM3cOq
EP+pxHFuIIBTa73JZ8IP5RH6M1o4KKXY07ZLVGnd7FXpKbSfr+hotuzWIWrDXF/4oTYdw6h6JLWt
5ZsYaKlMgeE10UDa5PvT2lIcc6FCxvf0H4RLNmiyreFYhCwS5Wc1QtxBU1LDsbl+GSGEqtkPYMJL
HLIr+Zk9LPnoUJ7b2Cs2yU2Xe3a/s2ELQjBXQlVQAh7BRONcggqFy50eHijkuRM5IuLH7Lxt12+y
o2LvmZr/xpAcaS6khY0nRfTnT+TkJmfWyHrBUP+qDmahgWDcuSObcP2V4Md0/DoAXwxYc/eyN39C
UFwcnKYEFnjN8VgkSCmcaGPXPmG8VhP6tpaM5VzsDtz7ieE8RPeOY7alo7W3mYPXDV1al3WB6Q+J
YlQaA8NUnGCxEGa/L5kE7aJkANc0Svl+CMYFZgvjc+n+kAyFNxRjeWdg1VoNc5+4sZYrUoQdpZeI
5mRlKXODGKabfRvlTczbpCmGCZtkObR64PfgShDbXLCQGCukM86SRpjCble/Ibrm880ZABfnBP3T
wLKW4uWRSzkHSNCtXjNzMlcVY5iasgkty6zTY6jAodKJNhcZYfdEpxckHz28/qmg8RS4zsNXWIi3
XFWvUBzIb3RQ7WhfiUERPu1GGoLSti7zczdEXa1ZmNGtrR5E/pN02/AyL0EybNf6PvKxRZ0RCoim
FaPwk8tYN4UoUtk5BMF3j6oHl+NN3WWl+I5cxNr0cqwM4s7a8zQZ7clzgPNAZhOSx4238DQlfHy2
63K6yM4vK7Q9hXMy22BIoR4ydnx9n8L4OkQQY3TagkeAWoUW8IYAPBJ/F7C6npVZYBZayF/J2d/q
mSZKIiROif/bVLMrbu/lzk8jI1NJSyHxTL9hW0w96C/criCpA1pmyApcS2lhw8jROr7zTg==
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rxFUvTE4tRLPFvt3N/9EtZyGaw28oszmausBGxzr0Rr+CJEY6PxOH4QWW3EfDgwZxM/cOUO59lHU
k5PRvtRJp7D7trqmZqxv1DsQpwTt0ucSCDFJUS7PLNW2YwMGZ7R5Hsadw1j/ur9o5XU3EWhO/xSH
MYvvNrz0alfSLxREzXW45dpanNwD8vLBlmeuMmGG1QVeRbVQEyt1ZzkgToA0bYXsTrbccOKlphBe
N+zWGUKc0NOBNy+77gQI/FcP36nBU9PM6R8uqEtTKQhWi6nB0/kKbMBEDT+KE6/M8NdEGZPzLZ4O
MeSDmoaxH+jUyDVjJAOr1z4OFi+dtyv8NdBuaQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11952)
`protect data_block
cj9cZnWsv5tsjXsRrDz9apmY/o/tj3OFqqgF70e/L7HXO/Oine/k22RZ6Uy2gR/kOMKOVb1FYmNn
1+5+1qxB3Jztg7LFiwQAvEV3AweEtQI+uht4rs4PWgej8G192N5GB+912gxAq612dI1K87UVLF5H
5VtMw8RIbOznSgzUFjt3h6HBEGuFnOPyyXu+waxKr2dKbqI3y2J189q4ELxWfzCHUKWYfq1dESU8
m1H9q3iU0kbKBdT2KNd4zmqnzC0vswLTrBm54iEtsCEZ8Zy/59JZBWJzTNx1EUym7lw+If/I0O/c
tVehaiMA6p2kuwrYSx8ZXavgEOx25VUjrkYaZBnq+Gv726SwWDFXSZhmHhIYxFap4OTAv1UEjT6j
hCXdJtoKZuphtLH9oIYnFHomyG+NX9u8cw5jru49bNdeddOgTnDD+h8l4fUesLd8gr3C574AX6JP
VizV3oaYY1tZ7hm/MaJGeTJ0NXMA41ocvYZ/S33zogbbTPbV70eOGOgwmb+ZqPYRybQe6oeH3GGh
y2w9i9gCOaw5ALM73CuBC6CnWM9V5c1pvGPPMPu6G+Tw5r4Wpg4bVwXKsWKW1XxGsODtnsFr//Jy
RDlPv5BBH5ij0gm5YyWE48j/V6GVADSQIJpHHIcE1x/RAiJQRQF2nb6+46jchT1DklR/1grU4OCJ
BXCzt6BnmBxekv9uphr7Ki/Jr5eK8OeMwMhn4CyoPvXM/isjC0wx1LwaFX8FIu9OjaDW06/RGKt/
6eQ6GtkoeZfGKDOjH2YdeccTDnGlmbDe8q46Er+HGN7RwbcEWplKiGrKUYio8KT08s0qnM+Btlsw
c1tO64k/0IvFsjqnHDTWkSARh+zKp/y4AbRr3T/hCS7RGrXFnfpKhPQZgtxR5+qss/zq7k6uvxBc
gvkPhyY5s4vpnCmJ8hdTslRIEt5vynEM8VhVyY4+FCkOjA4fwGPoSlHKoiOoL1WXjUYVVD5fYUE+
gi5Te4KOfdOKMpWvtHIy+88O/A3r55LBdYVJWQksft7IRV3F06ze9hEZAPogYlPVzGFSI9EOBdtF
9FcDtr5qX8xKW+4DHU+4n5HJFUmS+xuQk9ZjB7hUCmAO+q7efLyyv2JVEvxdtPq0oZEio458Dbma
D9S/R9R9Kx+GqmsBIwZei8wr0fx/Q9B9L6aKzkScceqnndtwjyMujhcB+9liDSGeUUsMQwodG44W
C+pKmNCB9RI02S1Mh5b6EzzTmcYqjSQgSJ0dkssop8g06qytZhgRIWrSdjNYhfbsAR+aKIMYt9jc
MOW+ehmZhOBBGhxvO/de4ewbrfTWuVy03So0vhVVADnwC6Oi6C4U+HO/9cdTe4f8wovqplC5gczp
B7/W7DcDi8Wx+5oMD05T+GSG/iVC8Ga7TIaQQWSz3ShG6qNt0yd9buCwkLUKY6LFretItv4uXrN8
21457FZtXwv9t9Pp5WZGM/AWvEkHRTPcBSnQeCQ86p2TWyYhZSpKO+RgbJF59HT302o4CuLSvYm6
3wbniFc8KvrVa8ce1a0qnfrMR/ujSP1ACwvHVPPswu490DF87k6TtFqyPwsjAtfP6QvWOLTbQYId
bxR0hXaR7DruCu1VZdJGD7HJZzp79HJOPM7AYgSeXkkgAufoqgH6d4VZhfP5kLRtmSnov5Xs8Anc
UUgJ72PnO3PeagT4EjV7T4SUw144uo1p9cZux7tbl8ckVQYALAOYpCc8tf8gL+KqU5KwiR+6EjOa
M6iHvvLsm6r/KfE3N4K+zH4w3WQCfuR0qwlnT29zZNQoOBEwASEtBqT2SAtuBlsWYyqvBdivk5I5
YqkWG3CxCJGiimx3tXyKRMFjTONt4tw08UkxsVub4WVDsfehGxwFlACzv2ddxNufhEGGNcGyYfRh
BRsGl7XNxMXE2jxJURwuaModqTW5vqlecQif0hC3DJGyoSg/LZYr+NXSjiFuJmQg5ZZ5hnQEyGcM
pPh3qPq//V5o8ibJ3CFa9YSezbpPn8dowE/dTql9YxjH/7kEYGGn3zXBwmu2H9goce+0iKTe8nXm
Nlzpk3V5XMJdmZmKX9gGJ0Wij9fj7z4/zg7j900YVhjxgcLgRtv9wdui8MgtVvK1yZXO4pEj3LGd
FmGS3xiVLYXgVGR6JSRFQ+2INld4NRdp9ZecYbVakjVm7Es0vNJbA3Qb7UAd/Tvo+FNZIB3JAhXg
w8IbMlI+wflw2kVTitPf41GLYOelR6jcQXcMETb92cPb6ZoGozz18xcQG7jVUncVwJjxCaY+ngsD
ZQwpY2Cuz3XpVIDphRcmL1KwjMAt64O/SdwZm5uOWVJIadoXE1dEgjYhlEWOX0EbGyaR75b0Zix5
HzsKlKm43YTkjKWFO7CIiJTZDOMX5LveiTSkgLzFOcaSaleiAitFFjCBPWkCEQ8AKlf3GFloXYw5
jkdGDfb64LRx6zHIYnE1oP5hXLOC/qp+U2n4RyboLdtfG/L+9ra239bRUlAmpwr852x3N7E/TTtl
gew5YONSl8373yjNIDpwHNqyV9E45oXKc6eCOAj49mSOGJ63iUMEr4PA/hZBBCxLgX37Qb5OfW1S
c82Z05niSJl9f/WAaP81p3/k1c3Gbw/RrJp7/orOX5fgkTKJOIavIW6aod8bMRW0uKToqS/w4pVI
1AsoeIVQGS9j3YPQFgf4/gTn0T9XJ5STFS7bLUG1YPypn2wA4MqbGFWIHRLDzGc3xEkmMlrgkUgT
GAuunGbXkJrjXc/3cWQGlKkUBn+StUmXrTZXziWJcYRoan70VXpmd2+cs/eB3uHDNC+C56AtpAUx
T4rgOMChU2eFn8NTAb8wNr0b3BrZ8yUYzwMdPufd90YHP2dvaVdY0sDeg6r8FBsSBjIDGWGY8Y1k
Vwq47WNmoKu/utUCSdWbr5Z6Kpmm20SzOjUNpZr1QPQndZF7wzdrjfB04/0icbiBff1yGry0oBSr
H5aaHQy9p4SUjSC671yZYKYv4e/JpKthRtOHElUkYWhhNKxUmD2VWhpWcuMgXaacpvodtn+SX4Wg
1ztILJlK0Y4MQh6npuS8sEnJaG4NNx+fHo+e+lKycFbcs4kRec6cOizgsjhdO3GTK0jVDW+JQ2L0
/+n3GzEoUONsfOHeGNWyWNHTjvkeHyKU13eU7xpyTPXp2QwfVW93yMolce5zuuqbYewMATuMRIwN
VKvIadiV3ZdwePP7qlAIGBluned8GahdBTsISRcSkhON+vCUkMiGqNJl8sAYdSgcvXAsJsTizfpo
CBXxxRoy8B+O0UvhHvVuKeAkXQHLAHK8I6WT7DKpgw4i+upPSqJ0MBWj368Zkx4oYzGJOxzUCFwR
x7H5Sr1P/T5ifDT5tsAGPq2SkdqnPYdGImX1IzO3+2caaeYEFJy1SWljvTspxQE04ai5OMCH54pr
kcIlk9ClULogED1uP31JUEx+VUsBFW/hx9WZE9fG94s2I1hn6aVXEKOwoTpEaLcxKxDkidpSD5YR
M2HRRsVD1ZTzGPxSVg1JSXMsTmEQ88NzhicfEjzMh1G7FsxZHI3vpU2CwGLWqZIPbKEyyaByqxKa
3iSm5BQlA5Ez7WQ4KWnh2tA4hFC7uBNecmROtSt0zgXlJX2uDXWluPgRNd+tV8gnp+Hv6Ua4S9sU
9YGGNoPb0YNvN4/S88L9XTJYeGOGjNrC+lFhuWNzo9eNOKe6LHMMAk+jL/1LU94QrWHisQv/qrSK
EYvj0XdsnYqVrOoe+IX9y03shDGkitpt1HkBeBki1Mp53x2VlxLmlMe6GQMu4KSKdSQ0CHLD9UZi
tdzNH/2UOUBVzfPy3GeIWqsoiqaJh5HgHTIv55DvaatrfUya5uxtSeUBN1J+uiIuMGGOiS/nKgk9
v2jlPVgxzc6vJizjol6NsA+23Ys/kLnGhOKzBVRHmol4MjTbndeYk2GP+0JpOG8vvpPBXubY/3yW
z40QFXXB5hhgKRSsD3PJZ36ggEqOCWPpdrc7MOqzoSSq2IkwRrfTLTOoK5YqbT5pD1dALLKJZzvd
Y7JhnGRG7JCQ3KcWA/TTC/Us+g+Nw05w6BiQ+FEor2r4Gdtdl6Q5UcK9XRnaZgHLcF0LUG2ISU9D
yhHBkzzprvh8nUOd8BlN9HGSWMpyoKtKlMShB9U2gASdRKDa7IraWhHYd9lDshttAxG2UMMD83Lt
ZSQZcewQz6xcsCCSfUmKAA9YkBieVWe43IIKHDepU6Qkx6C0tzO6BD/JuQR8CTSYG+kzD3GRmUle
Vk4dCKMK2o9t5c5aNOl58xSQ3iXDkboBfcdfIBUmEnAax6lcOpjUvoDcQJU4/byHzsNrPHMkCiCk
ydv3NlSZeFV3mBK30kr9a4COFc2827OVz9cKcmfj+BREM+icwMnADYlJEUVU7lExGu2gGc2vXT0O
TvVz3eSjtRg/rRNR7ILhyy7N3jWGtGuPG1QNKNin+/y0OVv3rf6mvTyvxyVVgjH3B96lMidaM3b5
PS2B+jaSyRZbbUNhO/9gAWey0ODZy8CbWN4BNl7GfOdsMueS/o71jvQrIsBH4j/KkBo80dVxrtXz
gPvxxZVQxAuvv56Y8cSFfN6HzWZGyfVZ0PydklFoYpWpJkzbF82wRya3N6aY4tXAZkhaA39LW7PB
0AJPBJ+MGmI1sewhUkJ2vtHI1v52s5feTQf/zPg+KsyFSYv0b/wdwEuXbf/hP535qfWZNOgEAEQU
Dt2tdNRlL5TsVi40DPfBJgLVwRfl9cp4WPt/xLfSY/B1Qx/qeeMPbtvW5bue3FjlVUjeBi61/Ew0
+ml9pJsqryTRM3CbVWRH4JKpzN2b9Z1Mjpmb9Ok9N2qVMZi+WHXSnofYtLiCDPbZ4GhP6UC0gd8D
+NWDxvSn68YWt1TyiYkPOjoRZipY/ZVvF6T6KT5WX3uJErbth2v74S5Mecg1nuC3521dobO08iF2
BDgX7QXrPMIfVUcC0ImDwbQQ1sKpj0lOQO7x59jlnrRMzB5t5cCkPtOZDfRl3W9EEF60WIycUNcA
SJme0hmteUFiLZwd8Hk5KakuVBD/1sbZmbDB7aqpKXDia9sATynevqYOX75dZCe7EhLteK8n2cqW
rpe4Olx11ooGhhLO7Ve/SbuMQk6vqbwfgVgSEhkiU2Y4yvA/E9jBK6AH911M1QnnpdIQYkIjTwwV
Zz6z1cVuhmMoYYGHd4G/dqiOOBkH6nLY8y2kONqmgpmJC2+4SkGU4SLe4smdrkuew7HbAM8n804/
HUdSZORqfahiQXpn+8EeBcZHGuLTvUVdeJT7pw4ZQScEOS8VqZxPQ/3amhgIuYvRodUrYYKumxX7
OCp2Y4iIQvD/ZBGe7CoTKx2BlmJikuPikXt9TBrS15vSnj+9Rz1ESWE17dp4WrLKnmy5ywjhCH7l
Zsaic8g4v6YwFYXzQJy7QlPHSEqnbXyoKpXNsRi5t8fvrBOG1ZKyl/M6cc9V60KnElcdtKREv1bH
o54zOnEdnvcOkDjHDB8q+oB08crsyGdZOYOjwcZkpINLdwzgEg/IW37Un9fe9TpYV0VULIYYFWHm
16hgOWVpXXvfijU58tEo+YXcZ6OxkxLxJed6vdptm3yreBx2Avxi94iv5Be8QJh6KpDz0lVeftWK
TxJFv+DLkWT+Mn8ZKWQ6Wo7xeoG9yK06YthmKgO2p9zpkNBUyYi8sUvX05P4uduqkGM81DNP1Ag2
Eob2TueTDaf4lrrLMMRSNZ/jtr/MOYfFiG5DZfVKtRfYxmAtvJioUUFqtYHPQm1yWwDsNgjOWPNx
SP5qL/BkNO2HSQKOW1cLezM4sfqXXIrCw7at9gHnJawzmZjcNl/LuGCbBV3AtmkI3EVIOnR/jeu7
AP3Ezs1117LiqIS9i4R2sEacpzRZdaUB+jAmZPCf3CVaAetHvUnyim820SEPtwnaR6UNTyHglJjt
mFD6c2GP520AciTABmAG4UOj5g7fRqu/dRraEKD8TGasbnJ0Rm07dHwNLbC8L/ptVIY/uE0ExaAc
M9Lg8ZjTA7wEB6vYOBFehVG+G3QZK+W6uc1Lf2UxBze1DTmALpPZnM0QjOrQW9br80mTyws1XGmr
ZSXZXU1KLYupt5jYkHkYd078rGzLaBzkRkKryLQVPm/LKVJLepmTjADuU8J1IcBKJ6Rzol1hpryx
euqsChQegmetDgTvfvZd3J+dwHVEzN34Nig3FyYRCnuu0kjhhmqtzHHzJDss9yl5Rd/Fv7HKG0Ne
37ObgFSEKyQNShu0HNCLDsSpWlvWr8f5V89h9fJrVQgTs6bAndS9KQl65I1JPiSkGRJAozaSp/MV
0kBIkKlWKnbt37oSbnuOf2uZ5ZWBg76Uv8ZaS9o0oNv1kZHkezWr9IbYEx+GgqX7tLVHQl5K9SC4
gV1p8meE7YqxOf4K7MqfXLEYDXLLLDqtQhTi/MQIgL8ySpZpjUdzFLJfljybQptE6pkSsCH8vsoD
OtFSsLQ8jZ0sMMDQDqlsHnv78LLPG9D2bPkfnZXXrOeJp3T4JEgvph7iorj51S1Yuj4Fn99xLzJH
6AXwbQIAUzxjVLenU+WmOjVYEbhLpM2+tGG3t+oyPEoeax/V3dyHlG3DHFOOaNu/k+2948AoVsqv
DsVhcEBJL3WeDx+GcuZ4P/zLFft+wljB3tcdeyJTNdwjIHTO4KncRbXKVNAQU8wyPQzmzslfPwqC
CdITcv4HWByb7xyFLbEVtkoLK1ZtDRMtEwNAYpQJJW+MP73yQ3LiCWbh1X+oqgNkMguQqsM5TAuF
3DeWnbaGy9bjGyc4eax9YMPVCCSZuzUVCQJhcBa5HCXfGdXmv/9BzDuVAo262/Q5Lh93ty+8gvzW
w6vemw3Us+sm3Gqo0p6Qig2w/3dDZoZMip725aUiB8/Yef75tJiBYSJoYLLCMnAIRiP2RoD9aDuR
mxgzAHSeLyLh8NT7D00GhBbxYdDfd3Bnl9NXS1ZMKihXcy3D/Qu7TRk86adHhMzcl7RaCTFx/4OD
PcwvCOWcds5ZX4VNVxM65xeKQCgO9vlsNUyRGF6tLW5Kzir5nucIUemvqXwoyZtZApCQ5VHbcW3e
v9tDyqGz0CsCm7Ap/fujvvvO0NOcyvbn8Tj1+RCv1ySueNCt+1oqyPPPvPeIzx5FqGTgcZCX30aD
3bdUoX7IoUh8SGLp7Z8/fld8JHjgnFvrckLXX/sqxw5wGHB9IsYVIxs9FOgZlOPEn7ka4FmUaJpy
5Akx6Iivi1Dt0q0LBHdZl9rXPTic7A/jAeSX05CW0BByePxyDLgAcztfKQMX4DOkQO9uPD9mfQml
AN69EIgQzrHdaJIv6j7s/CSn4Q6A+R9FHgoQmRLouoz8yXN5ElXklJcEkbX+ezBQRghW8w5XGA+L
zhONlQZ01efdxjuLsS7I8CJaAUgiaW4KyWTXZY8HkxMvPISRE1oa+W6CjJtX3BBoCadBIAGYyZrG
Q30c5XakpheUx2ySt5WOqALXr4XoxooAmhWNQ9tmt4PlKtnc+5p9H4jwJpGA8k5nkpQh2Ymp7Xj/
uepQivWQcZIO+nXb04h5ZvXiImVpGvrqvI8oRhmlLnuOxgY/zeoKqefcgwVRXiD6Fe9rt3PeDMIM
a2KhZ0JRecl7PKuRkavwtbHjlUhS2TeVZtaIOJS+fRI7s37of9D/RaV5e2sejsyNDfAoU6AZytYB
hw5/OA15g063cCtYzUQOv4/3nEUEj5XvcfnThBFrhEk05mh/2qQiEjkKJb9h3s23DzBp2Py9uRRQ
lXnkhIcrt0Ysg1kG9joKEd5xreXIGpfGVDM618jLjoATZz4ymnIqFXyK1FLF1xfYSzmuwflhnVsS
eP7ucMVorLcnPwiHH0dEpBWsX5XlQL6jQiz0nndYiUFjgC/4wbrqiR8CCzjRoNi+YcBfBx8QcZTJ
hoLm68g4A0aWApvjknLozzFrNIm7vngO3/1wEg1nk1w2zwP84zIHWQ5XL8uVvig2nmC52QKQwD3m
tCDdpVZLGlk+bFvY791HOYYyInWbwo4vZcG9dyRayS62M3m5iGEzZTaxfcHzPw+EOm3aDh9/6GbF
2VgV4LNYTVdLjYOaTxu6v4j6c3G99SBICjDDxJ+7cI333AFQKuWrAgqlh0qbY94Ofex+xSgTwOXj
J1g+56xBTJ8n0am+G2ZzgizGkcUUT5eF19Vgsl+3dKsWUOyF4Cs9chvnVe59VYhgxk1UmjGIYO3c
RLPXDgMP9YKtXmtDOyBIsKaPpxLdcAaApb+E2Ow7OKRSwb04tNjz259C2WfKMfpnAac9EcUbeWtw
kHgf4Egd+F9V5/CvNX6C3uEztVG8gW3rAjWykzbjMM7CmlO9QmGYG3V0fG4N/15YQMfdJwBnF8sp
qT3jX3vSdAahND4qlieubNREiD8w+phwgaSkw2/vNgvNkFA0lzezNlZreelyz6PUNbIeKdsseodz
vnOVfBV/P/gVd0qBhTAlmXI8uLhYBWxBjrg0GeqANTMxNqaY8ZU5z12AwyU1ZzDKvsGCajGgQLNx
VtZvrraqyw6k9DnH2s2kVN70uwle6K/nK+vZZcV1VpaC3EfUb/Suv4ynLdOyEbU+4EzvtuNjQBDD
jtQ9xvtXGDTgviT5RQMz2oaNhi8XspR5oUVtLgIFwxuaIF1d3Csn3vnkCLBwLSF/LXyPFE1FPrS3
HXb+uxj62zgQcGX9xPjUFTyHBAVIeW2U7meXwM9CS2G6vylTV5qGJUa1dxZ4JrLlNDi0dDrtxUlI
TL0vJozZKagq8UfXjOV+TliKWnCLY2rlBnzbm7w2kxdQkPBEkfIhpffuNt1iJb9sHNl8toaWouvI
vWJ1ke3mrK3+gpFZCfnHaJ80wgtZADzxxmp6fvTCZvISnKlK9+P6DIp5SHcGy41QTVrVULxEBdL1
11g/FDksDkbiCloy+mxnb2B7xJauki+N7d62/2WHKAjOpNxpqhvUT1qpziKsdcX7Ej2jHorxMDh+
xot/CmZgLb2jtFUvc/XTGaqxBHuCplAg1+WO8paGVOTIlaKbFRBRjBVXyWpTKc7Lt3tdv0PNl9qm
trVq5zzOu2f7zjg4BViHqG6Q5vbqB2miu2UZWCM2UFzIMXbmgO2oIMskfRDck+k1K4iNS0Q3R1+Q
awH9F2lpB0bAILvmhmtmVWaLNnhb2unTigxu9myO8K6QcD94ksEMgzE73aP0DJhgZKGw+b5X4Nqp
jJDAce9eL09HxttqDpAccAPPRo6Cd/t4u3X8MLYS9J50tlc9W2Owthx30s/WA4kj/Lg+OliUdavo
stzAfkNScOG6pBDNI+ZJzhalJFZQV6WZ8BueWK3nUwU8X0PwQa7fmCPpFyoS6jxe4uZGffZ+dO7j
6OCQiI41JytOyITsOKfNlKZ8q49koHqO4kgnkHD/Fmf7faaq6FiQ9MKz4midDjAo6DNGpdj8P59q
/98pH/t/jSN5aLoP3t/r1DDSbPgetki7BUvTF+YIS3cPIyX19eyjpF5+Ffkdq9NIzo56zfWFP/GI
EDzhpzwA+MUYY/Jdv20Wv+s/B0xZyRdKin5xoA7SRZ3mextHN/PylTjaChiGx8zXIDFh4JFpb3sk
ntXkq8Hi6lJJX4aV5QSSPgW1OrBdV8NFvLMVJFFDoq+E8mCdmxSvpme89GGi1q/QKiI0i1mv+M5Z
lz2UVjo/RxoAyvvoG+7+IZwEoAq4ijN3kF3smNOfcWcsMP5VfZsUMRYLXsJWDx9xPtNDCHBpyM+1
QfS8OJpCnWk1vIFGl6MA5mCDifXZB0OJBAgD2MNnNZsB1slCtsXWVLm1/RpGUUdhWZyJmLT9QFKo
qETZARGq5k+lnUVaKJPfz7ILhn+JW+jgPtyG55QG/k21tKRLxW5OQIQEqFFPw0iaIXqE097NRJoH
9q+pbUKmHmSH3fWkv412k8bjtHaxyYERzISh05DUmxk238j8yEqfanemTt4Ld4K+Yz5WBd7aqv23
Y5fRt80ib2zjpt6y9bkjRvfMuKCLGH7rE2888moe3ksTKzMDCEmZqUxUgXVEkSeSuPMQOoxq9VTX
z5EN20sGBBLfF/iEax4FM/Qrs2ayeoDxb3qSNLG6SLUl+RsemVnhikg/4yynJGfKvCLlVVJPt1vB
cVJc7oTPtzHDoH5OIlZGfxUVrFhpq+378JCylYHaxCBG6DXSFFqtsp/4CTQNPRVOo8/h2j9Be2BM
HoA579Frrn7hnwUuCJT1ofEmdsV1u+kETGtGZILJj5nDh4tnbykk/7moVBDF0ZCqhLgXim6korrZ
rTIadLbbP1nECEqB+hlgKNAZDlUK9XatT9pJHRlnfujcrOCbAXHEtVKpzOf31YOQcQw8wiGtsg+l
NYOiIe3yzyzCRwNRtO9QlE4rZXK+y/FQQD4YFnKZc8Nz0ff1y+v3uG9RX1LOdDLc2hGajrInwucO
s+zKdGWEY6RH1gniSUmMHHQV84+tnmvGlMkko4tWK/6azKx/8XDITxUaBDDu0W2XysHC/eG2cTvy
rLGGN4DOjhPfoZXG8J2HWjt/RqOm/FW5OXP5NsEwMCvBDiNdbdCf7BvSjARzG/x0V2wdGHXEjbQY
4B/nKhhfqMv6XYAattFVniNTnhm42M7RrcWsSfwcg/X5c8u4zYiT5UXt1AiCIVJgpHs+gFWVpkTn
f+aE9S4NFuzcmqSIoUDN7uILR1u2P/V5leBArcu5m8FnYColTOu6D47Y9h6XfG5wxLrVzPpFGsX+
hitpoQDBt71GjpdbhWkiAa0AAR6L3a2lzkgdEUXa6nsFX2s0PcwHrVZlu07gIEU8yUAOOF9PgzVT
qAJxyH3bgaq8P1/LFLadqyxKRmGYT9jPqw0nY1ZgFmh9VSnaqUaeQRyVwMdqJjXMAiyHf+SIpx6U
Ph3QoF5kdKizD40QQfEs56psAAJOW9IxakOO/wenRHVJ5aMMvO/smtYtFWdd6jQLknoyKeK9S4rB
UOT8HIOUFSLCVYwaNLWvs/RfHxvZtzKNca1LfvaMrjZGValDLAZwQVYF5fVYkvlYVkOQAuUzer+m
xG1JDJkLUR7zdE44p5AiSNu/SWviP5EmLyOXIrH0JD5M1LTUd07uQLFA55DzX8j//ORjJT0nK5yM
6VCk18GwHr2XaGdVkMufMjBWsdTIx/NragyxYgvWjSpNK3P9/HnBn9BI7/181cjvtW0CFwCPbAyZ
LkI3wMUTl+mKLwR65I6kV786aJdotnP0FzsInkbaEbCKcpRqGGjZEB8j1ajlUh9dUMMvSEvvc1n/
sLuWQC65X4j/nqPrp4MZE6YeHlNy202a6d3w7LIYS1fHE/2zt1tI5VysaDypwdYK4Xg6f3jB29O1
WgyM85pgeAzJFNL6rZ8llNtJIYTwlTEHF0/DnpvT78ShhTGz2shs6mz8aFkdUnQc2PhHdpUgflIz
CQfGtg6jKQ6Sp5oMy+yPgtpEYGvk2bKWHwuJaTtFtvMmU/oPM/srqWBQxLMiU+soqoRVY5hBsYbo
Yk8hu4Al20wdv7VZnDpdA2s0CeLHNJm5mIX/+SWSqOZ+GfPCJhhJeUtcu8WK46tn4LdlVemuZPt0
cbA6QKK0O97qDLmAfDyGrLmp3eNXhGT8tgmX6WH+pvh/L2LaLGdjcCJSt9fL4JmhmQUQnFeVrVG9
oriNJjSQfUa4n5oXyyl2LhUHCgGYz/0jzV5V5Djc0M0pyb1ZD2ufivWgaudgn2glY53VlkSwjdGL
nTWPL85HSm0Jyjm6nIounj7+tmR+BwqU22acvl0MXVG0W8i1bXdQMLLrZt8N+LgFlgjSLrvtvjk4
flbtMuuvQWQHvgCmQRicCNY8WHmrameDW25/dqoD2lYXZIwPWVm08B/8U/IaskM9ANAA9HQUo+JX
lY3m/u0+Wztu0evJS6wfMUPSBc9oe8aaUbXkha/Xrzb5Ikb62u3MW7CfwbilgJZDvfJUfVAbXoLJ
7i8bS7+8yAAQK54E5JGL/mnbPFXgwf1ne7THMZ8OaQdBGgsSRYexeU1I/dwbiVl8x8DytwMwr/wn
v2OjSyrji3sLjsb3T2cwFwd858E8Bty84fCYgDLTvHRxqy/mB8XSiAA/Cm4HMf5+gY+dZDn3Bw9n
NSrvtgZfNYP6yYYmuVd6a5A4AkyMslvpmIxa5gWiZi1R6dXbH9qFa7qpyRZB0JfAn5W2zhqWvOFe
93nR8+PbxUURGbk0005ytbmC5uesc8+5PDH/8arqOFUivALIfwoCnET2zZ5463doF9ImMTLbcPxD
T7ROJyRBFtFOhy39F0jQ5+3+VwD7eAlMHAmsHToN5uUrikUbOlQYVlyRlKQVrqHst1PNdgsnp2R+
UC0J8zDBt/2PVobewV7uRpyKUjHBEs9Gt/hW75w9JQ9/pAAYu+nvkvbn8UXnPr26h1kwTn7KdNgq
JJ7j1uQS5mENBvFUMOHGKAqzYtalbq8Ra064LGHUYUvCy0dSJgJgGQ5Ie9lpslXRNAtzFClUEP0o
Gf/3qlrDmpwP/7paJ5tL08/2ozpqYQ/fgNnp8p+4W00BaOus4rhkVMzOEhZDYOLeQy5eyOwm0Sa+
v6Sl/Ldv1sBTyCd3W+kqNIFBq7ypuYfGhu3OiNn8qlqhBNpKHoWWsw3sh2/ycVs55IqT3JEZ1sYJ
n8630SI0KSomAv5ASWE+j7/1U9XyWZWXCNhFbALxnu0Js//AN1AXmrvTPjYrYXAMZu2v/3SFt3FN
b/eXLI1ox2ube5ES3ZQyAxSZ0JbmWh9ISRRp1dYNOx3P3w/SBFG9wQTlI4w4vbpcKuKRxZ87aGRU
mjNv0sYQnf3t85kdrePWdzGTEy7MZcWLWxbnUGwf1hqVABO2onvdapgKvsa4EvFX52kObT1PgJPG
xMxBhDAANQq2hHvoFXTN9SJuV3snrRVvu3GNZQ271ez6soXw4J00IX6jjVF3Vh55Fz8Sopt5ewnN
90hoV0PyatEDlrXZZO4b+xhK903ZgKXYBHPITuwq+V2hBjYvegkMoKN5SIGAc5dVyJg8N30NBeKp
F0OoGXkgKdGEZRGNH1xp4ZQJspvVsTpaLBbfJUabDqEanyU8w7uMJFs83VydaEzcPMKff1ME50aV
PUJYoDBpmmLIHD5SvTM4//v9+Vr8oWitiEfYrrX90hCkIWvTLnMMvq9ump0QBG4gsyfxXSToOT6i
jUMLxKPcoD177+nvYfgXNVI9sBHIrdr6+AbOpFkR/civrtyY04X8PlN8ZfCm84bSbAvLVUQICm2A
BrHdUuSddM0k/BdhI+6C/ksSSfrkwamYKWFqRNMdtyaV1Zl/MqLuMpUekPAuHPQ6oA5xrxtTrsWy
CIoN+NzTn8UM6hGXaWzhP8leKgoL6bsms9oYVG9vNCpzpDbFv2oMftaXLVNjGM1v3W3K1dcwXtyt
O/A8gwij9Nnlj1i7VYmIzebQ60Cf8zZt9Y1+q44I2I7OgUCWriPExmbm46ONl4BbMjfZyol1ECZO
KBRa2hvX3OpZDkvfoNE+pSnzyTzCeMGHkx5M9u9ELe1nJPAn4rgFT74cSxxHo/8F3GjA6yxpK3C3
fvu5XCACP5EPy9ieWkIzMVwUei3Qsf46pJO0TfJyOHY1aqWOSFkRhiFvsitPl+Fl+58Dnsz0Dy2f
fVLDZpiUuqovbtTpUQ+sHJb9nH9Qaypa79+WOCP/VtLH1V+BMel/5wkrEN8fyHEW8X9Mkd9EMFXa
ygRHDJJtp6w5jx2v48fTy8xLkCHL1E+5zTALOlHiNoA7VtZ6IyIA7d+4Hi2e+W13Hm2zp59zmk5a
DUAN/Jvm9cQnsrjdWyUYOhLuin9/TCnLCBjL2xEFC5ELE1mT4HIyerueGr6vgqYu3esIqMte2oMu
CbzIEk4bJ+27pS5Yz6JEGTEGXi1HBD76yAJ27hXFG5D6hqLvciq7EQ671UColCvbPItVNsUVf/R7
WmXitxnWpiVEpvmJ8kj/00UqAuOPSt8qD9DNT3k5JSbWXgDnC2FCjxwQSIVvg4vdVU+9FxXs7dku
dJzKotzaOZ5GSib11VQF0IIz02cXAZkcNqvkGMuUFVeIYZXNMhmz56XGAlbirqOlVRIdvi6pZS2e
09ZY2BIc53HXsl2cCc5FaEft0w3lJDoqr17xQqxETz3SoPnREBJEnFrIsNIcg41URlcWpblqwO82
ETXveGqENwO7gF4+KeJNV/UeJTyOtbuuQXBHqO+munCTM2dAeSK7EqTb+B+/1d9W0Dv8bFWB4WBC
XkcOXPlmMTIaby2nsUlQ53QMMAkhutQUHr1NETVai1wqyPKodge8ivKLERgV/Hcnh5cdVOl2WYvZ
h8/IVLgVDwYlupgaylk3mpVRNrivhdniamJWsI3DRqQa+n9fX/pOfGGkgznFO97Z2sh6Xs/Ox+Dy
XT6ZLqSqJ14RXFonxVpTjHsa0Eibe/igwurC60k/amiiyTIFZypO+IMTcp4H9YopZ8sGG7DYa8bp
JXB8x0FKXohSn13tzwn+Naa25dEnLaYFhlCgmeHvTPZ7ngFqMI6qbPAVhoIcmp4VAdTglo00HSjv
Rs87b4lrzcDEacAeprE6a8koEkSPWYzG9DVKSCvRINZ9RT18VrRz8KYfhqoiRdNypViB//haZ174
Kbcuz69IsBwSb1vzXFTvwXIwZqxMtber4BKhilYyCadDSBM8p2X3/Cv5c06l5FhywMrsC1l+eFH7
QlQGtQhUwOrsZgDNT05mQ9V57kSm+RLn2w/z67T9oTiHpBKVxz7pZy2nok2kLeUKT9ICepZIhl8n
MJZrfBDdzc/NfYGUu0HLGdCB7jbTiAC5MrKg2Q/IkPcIUJj0/a2/YlNl9O/BoTzPhlegifllwKPK
oyCYyI45XHCVFmL85hRWJtFZfz8WtQAVEtiTkxARe1RdSGIdUCqbkH+boZNbs/lHoiBmApLbCQV/
Yumhzsv2UZgbe2606qgrD7Q/Em8k+U2DMisfNdk3nFiA6NhQMMrwAEJf2u+Kd1Y5HZbfTEkvhK0O
DbQ2n65MmZSlMuFTgjuKTEkoru7ZD2ohgNOzUbjU10XJ4pabzFQSxi5EqcLU9NIjzHAvRc1364s5
mXpoJjBfRhafh7EnoLJpW5ptEORdnjxGvZRsozx3/74tR6xJewP2wEAqnEnlpYcSgGFBG+G1rYMg
uoSAACpwG3f/7ts6diNvlatsAfqIAFXKr/3eMfp0R1sSzFBRRDaE6syeL6dr2rNW1oV1vcaxl3o7
hrTowUD1Rt+U6Kfohu9mvEGMSaxfjcKdHPMLyRX7Lj9IPP7ssIjxo+m9KBAHtiybJL9tQbaW2+Mu
lVc/f6dZ6BuCUrNEMSd39id8cP368f0VVzjn0yXVHqFLWuvvMLM/Yk+F9OsEjYY3wKyvSnNbGqda
TUJ8RuzG+pnYNavCvy55TyAui7jLjxeC7WI2jGAIBhshn67SOP6h0elHiEXM1raWWqSTdRp9JSWn
nRP5fk9RUK3JNLw/uSSMIuLEABLySFuqe64IMGz93i7DJMK6E2NKeGBWEpsnrnDFIYbN+3mh1Kh5
IkYrpYXxRBDKf0F3KNMZ3qBbyRsJl6twk5ax6lc4iZfO1z86g0wL/7qeblktxn4cdkGgEE73DTu7
zT4tTSyLpInr5SSZBp9BaRX47DeH2kJxqBdNb4vcrFhlTpbc9iLfv+69cB2tYJNvJodEDRZt0VF1
pHr4eLeTclYLKHJoWGZdKFgsfzwcM+AbHNl1aAOUlCur5NjktyYqAAEfVtaRWu+X6o+zHH48t7ue
cTNUDijsb6dwoH8YjS2UbpK2QIg8/ND1L3lH7oMxwtPxbeNxdxv9vOgXguhBDVq8cjNWxF/tqxoq
/oyiswll8Psgvf9wznTxxyO9LBpL7xQQ4FuWezRRS87gRwapKZZ1+gRiNeNa2/EPXG5DXsLVe01i
tulbBkLZpwgmoFKEJ6RpFu+Gxe8NeAzN4nmuIuABbP4kDfAfsQDc
`protect end_protected

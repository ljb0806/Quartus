��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y5���g�v�:�[M���y�?PD�C�c�4�c�������nPH ���3>�M�����E���H��zh��FX�I�:>[¼��c�C�.�lv�" c4m�\S��!j��6)��u�T���$<L262b�k�h<��p����w�Vq�����Qu@f�֟���f#ϰ�rT_����'�Q`R*�����^�1�ա���)�S�|uz�����@*[!�&����*�����M2HE[���nC��Fg���ݼ��c��u���	���X=���w�r���k�^{�w�;eD�n�-H�e�Q;@�nħ�c4�8L��#�����K��@�y��i_ȋ�Ie��������d�9Kl�gI��0|EI��}��G��"[E �ߌ{a�n�a�����
���b����T~�k�5�F�j�X�HX*��v6��̡�'��Z�-$�*g��x�ɷm�ö.�k����{σ�/�T�lԳ$�'9.osu?J��B��=�6��?��Ǟ#'U.
aɚ�^^�-n���~A�
��'��A�UJ�s#�H]��f�)��l0t���2� ~���������|T/Lw�`R���� ܟ�+4"'2
&{q�*��B	P����Ԉ��Ge���K���R����~�8�P���"*�D�K#v�FM�����-f�uF'�Y12�-xi]���m��Z_o�T�ĺ�l��(�q#�C���x
?��A��C��	�^�78������J��'
Oѭn�% �99|�g�kH
�w&����w�L�t��@���u���޸ȅ��lP>@��Q,�۰��7r�~&M�\#IC>�{�~�|9,<i<pѥ��	 ��"�_�i|'@��l�5��5z� �k�ÃL&8Wk,p�8�3��P����!W�����/p��^n���^�9�����n��׵�Ϸ��M⾢���p$cԃ$��87�n�al��pK���jɃ��Ai!]5��a��z<���of��P g"��@�=u��
��#3��w3D��Ę8HrFp��9���"��q��`�_(�d��ND������'qe��O�9@���)f@��� �zxHE�o�+v�X+��u�Iq���3���ͥ�`�a��|mi�3#�?�2��p�pv%bk��j%e���jn��l^��JR�s�[*��T������N?��)��eM]��,��w�z�5q��ןm������}i�P��4�#�P�+Մ�6]&��2Φ�z��I?�z�2(��z��kD�?oT��҆�#����<���a��im�÷]���Ɩ�Í��X��&4a3�ima��E���łFX��u�L	DL�Y���\����B$����O����H��ѫ�-��-(��e!���%�!%�����%�8M�`��U�r����MD3�Sz�}��g�Y�M���0 D��XV�Ê�_��g&�>l7� M���~�*��#-���K4������,lPŔq��V�zES���ۃgfŵ�; 2� wjk8�dP�3�}�ң}�x�!&{a���:VB�IIy�s�б*.T�v������⿪�9-:���]Z��T�>�Ƌi�4:,���.�{��O�{�L�L�Z �����YFZ��&C��j�wsb��Q�aR'X~�0z�M&��|�p0ϣEa���z&�����#|@��CR�7�" $����.{J*S=1��: 1m�<���	Q4�'���"ڡ�o�F8���wI�Xv��`'n�L}<�\U�t�H�|�d�I��CzI��'g�q�/%��>�>(?��
����`�-�մ����T�1?����}����n����
�0 ��֠ٝ��������?KU������Z���@d�e6'u�&mw+:z�$�ʮ�tRS��"����H�,�we�YG������+_��b����b_[�z�p� WZ�_����cПB�8r�e���k�-6O����*YA���(�2=�C��v^o���'�?�,�j��M�USǬ-��'kh!<иB��2�
�YKu�|�}����F*tm'��� t�ӫ2�ЛH�n�WӜ�]-I6(vʟf�4�',S&;׀m��w�j�J�D�y1Pk��a*!�j�W��"��b�ID��� _�ͼ+kL��@x�PC#Y���|��ʠ瑥�(҃����-LZD�h�������ٵ��~�8tZT]Q�N���d�I{�UF*9㎬��3������<��ߗǩ5�j1;[��^H�;���>��^��e�U��]ˮwu	O:����%���������w���D����)V��.M�w��}Di�
��6ɂ�*�J��g���\Z��ӵ9�a}�ǿʒ�D�1!�h1飵u�$Q�2�g"����G����W�ݺ��qI^��p���<��Km-�#�r͟p��4lK.��KJ�}X�j�@3f�	��T�0�A�8)�輇��X��E�?��)Ԡ'�hK�e��Z��E�Vz�D���*0d�hP*¡
��F�Qٍ�*�BU�8�~��zǐ��ʨ�KR����g�Ƃn�A:�j�KF�i���Es�}0{��i��˿�uIQ2]�s�i�i�<��Mczd5�(V���I�X��\�+���d����O�ْJ��0y%M��%��0E�k���o"���؍e�Gӆ�����]Ƈ��r�#��V`��^+���,��8�FVx��cr�T�8���_Cњ�T%Y���Y�{��?�9Òv����X�c:���4	�W��AW��U����ʙ@��mL'H[g��0*��b��"��I�4�k>m�I.�G���(E���s�+;��պ��R=%��P.4��a�'9-o�`	�Z��o��������B��r2��N��4��+�d��r�̬w����Z���v�w?��|�'9|dh�V��K�r4��F$�n*+-�Ա��J�,���~L?����to����J��r��T�\!Ba^��Y[E���.iwٕ���J�0�V��S�O��Wz����a�q���}K��������N��	��4�0yO����q����#k�Ӻ�Qں��j�]Z}v�B�z�G'�}�Eg%��\߃2����+3�����0vW�W9�֣��W=Ri:�`�x�� S�eE�����qg�ׂ+��w?��c4r�F+"���y�-��d-�٢�h����*x�G�g�JCX]2N��ߔB��K�(>l݃'����5�u��'z���Ld-5Fi��#eX�<=k�݄		��0E&-n���&���b��菽։G%*��(qIu�(Yo�cS"}+M#��.�4�G<�"���s�u��x>��x&"�r�֑ k��@.�� ����,���(9O#B"1ߕ/���a���E��H�����H�ஃ�÷���%qO�<�
�=u�8#�CϺ3h�wlH�K�gNs܄T>� Gq������g�պ杋X���]}�l��:��7ƉM��h�|�GH�)%ĶH��=�p�����$
A���Uu�S��.��]�[r����� �5��(���v�`�L����.�U#���a���7��~���r��l?���NgIn�;S7R"z�	Ce��@Xs)��c�Ã�V��N-��3�E��J!�d�p&gM�l�a\���+Y�����Pbr�.��Ά�3�@�a�w�tn���=Z\�7����nM=ӣXȬ��V�z�#����3]�}5���[�q� ���q]<$�}`��;��^��1 ����{���঳�����Ċ���Tu�q3;9Ź�zJ��.�5Mu3W%͒�H�1�����IV�j���f��EP����E�Zh�����k���60&�<Nrܿ��A��
-3�ȿ+8��TK����Y�9K��\��bC/F�1Vi/"�I݆T����h�gXшhY�na���v�'�έ����d٭S2��!�I���	�xC����aL���*ߤ��żA4&�p2�GZC?IJ��C�N���N���PH�	�Fs�,'hٸ6���e���K�}�N�Od"u�SlE�����w�Mזb� A��x���+�2�[�C�]h
#����N��~������$!�&���JA"%�-bu�U�ml�^��}8�J�1z�̱����<qɿ�l��+鉊_QB$�\A���_�ŧg%�Rq�ok� U#��A1��0����n��Z]1�^��缼��)��i5�d�:h�p��ec���$�Y�L(�������YƄ:�T-��zk�9���M��=o���u-E�|�F�ҭ�d�:�M�ᷜЇ:�[�_�ǄE-a�z���^�m���!y�\y��ap=O�C�$�a�K���I�����Dr�����[�;�}��D�T�[/Qa��Úp?$�
�E��W��{��;�]�{��i/Ihz_Bmi0���lM�x=kLm?�P�pG��C�_/>�B4O�)Z"`i:�ᨶr��y�5��y ^�<��X�W�y*a�-�i���_�
QU��G�[��͛�� ;Fj�<6sT�Ȫ{#���2m�VZ���&m�0.U�i'�ф�^�J��k��8/��g_T]H�r/�<h�����I����\hTL�F&��g���˳�S�����Fs�G�qW�u񊀁ԕK"MٌZELpu9F����b�CZz��0��t)�B��'qJ�g��_x�ZҌ*���^�^��	���b���iF�^��Y�I��h�vG���d�
$բX�fc(Y�̩�|�#͛�08����kEKHw���Ѩ���iRXe"�kT�5T ���#��c6x�� |��Z ����2��II7��?�B6+=;��׆�dD�r z
G�c�V8DZ6*����@%;?P��,j%��H��_���RN�����.�7{;��Q3q�����)��Y`�_��n�qzI�Z���Ǣb�xWB�a�"	ݹeKb̚���qy�΢�~\��`�f�q���k/� ^Aw�?.����YPoTY�t2q�'�Vbސd�g|9.��ց)&�mG"�^<�T4���CD���${�[�ؗ~:Zv|��;*J��#�M��0�vX{A�j�r�CZ9�~%K�}Y���w�����f;x�I��V$vU��Kd�u�K��ƷE��V?7�>Lڸ���Ռ��	�$��^�ROx��o3�TLAS<�}����<���q��Z ܏%2!ذ�t�߮a�pa��_�wp>.E��b�ɸ#ೕ!c������p�3��tC������&�R��V��Oݚ�r��j�X�u_Ps�{D�J~!�b奎���!�i��tls!��v�l �8ix���9s���"�חP�?�P�-'�xɈp�Sm�it������橥��߰�S���c>&��YlF�ej���>�F��!A����y�/���J��Ȇ�̗�`8�>�R�K��P��yQ�{���ň0u����3v��	:2�PE��o��dHz�U�Ӄ!^?^`L�4�vztk�� ������o~�J|+�zG�N租�խo�U&&��>�s�g�7��=@�ځ�o3P���0
D��;QX����.a�d?]9���K4R�O�L�=e��� ����)��<��H���U��l�"�;Wp��d!K�f5a�B�gg8z�N���X�BF�=��9�*c�)ʊ
���h�%��ũ*�3EA�T�s�QEX?o�(�I�n�7��'�&!�d��X_j���g����4ޚD���HB��|Z�R��mWz�M�h_��AXoN��r���os��tq��`;���o�D>'vu`F�pVDC5�E��J���B��5��yH:�^��*�F�Ta�E�#���,{/O��m�X���Ng�>"��,�#z��'���=�K�q���$�
-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RBLJWtWJNCYlWmzyutCdNkGtOH/hcVqzy8hTFXdpbj91FIHKABTjBYiwCpa8P93mADZKrHERDweQ
HKNMqbbY7IYJI9EDuoWB/0cAgkTam4JxeG/jhf4+V4XuqdtFugRdRPAMlWT8MpDiK7azv2bw3u3X
5FA5FckmqLEV6vVYgoMXu4YQHXMcl2oNnR9FMLJptCmufAPASqV41pPXhpoSMz4Os0O48i/WivLe
grAA5kk01j3seurt4qJfShsuT5rjE2jMFy5i8LQccbHWVx55wo6Xx3w0IxhW0FJDycQfi5nnGBf5
OT8GFK5nuamUGqnewORISYtFUnRb2vMSWzEJZw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12400)
`protect data_block
toZLirAX+/QDOUgTOxggQ25Euf63VZYjNgh3YDO+F6PaluO7wgagvg4aDTPYz8v9LqKITsFhNYd/
BHfse69nUmZo98wzU/ulVwYFwLCXMESIiwJaq9nGeszquGxy/5iqw+enFjA5j9yT9/KybyEwBP/0
JQ0RO6Oc/rTyAoao/jLdtSGKaMaSGVisYXiiYwBeFDTa6LNcNwAziI4mmht4c8A8ipqXyjBP6jiv
eVAjwWnp9AfGwoejqZQ2yqCn+EBPusIhkpq65KEt7msp50wJsEWhdUOfSayP8RkwONhBaNKHJN5h
vZpqkFGWE1Cpi1NFgt/gAPAdcTt3DVIMqDETNvp/h02JvS5/SxwSHFEtPwk25NqdtFSQU7K2xVz7
kL6K96DOeWz41cq9bCUpdlCq6ZyiNYnZI24Co2q6nSi8wxCgrUdbTjSMYyyPqzun1svKnxZJ/Xga
xXHMM7BaG+EdyvuZwKS44VE1EAOec6AHrrD8YJIHf/sxtY1uVr8wHTxh6ERYHEfx4nG5RCUIgO9+
owmW/xBxUZwh02XMZAQIN8p7ke+2rPpnAPQYaveXTph9PG9lp+X+OsOAYFVsxfqSiyShJGvlA7rZ
K+DnyfL0b4oAfIz2xpzn8zYNyJyXA8gAjSZ1Mw2BDddqsgNgk+GoOeA4jF/bPCpIVWiKhMFfBdeL
/kqFemS1c+LESWwqRu+XW8GCdTNHiO7oNtOs5UwMXOUnGQJQdsAEANFqai+71pbdcTk5ienxqukt
F+HsvjYLFVLYWKFygnTFMVzkLrg86RzG5a6uAofJVqU2MJIdo/Yt97Hx6ix1/5xR7UswymWXUTds
w3GBDL4xiyzEnyiDCQgc+6hf7kYN3db1j9h5+8QglyTX4daka4P1m/1lFt5vKdVK05cXQ9Ft3jJW
vEyrA4q8Vmjmf6656UlrfioIAaMabxe25ZLIjaxZC00wCe7s/c7Yjvp0/jVMyoFdvLHEMrQpPGbN
DmWsCNzsAsgpqi6mlTOq30rKfUHLY2sUjm8I+bZm3+12Q1HHfHHMSzRzjVdoQzfKyiaa+iQSH+kN
n7ACvRHTR4Z4me3DZLA+LbKFoEioeLwRIoHAzjsY8uhAT0umfNd7p9Ks25PefNKbKhgpcwBYFMkS
AQrU8IurShpMtjI3R2Q/ILONbvv7k4qH/DvNr/G6x/MRXuwGpU87lT3mR+IV0+66dUpYZEHFdxo/
mEhfX00ToHt5fS/NelUwJ8/yDNI0/p98/Csrw/O/6CiUGbrp9+BzHLGRW4nxq8LGBGPshi6YHh2l
mZ5ck4vOqogC7y8ja8lWs0tbg1/QX7mbmEvhoFQ4a5b2Kx4/s/KpTKHwDZgtZ7clqQFniWBmg/xh
fHwZkXHCNWiTXi63bNtSnQ9vgChANLy4ip7Xk5uwQFqO/g0l0Xa0U7uBdZ9NRrDaL7fZFHTSQPSd
SglhIAL70yYb5HpK8UtNormByqBFobAaIITlbRdV7ek0gGKHBjPKSEVhCZqAANBunxAMXZ5bQTsw
xhGWo8AEWZHQZ0CVe3XJIx8fmdaSoz8h39wby2vmet/Wehp90GDKIz8/sbhYMU2a/P3ylQ15Gnpm
WyHRnRPOLMCWl3hl5Bve0DrfC5UnuI28fEtGlFZoXgbUo8g2OKoiqeOFzTMvy0j0kj4DhrV2apha
Y6LjrFr5fl8P/LusuOpsKGdUDcHSNc+vDTJedpgxjVvdtYkffRYSDfvFBM202B7VRWXHMmYNhm7O
c9Rtv9/bgZm+NwZaM3qdy266o9K/+NXvZFq1h/FGnfRNyUzmu+zgZrHM+5s7+VZ/P0zQTiOKcvIy
7TQ/45ImjMbjiLMxEeiw8WiWmArcDRnYkHgO/I9cOOEPnnKyd0llziYdMktjSfRLx0NhnegA0dON
uKHvxZxoSXUmndT7DTy/CbMcuoB2toCx83cuKOiCxyfi96keH6ax+GUwH/blIA3rRhX9RUcMagH6
YfbKtNIMYkbhyhpwR0zrW3f8hpJpYkxyk46sH6vb7uGgoA41RXG3Wi5fRXUjJfWN/GVn2Zn0Ga4W
qK1b8M1qvVdaYl33bg3DCHeU9CCTXDmgjtoURVPadMou2fEzTbIVYc139yG0W2XmSkpI3bUkOavp
60yjg2eg6aw5+YxVblFoXAMF04RIE5zhO4xOu3V47oeJdS+Oac5EgbrdA7QtgOKPRrQmANohBh0G
HF0+Y2g/GcaUdFgzKsjIHBHmKvNOs+qV8ZJcNkl7HIxKozq4HcsoeWIV7ZDYjRioXFsgn97Mh2kW
lLrjvB+c0No+TJYqKVcDrSnn1W6dx6LwweSTaTwTsOWOhPXy9AOcLHLyWo8i0SsgJT0E4JaBGLJx
r/hxigTY5nk/MHqf9O9oZ0BjVjD94P286dcbXjmBY5WWFg0lj8W5YwNEfUfIULaCzZnbluCDFmqL
x22A7mtaEIS3t5VX6w3JpFUSpw7joj6EdkdXfn0l/fBdIyf8y3jAczgc7Xb4BKwldfkA8wq86p7h
BWK0gETQMk4OaDEPJl5ecqZY5dSYvZUljFp9KZfNGf03uRTDuU3dkdw+5pyYlCyFHR5hfgtYTdDB
rkq/mmvHvDTrbQUyQGIqDHbae+PZLVyxUkVoSs8mSxLalO46bb/kbB89sO9+Jt9TspKX7VHsM4p0
l6TeaniEOtiFyxU64i3PaXmQ7uj2dAL74TN5DoY6+IKvcJZCaa9jL3LlvVbs9+ExP2vzY9TiQtZA
VevJxtdTyTyVCzNpPSdLl35+HiaKIYEqo2MgKcDgIT1dA5Z+19prc7vfljn1ePhJ/gGlzVzfS+Ow
wLr/IxT3Tc5rwIETpEq4/VJZgsRkE6xkB6xnDuzgUk+G2OqdB1+ovyeI3yBU/wnCev5IgpzSSERo
FGA4uHY9ZIW6xkLaMK8aC7RhYsNdiwXscExrGi3y7Nl+L7oh2LBJa5CYGt64mDeuAD6vpyM8OEQR
xB1lk1p2L6Od36VIC6J2lsvdCPaqBbkjgoW1ZHRedRd4cywldF7dP3HFcEfUooNitIc54kOeGir5
owDiW0kBh0oiDWvgZ8d8YZzuKYHpF5XGM0+D54LFWwznP8MBwUbbiu95mxosbKElmOSGFOdftkir
UOgJdKCtkpITIxG97o98ae+tpz9vwuonR9ZFNG6rkmCFg5Ahjr+7JO8LtIojYXzofA/sN9VOWf+p
QelfpFN3XlqcENXKab12TaNfoNlzmppmpatFyWrJ06dcQ/0TbIVyJ8lPum7/2JBkK9m5606MH996
xQdVqIeBRS5IMIIxMfUsrRGXNRTj+/KgO1lztAxL4xZkp1tXIlNMoY5EB8Xe/PUwjMsw+O8hnkyR
rXc3JS2LbUeTPcnL9x2ELvzEnZ5XkXtYg3liImqLG8Q6mbdfbBkEgj66TCkBBpKh6/CJRYKDV8Vt
1nv1ajMImb7zJCyLQn2IDkfq5tqhh7Cm11SnwgkqISfqlWYTqNEv4DVLODmcbqJ/pbdmwXcGkVLr
bKjL+oA9YnQ7HzWWSuAxUIuqEn2W542AalUTxYNSqtapHdo+u49vdbtkAm6Bmvvt+2NWNA0pehb9
4wevAHzWJoe1ULBHpP7d0Z95gxQBJCKQqX0P9yhig98uTRiVQRt4yhmnn4vLAM7lFLe6AwgpD28e
rmTON0JZWIP1JuuVn/eisqEzGgyXtIGKSGvualuvDR+G3w6L22dGc4+ljfoqY+LM1nUuL3VBGIOe
2EwnMEsTesA4nnNYixs6ctt33HEMGEb7JS/SmjWZbLhUnmPvv/eeYKWiBj9UzI+B5lxiV1wL2UG7
tRixuwm0x1ZMsN6UApI3UQu+GlE/SjAFhevkMTJ8meyYnKSRvaogOr1F3gVh2WOD1+FyHM6+Jcqi
oUKY+gfRMOnEvEhjmBpQviKO/0mwUi10GvT2/47u+YdXlABgXBpAFPeCOmImlKP2QxPvYKtHE/y+
qSp3lSnoxSVQrBmc+W/L0gCDl55mMuSGYEKr6EP3HbVaI27dgEIlhpbrIC/ljlTEIdxEKNPRpmX5
wnrqqBL8HPvhVupxFXHSeS5WROd50Pcf0tYWN4WCFRiakqsse47um385D+uLTWZVZ+Yhu5El+utu
pCLH2C56bg/gjdBIbuglcZhh6d/rXIOqy+xTQfa1tbzOajSjKZpretfR/6xZxwNUzfDzdluWXGTg
iyOXcbhuXbPLff2duX6OgS8bULqS3YvKqRHfBlgIdTdogjvyenIKVvtlM1mw9SdxI0BafbzSwFcL
IB5cFY6rfit1Fjg8X4iTsN6C+kF8YjiGCPhkNttKFI4MKQbaj6kP1oAqMToBl/ZKdwnqZ3W6cdnI
qvBYzMBv5tr0+VHn+59mMSokNW5GO9IXr1H12V4kzRlCFgfyrLyd6cn4nZNu7aIMifdM2h3G39Yh
3ZOAgScZdBbwPFEJAe6Bcu0SCdPnsWGCraBkySPK6Arp7h2TS/ymmG3Q005T5Z4mMIdT+6VUFV5h
fPMaH+H6F7Z9bGIXXhTfFrJDZ5JjiQ1CYEEclMTidNSlYm2gjQ2sJpLvQ/BQDk2oOJ4CX+bsfZw4
MsbbRJYsSXBoIH9p80yCEn6gEm5W6r77/6nJ3bi1RIXlT1LalsHqlYPKOqAMA3/H7S8AVf+wh6Zc
3aA3jZaG9WuSBXbQ8+YTSRlMIFV7gqyvb4RNesU6pLwjHaljXoTsBPCnIS4xWVABtjc5kqbVJe+8
SdPy/2f5vtod/xDfnKlGPvpzgZatzApmmRE86nxuF9DcqM9kLIJm4ECOTUEd2Nts3NsUTKa4Z3Wj
PtQJH7D5SlxaeF4ezOulMIhuJF8KY1+EotIdCFrKy9cd2EiBXQMeT0+LYBxAcYH5hW0Mn2z1zK94
7x/oB6qNS+7ZUx3++I41/Inry0AF9s9MvXF8+D8FHG/PvIH3weLkenQusz91VUFtwNPBIHC7V05P
rhvwjMu5D/pf+RVEIoAW6mFWnXavVh/y4paVXFU4b5sc34z4DTGNnDec/Qc8cBeSRTVa7vJohLli
uMbRdeTqkiC7yoXp0KdyGdIJ4h/TjYwWrJp8m1o4z1SJMvHPoJp2lHFQWQZj5m+QongMSDRDvZz1
aPAWO+jOtrfSlPzkm4MUSQyy/xegaSDh8/tXUai8hVvyIuO1PfAy7aggrq0wSMOl2ZIIOMMz6di8
vavWz2fVUVDyKl8mXFGOe0f9uoZ8uOF9veyLFK2ylmEiUsjZg4hCzYL9IrgWlAV0yr1n8wthjFON
VbpIqi49oqxV3e5tDKKJzNjolK+CGjpF3h5DyAa1KWmmUZvagm/8BHZtWC6f0fe374pIKCDUdipa
Cz04w1FC0LznTQJ0IDXR40QseG2Pb8IOPFFbr5JOkI3EBil0M01EGBA4b1msorA2L+HrKLA1yx9G
vy7ALpzhn6+Vz/0Dhs+dAwv6XlZWFLm5EaqFenNzn3zxrsullrDTak7KFTIzK0BvSyxsVOt2Gcs5
VPPoV03Qx2CM9s2b6PJ1NMSn0AeggfZFEFeuUB7vmPavYxtRzIZxxAuDgQUgoHgHxs+EVkk9dB+a
m6IxOnZ7SwnUgIDd2a7BzAsM750H26wQA9zMZcvHCHpZe56HF8EYxzGkcdlleG9nx/ezAZCmFJEP
2NxkmrzjVQjI2Zuf/w+NGzXf9086JWPBfC8gAhH1Al7DhkDZYfEB1lqYJXFsXK+3RmLi3rppIBwt
0fcUKZz5ARtUWGDc0gU4O2zgByjn5vKY0YSa1/ARLaYdjh5+4kBY4V7k/keGIMw4svHozt4gL+pa
/SVSt13F70AsW8QLcfx5zrzYfxI9z8DU9VDvjhyey/L9yqLbgWQLkeuBLqwFZ+1UD5G16h5kpBMx
RpVYXFoppv5zk7Yc2vAep2Aq/lEBkjUM0HwlqcOJlNg1WkRZNqhdJu8vVhq7ttroPozxqPrSGuVA
Cy+FBedY3XCOZ+Oln0+re298HVX8/lXwCCp5Yd0f4MZhhGdrlCJh323fTWNERQRaCh4dzYWeE7OV
qTEeW2NUIZYQQq/SMMsERe3tYbr5chDikmYIo7x36/2xqxSCi/mrx42hdeTDuFUY3gwD27cNDu4c
ZqlFL0Xbl1FsUY8qClY9r6wQtM/o/Weuz2j7FSL1TdHdxAEA8Woz9bun6st9zkos0vNRus1sIf4v
vQn48qtfTh/Ojnv5dTMLP4DRrzgunoIkcI4F2DWgOctWvOBvBpHHKGpoAuT+blG5grvLQJuJrf85
ALML7Kz8d69K4bR3fW/0ltYk5Dnn0gzhjN8VaKKatSmIemBkPscPRQ6Rk9vlKrJ3V11XlPAQhewI
Xvgd/vxFbsjPFMwVQzVvdw4coxWe+2sTB64JiHnPSvQpPNXCe7CAjcHf77msjs8jVow3OlY+C+xt
VKFboHuPQ5dc8dYIi/u1Aa5229W9pNCy/YEfaY/oU7d8rF2hBPatxcS4zrg5GnpRJac75P3OVYCq
vcj+fVcTAzGszBWHnoicBLkSG8LrGytOmbk2MhzrrUZUFJNaP7ew7LYpSf3JokByAPF1DRY87035
+gngliVoP4P1ODImmwVrtrwKplkC4eCvQX4VsAievOIaKZTaO27mmiQNStf69y2yz38tTkoQLKEW
JINsK8/zoifdgx7guLUw3g7fZcXtQFwv9jSTZJokrex5GPwF8beTYcqoFeFyrlKHk3maG+/Dacnb
lU1t+tnYDfelvrTx4/u+99sJsL0+Vh0XN+fdzrCPxClGgeBDgw0RcgGrVrGuH6TDxrfyUCOmQ0c+
ZcymaEhKAFUIRQ0VPrQXTIFn9oGa3b97YQwxqDkcwMsMHVdDejW9s/H5S77ZlPMNtUASApYRvjmL
eE1TUVzWCZFasvZSNB5PdlR8Y3U3GjwtVMWx38Fa0HfM0060QCTBLfarra4Y6qE23RqAfrABEJDN
t4pVnTt+1Sykjpx181dO3yH3t5EsMtALp4K91nnxelou4QfnTmjW/hQmW0DkI5bc+bbxtBa/wPa2
Y/DGKZYppA3wGYSJZa6D8Xog8FNa+5h7+Uo3ZauxNZfFnDymj5oiMpWig2X8zavN9/w4Q070xd+e
Elqb1+E5DveUAMTYmzfU51Jp3IuYgnvi2WLpk5f73tc/XcedBpeBtjH76nCLE5bKRNRG3T2Fs/eY
s94vkEAGn7Ko196VVbOTuggsl0LN2Hqu0T4VJF3vAEEsaO60Vi2hFtVumdkcL1axdHaBzqmrdsqp
bmAkNl8aXwCbcLEogsD+DOP8VnJ/zVEDQTbYCXENgjXsLGrqhZc37u+T1zD+HkusphOCHBz1lhCs
fGMd4dtq9y5ca72bDILTjeONdgGwWedWdsJD7NliuZ3OgNFRj9BFZe2J5AZgnDWt8fC1XlEdCkWj
Qqd5ptCTSwq2ga8Gqdf0K/xdwnAyOdbOauwIF1eBat+vmGHENlbJRFsJo31/rMpWmHze6ecQHjpO
7GFbXZY5hF5WP3tkXd88Z175nc7t7xjMJs2Us0c6LD+NDb/gkvO0T+LarciucH9wYpZzFVKlG5gV
xPYl97ewxnLZ+IA4VMyT1vUG3HCic9KZNf0TOWDKt9fRS34moyrNRq6bxchACJfBjBs77iXuGiJp
4aHLRDVdp3eT3pIuhkC9n7+f2FPThPBepKTBDAsQwnN9iVKHxFJoVGnf+5LIEOVyuZNDqYoH8r+C
bDSQAYx1gwuhRglqIS7qR51MInGztsgtf7VUC4CqWHqVKLvl6bJNG3EurIf4zeP8ATTCySK17G7K
exQYYolIFrJgianlc4QXAXXpe3lC1XKVxXGKhq0CV6lDr5TLHJBrF/PcA3ptODGaaONOcshtpkZh
1ls5IQTYDulDumH+Z6zx1LEydasWaHkUhkN0rcwRSqVPWu389clf0JhSB/6ec72O1lJc8oS23vbX
6GW2qQ4Rtm+tN7rSiPwbbplfqWySorv3MevObPyXLhXeufWSXdYZL2y6cu8C/QqfoJB5Hlt/BjeQ
/GimnyEp1JMcfqYfe1jRqI+9b1GF/KyyxiR9a8RGgH0CetNddXC0lMRlaj2o3Rf+WV3EFcjHS3+z
qlKXNwCmiu9DBWYZ6+/cWVH7edG5DNOWQ/MIDPn/itA4GKVGtYRtfFLOHD/gj4JFFSyi7ioux3gs
I6qW5KPZrK8dQir7ZW3gWJrui631gl9Jp4dPmNJV8xcj2c4ApRTfQfxU7R+vNhMF9nOu3rq+viHJ
WHfoESb5CnvoMm7Sg6V5TjigNws8kvxlTG+13UlXNd4OZsmUwPjNPsLy8CcUAGJeRBGvtrwofPEi
FZ8S6P68C06ZTfFa2AJkAKQjXTi+gPy/lCr6jcbWMHMBnAkrS7vmfNVtcuO+yR0h/T0PXH8MD3bF
OmSX4ZkEcYy1WJNuEQhhOMPR+ldM4SgOo3QvlTEhV98kAU+2w0WoIjycvj0zk53Y/q8rAlw6N7U6
LObH2Q104JDBK5YQbCf6Xc4WXpCFFF1Q39X3CyyAFYU4lWCXuJp9eXj5pGXf/BqLAEhgE6smue2X
jWutwp2OejcFmOEHqKG2RBr3gdXq44zey2XwqvAq3tef7C5+0gr/Kef9gSr8xB5F691PTh4sARz3
Gm1qk0zCw62g4PXHiJXb5BDduSx9+sHG8ztkKCvZvNxzXuoh/k6eEazkYOIJBkW51w2mjEOo891k
Zq1jTf3EU5XhhNIEifPrCvLwr9GfjGT69Z2W+blFYfZs7ZK5Cd91WKDVMKb+yW6kRYO3jYonUmXP
DZr7zxIwsL6g80cYRhMp3FQLzFWtnAOY9RwNeDAT7HQIPaVOThSk/oyl3uHmsq0PL2Y14NH2PQS4
S3mRL97PKgi+wS8TK7i0XtpHwchiYAU/5ZfnmHJznaM07/xCCHfiz9EOL45XM/2xcPPTfYW5kon3
vwkuHVhZeGt+q6bhNtVfrxK9L+tPv0hL52fszUirbx1t7EkwNJBr0Oi76hR8fLylPkllBNS07HgL
VpZDKXlQGSARUy0JkpMSJSKszNKUPvfDOEFn9oABmeebN9QdOR1Y2QZ0b+xdpeCfzFfXtlVMv4V/
12xyEzDd/SEEllb1B0ndJJZzHkh0sgWXaXJ/rnPQLJW/16XhTuNJI8tSYrmvNWzRJGwi8UYiwAbs
keSJi+78eK6WwOJRdHf0rYKEPv8gyH2bySSwD9NABddYgI6Y89uCcYji82XEIRHZ3ifqADMkckAD
uSB0KPYpWg+D2Gns0qJUpPW5BqbD/gTxHFqObf12pyaNF1/ySybdWHyZd3KF0RLZol0Yfv7VfeiS
8QbRURepfOfNAsPrxzPjHsIbnDJDEtkq1cmRHO592gctuUBx3vXSnHo1CIJn01TX3kJVxBQnuXgm
2ED4J7URIdlukuMyySN4hiPmf03fPyBtUljg5mtGwhwLfKC7XDj1iANSg0BCuUJPhDARa9OjUUEA
sxDS7GT1bONm1dv0jf+D2bDE4UdxKL+fxJboZ0N2+OjUtbogvA4JgCH8zNACyD7ccisQswE/cMYi
4i+HYR/WsvVQyxuSVi5t9JSzzWMvj8VEMiKDiBMGY+0P3Oqe4//0qZAulZ1bfKHK93/eh8w9jIc5
mn1ukOm2Wl7Hr3iarU8mW65RmDEJ3HsAeZ/3WZGM7LUUfK11zcm+XW8/7ZN+1jFDQl2pW8cunPV+
yY5u6GbJyy37Ls3GB2u4ibWnZefv5L/c81od1agA3EkjDMRFgx1fREzm5eIDvGqdht8JQG8aJqkn
IovYGXcfaMk0taGDBVvwgOh1Ib5z1g2V6Kj8MAtYn1Cyx+DfbSbsT78Nx0+erUAPD4KG74ZOyjPs
Ak5izxXeFD32NN4NI1bBcp8kSf10+L/LW92tQGaXCnLVGQGstfmeSkScRPUrb1NlVvHpsgZW3+5j
L6XAKFrgO1VdnPU+Rxr1YHNBeM/waaIvNRxwD/nHa7mS8qHaKDREaN0fjA/Jj+BniO6Q8w4JHsb3
CWnznCTwvYuy+g6kG8bZAwjIov9JpYWx+dnZ9Of5E6DlsYH+xu9be9396vI00iF5aHVVZLnzeCmK
2QCQP0TDRW99SmHXX2pkwgq9B/ZJ3WDvuVm7A935zOBL3eb7MS0nlWfP7nLGHKz/HrypnmCo0ZYP
RG81bWtuB1T34WzP4KnGVCpqkeNNWOV+1B8g8Vh7j0nD9SL0j77aiIBucidtQQn7gvGkjg4tLn06
ov+cJPS8YQTtzt5rOnXD7xu9ej9BCAJ3LAU5uU77cI1VU9PaiUDKawd9yXP3SDgIkN6WAi7hXfDq
kVlIwzC/94ieFJb3zP1dNW00EpGe0H+91j1SDjGiM93v8auHRNZZSdMI2mP+K+1yJKk1oVqGFP0G
2OaWs72YSo4BOTKmm+WotFX+Fn9cgCeTVy/sMhiqc484oDJWk1kHJksWtCoqiP8tz8OG19467QVX
rC5eDC5Qnd6YB4DzeHmoUS2lqVMUjyKylhLNqAhWtXpuHjuo99pCa0MWc1YOxB7guCOyA00cUlxX
Y7RTcU66ze9vsbEedJXjwojuYzdOoNpY87jr33hZSN9ESIktKHzZBZeHUCtUpLEi7GoY7D9EFfAv
s2w0600zNSMnhrf+b0yOUX7IhxCtJjPXf8TB5ztDwcssvybQk4D0ohVqEleavmjqEgU5oJT7TAIX
GSgUth4HsNZXSMBCWp+6T1SAprWqZv3k7a6mH5/X/87eEacFvra4QM2+t6W5jdaYBVeorCq/XqGy
CU9XZW9m4zDOb28sICdLQcJlm6SVZtOM38YjZEHfXnUE///a1YpF7xHxSJdh6yYECuYv4LF4iqb3
bqhawTue3Iqlg0T/QBAHVQdWC/+9splHoNjfdAKh69aQECTeWr6M9/zctGL/eimuNvoSpxuQGEFe
t4bVJVPJEyIgaJ5wwT5yzFt9+gOBbKinsk6951ckIoMphY+0m4KPXXtKL7uZ/ouPyKQe1C0+rCXK
kyZAzisXsCUsx0Ed4FYUmSsojTfxXTrHadOZRk+NAe2UAN665Yz0/8YUD5hHk4l4BdCnJGcChCYU
QAKevfA0Y5IdtSilctMcpY559iUPg0guAmOFleALDGzO6WXPdAaggFRPH1mcnF7K+rDT3eZgrIOW
8eZ9fWAeCvvSNEclIKHvBiSzPTLGwOpvtSI3y6N1VLd8sbG1YK5btSPWLZh0hxeAvTTjRhaox317
HK0ysD5cuynOuevbL9SD+ZwLOpdQKCeIf0dZxVy2ssfQF2grNdug07fE1IX4OUwnMHgwqVmNltsH
P7Z7/ShwsD0wKsKumu1im8tvNPuUx7ntwYin0HgTrihuOxnS3IHbupyQjbE4OHdu3RqSpcbjt7jF
WieM2T1IZlDVrR6lRp9lalCE1iEdJ4veYQTiWigYBRkYbRBCjurtohJi/e5LdJzvpebruHlAzAbr
AOESzcZluz/Ra4J4PCOgt6iRNXYKWz5iLIN6Z86MXn98Vwx8hgeJeO3xZomS32D0DVf93SCiXXv0
o3hh0i2aexXiCzY6A1UZeu9pB7BQTEHyMcMebMa0Tnwkze1jLVjTzpWRAetW9SUzpNjDnLFhyVb2
oyqqawMxTjJUdSqr6MB8c4wysbSXNHm2FZWHTlKVrw7eTg56h/DTz5HxPJ7FHd/UU8JV48bygcTg
agnTfcxZY2I0QZMSj92qPnBqU8dlOUBR1A8d6gJzRCEHSvI6ZCyDqsC6rLDSIGJ4HosaSghrQqPd
fcugPzacuHX4wnLy51UzGUmW7Nj0Ex9RUmztLTZ4yiDhDvCo3D+wTQI3sBbBPzQkjSDO+Emn6S6b
yhy8lI7px15HWavJcyDydaskukpXq93VEm/8tuWbPtbizaP4mBfFuwh2/tGE8xgEuxQ06bc0HVoI
E7IOonQBSYwNnJ6h4e59XZZ0xN7UpbISmPJmM136NImqWiOoZWDUIXQwptp70irIRz2gKgbEp6Z5
YiXCsaVTOZi+ceOjc6BIMNJvBeuJh8iusVEx1Z6m8ojBq9d+BgtRO1RDgi1sSXKzh4LWbVXCSigZ
lOUnq2UTbvyHUJscy5jR9Au32lBTkpaER0QpoCex6Qhwclr3CQd3lhomfCqFpkGDcQUCT6nQjobX
3HiKABWL5Om21xrdBnYpl/LgtXqlp5LqWYLNsFbozvKQj2lQ+SgNczBXJhnWxeC3dS9+RquAkhkY
ZxM/EVlNYHA9WX9w72iqWz70cH2N4E815kFqtPdVqG5vT3giPVZl84t30GFZfUfe+SrBkY0XnKtM
qVIBajHzLbU7qZpxAcKskBASHa2GJKI4bac1pDuTrZ7ziSWx4nWcFo1zq4NvhDiccKW2br0kwiV8
Y8FgF+R2adZErM9HzBHS8FvcdPXkW43PHTp9aUf57fOUf50Hp7+Abyr3qjxx1tZ6mqT4/wblaMyL
1JVHcN1UNej+uO7G44Rjg2VOmSthgXn1qo1/8DqVjR5wCJBAEidCZl2VK/wZjklj7IQ5FVJ2+kQX
dhBb+mp4kMPqbvPj//cIflGUxE04yEmhBK9A99OpHiTCXc5DLpzRbSTSURRgMetjszXNAHfqZUe6
2zo+QPxJwL4N0DWzMliVYMiEj3xX2SDQvCTrQoTM71WzzLhnEWFqfe62D4rQ9o5U5nwqlTqE5BIZ
6CqpwtSU+xbcS6n+/2ayyEJYJ9HEN9/l/vvjHAXSkLnW9MtDVkGZ6SOPBqRfgCjqtzfV3XVtNyw4
siJrLqtFn5ZlMCEPqce0gCwU/uQ45gtwX+10GlGZm/et5VEcQr2NAaAutPebGfIBEQ6rzg3ohR5g
3pLnmxIqC/6jQb3dZQw6krdk2FCbs9YD+ZA+GaseaXt+/4Yu334Ewx6AD4dF1FLNpNbv085Eb9W/
pafBtz79c7mHvEeW9cYf2YBle0UFXmfnBgR2eMAy6YNPui2SgulRChlyAxfoNHMKLCNN/nVohvCQ
F23o/eceefiNEAya8Bc2G6hpaPmVLAzldq0MYUeV/483xrEF1/9/252wclE5Goy9pmHZjIv1Mzrt
6N6Ec5DmhLK4k0IHH1poJzGDbOV/no+adGHBJVrTysDzN4A8sOGxEraYBDu5NoXJ3QgXAD57rwvX
uCGGNUYLXnON6mvuhXzttubhZe6kPfePPftKZtW+fVjZE4CQXMvFylgMQzWtAO2qUtbDzEVd6CY4
0aGwmyBicAbgNLvObNp1tVhIwgl5x+1MGfCLTsHbcJzW9s0Loz3d7KTpJcmw/t3sCYdOrOaWfLXM
jQYE1zyastjpHchnSwXnLVDARaIs53Y0zWy0zcAa6wf9BvmiVz2+o3MF/bXcLWiF9I1uRvZTBnSs
dyWZpsr8R+eUHDYzniW1guGqh0ACp6u2n9+Gxd5xgFtzTZcOO8bYG4FNlFqjx/gUpKmYFXZj74jC
VTKUshRIuoOSih+9Mz7I/Dvcl+Y1Z3vFuS5fDZEdNUQUbK3oNyI7mkejrKMEP5cVl+BrdqoClkIA
w/W3/wgeKu3PR3zD64USMwSrSOSOvr9rZPlYKU8sSNh08UX5WDs4GxrwXAQdlO8kkvL/i5OVynEx
JSzT1nto1SXrymX85rpF57vYAv5VvY3extCyjqcEK6IBMU/O2sGA7Pm7Cg43EbnjLKz6tXmZqF8+
3zrTmr8CDvdwj3AAkeA8bSqgczx6YDWHHdQzs2IelOtEB48c96p6Ictq7mRfKRyUB2SpUJyQW3o+
o4NdRb+vQlG/lsJPS9dpyREFOuJAtaIMJjW+kxMVvZfpcgFadtma5YTvny2drWpylVEiDt0n2eI+
dvx4ikq26nWrQFkJX1qRUZt33vjBCEYYI2dglWWTWP8i0cKvWEUBsWda+0m8xPv2+KQ5oP2CUTFK
Yd8Pf6dL85jIbVza6GqqlX+CewFb7+JDLiWED2MjlcJxcUtEEyUrWp+Oi9qIfLWM+1hwQh2ZOJLk
nyeUhfDEurbI/UU8yL1tg7k4RTEwnmHYaatJUS0wquT5BjLcJrol07v3XAipJLFzCfa7i8/7pu/O
TBkVFLnUWK3UiBOUKUFOU+LlWFkIe8l/Q/r4NtetXKgqNSaIYgukr1WJrmR5WIKPDPnS+m9iqhBJ
yZcqwG7Jvzsl/QqCK4E36bqUxSQAEulbVH6sCQEmK2KhUYe3Kvbqs/hApa8PrRiGn0mZd2UWw4t3
XU/RZpuR/3WgeKmiBl4Uw0MLVJL73a9ztrS4maYZOOpBPmGViqfcbpH0FUL62oQ/IKBndvkcBCr1
BXnfDrpCU8fZ7+nq0DKNq8mwHRvGreQG2IQC3B5m8Do/Jx1Wi97d1aTb8ER9vQoo37O/eEaFoe/y
hTUx2iZYiPcG+Nezm9ICcu1Ks203VD99mEGN/tgUIMUBueSS7VND1Ye1B+88Qu+AaMQmac8UPGUi
c/FTRmw14SzaOqJUACQhA3kYZXLEsx/23frw7o5gMj0xxHyXdn+jlK+sMnjHGzX33ROZC18hPN+m
ygFixPYk2nhbMXwoV4+lb0RNbWttPd/YRleSElPJ3M9ibvpXLDtzM6jIXX1bLk+rhf6/fDX0+Fx3
Zs7H0PYW24e6dC8n9DDmbYhyKJJZpqwVKmnA3fs05AeJTFIHmGQQOD/ZWEqWiGtcl7s9hxJl8VWA
ej8AqBlzyzEhXtLpZKwYk+YSuWP4YShLRmlbtqyogX17zc5Z+g9KrLMevJTPfS4Lj3TvScBC0STu
5mAks0Og3oyl55EJw+s/wG/v5ACCxJEZ14QSGxaj8gP97VC8S1yZO9hahqj8/o54H0V7vLZSEtQZ
z+Oqrovt31mdVbMqDoWwkERtK+cDxnKgU+VgIqZpdhTcSD8wPcYRdz4MzT3E9JZidjEg2f+Ag7z9
3sjGgPdjNrMByCJgY6rSG0/L2450REvytJgRZVT4zBlDYQYpg7FPYt21v6IfKEMAsQItm76oMvwL
ZFtMF6qEvQYdDpGB+LTrMYVaPykjbKs4zFszN0k4ETmnZeCcf9DCZ53D81R7jR8lkcV5OEBmRhaq
LKJwQTdXHo+aoSk90HNqHD/LVIA57QKDnwQsSptQkg0hb+DBYXO7actJL4jgXgLL2/Ik8UJIu8hh
uThE/ZCaPrYRNvjW2HaVr5oUzXQjig5HZNAu6ybm9ke2QqV+EsEZlGDTkgk0kxaFCfg/t+e27tTU
9QJwOGh76OCwBOUzCigZnAcTqwWdgV9fhko5W0Opu3dNYPGY7UYmcMAMLC3Pg60CfNErXs6K7shk
AUcZxhL5MiWWdWW5yo+pSghawXCAD+tvI+p1v+bDT+iwDLNyNd/hogu7yuUXrbodRE+Hvk6fqGdN
WnZb0RFHVCQBzUNc6xU33sCRsYn7MFtU2ZjxRYmoDoTxsfjXE1oFWsfjbmaYSNiTYrZ2PwwKSqov
H19JL501M/FcA5PgAcePNtjiT+Irau5XAJ7YbQdgtdhL24txwXGpz7iWfkUlwbVzSmLY+CEtm73Z
pzKUTg1jwMl2FDlY1liRsLqz21NJ4GvPRE0h8zX78cOu25AyHKGeT+NVze4vmz60JIdDyUi1AxZ0
zidRyTVhIxoGLV0v7LmqxpvNwTjkMtPBYzivr0uK4cSXi35FAqBSBCzlD+UNfWzAUX9dRu+fxnne
1RAvY/uL4FXOL5Lk7LSPX7qY9Mmvrm+hL15xb95sAAWUHbhsd6ghgUguSS2cEfNz3rN5RGMzHWN+
KKjn8BwP6yqul5XU59hooZLumVwxUugybe/WK/WjHmjevx6wXH2DD3qOvtHsBcygpxsWlxfFL8Kv
l2OnZzh49VrBf7J/pWhcQYymS5FV6axjqxJWfK3rl9yRy+J/I+5mozj+51H99g74EC1eQsj5fOOY
ZOm/jp/68FokAAhoSEyRrWQkcEwTmJpV8HZhyaTvOKHOff9o1P/ywRn1qN/gLWjCEaBdQbPTUMZp
O85sjUd+ufd6jTkLMRfRq4E266RnEM2+4TZ/+B2okBhvz7SXu1uPV1q38zxDiF4HvuhQbCWIW+HR
WBqnNHcdCvFu2jIa69VTY550mDQOL4EK5VUvtv8ffz+60ushZfvXqy8+0WfnFAVPZkDoLuQhcopQ
BbrVybM08wUYBMMTAzr1ygBo3zuBCcZ40tgupJG5fQCvr+DtRor73OeTHVkV4lTJn+rM9HyKD5J+
JNzd8KZKBErVT3H4NUl5i8uWm8JGaQTsqUmrs8MNiZN5bTJBi0+/hJfUs8ynCtr2JJA+PkJqlUVY
T5SOI/p7GJ7WSGjrxuMQbbJ/hjQ64h1up3bSpA888yQJbLz9ClvPJLdaOuChjSAy9J0NS1mPBw5a
t+omnC4mtPQ5z3yVuT9asdWXI4/s/kxrRHelnkZygdyNr8jZ9heM8DF1xkRB4kncq940RNMAHfl5
EPINJM1KMHwrkDFbbrG/0pvtQkSAfMUa4S6c08o6QKa8jwE3YSr43Ue7nuygDipqrsl+IvMlduj+
HYzPsJtseAnIXZNwlM+/DpLpOW9Qqy5tjRV98evmtErYzYF8QvX/8RjX9phFXQAsUGD35Z9KTYUn
V/bemJzYvKjuPNg2gKewEuqFCucI2cS24NX4v2w1xw==
`protect end_protected

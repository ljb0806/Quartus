-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FPcuP3pgQx9O+Kl01IIdf/Ga3jeC7sV9n7Tnsx7HkcgKTti5S4oCYUUnJCqgHusO1H5pRp+sCd7m
okEicY5vScsNAPK3o2TbK7j0/vQ6L8ZqPE4syZfTebGt3YRsc7gf8X7GgNICgPihCNFFv7aCupeu
OdxMJlh7mStNKSYm1FseQk7RlfL6H6jw/SxJVgiz18QHCNRonDVHcvPAlgJjBxVHxUnUsy0la9Fj
Vd8VCt1nWtzYBZMGWh3vDGTPyhjki5UwfM8nZdtU2X6xhWGY7XzeK0ZMrzEmjUTFimxjWJ6gqO24
wwZMj+XjWOLqBiULcHkQ/Gg3MKwbRf0aZipGbw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30528)
`protect data_block
/CELs1g99ucJo0p0GgllFBET6Hux4q9IIFqo515uRxLwa3HUmZUCp6sDaEK7Z4bVsI7JoId+l7c+
nYCmb65gDu5QOEMrKsNyD8/jcB58He8R19gq68R6SQYK6rTJkTeWYWlr0L64Ak6qIhD0rP2lVoIg
SZvMWDn1SmO1VGEBeKVfwNwhf6YJRUf2gWXDjvW7D2gGjutE3vZ/BV/oJYnR8VRHkrpapgxz0Rme
FFK3/3iDXxKuj5jjggwx3p7ZE/Ma1fmhm8s50B9lr7R7Q3S9iejVH4fCoxHLe9efV6k4KGGxQ4LF
MzfXvfH4mI8hjPIUf2M7BFooDb+iofNDhR+9Lgu22atvxydVIktObDCuoJsTjTZBUKT5RY+BNUo8
KWzsKSoDUuX/BS8NGSVnIWmochOWnhTu7HecA6KXqeT7b97QBTQLeKXo6xhGaBozqK9jyxucprJc
FlRK+gwxI0EhIT9cHYsRcOj9UZ6qZfKfs1/2NpUB1cD9jBOi5azm0ZaSHzKIvQdeEMT0Po4HK72T
uD3HPwkSyGg+W4xA34xHn4S6HfotXTcarwbfPeXEJPB+mlePQrcwvEYVgXiL2KDz+v7osz3yHAVt
pJ+lGro0Vbx+W1QdYH4HHxLxsJCm2Mt2EoG/z+IKTsxznzK6E1shMfphSt/esLoc0YeWwSf8jkNt
KG5ehjP0bcU80+DtWxwc3TmOxVo6h2vPkzAjqcQCaqB5RFw/1EjTI59pSPksqofYSFLltcF8/Q6G
TojYyEe19YzPOguI23Thf3ucZNSkI/poJ7Um2iTxJlfCfMxE0HJCC/aM3cX2A7aBmOduNDBHWWnd
MOrVkwBL1fj64hfg9SnobkCbeGz25W2JTB10SdIGX562p/etOt5QbWbDzGdtzt2ewnM0JaZCtEES
iQHMFzpv0PsjZCmaXMKG5df7qiUqS54WKMgvT8af8qaPNBou9VZILW5lgTIcKTOGx8Wim6pv5Y8G
AU3GXv5q20QjIt+vtBrqcZ/vt68zKR2TktMPmLcEpaVA7rIjMuBdS1qpwK7VHI7fHq68mBGlW1Vm
q9T9eU9SrDdB/cl63Ofm3Kx/zWdv314MUhbRu94kLIFyaKqDo4cmrVnp/xRGNgcKT8TTSjzYnqA7
J/SKASRP7Wz5iW+kjJGvfxZXZqMZKgtnSuvRVtOD4jRqhFx9j0MaZFjdgc2zPrA2fOXueIaqUc5i
yKRHGyApbGGsUTlA/rTHtTDXxY1k0jvBI2wYkigQq3DDpgqTs38U35V44xTBRve3NBTY2M5yop8a
limSo6M7s8L7x5nXxNaRsTTs46Jr2OYZhZvcYbDUAtdcxe8V/o18BsXMsmCNZPy2ezFhoQRCOXKY
2urDaH7bGRcPR2T28v95lmVMce2CuuELbc6iJWzcfOsD247zjSFqtv/TYiPEyG+hBH0B3UTp7mOD
rYUcyzcTKZqv02ab2QDrzQjZPuvF8jOgy9i/bWxndwvdtL0/EBUbBQzJrXq5bFK/vB2EzW4eyh4f
+jRLvpqv2coSxrHrKhd15QJsIcCcf80kbsnYNJEPqh/UF41GZ1ldyIeQc9/SQi5nWGAeJy/jcI5h
LTcxgK5PfXWb7ubl0aKTwF4FA5lF5Kjlkw41Dg0wyhp4z5UA7fddNHJ1DiZpN6RJHTY9069K4c5n
sUTZwK5emy7E8cuCEQ37xrBSjWYw9ezJXGuhCOZsVc/E11hS4NtWIcSCbCRvZGLzMTxT5y9MtiZK
+8Erp3NPc8+NmTgUDJ7r3tgaQ3/ETo73B34jip5+DTggi2r5WWGHEF8ljB8+kqc9YKCL6UmzFBNc
ZfRjeJ8MElyydS8//vDtKiBMBAjrQ0V7xRiniREC+Rie7tcx+Z/kanq9NhFrd1z4fBsbQSoeQJ+C
NJZjda6qVRFmJNC88J5A+f7tlB8xUIi+2QeULl1phxbg5b24wY4j5hkzwP5jm/LhDHzu/RlW38QC
SXm/Kl+RqQeK/GAW6UMzYCrQQUOHQdIlb/T0c2zXzDiXnRVfZcr+34653aVVtxY0ozdEUG9BNnQ0
yQrgbd+oAofAIZQ3YODYJI/l4TqaPHANy2QVPByeVXQ3rz78pCNOJsKSujI+9JQCb+KEBj+m33x3
rokRIW54EXgeHtQrcTptQWgfu+wiDY0UJq23TB0HbHgBi9gZFQ+t9d6UlgLxSvkViWvQpl3w6pzb
eHZGNqbrex7VCnBf7SieynUv/RasjHn16xVlqk4rzlwQ6WEOS8YZhL3Y7Qf16LTWMEGPBhoQTreE
ySb6N8VLI7F2nrKI7zIOBFAhigFAUZG0pjCpLlTQt+zsHW9gTI2Hf5vp6cE2Yekygz64o9qu2GH2
TS79vMK9Muk3CKxQuZcXNLAIrUx9cTtmqEqAeHMapfVdUaJH9LpWOu3yX7fSLprda0e2goMjSdz0
fXSpCJ0RHlCU0J200dy0vDQGveTPJhRyyHo3SDYV6cbLe6Z77p7JDxVXdMJ+FKQWL5boGJVoth9w
w6LZGvl2LPhKwLMjlw9S81JfFJUqK/Turh8XBUiRnBO4n0/mTQJWxeag2L1ycKDPc+JQ75K2+ZCO
Q2kJR0EXTWfZqxGrZ0OQWjqtKO5MFP2njQz6/V/JYVJ0uuMVAL+Pivv7cmbcx6KeuSBhEK18smK7
OmWCdFhIPZlQhAQsp0aufbVvTg+AxKPfuaLiE5jHCXt/HLAvLCbntPFCoQE4PxTzlPQZVS33/xVC
IBVu75RMazFSWSl/otQnisucLOGvFXva3vqibZp2jzCngz3x4RD2DSRR2nB8GN+nzf3vNqyKv2/N
9fDZwHdxST+N5O0Dggbgso1rC8j8f0oU41fFsfhxilCTX8oKuu5MFaQF5SpTjX0YGbnfFTC6pOev
UNEoSrMzp54WR7gqpVgJjvv7wvLJLGhhc8m2e2gD6kT3buY/Ngf47fNB4egptUZyR6SNEkNe/4ls
VSb9TuC34itY5L30xHSpAraLWjCxJojF+9imTBamR7Tvj/PJvUXX2O4KNlB1corq9zhpvUWC6nW2
xk9BPcnRFL/W5oovK54Qu+ZyxiFFKgoIPInbkk+as6aVscZLKmBe6Jwj5KD/KZFuTLaOXsex4uUV
CyQD1aa6x0xtKYwVw/V8DvjiurprVFVTzcb5sphPk7tb/407Abacl+6Oiwwqt5ULroqJB3JeRm5C
iVx99nf39t7bE9xCKK9HvAodsOZtnXqdlkC5dpAlqmZAW3imhUP0IhHa+u13PJMQy9z2L6PcDGps
/mI5tagHDDTQirap3ks/Es+9nVvkIIYRummfZzAjokvhpzep06H2E0LrOvjpGdqhso/b5BI8Gex5
WfSX+FigLUPCIpOL6bzAF6Y6sM2Ptv5nuMnNFZCKqIe3JDFBjjUcMXnn/fjSra4PNr0rtV+KTJz8
oQZkG86NNQblX3q9DoAzxhwgoZsshxdleFVLGJTnKAvrlSXNx4GyNXBxxU5z2RNh9d1cI2bk0maX
JdkVd/sw+gKMWlwKom7TTPt/oC3XLuyBCKFdf2aUGBxq8g8RybgEycuMq8xs0bG+AkuavqHbC5GL
GbuzwqSIjlN81aNviEYYjdKC+jiIAY2rDIkULKcdnyJII1RRTz0LZ1Kp6P25F2bo49tVaLJcMMea
wlw8ds4RRiSwUpU6XTOxdtU6olRwYMSHJst0rX01zFHHR6zB30+ngd4wb+RS+jK+0VeP8CufDLNb
sz6jHA1aYIjIf8TiBhDxC9wMx3MlxNDqBrpZOnhXjJIyR9b6vnDpvUXhFSGDrHuzge4DTkR6PpGO
oWqN4lOrngIzYQQDyWjfgLDBjrr0t5fV+llxIsVfDzTbcKGLwyBpPrsTR2ltwIcS6oyDyKEo2RVv
2JlpdJsjUgxXVxv1MAEXUW/7CTHxP6mEbHKNoQkY5QJx2PDyOfrFfR7eBiicsy/Xi+FL9m+GyQuf
Kfrbw/bVLtnweo7WNALUOI1oXTbiV4E388cN+BEP/ySFQlw8gLDNP9+pVNo+kuDjguUjOwHaX8b5
1aJQTwmvhAKM2537mSFUczMw6UVJBJc7dYkiFuTiNeWXhQKAbes1WW4n8/5t/A5TvmBG4t3IGoee
4Qu2TXoSmjZEHMlpQmejWG5YlrJHUyiOsoN20SE1iAwZUPL1Ew0Ul5Cp/sd0Ce0xi2GgG9WkAsNy
XHFv1551IVYGTeuJ341SAO6eGSvTX2a89UD1cYCd31sjuOf5evUwb7Evhn3WP0N8K92vfS+o+SF7
Le9PH7LndlUNQUmCQQW6BrSJX/7T7SAMvINzLDoTdSBAu8bFh6HlweGpb6BW9Ezu0duIyAdVBgwD
l3xr4C3mJomU7QI3iEo04KZj2FW4Ih1L600UG0pcSfY98GQ3jaz3oEy2ncDxRWJPnIq/k6YhrYfh
tbgVwA7LMyNNoLQMTDojHmdmhrFynEjaWRMCUqD81fKqc7a+fVfBR0enFbssHAExs0iFH8t/LueI
/Wk2wECVjOKHFbQTdxYpJBJDTTDPQyo8cEaxD1KxEoWNkrlFL18GL2l23beXCbYVK0rKkSmw7Edw
LPRgOXzZHq+xvT+I5fggK5bdTvoVxnwHa8hytgJXot4bVNwO1zO3NTvznL2WByJMcL10LWPH+bzT
4nG9W6oqU21KHCuyzYijohUAF6+zSnr2uaswOVFAWmKHhta9ACnSMVI9M4sHridcRR9m3u1jeaWN
/p7fjtRD4ifconOW55LzVaRQ6394DZvLaWebIPKRFddmzeet5Cm8z4wqURm6BZ99BQ2sdwTclYaH
sE0vfK5F1l7HN9jU7y+0wtLMEum8xX+XRe3xvvAQzgXk1eTl25g58pIinSdyCqABkeJwjfv2FNG/
cH2pjVlQcrStkbx6wmnzMJFTO60qEpCI6Sp3gH2cyBr3aiLJgrGz2xUKXp5i876LZzgoPGAp4Y0n
sk2R4kmH93UdxToAZW/8gCfdpwAPnCrt+A5c9Fyzg5+L2msYIX8MzA9c2y6QF9edk5YUSzmq6T9z
h056Gd+EZmrMiO/omke3pYBNYYBy11ZqDKacMvVg0iUyab3EFnArXTXlJceidiKqcqvrZJn6sBsv
gKOGqjwDn3p/JjvWuB+HdyJO+MMO4ZxRj8BYSB9gT77Cl/A3vqwIc17+dk6fbukjCBb4cKevcm4L
Ghk/2o9CCtJdJBNbHFhdfI7bgoWyLx7F1AZCKge4xLxt1sz+HAt7ImwQUAOvZvK/jOWiDRgZhSde
D2beu+2oeJm4Yl928EwVrZOx6kzzz8jtenj3VxYRUwObvscdeXx6uboSsw8MLFoKBpPoUCwffneB
M6dxqoHGcflwSa4nDvx7Imxx/8XopCX7BfknaqzuIJ0r4k0c+o6RV+MhhUF9MAmOWX19VauBFs91
7R8DgnA9MK2diD4U0MBpc1+OrAwJKiDZtRjcRVWil1RBDRD31IEkdkvCcbK60pCNyW5ysiqczoVi
5Mtq10qFYh24xe2G6esbQOEHV/ZxI91RO12xeKDlOX5OYDfJbM+R6KaIUNQpvfyIy1EBPbpaivyF
G9sAhysoZPgJ21kbaMwNmivyE7/cCm/eqEyJy5bB/9chBBdXNseUjgeMsrw2PEK9Wn4apZQ/KWEV
DbCMdSlSOs+uoUk3KJ+Z4CEkaRx74cNxz2xEAgux/cxvLhCIomA25ly+Be0+6EgytDZt1uXl1kme
6jpMxlN+0bpZ6BX8PTQCoW1ikUVGDLqDNCzFsfffErUyCog/jkRJgyVugRKyRsoJ1x4r0ThhP5iQ
s7gj2q8dVZl58nlMb5eLBow6lN+FGKpwn1NMzFJ/JENwXqvr0o0AnpYEnMNgXNDwqMBqwMwkTFMF
IXOH/SqYYs2NTYJhezNlDkXz3YiR+ZgA+NTHo7EdkM+XbbRvS17v/Ri7yB5Aoy0DXbpKXkVPlCzY
L6mbhklv2BQ/NVpFqZk4PCihDyqBHH/IA8kthry1vLPMsArhqVtF+Vlkvg936n/HFcCnvdrWGuxM
LdzROuxnyBdBRs5M586l6xQFzzrAiW/VFnrBStPJdTDdSsSPCzUmTMj5ruFmQc2569GR0PmPY+cW
Wr4qlx0lUM/+gvjIvxxfQCiw2Qz+xHRgwa3rur/48bcII5+ryYv7Dcqu2RwenbFTDk76g/p/UvYo
4WjFhYqvtKkVoxRY4Ug0nnbhdDP6MG792XsvTSNeNCPIDtMCrrDHCNAb2MlWPBXPSSt2OxHNcWGq
CCEbpMlShGnX1RSXPt14otZbdF5R2KbOWsYJxMxdn+WlO8nuZLQ1aRAUc8T2IUfjf/MnC8ajr4m1
rfFkOt8w7VRH+7HlKtFfkQ2x6BrjJwDfubUzONHCHkszGy+49NJGa2ImaeFC5V4EAejxVXgSftRR
X+CcIZKKCJSsMsxG3ZkIRHyrqvFB+7nKeImdEW+PGSmJCWBiHaUgYikc92BEW4yWAOFZ8evc5TTf
mIjvu1fgVmmrQmvadgPXz0hRbR0KsDIxoqEttrg0nKZZnGK3EnUDrk0ZAZsOAiTQGEV9CRcg2Kke
hoV5/hSS8SXPFBNk19bfBlUmjcbAFwP0bj3LqSNR1/nudZPiI2WEsp9VVNko+Ci+uCDLgsieHQBT
kSeZmXmtPfH/IzmwfHKm0HtTsNmr9YdukDSHYxZWAE1lE0SydOCjj+i6/U+mYQqf6boH3pjN1WuS
YDGy/OSXB3LNbH+FNZqfHdYTWiXr+j/awjDJOwEfQLeBgGO/lI0CVFhgcGJMH0kYqoama/kWr9/x
oyk+pjhV0OQYL8bZbkciWRwDeAeN6Uacoe8QcTLGrKoyF8EOCJYGuzdtnV/3z8wFosFQqeGCyGiS
s9Mc60b1L3Ng3wXqmyRUCl6oPKqx32R3MkiDPwrkPwiWUuf4c2j/xXBLIy9kFvENfy1xlo9cAuHp
mMLDeCt/sIRlyNseJCpBF9KmPYLdHWQ7JN/NpQDYyAuPbswm9SIFqSAdPNZ8FAIGigIBn2TDiH1U
tmdHS/xRwoc5NglQIY0YQMcAru1+NQu3AfzG8NwLvBzT/vWWLPCRYBfG7O7kzzn60USNFUaAk2zm
MvUYzibEWvhstKKVRYpk7NX1cPWKBJwAzXdhFH4vOVxOcSWCHqH+Zj/CNVXxtk7cHQH/BfbpkB5M
msSy5JdwA4jrrnZMG655hyduevb0E5IiYi8WLPyjTz0uMaoHNHzllD/uKheyby/La4JWLc91+RUF
iSdubPtWSb20Gk3XHtkX/J9XJZU/gOKZekkEqQEGHWlwcZ4Nq4xAK40QcGgxq1KZUX27wn/mHpcg
TSvdimDsFcOl4ixUQVPt/M5K6Ln8WwmG7otCdA83tiu8tymjKtkhvF4JpBX68FeUf9oYFirqd1x0
55WpzzkfyjtUuVMU3HGNk9gDxGSdLB7Uj/dshnw0s21iGiak59ylWBGWbNHJNq4l6C79GdCd/zlk
Pl0ejehxzwV9CEtoe1TwYNjd3bjnjgMiwwcjc3Gh9nMnrgrVuFBrLSpLUKkqw/BXmizrhrDeRv8G
AYeYtHVTuEuhCsurAKSxVK6A99xXysgLwpEdLcybXuFgQ2Vc7lBgFouf1+d7K5oZZXA8/Jflspjs
RD81t4iq5SqYhDQVjo3EWXyjC/BXzv40fcZ4Tj6YcxkuVJpWF1LRE9kaRSh7Idp+8oAPbbaocX05
XvQXkMw8j0kXLd6tvCiYqt7KFWqSi7iKXsEV3P1asGnObjFyqyiCZH5FjNPNUfwUbm4TH9baobKo
uKUUORke+va8fnBz3tQNplcjq/Ay2zyxknxv5LbJrgj20gGeAbdygr9YhkdfieAffbNycr4mcuR+
NdkG+Rp9CEtw/pGxaE+vtBt4gffcM3xZD5Y5prW2bjrmYKPjWlUiSH3LAafF+e7bHt2PjYJcPPW7
RuRBBaCD/lnxLuGoTQQ77nI2Bgg+Qhcy1bJeZEX8VnfY27s4C37Ya2qebi1f+ybotcmLoY6gTxwq
6EgOgsvXnmc22rhIHYm7ePh2tquFQMJcC7z0DYQdPbHNZQ9RK+0YpIvRRkhg3VznqhGzyVpf8oyv
WxETUmRcaxYkJOQiycbLY8ecONqRf+MlGiq470iohLakxQ3LMrHb/ZbLjGjPk3QSb4v7zT4orspc
U5+5La7jcPL4ZeYFsRD0isLrrOagpH5SpuFGb6tTwFCwyDpVrJnDaAF8niqH/KXtJ6uYX8FbhAe9
1O3jnIsxsBq6MAkceSaLs26tryYVmLoMJD9HjzzkGKLaqmr6MpNe58LAvhUB0mLGKN1I3imRzyas
wHNWMpWHPLgYbyq9Owi/HEnSNaCtZkjBiNVJT5kNJqazqQXzHlHTXITAjAxPICRkZDiR06yxB1yq
I25R2rTuzrWZa8kjIdzhYQrdBUnLz/nfeS2pkyq/QlSFJNvz/timydEYTiTo52Ewy2spY1d428z5
+jSbxkAizmSYwX6BiQSjZ8lFTpqKtJa4BwAs6x7HNoSGuSlfIztjAOO6qoIYIVW9Xngf0rdfIW2i
Ysr2xLCZKjtv4nwQ71YYAhsGYmZEljuDVdCV1Vkh3CrBahuvAXZsCgswqrtOYSCt8thtQCLARMPX
MDxCgFUZYLCyUmsrx2l0IuxkSQtGm3AXO6QwneT3SKTi8ADijyevU6PPOp71sIeUHs00f+zOEPRv
fVYTE/JOR380nDeLASI+nsqFMTDqlUmmU9Xa4Hz4P5Q3m1gRdyxN1x5PgC+hy/BAlc1trTzAJLYE
Ba5hFcVyc2ARG8apIGGIZyrNdPt9O+eFN0Y6cjk3vJQgyk2WgVRCk/XOu9UumWIF4Yg2uJKtxCO+
Fv+Gz9qRt0mKjK+rqtJtGRD7MIR++kFeT25Vb5FHzrhQXoG5PtIiXdofduPXBX/fc9YS3/YMyjGJ
fgkOEW9KRPwD+yIdyyY/6+v2ZQBrYzX2chKfQlyjCCdYm7b5qHnDSQz54JbJdaFCPV4LZYe/lddi
j0zR7kV5Sm6eMXTXXx20SKjZLRhOCQ+v6vlJdnNA4CjRHXQAPNKvHt2U2KhSTcRRencTsn65O1C+
YZJtUR3uy9j4bZ2Ou1IfTKIYl8V9EQoORnglDeFqpzWbI0ajc5rXCISBRcscc+skbl1Lo/Y0xLs1
52BiQEvW8xx1gedvcMRQTUtJB64gCrVQ0rJKGWjbmwsJB/hd+L5nHVDrFI1avCVuzXxSxOdbasAp
oS1tepEYtZPp9k9TD/YONFmqTW80aDU7+xDWkOVVJMMGWAWz//fV568sjAZbBSDatd6oLiz2/RyA
VYTJU8eaSMHUVbW/LI9jfQN1uU7zZX+a/fypr9cykUScAX5x5Ge7EacNwbQLuyH0kRc+UhfbHbEZ
N1rMmEp65Vys/qfZYxFHWe4Rq88647Ef0zryxGetAlqlFPwTte+51PI/luwGm5GS4ERuH9T6iSYE
VjpJ+aS66J8yW6BKDHuvShWfzSnsFk3jZitZmG36hT7EAs+wrQTEjXYZQYb4GsaEODFo3acAxksA
w2DKte925sktdVKo1JP7XSyvfxJHXs6QAKf5Q2aFXj9ivcCJ7QiVgQ9KfamykJPrSuwh6YTR4yff
AgMZZC7qMXpCBLM4AIPrVP4jItGmRXAXOTQnBwThwyA9yRhazHynRFk4dUF3xZkpAXwA4ftEoMTQ
0EAG1muXIlJh/DsaXfyjC4GmlSzdxoYjt2w6Bwj1K6s6DgKHMjH5SRJ6AQxeOtFwseTAsdMemL0s
Z2cSojs0m9V3KQpOzXHVJwTUnoE00rrxjZ2iXuUjpyJbSU4OqkUs3ltfa7k3s5kWJWzqGIGIyrQv
doiTCEe4PzlYCuv0/VKC2HG+OoBH04hnh0BMOqRzhzjHflhTZvzQgSpZItEOnmBaTmFzUJKiWP3i
Vu4gULIh+77Ykh73pV5D1JFMhZhVophIXanAujNhguzessPLM4gz2YKQ0vCT3Zqwb7Bj0/jztSwZ
a91ISk0LYOzNAi3WnDsGWIF9qxvzegGhKDn1NRWuPdC4jUdwrltl2IHxH/2Q/635j3vqBXCkFARq
nuyHXm9F7ZQh2Q75TTr5qoVfKH66WtpHssAeiOFaavagXY41zdK7kUPxDe5r7mC9M4QVbhM4hHnX
HO6lt8bQMpILbrwNowXi5slh0AhvC58BpV6AwjAURJz/Ixxc8HoKDm0/DmLpxJH4PizCf4rbrZBc
k/Ce7gO4MUZFjDnjFI85TvKzCOTuydmo1yBMNHVh5pFDL91ZeWwAbdIptVQgVfstHVL0pfX4CvR7
Tn2DzOCpc8kasos6TtsZrM3Lm3CJpg3bppifUoG0X3bTecttROjlIU7dv61qpRio98b1bVF4uoJD
wYfFsaIrIvrRjCe+EMk4C9kvBSBE4fXw/ek4YNj+A2XcKmRrx0gOcCSUExt8CWm/Bec+vGq/qMvx
pleZbjaCv0CbTbBgrVc9wrc24iqjTCf7dCNNqwJobGYXjD2BqQQi80i9rXVR1ak307EM31OnNuoP
IiLak4nh1WhhLJgwXKvsMa6Zfj0oQL5QVuMGVW0i9MROlItRYMSEnEgXikAEuAzQPWGMjjyBZ10/
O/dri+6fUikSm+gSPY9JvhF9ovUNJ7HK79XR3L53H2FtHOCrljvckITzU6RN84/ghohspe5WvhVL
ESbEvHRq9F8Sx3FAZqueudS7WlFu196OSjo5bsVFQYFHfs8uyVgrsiJEw6OF2NzdEpgrbOQBERMa
Zg9VCqVYy1LJBZQg3LUtGpefW/NIPUC0CiRiPZhQbFQvW0Gh6ZFs0GmXA6GUd3fPpNDSYAhMR1JO
Qx/EGaLKCdBEPO5XZIuVbG85nLVhElAoMSt0n5NCxGt1R+HnC1c96dLeQGiqyuxIqWDqLiXsfoO5
bif9Ao8mOm/vSwPFav0VfTaRUq4F+bB994ed7npdprCgyC2ZmSNoKA0TuZ8EspseGuUZy090sAzd
Ev7zP84C0fRpJP2ObhqD3Sg5AvviouR9Z0KDVS25sZ7wVblTrlWKzp6G41yR7jpZw3Ru8Px3icpy
kcf/xk4X+PFgHc+OOCeXH7L1TKy4QnERKhuchcFXejP2SsHHDqZBtGWKLlJb9EhKdGakQbTIaS53
1GnOrcfcBkheR/4IfB0J4Y+ExFfYoWu3vk1yAFexfWZ4il1/M7dtpHVjypIEEFfiOFKDkrAQ2DOz
1gvnYpb596ZcsmdXEdR6ZM6ZaiuvhF716OjZ/On83HTAhiwEpQwX/hl4gWCGJgsJwbKqCzFgM7dE
vLb08nnjUTPpjpuksyVLeJY8cKt30NrNlhHcNcDoqHl3ScRKwN0JdH3u9WZ4d2vYlLVtlJlQR46S
mSFAmSIxtNSH4x7Z/dI32qnkkHv/yQfa2s/WV75IH8RCOjdOlH/U1C9w4NsHgUZ80abrE/JpShsB
Efi5qqWtANpAe6H8rRJW78hFNa7hZR8DDzKeCWdXK+dmS2pTR4Uhy6tv+9jb7VNrgaf4oU9x8GZY
xhmm7839DltU6efbTaKxC+0Gay3RzSZwA3PUlrq5peBVHfo3uuv3lFLIeZFIZXir82nvkWoekI2m
IVBhvbr33wmfDHkpTDsoZmPYMWLvcGJQ33XFZrFWo52/nsm8kT/uTOwQOkK3zUugXOuQOXSFJyLS
cB9a8YiSGdRDlBWoHSd/2qMc13g9EkxTvY3vbfkaqhVGFUkGiTHxxfmNgiCimWLRePgE7B+7pBkt
EaASc+AScmRMivOdIizN55G9Aef02J9TYktvuPer1h2+hNsB9WNtBVYVcmv7uaJuyp6hSmehBsDb
zBMjnLORZoDJYOd2/B7j016clO+FLl/o1LGz6JGiubv1cG+QIsVDDC0YnqenHvioZ4F1/sMp0uUb
ijitzl+SL4HA2ckbe/H5RpsOz8CkvUy8TZvrOEwCwBEIByihPXiwmcMCR/nPSQZJwkAROahOfAzR
HQrOTLBKWjtKD3I/Wiy3DyIDQ0C/8/hvZbu+oaTSNoBexzYvruSDflOPt3EYmrNZ57AtsYZD1VlV
ks1WJIA+D03cwj2pqrYagAEDZpogdwVQT42JstwbaZY0eIaWrYOXrm97Q6kQIdg3OD7H5HLOOqBL
uY3+Gw9fei3F/YQ6j3FkDH3PtHupv4RnAQ6CKnHBu/T5EsOmlDgBPqHXzrqFegOob9Fok9SO7/G3
kprSYoiI7/8uQGyU1n77+Qi2bb1IKWge4PO04F3SC3hGP2yCA/lRYoTY5l/jwLyK+Ga0DloivMnb
0i+z/4OO8bfR+uM4sD81pc4xyr02ApLQdLLwU/HS2+wiP2kc+o4EEQ+Wb+x8/kS6EaovQ14SIoBq
xPZ08um3o58LQPArkCCGMRTtelxCpS1VYLcy2NguzVQehE/rEgpbyLnP4ghyUPOw+N8AjZ/k2S3z
UUby/8ke/4KbJZiQMVLlZC2O1JcM/Hg/muiatS/sCCdcGFYFfK7Zyk4cOnENB268udcg7Zb5jFMh
fsm66FKPtEGY5YMH+Zby5sowUEmz3KONJQjASpglVk1XA+HxwdYjh0uR9WATP2dRDCIDjCPFwRAm
lj5bu1EawEH+sYrEJQ0EI8lTD4Ea2aX7nOc+GSRLAyGqDYlpaA92pgje4ftBbHrNGaFcp5y079J4
QcJIjt4gJqqNeXnEqq+M7gXQE0+VM+xnIGFLvWfTzMbbuADxqioawLQoa5bbu9unxMu1WfCb3Ehb
Aps5gE56q9Y92K5bBJ+UbeCMWMeBA9eVsBsNoxXd3fAQVs+LeXfHxKbPAxuyKjyqngiS0SVfoXt6
QC4DMpHFBUbgVCIyAfgpNztA9FqVFrkL0T+HHgvjgFvb4DFNGoZztsaVJMr6MSr8KymNpNuzkOJO
SnCjpbX2WSTz4GKtcCff8Xv7clsyiRpZKRBgEuYLnPRc0mo/5oisl39MUb8UoLwSPIcl4IxHJtuf
brhDG3z76O+qh9fvbSI0gfwMkWSdi2arkRjVSsGiR1bAkR4equbQhFnwmXFppC0+PEn5Gnzszfs8
3gJ4VEC4q+I73T962KdtK9F7FaQHPZU6cbVXr/Og9HGChwNlZpJcSlEzwbmKEFi5n4WJ/Q21OYMC
C9km1x8+S01lZpssfqosu58py4MFq5HGslIv1DRyDvLuniFM6VcywpaXdpO7Eh2Ly7Z5cc9cArLE
w6zVH76UxswbWl3iu0i4azJAc3wexCerPix6arGwNmbsUd/O09HXAfeOcPhmq7O2mTntliRZK5p0
ino8GJBZCwhydZ2At2ss013Wy2UjhmommWW066rW8b2o2zlZS3CZuyB+yNaJIYbDk1qLHPq/7std
/c0paVsJ1jC5TC6zUJ2HWlLkE01aczUbnlhHt2MTA2lyonMUapgQhhzSW+MNZoMpl0yrqevKdAyO
vtLqvizqNviIYm93hYhRAe/0MlpYTNJ0X+y9ReAIrCENAWI8soo6FNz1VDyeRbvHJlOTCSmuysA1
Y4pxzyIqXMspgngxhWp1cDvZZI+25Vn6b1NnLdx3wzF2F4Xh2U8Hsi1ehyDDQYD3zNgNyavbrfYM
v+3N5S6WRcWXwLMladki2CMC1OprGGjL+cUOpqsCK5GoEiuAZoo1reQgdNnJs3J2KIuMTnfLCerO
ZHlizV89SWgk84BcVQb+WrUrTg7tF53EhJE4qulqi7pMoCAllj+NjjTiXvqjs6fMl7ahMFwyA5Kl
7OXidNplJxopw+SckIYIO4FGl9LGIwb2Rb/GA79cKBLErccv/g2sn0/rOP8EnrB4y3vXxYkD+zBN
oDnZCmMM1RItPsSO33WYHnIHq+UYCaT5htQup91ObtXs7sraTZlJwn/K7nfyVUPikFcLZ2m+73Df
aaQK/bqV4uwTgoFrZb72N6PrJct2PSKVayIOFMHiGyesaJuCyGUxefQZUp5xQ26fth7TOyLzqpMl
0d7gvUyB/zcZUbJSeM82pGQLfbG3aweqQ8Dsk+Wt7cJ6H3aex0uGE3ffYM2YuFoq69YqLDHeBn9F
+pIE3BTVb16FS2JZQkCLCq4gqJPv5p039QVIas2DEz6jTQC51JRTmMolHPpwnO5F4WzAQUuq2P23
kaHI8oApBLZ++nNr6EjetnxUjUyLZP4Joyol5nLAPon6G3ooPArrxK4tZa+Fs2N+YtzEOrXz9Kl/
xH2R1Rh8B4NYNl8X06vyLmV+t0AkzitnQxz4kP5yb8bT4LuiH6SuhyY5Kz07HPdX4gThsVyQa2d5
DnZndydgLRHJvXHo7c736OIoGzZzoP0teCSzNkfl+j37/ZPprSHAuSLZ7RxAk9OSCCo+pBftGs83
3ztpjM2tVDjEw/2aQDLmptwuz1vJy7DvTxAHka/yNuKmy1KV4sdcZuppC9ZZsk7IFWdWwqgcFgoP
zrBCeJEMIGPgJlRKC/Oz2a9fKvxKaMygqpEhX8+sVQkBtTZuEoFLUoTdVup6KtD9JY8T1r6VYrcc
L36NRGvor6vCjUl9xyo4S9uj9e4jaNbpSWIRCVuLeOnz+ogtcIdcgr5e2riyRQaK9V6opae/lA9R
z74LHopHrwVWZkSoAs9JYnde1GG11TgdlEmdZKhJrJKSgGO0GdVb+aiKpz4+WBfrVZGOeBLgxQH6
zXR8MfDUSL7Qdr8at5KIeOzY/V0k0b4hrnejPlWc0PHTIePqcFGoIDlVxHTv7gM3nz+ymiQ9tkXQ
7IAI6xsO67sa81NSHe8S382t94uXQG+Z6mFq6GD0xcp+s4JiOO2X9qwhV/4JdtEcjPNj8FyHx17t
BSgYnrp9HcHa1tMxOpcjxt8LoVRIxPPS6iN3dY3MsIlVBvxeO6Tvrrr4MNRMr/uWg1LDWwrA+NA8
uCD14DQvFvhrDgXQ784U6Iv/Sp1CQFaNnxqxIZpw1rr/LiOV5d6TSZGl00TV7S6C3BKDflsznSEm
5fXneJg2Fj/XI0XGwTKpSRjnDqdLP7cZFz5EwpHG4cj7Ei+Fsp7lyZKgfbb/5N9Oy/iBEuWj0rZL
Eg48i/fCvLNA32xAN9yKyMXWGROQydM9Wy27AEqo9WmwRpN2dvBHT1uFFqxX/OsbCpAUauOLre+F
uEMhbmfjeti+kQVu7tTOyzW03Is6+QAIaMkZ9PuDAiHVMp9g2EQDZSGYSnSwLrd3JgmSvZsdDGek
gdIFOEV6riFd0eXnkUOgl/HSdQVEru5+0H1RxtSwe1Pbd2zCMh4QR3uwCFfukRV+wcymph6RjQfr
YxYfjurm2EJBjU0a90ShCbMf1I/UcZ/Lw9tZKvPrDA7gCUHjk2lmqb+rYXVAbuu4CvcvyiHtfgX0
SK1Z0A+4cSLUO1JIBwyIUp0EPwtSakrOACz0nIYXGBZWd983Hn5KQ0wCs3ZyX2xq4Mvye6MMFrhz
XcWIqCjW8mFzDFk2MaGmRVZXpeDhPwe6OkRdbhGbLmKGU1DlVla4TgJisKzQVKehaeA65atjI8P0
rmTOgYuX5fvMrEUC4/tvLDfwkO3nLFjPuQ3QTTkrctH5dyHUCQbI4bRKzm1fCan7fkNpVOwcACU6
xER1Giv6hzqrRRbb2hUIRoNyKy6ilKlDgykJkj9lO+QjlijIzRm6FAnm9t1hN92UOUyVEJ5pULXb
9hF93Xch5pAgbXG5T7mFV+PBqwYJaMRJtfUn5/bnJewpX6effP+xTrTP1i//vJN8fDeWg/gljBXT
5WkLnY03OJgDRzdw+P30RDsgdYZ3ySyggX3qoiEunfPQ5eRb1BegH2WSI6c99mM+u/eMs6I6QmDr
TS/DVKWvYDlrFm7Tz5ZVon3PHn3ZUM0bca8tUTbjtONj80YwTUqDJDVJG5Ihrlwqc5V2vKzYC5pT
HQa0DKauz4fOX0NOKUoSW58pVFZergestwWtDzDP1gRCfRCp0ToESCX9od26jKLm2VTbZlM4UBBl
ODZuKLKTPpz+7Tp2nix37AQBUlAKLxuSHm8e6H8wUFq+m1+tLQDKMSMw/pxuQM8xnOaOo9h5m6cF
G17C2HF+rzv5xwb+eR+86fieTGA6a6GR2MuxuJq29c8+xR4PEJfx3pCZcc3WKlJj/l4ourFetpa3
l06AXSeR6X9ESElu2hiXomQ3xpVGoOiZktOXbRtDH/USIfgHreqTZeKGCoVtCd02sNKTMdDDeZ4Y
H9xXTvtqLzikj8HDC4SNbtZZ039nfkxqKOzPU0AuzWcBndUVczcG/rk+2GIZx+PWfwf+Ei/ewI7V
NH8kS55iZa6mGur4fNO02z2YP7yLOiI4O83FInMgX7DfJk1h3sbNENTzNgB6Y26O/XzaMOc3nK1C
veTYyl9k5jfKcPIfhFFpOuumJhgLpiGL1vdYQO/m2i7tfxl0QqRqVug9dyXaWz+uB6PGMLUgKU/0
DdxIW9fp9X+YWWFNnfnGJyoPdUtMPATlU16fu0QaI6Tp8qlqXVAr6N5TRC9vevIEx3X/KsNTzXCI
OEK2iiVqFHEwvHWwqvUIdbhbnmm9oPlu2y7LtVq5GVo7Ayhh2BXuBr6UGU4pA72s9AVoD0s7+LGP
bVrgOgK3dx5TfHc6oKhzFS5XfFwmIFkz6AxrAiBWhHLjehmOeo/Y5L9MQ3qfVY6ySV8rmUOnaKOK
nxpvRz2dsxC82ghGWUUDx3ngzxJ72ajzrM4zvgRYU8HbJ46JwnJspV7EDyXV7nA8C0YKDncTZxu8
NLAVFUpHV2poXC3r+qAdscVAvO49NvCRbO5niJNPViU4z8C6GfuE6Ak3e8DxZQcwO4tS6d8K5v6s
eDazE/9p6U3x6zA7g1hpGIqlpZHkMbZU8vWH17wKPRQKAF0Xk0sCSpWy5DqTbOUi6uVSE2uavlOP
fHB5+leJse3+rp0BWGrb/PP23erfKTCVmQAekd5Mq/07jzu5wUtYb0scrajseFCuhFhsgvfftLYG
NuRdx9cy66U6xlaVHlIRCWNHusbYrsu80/+Y8o3gTuKaMPAVYSjPmAp2exSpmXaBYnQjhQ1cEvvY
0trm99pbaUrL4fFHJeWWTkQpos249lCZCYCEf72bpmyE+I3gdi+Xgyh2kGMWghs/d/efQydL37ln
SC494rQfJt2jG79qBU8LrQ9T3JHtnP+6GdKaeIbZtxOBl+9AgW6XhtIb3efujeGSlo/WultY9gew
XqbnNt0w885RNkT+3siPqv8MGlbNhibq8awo0zhQyJSYENtwpX0GPxjIVv50vuGaJcsPyFKWZnLR
pjMP/no6gwAZw+WlXCZ81ugRaLL19Jla5h6Ixx+wQkKlFAIBp6epIHSNl/C0ptUQOmwl0EBUg0ID
s3sTYDJqf8gxaaeu4EGVF8zvSonS2a/cOGJasCZwMBGxVuA7lnk6v5el8KlakMXrgxs0XGkZpVU9
uTPxGNJlysq5m3eXqbdbKeBFA7lRgDFVSfeBp98GoP76YPbMjgPSq875oHFP4TiWVRfy/BlDX7jB
cq9T7CHI17h/FdaZ4JvJ130xebE5Xh89DJza6hB/ltIznRZLC+/4MP6wXVK7vDxNJ9l3VSuQpDFl
L37hjq6G+Zy5IhpVmb0+a9wZGem8GHwxcaAori5vjCvx8v+FBpItMCCdJ9j48HVZUUvuwujlsUAx
az35ASilll+tI+2jjs+Z4Y9AvyrTC72dMHjL43CHTBOCRtKchxgc7FR2ReCj5bpeX17wmOvc2f5r
31xUEVRvPWD3u+HqKPBzLOKiKzXMCvOzjYX21QqbrCAEoOulVVA94I4PCnKTuXK05M0sF4DcFQci
we03/WJjKutONFzkq58O/lmHdQOixLeblxgpTnI08sU9PnyIdea6u5gDSleJWoP92bx0CWUKaLOa
hXKead0c/Jm63+9inX16adHChRQ3wRHFrKCRG7bV46ly9ZrWUeVoQ1Wxf2x0ghkAgfsLDVV5LEb9
U3MXVuYWRnqHdgG5FvSHa4PtkL1owJz/GJ8Ixrxv0onyHgo6vf7o5CadY8dvjviY5qMrkrwoJ2fv
Y93mnL3Gtw0egMJ1F7mpiAdIpdOupGIRAX5ZGKbs8OPUb6baIDbQXZ9eMaPJj1U9391oBn3A1vMp
PPSn39pLD7pn6cR/qrWvBNCFtRemxwCYHVOMO9UroOo+ztJOPDC6j2Vi5RZP3wB7FS9E8kzyhJJG
X0u/7woXn2DqQXIIRu3p157nH/YiQ1hwgK4NRlTlF5TGJLjI9ZqjGiaynHpt8L06sKgrCQr4infZ
RvKohXf09pMAQV2XNFGGqIvPDH37BSIe/io/V80bNen3jPbO9AZj+5duhpoMm8bpVj/fpCXifnlv
tRiKCAIAcH2KHgbB7+gh+hIGwGA+2hUjdCp2dV8yjywa5k7VC7ApEEocVI3v4Vwj2yu+wzKbrbMS
iEl1sIe+3h0NqSjU/zOtQNpogTTRUHVRmp72SbKFed1be9pc4AGiJWpMLCpQMdkREkJ7dgxsMFdD
kVZCJTbMSGQAOetYtyVb4txdpvxSvvoLyq3ooLvc+QRAc0CL0SaBhlIX7mSj6NFWy0cdne509HFv
liLyJoos26S+k3vCSj0u2rdvAS1yv84Cb88ss2FEsmPfNZYwf+y3gQX9q3xBIKPXktxQ5z8PqEI/
nN8kJTu/fP3rcsz+uaHESTLcTkDi44GoSWJOHLt6/wHUHpRooazPHP6qf6UHe71d1Nif1NDsMArJ
roASCYFMoXmRiVVFFr+bPKCco2sAPyzhrENDYrIigtuBYQl2mI4/deUnWQG3qBr3kORRE6VYJ0xU
fY709+7yXLKFOW6ZGK4KLcHA5KIjZigfVLkYW7J5f1DkKI3J7gMmrkwYN+QO09KBB4wBr4/AkpMU
u04RtNSeykWcVlI6dRDTKwsDorugitVAvvpvqhJ1hk0hGIA7XK4afZjF5sWrj+upRIeHwHCJpc7b
KYpm44f+47FcI2zGsvLtQrE2GENh0qTiKkULBmZuGPiXKPXFUHYnNCzZog1PANxWdqO/55pXk4Zd
eHzk2r2L+rqF/XBtiubiZZMCFvdfLvff1Bycpb8+jg0tiQQJpCQ7v9/v6URWzRmzLh9Yjl2bVXbF
moU7zsxLD+9EVmtJ4mEOVAjKsw2P8nWuMkxzvuY2xfo7DEWTu1KPj7EYtYKAJmm+eOtm7cDNrFsc
JD1L9MOGb/HU1f6Lk04Uqw/tLOPKUotXtsQlwoaVPuQixuwXmt5uHfD5KGYoSAN9GNHT1oemDttX
SoXOI3HOw5j9aHRiPtoNZaHkzkcFZ30ySNwLL9ix+mkQYdS8nAD+obI59PYBsFFjhDD14R8lwNru
hOX0cMpLD4f3oj873rMAWFYHbHa8mIdA5i+EqMjwWj3sh0ngOlvHvkQCTwZL0bIT2H1ndU26lWZ/
1ux9/a2S7ChXjXGbtGMHbrrvzsuPqiIINlbAUWgxNZJJ/aIqGYCdEl26w+zJz/QzhHZ30IMPPTlv
kakzglBAD2KOIELvg7nO2iq9v/PDG78B9gM4rvtH3lcRonjQgJ+mpE3+OWaCKJZOG7gJ8pyY8xcE
Pp7wsYQxQOCI3F3HQTNMCjnpdeH9Q6mfCdfXf2NRZSAnInYrp4tG+oXhusWhPGbdzS1Aovnrc/xa
CUCdUgT5QSm6Apenk/rr3GASPgxR9qd7UDxmSR6JP4pkNM41uWtGFEDk6LxTz7sudXAguuPqhbkS
LALX2Wu/yJmRfHipf//hNsLmRE617Auz52tkBuAfcEeg+b3001WVbbga5nWJY6BwF/LwTXqYcDaQ
/hXIBHNomnQWkje5e24wkNOkkHRIuotbnVC81r41k4ah/TvuM4wg/63sDDI35cokI94SlcejA1tf
mwz0MPzg5TODN493zNCERGYksvaW7YRJI3eMav5fqUqf/3e4LmqOn1kKMBEDbVKp2lsCg0uqFlUF
w9FopzCggI8LDKZdrPJkWANy7qO9hzQynLhZ8DuYK5PWaO3B756tzPNMAVh8rLk2yZEMmLLq48M8
wSSu8KiNLZLOf76RZy2WgcdQ11jA6Ohi6QGnt+jXYOUtO/OCzHpngsdYiegydYES7tj5lM2g3osA
FHO7ROYydwJR25mFjbysMiZZ/zMn0mr9adyofryvJJ+koMDm5wRNQHJ7kYE462z473fbG7yYZhNS
8KFV9zq/LIRfHIj8emHhaokB/D6wbg7ri8613Zw6AA/SKQp/foxHxH2bZQd5dWRxY5Q53IKrlCa0
CIr/U3fS0IzSBPOgmICS/aXkY/hTSl+gQhlfl8fj/3nGjCSN+GfrRSVNEbnBa/NyGybeEvhmuYLD
PiApJhYCUXHrJ1gELCyKv+yo7DQafJ17JV4MEiKmZnv1ZDh8+kD6EsrkVKwgVhk/GB0T73B9EmIZ
bY6aAGvvycrW82F/yc410gufVyUG6JxsSa+lkYdgysrbgJuw6Nxy2tst8uDy35Y7C5lHMrNTzd3+
QNNsymNF0Fb57fwLp+w4mzD7nLxxOuaW+gW+FeCdOsbv9XVS5kHzqm56XswnuVs5HebyMJ9iJjZf
14+sKKff6FYVuaYUzc6DeNcoDFKWh9LnJiYrxAodG3fYPp298t5EEADf4B76Js2Y3Myq7+YKtROn
tdWOnB4I1B15uU2pAYER3G5VxyR09Z2++Czs2WboLdnHa8a/jT2kMupV2fbnEGW3bKdyFTXP0B2H
wJ63SQr4mB0jHM0Bnz0xAyNQO3LoOqGtMv2dBj91Uc6rIIbUBckC8grR1fkNq2RY9CHyZsTu1xTj
VoV1MlSRZZOaOQp6BfDfeyr4+r/6xuj7WpeU4ZrarPMCdnlKARcbVRrupz8QVzfFo1enMVkfKdAm
TQ3txBywMQlqYWh9uXmtZIfLW8hSyDKiSViFkfgQosswQGaE6UnrHV7WuKgio+Ju7aRTmeCazo/P
vEPRlbzyde6IxbYNWAcqHSYsZN+jREU5zlOBAT6Q4O48iop8ma1fZjDC7vnKLyDt0tkhq2uhA8UL
dvjPpYxdAusPsOBbz7DooLSDMDXfbnwrI9J4P+aRaPds4WN+oM+jGVdfHBS2VKFXxryQibd50HWf
5GOO9wQRDvo5Ag5g0Xsfiz3drsKh5Q2r0A8n1tVgOWBb5mDm03dWGa8h5jTw/J7PTAj4rDSp/aQq
QaZvURdoHeBahQP/rLmqwcy296O8xzhB0OltJC88p06+O4spzP/RmX3dgFPItyM9GPpZdu0jGTNt
QhVq+GhzZ5mTKeV8z2gyURcKLzVWjPA+rseIFdMLxDhEh1D/c9GWVahxMukpbGiPwp3P0pkPL77X
KxG0Ev68qb51Wl4RWZuR127EPIRGFvSHaxYuX166e3QVFs3FRjZkIzwtUdqZee2nHCUFRnvaoYyv
0BPXpJxwZN1mwEldl9B3IW4N9XXGKL93moNEcTQBZ6T9kFzdLr+7WUXfY+3z7riutPAtM4Z/wnAp
ZGk0yn6v3ALCNORHyBgYUpasyQLEAWXXkVBesIyqW8Cssp7rLfOQmxPpX17IACg8Oc1EM9JSzR4B
rVNrSnkadzvsWH/QC5Fo1H3MtLd7/fpGPJnZGy4rEPMx7rSbmNRpL120HYAbWgSYLxActN+PEJ5d
0QLSwIgXgKN7vKY/J8s7ZpGc/vhn27D3SiUuNRIg372d6lkrpkj7ProF7zZGGI5hPJyZ21r3YSud
1XaGKgiE9RRfNKbneKbpYlQ2kDik4oGTHixPzhHQMRMR1LSgmNzWI63F8nGCzNZiLNpk/lzZrxLn
zNFnCTAxQV93E2ZYUNdoyTXvnP1eL+oih/m7KZCL+tyzaJK5eZc3YBn3vlhnG2n5B+Q+YYCBwFDU
C/axGP2MnpUEtb6CXU5fbXNq95Mf1LbcTJA8aOoTaH36miad0MwOWT/LLBy0ZOZBUwP8wsqd5yDL
G/1T/0NTIuIjqtB7GN8rH3h3nBluS/Dbp2s71EFRMXrLuFV4mJq3hDWSQBRiZQPGRSyGVpychdMg
vTvEsoh1GORjhl6F2jxrZPYT5QUjwn/PYMpJPMCYAMTV57mPkKtzTUBia0kHIZgNobasas4oM6tI
7f98y8HwFrlFdOh782an91adky+5DpWFDDv0r2KaH/MfurlUqiK5J8QkEoCLteTIK+xrSNwIxIwV
wEr33nLesCqXzzGlUaRCGp2oVWK8Q8Z+FiXmZcGsAnd0Vp9jLbbmCJRqKroZZ3HDi3rTMG1PVVQ1
LB91FgAfgz/zNomFDYzuhdZA7mdLOwG6JN26ZCp9gQwLkODtzqTByV7H1iEeZ+F/6Yd1XX8RAAFa
rc0jjCox/2/a7eO20XKdXI63PjihdTYHVDmrOJRDUwtmtPxZpgiq8bAHf/IF5nwKC/1RmcqFneN+
BRtV+X6D2SGtr0QSUYjCwrRLRC2XZIy1DzpLAD0z3DZQ2zinDNhUVLEkjLLeOhiRIUroVhBYt8J3
lgxmN2CyxsD5cdcbkaB0JSYWBvvwTO3fsq4g+83zng54Al0h+xFF7D0Ku3SQFH+XVCNX99hhsDzz
eLh4n1HcmSyWS40aAyr7C4+SGV6rEMDrZQgVSkQ76M3pRqC57bdICGKgXg4yIPtZv9iQ4jxALL5a
kcWKRnmjAYJtNMEvnPuCh0aIGqQnWEgV8U019BP6OE/NIKk6vEoUg9vtxA9Dq/Yg8Br72sd8tlRu
UNukmhUihDvgUv+AkSpBHyLKRaRRsleJpRZoZ7UPt7a7YFJi4ybmDxYLvtS6anDRgshkZ8be8M9C
kvl0qcJGf0OkNL9wq/yR/4uKhIpc4E9FV8cNgpDjMEyj5R1ZNKDxXFF+tLIxCBf3JTaIWwVhmBF+
rnL3ALNouDKTOV5r47DxnoeAJjoneGn4hQK1ZkKNM9QLxt7FU3GrH9Pw2g33t62JRiMncZWXp2/W
/4guDUz+Ee+uQ0QgKRyG6+P7jQA/qcH4BsEc40uEDTH00TA+q77Z2zb+U7CK1gmdFI+5Gs9glu1U
4zNzrtaxwQx73wNFzs7fx0eI/8zfrKpR4IkhYUoYxVIX+G8hJc8cxFW7uqXHADBaO9qw14C1HNcl
X2qZ3O3OqVNlSLvFRy1faiCyJs0IS43aFCE1nYg2NdZU7H7/H7vJcCHPdNzsmqGzmo/XaFwYY8OQ
+qvzu/or9IznbI0ZpZMR3S/EQRgRfPZEGVtL6aX8l4UESaqPWNdaeAqvdw4SEZQ/wrzY/anWAWz8
xbAmVRAgafjwoPFLSLVrd0qvZHA/l4Xz5Ny+dV/7eCe9kg7UfDTgDf2CzodQrp+jIW2QGpE3e7F0
v//6s46LAbAkslazuB19vsuqaNqllvHTa1TKVUsdd3G206l97If7lpgVcCHu5o8xEcZcmeCceo35
3TFjj884yPi1Sisi8eZthduQtkzQwE9csrg/AUHVPlmhN3S2G7rFfRTCbTt0orosh86ZZokSsGvh
3Xaunohi3/oySVC4Uj9OzDQWBGSUEzSt1VKkc/0wkcuqvfPS7CZCH6IZiZrTZboCWCeRam5s5SMw
fx78bPP/aNI7VVOy3UzYMZN2d9iMWWJlx5Eli5b19B+to0rgWBsoYV9SoXIBMySWXgDDNr8ebsAC
mSAeTCesHCv36TED+qV2gZ7c1d9kJXp4WlQSrj+4PPOygrb9apC9Xtbgf4PclsqMnDuRgVg4ByR2
n3149q3g3tuCaJuJTjkP8NzQsE63F7sn7vgf6gYQ3rmuuOLYrznb+eofucwkFCTwENobFjHvm0W+
dU8KikUR4xka1mCSe7Wb/ugKEEStfeOTF4XAAT7b+mD3mrDE1JvUpPihKw85n4XyPITJ0n/vf44m
c8XkF9tgG9jQQLG/uF1cych1l9+Sio+7yOoaq51xTPFZoHmDAOaTmoekzu7kBNCrGdQCfSH5/mqc
stH4eLJeQdGaVH+MkSl+u7OhLR4YCowcQTa8EuUTEiwvYHmOPMYWgkntFy+ojydExEMq6nsUkp6h
ezq5pDPYio0SZ+yPHYTfQJC6PdaBrR23huTAx5j71WTFxsMggQtSupCZdsx8TZ6qw+aRZLH+mpF9
GIA92cCizS6zElRQnTJTzmNjMjGkaZIryC78GdvM5DAjbi0GqVvPA28o8p6i9rneKrA/hapac4xo
6jdhtu98ZLx3dDktDteSLpw+UNrcJarioacJamkUhwj6aJ9+06kifo7Uivm4OBw7Px0nDj3HVGpv
XIzHe5aFnYfZTwV/o3Zp9g3lRlb8BvCb7qpA27klYOkBtYAixnRNezJwGut3F4bAmgQFbPYveJO8
NqHE1uzYE6nP84Aq1Ay4/41x7F4DMLZqOUyHBoEmgXvCLXJilCxND3QVgX3jQhxAnx3PjiBqBV08
F10UHcNct1oBFCqkkyN8ydDuL1k9bUtdWkSzQ9G0InlZkTRALKTjUtpL2dTR+pYxFHZTIeBE/UEz
I8EiP+KI+FGDk0/pUHKWK6eDIkPKwhg1ov+3EZhrKoB8nqVs9eeRcoJnWvRJv+fSDvQ3gLjDksOw
nqhBANcEADlIt/R7Ea4TSwOxBCwTh4mljd2BC2V1jEH5GuF/LZHn6tJw3N3dEpXBE3XnKoDhh62O
etZD+HH8Q/b6MVdGyzvGNonYaWvOYcgs2ErfHfr2rWwlzeup1NAH3+3c10NR2hTsgYKgyctiXov7
WL4R6WydHAtBIFYzaq0vTVLtC+dkhDQ+s9/Fgk6FyjJmwHs0EAOf0S/Iia1g6bCncYe0YbWqGJCg
S1pHmhVy6QzG6Pv4w4et5mkFrfG5pY2PwEUQ9Y01MiG0H2n0fOy/UP8QignLfG41DAvPo9vCDeYH
1d9pRAdp4dkglwcV+p1KLOaoBla7tWvAgr4sN+5s+i4ztuATu6gB43mVFmfdNE6CrxguAHqFbk/q
BXKffZghY5pnxLqSOAacJb7xp3vnD9UDQk1bulzUKa1uHsPVldRZjvQ6rCeY67TaLAmMRWWF1v71
RlMdS/GpAM7RIsHUCvsKFNj+KJ1ViCvqessBh9jxsXcgf9s3FYTV6GZaX/P0R39OBh0CYbS89+IO
YY2t+zZYhr/z942NexMSpuXBwSfNEtX+PqUWAVEaBZMtdbXJtmb1yusRHyP04mJXIu9ZJbiFTsUo
bMnFNHCDcMZyMrMGS5Mvgt9VmeWifjohFxRuC2N5NsU6Lsrm/D1Q2wZHyFKFzAjecNwW8NifuEhB
zLI9gxFI5JuJD9iqQ1GrZBJ25zSf2Zb39GKZze47oPmB8TOZqnkvEe9VYu14XadsTaNs81A5VQAm
keU9toucy1JNAa3ekr1dzqt7xwL9UOfb/mwlAie8O52GAMiRyUY4u0zylKO9RmfpcLXBw6/fKfw0
ODRDbVb8dpGs4Ef/lRiTwr49A0PCvV2uLxjN12Jp+36jjzY6sr14gYXaftnwHxiw4yJQqmoZ30bE
GdSDxGEbLHW1azHRJnqkDAoIWh9U64Rr69Pzbiknl8r66BVyYYrVFgGw3BgSESC8vsYvkbbXWS1t
KgcqoVoN5S9e3cUvx5ZuKPPv12Cpu2tvCQ1XfpjY7PXDekegZkbUwMj0WnBsItaQDq0bDwXcJXzF
Rp78sqSdFS3TlgcA8ZjWA+YKnvNB3TgCM5/AmphZfhtsZAbCZ0dur9TghuZ5DAI9nKNFjO0N+01W
mOfM+nglUoC0VSPme3yN5f+YwUvd6OsCnonRLD2tnXIYaCS6++eCr/ajq2dhZW8K3lEG9x6/olpB
J/t4GeEfA2BkUz5pCh2wv+pQ98+VbB2o8Vew8GBu1ycKcVloQ3Iz0rPqNLUUrPACsMjd9bljbxFg
hWQnTwt6gNegSry5thWjE9oFNeK9usaSWYkN3NNhyy+UqHUD6ndNbfiL7wFXAmTXUVq3aA7xn4r5
NYDSh1DrjxJdJFEh3yocwE+r8qDbqkTHUmyFrPZPJ0PoUhrWD5RvNInaYptDOJsV+dJzbrKJQ5KB
LvqyLmaUhp3vUDFAxKiGdKcx4ZRadA19vvjdPW/ySQR+bmroM4Tfh2aQr1iNlPU87W3jik4Bdgj/
X4CmESh/0YRCkd0NVCal79U0/YXN5RAONHDl1Yx1Cfsi4vvQhQQyNjiX7brObAhTrem/X07oirgx
bUK3W7g5g6E58d1g44nihrlVuOxB0qRk3aWHJWudrMAUBZSmdDSELQMAenrW8Z88nbBoKuZGn21b
Tt1M03i8B0zcMgVEX1oubf5BNmwQ0i7Bb390k8gjqEOSgETy1VWbi22qjTD0P7BUPoikBbJVOcDw
ZjmlUVyxmD/NS44SPODfnTvRu0ltpUl4EofiWT6dLVJJ5uACVeH6n18TEVtWtPCdqA6J8zbIDYD/
2d1H8echMYRb2jdR7q0QyYP+9DXptkmt1HLFZCInkVft7+YB3Rg0gyB0MqgtVkJgGPGOgrYgN/qi
u0adViFiKQdK9Y/BpEdA0TKrO2oHz9rVZKsFpbSQq055jDFGXXX06lDb7BQztv/6kl9xZXxynO+A
cmojAm6ajQ7fCN/b7jW28Awfr1U3LbmwBTf2VM3mLSZuG8KfcVW9BLrfjyPo+Ov9HR5pajsoCnBY
yOuAt3d8Q+62QSCbp2vp3bQIoO2MCeRm4GackiS9iL5PNZBP8HThqugPhbYsEcvr20C830AtYJKD
Tr0j5+fGnDLTIBHfx+orMgMF/R739w513lOBbC8YV0KbVDTuCb2AkqaWTQF134k/CLTDDtiyexLQ
tvr0iRAN1QBmaq69DT/tDUDqpXfqfaxi1f3XryGG3JzljRPPcBxPs+pd6q7FkOqsrtGk7oDeA4yS
c1j3CMUtCaJYe6lRWJIT6o0JXJJ0G6IxaCyA4qnSuabjWciGzNOwLpUEXuM6L2tP2EvrGQIPamVV
xdmOYsFF1LeL6PiGAAjjYRlyD7xnrP+VYliTOhncFDSk1VKgRwzZb1hw3lWhNTIvsHz6Ld/ivEY0
WLJWCXe6a3JRfBgOHHZ+aFtwF/5LC99xC0Rrqgfz+/9vO2l8tsbtklCv8XAtPNhydX5zns8CGhMY
8Xs1ZE+Ne5YlHzmQjnPIXY5TdZ7bKbo2L7Kij6yDHl4V31TORK4Ai2xNIpwcfYmvJVcttCdGpakK
MxKp17zxlhRZARp0nFSIJ5pAlFoEwCPN+DRpxYUEaeNCdPvBv2B8xivgmMtFOBfmY8acE7WWyt8V
54Rd0PEfWaSygUwOg+//Qde9WguCb0fmvykeYFUcEcI3z6/WH3DbOju7/kVMSLXH5ygLSXWge5Ks
KHbsDckVGvS1gXmyZk3PQk4om+Mnb+wg9DQA6KXLsINWTUXkGMxXT2dkgAyNGeR4h9pK/HVa5WdI
+8jZZlPcsnAM78HLWohDrV7cEl47kanNlfn8diW+C3nF24SSRUmmYvVzu3t6NWgit5MRFyy/0gY+
H9diwz3R/4cxbtXyzWw8k1cKJe3YFcEL6EP7wC6A73m4jIqN2uFG0o0N4/s1/BKmwr/XEmghxL70
1JVDb1P5neUvoWLjr1WgBDrDmW07xTJHvPfgcNUiFt+jEj4aTQVVR6nD73yYyj+sT0pxhcdpP0Bq
NDFe/Ar1dmnO2WhWD1jpPE0vk/JDHZ7+A3qJytgjklcL9fCtRBOIVs6o+ubCvxpa7SWHFvprvbCL
+LSym3G6Mb25qD5hHqsRqBKBafdfULGmhoQLQfiEwztIar81v374K9wMfagQMvaqmjE6FdCUyahz
yxrFHErD6FDLNxpf4Bkq+Yo7LOcSAL+hrfGE/rWJV2l0MXIbDLASV68bOCE4A7/uX7Ebxtd/ayK0
U0A5VozSLNEfe6IZa3Xhj/h9Nl3Qds5ccIIbMZpiyo8WHchMK88sm0Kgsa+LXJmbFsfbpOh22pgR
/tJ59gTrgSeqzpyOWtQ+SMsgwZqOx8zZrc3XyymqPcjb+Yfe8I8qC/lEWZgPDScxtN1eh0BcCThk
lClQmdz+9BZjHjgO7g/mCDLjwpCZPuFsKpYJL38H9qSmYUcqhsnV3O+91BUVlarDz3aJN8EMrblF
bW+Xn5ewxtTw/1aH1NYOsXQOL8Urjt+Y55slG7oBH35tC0isUZxrYAdiaO68tAL4Ony7woCnA+pk
yZgnAuLFzTFxca4RZCm7U9ytyB9HnUb8IHbQpD3dTTglykL0cErfgyU6mOGPg5Plp5DanOUjuYFZ
IejHAfbsjizZASwnn5Cm+zbbn66CIKR3Cm+nIqSGcSaiDAozoJBIsCXrmzxj7UNcs9ZdFRzTLMsw
4LfJ0dF6ddBuihjCzp1cby8AsJQmJ/7uqWAqt9gQCS+1D2ko5h9fWG8wlYW8uXbjRAO+LgsGQK7/
BTjv8aNIx6w9i7uj87gcpxo7ZgBd6AiFEl4I8H7b/PqtRoE4MiaXR2t9CVMxfETTWpuQMOk0kku0
tvYyflVhs6Q94sl2iMVKZIR9W6oCloYY1xpJy4i8T1CQPcOIRQtIU/jIkRCnj7jLaWa7EF/bW8ff
j6aAeq/S5UaVk6T4ARQKz0c5cnF2hbDMjttbj5GQpWHICABUFf8txIILXV9wzp+cCENtKEz0sJE2
fU+DRrw0+mHjShQlvA/dLy2lzpq6b7+bl6mO84XKjvoQOkdWjoOHlv0GvgRJd4sGW8j5DrV9aHkp
BLmPcPiYT1f6qgMmR/kPnXXSohCcBkwpt0/wlwQjFXPqASYv+wKw5XthoCvaOpBSMIoueoPhqWbl
qPpkGC+I/3M5VjrZkKDmo4GA/POxkySHIgWU2vPAnIk+oONY9AA6Xx4QtV50l6l3cRa4ms+S3zvj
muwOEIcXjFCixFJb1PaIoYm+0cKmEwP+kep1GHC1qCRI6zR0YnsI7TkQpr1+hDcbXOZ/+E7XLQHj
og0cP84zGGLRfK2JzKdhFG0T2eUu2C2X3KkT9uzHlyC7ownrVWWvU3TUmiGbqS4PltoEmJSxoXUy
Pu6GbX2j+03fLixMKA1ZCwbPTXvsE+UWt0Of8Yi7YiRU2I3V9djR3lQRJVmbD0Eu30grC1w0U7zp
z1iSZ59TgX/lq/OFX/Ir5w2ykrtNI7nEQFs4F68x/cDZt0hjlmvVS0N9zVkweISqFBl9haU/iAOh
DyJjgIvZkEhKDRKPmYgOJbQWekh48HAzF7aJ8lRMYAfwtv3ki8VZ0lewKzZh1v76nR7e9kmimIOh
+LOPrl1+C8evv1GRMwfBC9dQR6PURT/EKEBfGGyPGkSt7s7Dnw88TLZrkBw2djLy/jsc/USXwZCz
iPeCHbndTPzEWWvoB+xGdyO8BjnRcEwqnnCOzdkwd3BSvBr7/elW460Ylmr+InNu3IAWYlGIdKP7
Dy9xmohAyADdWdLKJhkxaEGcbBwgb5KWLbAjnBzlTthXEA0OVY+9c/qTwTvV36GBQtxPNPSusB0N
y/mWSwfPuvh71GQK005Aslqie5cj9Qv++OpdtaBMRRCyvGBCtai3j13pmD2uSdja43rtmAh7Cvb9
0sjSlBr3IbaUaoXhWX9tZJQH78l9qDmmoOgMsh383xDOATVPE7RjBAGV55Nb8atydm7pPOkiwf+c
bX37z5cRMmXAOR+xaCavv+sBibPUXxbJboeLN4mo8/f8K9/aOSwinqAUZE+dmvmnHo5IhrY6M2V7
xp4/ZcwdeOCKKHpoPJKbaJsq1mvmhuMDxfCfy27XDWnBgXmEpoaOakrCEsHrzzLgAFN+Jwj6o3Z3
FHaOhmBtPYQG2uFssOkgFEkPi7oWapqiYkPpFKJ3iJvjVC0SQAxGr0l1Sk7Hd01V4fxYJunUs3I9
iuAdyWEM6azGSXawnlonHmBUajpF0pDYo4bBSUAmu6N0vSFitS+MDBUVg0b2rYimZb0WwLULP2GM
lINtJ0wGaOrQYpt5nMXI02MYSGfHe7Lai37qSsqcp2w8diUOg6mgK2e+dRSee3HK1/jsj6e/uKef
TFv6eOU0/QLwrR11KYPSh5FlwNgtCgG9m/YNMXPer9bscyEj8uG5MJKP26/1v8Fqb+qTViCfRSOU
0zZwjvv7pxy+0XNm+i4wzDFHPCT6AHJTPu6ezwN7QynHq7QIzkllYubhqoRZZbNCl2lWdDPDb9j3
3r9/k338b/gm5sICGvLm9FOdlKpvcWdDeonzORb9qaaYPxyA8zm2qEEp2veaWWCB9MloHc97DFeR
VZl3DC/pOUtzxCzlH3/MBJAg43sTejKBz6WUbU6xS3jJIPRnZM7dV1kPU/EYJfWsX/wjolmo3Yt9
mHFfqKvtM4jneQD1/iV2et9EoCx5c1lVuV9wAQiOAlPEnUcUOg8vHDW8hzkwfQn8iT8CBjtjj+Ob
4XmtqSqd4VQVen2PuB9lbpmhITTj09KqGbtahufa284yaCWPm2ix1dRzbY1aNN/3FDXthts5Hl9v
PBdlFO3snmwxLu2qafNkDEHAVfkQ10DG87WiAwZTjI0C74kchRy7WdzEsI4PJYrsQSEXFkm0TF46
majCRN7Gx1bD3ZhIOvcK20QrkqlqxUWZ/jbfuDa5FXY9RF/VeqL0B32GF8/dlXjUaR6uGD/XsklT
e3v0aT15TIf4eeYM2L3sn6YMyFt+CcbAKfzbYjh3TF2ScsjQKiU/okljqHgBhGetrFhlVMGCUHgb
+C2jyPnmaEufdjtoVG32ioTh9hc84xnT1/h+hgtQpbAOhs8idMfOdAf5dGWEx7wEETN4j27YL1hV
/GeChN352t1vL9/5YTtbU2IWSwB7P/FGdpzGeUyykhXpvTqDANwhYfzT6qicDDMqjAcpz8BFoedN
ATy2Uklh6b/YZrFbi+BnMUASqHySEiD8QhP0T9+E4zcJiWeg92XNVZq6pWDBXdCFtXCWIKnLGGvb
soVFBYxoePw+kM7uGD1nfDZxdsvC77bxzN6F6zzP1g5EVFweFZri4JLvKxy3KLIqTgmAHMyAN4fB
FtUzsKtpQfcsuRQqKYyUrGgr9hHv6IQ0RcvjILGX9N5fD2QOWm1GPAARmumU61gF4zui4qyaM6ig
OGUcbHJ1EpD6zk8NRirD8WwOHiNXMY/AuPAoxyBJrA4FqYFIcB1NPsYjx6lCRAGnXXHk46ABSHpG
xKVxEDooliLvCZSkdNtWUnEeO8UociEbo07OQ5JvGoeSuEc8Tgs+SNc7RFrSC575vA58QE/UaQuW
0ih8AWOwxnlsaBqJlZQg4iQm+Ts0telAKDZ9zQGe7pMjw7us1r3Nmu6RiPmYLn13hIGwzgVBSl3Z
3T62W1hQLhHXD9vxckeIvycQ/BWAlnr5H3gz/vJ21RMyB9cVQmrEqO0/RKka+Q/N4SnVEUG+rLHD
6ofk0UZDDjb1GWp3GdJKSlAhn1fOK3Q1d6cx3Fs8FbkJ7IICkkMAiDucL4pBukgF4dK3QSEKGmwV
+NG3sjTTZFQ+JFCQFTwHDT+hgDWkfIbLmcUwFsa5Vx298ZbkJHm/bmZF31gxpQp9PdJD9crY84bv
iv4KBc+DjNLfC/iGu7XoReqW733DuQIFYSqw2dEAnXM/UESfjO00qp1qILc9I7euUB7EndishL0H
bBT3bwPffPpHQcxwAaf+fyxR0n7zVhbtaw7+kng4llCniL1M4co095FMA1TVPO2XU+n6uosvKsn0
wZa804VVf0OqItsvZE7LSAfZ9jZ7cKwD/kGmLE8NTe/fT7lEHzwKxrUlgE9Wus9gvywJjC29nLlg
3bvLRWAgwrk8ztmnITvdtAN0T0ga4vneFYHM0GVQiHE/Hsv3exEntgSgXD9TcJ9bv+7FkeAhAzbK
vdcZ5Kg5Nk30pm0oCaB89vCgl4kpSUjqlyo90xRHFDO+FI4XTKQEKcy2i7VITPJT2ndWjhRkRAwU
8UFRLV+bBXDUKlRbbezcRtss8FfZhFuze2sPdNOMqW0F+iZtOmvDg5w0BbzBeQeLDWFz/BhUbJL9
H1bRrP8DftA/WZbU7fWGPzX7s6Q6mr/UOEyNbhBo1jhbNf18ztL+CZbP2W9sBHFb6Kbc+OzUr1H8
NW2qo7R0mQc8hQ3IF7A3OeA+YoHRq3uYpWTaotXZw8gKkFoAvRvsImS7L2F1kn8uGMzx1LPmrtKm
ZHUewH/P2ravWw5u2s6RYPorGUzeuC5AwzO7c2L58H4hSyoXygFFQ0WCLVdsuixjLsXzRsd2MyEp
tGJ6PLl308o1SL3OM1ZfS1HT+xQg49yelZNqsE5uK5NnoKAuFNr04UJJ8+0ORPVVMFoiGfjwsou6
DDAwQDOLpz9FlWDS3F6K4AKxN4rXoeVK4cHAfe1cNj1oH3ZwqHjgj2fb4adPXvnJUrUB8devd74C
MKpCB8P5dmy1YOwitkDH4wGnzBCNR+UE59loWqgZHkV1GXMiPNaq+NETJcbkqqaSOO98nX2E1gSj
vv9NhJrE92RzVLioWAnAbzo+WaVfiQJbWhAaGj61/28NIppDmkkWLj5xy5OKLl4wRcRusm9YzSi6
V0nBls2lbCw1BlzEOFp+xhd8c9KOjdO9NIEu2zgiDndly1u/KYioElOMeXNureuRyWVv/SG6HwBY
8XjhZ5PttWiUbY94+4DqeCbvnxq4R5e7LogULGFzRbsnIkmyezhnpOAAx1EUoq9L1GM7TgqnumAR
nd6tHzBAW0fBhBwX2H3vmP80Ik/fxoHXSbHdkano+B9ISEsYCL0DnJGjMxWQkWHjwhiYJBtcG2q+
Ibd6vZeHaftHiWKsGVM7cpEBimzHduyaw9RPcHvT0eAmQnkCb+R6or4ouRPdTidNeQ5JVGSyPSJa
KsLnSLzfVjzivotfAltWqUxS+QAqFwY39bY+6XR6Z+FCFW54eVVN0N+7IH0eiraERak4CFUg+Ut4
zbQ1+Oyfmy5mxn/Z3TlNYW9ytCVTEepy3awhwL2k8RF/8AZ8zjr/ifDQ0/u/zWsUXJdGkQ0PLlKX
PNLnEr8LeduC1W5BSk5x4AXJhHB7plHfG3Y0QV7Dlyigysa7IpB00sxQD2d5K5ZryF12iSGiSH5i
0IqB2M6ngUu4E8Yi0JQOEhFKsmZq6qimEzJs1TyfjSze2bCSCmV/LOBxrT/u1lI4mQuqtv3d33lp
2NRbzZaTHdHq9tqBvo1rzQ9sjjtu372G27i6QbvGzdLFLy6eF53eS67kHFiwzZ2v1b/egJqN9gWw
sTNyeTbNgQBwqA3faeJCl/RrM5vhSfG1FAeMYckx1Ln4y6ufL3KmKx+N6OYFr9AvzLkjoVvZUUAE
9e8zLXSZUiiNgYwKv6seQxALyRF84VoHj3SkeG+lBlCMNfIIoj/3kgUGlb/HaXxmJSDtGYdY2dT6
uyALEdmGjBc6IPHjON0gRirXphn42uQHWsWtZTMSopOIm9OBHGcYfJxX7uFUx0oVWidScySydWNL
cuyNY+bUJo9oU+qXePMypKAev0GdRpZgFJCFqY+Tfsver1lKV+qR1BR/km9oi/meOSLNj/pOdkwg
whHaJYiO5CMgVO40LmKuDFU8PXqsz3PLPxU+udy8DCL+Ch+VipI3gkMNYJG9XaUg2Bq3dr+Kl55e
gkYBC1GipnGhwANvn9tk+b+hP8nYEUyz+XLzlMgAOEb2w43XIyIqk1DS0GaeTWVS56pkofhImvDj
rbegbzeWLmEPyfmegF9PBJ8w9G7qgav271J09ltlCBqNFX9/7ZaThIHy1qXoUf+DB0Cin300oKDN
S/4MzA7KfjiRkdKITbl52tTPLgQjdqnnrZ7E73NFLsw0W3IkLTlETPHUSCbzjmpfjKyBtkHa4yMz
SppYy8Q8RFkMWgoBu1oWpHK9P9JIk7INLvgpJdyMpBwRrWoQfO1+qxdAugm1LD/7mWuo97WN426C
lWcWmhjOBd1T6nCPAKRN382zc/4wYGpkFYPUenQUndx6u/1mjimXqI9db3Iv5vnfXyPtjgAAKjon
M+fR30xEgsYxVkLg9JSDUjjqqFdANjKxGczwkYRaJqKYCPfPtTz34lEpfGqeESU47Ry3m+Wmv+oj
yNrzaou3nxEO7ks1Tv9T9ZPeepV2+8FQpTXrS/t2BoaldH3UAhDbBovsA2thwzACfDZ78cO7XC4O
QPvObju49RkQkpS5Ub54TGtnq+BBECyw31330HNgsZTq9dG0nyd3hpl4EaQTk7ZfhAHzUfy95F9k
Pc4ADWaI9xJlqghvDEyKhHstypxcog8bQFyh/crM1I4WyFJO7r8JuqOX6mubjYb7YEkeYpeziYXl
g3zzVt9ze+BCf6SCGIRBDbRzjxWO62CBatR0RDLrQuAayk2Qb9koVui/fyan2UTORK6n3330u8Xm
t+JwToaJijiwaMy50TM1WeA/fGgsiNMuMeoBKmthzOJpMz85XrZJ+xkb/vMeZt+BBFzKmE/DaSbn
NJHhxM96f2n73LuIXQ8Ewh9BjlmlscibRMkljMtJKfUaf5sMgxG4qyke3uNoavqN0/A+RXsmkkXi
1s/V4gvAypdt8Hc0YdrXD6QQFVHGGfjHIuQC4lb/d7Vc9FbE47yVIJvBGCgnjniLscD+6yaPOc5E
w/mhDHhNoy2JIC5rYDkF1CrXPxycA6ALLlkg/J2VfyH+ZlQXc9vhmdmbNvZDvV1Hx1hjZB/ZwJ95
NruC32UHXx/m9cCTKlKD8wGabvXZHVYWr39bQxK58CMWNIa9kfTYK2VuQ98pK/NHNVSfSIs6vpTN
omKnyi3uFUPwCCIpoV60cKDUZMreTkTNWQRWNMHfwacVycnUfFWnqtLpKSEhoRqUrRibTSCf3WDd
V93NgfrlLHQ6oTY67YFlxsZJW+iApmRNblqezqnhCMwiHeP1RzdxCvVJ1EqdtvHbTURwG3eBSUpS
tmStC+IDm/UMXRO8IZT3GYgf9ugVFhx3LW5Pmy6WPBsv5rRW4RQ0Z7q1LG7TigPxYj1Q13bZ900R
AuQzd8zOTWfcEAVv2+hPQ19fNX0yy2NhDiBI9O7e3NSYUb6CYqRdDyfHHoD2JRui1yxSUUOXqJz1
Ae2ARrEPd5/3HWusL4t9eHj7tE/0FmWWcZlGtu96MNJyhx4xPem49AtEb73Az07NZzDqinYFfNAE
qJXcnodMjnqip0nvvmLFueU83Hq5F7g+jRhJWhDznsB3wALLA7pIOremVDl8uVZft4b82vSSGB4d
JvAM1OvUygGRfNZ7mHsgDE4EabYDGKDUNexPj2C1Aje6mo3Chw1k5u6vrmCTZRgdatVKoMBH6dcU
9QQBfx2MWr++ndTTVN5A8JLW3ckU1/6E0jcpcX4rcQ9sU7hMDa1ankL28GN9ts9yBXybZQx7izk7
geX/QhMnh17aTpWzRZtOsJN+BEhEImytrrn47XX0mcGXFaWmvBgcZ4pKDzwwMy8fpwg3vOYIFIAP
wUjbUPlTJKK/R0YKeV45sThgHkimOD2TiisLucnBY9/sfPWwboA9jsMsHCUDe47yThWaSN09n+4J
sEUqUGo+CRA1AwSBMUDZghk4/RVwPrvvJdI92gMlNhx12Ykgr1Ebro5Lnd444Gb5qF4VDgd5M++A
kdwNMUaQtgGjB5R4czf5i0IwpuDpFDFhxXSPE5MiB/RVvDKP+AC7FPdTgq9peoxbWjQ0w6g/EMdv
xjLFSkYHA6WCTUAmmwgTnBgVWM40KoYqCF1UVuecqsN5QNknF3IKdMOgmrz+Bm/LhIdx30IkMV6X
OSOblasch4qWYJE+GIs59+7KUV0l+K1N8KqN1S/y8crR2mpcoSvAzKf41awgAKuBAf5mNrvfmpAE
6KDYLvCSirVs7kQj3cnCJekoDHLOBEt+MpSCKTKtzturg+dx20BlOBDCanp8FuRhzVF+ZQx9I88B
nPR505bdyVddAKMXa61BHwKhtwGUiAuPPbS16RT4JBQmPvtUHt5Ik0Yl4S0i+ViGw6nx8hu6FYiK
X54HOPfy7KbCUC13V8NyElvABgROZui9Ujs+oFiGlh9kx+oh1n5e3lC8zrcL39QBXOfTDWHDc84T
SHDVYnN4s0R18KquOn3+ZOhgL74p0R0BUVJc/ymG0kdLXqj5VehBg0uGJVffrBQmwU9W/5E6PyOz
2TgAhAQNZ5xx2tiLSoRYW8CTTk5jjq0Vcymx9l154wrVt8PsFPeEAqzvi9yIOBZ1pUT3k97E2DNY
KC7XTrSMOMJ0ZZRBY+PKpcWNtw7PJvbP1k+mVU/aZ3TZZfaBzXMVI399P1hxYa3nkW04ux4wIJzN
GKaaHRs0syFWS9a0LkoEGcg3Zx89V1tCBhJ4QzjgJqCNnp3+5UhkhiqEybMHy+Z+TZMJqnsP9WKR
lkoGYyutiKxhO8yB5aJjNdVv1MW4ax26Yv77gyYF/2LZLBqpLwqQiyNttjBvP+P66DAEooj+p8l8
aGGX599W0fF7pnhe8OlfhJJQdeDsn21RtEtm/6UCfnV18PUmd9vS23j2cAsSnnq59HrUJgdo5kjQ
uXOnoqw4+YrCM3Z10l6BJ1l/muq14YnyUDGqJoqh+gI7vKuAypG1gSX9ZqrW6fHqXvVSHT7rFduu
ateAChPEIpIcXnhY1JOgpYV2krQrmFSyz8QRuorl509+Vl4ChAaLkGiNOWpLuahhzcT35f6AkYwM
c884ruPmEW8M052rh5aymfIQiUkjTAlWjAWjQCx05C8ygAYjfoBbFyvuh0UcDL7mnhMxCoiFQjDq
yzkvaImE/k5NwtLZpK1QFf5uI6l7238+KERHln1Uc4n0kKR5fllguK9ghkgoCZsJAz05Z52g8qjH
MJ63G9GvJd7XKWPw9mstO5/3/NqjG5l3nS0E1myLtvpuvgFGjcY3pN8xV/DZWX5iiNX9W1BWtjFG
ejjZREfo/lTcVND/NIUlSDo9vVJxIZQdE/fSFtsYr2gbviiPL8H6/KDi55YYLYh+69zI4eN1wHh8
CojYg7pPoLS/dHtHEuDGNWNunOZr+5gP3Gpa2aR9Grme6dD/6nCPmmUruszbo8/gUghfpCcSiXmh
XIM2pK0VDcNY7bfxQd9hoXqX2z0MZaEqOF6gjIfPaGYjZHSFGuAyHagXSzWysjEHDJaWvjweoLlR
7gvgE1fITjPiN4++k5O/GXS7GyLnJ9xtUGULy4Dm4kTgxYkUw3GBtFiu2UF4Tnu4KrtXjMHvt9tn
i/zi98pnQHLYnZQNMuk3GxbyHcB77qoWr9IT3ZlJKgBr8TMpZ6ZRpwhKSqkGaOkmjLb/zIvKfBcA
e/qTYZiisp+uec6f0b5dNgI44nlgvNHYU4qY5ZZJDIatunHO31WV7vtrDmxVWezhkKO4+rs/tAe8
KE9bTMGpnlmKgG8D7eiiLA9UyPqbLH+va56mBFu7dBY4mslW/z7KyRfzoeps4SqBk8leKTpWgDTY
A5ktJaVX7SOvE/xohED6zJC/PLt3CJElFh86PDdOaSK0NfPYCD74v4/rA2rO5FAwlnNGE/TkK+1G
h5EXy7MrdDmQGw6BmxBuxIGRLH+jhqpQK3Id8t9xqdTyTNdVv/P8oIf/MzVy18Qs7QvesXKIbGP1
+eaCvmAGGkz3YtAI9OYIma1uhu/gQ4PSaUSpa8RIIWjIR04I/WbPJ+dQloVlr+7YgvIcamW+UwG7
QWuHjgKbwOl8Yv8UgUU1XVt8RnJ3ohBDN0i1xuUp1iAwNWbjPFN/1adgRyC+cP6qyrgQlzaA0QX7
1vcQhlf31frYKlIZxGhrM3mwR+V3T7p9rCFJhSM/UQ+TeHXv3Ns5cOytSQpkbzwsndijBGlqOQJa
YkAWRjyEplTnApgCwSGNKOMv+0vhChXcrbXCwdnJbGFfHBifC/Sd19M/4YdUnmyIdAWc7EVPG4K6
lxwLvCyPQeMMT2yJmO0iBuBA4CWXT6cupVHWhOQtEt89Cw79FwgZbvsCDkxHdmT6vPPgAaSz3fRy
jos24lx0ZXZqbmGSzmqPJ7ChlyX0jtXkPuAlMy/wNnspacexuWYJmS343HdCPul1C0akWtgxFS8q
+0+sim0ASCRwcLTExTJAs69nZFd4xDKCj5fsZX/yfDPF7Ci7liJtm01+dYYMCo01VziWrOJaIfLl
PLYTn1x3cx70MDZgqks7FzcOaX7YZp6KXBF5Airfycn5u0Znm9rqHqG4YC+2iQ2tVqCm0B329Ax5
olazqQ/8uQRGl495oDn2KvGxSHjajxaprpWUO3Q2aFdSGUY4Vie4Sk8g0+0jGdwIVqd8zwZrNh6X
X0ZD6lZkaUGgDQJIdvDOC2DpOChZgNrNiXdxdv+fuSlII0CmHDPGyJvfZwcd3m7L6inmkEc4Ppmw
Nf7JojluLqnzFJKv6E2PtQFYMKvRqmquJXRiLVG+szqoOTW3XKzlJl561NsmyqFjK+26jd+id3w1
jLYsYFjsNJpAmivIoKwUhvLs3Z/qafjX9MK7Iciz/lRqLd77KGVN/2gFsuD6GY7N8a5aemcX+/kR
NKH0h9XzBYYJ7RChgZTNWy0H9YCy1/HaS1OYgD/kdy+38eRSiBr4gSWprAvdfNqAp0tVc9vv7onO
3mwV+0i80g3kV9qSsBhNnLDc6JwaziVgQX/u9RU2gdfdanA3H3xX63Qyj1NRzIdEU8aETvVG0Jsd
mv6d0rfJut/eL1YfIb28gAM4TZ6W812ajE1SHkLPM2wu0+AQx7YuLyTGgAvtdnVoDgXkya3YwrRH
QU/81wvOn47kgMDFSH2d7ldYo5tPJ1jcwGWxdCmw7zbWrL8pvFxq8UMgzl7/lXvAkWL0SeYLDOoZ
g1L1e9GQ5cCD6iJWNM2jXXfd3HX6lcDCew3bTduhuZ9bPkLHXpd5zb+YUw002gWnMRavsTmf4i1j
PX1YgDDtiOODoxR4YsIcLCyuu+tosROo6SjjZkIzIrMqfX7gtC+nwrZvekuwGSyJPAmh+l07iIvG
Fil0l2h2PhHydWYQ7t37VARSKszh/V3a/YiL4dRYlborc+DVFpu2rpAMH7WN7GGRi24ed0OiLU30
iFVY2LtzMAXZ57s/Yqyk09DE0WQpYb52uVIcO3obnIAZWrr0+ftpKsYIeNOAsRmjtsWJfWeZxSGq
S12IaPbRZ4rzEOayVzcezBuSkXdScNL8aG9fD5NPgBGFAucF8XcnjiZWJ3OTz2IglZ1UH+U6c8F2
tSlxHYmatZZHfkvf3v1vBhGs3Y3Ti0SaWQ4O88uMWuVnyRV+7RjN+i+76njkOQya3yKpxz0inogl
fbM4gn/l9VtlMRpu+GsFUt1t3zdWPv2ju2qBFYx4uRAuwYUCK/n9mNXQvZS8XmJPd/2KFbaXHJGp
lda+SLl8I+9cik1EFoN1JIxXwbV+lD47sSDOgS8c10+cIcT+UkD85kOcy9xdTqOh1kyB6If/8/iV
KDO+sgsDpoILopPLbJ7k36iBAWzm6pgQylz04x/986Se+ldLoxJRn4E1jVCjo9iv4QdhgLaLFDKO
uuILNox83BJrcLXFEr/pfKWmT1AoCQJ1D1IhDFx2BFub/Q5SC/jHq7t4djYv6LJA2fLwf7pJ6PF2
2Obrytt3ffuXqPtwSERNW8D+6437FeiDxzo2ofNorbZ6v7nWO2XaM11nxc9v7semwDOjycX5qkd/
Q+Gm/5fi4iia4PZpjoh1sDilsEOlxEx9nOI6VUTbGUvOcGqMesUhcQwwbQ+NwygNVr+Po+Wg/yob
bN9iZPyAyN5uDxq/+Ut8iZtPQtXYNWlgCjpgKC8Kl8dJjF1uR9Zgi4JKGglqVpY1ZMG+ENJaTILI
16y7LNnOuLP3fZAD00C17gtz5SAA/C1ZJIbY/nkzqt6nZWHPKxz3+lDySlqUQJIvv5YxIkioSsat
rmg9n23nE6tDY0Y/jJfn1628WJMgz51G2fBEOemzaDm8m9DJ1jbGfq6THzfotT4aPuY7xLE1eXew
APbm2W95yX5nojNEdPBkyjWB3Wk4CpqXjOzvamiDCe9PND4/7JWDi4UHoIqf7diaXO+lQGLu0pEa
URfaY5JzjpK0KqNypR7V/KGwY3bVxbssMthmB90uAwtaW1r8/6QM5P++tiLX2qP9KNdPegxgWA+x
bx+SwaA+PC9b7dasH6uQUfkXDXcaqWyaYTbLxncjMskE5p7uG0lkklZBd+KTLsKiDLGWcA9uayqQ
jjrpX8n+ZCoUsdX1DhcFUf0oUeaFHjSKJGfalI56fVtFyahDWIVlW6dDy8DofcXw6+bIZpT9zuQg
qeq2U9IuFVIkjxItp/9odISvKM1NhfW2gJeqsOuaCG2zvT9D8LWfIn2F3bKO2Dc086fDp9YCUp8u
q4f1dmYXwEasCIl7q6gqoSZDFe+0w0MsXdJd+qFpm5WXTbWH/0CFlr+3XffujJ0AN5Hp85ipEPat
yenctH/LJDH/rwuiBiHueQa45bw1PzYld78IihF6cn4s+FP/TjphU/ZjAs2cEILxK7jSu4pc+03Q
9c1Qry6sXAvytY4gc98L7euZ6kh2Li7dXFLIfHHyrVfrFZa9YDpd/KesrTwIIPhXnEhip/lYz0WT
Lx9hgVyYy/mYoJwxc2qZ7+sphTdgZ/JioXaRfnQXxpWNBkCJvmBIj97ahFW4bYLlYTjZIib/6LjC
keM9nUB2ZZi5SqltSkRkwJLMc1m5RwMjzt91maLYCEs8ArbXvLIw0ETcqLujOgYn6bl7kjQ8eQU/
ZcFu3oOIBQ+pcg35HmxhyKeuqmH42Et/b/nGqyNVFFT693n3N9Ch8CIsqoird0ob09fM2Gk3NwZX
CXM8o2TPeOKJYYg7XRuTQc9FYS/EtMBk3qpxmNsL6L2eOvLNXSIjCMYFvFRZtScY/woLDijAtQeE
VbXTe/3RYtlW7B9CD4hDVRbhniSAdBXP21flxwMSzLNj2460AWpFdbK8fbIlLbamgedaUp92s9zv
A4XKufQa1hir5SDfbtSKrj+W1XgyEYYzAmR4gDV1Ruhl
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
f5EEMQ1ZE5P4p0QLKL1u7BBcvzhv+n/czwptpnno33YPdcZJSX02Mpycj42OuDXA81rMSpWIeLxT
eqpMG7Ejhp945PfgKuySmjCVhwpeYCwOOkUB6uNgIdIBPpD4Ec5yiSopy8Z/+/d0NyIrZPLSoZ6w
CrSjUPiYTdf9OEo0x10dYkCrQWZZYApuSVq/n5WeWmeXMPcvna4qmU7KFS7gKqv1lgvLcADxPt5z
ruo6a+Af07YDmTzjeSTuxRIGINHjgHxvW2YdxOdROBUWeW1VhK0ksDhwf3cIhkMHHHA/BQv64/Bh
dunpv57VucszcmubWphKiuutoxMWrZb5pIY9bQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8352)
`protect data_block
NfHGEL8SXdsaG/U4n1y+Q2uEpKO/DEDJwahFDxmijtnWVxfkVVf9giD14vb6pAIrlxrmHoeKq7sO
izApVOL8bijS5zO+60v9b5/3mAo2rt8x3eOwUCRSkX6OcaodfgBTAZqdlar7he/PQXxXS1X3AIqR
1xdySFKzLYEiYtgw/iVDVpMmjCCeNw8C0LCh8bQ9OY1EkweilQMxxkXnOpJR/+dcRYSzLD6DNegw
8+O9sCGBy07bveerYj5yTZIrTY1CL6zBy2cizR1LTwdOfg8cIZDCKXNhyiHDmVcnXtfZ/h8fLN+c
ThTzlUceP6rso4TJWa5wRJ69/8MwWeDnleQ4VSLyMKiH+rUDTw/hYmv3s0vihavT9usJDuI2ro5n
eJpS/0MAeY3x9Eb1+pbXpBsPFMgtLQp3SzcKMdMq/mFRn9gIwb34OTGQiQ8AJIA749ukwJAgzPXw
NZiJ7QExOlM2+wAvT+fMEMKeUDciNcNZoH3iuxjXMzmbxgFEca5iwhQlx8eZ09ugJlEgNzq/uZhH
J6T+A5X+g7lf7bWZOszLV7QPbO6hRmIXOFwsgX2NXkqTKtKfNX1NcapxLSt2VbDyEHtkD+sNnYxa
MKrfLMQmQLDbBZ/7gvEPmEOnlE7IB3eHzXVTmmZqsutbQSVTLPPze9WdD/gdR5cHpiS31BxC5d4c
HENnG8lIARuKkBMT2jr2QcA2pnGk5q1ecZmtmKqA06LpaJWpGkbkAHfuWgObi8P2XBBz74xnNEIi
10doRLrAF0Te62QkMQZG9ui2bjwuuS4Yx1QC8+zP7Ija/iVvmzlBcbWQdwKkHM/+Ec5WlMpb2JuS
8WIZhX9qES8p86HWkaxt7YbmgN192rGINicr9BJydHIrbCJYfL7X3LpXKfUEY9UQcaEuGijS5l59
OeMny/UzIawCrFaj9TdPF81UO7fKLpZIHruJCsjZ01R8qy0ycFNf11x2p4OXWGm7x25zDWDo3O6J
f/bmec6/+/bTAzs0Wod6zHdfV2MW/QNIEkEeH/0J009tduZkU7rZLR29M0y4W6a5wQx7qUQISDUG
TGuCjZRzPE0saYoHxvU+yig5gB45+I9RdbEX0cTMKvrUTbGUo/PflQAwSHOFgZrSN6/BhjCwBgXb
+VuVJ0A5W6MM9pGTQKJ5fTDo2gISSnLA5/OsMQd7Yc6kvyDJ9H2mmUwzr07s7CFn7QI0hTZkjMk7
XaV1Nx1/wjHgr6PD9XNJoQPsZ/7cLyWUhyEazkexy3G45AN3TE3/QKg/W9Xm1uj0oDGdBgZazw7R
GyBcKu2UOvFYHkhD3mSKH/LXgnxu9hSgwE+4RcAuTo1RZaFNG15YBAa1ATfevEHFTlBWttNsFPPw
YzSGzkB30yeaLiY4aH/ZyptiIFzcZgfX37esQie1mgTXjEIN1KOGZevC87I/EKPSbXvPb4YMuADl
OyS0dyPL+x6zFr7wLDeWGlHLj4ifOT64XamkuM6tZq60V9D8HTgOEXcN61jDMEgH1Ae79NePddZN
tV+5QVyuTgq91jwYExn9VQc/PaCy1ZFzUjxHwK+6qkiycs0hETU0d0MBRUgzip+ivTko7n0yqrcC
rn7WqsS0Cr70Oi5eI4pnZPxFCJC1toYBiAHPbZQDlpdTPi+7qujOEJawkwJUojVBdEzA9eE+alOh
44MqJ9vELQmYtCfxQr7CKkIulJnAFKz19BWfhhhzJkiHJWDuCSML+ku7U89MjLWK8WFQryf+6xLL
MPe+mP9Hr8TN+kpV04kyDctdfcUPgzFpMzzhg3caekNHXyI2RQVY/nACx21XdkwhNWBxotq60pJ3
CPsw8JKdipo2qyOSs3EsqkeweAa7nnXYcfni3XcNhZvi1qws8KUlll62VHot3O5Rv7Fso9aZeIGv
5quBF107AKZ/ssEVaPlWGzQ5UJNBtZw3/N7V60gWmmjg5c1AmAgsjYzyaCA91Ri+7t1WbHtF9hXU
yFybVImPOY33hWe8Z4u10tFW4lqpYtltspuuZpt9jnY1sXCWSV0Ha0WgzUuGRppEeQu/5u8hE0S3
ZUem7lhF+9xlYTP/OZvAwpCsmnXr2DwSz5F27a955MZox//QkPrr/VBhr0tHL3YO6zwbuj2Lh6gF
hFU4YA/Uac+LuS/rWN309OI5K7MeYByp8zXOb4bywUL0/Z6i2p1Ms6AJDMJL4OrkCZS2xtsrW62c
C/QIGf0nigCdZ/I/5VTwIcNJyXDgGHBDjSOvydaZdVeGghpLfnpCBcr8e/yWE7O/xeVCBU4Kw8m1
7S11h/Fp8jOQagN0Ekzz2tTepieDwo5oHPB9qlj6g7Vs9M1Lod4nwdS0JY4pEPDRXovDEYZZhfLv
jdiMh7yJkWn3KVK2VZZYVQRNhRDtCfU8Ev5bzrVhm+JW7VxUs3IhGOppwJDPgyP+vMihb9iapjrm
7mnYqNVzyk8uwBgWJJGXccq5o9emT92pH60ILSwoWuNHBWNYU5HhlohLhsJEM0wcyhsQzbAtUuKn
Fu3H/EZFNR2f9rpBeGYR5400Wl/17yofrUCOmSf1wC21Zx7LVkYK4QRS1PuW8dt0e6GtjEnxc8Hz
UzgbxX+nnn/U/x3VSnO7X2oZuTkVUxqz+NmCl+qPIsFXYT8N0AfZev+44IQyOsYkku1OukIC5uo7
VovHeVM4I3zPnTgyn0kyygxS+qwg0HA67QLzGyXmVDTDIXY8a4xloMafCiecOVZzVngI2S1qy81l
tbau4MBg8cqrHxCS33EY1At7A4OL2QG/uOKYGcrNt2R0b2O7RxpQzIMapvIRTOubqQX41GM4iIO3
Ke/SFDsOUv0QCx0dddISSt1wE83gvxA7MBvg3frHsdY0esczPwVNv4ifMZYGjXVUJc4lMVD2f7Kw
GV4K6O+SSsIV7fX39njj77a9hvpIgG2zw+pYlEb3626waBpLF0QuMZXKzzBzHKzBb0aJ/d2PWJNs
d2hgRr3/G3GZCn24EQiit3/vDZr7ICdJp/UHczudgoSWbVCtppSQZXqR1EVt5wbKO07SyURrwmNG
dTSJvSrqkdTBAsJUYw1k9Nb95gYC7TjEQh3xjk4V1oD6989Vm4wredvl0Id/5EkAFE8KEmX+NR/9
jYMTtXh057OhY5HMw5jNdaUkwcTdqQhwGMsQ0xfZ47OTC582H2u7ouzI+CviB4HkdVrRUSRn1Ix1
+lElXCnFTQBy0UD3TJJs9OTX55guph+gizhOvowZvWa32dcroAIZ+73kM2hSh9Q+EIYwx/Lz1Nbm
BDpNJDHt4bH2OBOdu7WtdBe5Q7WY6ekVO7ljX3yA91gQshEcBRS2xShkaa9eupHsNwpK/IKxucfU
r8Z15e4/XKBM8YqmJC1lWvQbx360/nywvupZtFUMx5DB8BreG3jqR6E/8bKFmNmNGo1+j5Yz028K
1JvbTkQo61OqRCK8etYxV49S9oY/mlAUYLDqy5/8xrv9TRF1kdFtIAnKK8gVlupFpUUhcNbC2+GW
S3+7HfvUVvBBUJKUylQAMrDf+Xspu3U623jIFIj3ffVQTx3bof2DZVzF4b+jh6aoCyRjFlf1W7V3
/hxzsduoZMADLyS7SOyOG48OKOnaeewtrOIhui1gFGx4UC8s0sqjv2u7lVDa2hVmdNERXUGHlMUg
3qoJ0uLHHH4DG6YbbNptrWHjF6Z7jVcNrjJCZN03zaB0bUzplm092lbLKOmiUdGr8TUBtVs9LuDm
bmNfdxAv/k3ynblzv1UkA7yhZhTPMjJO8tLCR7KAVIMH0u6U+S5OVg/Uc16oZaWHc0hfGBYUGkmB
3sZb9E/EroHyYGWDbU19ESQomMvsddxlgFbcq9zW1O2q5C7Lh96hXm57hxGc5A6btOmwBrTl+6JF
cupe1E5r1TGAnQpXG2MltAYycJlzgrG7Y7ZAKRAXt8us1V5Ld9s+zBz8xlavSpN1PuH24zGWWs+Z
2sxCg2jf0LpOTgak6Faax/d/Z5RI1lIyIEJBOGzSsWw6XbBvhsMm8KZsa8IDM+FMeTg52LsUKfco
P/m63OyLU7mKU9tDrtQkEmbSZNBSL/1VUNg3rzmZvM+OpkzU3l16oe9h4M8Pb8ID4Msxp360RO5k
UMdOPccoOBtaaQSPjozOio+z+GubKWD3+oFONwCl3UKcEaRXapoQuObzbnSFo7RYvXvog3RsmRWL
CS3KCaNagRgVltSKW/VKVtZgu5hokqzFV6DFNqw7PKf84hR0Nqmqv6YnuilS/as5wkQam+1JVltC
6SQ4o9h5oBdoCPnsMc8sN5gQWWqbFeNwcHIquAsnD8XP6OA+F8RwjO6U71zDPJgOrESoZe72k2il
KP2oUcDKC3bymYt1psoQDutPcf3lpvIWNLc3ntgxKEicVFLl5ksi3N6wjOfjcTcebVm6cEoqgDGM
mnv+83Dh/8OzBqkMVzYXxEtGVGf5bUztQPaauF9fubPBF6kpRoOTecxISJILvDXY444A9rXOnMGj
kybm+fhwFUB6fB0nvXcji5qdhV/m61gtQzBlY5Fr4mPQsX3rlcYSJsjBRCHIFG5f7HF69sDDFQW8
onYjTryC3annAf8ex+p+VLhK/Z6Cm1fv+lZgaN+RxejloJSJV1CijRFOJu3WG5lBAu1On2DOJZJi
AWNPVicdL/8MuwNRu86cjbbec4nXJ+S5he6nz9ywvbWucYKASdWjyu26SDYzc/qKVgsqClkQyxb2
464X9kwxbAA4rPQrMQhNBnxqN58PkkgMwX+Enp9BB5/uLtEcSBTi6eVTb5E4Xz6oy2uq/43z9G9k
KVhPvDrauuabl6aHbeysRpb11AUeMpaOyv7IaCBGYYKdsN2EasaiRqtQORwC341Q4t7WSxSxziKY
sY/4KmSNM3IMoph41B//O9urYJZZbE3dq2lmvNsFk8zvHBLTROw4OADlPy1J8g2TkX16YM8A5ATq
PMoQql635oMkRpdu5J37Zs8KzSLqeVcX/e4w/et+/FOS0KLHpt+gF+XyPQmtxIvZEPkzeBfYA5Mf
tfjsBuojO7ayVWMq3spHiwSZh3KVKgX47mC1BkKf3WaW6XGfbxzk3SxoKpvonKYopO2vvfbwPvNh
AykBsVbkxhA7XKyTDO5i84ppTC+2eBS/v9R1RXZvak1YjmE1sYlXghbzWS+gjkivY7ypOuCs90gh
zly6bxjT95i1BNN0r6INK1AwkFrDaSkt94sxZ40I/9W1bR0hMwVEsqUmX9ky5F/6/Fj5+V0w61YF
lCq+twOIKt1w4h9gQErMMX5R0bKGk/kyYtLXVZUz6ohMS1WlaVuZm0rV8Ai6M+k2zdGoYLAMqB32
fTY5TGjDYSvBQ67z+JQruHqBgki8Ad08Oa7E1hJvfXeEJkoCN/gwurZsecznWXT6GIKZm6EBJnam
NkkL2zC/vbxYeiuROuv+wBqEcrA65itHogLn7JNsnapVnRtcmnGO8TJwfh/P3TnbM+LQeqDNbF2u
gwTzq6Qe0SSnqZkRLjSLyVirppJm+K4ojJBGPlETbsE4hAboN0L4sMeSs92jPzFHYDXpEglHXLEH
MSiprL37AEdU48el4Kju3usJ2z3BwBKuRPPaAXJOENHtRbtc5vxr8esXtlhcawRUIKS+9wApq97v
4UlCrZDKazYbWh+jV7yPZfVhtZS9Yq+sElABh+C624ZKQh1KveCfUG640NOD0cTTxipRhdtxLe4j
8k5Th+vHj8YC0ym4fJgv4SAu20Cr5YyDhSjWtq63+MBaGectyTf9xG+zCnisw5GBb6qqk+pDOzvG
QGvZDE0Bt8hm0oonDeAoa+oYDffUwiT7Lk8YMzphsul0R2gyhfDvV7326zsYPfT46cziEfc9xT8B
FwSSjOXJ2ZueYULcCe+ex3iefDwflmkVQwVaVHDTrBRwSjXhP9/Ty7UmPntcCchvRmiNSC2o1SNt
LOjaW0V4rIkwOieozv/XNJZrjxn/l42TO7vq6f5OsngnNlW5y2u5C4VWwv7WgNPtzWaZvKbAZBIN
H0GUqN72NgFRTAUkAzfRuWtMcYispC+WlAl079MN7pwHCCznbvVKN/NENR92V8cLrEMG0IXKr2oU
ooToQipxAa3HnxMvqUdYxI+LwaEonCuzxgjZDhVhX1B604v18cy1TpjSEG7Jeg7/WwvwF/6dYOkG
Q0TaevBpTmC8nmY5PQgtwdLplaq8YLOuhv/ESD+oXdzVQ7DBaZ7RWDeFlw/6ZwYf+VqxWPpfWZKL
WyR/zCjNNfxDCYTVCSQjHWK2dY6sqyvDG4+SvVXt1zX5mb2r+QBM90wrduBc31fq0CmaeKbUam4Q
rt2Js0Ngy/1b6/nAJS7nINSWRZBhd3DFbbO5WXSohquDUwKBLOslR7wChsYlIODGB5EA0RGnZxUo
yfLgsJRmNVqlXsI+B/q6KgdHRLOvTHb2Nkv8Jg5qniM82XGIcmb39pO7LJjdSAVf/eDXbGsZjjgL
xfI8gEi1WNBy40nX161C/vwlva0GBN9Z4gwPb21Vu6RK8HIhwal645nIQg7LeSHA6qd1+QCgIn1b
M5YM9aUuLjafObmKxZMr+/Ql4uLdFdr68QyV/TqWzsV9NDT9msDoXmQftA9rT3XnRZo6zoXXGf4Y
Ecc59MnGQq2D9p9OGOYxwztbUuMBb4K2vX5B7e6sYPY3WMifryuHzh54xw3lOiEJ6MQCz5su8+po
+ptzNN8D3Urvk6n7f/MP2stzzsZIo5cxmnLPbV+StGFZQ3hcJ5PdUdrJQaEvfSfMNzVuqgyxyhN9
6VkDIKRTos9FStbPT9ySSl2+JVK3f+kLs5THftRa8mMDQXgPW3cuoZduRy/e8vgjkNHVwKfOZ6qW
syp9cACQ+jHKcQadvuFaccONWrSU7bhiePVotcSrvrYmiRb1kULFvcTe2Whgu5871VZ93Bjb4DTb
TqFyBOTkrU86UL04S0P0+pDGL0TtExoGO8215CzaRDX0WK177b0lolHfTYmYXnd1SuCxUlPFPDh+
iSpoTs9I/a+3tDEH9s611xPCv6US6eHVebIo/NHZpZj2Ha+Z5FzAwtHRrrH+2qLu66BKjiiHSeju
8RbAqgqOvgk/xPhI3pA0TnaxhwS79ZY6mik5NZkGuCebTdjrx1KkWEnClrULvPDZKgT4XPnQjNNE
H6iCz3i0TDLCnBZ5oHJhzlPnCNUg96HuLPxSATlUgzjTO6GFYIiG7/rDEqXqn0/aoZRWzfGkPfig
YBxeoIgTUIimJgHyav4zL8NBm0Ke8ReHQHkaU1cw8ACwqgSrmxJ3bG4cx41LGYuKW42qp3ET26LT
gWYygxzSU1f4/zl+0Z2TtWLG6+d9MRDpzvE9LUpyU8XLMf1g/sqdQACmbkDaKRJOge8xvxOTXsN9
N5FWhKIq3xo28p3T6yZNDY801Eid52G3Acn4UjUfD0oGaMUSwLvdhSWUcHKbJCx3G/BRWdw9AOPd
3ZDXUrl16gNHr/C3OfLHFlrWJ7aOMI6hPYMz5qKaXBvIGNEDNut/J71vYsCv/hS9TrMaCrkhtAPI
lXBeyPdCVWG3swvFm/OD2AKVojS6T9W/qCa1RXI4GqRLt1m/68q4k2zH2hxa0sNb6DuAZTCxVi6g
wQlMBGWvEqJi/adFrarKvMeXkFIZKlS+dkdbA68irwCTOQMm6aRF0LppQZMxr7aiyZnAk+ZkvaGQ
D1+9doWSnAN/p2xOe/uP0QHBXn/pG0y+76lQM78J3kDKnaKGnvTqI2Qe/ZcriMTDWSqBSmeEPu9h
Wmn0FT8XwGp8e3TnYViDNFz7Z3z2s0oujHBd75oyY+JEFrhFbvgEiy4AM+XH9CTdKitMvvWB3syN
ppICVZBWGLZ+tQ+4BccsZVAJDSXINy5XftQTunbsJa6V6RSCFnHO/3R4yMpjtXbHGLa0mdsSc4vI
+6OqxaHym9FhuepRZloWqSTdoJwg7RrsG2Mi1cEgdZOUQOMaQUD8rSQy/VK/89tynVcL51UmFpQy
WmWEduyRiPpFmRPax4dQmdhcK2uuNG9w/yg/jH7TCfg1LDaG6uDnf2P6FzaqmBAB7jyJUMgod+be
t7rswx6LUr3Eb/qzoVzEWUH/QGsW306UfXykVfeJvhI02CNR9XJJ7YGpkznUzQX6HZu0SC8tvv+0
RfS8FmT6O4BWK4D3fYf8PLETOoL3EyCSRnZDT/PbujtchZXC+RkfbN7vgwNO4UlnLunCvn9zbqE8
4IYBZB/2Uy4WWjX4JT2kclyQ7BntJxqOjMf/5Z9VWPhWxAc7SSkrKwtYlrQDyNZJM3g0yRmli5NQ
x2EZ0vS6/030STa/RygxLt92WPCjMCxDL5MPe2Ef1Y8gK0HoWilpnocq1loisYEs4ncZ1lfo/ysK
B75sOBu8vXiqG+2dl3SkYcaL/YfTxmDosiOWTjf1B15akLVWNRZ5YLNEsDk4SbPNOdKlNZn3tt8s
H9eSxsdHEDaQJcCHyH43vR9TCNkd965/M54k+iA9awBopZG+4Hk0DonrxyJ05kqujj3ViVdTDAWY
o3/k0IoUrDDMYlMKLzxcmU34EpPjEX2Cj92ptXTIEAmTEzr+t/MfyPkTxZXMND7+o3u4CYLfHDOA
Bs+jHyymvuV2xsbITgCnmwXLk9cdo2FPhvVD6lZOlFo64j5cM0pXy1a6FIwD3h3nYLbUbQNuMeAz
2pree8veE6aOArFKsqNRTYP2u6lxZ3vMT9o5ALyRMHpPQ7+CUyX1nRStWhKPsTW0SwaRzlz9lMtM
kPdhc1eIENEQpSZgkv270OMWffPKdc4oYMF5zEmmKs3ArQ+FZEDEsaa/B1H6KwoHxRKS6aPb+cJG
9Ipq1m6++YQ53Eb6Ii394dwbJW2vQefhkgdxqFoMvQazizIKHr9PETunAmJLD9TLfIrtzSKMABNB
0qi3dAD/7VNBKcvFXOTbhbJSzfP3Jskg1zvJ6h6T6ost9xJS3hPDCWqa2DdlvHAcJH2bEkpS7wdv
o911BRO1Cz64lN/c3P2oqBJK51pUFSQI210xEr6jAD4FdNyExzxP8LZ5eRXJRLJzgUQta28m2Hmy
ffCJQjWvlFtPIHz6OZvq8R1OLbHznpo9PEJ49lKRyW4hksnDZIzim9rgejAWlTfyf4FFAKQJ6Hja
nRo9zXXp6QNwl/rWZ2dZqBPWLiCNFMxOzpzuimkQhsbg3vxuvRiz7AGfYgmU4f1Z1uki49ywhfkv
Nvjwey33VAcotVeOm8kTzOobNDRwbgtwLRBbj448J6hfBDcq1BFky8qyuNs4VjhgLA6MRWs7BOER
d0iMEBfzQnAFRANbdEfEhHMKfATNrRDsPeWfF2orz3jl/fZCZAXjB5rOzK31nZKH0zR69Drur600
kIOqIek9tijb7J9VD0BQa2iRtwmNCxzs/w78PcDGDQKgeV2VuJnK4XJzioXGNFh21HOqctHYl8v+
fkUrU9d6FhnnZiMaHojUxByhYOUMWasYaNohEQVgOfMUTuz8h2AmT2IuR9eHkqxs0PNGpTqopELI
YlgzOQPAWAIm77PIHo5F01DDjOG0BwYZH/3ijVhFypw8Xhu4TiiTDngFR8n6xhqDvImUn5Y/PcBM
/uNg/tibgTQyaF7EPo0X+0e/gDlriMQeh3mq9zknEejdMbtzL4eRUcmznPjJ5YIk3jtfgpf5T/Nb
U1lfVpW/twmy24w3qoJ4FKAc4N+7yN0TGKwndT5wjmTi2HBpCZAjrkMnCP5NzSVbNaiYeQqXnl1w
6xf7nEcjYtq09cAbgLbYxrH97/dVueQetHahj7P0cB5wqUgFUt6fA7u6KYU68oaPkHMsWdxSLJFd
lpXNu2O6ZlYkklk/M4qvb+w6h+gfdh8M0uJ6BEOqge90jwWB+94vNXY10gASHn5f+E5cEil1r4dQ
x4DAqyk1nqfeXAD9mvbeez9aRN81rfvkCO7RHVCuVxqT4q/jfXN11QqsuboCxhoGDhLbvLCKoxLD
65+aTI/+0exRnQ/+s3Rrw++qiLCTfbctu4DHPdrmrAB6Q77ps+dHiJhcDPe/oWYFFa14jwtgoS7X
acJYhOY5BoqLvXv6kcRAfzFWYTKEpn2P71uQgkSZztTO2PdaH28anCyM06OwL+nMa/9EL5V51lbP
8Jfqaz+wuI7KDXQrdrGrqxan3lY05kXTTJnqTGpvOfXFtmWyS31oZoi0Bphy0QbZ9Lb2Io+feyGV
+eKIVKqUufwlitilb6ZMGaNAY2crJm/MIKXs02idpuJEYKQnyQkxyxUR1IwOGpcw0+d6XrhTbVVt
YXrYwpRgZShef2NWBmmI7RhpFwzyobB+augPY/S+fmz0OJWaUjpDrqi8QViK7bYFDRhXX5l1OjEX
8vLHWS7Ql68qWSxnkcI9fCwzUontHaHTjWQlIObO0vVgRPR5mAUhwREEtZrLBhvJZK2oTrEh8e04
Z27b/RrVgHtmgjwG4htHWWdba+E0n8Q7uNG25VW93cAJnjD9PwKogg7vM8p1PmeNbDYO9AKvOUyN
pop5gAssIpMksKs5uYY5Cfh13uFbfx/CPNV3T6xkIn9xjfQ3M3cjuaUicfIcqaN3oDh+2CB5YHen
bnJY3C0/Sj7sd+4deQVfeqlqgi0TD3Dc3rLbwX1JasrF4K4dHJYcWW2gI3DHFDFvckOvnoKybrx3
r4dxx4QWC4WyoxGb1S/0fm7v3v5Jk4qplwLOeHfam5Blwf42gRcLIOWSpqgcyusnPhNpHFRVxWGW
BSn2Osqv6Y2/0B4n4oKV7WMhCg3tDiSCq2/MO3HjjCv6Iwv/uiENaQgG59GN0H8MEy7LxGG4pVo1
2ohAtU3ayT2SeS+7nmwewWXX81mA7wjy7k/bgqopfNlX+Slt/dxh126Fhh9nBdp0Taqdpfx+zdfw
O0zMaRYoFAwGHUpx3vAou8Cf92byFtt5iye0KpzA7FMJEiMXNrmF7PyzRl6lQepuDx95B7Z7TM0Q
j2oP1xUwlWuNX7PJgxtsNU9L869IY+SQI//cFH3IrX3u+ri8iaWBCEfTbPcuJ5RoDhJdZD+7FDr0
cey6M0PSqyoZ2LWRhDEit88ov9pCE1yVwWshxdR6XzrjYKIM9Pxm4RxBJ/FLx3N728BpHCq0dJyV
ACnF5LAokYYmZJlcZ9e8LWtWFICg0i+L9/O6eBXV
`protect end_protected

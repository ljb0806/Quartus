-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YDk9IZm8i4s30uO8VZRTv0Tj0A+HkQD71E7P40wMlfMbJPPf2Yc5bicDw5TondzxBTqGqdDp+E2L
2JCfNf4qxVHVbJ91KdbxW/lq2JRSzW5M8+p2hJArHa3kCYKKsjhi+mK/LXYToFvMLa/7gugl8rIg
xDS8/9vB/Y54P/MPn182SOBb4BMrSCMVnTW1nBEtL87AO3nWUJaPcZzXGWs47V2St/qb6KBDAvJ5
B1DFTE9WhkUzG7oYb+vRohFDjU5ATiM8v95Ft777hAV3UCI5O40vpi8BIm7jqYSCBM2CGB+Bzmzj
Pg0sYMfNkzuK/l5PFzMPuPw+0FAfpOiAKtpwiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 40224)
`protect data_block
3jjMBaM2j/E/Z034pAP+Z9Z6eJscfQKTU6JX5FYCN9EExpUiomqS+Q0CwXBrP2UaWksdiT1vdFFb
CcQpAUzd6RsngLpQsynBeCsJ+H2FSh8KjsLUREbZOVB1vdjL5PULNG7ihQfzxd/4KOD/TatOox8J
pLXEdXNxtv3JrGeDgsP01aR5N2l0cQCEaRPFxN5sewoEnVBkuexz4eUM6TVKQaZQbrXGkfxtbuzP
B1I4mxrxzMZPCdSIe2Svn4GwzluejdnpqevBIEm7Z/589f4j96YCN+rmitWY3dpXg23NlsPhj1sI
+WssHvjtQA0sVro7P/GgIwrru1kEBrf7NjWC4KDGzGyyInqdAOxhVHdgFhxX0tNcvXdj98p8ZS1Z
ZF/MoBzqkOmN1UYb58gmVOBF4nXfftxcB4Pali0vPYYHtoTRjjbIvYovt5UrWR1eB7aB/1sKrgcI
BlFOUlHIV9t7p1txLB6j93FOjqp+ucWQpgjI+4ym6FAD2jFNBCQWqyygkGBvqzZekBglUd4761Yk
fddlTtGXE2C6Ujz4mzlP4Id1nPoSF2TEPdwb9tDYr3nkQ3nz19yVrRcTZ3jCgHzztKExHOKJT6o5
7WDT5gjYOFUY231FOedUIta1XSvzeaOqfCapF0uHLXKg4Fcch6CKyq/3hYSh1jvLwcrF9MYCFBIv
dBNXJl/t9MM3wQH8FspPuUqtMHX9p6qZoFwKib4uSgL5LbICGuLQdRd+TkX1PbU1CjPoc0SiZq6+
F1p7kOePfD+8lAbGjKOn5D/IW5Vxlcltml8IC8yfyWy7nYcigyPyQZ3HVRvN+Z1RH+Fr6Ho4fI2L
49z4diRP7+vhfhsS5tMk40qBLk9NU2AdlYQKppUwqKHHYNQgHq7zDTQAhJ5r1KyJAOCXq4552A0g
HqOz1TPRcjJ8wYIAFgjbMk9GJc8qeoF7hC7/BY5adNPj/1kSGJtBmHdotHoCOLyZDLEzUzNd80lP
FZaFYfOllIYCqUGTcmCl6k0/Q1G5QRebD468BL80ZZQexWVAlBu2OtnYwq7Df1vhSVWi9hVdxXJ7
sjCA/VaeTGST0cemdufOs19qZdf0frHeMMXeIm8ysR3Zvp6kPpAzxaNMdOYqir8nGMQYRKGK+JQ1
LEVFa/firJGqkPyO5FNDqgcOgWa56pOxfXPZjhMhZ+A6ZscRbX6S48JvD7imH1u7Lv+CkW5jtzRt
+XVSnmfWq/my5SoSOqkNYvvwXHLgy7c3G8rz5US8R3RdSYPwV+tbJQYaiaixgTs3K6eIKaurMsEQ
KnKEACS3xNg54l4RHDyYHHpe3j6XJi5oSyyYlFYad/a/2Yz0EMkxz4hKzM73ow16ZqQ0uJZZgQWH
WmyvYzPaRAZY8F42zMZMuKvsqtBbn490h0j3FEIkjyqDeqyR6YmQpGuaoBmQQF/CG6lKtQIEbZox
F2CI9TVNbjrIDLXR5V/WZVfR85fyYE9cljjlM0ec6A80QP5UH2kzydXDhTAKvBQob4wKn2uUgwyc
X10q5sJ6bYSuPOaMvfhVMlLoQW1gs/VmVM8JxtIrgxkrr8ZCkXaUSc4yi2oB8iUwsNeHWxrKdQvj
VYSsp6cH2/q7Z8fI9FrUr/OP43ImjBF3zePKoHeiwlgzZnC/DbqbSikInH/xrFfu4DbBMzlzt5TT
tXTRZqJ3LlHSyxhaaF7pYbmI+Xhw90xlFIRVau4nS7LM5HJoThsAUdDb7+JQi0FRP9XDKcKLZ5v6
kbjujJM7FYTeddJoUrGEGxgnS0SaloG+zO6/ZeQac0cl9yhqoKsBbqwec72tYcZ8o8OvrKm2uVUO
OMMyx5UHssV2Mf3rSlvGcBfMu+GtvkzGrJONWL1o3a135+VMfZJIHlS2sASdsRvhzWSfOQKxwPcs
5wxTRbss/wDjU6+rxmHDh365Qs+Higzqwi8riKvh0O2MfD6veS+r+vRySGa/8WwUQQhbd0M8bF99
6Pe5obf1rzRlpF6caQH4qkMhG3bgiF0Dr5MDowrmnlyEMhwOgY7zEazI+TIfG2SZgMNNb//T+wzH
IR2CY0MTBAF4j9NfoTqUZnycceE5+l29bCMymYFpQgtKR/kCusTUL/f3LqinN2Rz3RO4+UnJqCsL
J29vXaQRrIHfUrE7Yqf/n7vRuoPq1cCGXCaD/fv+qmVGxNnZL71+kWW2u0c6kVZbaetpcXt1rt8H
vGf/EQr7P2G5PBdi44yUuME95RF9oCHy53DFFPotxcuhtQO9nsN7sUMWUEJvMbzr7zD2r51936Az
bfJaDz9nU3wnc/ECKuJR6t5tI5G7sKM/eKHh2t/ZFh2O2R035TK5KaR4xhzuWRb02C/NaUZMUuwB
QKZ+Xmu19IFr9bZfGmVsKvGRORe9VzX9bTZ5hpSh9CP5tnFdhgguGf380CWwu37MLujghMjb7LKM
SFsbWrcLL0QqGBiRrrm3T8Kr5feUckLTtFwPZW7YoAqpJc2zk4gi+sEptAx36khaL3wLmL0By6Gz
b7wsXmE2q+BzHsKGXmdAo+T56PPb0+XD4bkhVBAYWY1+ikJn7YuijGRniGWxmI4T3Osxzw7isPcH
o1mKQ9TKc/OzCHyjOF9LyEFCyiprckdYN8mg4JxRVLIYqIn8FAudR+pTFjQe+prcMrakgJrgVcnP
UPsBy9Rno3uVV6tUyUJaw3o7g5tszvUc+AgNmiDt+ivAedlnaLf0CaPmsUKMmRcGtU5zkdnfPBMC
+AI6P/mwxD3+qQoTPpmoDcrgBNA7Bfkl0LlsHBozF3ZetqD0sl5KZ8M+VpOSSFgrwHawLjwgoUYW
QCKfQADgLnEjkncNhBk0ZLtX7+scAdji4Y/FBfys/tsH1UL8MM5E2BbJFfpYgtqhX+Z+darId9DF
+cEzWZrAYqqxyBcpnyuJ93m8CNOPyW1Yu0d1ive6EFpiQkQoXjLmsZHWH9S/5byp7s/Sr7bV2SKy
FHA8EBm1ovxy1DDwLYWr1EoqSXi8Rg/5z8kfmEa0EYDigK2z4k3LuhwF7tJkBlMIqzealzHzTdoS
5Z2NGtc/L6kQ1H+PBADfL1dipaXn+DGi9Xt2hBNzjRHsL/OnMgMtqhcwh1Tin+UaykOKMx8/Hi09
9XRsC9pVUBsD0Zvaqgtw/e0zeeFFX7Tm6SfG6PGI16QHj1JUu2OjZC0Wu9R6Ti6bTDmu3q4cVuDk
ATIOWHtgtlwXqBPVjizeLNfNDkv4arqMBHizQ6HScBpA44LY8yLmEOK9fVr0or2W5MnvCIfCSh3b
fl2xWPLmFzh+59S7T2TxEQCoODpZexhSHNvWSx6nckWJCPRlnaZRizcWllIK7Vkxq9mdEzVBlNye
8Mi8Apie6rz6gNEWj+CYaw54OdyApmi0m6wPvm/22ym8OKSUpeWngpIHhjPOVm0LVnlewaL0Q9Zy
18TtP0OgQZeiety4KzZUwSpElXO8vqI7YkBN6rBVfZVREZm6z4FxFD7vf8W8XCOzHJuzDE8IkEjs
z5nczVJzs0WWOCSysfQfoFTym+BtZIfbFpM1RAgdGr8bK6sKCoI0IwMCeZFwY3g/N+nRMGJBmHg/
LNOJD6ApJg+TEsA+4sI/6wx/ih44PMsFMdTB1cPSexLnZkqD09QsPXZVIEv6ZWrVdvdabeZ14KBd
OiL96boJ1JwVKTukaAQYg9x5LG7N+bzu8QsCmhGinleVhgUJ+vYLS7/uYOIoh0KPBfGdBTLIqbou
OoCV1zvHiFeSbtlSOe/aJjUSz3VxedAAniQDtyQcpv4AFKjyJqJAd6E6Gd23RCTshRsaK5AD7emg
ekeyO6684wIk95g5K5jdLVD/WU4xNxwAFaVvm6yUMz2Pa6DKAaDkwcvOTBQZhdOtOcZlQRlptnlu
X6+KS0BRB4V1d1vYa8nOew7kHyxTvau1aNTjSl5upec2gUziAbhAY7SmbGmZKB7pE3OOJ7QcasBa
bRj8HngcKehciFdDTBqCquanbhu63viGEGfRBRdr/YBtk0mh4jYUK7FxsXIVjVATKslUnLxl9/yY
HKipD5GMf//HiVT/WctcQ2JfH6AmJpDC9RBkiNTrYOiscgiq0Mtin+wlZ2gV19ceyl6VxFYw1GyT
9J32CHMXhAuflWTeC5Vt7jetRxn5jToreS+d7xtF4yuGAt5wuTkzBeH0eBa/+UJ78hV2moiLA63q
FxrQv8ec44BexA0lFGcieZImQDlNRdkAU9NlE2mwvS6a48aX236m58GQTks2LENW8xOe1lWNJudE
Elw7NlhQbjM256pYu97fl3rCmyBvU0wATA+NB3g/tKBXD8wtXCSP8xIWnfo0eUAH+I4SOqc8SJBx
cHmQJn/Oc7ADg4BE0H7ulD5cGyFny8FIAepAf0s2HT9GHMmR0ZVpezWOSxPRZjyJ6Nk6gM8xFwGE
ValiKqd9tKlwNyCve+X/6Y24JsVHO0O8gmoAPiBMoh67KhAFwG+45ybo3bVm/IyAuQxXKF1fHbYw
9RAChHjR5MRGufVjmvjmcLPYDJ00b50x9sspnSMT6z+WyIhpaFneRhUWcJko1AkJv9bqBldyl4+3
8/2uw0VFTVhLj+QFfEOnwIEs8etIb/U/Cd3KKkZ5wh1K3BeE08wz3q2rWBIBpEOdgF3KVj3CjqBy
9s43inUHXNM1hkfMQEdjnmbgYCl22Cd1qTj0S2QrbOas8eURjyisTeu8qaPqur9bjkwZZJUJKzbu
IX5T0KZxca6p8gskjQ25NbyOwP5U88oKmMaKOcXnWVm5AAdvsYRAl1GNcb3+m0PZBRFkbO6WCarx
bIPVflQQb+FWC7+oIBbJuqRGOs8mtBddiiYyi94y25bvadwXJNfJw4p94yY9uC4un2vje/cWwZ85
t/gfMhrgafrSFBgjuoT+QlveMsB+tCFC3GekkWHem2Hc5+OLFtsXYzkYo3iaTaQSQoVuO3PKrEet
1kR39iVswGeWceOQlttPMAReFtnYpqvS6W50DFiFGIrWPD8tOpsZAROjhNAUWWyNRpcmYvFAz112
S1Wdiq4JrU9JTj7oVsnNgWPOM/hOhJeYywWvNipT88KRsOKUqfFKTv5ZTJkEvevrG6uRFFuoWgjp
WWbUkD2eYPWuB86Tmbh45aKUAO6brStj8HXa+NmNH8jb8bRt9xVnLWFrfI08Z2GlbNAVwXecBKsf
ngY9ZihGwIqGKUDmQBMwQ+ty7t8atOcMc4cdd/i9xEUvkOqj3b8KiY5X0chShSqiMGCY1e0/AGXr
0iwZfIxQXqBLgGGaO2pt8k7e0z6CaPIBoNdV6OicJaNjQWH4iOa3tIdAGzLE6erwByWMMiv39T4E
aesPaCMkoeegeUbxhs/JxdrJv2PW7GgdhMA7o3p5yDzPPBWNBvlLCQmh3PbpW9nQwJN0SICbe+Q9
4ufAzBhGaeRQ7J69K8+HbbwPZZ/fU0GyyeviLph96QWor07HE/JSoJZ6uo7//XYRLaRyaoUja+aQ
eJYKmf64J/VOOR4JMz8oGdBzTec+5a1KUDJK+vsC65KJ/ju7HvVI7GTwEIJkh0OX8hpXRp9rsJOQ
zgtsTT1ziRJebnu5CKsxcb6/d3pszwEeCEORTq83/ceA4HHMngSy+gtoR1DFiuSBm9KZFEnu4OIH
63g8fy3NvNKBENJH/W4EH4kshZj7gQOLSFCQITmu45+hZvPPNsdptPLJmC9k1k00YlnrlGxj5r7s
9qwnDFa5qHK4/kL1jVhKumy3W4a1mHQI40xmF5sC3NPiR+T+32MBmwJVkplbziKR7UZyN/Xk4KMj
MW7HccMiJq++4GPwd4K0/WtQsTGlMvOn5WrFW1UT0fDz32PLDhsvFRvGb0zyIbzB23pYPnp5tht+
02FNY8WRr4XWqL0/lh5NkshuN9vbOfjttY1hbob1twJL1D03Drs+8wY5PHjzDWJr6uq211KO9O6L
UverycMsvyoo1AY6Zn/ybrb82OUmpG8KtBm2frkCjgBHLALk+1Mb2p2ctNZvq6BABvR6UJpso5YB
AAVhaC0GhYHKeJHtL6ln7wFY6Kfk1cuNU/gEDmHS+AEDMRsLentUxd6ETdkHvkKeRZLrXpiFDmLZ
KH2AkjBHDE6B/SnmEHMwnr4XRPFCkcQFckMNBV3bFhUAYFcmaxqcx0tc+PnxCq9NCOEBuM535lHS
Eayxnl6EWmTvov11kSNUu87k1QO5tNq2KFLOL7fT7yCSa8kqv++4jbcIBZ+trtY4OSiF8/kl1d38
LGxQVS5p9/4GbXpHl/YaRa058B57ND6Ph76oTnkCsP31d4pJsUfc9cZPzId2o6/pjXmKw2C+xHlV
Ni1iT/vMWffZ36AKRx5sLMy8U9lchXUaOGmsVGmJRObKQTvD47fADSUot/3kgvjU+oPYtgyJqIwm
ahl9fmfLLbX8fLtA+Oe/chYec/NKTh3ivMd7Mn2nIndW+otkBiw7QIeAtIUk0cG6RPA0j2CwZsXU
sZTJw3HwaTqSwdvdNHolp/mm74WFQcM6KKteDsKlf68kWhlWw5Fu/K8ryL/IYuMmc5rMidBj3EG6
AwC7QXmE/kqI+5/AEj11b1fwNwqI2UXSZfgO0ACt+RYlxwVXqGRasGbL5Ymi2qKnEx3Bn1GDH85+
MXsQnDa15CuNmxMJlGKTenmUbAzSJy6XpmZnd520XE7yUasyqbOx5cY3a19SXgO2gCoRB0DgUPJG
OoO2vU9ZYF4E231PA54KwFs33voWTqcPG9jLI3a++VyckdZ4PobbhplAVELg87yBcsWFFDS9O8K1
fmKqYpjusaSbZ7zT/nkm0z90KMgOIunRiHXdPCqiAy+hC7yZovGzuVYdR6P17sBET2+q2FICJKRs
6fKzDhe+w7At27UHyQEEw7f7AXLHVm4GTkf47XyS3hwzmN/4ct57o5GdZiQdJW+taUsTfbC/S3n+
jPzd3Jip7CKgIuyB7/ex/UhmBX0bdLjzjPvUC/dBvzPTU7WoeZ/OdAulSz7SGRvYTdNsKdTSUS62
3lnB+uCeApqbt9Xf5jn3sdwbE/ebfGLFnMVVFBMqvyM1Oz5e4LdiW72d/sna3zahIKmJOyONxkOs
J+jKTpeCvC/OHJaS6RX9XXnfZOQNjcbRmPbu5Sf87MK60SMEOcAIx9v3s8oPIUGZhW/aa0aPxJbo
JRpPqDX1svVwNFjJ0SQDo9RWPQ35kAaaMzI/7/FZOpFkn4OgIqFJVeibkK6PHDpcQ2gf9fafjsn7
sWlKxQ61d/ZPiMAz90DCFsMA2kBysAeRTuwwvY/Tmmc3RMKyHgosQm0sr9E8WGkYGRLCUbF4CyHN
Hm4LUjq1/m373S8HwuOyhiwIQmP61zLK+XJgIjr6dZcD1rJQn8SoQdYP1PslFj0ApL92yO9QeYmp
Biv/6g+F8GmNR3C1+ZRB4Ey8NdKJ3Ma2lABi0KUT/KBzsN3UJKpBkHh9Vcu/lUv6TWSKpeng2XYk
i6NxpEYCfqMqAwkTooecXZ/7bDKAMbc4VpRcP8nq/ih85w1YOoj5mDqnURRDad5+ZiSi7dM0Fx0g
AoDP84fK0550lL1AD83JCPJPofEGqHYYXLnDBFFvujHrIE9YhCcgQv7MN6L+Nk5Sy9B5n3amd5IK
ydbwMBw4ar5PACBfnNhwMOO7u2j5GhNTbBy1QThTXNp4oheMyzMuUnXarsxa8dsneEvrZr47bk9K
jZMrrP+AnGCpJ9wdYeKaHwfAp67W5hvieN6cN7blgzycNxB8Hgd89m9nG2Ru0F6iR56QsH44QokM
QdXC0jBE33EAL2DJuuwAp8wjQAu2QWvdBFFi9bzJ3rkMB999fC1wFxMC+hLww7oUHVGD2S4atG1S
y8o6UBIsInRSvZdkQCBa1gWd/tZM4xaxJ8t/Z9M3OSEF7NbUCkibzJoE71TL8ve+fLuPDY81IFYf
fxD+DjiRjsszZzhG/jVzv4TMvaKrsfMkMyWJVhq2SwYlfW/7nDvavdI7JgjH9gs3ALe9slVVappY
dm60njVRxXEp2lGpEOdp8c3yBWpgxuL1jY1MrZTz7G2MVp+jSI9D6bf/Ea/GRs4w/q6YhhG+5MHt
auRb/f9bByH95BGG6zaCvLHR60PHPiI0GdJZdbhsV0U9a4VBCNyu6cfXAhH/daaHKPfif3oHzznQ
V6YWnIHISAnDT/ukqwyqg75K4Vcp3vtR/bfq/pUMu7QaL9YMn7qpqlcRFFgI0De0Qrd5EEUWcpW0
u1QVQWqca9fu2MQxX1Q+cwpymkknZ7w8kmyE32kXuLo7DRpBaT8Eh/TXyOBToNcqhsZdqi8o3JVx
ACqt1PLErdA1fLEa+OdCqv20onFrqPzk9ZIK56gPlXSU6d5fLoCJfPsR+Ca+sqIGTPynC3TCDsa8
u26zfAFwkDEDWPvRzpCFaHe1eQJMiewamSAYgeobdTlLzaB7xfyVKV82HCL/kSslfsvW36yxi5ak
Wmz/6da51KFf4aqb/rWYNXXMEbLf8wRr/i/lK0S1Gp++FKDSMbnPc2BC+pc/OIKcB6RfCpA/g6xT
c4x7P3Ns7sdaYOZ2A4OOFJewsIayljDG3LbgFRNLSJO1KH/0JmXLnqBTkqSLsCC2L4eFYCFH4Ble
RseSCVOaohY2Dq1l6G+KoFx32fAg/WfaLW95CQn4CASXBc2Duf2HDQfYlTJItnVIelleSnAefYwS
hdPxRq5pJOU7Wf3nHYQPcOfGv6/X164VXa/LqtVuh9ovfFIe2eGJfS2jnPRRFqsl4NewuH0bHgEF
PmfzrdnzTGTc1BbVd1AlniVo7IjOSE5vJeOCm2S0l3BT4I85sjbiqigcGPJODI/fqGW7j0lCce8t
0STrTzL5GE4/61mP6gXT4LNU91j1E5c+/gjMrYsrISmbEiyP4w9CQqu13/Mm1Gm5rde+nbWASMDr
lJbAHQc6fCGFcwOSTw2GzXkWIwjG2jymACU08RLSxwSrQM25jIZubhcU55ohJUhpqTuAWF12i5nR
Q6JSk2F9S2RP/HclM20KEdkljtYCCtpxkuNZs+KSx5uwJLvvVpPp4Fw5hxdk8suqLOGvkNGW8jsb
XcS/FLjTNsRkInF5Zo+ByjXSfR9S0eX09q7aKxiS85vS44b74b3vj5EWsei8nrysWsiH8cqE53mb
sf23uCZ5LCx/VeUDTqwC44HsnCS/SneknUhXHqIZeKms7qsWZAWC6M0MuVSAVpzVsXmCaRmfa3cV
TtE+ylAPGluTf0b7KtxKISRQsqAdawKeOX6yNRHxQf/+Sn2MuJgvwMtRuwb6kg6ISzrm+aoweuEm
7UICMqu8jreKMZmC/yVYhqKuy/UnbBJ3k+ouFOpyfvwAAz3XQJq54AIUJF8CGhmYZj5YrQBJZsdj
jZzuQEMwW10VEE91tLlqUH8m5QDePbdZSCTMWzRTloxe4fb4wpVd+NF/hWJcZ3crhySosO/wi9tu
AZ4MgEHOHYpslYftun4obU6bkhbTYKPvsHoaIJlzU5H50kLKbnwXH/gHIxpJG6EMsY5M8IxnA3mO
qOKCEIqjDbfWwuAmcJBNqT8//eC7tHVvtQiYpt0WGRHxZbwC8rMBpWhFx5qA45TUxdOmuJaWVNpn
+b8lpQbwTjcpWt1gvU6sSVDJANqgP9X6NwBu8QPgxYlSPF5CtT66PwWHUIe0fMUtbIfUTPxt6PYE
eESNUHW4dWwMm9e+jSTwURVj4TXZpJpWLnX2rsX6x5YRf9jRW/yy53G0zfbZ8i9FuP0/IbSqHjiA
p3zwSp3NmnbpznaalVOC8OQ1J/rRN49Xn4efpVugQG9sW+taZxZw578i2EEtdqOIj9jdqf280p9Z
t9n6wBhTjbLkbtzEo281ovPKKHfm/v0YIeOAnTpiwQ7IyPsi3eW1PqUDRfeRYJGbaNJ6a6PwNvUp
oWCcRnZ9Atcu5o5O3WfbYkD1eoZU0BooUByN04hzden3/yM6hL0Mi/a5t97rWflhMmYbVT+F/Hvp
bwNmocWQTM1yKwYks/UVvrcuhwz5ZRFnDefh04t0Ic+y2DDAeKCSiSjuwosWGV/j+Lfu0g3nu+Gg
byuOzmsR3DExI7IlTcPkVuv/+BRafxiBgpPg5Zm7oALOJHo+qn3APKNkMm95QqesVx2mVAzJOfmC
bo0MPL3P3qX2JAUNhXaiaB4hu1KSAwj/nKeS/K5UXRgHimLte9REnLZqYcdMme8n2BLkeUYRjtnw
CIcOsBanSDsZ8X/wqYAC2Mdkzt2Q0jip6jIXkuKY1GD8DUQHQm6DlBdV9X0pUk1EUDciD20OexhL
bJwmb5A0WOjo8FIcv1Hbonbp3zERmsvQiYpAQzSqKT+u4c9WJSVg1nMLdEo9ggjeV6cTUGynuAA+
bc3EFOzGuTgGhZ5Z/xG3JLI3gJvvqETnOjnw/JWdURkFXe9MibwwvfbbMMdyeYqz9gn5yu3fd7Vk
4GXO9z1yikhdI33AfivqZiQmjzjEkfwBg1nUb4U5tGJtAimVy9KNIq0fkS+YfT7cygQ1je0kONRF
Ses+z+A57ifL6SA2pjS12oKnmfgMuPdXf/42P0PvyuOfg4WGZC+4biG/OJc4MtMzwk8LcxSjQhna
QosamnpCapreFfmU4UAZS+MifX9SRMkUbtrknR9HdnNkYRa2ln5kWbcrv914VX6m2XpEBMYZTQjj
cv0iLSc3HHqSejnVVJmerk43xKot2wzyCnYJoQas27yJGIEelimxP5vtK22esVjyaSisRlvsVXNl
tjswECIbhKfeJ6eHcWDX9g1CeSN50sYVd7R5SxrBjIulZyHL+nnM1KPpiBteNxPVY2dyFRqRXNb6
TZBIFg3T3h7USZb9QmdnzT7Sj27uLsRXlE2xUymHVLvJ7RoZRJYnMkf2N4RhJnldkZIEv/RHatC4
py1OdEhhEcvlKrI2QimwlT/uBglNvleHdqf65cuA/0/S7phUC+PvC0zG0aOE3/tHzrcJK05d52jy
7xP6+PMPO70ko+/WibzQDLY8mvjiBiASxTPwgoTduEQ1fwUlyS53traAbVzKUAI9WBBY1rnX5C+5
dwvGEnm76N2UTWZd4qJ5UnQRnshOtfOmlyN4KBkMuUy2S7ndKvuN+CXzkJ2lVXZPaZD+4Yo7+DUv
E/gEp5vdwvwi3FcGHG9FhvsNJ4aZiTuZgq5yQboBkFBrsv/zRr40MfQEIUb9jrHoSbbGP922swq1
rXE7tPeLFOhIPMAmoh91LyyDEsjgj9aYepuMQ2UGGIfh3ycBCjyoRjOXuHq9NXcyZg7bv5R6wGpy
a6g2fWkaIHlnl+wzXUmNiJiRjKQSzM23f5x6+AdZ33y65ds/uO5XGUTNwxNB8VDKvFR7/TsLbEMU
VuaR5ToeNkTAnVi4ko7XTumzSWxix5ocBj7UUdOyKQUolK79b9c3pct/GqA7o8S0hLA5ud9NqHcU
qM6eug8AUXBc+GmDXeodODZWE+NyGzQeEWbhxeqoMG20x1u8MnVVwVupPye9inTg8iDAtWNA1Glt
irU7M/pnQ5TG98yEzD3YXCHF5tTjOtbpeZiWsmmRVp1G07atY7NXaWsipdJL3oy0S5BKEGQxSyg6
2IyijklhgXBqJyXCCJJj8dyF9MEKKeDjiYCy9NUDokBnTzReQeJUGzzaGsaElPs6AD5FkClhRBPE
QOa/LcvAu4RuSVYJO9STPvtC0hRMqAImFeDhPDBdHkKoYfewYJS8DJY2sJWRsZ6NkqXUlOM4lwfG
cyLas+4xd9q/W1mW7gKHr26zulX+Jtc1Eu9gqQNeedtPYOnW6p70BHtAMzLhwuiMZn5jEPYKSwII
KTTpCJbwgyjojWg3f75NWlJQiCLYJHgWtsqWpbpP8EVwqviGgQQomeJJSLWHr+sXK+ODiLvkU3Za
0MXkt/lBMYO+o7SDv8+xu7tTBZWwfzLvmFaDbEqcZY57B/3ECJFOK7d8+fF+0ctxr040VX8JV4OS
gfMFBb7TZy1KkFxFtndd6I1CcTEF0jpRnz5uvyJerXXLUlPF03GFoeb7/+3jWZINAxic9b/4f+0Q
nuhwSKmr1gCY0oDEtRp6MR+FuYrR5bKeG2u3/g6IiMA6MplSjyAPxEsN5mQEHeK+KgXRnMe8WEyz
K2PzYULxUJ//Jcf4Ux5aex9Q6ygcXpXmWlT1SBD/hL0ITweLUEzwvF3sJBUD4P593usb+SzzQBxY
5D9hWg78xURifEn+lmGerB4cRkb12OZsmuy72nf0UyoiZtahCbEhb6Ap5OFQ1WpmYIArZKPs8xkB
ruHfjDN6a0fTJSMA458GVGGzsQ1cCmjpQ13GniOimef7LmBwOFRlY+xnsLH5cKU5l85lKOCSfQWX
gNKKNut5YvFCRhTur3aJSCnS+nMVGlaDgPiybhFpf8M4P/X4rmmkssXZDIZpBQdqvqWkaL1DUbxr
x5tPZL9npr6WrCyVPq+JmddqOHLOPH3M2q3UHf9T51+3Mm9MdmiU120lkRKghNulDmgayTx3E1oE
/CCIR5UJTKqYyyIn7vOJL6eEm85Zs4VyYPDSMswgsTPvJJVazOo+n0c7JTz9JZ/0tEH/PeHlSgLL
znHg5sQMsbcr/lCSFcjwHSCZ+VQgm0W2nmXqLV6FPOs5wvN4/ntfGbKdU5EZpQA3Lag6uVqYKgyt
DPiFFPDmFbUwc2+FxUp6ZRIrbZI6pNqzDx5JPv+4Eub161tSN1B9dC5Bur4RYal17BKwpRMm70RJ
u8qJ2NWVgjr14GtlIQ1xPaiXd6cwavdRxhSMDUD2NMAOrxr2OoCa5NJY8xVNwrGk6fsMUsNour7U
aAXPdZ3PuCLqDDSqrf75HoMYeQHWiOunujpGccwP2IBfEC/kt3AFFstxx2VSLExUYwKzMQUIk34/
wOHWdQb3cCzPSbm3svVDSQ5Mo+Krq2JtBll3qi1RgRQCZlyi7xcDqNNqbT83rnZRNAMftQ7VS/R/
JWM9saipwBIWW0As1ZwiUELOuFWiiNO+5rpSBMKSpTf7bRtT8PZ3z+fFMpWtmt87TFN3wMquPZ8v
jXYPH12jqTyJzkuqJ03M3CC6sf7HVdhzHA+U0QnBTedujArIW+9cXUJG9hZng3t2DeXnY0DEV6rY
wEJM4Nm8XjL+h2aKPkWUxEYG9cUham8V49dvbW+6JJVKcRo7D4NfISwluwX58TeX+h+BGD2y6r9N
ZGdR3Bn/oWc6B8/hYd0PJNy8OL/DwI4TwX6u0qDvVT9+mCae+ENixK8KLAPBm1y/aJzVUo+F9RjG
bwSnUkFlWK92WivM1MK34AKgrOfFBBny8dZdlFEXq4Cck3S2lgqqx6/SDQe3YQ43IdEfAt48ahYI
jm4FiqWUg3GyS7TjboJTXe0UZBambF6SV1a2Z8vwcDBbqydl8bArlv48upl4ssHmMZ2wf1n2030x
WzvaJEZ9TWlGSmxZ3nZ9Zmckqmeeh2pLc4Sc7wOydYEZLVeQu7nkQh/5PLimg+BcVxCnHD/rEKhF
3HRe339/taLgeydaDdysAWReUx2Cj55Qe8tjBd4xyleyFBlj/pIj8Tk98laK7mQeiDLmqlMMY9hD
NaqhgBcB/72j52wQDkeiyovPhm0M+FISeeEXVN8uAaoT1tmaBjXHvIIahDKEWgC0b34cB1QQoO8E
dAOfoWGJz5iwq8TKT1jqgk3jV6Rkk8o9K2cZ6faVI3JVgJeYigDDlnhJR8Jv45VWHLTBQCBsKAKR
ts3SOr951puDxg+wqPCf27gJl3dsJnR+9PJlkpFcfCN5s+mHtYd1nLft9BqkqfqBFXCh8CZfiXEB
Hl9y3h6W8pKoL18bszYQ0/Kdz+Kq6oloERqpDJh7QBPACwMcJFMHv76WO43W5yaAVZK1+WEGOvKv
AP9MjA0KriscyyOApxD6gsm2aiIMXt8OTcoEUZswDo/K0plHgdiTHUzlhC2R6IrcAR5y+MrQL/4Q
UGMkYQnNxssvqF51Vd0EFYjhxqY3/rKQg64euwTx+1IvRlY3w+QLIefSSqTX5uw7Qeht5wxD2uBi
CyOISOYH51Tt4m3QEzhss564bCLZxmz5LfP0pfBwPbniRI9TPrees8v4Pjiq6gtIhDDqoBLhKLWu
+UpATlfeWrJo52IMjIRnumXLgdibotwu2EtuyYZIn2gHyGgNjXxuvO9843JipnUumO7S38ENv7ix
C14KzgK6WxyoJBKPqmPOQ3rjQLAr9YCbZj+513Ydf5slRwdn1+N70bJvE9bk8jwlfTCY5+SKiSQP
M9l/9hEWQnXL4Qs8JAmxxYQl7GNJ6K5UVks5ZOsigAdYORqJQNvcH0SU5gh3hOmwEx14rJ3jDuGB
Gh9RfINuz4t2CBedu1L6pNpWeEg8mI6XuFg9nE1WdSU2DIKcMyidYV1l4DVex1dCoeV5sxNTUQIA
QJADGt9Q9EfMienbSLyUAe9Dz6Vs8VcMZbZ1hFKufqJqy79TGd+0CeDMqreXzqJS/8T7wIHRO+8o
ekRLb3d6HOyNTv4IPebHaB6j4lu2j+NKnYx47GPPGyTw4HkIH+BLeF/oMiQedDoZ1QAvRH077gVA
n/+BeSjJLG9uYbVtgR23CXYGQHTK03Axw4K5FFWEY2f4RFEqUqeUFyipr5DCts38eXLXlCzPhcod
Tre5umr6gnM5llH6J1dkOx+pclIK7xujzVVdSFByllfbvD3wLEttYqqNSMjSg/yi+BGmScgxmR8u
ZROqcsdMlxMPQUSqZwuIILOBN6dALkAN50RQvHBn2cMCtN3Z9nsuQLSXfejF3zFIEg9UQ/9eHznF
HvxbJiv8Wvo/xz8rpPcP8F4lo7w2ahTfHoelBjWB0V4o0p/mSCaJFo2rebGvkjcjjdFRMUuux2DI
u86uqpoJycf8xHgrBNtVDMaw7ITg+TfE8yTv7nhgTYxc5ZAN/mY9F/oGACjcd/VnARnbVPe2ahge
CYDjae/ssLEHsOKdCCp12XaffE/+sFQSEZ/ibhFPBsgr6yzqAd6iJcWfE2OGf9hjBkCAc9fD3ftO
eEGV04SSRoFBz5rxxO0FCnSmf7JVP1bTXQVTiKwQqcw8l8f0KW9jymR8fWTanAq/kK0d/Z+iD01z
akHK+ICJjKgd5Sd/mCxhYDowXk9oM2/uvW3Ci7FptgeyyHBfEGrXQuszgcdYXD04TASZ/3kc5eW7
7JNjBInSf2kJa3yNcaKIDAvOLLSZ8Ag/r7v2nSz7jtck5NJOgRGm3lxn5r7tIaiqXB8bv7IVNgEA
JJOIj5LzS5WBVheB9589/K1JAq6EqJdBKKAfPzbErEUVADOxn/qbR3uHPsBS1KRqGfeRsiN9p+Ze
64USPuJshlUcxiAmiSMDn6PKVttwRRWAdGYTzM9bHatpn08cWwTm+w+Cby3f8wFTJcgJIpwta4VB
NRUYCel2ZMq+9P1G6BF9SHpgJa3iN7y8tXp5busA3zMhJaDjvqqVO5XO4t4s2XhYgL/xHDL0Kr7y
63ZX28g3MNr3V+UtocwJBtdi+DvU7B+Cy3wEGN8T6hPl/bjvLmaAdrgWK/Aw1g9keo8Gkilyt6OJ
P54MhHRNAM6JhchMI0AfEEr8JxRATnCCXia9FwNYKFzzPJxGHOiinqjPB0vhMKyuoHLXN++qagfg
4aiAF1nS97siqlN8Fie2BKHokIwGLr9z7nWgZUfuf0pG3BJakvmEP9Ryd41Y5t/kTiMzlqJZ319W
5ZyDst/A6BolV4l5ngHDqdStDhOihHU7koWokGJcSGL6GLsI2/+FgOCcy5i2XpRpcPJ67ObBT5Jj
TnLNBqzXDmD8fd9WQgfh9W0wrl5P6IA01jX2E8gOugbIy3YtTmh7HuRPLvIVQnFL61SyJ/HAosUZ
4QCwf7PKhN2LKrKYVQqBWgDCDKh68Lg8vXc5o+tDvhAX2myv16YOEx4t1lwhvpuRTsFldpHhLMCq
ZZcKZLolbseU+oV0PpziZm/MPi46J8nFocp4uxdfWtSdjGLya2VrbhjSAPZiOPAAYzrh1UBUMmHW
UfIyAx0kcXHMjV7BcN08ZHwlB1dPLdNZrXLHJcRGUCCDxxnHhC392XnohASf92+yf6TfVWX3dvOn
rs0VDO7SorVc5z74EeARi1bDkD0oNiA5qYPzxxjYCsSi/005Utf2IVAkiSBdgPBM46ByiNDd6AjV
eX4INH/xkQdmounoYEdWfnqRHlh7oPH+w9LBRBEL7fl7QR5SyrA1OJnob00+oHUB7Q3vi1/xxXcH
BPer1cBo3bFsKi2fvA/CmxEGVTV3GtcqXnxji7EKduJCpMF9I/x4z6bQj+JSwenI2+w4uWUM6maX
uV6TPbosgZg3bnR/NshwLgtarjXA6RxGvhncOh1Z18noLGg9JlXg3X40ltghIq+MfhMwjiNkzztg
oICA4uh5ldYupjT9iTcWEDD96DpRWYgit9JimaTT6J0Rq+0JltV2pVvjl1EOltdurvH7Sdo4s7Kk
QPrYm92j50nR3af3xm/+5MKzo+GW9XuiTf/7r+CAgzzfE9C8W4h3CD4Jj1k8kD0GglMiKV9s8c2J
etBUpSXc/R7uKQeNcJmHVvOsthoTyqK7VToetC9Yjr+lLAFO+1HYLfjO5O7thDoQYtkQ0n1/4a0m
lCMYBLXiaI0rUlFK4Odo5/J7ufYWZ3pcUBCd8QtmX6S+dPBLhgKV9of8fFU70n596tYgF9y7VuJ4
Kk+KlYYaTqxgpj5zX+eQM3b55cTQCjQ7bNDpuKyn8pp7w5BGq60K5869mkGw1HWikPMssqaT3XRp
TpeOMK7nL8XCWRUoIs1blwhJY5OwcNfd2dE5MNoJGH+FcK7KGb2DKOCEhqZ/ef8N/txc5Kfi+RLn
xq8UljPeCN4rkGyBdxVT8HS9oI4BIXmrlFU+9GdyWbB4W1GWBwlxAuHQ2Odu1ImezDW329z1r+Fc
rAxC5soVRBchSDk5R1CtVAlfIhapwH2NLDJ7QFxCELkkZsp4p44HAk7nk5lvqipUdZ7PtfuudA70
J2FuXjoiLmWM8dfJZ2B5pgigbTKtPO5OAsfLVvgiMNuIEZJ3ccDsQha7oP44Vq0uiuSehy4neBY1
uPhmGoM0ovdL9ovs2StzQEVvmt6vLG1hYbnZhSUf2xFgLjsfyGwC4Y0QDL64w3HfWarT3MnftA4C
1dWdvZyZzWgAzvPqNprYtye0DesMxXOoAKI8yc6HW/dT7TL61/bKDgenuzQQ5HTCad6XpCryDGP2
dRsUqfTZdTqE83X4q7wLsJFD4y2cJqwK5GUHaJpWgZ99ad/UCpnRwVAsfnCNAlaa/sMGFxRilwJJ
DD4HMVNc7SpBgCS3ls8w8XUlw+cytqzwp08SpDhTs/ufTzj6aiYe1sW4EytYDKwWO3k5muLlqeD/
hqRShT3IWXH37eO+00SMz1GSek3mth1IwgvH/12HBUkOQtgEiVWJRNBGDpVYvjSMxDnjlyEmvynP
pRvlx+2KxThjU3fIJWMfEPS43pKD3EvvORa0+VDxLWo7Ao1QlygG7mgP46kkMHGl07sVe8TXbv0g
1s4XFzF1mnFu/EyD1TN9p8SP0AdYGPyBGMuA5kHyLrZwFAJBYtyQUFVgSurR1TJGbaiKyCWUP/zu
pxYg7RHWVAlm/EVY2tvuxqbPIMehlnFYfqX6JsWl1TPhBnFYnts/kwOqTaHcMqtr/z9P5jgrHLjb
rLKQPpiDu7lGPCFE/rpfnOxN5N5FjfRsSsJEVfFNmhkPNoQzYv1a4fJUJy5OyGe0no8ToclE0EPf
o1fmaX0a/cIVGm/t3zo5eBBQoqw0zFfYM6VwgUcSRs0cVZKLX+U0878BP8XZGzO8nSzLcx0iSAA4
p8FTEmpfjds57iOiUGGWvJTZu0E6zS65AoBqq6O4dMsgyAwA4wY2Vilj3XtO/kryjS8b+2snowJn
JBvapKWmtjYxaaG0XbU8tv9/Mc4bl6oVRVdCycaurMpk0BTbiRZ9iPD1rM/XcxWtQmfUjvhwr0iz
hnWyxvDKpq5Y2A/5HH8XeopYKBkkFVpsmCs2p/vM6kUI8IAQAP8LA8vOqH7lNsy66QPovQt/1lsX
uJdYh4Ee6pb/MoLGw80XIeJrJMawAjlwP5S8fAJogGXAmw1vdiNhpIgww6ueJWNGIHz0MVMVvfik
Uzw6WAkmP+mi+mxrYwRz6UINVPYTHPhrF/WRYQQ8XJVsi+nz14GgrQ4aUW/iroIjeXRDvMj0qU5b
BnVqfmwy0UqxeMyfdN7RLExFBpeu8QcpjIrfzpxo72N4R1V/vXzQ4x7kE/IaWiYx27GZNfzPv4c+
ZUPvQZr6AkA3jGNQLX9XHvfda8SZXWaRgJrNmVwVggRD30QkcIG7Eh3uZA4o0uYLYXL0BDGbgWep
zFar3oW+Vx1tF5nHfVeelcgEpemesNSGlQ7P5scW7fej9YJmDHhciq+8yeJxz62r48vzem3xZK3S
o/YFjDLMAdv8iv2FapqKv+dWTcb7y056jHI/8GkwP/o0Pa/ZMfJIRlh8LH70hN6uld3pYYESK1qW
wA8Ijzlsri1CtqjsAZMBzOFfC7mCbLc+sHUOGC/bMZeOTQdZ1N25q7pIeNL2Wzou5RTM5MZnSAq8
nrvtxpkz1JIFMU0Z787tBGF9tYAwAzVWj0wePMZGJfanbmgbZ6gV2lYTk1Kw0RvfrC4H3KtHRb7D
L9ZFnWZo/zgvhtthIDOwQdMtZrnVMy6KRPblZzbL77nVpDAJakhir9Ts/25DPSuzGrcOe0RoFIfG
k/Pq5WJmHKxUjw38pwN0isyjRpcDKRqIP5FymzJUORd9vu2KjT4PEmwl/LLS09GeHxLrIkf9kNYD
d5mjzld6CobJKOJAwk7C+/s27GzhrvwKxFArdEwZdloTIzevgjRqs1S5JCruWStoWBzLNPyvoTFf
a2aAsqxSb5FigZGS6Ov1rhRHmgd+UEIZIz+xmMqOGjhZaXRh0SidhAXTyVQqebK79aaZDP7shOF3
US8OzM5zOaWvuehtfdZz8iFRk7BkQPbYJGr2o7a/em5c30KhnTVaqZoNZkkTzd4wlYiET5L2N+QC
uoGeLgrPidvmwrft1GK5m1fVHIMKtecRjGNiGoj3Yqvcs2tmyDeMPEkqGH0st2bl9MRddEW8k8Tb
v550ALOfr8V7QR6528qgG5TbGQgprUTYG1F4gKCcrlFflBmD4sGR8sRJoGRXqeJF+FZgzq71IjhT
xsT2Gka6GGb79YdiT+NXJW691aTJ1pbfBBuFOR3qCD/cicVVIfNgwMt1NuL1WGBACGM6sXNOMrcT
yryXWqVYaPl293YRVgbe27Un5YmS1crt/w8Qm/DY5u+NtrhctuUpuuz3a4xX3VNRV3iD1Sy5jrkO
nXYzj3Rv6X3IkgfNVbecMWcsLLcsMu0pJXAgfHfq8XIyrJvJKAnav1K6dBEeci6pi92kAYkALU2a
MaXz0/gGESwtJDhGgmg5EU0MwcUKdapyAh/curUowR6fERkPbRQi0bNouPTViTSmYbu6dKXoTaf6
3jNeMtHUb2txopo3lPUP4jKSuucuze4qq9FZfkUWCbOwtsyK2olM1M/FN+LtUUc8jKC2asz3tX0b
uti65rXUDmFz/MSZGYNJCeUMphKSuHOVD1vFzN47ZgSnNUTw8VktzHrsJS4CXw9LBHm++zprpk48
Vf6pScochH73Rw12yVPRWmzs7acj6F2eEExVVgcC2YM+B/LQJpqTcWWRs74WbDKkiAzfQLR6xu9p
LQ09hkzhw4bv9vwkJitMLfekPo+uVudL8jJz3IqNGJ52YBBZ+2JQPnASJSBQNhv1MPhO58wlcRy5
GVecqFXSwxumZQ2QwnZ9EZaC+VlYX9uPuvPBK2jSiree+tOlu7LU/xZii3Byhj8halXhT4dOmXfS
EVBgkXs12hniDtONYRNnZJS7PjfMC/9sL6LXAvR/2rTDmn/2xYYO02zb9b0xOR+hIThWpz927e/u
7q6t1qMa1NAXbkE1TK5oLS8a/t2crSmcijcaMGznQLcxRHFyEi4IpR4VC3hnuI4d2IcAHkmHkx5K
PXsx7RUCMWgL0O4Pb528I7Dc75M8L6k3YwRbbn5Vv+rtPhZFx8GXr8REAHTXetKsh3gga2PkfsfT
UmoUDn8wBQn1QH618P5tMgeiR0A0suGhRi05ogvbGIdyXyHf88h3uHCrPj7hTxJaJ4urKbvJeJzH
PXmgJElQlRagevhdOkCZJr4wrmuCB9qNKYrJi+Oc3VXYGXvni8niMMyu+xWlvRhuCseFcY6yQbsT
In+k6NGS1Nvd662IFmzMTr9EDgu5sL5TwLxSuH10p/9PuW8oIaZ3+KODde1ekEHMPn+zRfEUA7ug
dVSEyAkaNL+u391Tu2G1b5O0mnq2Fi9re9uXvz3/DbnSmlYu7r6htrr6ogMuHdSInNLj7y1eNXXe
Uy0RZjJzFCK6wBYBU85thF5zYotYCSAtlXjLQei7uz6GxXgmHPQFcPoaghULb6GXNln70yujtuYk
AEOwrvgnrEFNQywcksHiirMqhwDxZSMh33l9nc/tJSFPDtkYAiEqSXCFQolHbbOsLWgU0MECrW1V
DqjCktMutJAUNYf6cRlxFrQYJ96oajdCGi5ASLVqiSaLAOdCRTBEAdj+HrgHMRlbzvdr3OXnF65b
aok4oALJiOK4xXxVA/C9ERjnngpU6r6j72R3d2m40W7bcuMpzRyX1RpbUdjncxW9fm4bORlz+RXy
Q+anNBTQfA30sUcWZTx+0hF5rHCR/rgZowYCxfcjm8iiVEDJ0nl//KgPue68MnM3Q0Cpl4AabkGH
34Jw7QR3qydTAWlSSjfrIR1bxPINiEOB8MF4hc6htxYfRThlJctH4tjMVutQroI6AsS6iKeRQG8w
oAFnq1CIb+/10VYmkPMkXcSr54YBt3IQJjhvm/21r7w5mxfwGO+SkLaPdcxRJwVY5dtLtoU+frhz
nQj9nbZfuQT3vM5Gp3E6rh/RRyVS3YHrP7C8hEFXc0/P1uT/ik4p1ooqitbOjy86ntO5HbAJdMeq
+HSB/AvqA2BIxgbVyTo9U1JwA8mAv7ePTooB9mCkfBWuSWhEyA/LBgMcxQ/afNkS54kZotWOLwCQ
j7W+fE9UIZO1ffD2Y4cS2sc2Xk2UrBiuNXzqLSuIzah0T8cDEpaDkCm8PoT9ALGIwVX/SVXq69lo
Kxd7asWwvIQE+UgLvCwmgd03R170DKvGBtGebATDtmqVdLqHVYM8F8Enijw4RSU9mMqiPLf3XZ5+
WBoMwf0ncuzRs/zYvVKu9Y4D6WHOM2SJYgHx5W3VttfRl3imM9owI3U0baWO3UjQgmopEDiZG5XT
lpxn3VyAccF0RJWXDT8Q+ggi8tckzZiev9PZDGjgyON36u4orIOcR61I6UAOawlIxZOCk21vhKVp
MLnSpx0QU14N2kCychDOn0gOE4s8mApbfgWcZkfNQ9Ten2GO97PcbzL321fgeh+oT7kdTiBceIQp
gh/A9p20QEM5gtKVRrDZKh7ewO9Zj0bi3tTppk/cWkJvHOHqbuj4S5lzMddnDxYywdQ1mh0S+4Cj
ghskRBsvhKL+1PHrB5CVAMzOpcWuATwoKgbHKyhgSfbu2mFAyaXfVAzCxlOx9R+SU6HIBj7onlB0
7RoPDNOX92/AmzH4iUsdjIdo2TVqsJkGNcICy9QtZnNG85NjjTWSZyc3BU4qN7A3oxoCYPAbSH1q
LnyUiOJKWaTHF8GJ9ZfqSrYyf9xT8l4Q4ZSDGGU0s5JjhAIrPbD6pK+AMQf1HFC3NBMMQQQ1t9P/
JdaJmGQRwxKsWj987i8wc6a0s7eGJh/MAnWUXG9vDzSxj0tWnO+KU4k1oxArXComkVZMxdyct7Dt
i2L3/Dt5FhWJF9r1PRgSooE+U/lhkrHq7pquAoYp0jp33dj99YT6c/6CwK3i4oaTiipS5tw/R2ns
2iMU2Y5VafYgkAEc7lBeN9tPwuiAX5Dkvxg3v3wrj1m/LoK2L4C6pR/qI2I1wjZ4dy6gpT7MJ0MJ
SrnQMcUjW83dW0+apuqhdekhUlzyZfjTBJ516tldQxLP06rAX2Pi5b5X+Lrtxs9KzkEVVB3OdaT3
FbhY09ZzvvNKshhPipPOSPqLQNBxPWRmQyL/LJu40c942v4UDTXltrhbgl0W+PsUrvQzqqAh5SqA
GEQgmwuyUKnEvlzCeKCnkZoo7znnw1QIzHFCPyxVZsSrYTah6TCWelSraYp4aVuzR9S/11O7lBWA
QvATcaMALgMWixtFXCjdb2UW8a+S6JjvJIMCnCG4/lNxxGd1yHjcaFoop+moJAsNJvjh7Dmhf7S3
XLTO3LP8s3WoJtEFefnNagiv1HBpDA7FCdiVRr/NCQ6ZnUHLSAbD9fuZ+FTaCIzPVwDKMr7S7lkI
wmyVh0UKFyoMxD/u++GwzqKJIVI0nmCUY7uz0ycQuVciAl7ghJMAEIc5r1gpFxOXUpJbV/Z9FUtE
i4lAH5cCdlxm5CGmOpdqjq49R/YSBs9bdlwnJs8G2w74Ba3G8KJ9TsXQQ+3Huzs0meR+/ycF6XJm
o8meWgLu/g48oD4yQZzpGQCwMAOJRZz76KxQZ+PQh3qj5NX9X5288rPSBo8NrOWtwzPfSOkhY1xJ
kiUrZL7BS/linJO5w39FkKfDIJW33twwWtZ3Ns+btt8YyU50UlxNplYeOzAh3oGekLfFFQ78gdYn
H5JyEypLHN8BuZZ4bTXZ/J/lfQfR6BFThOuu6ONnULiBoxN4J5StsECG067qpwNNP0e5RmryjTxt
WDHfprlg6rgGGWuDd3eG/qhkdhDilvgHlM0pfL5xKku6bWMz2LO0RS1djsDxFPlDtepjAXWtvtnK
SoHqa9c2sv9nVW7IiyTSO6a/ZAxhJTgJAF2X6DPZ+AQoMO6OONYS1AIblnamvQUSVs9JFFe96cvK
q3eDPvPBnNDHVnIvwW8ik87bNWbQUKDFGiUostJsqvkoVsqKIv0Xt73EbJuu6uFDJRuXq8LXrwRO
BL/dRg8NvxBMfgDOp0Ol778G+UpowzdNtnxAaM/7lVmCCo0YFVXaZsPhsL/1jNfLySNX4bcc/Tr6
fxBoToe61no1pqXRrPfzFOR0JSlC+1GPi4S95/POmlQ5HsRiT2HPpmvfXswR5wBhwQQr7mulXdK7
AGNQpG7G3Km8cfk6eOqQJ1WSqZ3HhZDa/3ExSM1sIYXd5sCijwaeiMwk/82NuVH0S7tfS42MqxNZ
LRoaLofFuhn0OfYqUelsiQtuL2rFGnql72TctdbquKNjMTOpmq//5h2Kkkgj+c8J9fmXr7PqcdtH
at5twwg1QhwAvDAakCYRxLpHzl7gzVhYKxbeVNsz+hIExLkMKtSvTH8T0b+TdjDbwhiveg9QTyOl
zx58cRxqxOJRgGitCFTMca1fx/f9Nl5JGklG9VLz5UKU1ohLgAxOk0d66G5K1hJyzKy3C2JF4STf
z/E0uxx8CoN50jiBP8tKeSjuAiew08uDcG9H+IFei7XxxwHQ7v7YzFCtfzCwteMN4DGWPpL4ttYk
xn2NB726aVhqm0uAruY24jrQt5bbnVNfX9A7Nj9cJy471kI+wHaLVXjBca3Iv8bZAgoaf75wP7WA
6/KX2WWwe0yAm8/OTvq0cTYBy0TFonHAxqrzsR1/VhljrJu6uWureEXkom57qkMeEWb/GXYVUEvs
QfwHayS7oJOS8CgUyad2JdwAt6+BQ/zI15XqebxFuR0ZZfdKQwUhuvWqNNfUaafEZaNwO6Fbltej
9wpnfddOinejs8UWfO2lVk3g3dPWhV2xJtytshx1Hl+UYm+kE2R7rby2c4bUaZKLo/+9LsCbe/GP
dY1+lLPRfZ9Y7SIscEyu2Bre4LcZvfVycRmz7IzW6LlvM0Za5u9Ajds+RYfZmpej5gakP2YJsK5T
7G4Z1YbKgDsxyKmrIZ5Pyeze8crjGDJNLWc82tNq1zymN299HZW7rYH2HRBhyG3QtmzuUtyayUf6
gppWhc2QcGpvrlBFZZEFtK9wG5I/tvvDkbOXSeAQ3zM2qg2kWoBr7JwDyv4w+BOYRUgW33dOyyQo
WuPM7RYkTBoX9aREaZhANYLbZ3DQnCykDvW6yBsdDRVzOpsBvSbSgpSqcUc/ZbwQu0Q4wfhE24yM
mR9DiCBPgyE4TPDJ2cVVyyftkwdH4ccrXhmzOeBpZ8+79i4EA8XzUzxLulZDYC5ZwEVU7CdU67lH
NsaVQGg/wlzNLIOSpDr57xsxPSyEp8G6KWq/73q7q2TO5BhjbtT3WWnpMg6bqMiRjEpHPnOyE7T2
GdON1cCEFKVvhLRoolUirovOCP2mMJIkb6T8JmLTh41T8aIXL/UjxUmCdOXxr/0+kb4pUTl9UMRA
+IuUY1Y4EAa732tEAej3Vsuu70I+SEptcLro1fc/t05C+gtVUljmR0wOo8H46gDJv2tDseuohgiw
f1qJ6KRrscTwxW67v7wjXVrfOciYoXrkxanVK5Yuhk+GZO5ecVcTryCGhYEobLvrUUIf/vmudk2j
Vk9OLxwNY30/s3Yw1+I3wGCNd3t72R/8rfA51qbnRKWBS12r21iBtA7t1uNnnZj9LF1rf+yP/aXB
VBfwmwcjJl6/rCONsMrlpjCagNUcfOjjRz6eO0RBCfdTHi9FgRdeWXPD0wftYErV8KK1gHYKFw8J
VmsFMzPDuwanIz+6xXGV8zbpxUHXyAD5L++Lv4WXF5PnhmSU10cupE6HshE06WPlov4p9MLgsoqF
P7sXf+LwwVyOx5Wk8MmO9jouzLfJ4YoIlqGcwI2uelvX5gjhYElxF8BfjH+U6OAOzU6LW/ag01UC
XEbkJn0twXdiAzAFUBVoRWpqDFbpyblNEKtWb4NL3IA5Feym401ropebk8/Otjtd7QmD8hLZRgtE
y4WqVLGXUn8ynLOojA5kz3NH0toTTz03bmKSxLZyXKEUFeETa3GrgCs//digmPVrMyIhItdT9etu
Pt4uO8h16duQn2/VuhZYJTwziBIFqiWOVwZGHOuT1wf9SVNbl+EhF39Y1+EaUa/oFATrVpve1BTA
yd0mvrz+kJZWDlmZNxS+YsTkmOuL8+7beIhK+C/6DiKzU9hFhycptErPylyuRKhYKDsljyMCLbyu
e05Yg4u4Ao023WY0xRT8yf5gC2DE7d+bUQNjf0w09k1p6wxaN4fV1KbzrIkjQIG98GUoi5QbnQ7p
6OJRphvYj+QfY4gbByBlg4vikJs2q0kuZovQFUQvsIEU3AB5AgN01IhlcCXYTxnsP96Ctkuip3vI
aZ6UTW1xrwXzQMnqCtAlCjdK/roEB2AXPP/XscSykHdzzlYKGdYpnbTCeousy6ZCiISBAsRLRWm4
JzBjkBKbtiFhQhe8f12vXeg0gqaRHMnJOPgDBhOrCIOoCuoI2dK5jrNSpAWaSqrMP20YewpubKAX
4mEbTTC2WT3LBKAMf9/w2XjfiAAuKSjkeoZ+/L3eeEd1Moqj0eck4wgfSE272a6RL+6l0XhQmCu8
Gl0NXcvSDjb4XVnCI1xLQmIOYhzmudMAEn0+a2RKnh+2vYbfHL4WHRMmofqbyKz70Zhy+fmMZuQh
yjAH9Z76dxhqZyjbsOw5yLDI8WgoHr+BlRkUHs1004GWmec19kJMhh1ZEQ22iUKelgAQdUxWDCc4
Tj9fqByGI0Djy5SxdYJ/A5HXANFoua51u8utG1ksylnbdwL6o1Uqlpe1zruM6yfgLAOf76T7Dz2V
vFPb9O12qTDUBVNPjLLE0tsXcS9Ni+LA9jdvaTdUJ8mk6DK0iVPUu7iCuUL80XH7YBfzmMcX0On+
e6RnEQw/VkOGm3WaNpJuQ5W6BHPEZt5i4+CmuxO8E7LN5TWgbLJnTBUH+P3V8p2yF1SHzHEduZas
DZnxGzBtb3LE9lcGz8B8GD+X320nxXHfq91y7o7+bpCCeBSNMa3BE/xd2B/PF+DrjBl0CYJ7SxDd
hqXtt4jZsWT2+Fdhh/ejKtv69HMBmpgd30BGu7Aevw135emsC4Ax9DE7TmX1RgLaI9guyGiJtSu8
6gA4ikSCfAGE9rtRw+MXSCa0w3HcBWydFFA2K3LbZ8qjaI6LMIRHehdp1cN+plX78zyUn96eJv0K
Qh0If3f6pxhPB/JrZDpZ0T5WzCzOrWmxPz4SsL1xtRhBASr42NizWqNAP92Gu2oOb9IDYcEQ/NUw
qqY8tR4gBiKumO3algrTawOO4/Cl6Ermwxsj6UQW4eF48Otq4fwliNH/Bf1C/z922LcPPPDk6iJE
TVFwrjuFtHNsFwfQt07RuaEB5RwhlIohmlGCq3fCCLoSFykmznqITEJq+TeHqZmqjaocl36sxNqQ
+XtsFt7JjhAQ6Oka+qd3bE4hacuF4xNib0uWb3dUTVH8YsvuB3WrZcYmYI+JTD9rdvRXIgr+qStm
Dh9Oo3lxoOZWOyL+lmd/UgHFQVFiJ4Xt9TDDbmnBUvVZhGz3D7qQQhVWOkB3lZsDVsCRiHMEDe2k
SyLBDiYOZielSd9khyxSkrQ2Q7NdR/ln8fYW7J8VYfstS2V04OA05ieIjBx6P3LCH+kVut6b4uQq
oNTRtKtECLoTfG9ntJk+3nvKPv8ja8KOrwj+v6BEtURMDq71/Bwr0T1outoMU/twaYat7lLMl2kc
rU0utzFR0fx1H42J75k5+Lxiv3aZZ7vLPy1FvQsma9kWdq/IWdkJ1Co+TC3dVDJlkzo2njZsQBSq
LZj8k9DYe55Hpa9m3AFsfxp3RmMUjQzyeDxFcCIjN6Oj4rQeIOb40jRWtsEFFrKRmTLhNP5I1K+N
OlsVpoU6YaJoD8vd7xwHtR1y4+skKenyHu1px7USSU0nw8IDrbHLNaL35RCCgYKLnVWsvTQwKBlA
wEeHDd08sc7bG7sudp3DDwblhQRKJfu+QfV3FLC4YE/R0iyYgSvBFWxzPhV9pTJ0CCnCy7OMyeBe
g7GKR8pULm5i+QmQF20E0WfkX3t7unSI2KDIzyhSBtXamZL6g8MlcFLbtzNuqMtNed5Qowi7U+hZ
yWncWVH2XL/sLWeGdXc883sy6G/I+FHwSX1CgTtpL08LLAoFdRxyBYbUM0z+dj5IuHtPrW9GDHBm
s/hX3uKxB1FEH4dg8NSBPnx3IHD9rYxxg6JjCzrgeaNX3eGW8YOcpXXBK8k24wpnxPzmewdbQcbo
iXWHai5/V/NzoKQoqVo7il6pvZIXhZNrtjvFe1+u+k2uBUXz6D86xnnwOlLTwhV3egJHIBCz3iKe
uImXus5xV+z0SN4xdisi2D2O4rCcwqpimnXqldTAkNY/jyTpL53xjg+F1kZ8eTlQdsA2wcXfg6cS
nXQ3SaNdeodVLEGa1OoegXDin+IaDgbZrU280VUtyNIfV93LSfl8fmGD6oyXuGK9W0UnIXnbz8li
KKwPsuMx4WZQZBO0OrABRpYXpgnq16bc1kCC9qLYezjlu5AfpKXgnZ3wVneD+KNwoP+o9AiW/gHR
QujvP2k1dtpTnmr/FTlLqi33uAinxPHlvrZ+2DdmFUjSrkDgfTsLs/LvqLtqYoLM1R93pJi559EV
AGLKOdKABrQp3WpFidUsewG3R9H1ffH3QbHV9prTFaXz9Mm+vVoBcKXD5gv5W2j0oX8EzYbqIMhm
cyxClSMG2mfwyngRamADJcrvqf/7gK6Cb1Ii9/QJYGxty9+u1FWJZxmFb0DslJF7hII/ZuJfC0fm
KMwOsNTJjSqkociEhv3CaPK/vrKcTRRUtx1RymbiMIpaAUmNL3lWYYpmHCAHCCqPtAkuQBPUh3cs
HPlv291eNAgZKuSWHC+NaIQBfxdtHIREVTfYXB9HxTNoTzmznxzAEtM/jHgKk756xd8UcuwAPmqz
Q9HxyQygHfRhvXFRpwXqdj1rachhaQN2PbibGDEznJeuHC20ooOPISEZITwrJ8vPIE0rovHsdUGh
5GE2JpPFyz0bM2tqOFJp9Grr3yqq60mFaopyXVocD7JlWfJNbScLUZM5BDNbCdRebnb98NSUaQIP
rt0DHER3Bv4hRiKtH25sbRRlsKJugxlzPjbM/THhQoVoaRJdfvx7meGl/9qQQV9bZvRBXWBjma0x
jgtUo0wYF0oZz+de0UsAec5BUfSOpgmHgfHGDwP3jFmgfF2mnT2zeNwuyVNL/mFK2AsN8WvLRnt2
emCaYpZVyQJDFnWMeUFSUEI5j/Rh+8Rlk0hW6eXlmQkMMEMWT1sffA3A6adVkegBr9ktUUrfiUTR
CI/tTEYv4FE1a+ZxZck2Ef3It3DLYzLM2h1cNUhpi4HUIGOBCv9uPBLlx86+IseOgYYZ8JVI3i1Z
+39yAQPfPC7+lth9yZYExYkiz6zmOxtSABD7yOiImBVDBR+gbFAZgj7FF1CuGxHgdBMLk0GxHNFe
jL6T7DdN1KCL87BdN2+AgymtIOByoEUaNldJf84WJ34lOgX1nRW1Lw8cHPkgHmrnJUPuwZsyAF/O
uSFCL7KgFJgEPzZi9IMSbNRk9amzNHh6V6lp0Q9J+iGQ/7KR37y0e/ayAypNO/cdaIO+PEb99EnJ
kvP4ghjavUQnMCbMFkueOGG9a0yUkmcj+W4/Gp/fA1DhnMWOR3xGHYbbk34QR1pJ08DfHiActYRZ
K99DTb5MoI8HJjBN86GKriiuAWnRO2YsR31iiCh1gp/14Hy1WXuM7EMqZ4BdvlwEraEpWT+2/rAS
F8VFUE+AzDATubp/JY9jioHHm/9djep7BDw3ZOAKIgC5txZZkFchR7mJX1Kh3twWmjM/f5ua73mP
g0nNLdhSLb6jfIEUMv+pIGokw3RQwJmbHsYbPXD6vJ+keHU4W7H/qgFm8wVIxE0vDE22pqCtHpVs
b6LiwftOqSuAZfv7UJi+Bov6hkU00rKLex5hpzPxWaH9TzpLjZtZzqKjRTxHiTRXZe0K6aelohi/
9FR4TJVe67WQIKjorZv/ppa0Nen0/0Ms3IC0YjPmVHxyqMuP0WcsNn7flPEFuzdvDWziio9NBH1s
+tR+C+i92yqyG0N2HXa+LaypUrPLmxBLf7vyRPfvA+zJ0xfS8cCTVAINyY3WIvF5jJ/i5Gu6haec
i0WUSqOQ5DeUK2XnnYGrz94SybDbfgcSGAAtCgOzKWXhMNQaposkTKQDOImudGcgvbawkMDpkzB4
17xC+wADjN1NODhC1GRyzWCSjoCKc7VlWI68feoh7Qzwl4PnhT/SyT1YjtV/8Zit7s4LPe2ZnQFC
Y98BjLTUAaHCetXbZSONxEPLryVGYkYTdm88TvMQ2qIW90jXZF/gophAsbdHWA1f6pVGp9f21AH6
0GpkGwinFejMJWd8TFxXsoHWrKqTZMID+UQaB7kUpl4ir3RR5Qsu4+Tx4c3uKNr5NrrEu1AUelGh
6mUplTfoyrTzfrPAUHecUEcO+ywwP2QEWQKaKalNy5wswwEFNyTgsnJtIBFIXOi36pWwQTa5xQMF
mA1FaYFz9GoQzGSGRdiejuloaJg9YW1EcdMBinVp9kiWypiGeYSm8grTISd3d906GPIYmxlZpYKI
HAReeEl+jRyp747kbZZSAgmpE/BV8vDjfWWD3/y/LW3vFlboXVAOFtFkVpUvGK/2oSpkO4oE2mIh
WIsIA+cmRDXCvTB5Yy84g9R4Jn/GuYeW5brR/peJs+cDU+USU4Hx3RDfsRWla1evoL2GtX2X8x0P
EyHcPGxOFGAk+14YelqlRbvjnDk2Kb5GMhejIi5a+P+pXznJrbd+cf95TH15UyU8PxM/jNIeOnBB
DOXWNC3s2MN2hdReITzK2upZHLl1a+w3HeeZWRdXKqsSnaej4aggrtA56xhiqkQ/6BOKeGJ8rwAS
cYMwyVpCvDmBGe6/StmEMssRdFr4ckp9NQSZ3MCWXlxMUKThyJfenSIh51ZYKkBzOEPimSkGnCu/
5I5gdWOkP5XJb+OYFkJLsW/dDrmb+LPSlLAW2CyxbFD8mTPx0zaXJWFc1iy48gP8mIXyYCY4ljW1
O24sIiUm8OJuj2cOhG+fqrv8lHTvOrKrCYAE3HKaKN5DBmyTM93q829jkM9vP4b4jc6iflAuLDx5
m8RWn9PIYZeDpV50myu/LQbQrqO+2VVIgiT2fIyw6SUitvNjhKtea3RmI05vpLB/DdiKhV3nFKck
1PmEU+1TFbQBK0GrFdkgxdUfgnBS5B9+Ct9fNyymN2xWBn122EN1cUy+HpACdXWJfZkdZJIa9Bal
6oLTXgtSIf2TlVM4sEP98oN3GeITll4qqWYOPmeM9M9EaeX2bV2f4MitnPeA3T8XL6c7OpIQB13p
UDRxK5zTXsZByIzjldbykBN4PgCEaWARdPUB15YSuC2/yFZWBNwOhM56jBzi8RlftJUKtsKws+hJ
K8WE0BFgJ8rb7uNzCh1kYbsvoX55A0N96sUIxzinZTnuvK4JYe1s1JnmDzyZsgvngPrrcQ+tOcsY
8Ja0rOK8CTmaQPcD3p8605A1pMiJsyNuEEWh3PUevPfHUy4auA1zAAS8Gf+0rEHL2P9bzdRZ+P7V
CZYa1GmQKpxYFnkGet+KoOBWdCrr7g59VdbfrqkTZMO51uh0NqqJFxfeqsghHITD8StFf/KxUJ6I
39Czdv671wQ5oksBZm3rtSp3HWb2K9Y1XIYU/WsO3B9/Z+WO7o7pVMP3a8nUyPWn3mJezmjlCuIq
Ejxn/eQJ7uSTZ7/VJj/2mnDd/85ROMGZLtFdFVOEXEEli0Y6oscWTzhPPmcZWioEOUN+4oPbifkw
EoC9htCjomcNg5wEuh1aGErQwoNbruJJMF+2s4yhalWoee4G4kaoTxSy2PawI8jiBv9STu2PDI2H
9aoqMy/9W/6QNvAdfYBOo+IAX3A3i4sAicKTDQbAIyowe4q/IA9+hFU61p5T8CWz4L+W2G/i1PXi
LabzABopy6hkH7zN7LlfDOSAzja8TYCxqmT4kTPlNIk2nUfz4Bp8iqmlHg8d2XAVbRmGmM9Rj4Im
OOQSDMrszNIaPxGmWpY2tMHxacmhRJabjwyQKPgpq9kvgcE55/u7qj2nN68FSlp4djKMgxYhXAU1
bcv+YHFqRwtYdK8OcSHH0QxG7pHiZZTHEUEE1nXuH7ujU5LBbA6zeS3EyjLTCfwjc0NCOxTHfN0Y
seAdi+4GWsJA1DVzYSJHnK1oLziXTwAmArdzmqXrXO10Vg0t89YgjRte0DzlF+EsZGPJUFaPQMEi
FE2uff4daM2JGYUZJFiAIpjrykj1D97JBFAllms4DnxRHlruHdn9p/VINqK+E/jA7OU2uT/ZD2YS
n+qxaLQ70sY5wrSMoszjNaKxRitf3zjrZZ+8buL/RZEMxN0l+c6vK3hEgp4blBzQPX2W0xQ6hjFr
5pf0qtzH2C3MMSbf9NcwWjRv1bDL+H+1rlsWjYjfoxjwJAQWAAyD8RLLM4tF3TrnhS0cJtW4nB8D
th28IIVs5gfRxVhzSZuztlGI5fxr9aTZexIGMx4Mo25EW80cydUg/X9qH9OBRoNNEYVn+FzTQwFO
m18IH7O98V9KshadJtCLyy6MTdF6cAGdueaTBE0Yw63+O8Mb84Foun8fQzQC/bk4IVJS/sVwdeGS
F7OJip/zPzqc4zQfbgI2sTVUgGFnqXlh9XQxOh2/Kvs3G9iuMAf5wny4O5foIjF7P/j5hXoNx8IK
64y6xdeEx5UMvW8A1cvZOm/vmeTKT6dpBHVq7e9u5ybsmXTJlv7rhLoYrrVDOyf0Uhq1CZ/E8E13
0xV/WEAyLWag32wZwC+0koQdvEUCxexy2RbMuaxm0B5bd4946QFTHsDe+Wydi29gzyRs21RuzDy+
nC2SdP1UJNALUOJza5K0MYtUrfgk65jjIzP+VR3AhYKt7Fv6ltIANRGtD3oN+D5Q2njVws78Poat
v843KRSRg1JzpWp7x6/9BFkkagrOirp4wJ/NbrFOzaD2/PXYVSj+MV2lwneAET7gdpQD5McuMk2/
GQ1bLPOBzY35mFnYnvR8CsNmIW1XnQiezIML/UWWTQ5ibYbku8Dd08BVjQ7dlprbAnXzl1Pj0TlT
iWI8+3hqY0173EAIZrUlhpkcP3xxwfI30Rqq21ckY7imMlyVzp/0NMVLk4+78yveSXGbwb4/Hqtj
n8aE88YwXe/Li++rGtX/O/RyEVU7xNISpOCSpzKxcwior+7hwNGEXiJf4cXU852n7yevTjP3BHxC
yib+7/XUCiE9lSkk18KTeM3GcMzpRUkrELzoaADaBs3Jt4ZnX1+IimInhljvTLVBcFYuqWArWcE3
fLqTR84+fGUiGdTQxGZ500ZtT4xgkD3lNTyQkeyY8euSulG9/eHxjqC/B6NJ6XZwQDS+RH9jD+fo
+rtOq0F2NkRqByML87RVbyXQgJlcaHg+gH16HUyZ8hTzSphB+r7dISy4wCvjEstrCYrJinV8EsFl
zZ9Wj/Ou0Dn9NBFQsSkvHmYRYJs1jiQKAOHmGNeBcZ6N4rnCKqi9uzwOUzzz1cuCzeiY0yzR9xUS
qA+gB0bwbWXaNx9m2EtvAeGfM1rMoCbePIwxcDrFdbrt4YqAUzr7ir05PaDreZAamrf4r1IdeOIl
1oOTwa9ksiVNMK+BlPPm16UEh1MdwKkP7EQR6heVQdRzi6Ro5+Ss/yNAUz6T5rECfxaPuQa8yxv2
tVqo04anzynv7Kq57D0UgruoXZGX4mViy54Vf6NhTBp5xPLTn/VqVxg2WoXCFJCKh9BRrf4Wa3/e
nCvoTxfv6Kck+U8raArqid6Cu00dmV5rYigpWTm2Ix4OHGBZ4EdB2eeVQySqHWtG42y4vkKIqh0t
az6tMqARrd2Ofk6kvi/OGT0MH0m/zbd0PebN9IgsdXj3OUqa+Eod3J4vyZq/JeqOB/B+22yAgNT+
IQcsZ1sNUVXE2Qe/4mKDhxzn+neGvXAJB7+Gx5M+dQ4IA4R3V/qyweZdt/no/HGO+vDXC4ZUMMpV
VL3BfLTb9T+QDyuMyZI1QN+zPrxE8it/VYl70UFlbjHfDHEkcMTy0wfFgdXC1NVI9k5OKLtzeozQ
cs7amx3QdT9DwdhpwDcKLGqs8XfWDXTb7NorjtubEroCeAHGEhK1LmBBoUiTZV/VtdUpaqcTIoMh
Pibw6UtR0KwFzd3B4kgfisYAT0TTaJNGp6+7JpZVCl0bV3pQBdG4jsho8PFHKaje5jckz3W6F4+9
A9OJAmCl7i9wuwR6IU7ymaCZhY0vXwddw4UpN7a0SwwofVNbiEUAZSTg6M0f6vzVWyFSO1JjDNVq
tSSXSQ8/w8x3hrxiU5qP+BRJJd2QFOlfzyEnNuD/+pahZ3WSUTkp0opZ+8abnKJb7rtabC9Tzlb2
0u4qkhVHogckrkT3coW4ApKn+IFGaSWdtqTl3nzZW4JkUBk2JJ7eNG+B/4iDBPb4LK84T6CPm8fP
gBKtKxfi8jIxjMT0ITVvufiLgg1nTmJRpQQ+4JML8a39ofGnjgeiJ92mnpP1yxpxyOaYegcEUMc8
eW7CM1DaCCZM0PWRAYNXJ9u/BiBDvI2933jfKFhZ8fQBSQ3mMcFg827GZUUhuT+AjPvNMVy0eXrX
ZuFE8Y6S9VUlfx0W0pIzpv1jQOwCFkiw3b7KCFkSHDlYk1IsxkJjFhhPypBABD+Ew6MjT/0jKT6B
FJxkTy5nM6FscbkEmWpmQDW8v5FBU6fSahqImyeeBvp3ysJfoESxijuREj5BBVlxg5KPLlFiJAs2
wUgZ1pRTwhSAUO+ig3J22fNbnn5pHxryYuV4fdX5OQ7bnXu60ig4LCNkCC0nQcfelwbkS2esP7vs
dURd6Ad9IEZuKCRDQn0DQ4wzxJGF3+/WJXPjE350PntNdyS/iC9VgxfdT5eB8LXUoXa54B8lSPCR
arSeCN8EFODSN702xZ1SeqjqM6Ms3IXVrGSaK2u1gVwxXMHPpehmOcCMR1Ac5cs2/Kq9Wk0YiaJA
S75wIcQ1qrizzmUhT06xSjcyL4lyNRBACMDT/seql26mAz8aIY3GeeQMsFrK2sD1gOz/HpME18rS
Me2r+/eVP+rgVMMoHTatvuwZ4riplu3hJJyAU40+nonUs/qcZv7YUSwf0rpJp1dtW2fDBag1dq11
NAaWAReJtwzW8U1Iv6IO62DiZX6sbRS+IcX40++8EmdF4Hg7v/t7Y4pGHDx/q4LLC65H6r7kM2Nz
vCKCL/ovGB2iFQIXetmFqP9R2Iwt5JXkb6eW7lNQMILGwXQ8KPZq2rX5i7fIvuaBNGN+p65FuXlV
fT4BVk5kgau7B66hTHTzDU0U0smPfT5z02TMY8NB0TDieEilnI1LMkAnJF4uyvz4P+JRdi3jrC0/
ZxDo5fNNNR0uBZajcncOuTTuzKWy20pI8YjTO3mGWEQcs8vPrx7gfKqY58e24+jCnxUhaaEFGlyY
EYl55snBRFRSe6QAoMgzvqt0xTeDzf2+xt78xrgOn9vOdcfHl8NFmZKXoq9YBmXzs7px6Sz9C2ZS
+cHSG/P1vPC/PhLodvYZPtjZD3J6w43x4axjITAVUTqvsDJnKvZzEssFUmeLilDA6ylkV+6Dr5fz
q+mQ0n2Ny7sTrNUUktNRxQBxOWJz3O9kCKsuhC/BnDQGPBvMD/j7AYbxJVlVd1vEieCd67zEBhYT
qGHIaM7e8jbkf24giJm5V3B+9A6GpaPw1MkLimXRR3cFdkBvquKWHNFvCj7Mlav7nlEgFKwcGond
xm+MiVYPyaNH8317OGF5djgFSFE4a91F8Y3pEFHgABavwirZI+k/UYyCiLrqKNwH6ebPzVHJfDYM
3miwOSrtprflXxkqPiUS8uQ+4iYiAYxZJTu1gyLdSGmhwZ78WFIcAtTaygjaZded6SW+5obexLYc
FcPYP6Rml2hX8n9aAEELOS0H7/ikVq+/JTWGlvw/QvrXUPJ1M/FnQgBnDaH5u/aUB9TSh7wJlfB2
XRAw1EILvXEA3GsRPEj/IURg1JZq0T4jb+tEdetFy+8caUoGfqIQCBGWo9kIWLz2GTvDjsiVr6dy
wLauqsKvd7RqMelwavgRCWRxGdV6a29oNnMJR84jko2GlvgPl6wuz9+SVHxgaCeuRQpw+7qUjKFL
CZVNdArZG63yENdUdWBS/WC5kRHWNkMqoGjNiBZHL+G4dWeX+2VO7sf3j9oxQt0oMSdD+Uek7kHu
/GNI2KaxnN1AuOAi40vjXFXhOMX0ZlI+ksWQRWHRMrTinGlfRhWw+pyH3mTTrFXBibVg8nJDCn50
L+obDYUX7lmbFDKe03w+0Q6mL+xA6PYPIc+gI66Jn8GUfEYO3GhgM/tw7Kfexz5xMeU3UijFDSSA
pbaJLIUJ4xYhUVSRQkLtrVLaq3HCO9kpw4L6BQ4ZYhOaSMcxtstWdghKO6bLs/nWv6M0AJOEKiLg
qOmJG6On5dmpFZT7wbv6y9uUf4LoDrRGfIiJgjirRUmeaog7yG30g92vrK39V5KQRA9boLXS2UCJ
25O/YiUYeoWDNpwtJVAK285jK49c9DFnF9hMNxF0sZsPuJEN4sKTZgKmwn9zbmrCjWjZBHbvhMR0
SJkEAUyvl0sbUwL5CkNPuqzuMwrcpT91RK/XEwxFG6OiEuwk8mmb6tcqPIVo2Bfu9N4Gf0vGF/so
R33Z2cVOTqonnpWPRQMuwUmC6ZhdTIkxDiatwCIe/veQuEq8IY1EKFmHlXLlVseuN+wwfRXbQXqH
1OC0V/TKazyd4eu7Ihe5tCyhtiHVBUmF0UoIE1Z0qMNEJ5EEl/Xkk9VNJTicWAeO9qSJNvyHb7Ek
kDAQaQ4Jy+M93WuMhVSoAAPHl4BArXZ8gQcJm789yiaf+HRgTRNtr4ND1pROfVCLsRcngIIqMmKw
wX+8fI16d9lLlX27US03uYHoANJQdBBeCdqjaIOe+QZd4tSyIxEZ1N4srm9AfWSlSoZOwzg4ow7u
csAPTa1L+a3GZh3nAUWvldrq2Q3Y9nkBBJdcx/io1BwFxn6rVy6Vt83hNt/F5OJSK4RZ3FDN5XT8
ACoFpNy2bqHjls6FPpIXlyudhp6GoPAkeO5n8QZ7gnRn1QVLhwJ4u/iiyZ04UG6l3DaR3rjfcyle
Xfs38n9BDmGtvGPClB5tAkqy68YWJNN0UJrxRn1vTiHSsnv9fvPnHMZNPnC5cDuGaOoykV3wfnWo
dazqYlLgt+GL/YojPF6BO7TCxPlOiTSrJqt/x8Th8/aqOS7C0yYHlUAEuRGUmA3AN7l3XRrRJpf7
jfbaDMD8Gc7LLZJZFeYvw4R6xI2xk4fUw+uiJpgnEeAvU9mnYJ5pL0/fkj1SAvngAA4ph+QXHUae
P9MWfFpQXbemlQ+4QmwI88H/vymMAk4oOKtJEa0c2Tbt7CTJBQq9GSdEWi/Remcbe1Ex4j4t3Hay
cuW5zID2AH1zXCmD2+DHFofzPpQOgCVMT7okZ/lsryz0VJmIyoUU4RtxA8KtYEX2tIOrkvW8HCI2
FLu3F6Urzn9wsBHjD8Xo76uk5SX69zAOLz0fkspkiaxM4IxGadEsN+2+xzsplUMrW6x4jLpik67S
rwdx+QqAkReXPxMmXE+csjiUPiloh7M4T+lglXk/7RXWgEPR47cou0eqRJNIJmPjpSRE/saFQUWl
R4DLkEP9ZS00WTk6oC486sxHBRhCanjaOruevQv1YqlVS8Kazw7RM+ah7jAA7a3b0ZBDxDr8YUY7
Pk4usS2USTCreWp/RtGPl7L7u+9Sm9zEG/6ZVljjDvOIqYtIpM5guH++nkf5SWAAv4Wu68Jyv+4f
iskPAuS4lnoGq/AgLcOBWKq5G5C/RNdaiLOhY5cF3Vu3IBGfeKjPVIEphIT10nANHQybxT2NBY7y
SOTEoUZcX0Hrcci8RoLi3r+evUqh3fk2JwVgHTVtI8wIjTbCUsTxbP7UXTnvzgDtI2laug1fMNyx
Tk14tt/zTFMpw2bJYUA3sljRlEYdSZ1ANR7B0F1PhmpmHGJxcLElWf+yZH5xzy1N019X31qf78JG
zYLiGQcBIlRtfU7GapjrDGA3d7NcpoylQmb9wdo8w6hpqsX5rpd34z/cLVBx6Op1U+rkVIKz3BVk
0Cc16Tf3WnuOCj1L6gS29IPK9jnO9Pk+LnTfIsfu7z4X3/IzfpGMmTqC0JbdHgq8rlAIhoX0+AgE
0Wp31gOoWW0HvnOmOQzZU7S6fahxs6fSrR/CjIQaIKuOW1ZUfSS9ZZdUVzJioGz28UOjOlI6DWbd
g/7ermThXUnbvDLduHroVkz9Y1Umxx6puAIa5MfXFJcDlNeg8M6EDew19KGPjT7GeCjt+svHvOhE
iZ5zJOyp+6xcalgtSJnYwAHtvNXp0wr4+/22seq0xrDyOnI3kZQ6DxuuPedLE9FSBfLes5I8FtEQ
1R40DHBSYE9vtKtUQ91ThAXYUWFMwmzaPLoiIDqNimlaAT1y9njMDcd7eDh5Asis2wUqZY3Bv7+F
NHdzqw0N7frwvZrBoz6VMD+rPFL9bT1/HeRDN28drKxOH1YuET89g8OZ5wEMcuKrJBOy1obev1jO
Gz25XgyuIcWOas/tCj3cHdJ+1V4NV7uQ/CL7iONiHnhcfrYRn3HZ7q8yg8wwnHptiqHdyBTSHLzB
azaDoWoN+t+rv6/O60G+rRo6QMcFL8kYZazRdpTt5RtmRFDoaORv/ar5kioVkiiz2nxTtUYgV4cO
vQg+kdbVd/VGHhIXoA1SEWcLhLAtFaopVi4MX98N2twZLMP/AP4nX7TWk+kEy+IsOiBfM5g4nv0r
3nX2g98T2ChwqR0ShgiQlnVmZKTJGs/V4bKVmV5CAO61JxYgsy816odEk3wQz2NVmWKM1XO9gIUh
Jlo69J7uObcGMiIDmUXUfksR9oYyRMzf4wbUExtrtbO1MYZztFRLrBE66goB12f1rmQhQ0vKHvi1
p9JMOirhYhNac617sc60S0Tqz+BgdlxjgQ0qaz+IFpBmLnbG4eA2N53+HZUoB34WmwHWrtqS+TjM
XY6spMZ0AhP4SKOzGVZmDGcUN2jEN6KD3r1xRSjSs2ZjSPUhjEGP3fN46v8sbS7tfOqsT9IvKp0Q
twE3tvJ/fJ6xAzc3CMZYvnyJRXSMy2gAcDcngdVj3jXuVMYrMSj18aWBFX65rwzxdPAe6a9hSPtI
iKGdIkQBORzghanMDdkVnpyESNmfhdvUEZKQxS4wLNHEDlcWpq2J9x7TV4pc1k8wit4gH9wfcFSB
WVkEfLIj7eUv++uwC/4GlySZCkw+YLBHai1TODvAFq8OALrUy+gBVc4smT+KZwl01x1plLm476jY
HE8v9dnVVvMp2fdkjzoZnQGFVudOrCDiEtbP97rEQMWZLpTzA7d8v+HsjdAdju7OO9xyUItplH/v
jn5jEjArk0slD58zntJLGV1lNavD57y4LVi4Sqzeo5a+/6wYsPV5jS0HV3xxCSDiHuZw6anQWt0O
xXyd0dqHQNIq3iKvZA5XCFccyt4u9xD0b5V9mVHeigVaX7vs8vtMuZe3noj8/ThIg0fxsU+7r3An
SNFnrOaBaIsEIHr5TMSoDFAwF5fgVfV4o63YWX4FH9egJBSbNGQKyxQkXXdRj2eweMQuBOg0zaV6
ltvKGhE0EVhaey4LXDIF+VayjC3XBNpVhieiJ5TsQ9CkyK0ia4rmDnCZELjy0J9FflAvgWAOzrqR
h1EnB0c6QOVST7ZF/sgQhZmxvsEJM6LphKKhRNc5H1WpKfu4ydKaHnwiVTNwUuvzVSExojyXmlHp
56Sw0EfrAz+ecRwecdmJncqp/zwOXxS6V5NmtwLLXeG+7TqIspyQLcdDLPMYxzpaxXy/SsCq0TuN
/wrkZIXE9OVmBHTUA8s3wv0Up6CbzyQyHS6VGtrWYEqSSgunS8NwMyDG9zKzZdEZsZJ2S3/ySeqR
eEkVPb59TNNHDeW+PHMGssNqfsxhSK22VoM8fmj7plshKqrWCU1/bzekf6vctJRDLNFXt+8XQVzB
fQeNHRpq2rAMYVdZHhLAkh0/YeHsEMC86oX1bFVtgV0Pm912auq/s6b3pQ9gWZMImNPFg2aI5IYH
9k8F+tc64WL8Ao4I6ofLX//vsCVTpHZzZ2rFRDHKL8QRCALFkmXcuciwHjA70uqhANoQNz05GWlF
Xk2neQoGR+t0Czhhya47aGqRVcZXqvODQrii83H2ZlJ78rmRb3JOU7hBk6aYdMMDGzr1UKsORXZG
MxxGIMb5jUTDl7KARlsXYxp08iSNjEoVTwe5fHSy0AJS0uYAwauCbyqbe7M/9lKcM/Laij6v4Y5Q
uTBlhI8ZNC+NmYrfRv3a76aCeqVQnpDnq2uFi+wDuCHfxiA7hu5LCcgU5wyAvydSE/FbL8KCiQBV
yqMaCIfPmqiAvaro9BrONF2Cxp66+iLu5FI+gfs78FV30A9fVJ+9hhQeLbfduxfxgWO6XcERpzVl
vuK1VE5iA5uN7MaSNu8oAjdsMLMsawJblDfGocSbG0lMeGTlH4xB6wJNAAoYeFwhBT4z0/YUIqRP
xhCCHFt+fx6kpW7bYxm+MpRN6QysoQDUMsFUA4b7zW3LSS88XvHAGep2PEDaOkzbx1BNlByc4Gt2
2s9NGwsH6UcS8REJifS9jOQfAPRM8y4xKlkmyTjuq8i0uubXVt3cFO+S2Y9zjfru0rETNEGI92A6
/E0XoOGIsynWTJ2dbeAiYjWO8bECMG9NmhgnOFML+hAX4a3IF6Cuod4f0yElE8x+8yK5AK7ZT6wi
XxEEPlXHAzEVM136CMbB0OmL2Vwn2tfhg0Xo9jaws3A91lACWcgLOX/3r+l0vewwKow/xz1zQnH9
D1ChSgEcu+FL38TFbIaaSkwXNQjRk+0alj4QlicYSKwCaDQjmGwmPuaARVf4JnuWcz4srwo1dQyg
QnMdVel/HDq29h+7cZva/TwFthPPyCBDmskEo1msPHM4PE8IBEZXAcmqERhBbldIDwRHBV3kuyn3
0GIVB1TQA7GR5RR+40GYtdJvLz/hbJAcgm8NuOja4NjutR/dKN0WR+uFPcEA6VWaMARqaKsoWjID
bXSQWOQBjrsZbp39wRdtUDumqijdaL/0ukzffq02sINdKor5jFi6HWiyXAdyCsRv16sAiCAIJyes
Jl7/1bFoTk9p5Igmm5SpNvvUbtbCcsX02NC0TTvFAhcf8b+iPLofHz6ynqnkLQxu8K2pxGfLxyZj
J6HZ+GoMTGgdiwxT5ox3dsz8mcwkv9qh/3ZCBSQBNpXVhPj7dYPCJBjnsslTUAf8mlym/pa3MTkl
PnoAybnc1zBWw2OryB0QyAaTa3Xzglx0zzBTV3dRRgrSCfuvBV0tJcsckG+COY6vsyZachqeERrH
XizxKs6pAllQG3NBbns82+iW++vSJ5Cj41u59DLO9EpYlCt0IjZXt0n4tjpGQ23hmQT5/Yep8cak
0vqfbs41iV9UPruvuTaEuJQd4HV/wr71hZQ9sC3Vv5pJanAsfQHvMjKFQwT6wn+17TxETN2wiQo+
19N5ukLhYS2nIbE9vvChPju+huURmFw4VOEbPI8IefrEMrO4RoXjDAxkeHQUp3ucosUMY0FYpLpu
y4gX89n7OipqvB8iOEsoJwrGkPkItLUu+t07oCU4HDRwV3CSgN6JzzI/j3qbjFuy+2Dtufxuy/f4
+s+Mk7tcoue7vMAeoswI2EuADV/eIDJ+PFD0ww+K4EyvTZFLUbpWjP5/0g02iBvh4XyHRdg9h0xV
dUOiXkXiRWZVYDf7Z2cD7yFBBRpN+tNhuhuJPbbqcRiNky60DLc5v0A8NlohrJbN0Dw1NqH4aSWv
7fRUPji93Km99gpQNMeb+8fTMtP6yJPkjBmAWSkdlRyF0JDRFAPVFlXULeWuIK7Wgw1/raw7ZE6W
+zK91u4g/+fZ3OYVqrzasvsrJrtIe/vUgEt2r23f3h6fbZq9fimWfuBsUW94DJilt8prk9EZQZEO
RPrjA1QRrrpieTFwXlVINhmabCX4O8vBqEcsviQEXZVPH/P69N3AsABlTFGFwTFuYyTAq2JZhaB3
LmRwxi0nwR74smws0nbIMHVkBh4YxGqvVn8mLQE4tdxgw4dTlUr8jIQMwYcQuiDA5zoQbYCllPGP
lPNjTo3s6CxYR4cumz8TLCfDTfbgcKV0hgqTj83c0QmeMG1UMDUZ4BIZcCTvnVKL+II1lFX8n8cc
J2tCDuxf9GiSRgi7SW6AOf3Xy+ZeR9YZu+CnTJNUq/2pABPT/v3V7asnI6H3vP2m1P6j86b+ZSb7
b0mO5K59u0sBf0pkAbJWi5+fjTJ87c4HPQyssZfw7d4VKsbah/ZdHxJ9Rk1N1A0YhctIyvYjcWqJ
yniDklDoVETBl7vHgLYWwBGxi9T0gNd2jBmBBtn8DiCH1mNYI2KWWN+bm1nwCA/YPnrTl3PSfvBQ
83s+ygbO7zpwlDl5m0AZIwPq9yb+hoV2H3WhWBOnanX61dQFiPBVCWJz6xBoPwytEjiatRY5fgCE
tEh91dc1+NAt8sJQtthGVkRne3x+K7dnTWE7onMvYi/tiDJIPYlE1lIcxwbEjghZ2y7zPtEvOql3
e++UsvZQ2fwcfoF+0G4XT6mgwgy6uMjNkyPiaCuL8X/YLU9xSEdD3T26nOeYAbuQDrPg4rLVCzK1
H4T/sw6Rwahw0MlOjNFKZOBzMS0v90xP19rr166yN1ie8xsJ+XgNcGsox+cvJXKBncU63TJiHP9A
8iY5iUIl9pM/7WsdYE7K3U1UdYfthBUq9n1Jp3puhj6zqrMriI4swqWsKFMPyYy8VIcx4WGDgUOH
Dn3cfV/WLcWyow5qJpL/zuk6ZEFj3oT7YPr0MK4mf4IeIs09zwbcLYtUarf0vkdeLUuS4nM5q7Zq
q92jkYEkuAK1bGKWqMBpXNF4YSHygNSdV27a6uOOTxedVJyLk8Xvx2rYKuqZ6CfH+SzspEv5vwaQ
sy4GvNZwcSJXzFZHfacWe5OWoTsZ3Bw64LAXh4GdXO3s0r7H8g8mC9Jg8ICpyrmU0r5OLzWzB3XE
Vs3UKSKvWXDvy09WwnbR/dZL2Sz8OIGzHqKnmIbEBUowIVa07UWFS01vAGYL2vYuCzfWD1Ia0zhe
L5903EO/x084HeHKmvj8gRRNHdm6kdd4ClWBsnl0CB7UO+bkEm+mLAmwhxRmrFDgW1Ni2nRAu6vQ
48ObCQ2HoRD2d+RlyX96c7q2zeeLbVREZtuNW7Bf5W/ypiH9fZjcHinm4IDN4Cv8zUaQX1kkGlEf
XPty0v6rTaiUcgl6upjeX4Af23mmrB7A913CPuo8WwfWGm+8jyZCJZFtKyXNOQz7LUws2J29JsFp
mOnmJdI95juCB5YgniOZG6qftio6wwrWdvap+BgiAZNpsinBGwKgDKX+s9r/P/6LxWXNbr2aEQV5
N0NVOONH5ZlXPUPv+iVPiLWBrPxSom+Zr7ndEZIEj6gTuP5jpaAKapiPrwRHjy3ZFt/RxqA3k3+j
+GeazZLjjnFw4YXWIEA2Kc5pXFP81xS+a9gLYevWIp+hhQ/pqmJAexBKtrEgED4+rQNBA9P4oT02
1rKFz2dFtL/gj2/5L7aL00RV060z/sNmHINa1YnahukPuJ9a0qMexTjjvXQi+2fZpHQ3Q4/tLeBF
eZA+G3c8Ws3ZeTUIPb2ToBFOa4+2uSosLcg8ji+r6Ot2OEBiqeYS/Rl9b+t2mCowFVlmAjVjMhgL
39Fuu5x05o4krkWvkQCsaSphBrRCd37FGR/g++uZoCXBkBi8ZbsKJS5E+y20z5a1LWClrbl3FAPQ
R4kMNHOyEtCBj8ttEEXaq+C+7/KtRQ1klhTxvcVMdCYYS35X7wMpSA/Xk71vlW8KlzzeoF1fftrp
mWHJHK4vUWh5O+qqP+Fv1AKdulwOeMBhhmcN7bmWx4RlSdCnTZeHRubzkJ600SWlanL0bIHeHLxd
qRbViak5xF9MPJWfkOJlL1/HsBVon9RmQpazMFm+V2gxMBg5iXykrp7AzmjE7emH40+Bum+DSUZj
wbH6VBV0QB82wMvVMm1sS9PHdJSjAsgfsUEL2Gm0PYSoer43CLFQeteBi2gYwdXyGNecj347j3xV
UBm0DHjx0HCFjchiHr7i9e1B0uEGcNlFkUTLSiWg0FI7caFFWZ+Zl/i4UkKIfztcrVTl9hY7JB4l
AtMdF+Z2Xs/n0r/CcFeYs2Qxbko1R3QtaWN46IM+BRE7uzDQw8/UmpJeOtDrjlPYgKety2+seMD3
dmO1MBaTJJzKEupiTRX/4hwb9ZGkqM7VRth7JVyxnz1k4iBTftwEZACFX8MNriPZe5hTORgIJefT
dZL+elhg2itONH/Mw8kvPZ9c8njK+JrgixzFz4et3NjJ7/+l1P+TxXascH3FDBnB/093gwd3jaTk
Sa7GHN+Qdlbxio4+bGlC4OPcwX5uKU+/iG94o89lo4sN30giI29m5BFL2AYFkn7p66C7IjF0Dw94
xpaam8/W1xhQxEmYTeWhy83/MT55Y6JTm8FrAkUVvxr9zT+4ZJlJIAlAOlMcwaSWJxbfc1Aui3Iv
YJtXo4muJaBoNSUQeAkgUxqBgsJwoIxPFPs+PHQx84rNi0dObqaZy7dcmqoJU0GI3tWAkNoPnD72
WPH/5fdC5jg1OtiJ1wEoZS36P7l8C7HYbsSdDlgos6l1FYMpHzIP6Cy2HMBQZpZF+QpXICBIPPiC
aUxRNXbnaLhUrpy4qAYXjnsr69JtT4mykYahV5QOa4mCrByUIVrb8oknHo/bdXfyeDIocbAdSihr
hCNANOIUjgIwEEKoHa+v7J3ruEBUDT65wTwW2k4YQq+DcejdmlgGD3FCAuAaaglK6W9kMJVoZui6
YEAGcd573yYnTZ94gckip1fjUESjVwDzbZT2TqwbUmO3NG+3tyZdawBxssHva3EEFwhYGhrv3mXZ
YTanagTfurpwuVOMv025g2EUzEoSfk5AQ5pXVVnSXx8AazsCBxCqaJGNBvPz5tzcD1L+xdu0+BjB
PTIFAouctREuYbbsp0SFYLLqH3GP3OjHwGcZ3o/A7u4+ejnNM7wEtPzS7kWh/0aIZYn8UZEdmd0Z
tFz9rnIShgAgH/aKN3Xod1nZj2aN/XWDnCuqy7tWBmP24yWgrCITz4ymjRBgSOc1WnCF0ENmaH0E
leI3MeucDeyeXasI+xjCCoXy7CoKll4CYJevJvJ/nraGjZ2eE5q2XJgfe+FiBJktC6ShGb9Da+0N
TZICtDs9hwvlO+GW4UzVRmrPZw7P5t281ZXlBQ4dDiJ+SLeacajG9pdg0IjemzqRZ/qLm8HUZDg4
UIUAQYIT1WyXtXOigq5OgKM5vPDcDQnAytGW7T05U5bL5lDH8yzeHqaBfUAKstC3KwkSZwvVmxhE
qJRpfkuVyg4gcKGaRMTdjnl1u9ibKWKQk9vJRjJ+Qg8h7VEBEpRbXB36RVWftWFB2AvD0YkuxozE
+2mtEoqCyMWwNDrOO65TMQrfVl++GDkDgqRihJQVIVDi3p0UAtHjoxIYefCWC2mWNRKoNAfo9qfu
v1yKTuG7YWbR4m5nQ1NqDovDaklDfPPA8ZDN1uOEjpE3S1gvxGRZuLTZu3A/POH2PgLW3laIv42Q
o4bImVOMRjVl34YFtlCN0aKT+jJEx2YwKUHFf/MBYHByEXsU+d4RyKthztuPxahRtJ/cSK6c+l8E
695B4pJPtp9BmwhQRRhlBhnJTSOgqZs3shQSmZd7tjoh0zVUC+fBLHANXPfB/oRLXsrLCh74ip4X
KhvFlQT+RRJ/d+boZH4YbWOFBR5vcBlOcXJtHT4JVq6s5oRE5NW6qhqo589Lod3mijQ0zXQ2ORsj
KWUERtfHP44o8dfizUkIlg2P8Qbq9uhfSZxNyX/QoAd6qh7ZkIxyHEJwgy71ZEhsMcmRBkytplGl
BgKuyM89WLKJuI+bu2zhCxA/o6+3KziUPmLBpjUa163Dynmp4ef/1vEfO7qWrvehiD7pyFqfWPu/
+7aabrVhnGjTF9SUYqGM0lBVCi4g5h7y84zEKhY5s1CxrNPDuroxt7JSquO2W4gfGQjiFM3Sdx2T
MiFlMDUDPO9z6gycGTdasTrB1I0FzqL2T86SWMciWXTgNw/V72KzO9VPNJFwSXXwi4GUBVndee4I
l81sy8BzYsZXoWbxKXYBLusrleS8UNotQUZrY+tVW0Z5927LFEroh/6a80pVLesToSLCqdNfVPtf
vkxwJ7HFwBJi0HYg4oP5yFezcsk/invMYmykT0URRhdKJDcPPD+cs1yhefkdqwm/rLvS/S5/fp40
wDWdjRo9F+pFhuPWCsqU4e83r90TzyDdWiOUSy3dYqhMnEi0A8B+YBmr0vcjW7SxkGl7u4aGpnbs
1CkZHr/5pHl4zT4hhkEyUs52ZBoo9lCnB1cdBm5K3DXM5MHUiRuDcNxGaFpIH/+qw4Zw424AFvy2
eFopdK6mtAJNYx90PvoPSl07K78L+HqFRzSnvp3MOr2MueHdaECQ7ADbBOW1DOh/3horhs8ft35n
lVyvsvTKlIAL3tDOmRgqNsiRBZwMwePn3SqWH62yHEFSuMLWG3M6oDFCyhrtyH1TBY6FvfN83KYN
lkjEzDEOWa9aULh3Jgkx/Gepk+nI4qDOfOuL3DtvYfPsgHGtcBDTsUA1U/ytiEyF9x/ViysJbS0w
4kMTDPLFo7jz1a28r6rKIqcvc+qVACiUWdvDN/a1QpnVVfn6XnRvBe1YCFN5zckJo8T/HPidIK0X
LEB6EoFipCdGZP07YcPGjqpNB+OI0KWzHWme2O1ow26Q5F/JzLNgfn3HaPKARmoQjHzj0e82oYIT
VgFxAbT3eFUKbp4W3xkJnKlK5ozk9tEfZ8G/xyhMy+tYvtZymflx7ClwCvro6Q3fg8oYyGs5uPQN
l0oGYD3q00f0CDwylTj2QoXJRRXwH7BiT7TgROhKdF4FSlhSyNMp7s+Ks6bdl8By1Pvb1aU8LgWf
ZjCnht4aCwbfcfCSN8HV+00KoSHYV47qm0ES3x6hTMb28qRF0rAdw6WB8q2F+HaqVQnwqUJtRmz9
64fsAgviegp6SVrwVnQy98qUwJyWgVNE4rj1GvrDkBotQA5P5TWn7ChXwektcKYwYTxR7fsFTBGI
Mfnk74Q9I4QTzcSA9i6bfE68k7dwJ+I2mODyWqd2rq6nH8nqF9GgmNhw7C3vPmPuDs55RFNz5dfN
aTpv3K1rPOnxm8DFkEzvsXFD6ZgFtr9vR8epp8rUBiBFTG7MEPeWWHhRnV/unHdRMNXVzKWD1q3f
kuBMOZ/oKiUFvmOjalZuICIrgZD/C2LNj7VvvQgfHE779RLoYgNT4UCL0Ac7BNMg9rSwpzH91ncM
okZ9ee/yR2YuWCWS9T01eIPsrUGqkIZKtYEFPMFlNAlukzZ2Uc8WEUy24HEgqk3+YGQGmUBOhKlD
q6NXIADzIUYVHql7cwe9eV4XZKZtob+gO1cyYaXbUuG2cLx80UsX6KYhCyds6N5Q2pA/RHRDJNPk
csHVgLk9GAVq9LY0LLfnLtSUN3ThNyw9WmSN1xjbsDCjKOjuH+LXUdNkrK9deUkvquPFyeJOLszG
01uYqaoi2/E/Zuxh9eIWKNm7w0oW3PBe2HOg9ZQpohjFrMZsCCDX5r0smY3Fp6MBf9/oGMHN6jMg
D+/EtqFg8NS/ztKm+4aONO593YiVoLkWR9ZzGeq1xT5qa5AZy6V12gChyjF+bLXYD9GtP8AIPlCO
ZYnv8WZPL3LC2WypkWAvcq0kBxcL8Di8oawk8rdLE7mMmoogRdOr/kiiLonlUa2gV6LJHbqQz8a2
A6rt0ibY4D0jrC7VzdKVXKq9oZ1RuFtwWYM+WMjtlVeUaHJgbR4oGQ25jPvzFiQTXUq2cZWmmOBD
DekWPoJr0iBeh8ycJDrZnZG9tQdTo7q6ygTpcsE0Yr5o4XGJXPNDNlCEEbPnA3HtxXT7Da+Zx+0Y
TveD7rU0+bsPDDbuEKlzUrSq+5p1aCJchWdUkD6+HgIwJUoIDBWib+tNCpz1crSoERdSamN60meu
4zfMcBQMNl5nISz/KwVDBqM495eZ0t+MkEEcTiH6QRuEc5CCnh5mKEmik/1lvFPnxVsVMCrA9d1q
MpGnrL0odQv49uLI6kTiRVnh7Oxaslhz58Sgsobn1jb2P+PdFIqr/nvfJlOHPwssbULEbgPNTURW
PsXA0i5YYNR0fgrnYilRk3bp4vgrVdbrkrjDifx3QE1Nlc54+eYh7ekgR2Lb/m+zh4iuRhGJGRQT
w0tEKk2aAWy7IXah7qKrx9bsRvQtMJyIlaxLMNMAjyHMBCICyvaG10bibj0qdiBDU1yntNA2GIQD
sDuH96jOjoLQpSqDr8cSaABglo+jL+EjAQCgbaXPbpeURwEHG22ewH+sqWL763IULNSo1kwrKPV4
JPfgpqD1Fdw2F2gUwjTZY7QBm7eC+2dRx3CZemdjZ7r0I9/GcvwOKqKwyXXhg9rgMsBHo8ENjGSy
P7ss+V9/Qe7kgzCNcATgjwt1vwVAcCyECYvgrsQftM0Vx1eVLSYoNQjb6iHMMBrDWdmdk9R07zr6
C13MvUZgcSVZU214tyY28i/+6d4qxsm88HUicG+mX3PEJlLVyvWUBdNN+bAZT2yymLxAObiU8I3y
/G3K3qcx8I7kUslu4NOjN9et96bjA6E3SaTj7gDW2hkfPTGfHkpFYCKjcw4QpTnDWAubwNU2SNPC
bX0ZvDT8CPD6k8L0NN9dHh8jN+ovFOZ+3IVkvOTUUUEs9rJtVayl//oSgpOsi0DAPSaSPRKaZ74h
+v37vTBNbmC9dfE1c1vIkK/RW0S2bHok6uBruPFEsPDFiIVAxVp9oUYCvq+OMehIn7PkHLI5ZaO+
eykreJ4PKe1lxOK428ij9wSxN2kNnwqtnotl4K3P+Y98LQa75niyNjJtrF26uX+/8axvFF2CQcDV
2SRQ87bGDNml1yW2c4XUIiMs0+kQNL9L87fW96d65TWwsjGGTYOwH7KbOOomRNQaej6oFj16Geeq
Ind6bEiR5a3J5eCB0x5zCYmKeYCUdfqyqBPdJVMR86Rnd6DI+usCchv2OaQQKFjeSjPYWLsCaM4x
r7EFbKLP7Y+RduRpVrF+5k8REFeHmxcn+53gYRpqpz6gaWjfKGr/d4k0EUBbBwhYjeKg/I+YZGMG
TWRzTUXKMCH/Zlooi7BHQN62/NmipE7LbCcHb1yerjVORQz+r87+p8kkktPA+9Q9mc1SkmuaeXxw
f3lLstWyZwfkliGppSC1B3hwILHyrg1LVglDU54l540Eaufcq9Hp6Z2vpQQh1lQG52OG08UIaiEh
U4ugx5rtGDO3kncs9gxmrWeBE3Y4ospGdAVwwu7WHqdGbfJwofbl5D+TL3JaH+UjCI6qMFD3os9w
3taUJDDe3+PBYhMzzy6l1SqI7rpbW0vKIX5Z2heD8Rl3TrE+YMU4x2FA1Q6oBEeiULcQD14rFZTx
3qDaeK0Kr97SpBZUcrmOF8mlQFIs2Qu7m9leuTUxIGB7IfSuh7K2rjJ1V1DzKuOgviZa5M49w294
UxqSF66rUHWXj7/dgLJ/4zXhwb4sS+58P1PDQOVDYQrgcFjb22q6QWeEKMnv//gTNjPLk3nuQ2/i
pAF+dwK8npu2m9WWFji5u+pVwu0jHYA0qmjYzMzmzVvz62I5kifTkkUF9B2Sg9FWGfGYmGN37k1X
7EHZnMK5a2MTbZMYvYz4mitDyT3zQBWrz7nqm6brQqwPAbr8GsK+WDL0yD9wJSzU4C5xWHb0F7az
z3O814ZW8GRoRmZKRBnmG0PROojb7AaLLv4DmbOpe4WgfJ8JyS4y8P4s628cAcuIc9Ufva6ickxR
BSC5KcWgtNGxJjgens6THPZ1AH8iPSFAAsH3Y3rKR4VV7ePMjVVxl3/h6DaG728PtbDzKg0QYTeV
lg7vuZzveLqqkGw+Bg4w2461vz3MS+WTT/rUeIDxy3lb6GGS+3YmcnOFHkXRBT6clo1L2+lYJJ/g
6gegRLNrGgSZdyZTt+yaqvi5Y3oJwcJ3blHp8sQ0PwxaXfma3ii4Kms1Xyoec7X64wICnJdEjF2c
bc76y5/x2i/lXB1tntn5g1bHryFZvcWABf+yhvjlzNFpbvDG26thDLrT6HBqxqnNKJEuBWlpI+J6
F8YlhqlApToHSm9HKhaXtTeujS+K+OaJvPEJZSuoI+uYicfELm/uDSTgPbhWp5NA13Gp5DJ4lh6J
2VDNRcJRyGitJAPSLpy7pVJ/prdfTbzaQpEdLYAxjLLXRe7VMjbVQ32GimR3VGQz99JJ5dAJjMoC
ITg6FV9fwM2UfUJbLRkoAnJNAqdtcFJJByg2TsqgCIbwOHhe/j55NlljOoX8JBGNob+s/J8HSucw
yWo148pdUCP7ho2h1BvjQLYyBsOF5PZfWrlcH+yyYne0l7Jc+Anr7QxZlzzbv8fk3xN+KER1wzOs
fG0UGpCbwXX63xJQ9O79baXBPIoL5Z9n9Yp4dATt5fKU6+tGifBUJ3g8nautj3V3vHvX4G/HOeLL
lV0ZAadB62RnWuGNVFS5/PulI2MS5igcNQI8hzOZLt2nx6gBsArioOEPlq8mLg6xm4YNnChczhgj
d4olyKst3X2OZHw/oM3tvydR08HBT+KJrhI36uTBHQ2b3u0DfeHhnIY0dY9vxzZdwFiOPR8Rx44A
ZEmi+7IA511zcvipEJlEakN0XM0c8//Uhxfy0TGt9BINEnEpmcU6fXEbqSPBtHf7eEj9oNhJocQj
A4Bjp7je2jDLuiiiYKtUaO821mVAKlo0aEDcntr9K/BE4x5IeJLO4Nb7eLJ0B9fo3+pGr6R+IfsD
ZK2yzjKmG8WsslveyMouifFyPadVWuV+s9YLj31W4FquLXVe2Us7AZ3R6Gd+YzzE2JQzDuMObkxG
uSp1PfS3n0Iipyo6+3o/hE6wXaK3nCCsfvGXwyYSvb0nQwUP2NanUqnaLUiJMtOaFhKwblL2SCC6
m3FXlh62Gr6rQlHhZy+wXqKYGGRlkP7pVvg2cfPTXcJOaA8/daT9xT2/w+5GTTdqx5EL3W+Ltc1g
+wlI2TS3AgQVmqPPEy4tjq9V6w2o/bU4ceuFzPuGM/LxOweLkC8oxm46ZxaM0GHM3kFwC8L9v1Sm
9lgkD/uNAg3mUc5eIBdTPM/Pg5qMZW9HBp67ZQKygE8Gq6TwcYIDaYB5OQLy1WFmJ9iYF/gwXQP2
oJvDtPNZUPCBdOZZPN4WWrigoqrNPN9aoOjE9r75ZCBLrC8OZsoIceafl3jPh0tNoxaOVgqPg4l1
WKZCcVKsU1n980Yr2yi05gjf2SKaJstPMBspMJrNVgE609x8gsmrCtK00hE/1PMszZNMYE+nrQjH
UU+GlvyzpPQ9zoTJYz6Ro0jqHPXU4x0w16QoDCXKJpP29urlc+zUX8dz6QZfOKvAo0rdurPSNZnd
hKdSJItaH1AqE2xP4yXBJ/1KOdUL6zaJ0ITvr33gr+ckY+aNkzn9VGd9pSJyvkis6ZckyyMa3ESI
E1b1XS9WpNtI+eHplf2xI6mLp0sNvK62AFhXGJ4JrLFRQTwb60ZniEKe0S9qpprvhnGFoSJoLBQm
7rPQDOVOew5KKmRSooHi2d35dR+lzENZIG2jjWAoLtaY4QqHs1Z9JRHQhJ03kYNyop5EjHzdQEKn
i4lYcG/Gi9VoCtRcua34fGJ3dsuqarUadwjmSlwQrMlDV4bigAnrT2DSmpTpmgmh9EltZkYhx330
ikkF0LuHhRY2QN07Cr9Iv/Kvfun8BLEquttu/gUkgI84ZPRN6S+Abq/Z8VO+t0W63mFTbexFY02E
QcnU5ChFQ8JLbX8RIRENCxKAh54IkHvyvhg6drX3C3L6FS6kxb72KxN9fnYFgZLY0m18zBcxoaa9
9+lcDA4bAIzIa+VW3sqUNKISwqElLO4qJzjm//Uqwo6Y+3F1CObiVwbFfD+lo9lrnbM3Q1FgJQZK
17VJxHGvF8/Wh8q+V+r/jnOj4GX81sV/Ew29dvRMPB3OMIZ+5vPyzyvdqCZ0Cgvf3AqI2IOH5/yo
3wFs46TSNZTWjyq2iy3yxI3TzLm6M3SoEDj+UaN/ePmzHp7Y6P14g9QjCTPqqGFUd/1hu7knTsA4
K5/cOLqDjtnCrb6bkw45cpYQaTaRWnMJfTTLuMO9pb79tPeEZKLeKQAcvHlKudGAziu1cws/i34E
61RNg6dRYdn08siO372sE42TW2qCcanE4U0R1SAMS4KPzDrSas7avBvJLXUriJ2PzTUP7V2XF9Dd
A6SsCnkysJuMXos3EGAnh3fJR8pNo7bfgwLieYAWar4Uu55XTmjdM9Q11/6UVEasoV3yvSrMlhft
JNiRcGpQCKgAhnxtvbNAwPTDGScKiVgA8OAo/VFuQo3K1eD7EJTw4fMlM2ycHqqOj0mzMNxtrQ2f
2nmg1TQ9Ir5t1/ZuRWioakpPNFI4fZDZnxDTTa/zlttqMs9AP21GAsPMuemBAzoZO4ZtMDHhzD2y
2CNqfVDoOT3I1/cWGm1QNrH8mjc5tk+vXNWeEb0nK9tdQph4OzxhrVvUuEGKc7adpSeGgkUwaxeY
h4fxbWtSvar1tq6aHLsuMKAS81+MSkdSqxefewsQEZe0M909sQ2NrlsatZ2/UfQPNHoP74nwWPCQ
H0YtML1UbizibBkJ8KOLKV/JeJ5IKfjWkO2sVfW3oavs91H2DbLzn/6PDVJ/9Zq3VVIM86qUWExi
hDAHz8Z82ni0V23zP1VvwM532+dtcvoQON1ZPhEzoFIWPQAOH/H0IakdMJBcMFOdd6ni0XIDu/N+
RLhbX+c0ovCm+hc/9Vx0JvftDxh3uGStqhqlMbdG6bEU6A7faEwAarPbaNl/B6J1RJ8LE9BEdry9
6dQnfthy8oePl6NS0/+mt7YVUkPNYdBe0gTnNZ0p4ADvBNlv6NPfWqXkTlV6X2V/Jwj4IjdQ/oHf
7lCnMpe23H8cdpOls3tyxP6XLhiVhVxxvG2enjojIlEbE6gADAL98vnOkWVh9a6GyaQP9d+dtpJv
f5Yb3LvtMDXzhCzmli+507SOwNtE8BagjUmOZw3g/NiNozFwLKFNKefQ99E4Gd5JGbLfPIivbSgy
2KnYK6Fs0SL3Z62IYycr41PfnWKnzOtlANBXYCLHPjVBxUZ2V4/25BeOlHaZUMtAeXhhr+I1EGYG
825nhfGQMwknbYHV9KqysZI4QRgpcysBRYeQ3iwYTXwfiMRguMWAh9K+ZesSNXA4LYAmjpTBQXNg
RQvbX6Ytx6yKbYRx+hq0Pkf8nZ7zgXgtb70T7pDB+PY5GG72dVWKB3Q3CwkT/zLK3lyH+zzXEX2m
ZqDQlzHDBRGWW0lr2RkVdhyHoXJS1H/cO09h3Sp710rS/9JzRAzCNf4y0h/U/YP++jy8a25AjBkB
Du9eZbgK+qdkzBDzuhGvnTs9XJE4XgHe0LG0m5/E2XRJ4QMaGR2vDYUWJxc0m5JMYpQVgOx2mYJ+
Ua/xWzL1fceaqGUFbz2LsiNQTSlTqEBWTKgH6R/yfZslmtqpmofetJv5qQiA4tfi9MRm7Ehf5XKM
M6K53Ch93Hr9InpZtES1mhfnnYyFAPj1a/oy0hgcOIv4EYyBnz50/WJLMj7W9+hO9aKz5BxsxVjl
eheENymuoz0KoOIKyqEHn9hxLs2co9A2XTg6EMSVZH8R8SXHfZzpbt6XRIfRTxu5juYT0Z+f/d7v
cnRXdHUdq03jgR/X1DnyRq7fAd6osmDzE9gu+/wkbEQslV/Yc8aM02j/UenAMRP0gfUqjsxz1YrG
XQHIBNtPXiu+nkSfC8BcmDfMtL8eUhafXl7O/7rnLGgz7THgi1Qy1ViWqfidexwOujafX2ypRL7I
um4jlBFgTHKFfJQCat8bS/0yusDekTExrbgH1SpFUQhPssozqUfUoNS3lnGcNY/hgFu9MNuxbjXG
EX/SlArXyTcWcpe1mugyTfEYaxohG6jhEYKe3n+e2qTSsZVMlacdpOW/JXxSZ58o1ZBzbV9vwuVp
KPJWLW9OvDqKYxPph0w+Rd8ccHjycSJ4VFdozy+s1zYV8MHgh7R6dUokxodCxSkGbz56GlqJ9lUH
ZsBCb7Rs8sCGyVe73a22fFFU1avCZnL5eNrD0CISOa1yiICdgMUgDpQpBsKbXzoBftgvBYzUiy7q
re+QbDvt3+OKIdbk1SZwkZtfZT8eLl1eNifS2Rq9b+VbQ2sG90TMsLJEtCo7QXFRpFfhbyDjGm8u
3K+c1mQdt579jnIISbnq6MfZEGrk8EZhIfbf2b4peS5L64vF+gxqVtwZ9TlwuxzO+6yq5HQcjUmj
q/0u2qDFVtzQeCsRJMtuik16FFA8k1DTArse23nxypyePoC9qYJnSqVK++isC//j4GaMN0+xt9Zw
VX240rm0FyrLd4ki9r++gfG9pUyk7cdkMTcvqFP+NsKB+4dEQ/e4H3vhU4Tae/FVyEu3OxRIA/b+
JLxFOUxGpWEgUhIfZ0pqYp6TB2CcCAVbEnWv9i1fb1kpeZSt9Jq0CE13S5IKMEjIAT0JtnNDSHLw
6gk6DusaEdWVbb8CGDwENVHV87OO/f/LoDFhyWhuz9C3hmS+N4YLbOp50jD9RgRaz4+zEx9AUimY
X47m7X/Z4gQvMgdco3/vPOU6/vQZ4e/SzdJGFfWcYdqE52E8Eq97
`protect end_protected

��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y-=^��l�yB��O{8�l�nc�:�=UBZ�랺��n�	��A��>x�Ou��ΗEpk=���zCA�Gk0T
�2��K��/�9�Ҝj��,�q�/�4��*�^<0e*gG���RFi3-ē��N���d�'Ӫ�Ce�~<Pk~3m�KOi	u��_��az�d׎�W�Iu=�/�kZ��,IQf�L�;G�����A+wժ��b�#����:<u�����lN����ƌ�zZ���[o���X]�"r����:�FߕR'�!&Q�ed�t<�H�i���1Y'&�#�����;��t�t�M���=,�Ѧ�?�޽�Y6�I�����0R~��|��f�/9�a1#S{{�ŦO�n�/�N�Hʥ�>����f¦]��O�}�g\;L36���#�DAC��eβq��Z�^/�i_�&�L��r�۳�����'�x���B��/�X��Xd�@�G3��tc6b�8zf�]$�����F�s����6�����e���l�2EdN]��K������=���fy���yDi��'��ugE;K�!��ne53K}���>�3ӄq�Mvg�U�y��������$�Q��dd��e؃�=a�tލ{����p%��A�ш��	;5ꉕ���D�s�C}8j��D��#.괬�j�;���8��������XB��-�O=��BX�����}�LX����f�i��X�U�|ue:�7� =���qϒ���Y�=[6?�YB�GR��Ji,�r�YƋ����k��w{�T� y�0a��hb>"�=�e��jk��p,��H���q�`�6m&��+��� Q/o��-�2�K��pկ�f��p{+^p��_��)���F������n���oyo?`Y�#T���~���|���Cimj`�@��y����ᙁ8H�)�B8����xO���ߛ�Il���ܩ�����zqf+���ׁ�\to��kb�N�ϩ�,��S�mzvf,�R�i�{F�����,�C�Іpf4�R��c����*���l�0c��:"c��7����Ӱ��"<��踳M �>�O{�%+��\t2cL�A֤f)�HT�CZ� ^.B�l/���3Z.6*{NzԷ�U=�8� �Ok�J�9_��y�o�mAhs�.Қ�.=/}40���٘���0��1䛫T���ӑ��!������l]i�`�oQE�
rn�p$;���� ���8��EN�砵��@�Tu����Չ�KU�T���f��شdÏ~�@���{����j`+���p�"�'�H�����=��XS�������VX� �J���ݚ�^C2�7R�?\N� n���������:<M�S� �H[�P����R4x�1�=4%ޫV�.�z�L�����F����NBЪ�r����?���T�T�j�\�#џ�t�֥�OiU'�.}V�pȚ��VK�a���2��n�k��
���zG�e+��ɶ��R3
=R��N�Goi������ΘF~-�R�CW�9�gC���}�s�Zg^<k�&��ja��xr��:�����,{t���Saj�*^�YP�(Nݫ[�`?;��l�b�Qͻ�VۅI��7L=U�u�UݻrqPm���x��� ]"O��"��=%��V�i�D#�Úk�-.�<��5�v�|�^��)���k���Q�W��(2�����7^q���3Ĩ�4�d7ժ���z���d�űb��b�OZ��`�k;U�qE����kh&!���B�r�6�=�v$�V�VY�`7(�ta�����5�Ш�VÌ��� n 1f(z� #�-���w,+Z;r]\�m������棃iZ$���c��ޙ����J9x��L\������gL�����?5��d�W�x�b2��8sCaoý�`)%���p��1R��Aـ��&�"�}����?^�롙H��I�C�}m��ϢG�����GY��p&M��>,a*k�զ��7_(A;�K2a�f�;>���煨~���b08�.�GK"
[�˒��_OE�Xy�\���L��l�8�"���u��"c�J̑b��	4�d�����X:oC�f9?�\��R�}����w��m1!���$F����U�U�V\�h`@w�(�(?gJ�#	"v��X�M�.�'��4B*��s70��RxWn�,�}���O!D�Y�8�����辟����j�!r�O<��y໿��M��9��T^B���d۝$���e�	����,�䞤Ua�:�I%
�YfT�~����I�����8J�ឞl'�}��6m�m�k7����tq�ە��A�����r�u�t��u��{�;�q���(p�$H��@��GtE#�5�_���"���@�n,5��bF�7�`�_S��*�t5��T�MO���L�{k�j�"�`�����S�����Ok�b>��41�VW�Q�a(�/��w�����|�h���#��i���K7L0z"�ӆE��r��d����ۅ�ŵ�.1��w��۬�a�PB��?%�Gz�r���r�Hc$��όN'�~�FS��NWj5E�U��n/��`���t�Ҥ]�CP��T��|�)G�Rc�64�_w��	'\�ae*�b���Ô��N��@��-_J~����;:���ώC#��z��6���V��d�0	�E�	�ş"u�O�oVY��y�=(mQ�}�iv�0�? �Gɴj����IZeİ����N�q�4bW`�'�ee*���l��{q��I�+t�M�i��z� N�n�P�|�#$���X��/�//�۟wg��=��U}H�m�wA�
��8�H��v�LC.أ%��m��+�2:�f�_�nn�[�;��Wg��L{�����������g/˂0)EX��7h����c+W� ��t!8LVk!'|��E��3$�q:��+sٺ.��$��'q��w
�ߧlB�3k�Lg!dH]'�(�Q|:;C��R�;��ɬ �6W�8���|I��xw���V'$n�í���93B%ϩqC�� `(Ch��~�$��;`��.�{L���)[�py�~�8�������1J��o��d-N`���Z�=����G�붜�.�,�\O�M�D�J�m�����j��q#�0d����%�5�T�y�Kذ�3�#:�#�J+��Ќ%�4Är�Ո�kY��g�-8�6�����W����t�a�V4��'��Q>��)_�ꇹr��=��|�<����މ���Xq�C�ϴR�BY��:�,�d@����،m��π��~���Y���m�#���lf�~��R�a�d�%��Cm�qf��s~^N����n`��]$�������;´~���2�����f#J������~��1�0c�o�=����yo�Ⱥ���f�\�'ss�4[�_N�ؾ|�i���=5�o�%J�'�"���e"�d�<՗��w�x��}t����M)DC�YS������[��V#s�B �����12����5�y9�B��Wm?�=�p�#�J�RF�u]K�R&�F�qb�˫�.a�d���u>-ۄ�p%��d��rk��Q��k�+�Hln�qYt2�j
��z΄k�?�C��F �ͽ�a&�	��u�h3�B&`�I�zȱ�[��եUQL�*ɭ�r��dU�;:J�D��N���yi��u�Mڶ�w{^�va�63��,���O{���.�L{ݚ��-�e���g���`Zf*��w����6����ɧ���;�%�+ػ� V�ڲ�7G/�Ë���,��9���x:�6}�a�rL���p3}I0����-L�3��:ߤ�y�ָ��t��#�t�]����b`�d(��VW�䰽Nj��Q�T����+f�0�.�<� =8�(��d�q�|���.��E���ZOL����+{��{7RC;�?,(5�C!ȠX<��V�����,�R�u��37�Z�@zK �aon\Z��r�d�c�I�ط��57�Q8�v�3��<�_ڪ���j�1F��������<�X�[��]�����{aFl��XU��t|�k<���*t��U��K!Z��2~��=(Ǫ����"���[\ˆ��� q��Q<0��Q˖r��Ҿ5�4�w*d*y�b�^䕾p%�G�ə42Y�j��q&H�Cv@�B ��_��f۲�U�01|������kL:�����S�N\˫�~�g�hf{iڣ�����+�ƭ�Dr��[�В8�=��r�bL�].����*�EE	�6 ���|���	db������qՂ4��&S�E)��8l��"n��K�����P����VG\ ����֑,��[�Ǘ�bnT�'�R~���]�]��F����䤃�K	?��ĵkQV�5I�t�G�%À�~1����N7��0Ͼ�A4W-��an��(	�Ib�3�%Z�E�t:\
h�R�+y�����W� ؆$$�N�D�<aH/��Y\�]��O�Y�.;q��L�	q��t��ͤ�� �;oߏ��|k�]=Ka��P~��| .]ū$����F�1Tm�6���i�@�FB��I$����H��Cg��Ց�a�v��l|h�3�6حᗉ��`�O����e,k��H���%�J匏��+�M��p��RG�:��@�?��H$�I�����x.L�׊�]ݤ�mŝ���27z�I���8.�t���-P�LH�E8�$�Ɠ�ܨ �wQ��@1�y�CH�����lF٣0��C�������w�
B�`{l@�]��g(L���OPZ\^��{��آ��P2t~$�ҤNc�~,�>hQXC&J���Nbu����A5
y��1����@Ի�t�N�5�MViX�<���0���\����� ������L$�E����w<I���ʽ�� n���*���ʜ��،���G�C����FJ�ut�!��
�V�&��,�r�#R��C�o���GNߵM�e�4�+\�ܱp��M��_�? f<�<%�т�����0��-�	����Jr�'}[N�Wc&+'7n)��_���t��E�9�>����Kl�Ktt�7�����t"i�(P�GA��L��&�u �`�S���l�`���B5�y� ���t�〇c��[�ȥ�S����z��V`���Tg���(]É@) Ì�ԝ�W�cS���}
��m��,Oߦ+boc�ޏ�/&(ǹ���w<�sޫC�dA5i�f���^-r@���|�!��NFD�6.v���U%�
uk݇q.�:�4;~=�+ֲ�<-��N@��ǈ/@�^�FҮ<}��Q�s藒n�ĝ9s�%�y!�D���9���C��-\���u����~߃����<S��h~��� �!��[s��˴���O%�RFȆ�++l������Q����{v�0<���+X��9#����LR>�m��'�Ӟ[���Q|ʌv��u��a��m�#8�A�8�K�1c.��t2d����7� ���}�7}�;/N��ke�J{�ޟ���'}}�>K"�1�f3d$ Uo�R�Q���[L��<�Gz�e{ba�y���'��Р��5C6��tOeOvag`Q�PX���o�]����~Xk��5AIxt�HܩV̯y���)�;A�ӻɹ�4���o4�j���������i�I�d���5�P�?p�ϕP�NE�lf`?cx�=#�Y��~B�x��X���,Ώj�M���VA�{��X}����[rWs����|��ʹ�0^�
c��50�▄��"�[ N8�'��3d)RR��Q%��VRF�B6���u L��sB�����`��z�9�j.֡�p�'���Y/�Tv6��=kӕ�@Pj���Lm���:�3Ͱ�{�;����_1���,�R(�̚40�t�A8�ɞ�z��-��I	:*��Z�	�����)��+�#	fAs%�_89 b��EǎK9 4T��diYC
���� U�X��f�ٕ@��3�+B����[O��BP&�'�A����<��$�:��G�m	���3��Y������-�K�!1�e��%��6�H&_u�옐sAe�;J�Y
��qr�M�Ȁ�1���Y{Vޙ5���%���-m����>[ҁ�q��
v��z�,�g	�G��eWݰ�t�3-4X?Q"r
0��i��.?G/���sWތ �!g�a��k�9��+.+� AT h9'�sUcy%N�Q��G��Ht]^`����=�;��"�e��[!�1[R��؅��%��A^�a{mF�?�*���Koen���䀘�sʆp�JK�i�w�:�RE���m�Ѳ2��)$�<n���V4k�vP�
�L��G�&�9ڳ�a��J,�����&ڏ_mV�ݟ����6�i���p��M��ΰ��6�1��'���h2���7[CH��[T]�p�sR5~8-NA�1?[���u�c6&���K,.G�)O��F�[�,��G;������9�ʭ�w��v ��cy1�P&�''�tpfd@ˇ���Y�E�����|m3�2B��x�5�AG�#=��%p�	{p�ɡ�xm(2����܏�m�@�L���/��o@Ѣ7K���`�k��f��c*g��G/9XO�p) 6F�����}���9̃f�'��b���y��ף�5�/�+�ǥ|n�)�X*W���)B�}�F���K��}��?j@R5}���Ń~U)bB.��������G���9����<`Iz�9�cb m�]�����,��Qze��Gt���!�&�e�=�A��4b�-��r"�G^��𗶳��O�[�[ƿ�CQ���9sdK�T\p��J$��P<���2_�Z3�n���:6�}�^*g�42�-�� k�=�M�?ǿ����ĀBVB�gZ��x�K��TM���;�h��q�4��7mw%]�r`~N��^(�b�h'=�2㻋ť���:K4ޥ��R�6�'��&����O^�/������3���r*�ܠ�~��M��f,����m7/s���:v����n���\7ܟ�+BaODB1�a�)_�8���|b얒JQ#�ig���9��~�6A�E�!ס�{/�ĐȺ?�Vq�!�a�]�������qlΞI<�֙:��0fS�&|�/�p~��"G6]�9�DBt��u
(���\�[��Ύ��Hjw��Ki؈�,���c���0�$v	y���o���{*�!f���{�������Z�F�-z�+�mkۭ��BK����B���x��w%�8��|��(����{r�-��I?���Y�%� ��_$ׂ(f��j4Р	��+&�(�bN�c�c?ڵ���45
^k=�Vb��=.��`џ0 �92/����a���ò��z������sv�S5wr�U��xF֫xݡ��;i�:���2�7!=��֢v�.e.�Z���W����րE����f�ۆ����}l��؊�_�D����n��?,��ϛ�n�ťbd�o^��1�)�(�a�?�2{����C�aK��9�$Ư�y�g-)��$���h�I��.\�K������.�g�����ڮ/O� d ��PVۮ?)�L�A~}p��KѪ�0>Br ,O�md���U�w��r��Fe-i���@*[c2rr/�5�v�ѫ����I�@��L'du	���U�Mm(�O���>�<�-e���S��	�f��h*\(�;�	�{&j_�-�����j1e�V�o2Jf�Tۓ
A�Z^m��v��wZx �E����{b�I�Ԥ��t��"ofB=�fh�{���@��@:6�j�3>���Ӌ'w�%/���j?Q���~��_�P�����Ab'uܒ�:�drq�����ɱ�����l�x��N�6�Ӌs��H~,����bt���]s�xЦ��y���럡^U��pI�G�1�ʆ�H)��N:����V��JBɣ ]���Y�"��սmۧW{�$����*��q6N���akG=�v.Pn�� ��q+�9<����8���:�@jw�D8�3	�o�H���m�r^8��yB��6x�V	�dЋ��ߴN�ߪ�{����=�El��S��!X��8�UG�dGꘀ+�
�8��y���x9ޖ�>��2��w���ع	��#�U�G�a7@����4�����<��@/0c@���'8��}�Jx\����t�ز,������$�9=�����ԈP��hhR��
��+��cY��H�C%�3Ǔ��]�dt��ɣ�*�	�\qx���zht���ΡՓgTWg��MMU�l�J�M�)bZ�Xĵy�a�&��೴��@���8כGO/���k v���G���u��V�P���K�m⤇�Y�U(m�(zV3t�ۊ]��Ą\�/E��d��a��$���JH�8���ty�)1����	� ��D���3��1�u?�{!�0�ܝ{��}x��Mɖ�"S;������|Y!�"��	���g�:\4-Kێ=g�v�<b �.��}P�S�qz��}������פ��^�r
�G\|��N!� 	�@1���ze��ʴ��|���u�I'YJ�D��Z��P�?��7�H���.� Uh��mn�Cdxn�:��9�
t�ʣcI�q��Ih5P��b�!c>��q�M-���?*��S��(�!�.�s8d%�>@w�%��e�N[۳�낏'(�(�߶� �>c�A������-�0<��y��kgc��4#�0vs��^12�wE��A���4b:k��ͬ��3��{һ�Y@�$�Ju��%�v'���	[H[��r���>_ƩĴҴ���s��1R�vj�/��Әy��&T{���ʡ��e�#'ǜ�wޞ�vA%]���\9�r�~`w����}�||����*���D���ތ��gW��!�8<z���}�3)���~c�~��P��Ů63� G]cx<g���<��� ��c�W���>�%��u�x�$F3�>�{Em���[Zcɂ
�%ǜ��X ��Z7�R#�y�B�l&���|"(����p��`�|-�?/�!n��F�F�Ҙ��u  ��p6��������}��)��<��Iu���g��_ h�"����9���ELEV.�3�BZ�3�$e��󘎹����gxQ����?����7=4��,�]~�N�l��;�n=�N������6#VSW�<����{*;FSS[����機��[AO���,����[Ǔ��S�w�i�b�� �\�q��٠����f�#̓v�%������Ϣ~h�����fD�Vv�����s�&k�24��n��
�F���w��ҝ��=-�&�x�t���Wg�w�����ћ#_Y"�s0h}l��]68��3.FK�#�H�~I���p���o�lc��"ITC��@����]�Ě ���f�hF>Ȏl椔��n�[�W^���<4<�~�GI��#��b�y���Z�on�B��D�!��wk���=d��#:tm�\�B��:7<��K���	T�h\r7>��F���S�����1�����-�q]�< \Zc���{���e�.��2�����wW��,p��H|%����������1R�^�]D���q@��f�l�����=��*��:uқ` ͠n&�,#��$��T	� <��V`�ޙ�)׆N��a����,�L�$Z�H`p�D��q ���q=�?UgsaS���Qr7Ƶ 8땉�X��{����/&�ܺ���6�>;9O��<4�>;�ߊ��F~�1�4��c��u�����XT����s\���ԥ�
}�ڝ��[�^�ԁ�×�b��i��J�{�j`g���[�(� ��r��X��H �Y�ER����TWm�m��$�B	�l:�1���g������Qd����X(^�����b_�@H@���kg4�㚊�gK����RȵB��.b�	���$��u�h�&�7���$<]Y?&�D��Ʂ*3I�	r�8��K����Fn>r87��j�{9�2�ʷ)�"޸+*��G��S�6�(�R�
O��WI{_m���9P_U����5����'�|���`�| `���.�~�;"� ΰ��Ʈ�	U����Z��k��7�˕�sX|5d\R7&��%�%�n��R�>I��R��
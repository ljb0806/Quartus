-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wsDSYBAZNz//0qbUTYIMdrCJZce5H5c/F6YTQaFKQJU9NqxMbsJ7q8e6Ree0lwe6LFt/C/XmRIbu
UATVpB3Hr0TQqbyG5ZDnI+CMZraExDJ+HRbb9WENRQeyim4eQLMretZfdfSRtC4BGHCj7KWNWmSt
waLXfbvJ9aSNPU1VByABZa++w94ng+FDEtZyUsvnJg1f7Fcu6ePYSXF7q8YZyQfgYutcbwJERS3J
l9fOfBn5zTQQpPtfB64XCLd9ib7/73O1aoUdHKqfh+zAuQ3UzXjXjJWMKhR7J23YhTTzot7C3QMH
r9/7kQzi0wK/uWmdmLv6dTj8ZZCIeuetBfprIw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 56272)
`protect data_block
j3Rgz0OI04zi8HR+GGb1a8Tq6oHqc+x7k1nhmnGnxURmenOMnXUk8K372Fbi1c1rX2id1GDp26TQ
5XrfP+A1gZvjC7JlQQjREdgKnQJYYkLQ2W+ueKhbny5nx/X0eLFjX0FTYXaxSVD6UPPXByuDutix
RA85KSK6eMKr0LB4dILeiHQYsZDNbQZOBbRcFxacmG4t8tDPE8ESX1EPhH4GV5KBpi+L3Kprop4h
+D4D02uwZnROjBSFPdoHDah0Ih5ah4UzT85Ll8OrPztYaJ4DR5+1YRlvh08h4kU629ZXFcbFb+eb
n9qXP6Q06jUt/gxahseOm3kKXKPB8IJuPCQ1dCG9TpQKaiTZiTQkFA2gzfAHqUd9cnpqprbeVwEr
S/MCVLvpu9z1NQ/2b/FsATNONL23s0aucHJRa8lzbOL7OHWdtzZfEEH44EYt3uLejmzvWCjKbGbW
+lRQc9ywq8sJkc4sF6aeiQcNGRuAPe/ShVpVxDLj7hME8shPeo0Aytb6WsBQEio6d9bq6uJiE5OX
ya8+IZ4HRnG4xCthrTB7/CxYHFpO3L/vtjjeeMjHNtbsvzTcGutPmaA8KN6IShNCf/C0Ppwv9bv8
xPrhtX+UbILZLJnprO9fn9DXye59JPwT1ExfQZ+IoGmdliD1F4RNmCraLr2+1Z+6BBgMM2oo1eTD
o0SMshFJyBg/ClzixtgXzxDUPe4uAOCHpcuzXorXxcauD+K9yHJqNW+NPExVPNCENcFLj9vb+06V
kvenFPOrVbXsU7iHrEogiKgWoChUVWZ1DnazCB+jBmFMxiHbX7BqcBuWcIVujubG8KSHd+UTIH6L
J3I4MlTDabmOXCeM34XCUO2MboMAmZIC4odA3dX2beKUtwEVdzHEdsj/GJWhz+aagkkSZws3uRES
yJhmXTy6jS9j+hKx/BoobAxwljyu+T0SoKZWPp+ONa6dEhDCpqLMKIaaVjP602Og/f9OoJ8kRUm5
qD8lZLkJoPRP2uqXne8aUPszTd12xvJM064cE1JySNHfcU6V2tKCEL8Jcxab+rh8ORzIW41F5mJY
MzV5kfZuyGe7l3k9e9xdPg9C8BukAgp/qMGUkJvgWbEF+7VsJids3pwrC/zVKkdsXj2Rht0xcpnc
E4muptOlgHthmdTmGJt3aN6fAVczGb8bDt9gw/FQhNjIz7YqVqyUdTCIjRRuEPyHHwuD8bEma4tf
3tJuPszHJb368pe8Ols5fTFiEOK69nj4M5MWOW59xWbdFukYCblSo76IcB+k+TsDje42L1CPYE9E
sPxAwq3ZSuUSEkS4EPqpaQNWHwkC7YqLNjVkELNFHb+480+ng86RUMOQsTJRsuQ19z3Ws24E+6Eo
okIqi7rIeuYKrvQ1rv2ocLmu97l2UyhlR5ZW4YHJbRH3iWlQDYZdgqW552Pll8/y4N5sCMLX4RYl
UXgKyaPWCK00xwtqAwtoVA4ASMKciHp/PwkAdczvhw8ceuxtmGXrldUYGLnBQgPs2kcFCp+IrWLM
C05FpNVlYLu0Jap1uEn1VowPaXdL2qEfCvblwp6xZ/EuAnfISdjk7LJOZBPcRYJcgyhmeRfxv6mz
fSlND515BBqGk3J7Z7lxol242Of+4Y0gbcC3FmqXXDTSEGwoIDlsS/voCxEmMVR/MNbjFXLiXUsD
XWCArUO3PLJnc5hMgQ6gOX1A2Dv083bP1t/XVCBCQysG0i+jGZcfFfCVi7s5wQY6+GBmBxKbtv6A
CRBdKW8Y0YAmc3R285BvQI4FZbxasBlzT5ZmiT0evw9cDPmlAqWO0TmPYy/Li4rXh7oREzZ3aJw9
zaGCZ6220IHi5/dMa6AffqEFwFGWAoqT2F77Je8gMfRXoiypS8HtknB7GxMQppNTd38fj8pPlDxQ
Ldedl/D6xiKVbtruQ6eavibGNQGzaIZQCpEaZP41VCPeDQV0E0J7EjaqQNcli+acHWVyUHNLrhRQ
X3WD9OAin8Q5UVf2ec0KNvBtqXb9/ntC/f+z4S7Z3WlfIGOfSMY8lavd8c2Ynnrb9pMn9cdpWUY+
2JfrqJFJFe9QHkC+RAWn61xhHf0urYUz7SLrHQcdpbJfA6BCFn1oPrr3yHF3wl6zQo2ZZ/Q9lfaf
tRF2IFT+ZggVJ6PLg3fpH4B55jmE+YlfMGd4a0zyoRLZpJr4mSjrZFJykgzsx8d75Sxlgcj9lsMm
rA/c4IGqkFSDz4zaQb/rmSHE7MRswXR0lQSdgkGdxi9w/lQ2Ikrv5LJ1wv+/vShCcdq8Zv38QUng
ISk5BRLZrh3Y7XygiRKorNHBZ4gjye1JdM1eIkLneglTpeyJlCicoI5wIfl3r5ioU5Hhx1m2gCSI
bnoC50Bedn1WEF6YwMpfhdi1+dQts4wrhSlLpR2m/S4gRxVTiUCk0e+xBeB8/ud6Kkjof+86Ve57
QB2wdyyfbiFbCjicL4F8R+FXQeZ9OGhwezE694Ev1CBnUWvxz4IoXvIup0a1DUf3RLV2FX7nrUGl
oRMPEb/InI+0RUtOusLKK0vQBx2sAX5z4+goFVpsvKZiL0fQ2DqadcPdy7at2dO5Lt1O2xLSrJiq
/oz9D98YJNn2XwTnjPXCwB5HlGjEpOKq5CrdRDviJ6EbyLi1savXMZcy7+LYnfUXbsu0+U7u1Jq/
+81NCHHgGxjV5W3GmNE/goCicWUj05jZphe2/orosdLOCuhAgJKT8l154oXqOnfey3mxoqASLSSk
hRcB5dSOe9yJLpnF6MQOhKcjj0WtGQvHP6GWNXDo4BPfZfu+j6u5aDFae3zF5cs+4iK4p3Xa/LzN
oRSsdz5Qtqap36gZduzPy/4/0O4sNZsWffewttas8HRbB6owXsSLuILj8nfRRzoI12fMtn9DRzFH
nbZV1JI3qN7VdwbgTXIMlymXDn41C7YsPa2M5jbgXpV6mgZJ5Oi/BrEMmGVEoE+Z/msN/qqmWm8e
/6oUAthY4reUeUqMZ1GMhpEtgtKYhX4B9r+++ZDNUZXxjg/mSlHdgA/DY0emYP1dq8RvhVEWKoPz
bGe3CPJQY1gWwCdpnddtkuZT0K8SLm5vmaOR+pBfrg2YCp/G9dw7IeOONKFk5ZHC8vuUZ0gpK+Jm
9f5hBwfPUBSm/ILG0AC2EiT4wmzwGBrqNlT7YA14crKZkaj9OsK2GKbG2k04agJXV9R4Bem6NfKO
3jdU1OpQ1qWe0tz3EjoJ52ZbIKvfeBjYMfLdDzZhEUDgqx3YWx46KEZ+h4vnN2uloOa5F3GEjRVO
ki5YICc/yFQWHzFDytN8OC/fqhWKaOZInMEZhFB9dpsOb2Mg78uamJT3GcyOQxHoqavlc38UqC7S
J3rBgjKgae93lr0aAD6GwFixLO4B1rKxNzaKSEwZ0IWEFfBYi2LGI/aotQRpu5h0xvqH4rICxhLA
h+ufomagoSnQB5l0ODNZykjFUcVz+sQOwg8iJRcayH/2ialDTf6gg2SHOlvMv6tRpltGRludHO66
jpn2B0z2J3NwFdX+FPquVxVmRrA+5SbCcj/ObHyhRGkOTqU3wtOrYqdftDnKxZmCnYU9Ow5h3GyP
rO1pO0rUaz1Egmos5o4p/7T/RbBTWNRoPNWOvXIgDlJsRKIOTiD2GOghgCtv410WGHjxo4inZ6iw
AgyiYkuceyCU/Y00rSbM/5stSmZ42N+DQBfFai7HydswJHH9yBAxZNsCmpl9Jfns4sOFY0FSEapk
8R4ciBhp4MiJLRkNks2KPAYA/jD4HGdrWGOBNrczI3Q0eZV9DbnvpzN7kuGGZshL1XNsc5o96AV/
vzzFDdq5f+9hs5dj1WzDCnxrwKnSfevaNoF9wopv0G8vAzfBOoj7iuFqHjs3MTJ24S5vkKmVv77i
VeM9Y5GrWf5BvYHbpPT/lcxAbVdhAmYfQYlCJhyGhnkqzNNil5ITks7/KYGPWBQOATgy1nZlFF+b
E//WhMA9LSYPkz0n/iWhHWEW0Zfqzdd80hG2FnEweJARUyHp9QPEmCm5NfgBTfO8LSXVsOkbh6NC
CJkcFDLwCufWwWZEvntc8P0ZFgNph4kf/0tcn8ave+Reh3/jJU01W/lFaa26gJNFyrL4EecBkIaP
3Hx4iMAYFDpIKZbyGdFtdQ34XQi7sNX0Km4ZJ6x7JZJa6U9bfb0VLtNpC/PklH73WJMsRRlTW+5K
daO8WcZQhymm8wP8ZLGr+320sMRoqoOVYTri3prFFdLK4/GcMCT+2PCK/GU1XXO93Q0RAwNwhxpf
AElvhx8a0P7MwXsSKfGuQWiwcR//ve+QIgjel25O1wv97niFHAScs9ZXBfK0zq0+Jg9QA67juGnF
mmPfUiULnKNz0kMr3un/Xzp4XIEGY5dYTf2bMeBJRp4Cj7iBMU1SO8hp9LJWMDWa8f2iomQAPCTI
UciEhSBktsTGGc0oNXeKuCsSbyhit3hq36dsZiqfXy0gTa3mMbc++XuQ2W3RyfUwLiWQTfqDLmj+
RzXmOzQ4GOXlwVA2r3lz4AnM5hC348/FHGTQWnwvePL6aE/zu8gx1QCF2OvWn7up8h/2VdlNA+J2
4EYw7mBOHbMlevN8E+phbi/79oSOY9E3ncNh70Dec2EKT38tB1kXuUY27n1YlJkzBLklBChHY695
hx7m95SLb3ChnQwwdWT8HQQci7OaXuU9ztOQU5y18vtUkwA+WqRnxJxhMGOctQmkHh5k2V1Wx/fY
+0IZLQzwfHbrVI3QzdsbQDQi1lCJgq/kijhMJXyNRmRlfZ4tvg2W4PH35uYNaA+AYsA8AfQV6HDX
t1hyD1ZSZEQ8lzuE7UIY6hPKsW/EdbEp2/4l49PL2yHKgsDJhKwknTLhqsIyk1RgdqEJh7o2Z+od
X4n8iM7GBiIlVsphrDSsDlhSz1I0VD34UHiPofYGnrrmIA2rd5L7Lr9POhunTN2ozrncCQE6bf23
ivWWMc3O12gO1RJqcmwQWIzBL9wJbg8pPvD1slQnGWQ+dXINskbuY295iqJm12PmkEI2G+sq3+vi
UlzCKVqfcyRGK7RpopMtdWUSgElLwlTZ+YUlWkgzxpjtqN0zgE3T76C4wr1qj4bDf1y2yGrXCUyL
DeRwTkSsAQymMriGCww8sU9bZ+epo6eN0Hjrc4Y6O0gsKoLRX7JutADD48c0HAwT9GfDDVUJ1xzK
m+bXNUVCdqbqwLBw0amBXKDRLQgvLOJg/lLTqgbUzyMOfJoe2CFngBeaAVQk+xyHHFTAFGSIuUTy
4hxQ8WJ/vsEY0gQEs74Asw0dGIHOtsZ151u4xuKMAYlMflI39Jy08/jHOCjRvyUOQltq2FOnqG5l
GxeASARpRZtiQFR83VNMqxLsO1y53XF+lUB86gV+w+Qqlam4ubLFepIj7PzEG5CC9DafEN5xk36u
iFq9loTmMSWi9AY9dACkNkdg5TSmR2UKma/pDj7oiPw1BDUS5KUgWR6VQSccplghGW4mQqohCKZD
0ErrhPQE+QJDI0TcTb85BPwSWEOSUNI2RuAnZS3mTKX7rFO9I/FJvenln+rTMRbvloEJGrNKzL2n
nJeRQaYa5DaZLOm+2SGgaFdpiu3uM/PcYXiUAwe7XrDWzpHxs/EP464RoDmQeYOqVKpcAgs6Vctq
TuC2KUNvAVDtOcCu824xfvq63WtIQ3//Xm8ris7F9BkOQWG4Mxdj8+2XrybF3vZb1ZBv8f3pdt9E
w4Rz/LpFScsH4ddK6VKKuMH05l+pgHWjloStyvSlI3N1GB2OCwiXsOjxmMyFMOkA4Ood33UnnM/e
AjLS0mJOpJc5JCZGh0qLhdfjgzY0sIRWq7sZOdoZbo+HKCGHgwl+thQdO/1BzC6WZym7NO4I76n7
Ikg/6790Cd8js1knGwJtRF95x3RDjtC+uU0ByciRC/Dx7hg62v8Smsite4qtx79q7cGWNSsTD5VS
SLdbygxWmBv2073ElB4iXo7112jeVEbW2mYJk9f5FWimyFMldLSbuWEcpzf6JgpFG7rQOl9/+gXk
guecLClE6d9CtCP1ZMWf537HJ2vFXHs1GWKPfCNC0hU2WKmqv3mIKW4NbXcbVCu3955aOyGS1diS
Sq1bEhR/n1MZmwb+vzAvimMcadPpQDrMZlfdZwFsFeq0DaSSdzuyUOll8IImBJPspXnV+Tt+beRw
q3whH3ufsW53C0NhzGXuUmxEXbX0uF/Sm+7eZJ485cg8S3E04N1wAHpEFgqoX+y9h60wAKFPlQy2
RCsONlz7+kjLjfZjilQYspXAsNCbKCU0Hh0XTL6NLrURi4yoQPFKipMICQv5HSXXo/m0OLHGTi5T
2fWc7dATvfY1uTBOf5p1TV500I0ctbyrIxH5OzmgmVLQyiAzF5PGB4lvHV3juMPKNpU8aL6zcuct
3B7lnMivU5peculj4SvqAuciUKnLt5xQK/LmBuFxpvvo7v6pz2aiSNoyXEQT40ANSeXfFoC5f/SJ
YdelwjFaKttcd+vybW3SyQdIeA9Xskp9+gtLJjnlul/w1iG2YWPZj8Rs9VLYMQLwXBOP5AzL9HKG
3+1ti0JyUiFpmqnLVXKH8pJwwecjKybtmDH//pCpXJMtm0nwwvy4qW/v5t6DBxRxtPsHHl6DS7Be
jSFKtGhJ/sQQqLFfqIJVl8np2xPIQKI94FxJXI6lVNHM/6r4Hq2aG7obzGQeKf/9h9sdWRS00r4r
62Et0TKEK/OnC9yxxkEX/zou32UMd4GB45X/U4fAgMQHDzK4n6ju38gpdDNLavpsF0YCFq9YC/e7
dcXXWaguet/4dl/YiutNJ0KcbCS8l+L+8ZsnA9djD/sUkPjnHpgxsk2fDpW8Qf9BrVz1gvOoqTwl
pUsgVVCFxl4MSNpHeRY9pFh30Mrx24rRhYZVupAnEsmHcnZPKmrigrDQ16MH356BdQ4f+3qj50PS
rPy2Kvr0rOKaXoRMlgpE72T5tJzqxvTCFKrBqrICRb9dDTZmEhNlPe/8l2OTFjj58Ah0vpzCoE/y
02GzLzDMbi4XXJWpb6n7/cWTJuMTg92qe6SqiCI39pf4zkayQchSfmp6J+MNcpm0JQhqkglzfp39
1yxn9KOkZsNbqqr67+yGLYN2LoFUc9X3NiTTjGJ2MtqyIcAoaCxr792ZQiEJFZFacCE5THFjALyP
T/P3rQF4fAR5wJuDmaf4ONhTqb5+v6ywRCjgUs80b9TqOhO/Xnx1bVHZyQI9WYr1s51iU0Szc83t
ocd1TdAmPVXxKK/65NuxHZhdfakaROFFmXsrvSxW5ArdnY5CTwYwL68yTMaenuso+DSwFXQXdz+4
cNPPERT9A/9cSYWlez/iDGiJbKiRYH3qi1xeblGwFX41q7KZT1IHr07HYHJ9RMNktaO5RlUZ0zac
2H4ZWqPapLZ/K4kQPTCiNN1EEZP0CXT5IuUBXIW71ckemhyUXpJltxSdMiJOnvyUL+J4EeHdRa8s
tQ/9VyGwx/cogLesBea9iEAmYWlQFLKg1ZWLERJUzYrX6EERI+TVj8Rni6bHtu06SDfEh8WucbLF
/5LdGJY+G4j0uJZ9Y3iZOzX5AnxXvEFqOYc3/gzh2sDnVo0pS8lr4/U07Td/6NdWyE7A/dwKXW3X
V2+lB1/ltOyDZDHgf9QqJxPc+Tk2LGuOMIDKO40vbGXPEcXJu/RYLhH+LcrCN3HdIo89TrRPVWpy
lvOqMKZGUEuk5wl1yPMtCsSwFyrfmnFPFZrv5Zl0MsHcB30iPV+hWDFAQ9Retk+koUOuAiOwg9ma
PQqIAKhsb00npD2WZPAokUhNUI9jx5W36rZR8MrJeTcdxTgB50H3WavNdWBeshbz39aoTYqis+r2
KUcr/kCYyG3pwJ0PxChWPEYwqlNlAseeep7oG8pxMX0KcYwp+SUaHzHkVOw4237J2h0/EHoEO3ZN
4tXW5yMM8WQgjKs5C05XO511nsWpiRYYqlaVssNZgehuNxc2I9SK6pGo2jCA8nyG5oaGl9Rpbwe5
uOVd+cMC9HhuSJ8JUf7lRrJ2+hguE3Vb0eLhZW7tg598xaEi1o/ieq0usuV4fijfOBV7rIibip/f
zvEkDXow9fNAPs+SDuG36CgV3031epXGIZ8fv+TlQJ8+IsQrYztVxTVtJhk45d4ueOouo+kM32HC
iqnG5D27it8ibBby8826CWA2tBw4KimjncFLKLdUKjl7caQy7KfzJZ1WENkxSEyCr08/EN3LHNXF
qZic4ozX1sPockOz094owuoL4Snti/m8S4DO0tM3j5xFUTxXxzmuCvCVjyaU/GM7DyBgEh7qAI0V
jiLj0n0lNlMnywTFpaeVKng9C8NAbBZlB298rPnaM6rfh6MnFb2a4bTASZOWRvcOAjJlKmD+azDm
ywB5IvhwDFAihoeZTejMweKgBgY94Rptn7y+3o/7cKfl0jnD8ubli0Vz0fBJWtZFTLFJ4HCXcs2g
l0n9CrX/jFWU0c6cIGhA5Sb23IHT2yOGrYBJNsfqDpgyy/FRoIX8J9O5azrJGJ8+LLm+tI6M1V5n
rwVYycpx/jTquX76jR1OJTa0vK8lEY3Ax5Rm/0GLYHr7p0f7uSoHql979vJVT4Rny0ErQlh7PzdD
02E5HaVNVUb1x2BE4J7bX8BuzCAIlAkUeqVhhyVypghKZGR0HFWydrKp0iprq58ovk3vs2UfRMA/
Osq+o9EtMJsqucj1OJcOM+lgTBc6Wow8ndLdtfXiJUwWz+aIXsiHs2mG5bn6dQ7NrSHcCWd2+Uvw
NCSmd9zqsM4wpwKCioMVkeH5A194rqQkHoVAHnBFeuZsE0ugyBIWNU6jAxji7SnMYIXnV455Rdae
sfmFuF2pxqihemX2+98L+FGxLNKaIW40R8PiaRYe9mwBgpfEYwlmeyHfgP1sCb71OoiBKIkosAVN
uXy2FmzzkDhvMR1xthCUaLwZCsjU5FkiK+sVyRN75CKTsIflK5YoKquUAPaaA7puFro/ujYHSiw1
HKX3/dnp1RR6EQkJq3cm3iR/lE+I/iY1YFO6x0wTvaw9isBX60tsHn2LfoZDkdbcKVSunorbgu5S
lI6RTlmoJTPf3w4Nc3MEgLAQQ95hka78hiP4UUjr6DmNWyHhr77g0+gu2sqyZUsRnFe5qNfnRfSU
rpAL8kZwTRBhDnUwiHNPh0SSA6ltnqAX38xuknwXiBcNkqaPPqQEFRXhUTR1ymCS1lNpRJa4vVlG
pn9jPFlAAmwtkU9lM7BRVcQDfvSKSqSY5tlHLrV1E9j5N7BvNT7Mc8T0/kVWMfOCNPwQ9Ad289+9
nRl2TOg4/qG/jxkwwyIwjjiiz8ehfcJmRnjcukgb37jGq96lzgMBBKuopiW1LSWegflI1cbMId+A
eAp1SLqS7ylZAyei1XPjsC4Z6sN+FSW3Bsm+Vn8BWZ1iPIl2lIIunbtUxKmfn69uoLZFrLYu5tdq
0d/6hNlBpuKWgKrl/AiFKFD0lxPeOY5oF+r4q/lGwSw9mJpJXB+b1oo7NS2QFRqobYV1s/nR9Mnf
k14nNWFiepK71yH8uU3/I+O5+mn5t02sfc1MtLbFnIhfbRWj+hJ4moXp2paZh5hQWiLu5um71D1s
zn9q2tVr/H353MGYLVrddoPmMbDggXni08um39hoyZUvfm808IBnJzLhAKxk5Hi8JLU4sDFG3/4G
EWRgnos1Bg+zoWMPawuSzfn/YAu2S5bqZGoXkU5KOckPs0/Z0LWNPJofQ37D3Z7DecX1J2ZkxKLc
GsUfhPmqd2Mzwfb3QfgumIXAhFEyKJKTb4Zv6AxvRNUFU2YgcI/Qu+rH5qlQbYWF41WAm33MBcxT
taw1t8SBKC39HcDSn3TPMz7MBSVn6XRLiebqnc8tPEJjY2lZv9nFPv/2t4FEfCqwvZZHQnTHVU9+
t7Ekap0ZBqlaulM8MHzW7ZEeMJ1Dlgkhfz7gaBZ9Dgh3sdyTR82bushtetaBWSQmz6bpVfe6EQDP
VbjXZkhfWZK2leN0GT7Xg1jgjhJr4yrIkFWxcQ2Hbwn7/+qIMawFXtFxGapqElKAb8eyn/MheC5l
226WVTT09ttZZ4DhnhgGUTy9jVw5P865QHWxn/258RvLZr/B5KlchzAvEQccwj9MhI/XOzd8e4Ke
BoUCwtwZWFVxfMgLUteNKz07njXm1Zs7QHWFblXzTNz9GgACV+uJJLGIhmPD/OzRYJh6zqUmkOrl
Sb25xmMEDez8Z8T9A8/7aua01UPxCzKzT1IR7PDoHhnaZwry74EKiBZHq7MvUVbBCSGZjevWGuQU
xc81QvGaPAUvCZ30VoX7pvyS0G9tumgiNnAXzJE60up3qZybFe5E+W+8daXJ8lNF/1InaAvuUgGy
tY7wC2mHj6fr5vF9VD/bIK1wwNR3NEYfgDMQPGZ7o/Qaq19V8v1bGWv7hJqRs0tWqjj2TL7U2iXX
IkLS5fXgc2IRVwOFjp+KuHIwLp2LfZge3yYKQGO3ppFhiq9WdS7RxZMtl+Im7yRyywKktso0WJGa
u1/NauEkHeK2EJzrT0Fbd7mLpqOWsud92iaoIkQsxS1m8VdDZjzC2GtqaxBO0doKfYphZHOdOs7K
YfMtofuME4yZ8Xlh5qW37p12l4bDhk52cUQYMmr1sdMRkT+XzcyPIWqF6XVTjkJmGyFLGHoeXVlp
B+Kz+lol10pVOx/IxLlsrKLWcqmfJETADR8eTHnoM4ixKSGDSL2FLoxsD8Tpi7T4hZzfWTouk76X
f49iSzJa+3e9SOPI3cABKoF9glNQQOG/vuVfHKxYyv66i9z9bBvQx+pfZPE+OT0aLKC6lN0oEqtW
yVvzr0iGk6uU5g9R9p9ZOeVcKKybS7w6ARV3MvhWIthCXMwkGirFT9BItiXivIGuIm02IyXR3VHn
f1Lpd2Hx2ijN+Ur1lRp2Bk/WuCacVxPcI/IvOJl6Xr6X/gS0BCFguxnIJ6JGCG5Ttr7PNzQD0vKF
mKOh5pfX7BWGQyhMXbcEUgg8F7Jc6MoLQtgcDbOd9nv/Mm0xh7UvQVsQUWqu5p3vc1QZ5U4ucAlM
sIM9YIdhvCJLdxsr/dpssG2EMlbUfj2I+Lka9L7i53ILZ9SV8HJkNP469LIFgcich9m5Q4MmFVnx
zhS++lWcN8xKqQ6D63o5+YDJKvpuWIErAKy/o+LKKN/r3HubwGloTCHJzE2w744Kkw+rGLnqSHhe
W+NHEhRVBK1LAVHC3y+ZRFh+d62RcaIYGpwOffn0PXPLnxoXxWrcCD9Xjdjl9NgSdeIRKzzgVDOp
OIiWnsppjftPf0sS7fs6JLaeF9QF6LN9SZ3KHuiA3auSRunL/92zqMGv7Fzp2Tk9HIrF3dBOcJ/w
loZwMFL0lLuaaQWfPsWcc5sRpSlRgqiBLPRWaaR+mCIWBia6HsiI8roR+mIcKJyR3ZNVOiDqKHqW
Yj6eCwdyMQjxFrdKn5gIEQ64kn0lD6NzynIT0qdQl0/Zi/J8JHZrlR9CVnZ/FNQSSUocUyPeFazR
IywxoTJIfyI8/kKJgOyTA2RkGR6Q0izb5BjoZwGWA3IdZjYQBQa8Tt8vmwFayyzGNHtRCC71uB1b
tV7BZEcPZ4dKgJdvjjeq4dt9sTb2qyofxO6ZHm6tWGLgA59E/3U5D13kG2Wrdg6TSu/Rbq9M3uZ4
O333aNDlOuGIBBSwDyqtEGlcTeOfAbHF8yEM8/fX/pXrsEXXM/4RynXa0aaOzSANjbq75C7G+6n2
KzZW9qd2A5JMbz5YJgPpsnBFKvbvxsEzyxJQAsYs9zgxEQTX9StQQoIKtRHjKnwIQQRpk2v8Q6/C
2HMcaaSg12UmIvJr5N8E+RSEaVXMkh38Bjo7rL8E6D1F9ZMfa0B5ZvRKlCYgksRr33J1ZSN8cCsi
t9eSI/f0Iu5B2r1ZuXMQ7BKiNIsQ7pAH61T0EANtPbK1/FtXqiNAqbjZeGGzj2KCgtbqfUDqZfpM
YfveKYT5D0eKaFz+J6oIqaVmCrmiLs9TwxmSlZXkMtOqViPC1Xuy1xweh6DGQaF04FyuGbxsc9oA
gG3IdG6Da7tR7bEgGS3ovdatwtXVBolEyvoPQMFdJ+/9DgdsOdg+fEesfg33/5yz5DiGOYTRzdio
4M1C7GMb2k5OwQ6J6pW3p8+N+EPM8e26HieFxwALLANwKWdrWqdyIkjq3O2aZJd5Zfl6/zNkDqhP
CFRFImnITmTA2H2mBmpq68bUByDVfBQuWWOOftcRd3UBi1bxeyCJZFZSNYvDr766+cRbtduuO55u
5wfCzy6zNholCWPVmwEM3pDI+9IjnYi8Lhqw6Ne3CMfQ63T8N1WEgJnzaQel53IswJSzdPvyzWgY
dnMBkvrS+wPUwom+Xi6hCFt4BUjB8FXyv1/DOvE0if8/wGEHRzSpgY4sHVmJ9QxobB+GeBa36P+z
VdxzAM6ltO0uHpDMTF6lKMBzngp1yqJVERsd3mOZudXZSRiqN50/9Ty5BJLh1uD35oPf/pIP862Z
WKdDAfKDXtMxeTwz0RyF6OmubOs6OPbOQVpxJGvysotis5nt2cgSRxEWYbi1OECrC8KR10aGkXwl
sdmfKyYmbnpCg62bSEoSs9+cl4s6pKDYD9a6ygtuCCbS03JKgRpwk6DkRex3w5ipFms3m9F3zBAz
kEtPWi/tbS6HQKgPGx0OTwn7UBgfHgakFtIlozzzyUA0LD8bRBXaEPOAiG0rur6s4SB3BWgeysRZ
XsB0xGpvI4v4h2iLZAaisD9NVU1VVmQvdgJqaRiVmmwLPL5UP4AtCjqPXJakQUb6Pkoqka4uW89X
Ab7Y46t50RNa+4rCGhX27HWCLu49ewoV/VYY5CkEknkQGJCXTCV6lYGTdvq5MV6lV9gdcnn1VCXo
8L9Vfw1S+BQPip0jl+15YDF3uM/mFzDaFzoaATDiTB4WjIqvXoAvcjOAyhB/wioveUKFXWqMlX5E
NP2SsTYLvdW/PwT6WPIRM7tII+IovUsZZ69iuKoNfWPFj0SrsSpQVNvcl9sSVcGHKMZT9xyjBVNT
G0undSz+XEuKljHE0IlxrHWgb4MxtHOcR+t75c331kBgsJW3Nssuvik9KdOPiVUIUaTOfdj33HSC
TGaPlC+Kvjlcufi4NYS0FZOQZhnRAsV+9fnyzi5uQs+yPsERf3kWt77d3NaxK5gHGbGtHHmKVZRj
IZeJHPJsXbpZuzxGETrgvSO+OkzvDs0ItE366PHGlNHsxvQVQjWuRZgMEyb7pFg9R94e2eeBO97W
fKgkffThoyGT+gCxSHt2JbUBexydx6Rnn3M/2WmAZluSJEkqC1gh2EX4pkxGGj0DOaz5hhhIajrM
2rJecYBCqk6B3UHMRLzgqTeq+drdeG0G1XKj36NQEdL4DMg4KhBzNiup+wSB19FU71yJJEaR7Iun
sCHpcQFYUIpUxjGYUCC31kkw58r/tqDrthg7wgU/He8Ozvw9MZjnBxl5xLlWxHZjsiuJG2jVTj/T
BWo1T4uLOhYxBntDxC5yHKGK/OJuBF8FigmxzMrGDDBQ5Ai+A766K7BMEmzewrbARnSqB+vdiNmY
+4qsJFKzL4N0jpCXiy5JlKO5nU1V8INXCwGGT109K7ZoZjNp5zlpCOKJNcbVJKsk/NA7o1Fnc1IA
gurKQx1oQVQzcsohO4YKJhNKhRut5YVhTmKMnLz26RXoEaCW5ultYdsJWxt+92JG7hcf2wPhZ3MM
0RHvgvyZ5QauqTUKgXhbXraZse2fdKmxvbnZV99TSw+1bU8o1qsI6yalGlpMS0OXqTUufdWRFue1
dgqRICpIk+Ht8IcfqFanE0Cmn7rnIpOftt2Etv8gm55s+lhPMrzpIQcsgRdR6B8S7DFE3/7SwgKK
AR8cfro2zZZbgK9fbzrys/Vvp6AkEYioXPdiWNklr1VZILJzaHrTHygRSexFlal1Xx6UeLmtlI23
UujxMnS5SOw8b5uC2Eb1UPuTEaWV2nLOWJbnz7CeIYbrG+9ZFWaH+BcPAl8r7mZn5PNa7EIYk7nd
lpg6JdLB8WfL1fJk1amx8Zh7kym+S9J3Tsk5j1vAtpCYFFNLmRE9RgBOAiGzrD5iJ95Vj4Ffqx9U
MLZj4WhWLQ6hi4oNNpJ0wAoUKtyqtwha7nlTKRBs4nczSQFbkYtALxtTvKv5NXi3v1lYiJoEeHsm
7syP73dQqtnB7uIh1/AiIRwzuyxXRW/pzrrSfa4Amfb1U24PjpGKt4GOgLQPDCB92DVFmv5v6B0f
fVJ9IMz2IF/4AwmMpmy8ClpGS+tLXSbgQe93YTZbaXglqH7NKXQw12T22qKqmWiX19a11EeH1BVK
0YqN8y1tjxx5bb2XcaFhE+zj/DjT1vbttrJeOXck/JVDKoj0Lz9Xo/bXp/DDswuupjm4a7ZtzvkV
owHewkLxkAYQk/hO2JJEzEPerb7kD7fne6uAJc1pTjKAJpWpyF/IuqbQOc/aSGB2qfS9tdqZ4hhH
kuVs/qzXelIcauJhlX4+0BTWZAlc9nFsALKoqvH3j9xIMylnA2CB2+d3APCWv4320oTUlyiW4b59
86HlXT1hD9BVRt9/C7Tbq94LM+83IkphAUS1755DDERV4Da9o+I5YNI66ERyDOSuK6obl9H97Jvt
isRxVQ6WrxsYQXd9nReBpRxPvWfSBzEsC8cH3AfzVIRMcK26qY8i6IqVZQHsIf6M8YrsuRvOJck5
61EDiQSWg5PAKATfYiEFQFA0zLrygqysPCsP9WXd+jqm0V6IKcLiD5OqZVD91Mtj0NXL/8/UFE+q
NOkQBiZe5NdgFyxL4oxsCmBG8c8qBf2nXNY+4GBkmbl0KFRQ1NPq04gglUXWfg8nOGt+Ptz/Hacl
Hf2q5+n4w1gATqJRAmDhmeHzYI5hi6n3E45TNLFPg4/tv+CD/N51m/bgvY/IsgPql6Kqc9ye4kQc
IHECFynly5n+oUlmaeCBdTo+EqH724QUmv32L5JsKBadexHrvaZBui8XJ4TOdEpddyoCDhXpwFqL
SvEmX7Ii6sRect6fffKrLsUAxba5SQxEIN5l97QzRTvxHDrMvNaBucsX+J3FXPODqk6ewprGJsDy
r+HaF1p0cdJ0y+7tH+sg0zHGHIuwnaPRFpolKXca0t0As8h/LIzuN2DTd0EcVzkMHG4TtFaTbKtu
YIU89oTt5VMLbg1GpQfcyXRPSfSvLZ6Wp7gdXkV3lYhmmew5V1jmB1czTcprdqhJ/klLDii/fCT+
lu4hEDF43dStkgVGYxhxeMVF4PolLt1UMWhjw4s8fwR7ughK6R6gETar6xmJpcHyltuMdahqqWja
EldtDSFJrYQwNYF6+hUBhgMEXm8Hh1RBRZqrFViO5IXFlBq95B8qJiGZO5TxzjKmR8NPuVYFme/s
CynYqzTqJEYetD0AqzrT+OM5ilnq2Qi+6//hWlYYhDGZLvpvJkcEzbV8j0Uc5YAvQpP4DNIuzdZy
+HML+WGTOH/Tq16ax56NBG6bJ4QFuwUtVqzs/2sQUoxQtzJIbZYlACOf2QfYkAQHFipFkrzDaT+Z
a84oKyCJr8nzeOU6aAuFyDaGSF6yJ5x0P37FMeNYmnFMJL4z828wAstZP/3wy8h2VMiEVrUs3dBg
5moN26T10RqcYNsYRZTN32taNvwz0r5PEjJk6VLPyPL17hMB2MDgCYqhL4bx5IZeTVp6C0RWb+zy
EI5f69yRLPBQtJZXhfJFSM7vKDhBzIxSIuCia92sMqes+lN4SGs+cBhCiwoW1rbHghpfh4KbqC2E
6LdTCiO97y8YXkO1tp7YGyw8FRZIMu7GYeKIFn0wFVnJXDNVbxBkz1SDc5MNWWukz7zBgZFU4bBa
V5mlyaBWybd1jnieOdpQXHEOIKsAbzOS335wJZLFwiCioHoFO0NHoXRtl4p09GQuOOM7buMD7qFl
iX3Fp9GbvCF2n2fXQWaMpa/Uzyf7JNDTfFiiY5l9hD50/kCOI5iJpI2xhos47Seixw/LynLkB+PD
hFKKj21v4ihk32uEt8jMXS4/N6M2gUoOh+FlZA3Vx8SUfR/5coOGzrog9nfv+sxgZ1TkPzqG2SPo
/jqHfBEFmH1oQnVCT6fcV9xPcr2rtoKEqwJGc5ZMUi4X2uOmr0VibtetQPwtUW9Q/UfhXSRWiWJB
O7Opc+PFhXbY1yBEuJdw8u7f/Dk7M/RA5hX7sISBHtPOj3NkXImLKGuT0d4d01KKLIgae/qZUcRu
Rz5hfnHI4unYZcTDSD+2bL/yPDyZQ5q9jF4tmCivKx4+twMgBzkQcPOwtkeAEfp8TQjCIKF/CwOn
CuYigqestWskhRy6P3WxafeEZE6vFwN1Pu/ytpvFVG84Me11TSn1XD9qfS0pz2PU9NhaCSyDq4yf
Pra/cSqSrYnrZnhLlfUO9drsv8o7Tlo46eCRx8M93Digjs5+kbS9mWQTjNKh39++mwYwZqxsmtYq
nibQ9Kc4hj4mdu9zt161RQjTCAXnWYM8UiFaFZH3RXSfrH4168nbrG5PVl57dIhPO8jJnHJxcCfu
4JASObcjzP/sd1tjJEUPgWeCqPeLHzZNsyN+VHRdQuuunwsHRe2vmGG3mlm7724nFrcrhEk/PhJr
j7W+Qst8j9W4TAuuSlRB9wjwkHfAqTvo42eeUBzNFxywzHHLVurvsuIWaKN4q7648fJ6eJPRN4jd
JO2CK3LjKDx7f2DC0llzhu6l43in+oqv1OwEc9JMqt1cYkZGEi4frVqsl+kKdYKv8MJA6tN+IedF
LiqOatJohifoWQ3+xpKyoiojUVcZxE682cdZ77nT/RWBgq+i2STTNGqWkV2pcaraeakgWlq2Ry2L
zu2hEiNojRyrF51CJbLn5oS1dogIzv+yGyOMsSc3m7HWLJmQc/mHi114gh5rZv4bOIvH7v+SvTMb
xdm01onL6yrkNnSFyH6PtZVkHUYHj7y0UC67DooaZCZZkCAWj69StU/xBct9ey1RculJx6GvrJXy
fTWaKHiOW2JXUBPH5BIjUxaNOuZz9eP7S19tkVp/Y9DsgNiJ11mg+CCFGxskfBrhrv1JbKOweCzI
yOg+4bFWmSjlJMGx/gQhLuHXxNaC8BrMSJdDDBxtinQIE/RKOAWuLj+z5Xi8HVBC6WumOJSgYmIf
h3Xgli/HzblfW6P61KCQv4dh+VQ9hJYp+RiZ+uGAyRt/5qmxonLHUqgRn0fjv8VUYi2wExIHXei3
/kcgPOsCS+LiFxkyDFeHRTA0Vtb+6seTb/ZZXDca5mn6nDP7CR+R/Q4Li8/zYxUJG0Wj51ArH4hv
tdanByWpsRejsznGCJIxZH9Ipjj/ZGNS0GRm88wriDdXbmr3y2//2+k4M9JtWQs7Tjy+jzA3v/oh
WgoXxrw1ZfjZlQmobkE3GtHY49aPH4O/nxjcdjnS72e7g0G9P2affHBHXzdJEkuF2JDcetRrix4i
5T4EJ+Pd4PyAuTpys3mO/h7QhYf9xm6uVCOLwFcd6vTeB+WM+2h0QWMU7k+MiiFUhT5wJ+f0ozdz
F//lLrxOyHCesFw6er/9dTSVsQq7dfOYCEPPcn7jWKxu44plKeu54vBSeX+9k9hjZRJA7b13FP5a
OwTvEk4mnh3+9ex/tn1+CtnijSWHs1SfDu6B4Dusw2ml8sWhRm0NtY5zNDZE2r3MvQRdvhS4CaoL
m/K+Cg98KTs6OwZZpetDMPW9/pfzHA6SGvg53e31vMbFfz+13Gfsepwel77ORXae3lCbCITpj0cs
gL3rivb1WwpzFzHqlj6KuJqUIpteiU21kxPjrelJh0aTizI+5Q/CRjmJt5UMNtwUoETXvhzNARYB
Lt9F/xLfg98wnzjRlL4jzMTzehQatGYwSFOaBkkAR3Hos5eYCBffBQG642xRykOqs9o4JdIxVwX4
8lkSJDYB7TNLd6Oz7cZdxQVgyCsKE/jQXRQZlYfFCAjBnZoWMLpRRZ0ty1Zt5fbNZfBPnc4ZRRmw
/thmDFX10IE+ZeI30xM+GZ7nLjou8jToSmNQ5p/uIoQDAAyS3SmUCQ25iYDW5e2wLT1GRlPVVyUC
T0kbDnbAd8vg9Y5nXGSwh6wh8zhO2VEK7bEI/5aWWW/2JfjA+Fr75ctpVhH8Vz5IDXO7HMRKuQEW
Llz03p+gox9YTFQXVDR4lb9KAbp5kmzsKPdDDe3xIK8/RBu1ncWLP4stfqwDQ49ZV9NZ+N6kiSm6
JMNNcQ3hDu8n+JCKURCxbRRKQaMmHOBMi//ozlSdzOzqb3qfWxk3LC5mKCwtAMHxLlJQDcz4V86/
HgMKqUrlsiqm7gy3bTfADWLOSZxHIcB1Xg4ZT1dyI4P+YUUyDVOVrKFcvqk5DV+O5ohP+/3/ZATj
0wOYHZs1En6//ANg/1kYFwamAB9Vqw81BU2J9AMGyYOmbI3mgI67zLKRIuXD6ruYjq102Za9jsQs
IU7Iw8u9W97pX59wYNf5f50S6ztyO6NV1/WiupbdBFhVISXLh/Qtt9G1oPUC/JW4HYH6zalyArMC
5wSPZj45IpL4BaVmMwhEkk95BTFH4Q1+fG4wQpBakCfAIzrVsXqyQ4g6vJC/LBPQMP1NL2bL+kBQ
HGKsszNs8EewZ+k9x4VZhFXD/w0fEQvb77eQ4EcCdeEni5V0Jhq1LCc7kVlvfOGWYxdaQETliF+8
AohMzZ+GDFa7XwTT4/ztXqY78+CsAkRoIiS0W5aViML7iYo8NYRSsFu2NJTt1zltFggSju3f768L
YFqPpiFtz3E3C0G2B0VgYuQZaPnNFXq6DTDKzT+QFXwy/RThpwbm4A0cCtDqJO0y4Gp/k2iP9eoN
zDe2zC8VawV4axAwmmnMV4rldgrqbU/mKbisyQfVY+nCMW+dEEOhWtE4TUlyYmznQFtpETELgqjE
Dhe7rmQmVXse7Uzb8VcX7poi8mOg09zooGEpMWrKz1W0ZUAsvtyiD/1kjWuawuZXFV6zWJdAPYsY
fDXYCYGx7vWk7VJEkzUhY+z8MjB0wKQDPjTuwn4/16FZIkU1QosmY4xqxsCt30Z8GJP6WTqMNa99
gtyoc9w2/kHs/QhbLaDFeyXTTvabTIRtShX4j23pqYKaXBfEDR/YpTJhwC+U57rJ3Lr5wenGQjdN
c9M1S+56JP8JeD20NraeFYJiGqVzeWhUKJXygvaEgbEychy1xkewzQerzLav4+YS4BjnMP/uGVMj
O5jn9ZOvWkgflRvWZVByKem9p8KRLnDws0ucXpSfyw7pq8RTUIhXIoBwGAOoeZXHpWHe53+QaYU9
Ui+15ZDQkD5l855AZRzO/G9PByQ4Xyddd0xZDFfE0c4CScceeI+nXdZaEz2tY4fXBbbS7vG/13Gn
0wqlv/f0hktL4yYRPBbKlWii/2xOczqfMn7Clf93R+mjWwVgHcEjlN9+/JuiinaiU1HZjxWs2Cyv
7gVMPHQId0eoGsShe7xAmruwBUoUgvQw362UAWPY5XlslK+ZeUYqocw1mwq8pmXpPQp7tNHvD5tt
1upzPpaCKvYqoGHPnlMKIeIymgeNOkkMkUZMo0prKdDVo6NynN3T8cvIfaNeDElk68fLqQ6gT5ZC
HUMJx9pLf56MA/4p9mfGEGPXoOt9PdphdjuJbcr/B6kWm5UxErVWj50jfSn/f+AXYrn3ji74BlmK
A4xrQcy3MJeBC4qbQWaQbHiUY0s+JS6/YFRc+/2bNEdGTZWlIpgmRHkDywVvzSU+Z/fII2xezGg/
x+JyDxS4ePKT26zJu64Xy17IB5jNXsqy18EPGg0CbTd2IEjHxL9foTFU8/LPOxUap2HJq11Z+POb
BlWWz5ljZv6uMR4mblAjysMBTRFMr75qlTcFiqWRdPUkUNBlrvmSbGne2nT/S7fSiH9vyZqCnxFJ
HX38qgQyrFEfNt/Qd+Pm66XWXXPj7owBLMQLUUJMGuP5UYH5/ejN8x1aQgV6BvQUIZ4epZTC/u1V
j6G7XTO07YEyIS1I5qFj9U6MwAWNhwHwCIqtHwvtgP8qUa7eRN/I0qMl3nY1prMV8UVnOU5ZIe2h
7zB3yTMDKXvqpnuzOy4tcd+ychvMtJl0JBFYhxO3VYjVF135Tu82BLo6fKBZndYtYtoiFrNHqSk6
Vv937OMCVUY5VwfNKV8xqGicStsl7TJdynCQSLub/MT8NqMKkjcULDuFPb+VPekFZMb/WDIhxWpm
Gr1ymgitwvoAyuJoWxo0R9i0MQh79TOu8jcHYonhRABjCydnUQhFpdG51BeKA69PuuScZia46XN5
RJ/Ulg2nfeavVO9Fv7lNw7v23vhyoNa8CdXDPRjLKEi0SLnP6puPpiNZX+g3e77KYkaqGOeDR0Xa
cu9jJX+ZcQkSfEVvpP2GtdOczooVVMmI0+rwGtrnURXyvuHmK/S0GAYi3usY5lve021Wbmhi6pGd
EBrInvRZkwNjS000SPFtxYk6ZOZVjgdaq8YY96opWpP3NrjlyUG7f0OHB7TIyvnI7Zea+zxNLODL
eFIuMe/wlwoCNl7A9GX4wRVxWmTJX219HYZg0+x/kkJwnuJ4B9NjxGGKglSLtcjJr/c1CAFvqUpR
U7p9i3X//eV8KCY7Sk9JGNOim9J4V5HnLV9kqKahQ+W4z09tYMA3aAO9oj7bs/QreQei4JlRsoHj
TKrJRhONWN/TJD9w/jaLLBZ3rSC0GwK8YYELk3tMjLetPUq9VquMxIRYXLxAKnWMZFJZOXpgNZGr
HDCueo+UE6zFZqmALc6M+kPw870krXYZ58sfDHhgEiFTXTFTWFcD6BznuS2sRpLxIgmA81XCz2Um
y9lwWe/l+bthd88eMniEuAgrYaBkf1p/L2Aagnf2+tB4UX+BxrR1R9VgmwdRDAymC3NiKNE73tPM
e3vJb6JXbw1DWZM8hE60kebiAlvditIuXpaefY7fCPuBEhalxBqDyTUhRoROL84Wnxr8HbychA1x
B/QXW30KdmRkYscySBcb33TFxS7s0Rd42Qde9AZWYXEoMSO7spMuadRglVIw8UUJL5Dd7Nws/xs9
AUry1+Pp7tm8MFkVfxIeNwMEMgfOSVgujZ+Tofjq1f+EMfV35nY5dI7P5ZC31jK2dACtFmUV0xJ2
uLWIgyx5CAz5qWbNAnq9AMFH43E4hwcKIthUkii7y1cbvidVTVVQ78kMXc2+klrZYyblJFh/l9Ky
4T+OHkuTs1QKKR7UfKlqqpSA5MEHWp0MJgY2TOnclfRh1cxEsg1On7hdk2JqG7zudk7MBZSzlRov
4/408Fa4d3lyrblAcyD+ruc2pf4VKkPnuxiqseLbFxqbB0B80WCt9pcv505wyTcH9Nz/XBaEW0dK
2TDsqnlEj/22z7PxXbpz1EHxYTaAY8CkZDsOelXueU+Lre/ji3diey7Fz23bIBp3Ib0p0EG9Da99
dWi4avJkEV1cBv8fQW4+orli+mnsIc0GnNfcko3wx839PdTh4Hi/iUnFZr3fA5mGhltwoWvE19nv
4PJDRRbh5TnEoXi3OIJjjO939EEoM36UDt65TVTkTdHn1As7YNd5iSIoohG1Akvd7YvuEpvWJIxk
i/TZvy2EtpCpBC8XqtDFdPo1391NQuR2HKlwC/uUjzKXm5VxfEJqJic2DalWgUVf7k0Rd/AV4NTT
IKGQT2rb9gjTXATlMb3DI6DOD2jDQtqWPp6E6XuYnsogu1gFugROiEDRZpcls0t0oZpatNi0+IWp
D0Nr7H0ry4M35nqjvEiXnkUgZsQOQe9Yw2qTfHplj3I9QtH1HFMyv4HnY3QbbzcN62bj72tvacPq
3ZHy61l00/G4VwKINqHCexNrVDSyrD23tYO2Qt2GN9R8EG/CCRzA4Amyyj36m1g146o//V8neLmM
QT28P36sC38juf9Kyd557sl7pTtEKM4FW3fu7tc2Te6cpO256ur1opvb7JfYcQy3hCTIOazDhIM+
9OZQta2UwaWp+6ipIoi/f76Y6AJsIkND0uApsmzWTotpdakDIYnQduwq0ymcZjkBso5zBBBUcylg
FqnThyym8VMGv1BdjNsFusV5fSrgHHP4M9XI30NggdfzV9zDaMPUXSyXbkiQkIwsshEhMC5rdR4h
Bd9JwWlNhieV7TyXLf9F9cVikUsHTZIckUBZdWXH1MT55C5GBvSXXizmAQe2dQNXvl62PzQRjZ94
OcGM25a+sAJqJ7PxpTuviqRZ48RqN7c5yWcmvZvHDffYTrJTVAq/LV5zz0waehtRcwH9rza1rYNq
CR9RwNHRbzZNdg52ZLuZqvfdLeZ5oYB8dCe4FmRMCBOc+F0XPAOxo1YrPawPdq14BaDfridol7sh
7+8scJFZh0nyUI6k9lgBmJLlrGrnDGBqfPaInbxrC+IAlprL1PGKvr+KcRLKoBC8fgTLyfRI/COb
X9+JcGV6CIIzpcZ1CeFe1eVrjMBu6YBUfHhHkxzoXhIAIWg46tI0O7w7HV2TlWMkR/JHXzJZPT6A
f8HAYOELOcs8UztnKYd9NC+8TtVkVjoLlZUoej9r+9i7FwlpxmPGee7Vm9Az9C5kqlAGYc6+PKWU
bTjrpuNFUFapXTY1WOws6HpsvvTx8mKBgOM+78/VhMNRfMEbzZLcRdGu0bqrjfkHZ/dWfP5/viMg
9xjUeT2uJ2NvBoN8+g6rTi240iEAEIzcmy4bUNi4aVky0/CcZIC/xpv33NhzS2QEFXJKRRblalAi
+o1Dh1ygl91c0ZDYjjG1XfG5dXBF5oodU0x5YUzd3J3MCF8qImPiO4CLElN/FcCRYoPYX6DZPyrS
Wbw+0ZpAgbPKUcaHO/7DSqkHPyUVSE8raK/gPaiw1eKiR7tQKI0yLUf/Q+LapFh3pDdtpdSKrc7G
DIciiVpHDfhZX/7caL7BdW+1gHT8XVApiN2FhEUtf7dDc2FrjhqvQNejDvMsM4MWprNxjzEdzrdn
i5Lc54SgHTv82Bg69ryNJKTD8FJRoYPyawwEP1V8M6NVwQTjv/rQcIKvZCZRRkADqXHnDXPjWS2x
z48/MOKiQyF6otJScX9p9Osc1IxfleL6FDbltmjQdoexRojhR3zGQXQ4Q0uXrbPbK0aO/A5bHhes
rxIvGBRnQR1pwHwU29M2KfYqjhjdNwGkUgT5XC/GxvkREmMla76ly/FthaG/rZdBaTD2vvL+irVN
Ue9SHajw6TrHGyGxGtlc4tcJCn+2MD3mfhM97T5CVxoiCmZD/Rn2KQicISmAw3YqdaZOlT18xkzy
gJmRTj5CeZVLsZrPsj5BbIU5cxize3ZR1ToHstyaL6ShSd4M5Kg9VKmwSjFaafZZSGLw5nPJFCqP
kK38dTcRKCPYIZV9n7rw3wMhSd5u/OAPPtHTPPRx+jQYg7/fPeLyvnUenEsuBcBty9u57UeituyU
9eTAY9FMtAw5AXBNwvbXtmw2wjCPYvRVeVgCpqL1ogdYNXVJWCKAF3v17PNZMFA7LAH0POLUWPCi
t9/sfCAg/f3GfOtykKUsZFq4ysUf3fcbZPTuNgtq1Z++MrqX7fCNKvBF2aD7NsBUVK7anR0sCp6d
m4YfqyNgVC+0dE/puap30loRBx0NadHwt4nEAd7Yi/DcnVUfrGBE6OgLiv+e9DloG9jiyx2ongIQ
27XVceVzOaSXtULCinqlMZGCP48/BvtCyRyvDkqFHIAWN92nIzJitpx+hnWFdrNcKEfAWYIWZAq6
NqcxUliV3Dn/H5NDUJLSGWy/Oz5gBxOy8nw6vuFzhum5SV4eTzCHrZxWlfH/5yHPvyzaobs9PTkl
fmGJBZv/NV0Y87HnBsdAgWC10g45+dHNN0iegrA1blV/7YT/wQOaIc+vfDeI89/SjJBgFnC124rb
4R3kpeY4Kz0UIx2lUJSK3XYMAre6Cn/HTm9mcqCsHpASVG9fsQ/I/bR6OZ6ZFZsC99G34BFrHGFX
kg6dDWUDiTn/mFtsSdxCcl9iqs7LbCNLF1TqISFqvVDXv3/BfMTDaLbo0NuaR3BnWexb5qFW9IRf
ErNoQp997wI3oKtwa+5S/u8i/ydlfIEltsT5t1lZwwmZHIXMpYe84+IsxhZzfDLQ2zsrBoi2/VpQ
c9JFhMe8zkBn9YTRbN3nmHJLKHz6is34NaFbnWQ9JD/ywHKHRsboIQt1ErKsgUYAPMxpCNYiavKw
3HRvy1+z8kNgpmfO5n8eDEODzH4I9320Hgugij6bFxSAJJS6XNLTtbbDvuG6F3fgBkxd7nKLWMS9
MTqIpg9/gM3jViyg9zWTZdmAWw9lKoiNXA65+VF0DfQCl1fMuOkdHFPd6iXZZmbtZOtWsySWPzO9
3VDjcYGMDm6GlYhG/fKXKmwUYFGIcw+qwAOTBpP/O5ezZ5hkYfJ0m6G52nLsNNYVgNVQfSG0qHNd
NBfaJJMDRS1OM7sNBF6hYIWuKmyAy4PLLffC3a96bmBI35S6J9PJKjkpUC3K1fVn//aAeochtj3v
JkTTXDWNBpT7pzAtdsca6iDo6iaM9jUwDfGciBPGTewqxOevnTZpQ22FNfLKoJyefznK9Sb3tRJ0
TuE4oir83dKo0QaXRrxb/3JUlezTjBDbImxNGOhoKL1DN54bWr91/8/5xvNz9zWWqMme2uoZewEn
kea2B8ZYwAP6Ra4YJLnfZ5V7UrDuCmFYmXjpbNRltD2t7jbFLg6HeteG2804OpRqruCKy1hH65Y+
VesOQcxTthgoOp+uN+wizlR+AYE9U2MToOU3M5dSKiX20RSoMqCWrXnJ8oTGMtFyiaMoy2wNaN4e
3CEyURbkFANZ2ZOfZcIJHl2tGwNYtMRXLH2oMxr4f4EICbigH311YJS3FrqNqu5nvt1PNFN5ahf+
uktYDlIzJvDR8OVmABctYCnL1ajeEKFHz7WiO5lf80duqtcOcgF/h5ozZeWrwo2tXms5Kk1ANLYj
MGaLi6SLP+WMXdNw+oXL6UNmAkAUNTgn8Bi+Q9rci7MoxjhDxzaIPbLjCTR29OmI78P+SuFg2fZ8
DSl6NbiPzOU/sm59ulqbVXQ+b8hUsRw1DKvl5g9aU03+VSSncT8RTFRfdjwl644TsbdWosq3mUVu
1euNg3+82z4n5DIJTVrNkoWkasTj61g0zO3Owa83VuIQ9GiWH9SSB377ZGhufj795pYp6iKHHmNf
Xg35x390df7U6VXco3+iEfZ4qFYzWs9HagQAiuStX8EyOx6qr7OJ6P0RX6TenTcSnSzLn6pkLAfi
tjdg1uAqLPCvmhcIM9wOeCAuVJCYGnC7xHpFueUXPrn0a3aUx27cHeNPxo4MDeUT9FpAZn6Jvk9F
v0Cc0gVwCe0+nn9LkdkqiBoVnLkU13PxbA/8ZK7LI2brFbEI8I9rw536WmumKqywD/6+4rOSy5p6
TanEqE4RM8aMUptaai4lRBzNXLAk7JirQNfJHt/kzOpip7xudEqp/IOmvUjsyELlC1CGsJb88jrN
AO8vixP4FN2kdiQMD41r1HSi5QKPFWvnCsYkmI5JBAG8nFep+ktDDeNR+zhIBGGtclAcPP1Bnky9
3Vdci4Tgfd4GE2rxCmTPC6vhbM9efBaVsvxPepnwyoufQezRGqcXbYsjAJ6vENWDWXuuHY+G1xBJ
/8ydY3NHnRC/RIKDcPUnb2TTutSKY3J+BuijX2gTKwZLXZryXXWxrwkgnpo9JizpcYAmjvd4OVzV
W1yh1BpczBeTGXRN6HR5FxyxrYAyVaqoM4302MTH+CGNHaZ078N/sY20ueRNe7KQMeKdKt/lZhXQ
ssTJcHK/YhRSHnsoCHety/nNvjKQJVYLNCn5nVBB9Xucs2u2d9wuOTb1IqS01CmdvxfwA6joQxvI
SfcO1RzkoSHv7qI5B6OJgdPf/iJgDGbNvLECKGrUsLWfmDGv8mR1YJ9L42fg1rh46Ny3nnbBvn/I
r0bfDxQVJUUyC1pIu5+iUwpqubeupTfaS+OSatAJTw2Ut2tMAiaUqN1zHtYn/55LglOBwIJk8Yuv
XvZpwT8IL+wynL8vLRCh5OvU2JsM2OgeYf7PFUDfZo0ehDwSibG3ZyEjTvhhQ0zlc/qY8Nc0xz9u
/rfV/xKOjvy3LIklPiINhBNOF8LpWE1DpjT43SFz4AHQ47Rgp5RududxX3fZaYH8pohbq2kL5YR0
YBbD7voAFiO4OphXDK/Vmng6G/ucijXxEMFoUZ7o44K1UDDmWPdrHF/RYKX9bZgphn4d+IOHwDxk
vk9zP5EHp8lfCpd6r/kJqFR1pU/3/O1Yk42eXvGx5VOmKUGbVI8r+2cLZvbEAA5IWcAABNFZ9nYU
tA5/kZts+CO0P7rL89VHJ5nrVKZ4oF1RZxmH/moyM87NGkPLn0gyqWco2U5xpIxoCypPjR/4+oaD
awOZoINfokqMuWHStBcxsAsYuHPpYG9ngc/cBSBI3Wxq8H08+zBbw6pWRDUNJtGzKUr4NDjc06Rn
Th5HSvhpt/KyfeLsjVAmFanlha+/hf58tI1sLeVULaBdaA/VvOF+8gX+WGd2cUM23rdx9ktFqgnv
H/HjMg49DKHiQ6PAIDUIZy+ldkNjO3TQUyPqsAQ/upt0PACavsae1Gy1Dq6lpsmh+dNvlsDF2SZ5
+bA5XiriAKrpf4LR4VmAiA0lR7arpCcnNTHTjYvyYJQypLoAZWBJKkRLEAo8Ibh1Oai58Zg2VMHi
DS4uDwYo0jDtZvdw7EZUYPr//u3ZF1tGdO2cCFbTdsmOI5WznXe49qvTc15haWTxunmK5+qJWpTO
Mjzq0dqh+WcrpjnKCuRXtjKY1/pqvPFYQxBWBpVRpp6dnXsqnqJ5spKlcQgt+BJxNrboIgFgDQIL
R36bEDqpJRbO4gSuuLVunaRx242CnAQek3JhGKacFNQ4kC1aQyH0t6WRMbj2gSnHZYhLP42LCERz
8iYydPiyf96EHMm0a2MKDBsGNF3l6wEUrto4ZmIEAqU1NwEsPMjTKP/Nr0RBmQ851YbFDIZNLcDi
sCw/JU8BYcbeECwCYnpAYedVjEQ8HrHqhRwhBc0Aa4dLWqBfcBOXVP5bRkHrdG0n+H5jXIXtRnlK
qL5E6uyf/FZBwVvEc32+vFxbmBCKP7AlHomN/hO3YsenySjNiEuNwAg57WtR5PfcBuKNhLYrXiHA
FBlO89c6QUjeiQhh0XbvHk4BrwEs64GvMjIO7aGtdriLVH/qVNeQU73A+RJgUPgzkC50WBHM2+qB
yiV0KfAGtPHs8UTTFNqevozWgxT1izcwqlrA22q3I9FWlCWjipuv44NpUlOtgEHAEJI6oSdw6tl+
6+zkPx660P22j7Zc2Nd2uCO0xT6Vr7Hs6NCCl7Nsnui2SoqCpIS2IgRrWYG/LzrX0tEBIV0lxs0r
ht0S34o2AUUwCSSnYYVsvKsOlIL86k6vnnZ5pEchV9YrNr8Pl/NKxv2e2n2tJSG3jhbLSuf7uFi7
tAUEHijeDtytfm/O2/ZcNZrwWYGCLF8uwRsaHekW1s7fOKi9+7Yo3XVhldCDDr1nlqWt0+vv4+dP
TF+mweJauLFkB5YjANgytFH/mkfR4eI2Ep6PmigodRoSBsRGvcJXhWckt906fBHpMOEsh2q5mB/y
4sUbZ4z+rxKbc2SfuXqIfEG+OQ5oFvzUhBSHI9qLIJUWi9a2shT2tzo59r5IRwGMSNgQPH5rhfuv
UVNg2TT+XbiRx8SzHJjpZoMf8i56vsPbU/d62r0z33hV2NCa/UDVitqpZx3jlc/t5Yv2dR4yxaHG
m1qNKVlvIyx5DFmgpXAqJfuV0nlfFRY7ZfZHJmnxUO8VSjtVkZLZBJ6NnUINn4gawznH1zQ9ruiD
7jKijSOcRwyLtitAgxGtjtWeP0lKeWw3Xs8mPshtoKeiItt1zl0JHf1OUq4KSerVQ+Gy4RHbwzbr
sDwf2qv0QB+tUb5l8+ix3mUDzj4vvknHpJVhJxN0DvLUvrQhx8mRswafC5QN8VuNg0wK7EQpzTBG
r+kSJ5IxS+dOe/Ye+pf7kjv49oNH6hNjHGMKWNf+GJ9Mbg1N2bDCePG3KXvIKtP0AtJ4wPlxGOvb
rRG2WiYljJujifkCcZ8/7VElF8KxSD3A3l5Hoqk0Bcjr/76qL2WKneV1GLCGW20gM2/5HRtIAfYZ
hBLpGmUjJd3ps6xPLLsKg1Nj08Rqp8BXdZIIdwjUT9j0PJbktQFd1vkJWA3d3nzBXjzXw/A5DKiR
JQps+B+G55EKzuKSdtJMtn2XDQireanyzvfegSNUr2UAjSokie4jVtQNSVs4/mxT6Wz3bpOIhpgk
uNplE9GiYqNMaHzsv0OVznR/UsuyZzgMIFjFnn2KpEQZ0QjW60XR2nXM5hHRdyGfNLTV0Uv7EYgL
vRgm/U66BXGliDAqFZQxMvLz+8xEw9Fi/seYDwSDqcxObLW5L9ewGhoqeir1kmda+ac0F4Bky8Vf
8Nw1O6MzVT+QLeRSdYdSy7u8cRfmb0z7bfpKckj535Ft7o0nco5wxXw09EBQGQpNNJvBqZEQP4z6
1zq5k1DckEEDnxLGif0N1w4yYtPkdbTv6P0xSqmwmbVuj8hQxf1EMK7InFHEYS8HHmlvknZVskP7
tGvVAJ8rpzbvcxOM0bPablcP2FxMrr+C/R41fdDX2Cu6rSMmJx/J0M7P17LHPjpxCng7gLm88xYF
11Ym+4rQT6hR/tqJjIpTuitFebERsgoAAtxzMNL9j/eDmQKmlJb40f5ibCnNNG15dLMQQPMc83Uo
cc5lZiWOs35KKDo48A1+TW7QnMUKKoFbHl51UPnVF9ymXvIzmj+AeT11chD8PQGEBOW5rXsnG8AZ
rx7taWvA22qz0Itcx3GZs6+7shdF028srZKx5Af6p6TYTIS0rfYrl5MQYvXzPHpLifTD0f8Q5yum
UNNAjpmGPxdBqTz1zM/4HdtW2AL926Z4MQSU/4ynSMS2yGiDZWTnYKSDvUnXWtxNWYf+FwUQ1HTt
v6QP4+L3BaiZTcErM1XCW7CcRKlLWyyYQJV2YbRq1MkAcmMQlm0/YsnJ/Y4t42EvAPZIMFEDXglG
tnAA+hzqz2qOPsToLG/QdYO39NdU52ZsrrFY3Sp5OiBkNQXTl2UarPCi4mJ9l7HfuS06/fb1iaVc
5T1hnbHeOex2lgSWmUoqLl21KCFfFlsP0pYiHDwsgeWqMlHn7uRcRNQJy/pDwKLHerqpMnDqpmD4
ReoWLtwMMb3EE6mJWJxOutmNQxrVVz5zp62GZgiF/o/x/8IFmPNuc8OqG+pZXCxuJizjHiNoJfEb
yu69G3MtgN8Z1mJmfjVILEBVuMWwLycqBm2YnKlSq0NjxtGUYpTZlZX1HOrUjWszsn8TJgWp2t/7
A2Qfv8CMBhBDmt+lzweiNL8XHMU6BlDAflKLW5fJ2LXo5EwCZzUgTCZieFa17isnPrqV5W/ZJA8z
44UD1zRo3DYxyHit5LCRkUWEokwEV/WUgW3TZcWWOnaPkmma8yrNpO2w84ZU4F+JYhmqSO5OZyBt
C/szEPHWiHH2lv8QZxCCamDe1i1a2HmCZyHov+Ydcic494TLe0PVAzGCr9t0okhZYp0gpaleqj/y
fNrv3z/a2Zr5cwwrZ62buoHLmj4eRkIcz7amnIXBaKUeeJSOGkjZhRaAU3FaOd7GLSsgcwVLI5n7
lShno5Yq+ZoH17cm8dschjclAXco/0jIv5bshAofEuDLBK7RSnLOUjD2xsiBFYMsnMiAJeAi2hLz
m9AflxUG3U0U7RC27G6ql3ZqsS/jHoMrkpOVziVBIWxNlU66dhI2W4abIceb+efHlGyASf9EsSfm
++xTmhOjNCraGOqVXF/mj9lU5WPD33qgotLT6qWNiXVK8x9L6wM2s2Zeimux3HNczy1BxwQSLWyc
dEPUVih66BPM7L3sIw2FS2RZ4qiuBPnCNnt44Hs1hlNGuimwUWCpxhPdtn5lxjJt+OG15RsQHy19
BJgnTXp5HNOLKaUTKI7WykTf3hkHlqCa42I+tsf7JTu5ZDTk0mMh1BE/fIau80AVf1nDB2bPZw2S
Pkj+zKbnjgurZVIemPXz/fyDVx5cAj1P5g+/kgnZ0R3AyNrqwPgu3L3iO1TXPMVlRUSeB50HNIFA
B9pHm9NX6CodSKeMz7p8v46YF3MI1t1cw4ykXITMUT5mAyfJlYCBXoRZvLe7EgwMaiHp+WtNueZH
JU4tl2DE6Fu1zihsYLvv0eGhrJVdu4khJcG+maTWw2ptirwABrq7XNK7qVP1mSYcHP2StdxgAjlW
832q9aA742f5s1KfdGOcSb/wcZMnlwOG06P8dZPjDwTB4kGCbrWtM8u2h2h3QXIMJHHEEAV8f1/n
FeHFe1mqhs+l34Akv7auHwZY5YtAXSJlUjnqdfI/M3/wXOrE2zu5Btq2MGNRlBc/gRTbzEC0z/Cd
Z3hrdDYfhtU2k22RaNE/fOpjx21X3S//spf+neo70/3WdLxfuwLwV/dcfCkEswceTQGY92Gh95ia
zJ0VbAasUQ9Y3gX/Of9yPb/I+qyGiEd+DckC45uIAr9DEsqMjR/csqLA55CUSTGtZsXvYGgmetsT
Bcrr/UPuz+H7uyymZdTrMCge10uhuqPlrABDMszwzq//82d30eOQ6GdaU7Mautu8ZhLMFObt0Xn1
MySkCgxMscSIM7U0aJhkkHHFHxOFIRtLnJQspdo7MCzrLhHo8lWx1EjhahfKeY+s0/fuz4QZhMBv
O4o2BwiEJSyBk4U8O5xA75ai8jL0YkkTH1EQw0+zpUyW17rSCU7JYolp9ZdoIoviSuAI78EXtCnN
UzPuJlO2MaBfpyC0o2+086HQ9lrYHxdvBBW/y9SK4cOPuxRwPg8bwBw6LuPxMjgx4PEMGFS+HX/I
1ZEy+7bE6UwlrcvCnKuty8R+X2S1gZcfB5w/KbuniXJmnXwlNVTYhjRS3t7Zc8opAsTWMLJFZR5f
eGyahKuv9SoZ7ErZx3oSmar5p0xXJoum4NLtjbcxGPvSW2fdd44u2OZUfIQ2VyyFfiKoWap1b0FN
5fVR5JI8R3imBtHZeoeC/ZEEGPlJeQ5KJFGloOQzCkZlj7x2saZtwYDqfRTYDOAUdZ6q3rSn/vBW
homIOjH6JR0ow2pZgq3CT81fiTXbbsf0d8Yw9pKDjVIwR7oI2NSVYnmfPdcPw/xx/rcQxx1ODrDd
o7e5MNEflHF7OcuWdXhwD+WJJ7ZAIcsbRhn1h6H9JaSt++fRKK905l1zpt9Js0SON3gGhoBMcG1U
jrlHZaEJaTWM/REzhRsRnhFF7EhwQ1sLKA3/xY/1tPNLcCILrFdoWeCft+qp4d771s3WGgveoMPk
y6pOdWEE+xUrmWjl5AwQ30BZ/AEdWKnqoRWzzoJnnx0becHOHLJgdjGkdWKMevQ2lh65cePTvCmO
V/eV2IEbrZzootFt8dTWm3VBCtk3WDVO29W9nohJTRG4wzsR2w00Uf4/q8mmp/3+CFVHHq/zFRrv
KXxNs+XBnXqnv3eklK1ZNkr8c5e1mDVOOi7n8whtu4KnZff+3e+fN8975MF709VaSDF+tCmEOKhB
6UWbCsgzttHlygzofG0+h2yyVztY4QV11J0prl+Sz1Fgzag94OWDjcKObWOWgqaIEAUNdKO/TjOX
ZvuzWyNG5JjNjnpy2iz+X7l/UQPtZnPKbkWTrrxbWkvUwbF/T4lXT7IcudNsQUnLgn+xvryZ6Gn1
/JDbixUSpaUzesCYY3IaHDjdCZoIsbzkAdeNJEDboImcO+bRGEt0/YUcoKIgkZhs2B7qGmpFOn1f
ynumIx8K5LDIdZBZmLyP3vsYlJ6Ti0l7utpt9n5zma4DvZhU5BG421ah3FePvzmEab8968ULjn4g
86HyHqbGCelQlN/WdUJnaS2yjdmfWTvL7wNvsXYJZNJiY4grFcX/MWdf7I1aQO7Xic0WBrgFTEHR
zggMyqEfjXvHScNyY2bgLKeLf8u/Lt6r1cgDIbYxulirRSJezKoqwKgyWSJZeWzVKoser+MtLoAj
+0Mloi449OiliG09sVMKB1fPZ8RYMpJIzUCEWWCi08Bm68OhcA17ZpMNGBqqT85ruUvLXtyN/SfM
Up7B9o/EVlHmJZStChLHUFFQSUPRhc/3JinI5NsLJ7N6ulcnmkO6L8d69ATC9LB70WKLgFZkmoIM
pUZflGEODfjnkw5j2BXRaGn4l3cJgKxBam25hJVKvEKXF7g9CZ2HPgQ7q/p8zDRQ8Bm0c9Z14F53
cmtFPIulScB9qyvisyfi6azvssFzzBkGzcCge5YO7m7KqgeRW8JTGE3RhmMb5yZE++hLd6L4AP2L
MK3ZYnmE3B30a2WHpwE8czsmSVVlBO7B+nkq8SoxTZDYDVIqhEhx45YC5LsOKjK9Kfk+eQ4qa9s3
OIejTaAHe27JkVzq0ZNW4sT9gItUd2TstQeIEVrLI3yecefKRpfTm5iIupTuseTHRlwh0m9y6ZLf
FuQZYYZtUlaXMteC8gRwphB4VLrJOYxlMMolbtC6VM0WT9IGu+QD8HomI9n8zEBxDOhR7nH3/qpZ
d+04yWOdRbXv9zzJdVEo+ZsCubbvQQ2M0T/wxhwwGFajUCh6jPmP/B+s/8ifLNhj4IBz7cw/xwp6
L6kIEwxaFtWAFyH0nMooK1POSGNLBpdyvGS6HQeWi07c+zRigCy5Vd1usBdDUONqvrt7G/Gg+IID
SeTSf6UusLdLmvosH26rwETz5oiPBlGb7tNDM4yYHozZuaPKHQ+zp5irw789uJOCk+W+3nZDiPS8
bFvkePu66SsJZnzzh6ydpWbJAEFLGRp3hFuYhVdsxWVK0OkXwh+1Cj4dU9YnRBa5aaEIXfAl7WB4
e6JrrqY75sm+a+IbiCBv2WuKTzqynKVHpLgEOBnQxfPZRBOAwRzNY5m31s1CuUCOFj9pV0oHM9GK
odJ0q3ffjEDB9UxGktGizPmmqt2d1H1twed93ZnOuX2jr8Em8l97sjv4dSLe/kqUc6IBKdDLwB3B
oOh0cFMIM+WwR+YuB0km3NLJzYJv8Ttj3AEo+x1kpWCDSt3qVBMrOY7GffPwkbWxcS0tiX7hUsf3
gdN8kMeDo946AoKwNddHfRS4nf8Bm+NCqKbeIc0p2tL+++/7VS3YiWz/swz+aO352EdpryRk+2rs
pwbZ9lWfewYVEbWmdCmWHh2tGLaXk9NvbxGM5rZSiOfB1rVa1OSIQ9yHH9TT37aOsYS7Nt3mP6uh
AQ11NaNiKftsN218bJRjZqGqlDFB145uPWzyRql/bgeBJS9OJkJYx7jc3HCWerh17W8N7Qmm9eUD
wOrAg9Qt3/5EQOcOjb0hYWpKeyLfpB+HBPnddlQmyUbIwwkUbb17xAOayRc3NuOzmVEfkO3WNYYn
uTQHzIwY2Xfpp0aT7GPOtQm14nECHokZ5wSTsMzWeOQQeFFsmaIbaWxx3w0is/LoO8icEsQtfrx+
VF5It7QUvSfUoBTRMZexG0/qrP0VKUuhiQhWFPsgPiFQ0ofQJ0hckGgJXt+nojtyLK1HeCFdlWmz
o3p2bNV1ZqrKcepGJgPbVP8AZ6Lc2jOSonldHp7lr1ALi6o944n9ZgscZLHkV0her2xao36hkgaS
EWkHLKtvxO6XZ/uPGLGbQCNQ8Z04xLUnql9uhfhMFxNEdM/XYhuxiGXSjOP+HhHkCMVY62tJ6q0N
usaTOziBbqlRDCJ/yWNkI7yKnKa2qJGQaI4ZW8bIYcdZeOmQSkhV4KlXs3tbTERRNzUlcjl2T6BR
4cMkQ0zgQkIrDNPE5dIsCc3c46ytdtZReKD70LbJyOHvaLLXhQEmbjjz0Wp4MGMsyxBLOE3uNZHm
elWwz8tmXoUEr0TAwGpJo0Uzn0xbHvGmapMchw2MgZrP80OKryE1hizZNx3qVSUcJcYRTInKzOP5
9dBH+1M11MIg5JHpvTHkHSxS7l1kouU4hj+Qpfp86mlkkIUTCPKdyHB5uPo78E9+MMIJfUjRaCuE
oF9QCjHGtmPWzFrAwRkxRGYmdjtrC5gde07pk/GRClSgkvNApo0jC5EFIbThL0fojoN49vVWPM9d
3E9D9h6bKERLqf3MUocxra6Zh0+7PdNydfIebYf/WTYxQHNxvohMxWM+rao2dWlidvD3lh1PJvrh
H+HDLZ/lH9R6dSoVxE21EgGeEoN5djoPlESiIu8hsN21fl8DWqSTN6M8hLuHb1qqeyKscmc/00xp
ntNoJ0T6zi9uJj5nXAKDwOJIuRjvQ2PFTm5PcUMVA9H/ADJtix4p/iE7EFtmSPWTi0jnqo4GBf7f
ZTXwRTKNVnr2IDKns+I8H37B3ix5aPfVZHz3mEK4Z7KY8jDpolBRbOH6LxWVJvPgLKUJMUJxeZeY
4RuiSl2DWm8c5dSaqUiWCc0JmWGM2Be4LB3cT6YKYvCtwD4rwTXrUu2b/urjsWI8JMM9RKUeYiBd
ChJefZAFvOiJnnaqRSQjIotqYhtTYxqi47x744UXdrhp/sZ4ZJDwAM5Cqy2jZAhFqlDVi7j4eKDn
PCcJTP3s4UL/BAcijs+oNuRF6qNqWV4Qtfe+n6rJWAW69mRD0BKMy1lfIhkA5wnOcK9KzQe583Z2
tMm9DVQXzQDl1sHlVwdoV/qA0TfJzbfX1h7YU8d+U4V9mRD6zdCvOBjHtsP6TVHh97JxNhHn/zMq
xMjYZ91Tkae04UzCeJxTZdWvw6PrRIDP/GFL0J4x3qnBZaHZLvcVg/UvzR3iIxop91iQ0KVP9SFi
gRnmIzOoyrr9As8sGf5AMbCFtqez5b2sf+FRN+CmXu6Qa9deX25DCfDAzMguWnLZImDdLTssq1ES
BxXdL76/RTdfo3B4eS9LKi2tThBmGiFWnYYgknCIRoLYoS77H7z1mDDNXKyZMKntzbek0at4e0xk
/iHTALFZsX7t+6tAm/gcCdjaOzUo8vF0OoHLL8CXhcnGOOpkTh28KGVSe39odLZLjTpF12Dfk4LD
+bFenTq8+vmHUPEGSFieB1VHnatswulK01suAwxd2ddkyfkq39EGZFE4Ss/cuXfeE8f8CDgC0B0I
aFQ9crzsrv/j2BG2iGrAPZLcJjtWrjPgblgoodFZROtZUlnQ4zt/f1x1IN8AIIT8mGD7FTDhB82V
DNmH+AuOFXYV97IGEEEBgBCrUAU4qNq0n29Vo6BIJZKh+WDXbPpPQUoC6BWqA/d2ZiwxW7+Qa/JZ
caZrm8OxGju2z+5NnKa1RWEH67coKYEpfYEYsYYqZoiN9g0BpACw7Ege2Xz+aBvHCEn32rF4rmH4
CoRc+ztEAaQf1oDikOYBvR0iBZiFD2P1550wZaLmoilSLDd5/ipzDdttBgFPv3IblutMc9PRUOtc
N/tz7Sv0ILH17mL0vUUjvS3+cEgPTE68JkChTHaLsTvgQl+jXsU9mKjw3IoPV0EPPlT46q6wCgjl
mbbnyuSi66j6kKwAoZXWElmgK1156VmiMEyEHnRAzge6hN/DGhgUPdGp9Y3da86pCfbGiEAkmAmf
Zy56pnafp0YpP06bob4jzPDuolpe0ZrQKYqczwc9ghKh/KamQbAcV1tKScmtUuNopZtAAckUZZNU
BbL9arV2pmaV1cwWn2aTm1PWu54ppn4YH8fAmWnyUN+VCxyUTNml3gSC+fu6IrM2rIxy3ssxkzlC
j4qItfmEDdZe5QRuuPqCmEaEPj3M85HEC582gOLsBFZDFEA2Wr/Aeg/TucIEzFcFX6X9qlQNC5ya
hkv0dKX3SMqrOUMVv4yuyGddTYsA33nkbPkqy56CETrISdnMzw0cScR7Ev7gHTe8okOHshMdEtMd
R+gBB2LmHE5x9kmYr67tyBERjHOl80jPTKKxY0oSB75lkKmNF/N6JGnz7hlzotSrBgpnuCoYCC42
M5ZzOqtJOWnUseskGD5LpMkOHdmQoie0Z4ocJKCTIpLvuylm27WA3PW3xC19roxYJx7OfOh4Hh7U
1K5Q5hg3wGZeCPFfvLRcvRnNFFRCYMICR9+p/CEnBaSoaBcGJMNjjRHn2k5i2Yq1OcFkg58OhuGd
jJlO79riycY61P5fgenHXY28kK56Pt5hCVHv1xH5Jg0Ga+QBXOI6+d/VMahbFt2bk8WmKY6lxrqK
iyUV8o7hRz5LoAOVRtBAWfQTq/mzQjSYgKO85hHxd+cGkiboky0BvqERWjWCwDhp1NjGanbeaQ9s
rDLZBslSN9asz9r1Ugq/mi+3zCDkQ7phAO6MPAd/zSAxTddpIlZ2X1/UUQhXrcGj/8uydYjYZ0g5
k5CFBWWu1iunQJMJ7YR6f1n9RJew0O2M5NCG7SecAAWiHUBja0SE6NmM4E9OvJ3CGNH+Vbj2PuSC
nes9KGfytrylCv7FqWkrkhA7g76EEKF/kdofu2ofFwrdxVMB8UJJLNbYpUoQ9aHkX7l8BkdOq1Mi
q61/VFiR77Trb4D4WDedoooXDZ/0bPffer+GVgtKdfaV68rRZtu1PrWoI+1JB6am65AwEmve4vhj
aJPw3GErLhJ439gNsdpO8UfiaYnrX+HhrJB0KrIZpkZZT/ltBo9v9WWoTJryEFjt7N8cqy3dOduZ
6Nx6rI1gnq9rCOLl0gT4YDremiwwz0hOCnJ2/qXSDG90bjRpdxHZlr/T4RG/Hd99tWtsnSy6hCz1
KGPU2G87Rrw+mGu6+W0wVR7L/hD8C1PyIkosrF3mE+VD/oYLo4hoMwAaiS5Q0jTzKmr20bedMABU
S7IAvWZ9uDxAONos6K/+Ux5MEXbCoNAomd9aEIU+FoKG5z3sTzm0ZrsWf0aRVwRBYIt/PXFOzkcm
2FNlQ90zF76Xjobxm877loS7HOtGLI6wpLJAWiEk0zpfmSnUSdynhrF1dnHmIlnWwgn80FpS97Ss
a64zGt2DSe1QcpntaabNW2knPQgUpj3NIe+H2ybWojYNhZ7yzevAC+qHezpKSM73ehg+GJMI0Rov
Va9JZdIxWOC8AKAvarLNRss+RmkGyuvrFDxsuPklaF2c2uDNxQVjKmSHJ9xoGWApCgoCQPWPfP+7
XIbN5YvgaeDXsA9XpauRdh8ikUwUZhq92DjfXz2hqIh9J20sfAhuKjZmH6TkWjCmzfA/wRrQo5jo
SUMT+XRCj6FsBFaikadXrOC42ueIv1PnhbtgJUy+LDzv92rqlLcKVw9kDEBMGBgrUiBfKaPrlvA5
8e7jbrhQKWcb4F5VB4LXkdtz3vZbDQTQ6kFUPHWRWtK7Sxb0TajEpq26qPwovb2sinP6H0BT2Skp
R3EaC+BlApsXEqLxumwV4kjlZxXt3Si7OGCD+kbVAuVtM6EXfGqs1PdHQroSWAYTxn9qzCQ3l/ZM
GmwauWdYpSYcEmVQflkrzke/S+n5o/PgS2ynqgZPwLwKF2Grx+/jJAeiYWEgRvQnSmHAyYiXjL2g
I3yKyKoAb2rHx/dO0kdGCNNAHclq725X+waYGrtWMQlGLj0RQTyH0UtQ/uq3o5DUxQiSrYRnLT8m
27F+/H1dGUYqzCNhInlOJCpUtycMiFro0gW49TdWgY3Jhg4jJOKPccSiBCdkzYISEE6PbvBwVaZR
V01z+kRs6jAezmuvYt9kE8+WxuHDJeLDI8H677JfnqzMOGg1nJ9LQ/UGZwgDJU92U2ZbptTRbqDO
5t5oyjDib/eDLWWyYD8RtwmaW/H4F3iFZVvA3fT4X5M1H9KfyeX0K7Ahwfpfcrjl2ns9SZrbENXb
2dBe9PVuUOnJOObRDMd/H/7cqPgJdtS/7euzHRacUEfLgodMyUZRdnEIKZ/hemO4/uMMlWcQKs3p
IoEcbTFeeDxzww3cT2yLODO+gDGjLvkDLzH1lfUrrca0QjmESEv4m2ps3BpexNjh1EVHuGRNlwOe
zHikbz684VxAu8GeKBB8NygZ4qzXjY7AVOLVTKlAmmpYCh5cdQdDe51PRdnSSnWxY7mh3Cwtj/8A
9vmNPUIQXe3VcgaDblrqPZL0udy+vBEoqDc2gBUR9Zip+hvbKQ0NB4Bc3NONlLGIBKVnJNNAw71E
A+0EtLo3viep4giGVKbRA3YEii6w0B+caJ0IXsNupbo00mz3prl7RQA69uNj2NrVanWAuzZk+ICH
fLW6S9qVIi1l+axzw2Vfm7+pnOe48Kj4+EvtDunM7sF6eMBXQpy893hf0UD1pO6GzUTO7+aamUcB
/1MvtBzh9lzfu8zm9UIUOg2YS0g+j7uIgmckhf6TvrbPmMqRqshhGoRA2PzXCM9+Xze+KrnmfGgN
Ail9+YdAnNbqvOkLqFT7bU3mqt+abv4/jJBSYWI8AtBzl9QMQRYUxR2ZqB+rBeXczLbaeFswfHNy
A1gBfII02YX15+voPQ7lJiEChkAnzPCNAOxm0V0VVlcRz0AolONHofBYa82z0qSEkl5fHxWlrWEW
QOBhxJ0Yu3Xfs4k4jlqLsMTUgKl5qlGOUjT/YUjAc3TfCN+Z3Y9KT173qKfbISyiHMswr22FmeOX
mgphWLvAzsIjJoisNR0G7A5nUVnr1MD1byvkUswMJchBndJb68uYnIeH9cdku7ugzymUn63lIi2q
2711c4jQj6u9UHdlkCxl3oyIAFXd7wNoJFB0x81j7RZQWSv198+hq2bHxoN+14GMYY/oHfB6hwLq
1YoIatmaJ/wnX39Hh10sDidjxQdV+egehDwhpQudTrFh40ZIF1XNSffoRrT6oP+Yn+iMxD7FuxGZ
W9VQUkx88yS00zewDQ9I+mz3qFlJcUVKHl2200GbHjyPzFTi4vIxFxoh1ENrjQrEJyFSe1fOYjcN
m18/23ESDnOxttsClW6nueq4Gb4WOj1bUQqUoAKaR+gombwE1qZTOlblnuTeuapMf/hHdV2wzpjW
uxs9cy1tlxwO4Y2LAFzCxjG8mf2Qq7YMaUuMDGLRvMDxTNh3Ky62waRltKO5qzpp+N0v3xJUujfZ
T2Sk4agy0JgQeb/eOSGB9KZcB1WikNpcSkI6QM4DG5LRdrNz00W50C+WBJ6dwoiEpzpA79CKbpcA
8urwM9SPGhSug26PGB34wcIRL1/RUS8LswqT7lXDu22Tgw/dpV6VWO3ddaJd9W776iqDjncYVQee
HurAOumtBLLMSP6p+R2sIIjGbfEuTAT3bmLz2EsLWFasP1Gn30dU4dJY3imZxSgQEvnaGiXT7CxF
ONb1exUle8f8H7kFX6AxvjgUSgQu6UwMeXJtfSMQwl92aSMqoHZXBuXFzgMH7nRROb6hz5V+YJEa
ZDjcrmtuN5Cxh/dpTYRVhlKEOBbyvJo5YcKeA3fkxsy2VZ3RpkzRpbOspMejdHKgaSwi+nEm5x9O
JhNfQ8TsPde4tya0GJXtE3tmKXOm0gJj4JnCAvN9tGzDMALo3Qc7PaBaitlsybAVU+y9wHuKZF0R
XN9VNX3jaiDvfqC0KRq/gZE1Asx2XB8Xjvn1bY6ZO/iGc/Pg4Zd6AnR7XfJfKClqwYYzAul9LnS7
ebqAlAhKte94CpiGuTy+H7sWlPBV1mgBl1WoJkeWd4zsvJ4KP7+d2CLLNukA332gyJlRbJVbZYsa
CldHQ2H7eP15fNT4fOyeqaMcuJksRtu0vOwzaHoqsGlNMbDnKGhcnSS4NNRJnZ9zW8OgrJmMFE1h
jZdHBTgT4YP/Tv64R0DQHacofdLCn2+KK5waptyv2yuFGOlq7CG4PAWE6vPeKCysx6EjlnlI8LXn
qLSmuNmQoMHWqnRPvgXM1SI7jS279uEniVRIR4B+maaZ4d/pFihQZMJ/231uZYangsXWcqZeT4ZI
nIl+LUyWMt/UAKB/MHMBu9UbI3KnpFVqQYAZ1udFRXDdD3hGWU+Zl0EzjzLl/UezJPqG+SLw8P5K
avg04mogoywyDvg+g7nWSynvLPcQCQRGqoP7wkNRbuyLTbAhNne30NErXtQTlGu8sy34rLEKo7OA
ZFQI8L7H7haAZGp4q7ORzL5Q2XZJWscor87Y2HzkTyUQzTUW27LUmKgJbkyA/2jf6Cne54MJLsbz
CLix//O997WIhRcuY5ghR3eXtNmOX9cHwE+KoxMTLscyJFfRSqH3lLUbWkXA/nFJ1eN8Ba7zRK+C
IUrTMd3pOJCtUR6bLmB4r9lMum6NRRUTQjCzW5JdZAB/W+JyR8k8IndMcFxnbZ99/m4VkeYtEeHF
yoJkacaCqJ1rcuosd9JcroepHc/2FuB1ufcbcvHonOLbN2/s3Hrxrpkcc3T0a73+EjONhg/BcK+p
4YUE3dxfkNi/c5MJLZxogfzjqT2lYtWH8fxEMCxhh8ndrcr0bTbFwxbhUuTQ8cjjvij1vq0rI6TO
CRONhxf/kLIyXvvcXIt21ACFVJEIthNQZH7VTHynV8joY0NahPCGD6HL6aCC6cv6QRDOPoneQH0i
PLg5npMtjs+fyHZxTjCnJlyzeMYkzanmk7FCl44fhf88wMjwtZjLm9T7kLPVJKmw4y5VwOA39mcb
jOkXXw3V766GGdPEZs92Vcm0nN0NbH1rwhLkbcm2LL8AabI0NZH20vGKZsa37uxA5ZsR2o6Y8dE+
ufJ01QDPuIGoYQNNH/BFBe0VttFKRvSARYCmbJj9PQDVFG4IOpHzNOPiOSK3C8yd2cCLwZq8ATHu
wqsG4b6LUwUPz6+97G2VByN9vGBRVbrGDFUZrgR/oHUu8qTovhx74MOJ8Krh/DQaZswVxCV7/wUK
1J+OGe+F45rSQZTCifRVaoHk0jwHXQMfKBci8w0xsxfUCB2QWG4PCqMmi6b4x9l0gAuZajJZRqRf
Y/zjhsEPUsnniV+t1v2iii79A2NPtrG3r63Qa88RkhL7OtGssnkau+eSYLRd9+iE3Py3irU+eg/8
1Ox6Y9NgGI+0yPZNq5Sz8m6ptGI4S2hARiktAXKsz2G9vsX7iDvc6ouM+/LO3Sc/dMgHFRoNX6m2
62Y1Aq9Wz7GNj+HWmLm7NyQi6EWwbEEJ8Qtiw++eoleqAoKfml+hi5dUz5N7+STqLYFMBcwQBz0k
77qMzKBijtVOU64L+DOWqci0BVlbjoXj3+Ls8rV+QCsySj/kHGnLKtWkFR3kQy9qGy2FGLtfJzGk
M2xumUBZJldEju/NO+4VHlmYWYJYQaLn4n+D/cFNb79xZQABtY1TibvYs9DpUyWxSzPlglJYVyYS
r+URFuHmxQa2t81Ubt+9UXGWAFzM3tXPj7V1bKvuE/Oyz/nXyluJy+aRpwys369azPqtkUQNPyUw
VSQX+7DzdTdWg/8vdeU3XwXwbYSO1H5lDetpC5mac7yaTsDj6v3+1zjIU1SzCEpPgn0qmi+43yxX
wCngCaNOPadG3w5Xwdv8NZLF2ww9GW7CpvrSGteW4yGaUOwhp5poYdGL/9BrCBOnwYPfyJfwJJEn
t86mDSoM7FGk6qE7Iv5r8KBfm6z+gjy0CwLRQ6afcJs6fzYIAgJQNfZT1/qItTsyRlZOfe9cAYYv
I0wvtploIbTooNyczXXW4BQ50yKlEKPbAQL8nmLFKP7Fcg16P81arwJ0E2Xml8G6w7XvvUd4snFn
UyRP2kJdVxSGc9AicrpWEdaSZfox0vSD5pt2C+48NU8EUxcqZF0Kjkvk7AEa87IuTOrjRekT1A+w
usXtWxGPbswywenGyPwWZXKPomx3wqFdAOgfZDQPATSI0EzCf0yxJOpfzEzJ2VQdMJQsupddKpKp
e5uqRHQu/RyT0+izLSLrQv8DtDU98sjxGEN0rWSyTMWswqjEWLzaPtn6Omj3RLqi1B0GXpFAMSL6
GeQknw8xBE1Rk23ZDJPQ7pWs2f4DGPRkidYRvLOSaI4SPvupGHaBLl+p43iZqzdwmou7JYIboY60
qT8losXzJ0ocrR5f/N5cOYq9nVDE0UUOSb4UeGdLIAnkpoulBrdOfqFwHo/AvkaNyKMrOgcV1CRa
VVC/fCcjoZAfbZrqlNBGShikyoHd8aus5vh38ouEUdTLMGLuz5ieJS2F4uAIhVN3N6/FMVfklncs
1DmoDQ8/8FSYeB1fD+xQrrkGfYA87WvF6bjM1PzXqcJpsSP4rsjwnP+mhVilCep0/ZPQ/KPHhTGy
tM6ilx+OJfPKFl/NuEXfjraoWQAUvz9X72VycGtQejYm9Ah7m8v+t5MtZjd2WEspPG6ZMUBrzdIi
Eo+zqZXuFz5u8JKxAEsjtsurU6V8dYnFiZ8Z49aQ1KkMf8/85sxaackfwdYoWkyyHgZVFi0S5BgX
9wyugzeljS5RP1E3Fia6AVAGj0bIfrWZT3kXDbKecUa/hvDc+EHAgP6LKdJhyNhwGv0zh75jNeBw
uZiOuk/tuZy44yQnsK37umc0umNJSLkQlf9o4vviB/Hb7QooJK/vqenm+Nvx7WOev1nUrnu/JjmA
sgmFrZcwbiHM9OiBtcjFo2O76alpjdqtDcHnqOlL/W0FrZfUuAgTM5UYaEU39NjDyPvLhnGtX0YX
UM+PGCcTLinZv9l8tfgDgcTjqjdfrsCxC1GxwPNFl05G3YR8KWBF8fHxKK1xu/5tcDZ5j0YuCJ+Z
Ttl6FsFvGu4WErbu7PAhqF35m4/0pAPTcfQmnUMU5PY5AqbJHlsff1+N6SX96BO+Am6yhNKk0X+M
OytcUkpX7GX5vQIpzk2RwcEiYLr5RKMA6o8tejacAPkGl19gBt2S1QhvI0ZFNxR03nXuLepQ/Rjt
HJHa0N0qomuG/Da0sWvSKV3aS40CjHdCBgtD88BiM6xYaflvRhrOjJyBUfQr/+eayAcqd+cdnGdN
VWe6Jjvq+P7OYMQQyWZxz0vzfOnDHsO8AycqFQvKeZJ7M+76HTeWyU4TYGXM1PKrDr1+ukotnug5
kNqJjh5OqjRjl0PZ4K62NAjD62cmkYTno5ElY/HAdjvAp4UTRt4XtQM3KAEQWtAlMwXSemhbt/Jk
UtfwOV+ss+y2/qdtHBZAL3cnsLqMtGNRS4WAMpKnXD7r0/b6VX6cYprpDTjZH3D9WpKbAR4jTR1e
RN6QgJeph+LQbEPqsDJ7Sqw0ok7vc/vmXEUTRr4HFotFI5HIzqUKe7CwBs+0yDIWszYOOvWyFm6m
1R5uU7n7eX+9QwcSSQBywNSgSz9UEGESvDR9R59489qqDO7yglrckVnE61mQycCwt1yI8U7MF6+v
tEHW90y8V/r2FCjER5Yxuy/PLBnIxHAiZJ53ApasFiiXqQCkwm2r/ljj4nYrBpCsxpfWyD6TiGX/
11eAwy7ad0vHuAiIFABx1To3Qvg1tWptyzN6HgU+JwkoAvOayPE6DyvhdFPqxIAN0OWtf4MkNKL9
YvKv/R4pow0LBaucN+JUPCg6ghlEhDVmZ1StPpoyR2QIFvsk0Av3NHhNWNIhnk5pXCdzws8HUcgo
9O4l9iN5O+gfoVBiu2237iOBJalm12rMfhieE/xI3Oog9SmN3VUmcgUm/nptvD9w6VL3CQWDbnWl
Tc1P4uR1h5hMUsd4W0pJ+3aNXH71cWZTtqLX41FMoKe7sh2HIqAlGiYgKisZDQapSVm5n6Wrg7XD
fcECFRCHvIPNVjwkk34KQytR9BnBxCxMidivO2aw+6n0nBv6plwxSrd1zbfxvpRPLw69PHYjYIou
LKgmmfc+BduMdhBFa1K2gVee0+hwmEM7WfK2HibX4oHo0iaUhWNBHhWlhIRl3g2/DhJiosrS0y2K
gEx5naxm4ZL08C6mNEAniiJIMBoL9sz/gDlrS9fXhSSplu0qkTYCKf3gqnHzmkecXWi074bccM/f
XIJkRmpA8df3jiUETSZnFOqpyxrjrNbizDwzBtDozsSjQlnNIwyfGAlTe6q9cVUflfc8KCq7txRk
8JxHv1yG/Cx+8H0Wl72FbhGKiysouAroh3il+XYyA+jbA25CAdigzCmU5ya054577WPoYMzwW4rz
1gTpIezUfpaATDeUQsjgTp8WoBrgpA4hBUZo0TkFHE0r4hie8eu4WnuplVdr573sDqxR5o+yePLg
3zOOuyUCW5F7q6tKN+HKDtig87cjC3Zp4H+hF3ScEnpvCGlpNjHx7XiG58ZYRzlQLajJrzNmWv7A
cLb5y0bxZXQpyEOTjxL5NKxxEyd0nlgSsf5FuKo0mNgldlkV6t+8dUvpmoXhjMSovyRfLEuuwwRz
yEKhQTvuwbF80j4ylK3jsYWJCgJqIWUvZeWO9Gpi8+3xaRYimEq9aTN3f5kmzQ216DbkCgrRz2rR
qGRotHX4VyJtZ1helOfW6ks5r095oVNGxlI0EqPTzu5OkEGrg1Un0YInmOQJHtmKaEkUURqLK7El
8rthXjc1/dtg1H6RdMuJe8JT902xQaktbjbD+ql9HqG+BlbWsJ9zrKIrcyP9gLcqSRSXqYrQN44d
r4Ao3qo5gSDAu+y9o0JFk/PtypuVJ/nFED+s7ObbjvIetxXJ53sMQpcI2bd1d2zuntKEm9beJJsp
syS0/w9QGoSIfjQ1GJlU1q6NLk+PxLHnC5UNY/O8qz62hKVkKVQGMSubnLwe8mopAhD+/ttfPMzA
Km8ogiIetC3mU4zs7Ch587Z2ncw+nQoKm38y8Ni/ANE1PR/tpgAnhc4Fo2ewFrabXc902vAzYDNZ
rfhu9zGiHe0hEqmxV4Iz1NZt4ev5Dv6Nd1zAc/EZjEgLe+GYfmb9J5xpfC458JoZwAxGLSZPn5CJ
WyO4AF+L2A7IuEmdCHqpZ/jgXeIt/vDtbCMWzCuLMdoaK+nwuo1/nmZjQfyVo4FOz8s8n6XTLe6h
J85Sc0tNp4kPj4lidrj55g7LRokTHxkIIlMnnTNyhq823DSngkfJ/gbYa6NLfWOAIZSIVmwYwron
U3igKBrQuBPtMZ3zEiK+OHozQx6rCkleaSlBjosqkfl6MCNlE/hcC1qekZl+AjSIC8ejEA/T89iW
+mKcblmFq3mjHdIZQXMg8XtSilPozKn1+zQTW1RdEvyCsXl4pUiIVUPin2h03TPkFiE/jjCXKXsH
4B9HCyDph7rrOZ4rmvfUNLYaFhFIsXm1rMoQwhp42Yq5DcxU+knEqKYWF4iSX80VJj1oGUCuR/fI
terwqTijTj+8kw9TWm6kFfsFYnOp131lBzQy2vxMK8R+ZYRw9oqjfLwxb/LAiheqLPUMxvgMNhQ8
sZcgR5kin5rFbCkjGpzwAjlVAQ1TCIcpat6xsXI53trkOZ9j8U2i4G0LjhsIVrvqqfFWvHMAovbH
1BE+QoomMtU3jxFoCMzfGdfBrIcx1b5HxPpKf8vOpHCoI6wC8jHiswKfcRuqyl7mPqcJlLmwVLSh
jmDOuocAizYztwqObPPd2/dxfrBHCLrVk6dBJEArSoKVZNG7eW1Hdv6Sa/LsVGSOlZkNqMetWSWB
gdy9fjb32z5Yjixr9CHcbJt34rqb5y5QTl2aaLETKX206doUAdCBSOo6sBHr6PF4CZsF/oOscJXO
v84sQFbn6w4NwwLfITNqSm6/vwJuF1ug2EREHp79tBWLl6wIbqSY4cnQ3IiXjrDkVRgBWg3yA1hQ
BW1ksH7xahmkVNS/lD7iEb4a61ncMPbUgPLbPUOdGMixQUrDnPAZ79ifYyESvEBxsJJFNvaLOoxz
ZHCv6phXybZKroxIKT4aIXAn0lE/KsXx63yDsTiB2UjlCYNTvmYQgRlrn02/EvVQtaep+aZ6CDMt
Uj7PB8rS/d8U/SihExj0/fTT6MlkLPvQnWKepceVO1LPO8FmvA1lqQyc3HSrJTm/M7JpyBixKKpj
Uc3zQvnxs4FmzcDIOh5GLsCt4m33HVX5jXj/n8fInqN8EODhCiDBRIldJzF7O5n2h8hWZ1KefB0O
Wdn0IVqSBPXcM3ZE2yv5K742EtO1edXHBtDJWOQPb6YeT3wcIG+RkWfzkOvUt9LBwefDAljKINme
JSaa5zBev1OGmDDFvm1yrV6z+XqYWgXOX3A+dcpT8vKTKjmcICT2VrujsEWKdhd1N3S/7CoX/BAh
PLf8YKTg9CKGfQu5YVrU6FoZobLst0F8JvJwc6PsybbU8WiE6xmhg4dO8o3Qn4vY14pz3GtvedPg
j8DefAwI0PjC4LbWkkpXWgLSVu8Hl395NVQcwRnFKuGIeXXsbZmgsPiImqIEwqV/aH/9JU5RUEbO
OY9OCRbWG/eTe5M6Qq0+6iKzZAeIvtRuV/aNr3NYT9HvaRJ+VMdDm2eh7dhxrNns54NrI7+qO1MJ
5xCe4Q/Un4UOaUuj9rYzFSMSf8i82Kqj+8q4ucoWKj5CzZesU5KzGUreza8DhDyqb+cSQz462Muf
v6yBodJNmVz7Wf8Wq5n4Q77wkPbdA2GGqOSsS/ZCx10uSi07IaY5gB4CZx7wrNWOHFe5UegZVfAl
93vrRV9LfqUkgiJvcd4zGoBusu8nuyxOELqe7NNmoH6iQoJdvre9+xDhWj8o/Vbv53rjnBoDLCGE
arUnm1iRCiPZY67+nKp9tMwHfs2PEmHCaNGe/mZrscgQM6NOaZIvqj8w1y9R3awxwER+Q1yTgnSA
S3rqcyRjLMwyCb8aRwB4cH0aOkYg7s2cgncInbrFCRbu8p2D2DYYw0rbCCA2cAnINqpAhZv4oxXe
k83345XMVYQIH56lKZ2hKz1SF0MNeoeDZ2xdlIq3ShkAO2nKRlXD/ep/QIXh6stNaGl0c5AccwWf
uQ3ycmSfMzxKRqHIi9Po45PFeq+MpdKXteCY8Uea/ZHHOTwE0IAWgsBgIaNXvzNSZaLy6Y21gwNe
5/3pFQj3vx+nQr8qXsigDqW7OKh/HaWiQnTJgtqJjoWKFpnvZMqsxiNI+yMdm3DxmfbRoGk9EZbO
ygXvMLKtwM4u4i+n7t8Hkdtbnnq539qY/0rz175/Nziinn2JhXAYv9CO6la+dK9qA08OShqCl3/M
fSCZ1RYbtVb68vztceG109rR5owT6YkaAxH+k2IdqGG4MQZEUWPfFX3qVMvITn7PNPwg4CSEkeSI
GgN9cDvCpNLN5h9baFyxkACUcDO0IlBf9CxPwaGg/Mrs/xr/Ct3xhfF7vDmhr9pjgcODjHFTQ3AC
izju+2f+foYegjoQ6Fh3cvBX4na1yQr9mM9uQtOwJ5JNsOxx1WHXB2qefejGdHZsEEVZpaBmxAi5
mV+aELmN57dTFO3LitLLW+EuKmB5O1Pt9g8c50tjn7XsvU+eD8GEpm3P07zKw5yZ0ah7e8QsALP9
5t5P8j/rM1mqRqw/4fuSo2laISsqcZ7ZaQCcUQRaa4eKxqmc4eZmljOgPEhNrOw+BeDtnEmyuv0z
mXrPowamXK8jZjApR2IpfKODnJDcUfSwSUlknW+tm4f3DICZKDnryqqlnfMYqhnWAOj787DKSqiI
LhTOxxoPEXJR22mwiNU7xzz0g6Ve63p+K0nJP73UsYB+IAXwH29VaphM7R6G574MbCNrn3mICJna
59YqbW5lOPWdNjgM2Nq+8kdakEU4GpwAHjUsoh8ST+zHcUL5BSVVP91lLh0uVqlG0Bx6zjbg+d//
1GOMMpf+WU5ByYE+gOywn71+4Jv/Ok3qF4TBk13RwKpzZrqmXJT36WmVlqD66Gy8cmstQDXs+LeL
sY8owaoO9PCTVZD5hspFlfrEoYoQq0MJ8p1ZXHKwDSHZ1yUkrsW6qOmc3ittwToMPEjOZ1EaXp21
SM8aaK6QfP89gpSMQkzGCjS1rYGJOnaA1biCwpw+E6KaAiQUMHzXhUWzsSqMtkRnpz3z8Nkduho2
G9avMdSJzB+QRou2TNTH1car+I/3mEjOU7bXKyj0/c5uPeg+1yyDohcfx/+KSUDzZPzcm1NgX2MO
umGMAT8d65sSE0cvm3Vrn7wW5JgJTz7LrfNenupYhqEftoABOZaOsaT3hnLAObBRCHU2O9akFt8h
MyX8KH7A+ST6NpUHWWvIk6DGHq8YuhbKvXkM5SqGEccRNFH55qArevH0NBojO29S7AyQRcdflglE
Ok3FJXABR0swxoIXL+Aq332kG9R7w4jnZ0PGhywOJoXE0PhXnQtI1k/deh49j1G5Q/KcEKIXNiSa
r8L02Wlwxovo4pM4zxe+RyKNZaaERXUs2exuIcSwEupfDTHwO5CKXIu59okJSY/I48vNVaypab88
rPyZNxmnXKfje8NJZ/5Eqf4itRZEA6DrvRHz69viCzbA3oIiBt0WjU1dmrfgmw4xG1M6alEeRefE
vvLXuzwxDgJuknSx7XtUdVPAvvaMdSMJDwwmDYJRsbXYbfviIgXVW30jyCPk9y7K0TaThvrN8n/x
rcKcPbidpen9201VKLoTU5RmEOiOIV09GrDzuiPKNP2MjQbD0ES4OET5Ypng4ICUjg3/lsV0k1Z9
o4RJ6ytFCxA9j8fxmzMLcoIrxlVDgmPXJf/ld5ea3nTrk3m6fMQpYP+V8HQoajSeCg9gXIzXgnib
uLNr/N1G760de6iYn5utf05J3cbOdEKODYGUTKJ8R7efm3DchymJRIEWwmRaXl6VyPwVwvuZfBYu
LwYP4/1aUTCgA+lJ1uJMU5IpgWL20TKF8GTR6IRc1pREY2Jp2+fUfZPKO9Qx0etaTORJQqa+itB8
6WbgfC2jAzz4gmw7Y180rFpoT/g6w7qJNAYsYxGp9qmM5Dtrvabf5MtjcNGv0q/YtR4KgOyrzvfQ
1AX+b66tbcoaM+6p9+GWU2+AQ/7PGQ3sLdPBj0gzprOX+nTS5JPZoF3YSdmu9AwfvbZ62xI5nNGt
+7kMINpG+NmnC7YwO9jR3Jxacmj2Atn/FY6mlQrwD5C3e4ajiR+8BQlmyihAW52D0LwP/GHWkVgG
6krmFzYSmVmuEyOECUMUUvzXIhqs3VePg9l4ThchrVGCtKR4ubyZimsCGfueD4eMJfstfOEPcHEz
Eu6ejWxs42PDKBRyhWrt2QK+/f8jjZQW46+JQ69OH8fT3eW5bvmpESrWgdtgAK2ChRNoK5Cp5Bes
/GYMJns4QM1O5kDjwvQUlji7TyoiIn+lWVVN3oXUwgnMkKWboaQUWfo7n+3iD0/kWcommCIWvnIW
mQzHApq+25nYn8xuLIWJz95gT0lVCH3roqkqUJrNo9XTbbtIeGUNIRQaapt/3zX5pdv9ya0kMjHr
zyWl1G1f0o2OSwtSk+X5GBSmoJHDy4mEtUpkcPOrgaCC6n1FQEpcegBnDnUSciKIPJNP5XTqKqRj
ejvsgxqOBFfghPXgCOduephkD3tLumZWGRS0MAkliQX80UynRjylnUgrAkBD7Gmo3vbP+8St6t0J
wBIc16UAN/xHuHWcwtFdtsgdVUML2YfGQSlIQKQuK7sYX4lb0FV8xTIVowGkuVMOtS+lnOaNK2Jz
UqTX9jxyuXJcihZ+JXIZjHsHE5AjEIm5oCIl6wxVT0WgVYyYUjAtG1mSEmzSWSOA95TpHo/dEzVY
gjYKOFuhQbsR+uTJQHg3/QEwoX/gnIoToQxDNoMWOfdxW7S7fZMcCx9+KbTwXPVaaIFpJ9p3qSe3
WG9pwCJQGsckFUUu6g4Ul1LyBR+sBfngK2LEI75vzjbVM8MnbGzwEYf3KfpawioU1bJgLQEJjnTq
pCaZqqty14yQdKCfisQpNLYZsH8mQh0eGNR8A/+s6wDfZDHpEkpmson86JEglry8TjQJCIdpDEuI
96Tqumadv0ZhgleaDCx34IVrecURCA6/jtF+3+fVY3Fq5UthzPoz39vC7pO8sIB+nMyhMZpNu+Dp
/7gpYzK1ff7fEbForXBdhrEFW8IsWUnkyf6wsZGqG26TSK6nx+gM/h7d5tJKlvBZWjhMOblkrcpz
cPTBt0T0JfIZsso/I1zdNGnDtnxCf6kuvoqKzPzwddgOLGX7DR42Wn21WZfnTwowziDOvYZ/vlxg
+4FIgkTyFRE2tawJwovTRmRxFQOJ8+fyR6FKtUpme6USHAf4s5KXEvWsQyBB7fS7r53ljy5RDPLw
vI8ycwNFE2b9Sfs4fglq5kx2rJuHZJyhF7OyNZTUXopufGwgNJv3hXS8Mb1qC8XdubN7INZe3uua
SeECe69uXxUFpd6hToLmw5ypootb7raWFT2Ra/ESzTkBZfT1cu8nRFHJL6DrHnfHX3cmg/dplxMq
p6M9Yc0NJxrRYwBBuBUPcrUw/0jh1fnAJfZSxvMS0J/2n4+vq6POGFiNDRgHB7oJa1oh9aDi57l+
a5Kpkgt4pld0jRO3EUu7Fd2SkCsCMTUr0C9Gv+NoITN/7PpzayoPcZ0rDfTapr3FKGXlrlzArb6t
uY8FlJZ3/6915t6GcEs1pLjZtPlThYVH3akp+v5TeZi1Yjr8mX6LUc0APvhzW+nYCxjNmEKWn9jD
UQCZlfArd8cAGk++ZUcG0Y3xXTV7Eil+GnoHbjl06l3DrkP+hG9Q3UKgw1g3B+acxLoV5fYQvYwL
/OCX7tr/72/eXTth4M9yLipDcAeX/CXutgDAfVg13tChK6QUpETPqOZBOQoJ0R8jttSCW1nUtb92
HdSowNm4NpAEyp89colnZ/CTcvN+ISCY+0VdEBLCBzKiwwmFYnvDqcqZuFGy6KD5O9MIJ8y11R3N
6SjrunWCOpJkip0e+Ol90YAzqEJIBwflTgoj9tVSn1jaeM5OxHnhXctx3FxYHV8H7d1Li2KE40JF
M21lgxt8MPBrYnAUUKjSVFlD8IN5Auj2bhVTtPY5rYa2909Eibb7qvHoRLYL43Rl8T2/fKlyR0+a
Rh7qgLFtv60D5SDYC4GovM6CVykr7/JKeyB1fSQ55XOrL8WDTSNWOfVTA6zB8Jxd6cCp5E1twuvq
NwCcpdBTdH8q2I8GLj7HrMpn0zE6+0+5OnhD36Y3TAKSete83bBDVoDhxMXSpAF9Uv7hjidyRr1X
/nghIWoFyvJEGxKG1nT59wIQ5EnsM7cEvFEg6aezYif+DFzLBSHSidkIxrz9c6F0BUA7bBlM8uUP
m4bTASOqjRbIdkcMHm2yuMlmE+pIhPxgEtzUhaNfklOvLjN6Aor3qnyiZHSCFd52oEy4K2yA/g0S
UIwmhMRxcRkx4H+i5QBDTWd5kQqqfKoRcmA9rxoYB7DGqWxfIvZ6eoBNaolL4CGhOYXrfNvbaBue
kLdlo8frh07BwiqjXw2l4fT+AhILAVpU6iB/WtuXNwAW5ED6ehuzPHBUeHpE022pzo906/S3/fiy
Dt1Z6PTqtW0XCv7e1WhTyIaEFqnfkt4ehUH9EtLYffJqMuNhd0ciXHQjIfkRpuZ9W0fh97/OIaoT
ThpjuUQ5FZz0e2glbbvkQbbRb4cFDxlBiLZ9zUdLO5Ay3jN+YwHWfX9b6Uq5QvlpVwwW8/pKnUIu
Ozo4LxH/J1vJj2cqrI4onNVzXYMT8BBl1JKs/X6Fv4g/iui1Z95oMga4vcnyUsiroW6IOLcOmTzy
ci8EDEBju/2nrKQNvuI5yK3ioF7x7TiCXnIOKVy5Fw3EClbzRgZq4IVkhJUX+uyEZyJ8k4pIo2DR
9weEalSvNavWfc4vPEPMOFO0faflEFEhz76cUyrzQudLAuFh6+zEXGV61QeJbTrpMznzR1S6Ftw5
LXIiLacldxvOtppznHCdxByI3aG8FqTQvHWhxhEDzNeMnySJMZ6aiEIlBcVUPcyiLxDqc6CR4GL0
u1NLB5mlkF2dDCvRRvul/sKm8xeECs+6rZPXKtIja6f/uPOw7jaBgp+YKagbzAWdls8mfjIxXJdr
bDRtJQRd8J/y+Vpgaqif1/8FolBE2QlwLPV3MdSrvistU1Cyc4RBatqGAeuKo+enV6pq+R2J8uTl
oAl6K/7kIhQl0tXIzt9ixig/B9u4wTVhPXieXUVusutk9HgIt39uB30LcvgNkLwuj2X/CL+3wW5I
VN4jH4myTu5K/hHB8LXH9PuTAoFNlWPgF1xk7e3NDIMDsk6YyqFrKaLC9VLZk9izHTmWakIa6Tbt
Vhyk68DMwB2R5YfjG2YOm8N1HPgf1aPPdydwqriHalViFJqMqCthBHN8s2BdhKCgG4Y4QARCovVx
9buTwQQgUu33rBip5k2OXB8YIO7J2q9X+mydvWqQHmqbDQv/qxaUGASiT2x3RBOksYF8ixCWGTXH
Eth1ovFWy8A3KJUiI1U7i422cHkJAGF1wirf8h9f0eg0H80VzN4Y+JWBvC3IB8LZv/9VoN51rwhd
AU/7cufT/FizJUJhv+jyUa0JSIKkZ0PJTaOpkeTNIQRDGYcy7IKSuUghQ+UsXrSe708Vne9dNUPV
GUV9H4TghlC1BL7vs4qhlzUDQJfga9mPy/6VhYnDviULG9ZRCZkqdzL8r17IXeYj7VN+A+IN2cC/
TdvS1n9KVoPIPZcnMcNfq0R4edjyrOEcgORejB8ZeXh/nZl+LviUi3zyoWjodTaRwY6eqU59tgQA
Dnv4P78RnoHeEOQk2URl61yUKGcQtb3jHGwzqtxsv1s6rJgYWBaDxMd21cZiKxx1ckwu4SL5tSeA
SAeBSLB82jOGWifYI385QNy4whEIW3Uf4xlqsYtmgfBMOy4hHaZcTmp7z9GqhicX75D5GokY9qwo
SwAEMnWwCRCRWOSN8nYlbQeZcI8023K2B2Y22ShwfMtbbAtBYOn0YE09JZh+8wJM20UPBDEeXozE
b3iNUSF8Jmc/Qv0DNHSHfih7pTSwXCam3m+aQOGBnf1veVc50FxuJHIKsQlwzljeybLqZEbNDsWt
LEALXiwGW09Kre9LDn2pR8R6gqlVmZ4KWSCnITcKKe6YsX+2RSxZinzGVb6jbWuNNRzGrBdqiunH
zHw5mrU5kwjP5vF5Qr/X5iihh+NHFV+i2lAstBc+xvv/8QgcantXdSqyDxnSp5BpAaLaq17g+iga
3r76KFefhGNGL6mo8lqnzoxWVsnK7nGNfre/NRKVWFEQrzuoph74AAorZVEEO5LUu6W30/zBxcIu
AAkOtr1WT9/bqI0jub0kXQ7DHtw1HH130D89NUiYQsodcYb6iEac56i5gsEHuO0ijntp6yHLmG9E
XOV2cwOa3RpUMADoD73u2kvRRWK6YyiBVdR4a82idUtmlXWvnS6L56B0ZqLBNdnUAqBusyyLKn1r
5VjLUgtux8guahJTRVM2COWc+hR+dKYsodNgfVfYcKyNNp7u0LPALNLoLfsAli6SF6YFk4KFu67U
jEqfk4EX7+7RecbtbEhsw0fvrj4QC4YefwcRD4Jdmj0cc7jCYb6IGu6j071reQ0TwzAII6y/BxH1
ms8xyTXM2bRXf5qMqwmb5Sf1c0SlpzeWusUX67/4tFPn6jt5lMeCSCLxERmk+bm96e2YAt27xMb0
6pfrkqA7clBbbiLOQC+GyjDpox2f+hWYij6ojViFxR7Vl96viIEKxPHTkCXGD0g8W23e7zm/i2Tz
iUXqOdxdvJ8uipqJp4x8RYJ+ES6+3F2T9hCOPnPMMA7t4wDOXzD9eKFYvTnd/ACtMwixo5uCwlQt
KP9DxrKOiN8tz5W07Au5yGY8grLhbGdhZwUxkYieP4SCrQn6IUaLd9li4tfHPOLoEro/AAIV5bau
WpcehTnYPAUf4W2qnLOsAhrxUxo5bwCd0t1oNQX7QhhBwNqFnFyJw/JNPugNKbAyAu8/OC7Kxa6a
yflriej5MZgXW7CIF1XUIUNFJlOZ2SPBEOlrGnYaictFSs7stKs/jxQ0VaeXxDD/wwQitwtM8dcG
GdRRorLxF4EeXnmSI6CykivTB9KI709Tmc1GAM6TEfHORRemkkp5mgH+xr/55nyXy8TzFeyXoy8C
n7wE1vIT+KzBsDzS0HAYlnZSs+SY8F4zjsXqrOlYeOOPgW1gju5nE+T2VIwvPJG3z9VjOi/ZQ8vV
W7tOVnmDkc1tVoFCGqsRjK0/dUQTgeypYzn7OZffWRvfTflUYd+Dl6f8u8oRhObNUs3WlThCwa4x
qPPSTmW2wdkXZvLWTKSnHa0dwdulTvF4mgFihs1JJYLUmiX5XagLH1cf4puvgdvibznRKu6Beo6o
oqt512TeHfqilT0jQhsDMuSC1wacrmp1ZDiBtAx54QXQmNkC6cdn0dIxub9UMBefFkC2Z5jBI/hE
msakvhwOX2Xl4W5AFLNwPRgrcZ7lq5f810QyxMWx46KVTTYtrcNG0y0wnKGeFbbuLk6vpz5Sbetk
FMJr8DYfN4h4NRiinJnqoHOgwMlezORt75edCGmPEI/fCRbfbhAws3oeFokuuscwyYiKULuofeNx
Hs+MjjPpsAs12px+jqIywYxCatRXdE9QEcZ0J299vVqKEt3lZCAVbnj+3LvZiWb50Fk4JuDPtFEG
MIxfRhbf8jhX01/pR7ssy87wPdN4NrkWjxARzCbf7Ajyyjyuzb6v2NH6xKlZ3Hl64/sKkJOAwwCu
JmvlgiWF4yOhNXYw37lIDJf/hULbXz4JMhC/fpRkXW8INQTGlanCZTbr2rAdJnqeCv77zVU3T/6m
nkShqaRYSK+5tkYqcy36XzpgsOr+j626IcGXdY7R+piI9JoW3niU6G2FXl2+DIX7u0dOEjAEF1Jv
eLCdrNmp1RT3jf3BMpyhRmI+Ehj5P+Bgq3GmS52cdY2Np9qktcym6lPoG4iSlT5Bu79H10X1YBhR
WNnAzGqg5SBTgDYpQczavjzCE0gSfPVZROGFAsoB3NtrnQ/A/M+FzvE5YG0WtynxofSNOJ6ik3OH
ilLoM/TmyXghg4Z6YlkaEDMShxIHirx3D6O9AfNJDIW0o+10mEeW2Mbm7fX7SvOp5L3I5w1ruhhp
MSRzohDrtERdnGSrd9tbomX2nKDPBgSSJgxkkcme8WjvKyjX+GtYV+O2pC3TPUGTiffUUvOOx+HN
8DIg1iccpe7QVuYxgfT6YCF3AD3zFV4vbiTkdwphBYfO28cIdcrAat4IefncxO/9V9UyM3LyXomO
NGuYMUkIt9iQOtcP7L2KAePvwBwOrRCG+SPrKfUU+lx/1ZRUO2tKl9FrPfzaclB6l3/1JxQUnzRB
QaCRenylMJ6cn7TC0v0vPWnl+COoAKchdajmbEwANgUWU9NZJ/Femd3yBIDptGBntgOBYPvXusg8
KmLDR1rEJZxQZw7vjZqAKengSmxFSfTl0fBS7Z3KM2pdkehHFtRO5lH/VxJTXyZFSZKZuxOKsgjN
Mv1FxlQ7jm94c/MnxgKos+kYAP91+CIyJk97t8FuLyAVT04HACkRBFNyCJz6ptTJcFX5ldET/WYN
7XcYHoon/qlrvbKrpwQcJp37vYWXjZwPguxqwZWsytWhnKYry4PLqVC7kBhrjYfrTykL3H9Wbqe6
S7sLPkY/ZEvHenslgEQDFOyblM6Bg4FLZGR0GiBzRCqumrU56opXtZIN/kmYcwjM5zhlfHFXx6JL
omMaZZNQtSaq/cureR5nM+cGyLe4uUl9A2GkoKo1U6CCMQ0eijrOfA8ZUV8fgq5dU6sdy+1WEbYC
kIYmB+4FamqkbzWNYlgBGfWiP96M+ZGkIp5eZiST54EK17gRl0XSMAJ86vui81Poh9bMny/If09K
nl0flrALUPF7Jy6QYYjIod5mCrXZhGlt7tEiXVckTyIKw/AKKPLtyqXjZcec2A5+r/xpnpYprFrO
7J8tznaVQdx+V7YsXvEkqPHdbE8LYF23Me0uTz6urYf+dh/BHvEWZpF9xae71ujQcdSEycLehcPq
VuU0zlaQ2jKb4aexSR2ISYh42pqpKgRxGUctSX4tJ6hvfCzmJI4RaIc8XB4l+a2vscE6qnb2y0Kh
aDVpciEZfC/FdCtOduOkM3gBjQwLPMxUQglaoBMGaejQX5OpVZTKqbnFGcg19w9FCAtQEptPSoEz
s+U1qtAhdCCMXRtxDj5e9FhVlXVcXexDSjQXbWWrWsJHRDsIL9M8agi/8sMl6suZSdqYmq0u7oXt
IEvB/Js9h9tAmougcgdR6JDQ9ombOUkmr9qyXsCNdhjYzAPF9Kn+6T+OmpVRgble7B/UHrkTzTHg
Isb861jE6rJPlJl5GEGBbDHFiAO8enn2B88Bx/jCr0+PUhullK46tUm3eEt0pIzxxg430F7u26/U
i/UNzSPLQ69u1Os8wj9RoeOdHmhdcPP4xoouB42dtfClo3RB9juwWmV9k2wOMUypi2MGOtT0b6rS
NSXYp0+Okw2HqQfAsfwxi1836vYlWSI85EFZHcVDN1kCSrP1vv3VSSlGaFY+bTggW0qKCxVfwC2X
PxixI7MZ4/YRehrR1hm5Zm/K9t/Zs6JoWcBSFQJDzijNeLkS5dN0k5esbWbV/cS1UmDNVJMwUsnn
2N4pc6icCFQqfaX3al5xPulxxEpS6Rm4TT7S3pJ62Y2ah5pdtvzu22uoEm7UHVO/xXOz7yn0gjFq
zVtCnGJWCqvZ2BOwWKTa3+T1e6KRWfKE42M3fcQAalUwKSM9zXs0tAu9pUvlp4izilfkpifQ7KBg
XxfgopA7Kx2AvkWjScnj9fLYTmb2zA5rT6NrdtbM+8Vpvfesc9O73HsvVb66nF21YSaM9Br4QkiM
SUED2EPGHZ8xEohYSC++WShztWi6T0RJtdV8sAavt0gooTPJOM30eZ50Es7x2BT6aGqGkCn0Cwl+
Mp9RcrW2uy4Z/3QQi5cMoGD+Ofnu9IhcN+XPIXFmsGu6ZtiIM09IP8D+KENAedngG2oaNZ3+Mrlk
WjRdFQQb09EiG8STiDrraTcWD/iIE3vcQZVj/J2H6mylmmQa2qWytGTKuz6GyHPN04SB6vbHsVLB
inFuRX5Ro4VkHeY7iW4oJ1RGZSvE+4RppJmOskOQcRB9QlUWtbcOt+cU8eqKWR8xDCBGdOsQoDtl
a6lgtGt6q36kKiQx2+KpW/4KzQPorcUPnf5HGcG43l+L50lhUia/vyAxO8XRwr+mW1wtagQYmUgO
68OXmwCRxz5pI8DCuIbM+FdUuffNZBChN/PASmVfiYDAHnjDijpsozVjb8AIl4bMqymlswNWAUGX
7gh0J7CUqlhGqJFvRiRqjM3MQaMW2jAgs/aMtkGjQuebHLQP/u/ZfRZH072ydw/CDnGTmRhw3dob
1XT9B4Osyvd7T9LA2CRUCNM6LxJ8eC4WVH02nZaqmwtgmnzSRjq6r2LWXyMZQ7fkZF8kVOAhI4Lc
EzrlVcz0PgF3dsESAHjvT3los0svI2UAwozcbP7Xcw7Vkhu8ybk2mfkXuJZmpMgpzNkZQoW/BfRK
png/xqGH2VFdL+eCoPjmn5S5WPcpmF0Lule7G44bOyRFknkiTEz/fuuMDuz1NVvvpX8D3aGENavY
Dle1HOt0DQYcyPBsDzLmtCIhALM2EWz1mx/xG+2pNZ9Bw2VWS+pu1okiURzttGkk7IOlKxeY5sdc
2JPY0X8ASLK0k1dIacg3Bsqj3kcZDltiC31AJYTdhGGNQpsxfTJZs9i7FSuqSlE9IKu0sjDicoi8
OE0337RVn9RHq1JUk6CHIoI60ylVKpG9xGS5ywwet1BITEbqtF10ZcU1qdKcc6AC8h60NgO85whY
ZGIA5ort7x8GccSWrP5r3vjig8FdEyDkN+yShPP6u3+3hmjoMKLo/5xMdWXXA+xSWru8ubxuVwOc
17TT5Bdn7a2pRTJZfmzQr5EfHXSt/EQC+H+v9sLcwdnHghldyzjxtXb3xB7Sr0FsRx3ql+dyLJsu
1CUe9LuAebRgXRgOrVjZ8ktpPNT9vtGUoUCvAIJJg37vWHuE4jQE4v3wUFlRVhALyJDRHKFnE70z
ERu/r8wV7trto6pkNdT9tIbvwDFz7Xf7igMWJsjGN+MKdAW6AnaiHHAEgIpm/l59KOFnOcWS+6iG
jSyfF76rZ5hGE9o+ItLXxEeIg/mDu29MbYJF4DNpzrEYJdfcLs5UX2Ws/QhnKZuDGqvjulgKMSQj
N+Eq22GEzM2UmdZ68LDk7NnMbhKaLfDb5hRSNi7jSRLeC//IPcnmpnVy3T1yshGuk8bc/OckYloV
9CNIuK6zxqZ5HuMnNw+TwhOAUy78CnNUGaHAVklN92EtOy4dSSygJ/UFd2DdPOdinJP4qK7qHNdh
uvh0n1fr/L8XGPMv7QO566nHpmyQFpbY6VUC86hUvb/zxuByuhZ4LFZztdmrSDrNEcjw5JBzWkyM
9gNqaMVCEHI7f87EqhcmJ5l3Ga8cG2IrFXrlQ6UR91ByriLciuvPl16/EEHNuTEiI848bJs9vPD5
Z/f8viWXgV9Ua8okIj7x9IuOv1dqiTLZ3fIr5DudBpw8IsCovmyD3ba/XURsKFCAKjJ41vOn4GIg
pikqgojGkGA1oZsKV3beGKDoqct7P0h9QyVh0/DMzZqO5nS5+V0QPLCfmuZW9QHNGKeoW0KvGvkZ
nJc9MwJnE+6wv9os3ujD/w+BoDSiHsb1CE2oCEvNJfiyu7Ax6XX7B3LepnoJgJRitU6JIOgrUikd
AzL8RgE5zc7IHeU2BR2T13NZAd2g2IWnkdE2jxoLEYaiLS0+7Fu4rDzeSRF/vapYj6MTVjnZcut9
ulOmx/9d3cfsSa0Yr096ShMeaIR9+YawONTbRiQBbPBuv8E/H0XWjICXLVoNrLNAYPb2r6tzuJE9
ML5ruFWn7h5QLDk497oCiYycr439B/hlQDGMLf/AspFOIIr1sno5nhogclnNb3yfW2adJRnkXlt6
j+OITBpTFOYgdUxy3uhQ7XKb2UvhB0AXN3jfOYhIOXn1fPd+m6i4cFSdix5MJgesfYxEtHItsqUS
x1gXzgdz0VcXOFXN3huzXQbmXM7zCvGo8nFiMddLMNfDX57qgf1J2mlR71wKDkn8gJ214iDlqqZc
tejEGoNDmyiCSRtVDWZIqtIYN5lgI6ToAHbHcctgjwAaM6U3kU9j6mGSTSMoFfhQfDVTTnE03D7N
9c0NVe7vOV+8pybI3Hzlvl0Vb+cabUFhwe4FMF1m11YrT7UimBGnXuPoSVGSI+msnaE6aXjAYVRj
PKGnm/4TEq0QhVFrYaJB/zRFsG61iKsZPWcrjGQlBpBvOeoj7vCl9iC54auukW4sHW8DUHuazGv9
YKiX347+fcGPQ1AIAH1H1ewmmPgMBBSQ7PszV+LvIg9gwYDVCufKem9Mr70sfWsWRWvvDIP1a/V4
g9T3wd+W7Z9pz95153VowCK3UPtv360PQs7XW6/qiYWYGX8umFtAI5n6GmZyIL5Wo5ct4L7R8J/P
DgxitBTNyZwcaAvFNNwchFWY/Rv2dsWyRMoLGXYyGSZqapNTSswKsJwP+XKZ7lYJYXRBVxlbC6Ta
BRhAQDl7KG7j53E60xM976uOGF0LOHkjtBRGux5Oh9HKuudUAuIHtGbNHN3DmTiqeGFGGzpc1nOf
wQ6pCnnAzf6uLbkJMXfK4g0tTOyJUXCXpsjKGCWj903fFlc4uDVmbGyCRViognDFVrzTQrs+S0he
pi0a0y/8LBaPWZVmr4NbEI0vPOBEFyqDSQYJLoDe1KPejTzA2OFAxdtndDeNwy/rte5zCctEQpOa
mYj6HUNCpHepQXT9LQwcw2AkJlQC5ywEgZ7yJQYbKK6cnpyAKWSSmFNQAITWiCOSxQyhiVeRe9Y9
mff+rB0Kf+MiXTXyHZoyOxUaVKfVrCXJlZLhmER6XBSBrv0O1B8nDVzHU5vZ800YqiZfADibOEqe
N6YA3/PwEYKYgOar20GoBbWh7jF0quKV6u15B4vK+DJQLjiBmDVPEa7aJxrroP7gt/o+UaYdsU2l
hETPkgkYLsHvepeP43RUjXJLJ/NSjE0Rg5jhQ6kCzOR57vFjF16UMyWFOogE4amnW/QghoMPmoux
a1aOlLF8dPsfil3E3PPtwDd6FM8f99wkupXTZ7jiCUIXwSew3AmcAHn30lTfzDyriM6GZnWVPWSp
pA6yFladXvzXmXgmPlAc7Y/auw5EVCDLT3KOXbcf/GKRdP/BpGDJlO8b6rjmM652x2hIsSQWaSjQ
ZhqLkAU/rtDEU6HmsJocXgcKjmTPmHf7Ppm19GaL0lJHfYzdOjO+qwFjBDlpEP0qaDoH5Yxl9hBs
UqR3Vmjb7OC6EhFtcg073yeZbEk8xQp0qDPAW7nv2cn1fC5KHPBEAGt0SI8cXcCoc3hXxwbs8VSQ
5uw7DlEPhIxTzGF5vTWvggcPEJHuosKo9+CsVe58NGvUVS2QBeZB14f6H1UZxYja9PN4gQ2otJ8l
bulynT0ilgWIxHdbhUf9pIADoPI3LXcbiwiAfS913mu7o03LZ6GYgakB3X2L2hFLxqLiYf+VVoe5
zSIfSOC9MIS5n9F/A0hNTPxAYaVPwta+qkzIuqHJw0Ca7ePFvx6b4AY5mwWEEI06DCF9+IiSKtE2
kMJhSdn7N1VZ2soAb0FSDxZH7zMR+qV8gMtx2xK+XLQKKdIVhcWQKu1FrXDTTrGojlsIaBVw2kql
0d1bl2QYiKE13tuX51BeObN7mLjR5q/vY/flIs7mnPowlmJbTMTlyja7mLq6c1oX3qZ8lmW4VNz1
aDWGl7DXSc/DhtBMsYq+QX2+kJhGxwdDUdKOXW2dVhNDSMIKMRcGMEwRwUObd0SeK+FN6UppYz+G
fGdBaG5KD58g51ZMTDhXXd2hlJYXx4YfoQepuC2MT+0+f8+KgJ///giiMepiUeU70Athg+FDivIc
SGiUc08RvUymacrXBWIznw80X8e6Bqppwb3T1EfVYs0lmF5Ww+ZlTkZwI8UURJgK+yTA/oJ8ym8X
vI1xuFEbzInP0/TefmiviZ2QK1ikltJgO8lcNyeSIFyAiTkIPEiWAg8/cpNUKYL9s+MCl5k5GmZi
Ps9fxrHN5O51TM3Uzecb3bgBEGinlQOrsH9FqxwdhaPwJtFM0xM/Gp9015PlMQ0sZ270khfvQfCv
J9641n2l2wD7PrrMgnQHps1+/+n/TDqvlbqjXs4zghAV6ORKoyLdHaRAHaSHG2PCIfw2wdb63MfJ
MI4aijQDugEAph5Nhiowu6O3GwQTvW5Lm9JrA99iJfd52BgrhHAVsXqT9nFPiGPJAavnCeCqHOfi
wD1eV+dVdm9RJSwZfym5q/e7tQGmsn6orB708MQcgJIzS/wfmQKl0vhVA1o8u8rWVPpz307UTSs3
uK4MDo9/kpy7Zd2AUvNGgsRP0VGGyP8EQf3CjXwo5gFj3vK19V4C8J2yIg1kBdYUx60yg8FRFFta
n/8hv03dJ28sVq1njPDy80W4/1NzzRvKdMyyS55eGQSmoS9TdYlNQ3XcWXQR9yAG1P/6z0dYkskw
TZ9Y6Q/7kwuZcXt/SP66u3RqZO7dlTE1wbZlDcfzZ6LADOMA68akpjv2B+JGOrJV3UnsIxsU/IJr
wUIWg3+WVEyDO7hB+vO88sroTy6ZsmlwUQryJqnrnvnKmbUZ0dGZQRvWrkNrC3ZJJBneMb/I2Phi
jTtkM746UWJbnmVG250rNapZYIqw+eOzvshvKFVVxHNXaBzUOcMo+zh7Tj8dF6HPxVsN6k5ESsVr
MVLykdm30DMFeuDhO0QgpIxQ703SNXUUqWO1M3zPmFvvonX/Tu62vTjdYkWjEGBQ9ORRO0hi625D
xhWLNcGAuFsEG5m708sOAsp+BFNWyRGDDulYIemtIYtv+2B2iPG/JzHaXEHUSMdAb8Yhs/SZVDvr
Si3T8DRkYhdsR58Yqm+m8FAJRgBY6W4HJngnfgkl0P1e9oz/m/s8l6AOFyDTqY0lQc0dpZUlPCfG
w+SV93R8XcOPYYhogERJiGAqcJkmz58D2x8NBzgdFEhQwXvQNk/H5hKOlO4Je0IK4piU5+9D8ESu
RWU6xppzRIA6E8qItsGQ72tuiBeKhv2Xm3Y9/giqsP2IcCGmCIwu7N8bRi+v8JqlW6wtRb6LNJnM
Ta0yYb0Lx3hFLm4TSmxXnBZz9g4tbAwXGDcoppVXbNgQzwyFT4iIOxDeb3D7LdcOHVFwI77ThPue
IAJNf1u+wcEk7D2HSg+gO6+LrErIEiW4P/ssSqseOVk7H/7ATVb41zlnzaZS9GexM6vawBF4Lnra
Zgw+syHZkJm2ELJEXF4PlHE0LnKfLEqQU5GKIPiTE0Y1jNJ0VXfpxY0dlLoDm4ABU2+9iLLdhaV0
GRwBuCyBeR1BRfLIwN92tBpllFED9kRTsZNz2i9Tpb4RSzjJ/wz4HneOEMb8lZccNb3rfEqv2e1q
fCY3EZY9q84HLtNXhvRiyMwpSiA2U7W1TO93Gw301RJPIUXH036vTQxff0T9dzPE3kA9zOnrymfF
S1m+43drRbSAJljmZM4XjqhftdO0h6B4uI/YvTaubUwgw2dzXz83NHZIJ5I4fZcAufJZrbBDPT6o
BXXdF924dTC8keAh0WD2QixEjDo0Ta+bjCIrc1LEyo6k9ewh2av8A28k4plEwCao/4NTV8C+2mga
AVxKZeeYmyP48kti1fmyo2NtqpNuhOMjgQqfz+sSLwV38AjpJ2KgzKWUei4+DJ9K0xjieSHOxSzu
TVM9aTS5/WI50Ds8iN2GId9QRPdSDMSPfmdjdRL/Ov+7/TaBPZB2HsYJ5y9sHMsS6tPhcpnapDpj
T8eUQYOCkZ68u7MR76rYqvedLuz4y/XVXztPmOUNjCirIHXYj/FDyq0R7cEFde1pDmaiM+dl98wT
/yIKbemdZR+aThHWLYDvj+jwPul+WgqRLyBBLieI2MKkGHkOndrhtowcC39oEmg192W96N6DVZ24
efj4S+NvdrlPpd4ibREftmrrTdd/dHHIx5lIGCpWqCpEdh+XiLSJ+7rIvZeRg3KS+nHrYAjneejh
s4wb7l5qj4tYBUht9++T5HPdGHdIoAIl7ehEPgXgo8i6asACdmq2tQCz/IqpIzAjiCeN0m1rx+lB
r+11k9BlCxe0+qhyhctKhKqxtYUyMpJY041pzpVl79qW/o+x+oehqQXDjxwHpz/7Yj3rCYDNnAId
ggEAXOyKRXlfyTkOAGePLsZUQPyi7TGg2du31tbz6nSKj07abHXUc9/tKaX3kkcmB26ZArmc5AuV
73705eHovexGGtbPXE8RzUCfq1DpdC+mVuhWRzpLd4CIQXeeW7lU53Ib4M+ptiqtCTM5Cm1FOw/a
CplZ4cQLYOI7utQ6xnXKudfPd9DNJzdVCsQv+u5lkH2/mgRNIc9wBdGq9mEZhyR8AZn4xNqRuaTp
+JGx1ApLw5WYqUHnqFSRxBpXULKcCauXL/ODtVrVRFk7NfzYHAY2bXKhbmh5BnfNS3PdPYDuEq+P
8YfwDk4ecMNYfxQG2BoiqA6Dkbks4lYNIT5Bhcz8fgaIXPDqDe96a0QsDtbaC8JbG+TrNwOK9Hz0
4TN/WIOe4RtRAdp2T99UQekg6On7q1KNqHLgf29CWNhjxLDetEaZcVnRFBkM852UiM2ZQI19Sa2D
mIHT34+87bfVsiWmgIYEPpBTD0MtI0f51BsbbdNbJrMkq3TEkdyqK1Dq6mvOdE6WbqzFF+rde8f+
S+KTVKsx8Rw4oXmrdCjHuf7R7QbtKdQhqY9ghjJLiGM/OCecTFalHDI3cTgob9HV87HLljidJN94
HmMUoudIdCmhHeHHMKbUOa0fQ4+ljnU87YPHbk4VttPO7DqZqlIQOL+KO+Z2VLUcOCvW4dyFuCqB
JpYiTZuCVuQNh5v9kk+23KfN5PKRPxWtEimtcv0eBk61AMRpHrhvbU6bafCLL36MItNjGtgnulFI
2I7V2/8OIZyE8DzVzKz0pj/eULie5jpDcMS84YN71X2uKLkz7lg2Huy7hIbO3ympFGjsk+8nK9WV
CQ3yrU6gqtmdR9LvQgm5HlfBX4M0tNq20Qp+ou2uTJMoCAbh8cfSfDSOf6xZxyimJejGftRJjwK+
NNRqmQ/N0hGuuey+BKMr7QioVQAj49xGbJcFkUzJzhh6tkk+ZaCswc6+qZSWp2WifZ8Ya168LoQs
S/kKHL+I4tX/EDoELoqazDPOufz1f/CTOIzOsdDygpwI7P3/6DGhtXuLM3KaYnt3Z0Aqjvu0Nfj8
thiw+Yr6h6+HwchJwROxtRlqn4og5lHIauvWVEvGy1mEl2NS5cvuTBNaqsewN810XSsQ4MzYIs8s
7v4zoeFGAuW4kJUfo1Yl90sth285RhvlcnNCrYWH7giRMDFjiuCAooXPg+sSfaBXTBzINxfBoONi
VdJsj6n65Ilx6L2FDiLQAHGDj+muMQfIhN1SXGFId74xuD32i10DEhyYLhyS8bQ5qXNohs04NxXP
43Dk3+LE047rtxTK27fAaw6sp9LGSQber/e/ETcJ3YmREqEMY/0b2kfE8fTnvq3ncXTAuP60T7LN
fBMNBN3a5l6d7ypfQVF7xsEikxlIoKCZF3j+tw7SiOELnHdlorPUh3eFEVPGbzst9z5NqQzmvNDh
wzUf+j8pI9CSyQnSNicR10S9SEZ8FtwT6TBX9FomtYFyx6ZYImAR2nvvta7mQOYRRsUhnX02evo8
nx4Y9XXmf4x/2dOlqWbz3T5+CJ9bQu0dM8sWH1KIH++RCpIZY+C3d2Qe+Ty4x6G7N4UV+lDb37a3
qOUPnKZtqzNbb5SXx8V7iALYSjtK1dLhQtSbjdZdwJjxGKl/euYGwjlg09OytmenEMV+AThYCEuk
5VicT/XeS3H0bOVnrncPOP0mT9CMXgRF+VPJcesqLNQRJaRWwarZ37PUeunGMAdP8f2P+fvpODXP
7W8j5uZfo1ZbkW5STjQgF9fCHrI0qRONSpA2/u9sm1R9xiez3YfoLdMnnfkhIbeiGZ4xuN4Mvd2R
Krt79q4zitvsfGC4W6J8TAM9+d0E73tFSRDNekdxMSCnRL7R7rJiAvoJ6NwXIQroB+XKFyO8yxDo
x0Yf4Gq0Wwj43P3AaHaxYhOu9WuOrxFlXLvfIH1MmIYJfFIQDZiMydULd6vX4QR1Eynv7JMIX4Q9
YQq0LJX30ZfgzUY3ekxRHP9yiHTugmdbLOyL7+8S+JYUUjJZeJgzdjnRYbjdoLUq9x+epoLuOZ9i
area/jZUWpLmRP25eoYg2gpbD8SEfz+zuml5716ld1KW7Y9BzRYLZN2kksMXtKthobcWGjOI4a/3
OdpINfgZ0pVKN3syodazCP9AYDCBLZfb6olCXjiMCgxJSzDu/zWo7rgnSnfrWrI/tvgC1pbjYGz9
iqRdqN5rFv1AMm16nEdY9WeIKFtKnwXBjhjeGd4YEkzDHd+YvWYDPO3/5D/rYuOzhZJBeIc6QCmf
2KJ9Tpo2Rsp29zvqposmiZzxdmxV11ac3/qesgZUmchBC1xnepOdDbc8fbSd4Zla9x4pELrUrYND
JpgcA0t9RlGLb+BI1+Wt/9JC37HiCraJ96wUsYtwqJDvozwGIH8cle5zSQNcPFRBrsZ2aBcWIDZ0
zoyAuWZ1ir4EQk4CBZFblwvLmTQHGW1h4QhMOXxSH23ghIwBy8wI/tFA7aVEdb+Fhk7ES6P3KOMP
m/4HpTECDABBhO0f2ZQOZA63YWU8QCBqS+igJUVNL+4GLzxMhcYM/as0ginxAFcNpaLDwIkD0fmH
4JTHKaFhb6dQ1Jh/qfiK1YUajqO2/5I5atfddVqI+06RX3BCeLR1FeXoIUq+nTN4sfLqIyDeuIHW
f5NsJs4SU2U42iOmcajJ84vyhIFcVFv+fRdOUMyJzQYkXhTnVmofWOMeTm8wlTkzoaQ6EiTbz1Nr
Y4GX/Wb/yz8fjQaNaw2aseVYppYqaH1VrIjnzPMP0PciF/0N+4l88C28J86kxVOsmeioazZe3N1R
WJszZ0JUZxoL3L8DoocWtqNYQLlkRQSiI6uz8N1VEcDZkmg4yzCjKkZKTSxbCSvUIRw0V5P+eLUn
CdTs8LKe3Ugs9KsxlsqbEPC7XbUvwTTZ0UgFC9YA+nl41eAdMMmsKuwaChBIQMyXFyhWeFaH34lR
xChV277M47HN6/Dochbj7/3CDaFzNnwv21+f1zyQSutlwuqeyOBpfAhyKawzKBbq0SKHLERTmrw1
YTigVoHlNxBSD/3VzX1QZLB2RpI8SKoxbqdCxzE/7q5KrDJ/2phZgyDP9E51S+fA5zClrxMeHRai
g8KHpvN03rKVYOVC8Y02/26uxjPNoPV665zPlmH/iM4BxeaE2iAqae9SG7sM0L6r8Jhl2ZREUsAV
WSTSb//ZS2MI/evYaEHGyYK4L2BM3whHPBtlTnKplXdsdS/ax7QHyj9JNVC9OYi4vySbNJfuJqcu
mBIkIAU8iSsp34nt9HCrWipNvu0UIWBeeRoXGS++49zWuJrBhma/lDeiDUwr7H+LsNegywt7MhH6
GSVubFdN6jrp6aZ6HZPKWFpX2H1sxe7k6nsZZwLiltmipanZmRUuFhe6UhABPqYGx9P+TkHZoDKL
soAA82MN0yK7Yy8wFHppnjnmf0tKjrnf/X8avwAmugwKqdVHKNujoROpqs1IZ6cNSqNrGp4V5eK6
6Ykh1WV0Rr97QPPbLPPo6GQWoOmCvulOA8fEgncMMcZC+7OMJyLkFuwqH28IkvHl4myefgkmfXWO
2V6A77cThqD5yh3wr2AaaCCw319ch9D58f+9PRCyE1oov52zhaMJ4Z7eIXL4wzG2M2P00578G1tv
+urE/KdVAxFi0N5iAK2i1bM2suNf6jlygkGMfhFrJbT4SDxL0ooh+g4pit/+0/Zc/+wB1E+xwM7f
N+wvf07x5rdCi2s+7+Na/+AO1MJj6QR9DVdNF1WdRs6+nYriDNoemR3FCUtE9H5ZkEYjnegKExR1
Z/+EV4s6NvL4qfwtWqyYRQcgECjl4lxstkQZruBOJ4AuXrYTuzmgbIOir3EbeNJaF8PZKE4otBQT
ZDa2ONUwS91o6PU6fnhZyrirOSYPIqB/9sWQfaclF/78+xAd4fREbnVYi/sISkadkQE2/OqGq114
RINpgT594e8bWo90jloofqrIb1KR5FddNKidEiE2UHXLZWQvrx31BlcBo6v4qg8dnVG8vBIJV5Jl
1yZc+tRERi8gQSSSNR9/8TTrpGovXV4fS5ow7Uegg2PxVpdLZewBQmB0s7cuahZTcdTuj4RtVOpt
Y+rDK7A9v6Et19s5RAnQXDXSrNzZSoitV57V+LqJeuMI5CrvzbZ2qRDrEVGbVj2Ut50Dmg063SZ7
EqqTVZBZKx3rK6yvZzVG7PNsyAOr2XPPL8qfOF7yC7pVSAqNvS4LBOjPfHsNMHgNwxPIEHC8D+KN
/9k0hT70OF4PQE3EwEHfebUozFahVr490lWXUTu95QS0/ugxe4/WVa6vfV8nyJAsFc/L7yJ5PqBq
ybrCLyL7oXRDv3qed+knG+Yt8/Wg55SBN6yoiRGIz3vPo3BwchpKlTFv9yeKfpJw05xdXxEWWxcq
u3sITZARIuDULsWEKKj6xAAjgsajtsg8lwos5ZevKnc8ILe1XgxS6f3xz1pjQPD+2J/JW8hBd8bF
q2EIAuLPzXHKjKHzR7QGYjLmfo7QuSEUA7CtShqEyVkV30t2KxvdU5+83lQpg7K4sWyGuJiKZ0jK
i8m3Ws5m1PGzD1DqiYRVeQVLkPpTdJXM3CTpQcgQTace4l3FH3LSOpAhYo5gLnTlWSyPG4PukTay
cDvNCdocoq7dr+owLqdR/pAgXF0smetxV/pfp5YdUMnO1AdoJg9BC6vneoii+pe+UXUc/vO6Ahue
lVVVLoANu0yCgAjF7ScjegmVjLrxN7M3CGKUQENfJ2J0FitQFz/NDBJ0GFCqm6Ow03Y05ghc0KfY
j8XwxP6b6NMZXNq6kjP7FsSSzlV5osb8g2iyGMS6ecow7EpDtUiFPy26OQtGQxCHoHHTIGc8BWIP
hBtIc9AzzHyGSsnJwtWo3Q0EeuTpxWj41fd0PF3EpmgAbgut0Gm9ShKgA7OtdVaTMXA1XDNw4riT
S8apIAEmQZYLQe4GR/4W5+2CoVOC3LT9WMqxbg35cMywrZUFOK8ymNoq8dvGyq2YLWxS10cxHstX
YwEycCy37jbn4xdDvB/pkyWvUVhW02kHVJOQoCNQ2P+Otrn5NA73e3UMf0360pw64ZDYSM3jC8c4
kD7nok0JZhuLxYeQDrSVtfUT7r0ZWIDMF8DN6v990Fd4GlWKiVdOcz5DE+YSCInGptEDC6TJJ1cM
ZRdGgiiV1CMT1vJxWxTaQuYfd92+MCiyFpdO5G8fBuZOScGa94BY0UqNUhYOGb/wQV6rBz+ILjf4
t1XvzeXMoS8f6qsaFeUUrrVLsM+jD9Ikw8nfwIYYyOy28prHcccNej2z9DdHZ6N3W4DYCTe7GsyS
FDzeeTWLwjSUfAMo1oaDEfJRcTfjFFHmXcJSIgQUYaQzXF/GFqoSO+GFR6+YsCJK1BE75GzVMUGX
m5viKN/A0fwjOkE8Q2/RfUbhJGoX+e4snt2h1m2gLvnbAeZ7BG9VmhpoYEsOY8XBaESGj8fTrVyW
jIkEZP2q6Fe22FOpZp5tTQ4sRPqkOK71idVg+Dade0tW8/Sp4+VF/MTcCSnMVPtzKfGNMdWdhvm9
VZFhDbLtLzOKBdJMrKcG6qM7njZkm8bLAc2LIgYrktLSwzUq0K6ItMRWiIhicUyrnUL9DTwqbGcm
lfdiJjChp88LW+BsK/ZckXI2mywhP6jyMcvRuvErGBzLoYwdu1CD6c/ttWAi0vz5ohf9iuXhSkIL
SQSSiqvbOGg4q5d8nEPnC/3+b/4x+J3PsxVEhZXpDi8yOMHucHQiT8kZDXzxGNIUuUHyi2Sb+W+k
hRByOlRUqTsMqF8YZv8/Axg0cmR3/daIe/xHZiPBWz/UItCdGKHzJVmar4MHYOWqsPUDlO0rvwH8
JKcluTduRXzkpLMrTF/fyEgrBWTnPbp4qMsKa5FKmlUtkrGr7g70Vwu0Mf5LM0WSNM6Z+XHTxyQB
hGoOSRV6zn5AmHVbAwy+QUDcqkR2aYomx61W5ivBSDMr1pLkqXzkyMXFzaThoylcR8z6ApOVAhwr
9AVBSjqd8/YCNyNTK+MOvt8pgdXi0zg67RbXMTQtm3iU3/5eBhpbWzwv4EVeJTaMGUkOkuzBOPXH
TFJjPtZhA08BO0962f6k0v6LmYKGh/PwjyUsuZhwHkKlvadapB7kXsz08fhPkQWdmfeE8U3pIPjh
mIMoQfvov4wP/SnY/6zLueR59DAd0tb9qonScxfmTHsGE3pEYUYRP/iG9usUlfeJNIw86C+xOrrJ
lrLH3Gqt1UOu/AGsDtF9LH3CH53Z9VtCy5lkhgtaZe3LXiME14MdW0Hx5UQ1BG4uIg9bh1Nx60w4
yzbm6ey5rQGQadFun/gqFh4hnfhyyolD7TRq11xGK3FVXB+aS5iTCI3db/cbUzdAAIBbK097RJ25
9S282QBVJ8vS0PweuZWT9L6T8dMtBXSu7rvPzOUwIBmPuOOwR9Kt1N7jhx7hO1l1/Z+ODoUXnndS
rGY8vE54O4o6ZDbsZEhMQ7NznAUuPjHozysCFu1W02W3fG/J0atcaCV6DBAuj8npl5HeMUHKL1eT
Ix5q8AomRgyChzkyvqzNNPFlX47tpCxeVGDnmdAx6KW3UuCxKYAyBIN7MXoiY+X/704eZjRwDRCE
go9+s4IcFanP9OLoVVNTKGF7DER3E6INxEHNMQ3Alb2+TQfveW55pQPixfNKIYL40G2xTDL2kcRP
Cfl+9T8OT+f+alZRdfFjSkblJA3h3DDR8nSSe3VGwn/7/lv9dX4b9BCHJPBeF4h9QXV0CS0yZ1BQ
PWwvpfxB4fJvxz3zkjJTiuRLgg3pJIsN/8zWKYXtGf9gMahx3ctP7yHZ+QqjoumOlRL/64wb2Cz0
3oUKY/jle2ZPgJftKrcxefZgYJmsSw3mudHG4OeX4/H1+O4zoOF57q4p7/cjvrb1XcZ4824AVrIj
/Gedm0hcn8pDkOwvj1nw9pFPsyIjd6boFzpa+hq/jqIpfD+2yfSvFqq3XbT+fdixQZ8eEZ2eHETp
Ls3dDTZECZQE/EfYPOLNCcnUKdvBGK31q3RflJtkHO2VAcmL+rnYYoe9Xr2wqxLLblUwyweaaklk
MTd88VHhG+TQOzNpTmRhufSRtpjbWjwB0DoVLld87g1f0+X/2EH+9uyXHaRbUrw7nY03uW4FEvsV
W9uQ/rFfSEBaP/PpVSCEB9ltqFpWVOkDPljyskDHl2slJUfslv1Y1NHMF6yRNtTKXB7bMBWf4sVG
tU8/axrYA0I0v7nRGHyD5o3noQ7CdKDS0kMBchF+mA8uWp3D+zjJEdftIKVyspB+EpAhy7ieIeDP
pzEwKUUc/YDLtQndzSzWhlREG/vurJjSUdJ3i3iU4IyqSsWbTwGmuJ5zjrhPjE7tEmzO2zUJ6qAZ
oxfvn/ZWwkSGTa4oAgPVv6kFkqDSxDK1lf5jcRDuCZZwX+J3azH72IHDBlgrDNYCR9qXdHRjYLIj
t1LtirAnfka3dIf17mBlDjNB3gGcR8J/MGoLlGllnOIMKkCOX9VOqX+llcB9mh8kNpIQF/WYMxWs
CEYLOR+kW6skyidP71njXQRQZAjfmAbplYBpX3cyeWsXdMQFEhLngsjPrADyXMf0FqyJpKBIg8L1
WEIvKEzoyCKkYmQLZ/3R93vSL8qGfBBZY9aKMYEpxzKXSXGnmtuKM06wLm5/79RCK4uC/TP2llKc
Dj+SIM3BvnMFIJg9lCZXEOyeKg3h0nVzqtiHumK1lKdHZFn95J48qxlBkCy04JW3fV0lQxh0E8tF
oomzBpXQKFvrHpt72AWH/6un7yLQklvgOobRZr59dr7b2P0fMwO5A7P8UAnHTmp79YYJw7kYClyN
A3H/Y1WewbGLXXfkwaDTbyZJ1G48SwgNonoR9Gyqxmn5Z66bdN+5ms/19UTEMdn3o72jm8+qEWTJ
1UHc0UIjpMdQbVvZEPDCi+PsPcK2afnR89vbZMFcLsw44LJv2koEmnCk55F22jWmE4MIiOROfgp+
VJ8VVgiO6LTNPeWxGaqHhP4nHSdUUNQ+MFq5oW/sWopsZWVG2UqN58Oo4Va59Ef+jwBHsjSF0DU3
6OzYFhDRPAOLNsrv03UwHCLQbnF6kUcP+9wENjFXdmgQMYxP0axWLm2RrgAEmOOX+Q24/lGZeCsR
OmCTkOYhN19it+kQkp9eIYOQee9YTB7Sgz3/7HLC3dFLrpv/o7Fceck6FgLA5LSi/9DkRdtLT2DX
ZlSmK4WLYsuS7YmVRDGGdpjYebN1nx51OVHxprWNnvsqi6EF03O2jx8SBHyQAGJm99iZUkOTPCcu
s9dVDT4alB1FVRN1437bbb1r7hSlIyNMYxe6iU6pYuVfUEsZZ8Q+f/mlaGrsyrb8CDHXk96xD1Nt
0LknjPaOrzMIgLMhN6nLxN+Aq/y9kB34buEsWD/Wqy5Mq76L5lOobmdjBARi0579OWq1Z5MK6HIJ
1C09TfeynBYy1tw8zdFGKX0ypwlW+GV0DdrssrSEXhkoix2/mif/3Xu4hXFfE4TJhAhreFpYn13Q
Q3KJ5/OzD5Dmt6nbzI2zmwQdFX/ch9MZUG89fYY9KQd4WgegVEqv+p35XJsnxlcutsa7c9D291CB
XnOVbjmKi9bmankardSncRP1vu+Tah5QPmlGAL3oNtNHhzMRfuAwavXao9XnCIM3sYc7ca1V3afH
3zxhCDsgYv/+SXLbOJKT15wvq07ev3UUwJEuzVC08HuBxdz+dlEaJGw/jLkaaVXRz2mbmYmvMciV
syMCdkYdUL4EaZCmBJljnpLGW4o7pi+WgmoUXuIhfHvRXareEYHT71NQNpQmvIfFqUmJR8CewHRA
rdX+5d8/16tuvi602303y7WG4t1PhIMXI3+kZIOkDq4G/tZoGY6YhPoP7gIpsoE0yPcs5YfUfQw7
PsJoY/+vqrM9ZhDdkfWqykQP2OHRkJsUyqOmP8EnIIYFurkmdS5fnWFg0vc6LULmvwYwPHXtrZZE
KItc+Pkzhp+Wmkz25QypefSUb01ddHg28nyKAPBxROvQH5dmB4/8YSof8+S3tI98RVslPk56AJc9
d3BCY2GkBhRQQ7Kk6EpzD5pDcVmNNrow0NvEg7hk7kzjr4QTQ6emfSlx/B+KhqnUx/rmC/GOfEWn
GBthUDdfrfqADUOpWN44bNW6GTC1LIlPrhJmHbSeDBNh3Au62Y5XxafYad9IT+meZH8g7e64E8SG
dsGM8U/wURDO0wqA6GBQFlKh2QQ5G+k0EigQb9s2YwBJBhcoZJxwBuA2ueS168NMkbePfMMArmqH
kgCc7yUYDsYMsia6IT1eIEQv6d0JKmoCPdrDPHvzl5sk70K54BdEmrL8biQGJMFbvGuI3VEBje8R
ciPjoMbXXyCByBvqJwz5DKQQSj117cUb1A9Hn9Y7/J/De8zOmIMo1EmdWOEKTUHkpBXufrBBm/J3
9Ww7zPVIF6H9Se19gXWYWhSGSzJKKQ3WceZOPBLAuPO4sjX82IAAor6KgGNUUpTuPPJotmWkzsoi
Tb8BMQ4/lzuaBpvJmkyBKX5wfExB6BralvsUF/pXfB5LobTupu9MyZRkVudYBvCDROwqyuFmlDvg
uwbP1X+wfzuCkVyqrMiUmtF81QAHJ2rr36oihoiZ0e8qc8AtE/v+wWbEpGsnhBORrzjU1vXqeZcs
iGM5LI3035QHMm6yORotMy8sYszsfMaoez+zimpicecEKEi2lSHdi3xcDPOYV7zU6BLOlrWLU7FO
nL32+A0h3k7LHEPokwlj4dr2H58ThI81X3LpqdlexamwSqK1lG+Oj8Mf4Uyl7iVcwC9ZKv4y9wy6
S8hJ8vpewprslOEdqEQaSHQeo2i5n3aCtYn2VhQ5Sgqt3XE1HwSi5uVincCM77jodc71ak0XyLLM
zshVrBik1asqMgIfdpJni1xvlHYON8pr0BDI4YajHDntnfeEQjjkL4zZvnbZUvLMUpj1sjAlN5Ah
aDgM2H+aG7yhE50xjqkFvMA697NRjKj0AI+DYVYhSNj6z06jhWM1etC0h90g2mI80PAODMgyEagX
rJ3paq9svqY5m/Z6v+lTNl1XcZF4WxdUZWOAq8HnPWF8tHJkrcjkR7EXegXfGHVE8LgldaD3zcy6
dd6QC9NPsKzxCpsa+YscmqmBmOss9aZC+icyIpUWcnW6Gr4eLdBkwaDe86J8IUSNWCrRf/VAhU4V
LQYtk+sApLMZEPLmA2tookym7mq7bQTU/ex2i+G7223Q0ZT7UzxjNgww0MoXSK3cmpsBUPXGItyV
smAuDY8vy3hsTpc4HJCQrGhcg4VY7WcYjluNlXrfp2OsLwvAVDr5rU5S/nTyqsW3AkephWFlDAZ2
SbMxtUfggnhtTCM062sCbHba43VA8DncsMMgoZrDDdIS9mfvFB3SkvxstYbhcBO9SDc8aTR9GFcN
fXD4On7gebIihEfLZrwOf34iwJOd1JJa+/e4nsNfQ8+sUYfyOnYGDDlSOYUH6AUpjcjJ4m9v6WAj
XvNjEwqSmIStBcss4/5YVwFzXBfEiTKl3szHb55w5QYM27srtkHQrFJqdZj2E0SpfkFVV3K5VAaA
+8kOx1HnuS0cWOUk4Kqjex59Et/1ouoYl9KXwSwHuSLLBxW+6evSj+yd79U7C5kbttCo3BCzE3K2
3gwSJbEUVWpBqOEzWsXiieHR8VvzxTUdWpspMZDTMVXaxHeuCHsMjYGQWL8VpDaSGP9m6kjwsQGF
UebGCcvFxYmWyAok2E5zfK2dwiNQQkqFnvojMfcPvtmyEH75JN/RACJ5vCPL7sW150w2QBmyi7A1
pXV+B12h2qH7VZoECizgMTr6vrR3HJlzK13BlXRHld412W0iE2djj8D4Zrep0z9tbMQ6KnOn0dgb
WtsV2d3IbWUhDFCxUZvVnOkNlUpj9/mRw7gP24ptWrEbrKsyyPCwB5YUKiWAv1v7fefHdbW9KOEZ
ShpyB+1G4JfL9s9XhRlXUttFwutqknseBjeYInyqioNtvTFzV766WGcxvmMR5wEDTu+riskOhH4f
IyokHM5lDldQwis7pJYD460nBihFTH6QFZAkYkbKJhoy2q/ZqYshSv8rviCW6gRP+87idUhgU7fG
mTD/tw7B3scKma2TK8gK4EP9tZW3TkinHdcyB4udU8CuwD9PKBqQpe5J9TkjsObqbXtrwW6Wf/rX
IXalWlW0KDliR2OLHtX0CumPCsLnugFyvJQ2twmIrOFMhUh33ounu4nerK11POfvIaz6h5hN5TjP
46arOAbu+TeFTYQKc/Vh0vwOnsDGTpgYe6zkp/avSKutIYehm2CmJsKZpljBcoDD2kwlBnaCD4iu
PwUB9hf6PLc8kfVj5zOw6rEXbMxdK3Ane2QBMahjB1ZAjbH8sAQieo8U+/PHTUB6h8EFFrKHARae
AhIi6k/Gt+c4ddkG6u9G4BLo7j50Zr83zP+5blORn8PzsJX2UoO72uzDahiGsB94vfWgi8GFu9gu
86N1XLCSvVkRtnZPf/EBDPpCOfcpWHteYMwyZddpv4M74BNFkAq2xtN6i7sQrln6+y76CgtcWVSH
c+RzzKo2e/ti8A80yBaRcBj8heu+ZVSitcaI2vjM2UFENNxxrLFIWrklkTbp2FGaJ5xFnUqkluq3
bGv4Nx/zWhn2+4/aziWr8+C3wf3GX8z92pTV5zOxzJITeWb9/rq+iB4iNE0Nc2AvvD9sfRPci+ZD
rt7UvC41kE0BcM3plWCTkkrT3l0ogjerTEqlBRiwBUZlFldiMCS/nT003GLI0Y0yEpt6C/4FKC6K
Ri8eAn0lvICQn7zruXW+Xx3MLh0pxXVW/DXJN+GHhyH4ONJQ16O19iWF/JxFPDVMcUJIVkdmhbtg
KoY9UYUDSaFZ5fxxMq2XZ6TgeywM+XsWgnBjDdMnRVr7LjOY851AmvjRoFN8SYOGa2+/wWdb8dPJ
JfxXzF8qoXyvFNTWEo6sEdSOSQ6bkI/i4UoAS+8qUp0sPQ2YsosVc1BT+058tfuV3rNFNDZBCf9P
O9dpw0lCguFhjFhQVAEDgtSUAqgtU3pjBvP7bU3Sni07ecfQXfeAbqyu3y68IVvRArowgZEgvVsL
6YqVkvfydDkVFB+SjkGqBkpS2kXf5DK/JlfzKFFNu5RM+8SLxdbrfRpBJqN/aWE740x77kdWLQYA
P2gvEfh2hpCuY/lIjT8fWiuVGpgvSgMGat7xZf4DTuqFQOGehbqBa9MD6AfcZcCjgXwoUzHlXMjg
Anlu23Yw2q1pHP7tQwDh+E4OSWTd5gsewhWe4YfUBGnX7nVB/x4Jm9hzTwMhBwdmoZaWj/76m0MD
cZOTo8+OjmTcrP4JDw==
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vAJ++Q625lSIUdmDU8xJbeM2cLm/unLDt+Ip2RyVI/8tB3zK0dztMrxjwwX3fEZOe40akBcAE4CH
kSHn6Qqk5xLe/2cFzG3B19FSEl4+esN2qikUHAq5F5KHEo+N4ixoMdd4WmHDurE0+S72R+irQE/y
q9QjW/pwe9AgGiy7jzzicBzDwduKlDae4kWrhvmT14tXYk+24Nvk61Ui54upeTEQ7jjmtm5ojg9J
EWWxd/d9h5h5dUcUhtG9V6iLp9v/VQOzqOu3yGZproZ02ekWCCS6v3nHqFE97ATVhYvRnHf2BRm1
QcCwo/Co3gGgxG6MT6dLeDbcWfGanRYy+h33jA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 100896)
`protect data_block
5+/efNlIjeXoE2ouRu0SnUCDvmWJnAAqZQm7g8speq4dwi0aYpwRlSEBtu2+sxLtkcxlQeSKIVlJ
tNYnCX9/rST+a/f/IsN1i22dswVwFXAkmqL9u/xppzBtZdMXMXe7m+q8j8wCN6RSts61hZJtB0OH
Nn+2uM285lj7lknJPIhsT9aXIIDmX3Vtwm1Ur+chJDMT7MYC5h10udprvtfpjccdAhmOfUPNCEsT
T92l4Fi2MliwoWOMsmqP/ke9dO56NrtoM3nKS6lnOI8I+2F/TvkU9QUCqKNsoLE5hh/X6mprnB7J
sgUuPhDXvv6kBobF5/WNauZmNw8RBXrHPTR9H8J8TVJRTr423Cd06pIaC9PSm4paw6cdEVMrJec4
mG+mnFpVouVU8SfbSRyZQk0xstIoJrnHNBHXKJnpTfbbFGVLeDR1zH6IKhce6Ieqac/8ynhJTqNW
G/qFUGb3dwcPqr2gw8JoF4WKNEjd7umoVO0InygVq/o5z+x16gOjyYKGRSQLYlCw4mhLpP48yJWy
y9+W/CRea0CbDnOsLRjG37k2wg6KfPZdcCWS3uZkM12hBTdT5OpXkGf9DGivYyRUOm1PnL8/zwmK
KxqVcVb0G8QrjSZ4NnafCD1hOROW8T8N0QtlXprsNaFJodYtM7fZ3JDruXfwD5/et87yQRo275ts
CTiCsSi4npK/HIkfo3A4N4PpO3DS9vE0wh7kHzT2XZKCeVoJFihj7WqoVBD4GTvDR3uo3G/Cqws3
Z3coeQYzd+BmgMq3h1ErOAOyKysYNh7Sfcua2K/yFL3WeevgS93eQqssxn71dbocbr2m32Jz3hTz
KDgax5AljeyxVSIG7cviwDVJC783KmLQoWbUH8dbQ5RD554jilLppbRFe7CHjsUtK+bVQwU48Ifs
j+7EwPG8k1s/+vqoGVP5tFkHIb+0feiS0KMedX0hv8NyntzWHQBLsrs2rxOjOIuOcsJQe7S4YalV
Qhsc337ktqksN/Dq0PpQL+Fmef9dlg9v34YF/MAGbGZe0W5xxA5Dlnk7Btzlir2qb/UW5o8UVIom
kA6Q3WC3TiILWFya3QkzA36ORJsxMdBALX8eWwEH3v9xOH4NlOpR6ZMVlsWbmD/i7dvkBHfDxFAp
eubrU3BSQxG6mT6BgJDnfmJNEhUDnMGwmlZIrWtvzRYByvwXzN8Wgik1RVs+9mQXktfPcFieNL8W
vvOsGbZWCZQRXjGmk6/a6Xaq7sDcib6HcCsjFZZw9Hc8iRF4g5VgfKRDGMkNIW7lyqYBsWxMHpfT
DeOwpkmhoO8OuTe8+WGkQnWVTnf7A0vW/Zd8GHkot12dyuvjDugni1hSJgYiOy1MMCEik6B4PszQ
eQkJmpP6VFMU/PWc+31ysPIC4rkoBbFg/y6hfdPp2K+UM97/6pIJBrRFsc5vs3TExYgOxiROH2EN
SLwkZOT9J51yjh4xvjqPdOvLN6zuQw0qppdq6m13KDsxtYBWxzjvOg9OaXzHDakMYlvJFa2eYbcd
CYeTo/Z2RoCBR3udhbnmKYfKi9Gx08K/NTQKfEZO3vl29Ecq9g9C4pM0WHT7M2YURcLpz2/0kk5Z
T/Wcs8ephkevfyEYqqyJ00eWo8wmLbXSiLJSEVlFz+fxxVwUQR6TT++o512RYQHZSoQEYivK7S+E
1Az6S9XxWKt+wndoMfBzvUON4fjCS7m3JBLHZeFPrxnxxrjUxB1X2YS3QEOD8U0+JJp+u38Of291
733VaQslhSSd4u45+L7iuyp2Lb5qRrLBxXxu333oUdfrQ9aSXkr03HoVA0UJR3hrU0OAHuro+xpK
OxoZT+RpexKoaQYlpxYrRfKfRLQLwTTppyrA8OkOkDIaRbvcNnX450xmaRfNTqxgIQjgxebujiaE
lTFgFVOttiCKffW+boZf9yZK/4FEY19aETcotndteycLW+4YZ6Iz9cmDsV36jLVHOEL3f0V5bNKa
goDjQw4c1AJOuIoZGEBupJ6vQaD/ck/DpFKzzs/BCus7/SOs3JJSAdKrzJFbaTSm6KADcJIIxyTE
uTKyAYxGrxRd7P4/JlY/PBVwxGU7MbQlpXflZ1U1SexnW+AAjWUzOGkKqD8ksltb4rlPOovsprPr
Q46GJgm/JEbvoAvSIwmthocTuoTlKC3PiATyVwWpDssM4zMyU0IltAJay2MpsmywMwzx5Ud11QC6
nB66EkBysSra6ZOk+ECJjrCbzs40S0o0GEKFWdMfkXCvDdChdk01mJfJVZPQCXkbA01yr/PXCIM/
hkMxL9YW1nAp9rofJVZ3gkT3h+mZ5CPhHF972FKjEFAFfYD/pn33q4ST1I7Dq+4O1jPo3ogvPOi+
a/Ey7twq8fED7h0XZHTSyadR3aUC+szX40pe/DnuOUnEW8vKMJBVn3TpTZ9wsL5/GD0mKdjAF+kI
rNXSDC1l+WlkNkGNHEfsmkXGjSxAuNT9ovJRPagAm9xWcMzk2mhI+YyfZRsiOHvziEG+ZWMI7Chv
VoOUSbqLBqmRjDaBmfmGfN19aXooCKTydcqc0Ly28OVP8cy2+JMC9IlLc4XYWmEjQR2QanMfxwl+
ns2+7srLJB/95gm0Mwfo1eUtxere99ZOy+8XGIkkSXSe4HNpWKgwlrV+bk0Hlh7pobFfrzBXB5sw
KcTCSMzfsmcsmDiLLojIm2lGgAefxFRXud3lfrN2rDepPmazr7igEHNw4OT1rcZllxnvpgPSHyCb
0r7+oVdbiogaX4WsYev43fe03B8GJWgUS8ey18V9Zi/POX9fnFroNSoDNtGYKrbzO3r9Ur5ji9Tp
8U8I8rnizOm8DJOViFlOMp5wHHw/5drgyCg+RchuGi0QvWGrzHePpypgpWNfTDZjthdE0DnX6See
bL0uDmKi8mSR/pdRUmFGnnsqLtSOD/wFUyFhM3mW2rKEgxiS+dq+C17gR+avRWpaX2YYUr6dLQEr
2RM5C1ZVfUcNkI96Yl+UeptiDStgHT+d9Q8PWDsBRxsMmjsHnIGFdY0UbWkxJL0zTuqKSkqMl9aD
amcuAXrxjCoUHzB1487S20k4WacHknv/QSVijNd/y+b+629QpmgEIA/jjWp0ZRfN7biQXDlUqRTG
WMW1cXcvrfnjmpVnW8KhC5FItQoO/AhSZlKtkXumvFbW9bgspBt9YBF38VkbZgMAMCBqMxkVsrW7
5htm+5xMCHHvBY93cxSLTHj/Sny0r4smS8QffseOp12GzXrrve161qxo1zYPvJgLWVl6EYdO+zpG
LRhVLaUXmRljVpqkkFHFlfKQVmnZCte5LQ+1Z4IiMGOzztma/E/MtHAZacEOqBU0Z+ki/zVNYXNi
g1Z6jhglynkqAB/zo5wbDoxlpv808e2RwxXMJEr04emvMyq1C7IQ3rZrqX83MSrYCuoRobB3C5oN
p7CEdX03jJ/rOAPxZYgRPYc/9Cd559759Sxnt4PmkOkWuT8ddjk8L41UR5Os/sldNK6FqO4UO6IJ
4uG4UOroKIhl9VK8O9J76SQhuu/OKdNtpRTzbfrXoZXGWPdapY8sY92JTGVV6sOgoReldyHUvn7u
SXJZ8dzlYewLZLNHibLN+doJpJWNiSy3RsbFSczii28a+4JI2TTLtv1vpjW+xeUmKU7mLlxo+XCv
CCkf8guV83nR1gVEFil24zqBoYSUUWPZdc2oTlpndpaA8poHZmgpWUWMi4ZqKvyg/bk5lQHC0pw1
Kn21wnn0VRRqG3jKrCXjp9iR4UmZOajniuQsm5uUoFQIwyIaYfpkq/275mKDaWy8QLZIHid863X3
R2JMqn2WHmcLVqEZ41KS/7JAv6hvfR9xl/0sSaaDFKosTbWQJJDqjA7qJ12PGDHsFAvAKToOcVG2
J/2RU493pliGUTBdYNZSNkp+v3aDbqW/g0PgEtSvFguGP6NkfsDvMpPAyC4WaRAJ4Chb3S2gGooM
y52Usg9R/u7kig3ST7dHNnMG1Ufrwjo1D1uhiCpKgGV/5IExqh0cvj9CIhK+57wtAY9Gr/NSAtxY
48QIzPwaVuItL94F0C4PozU7na7rnQDiL9up3E0R/fbuxI7qjY55oE+DxoAiDTQRzj/liwNrawJW
9jXRFRSiv+W7/JW4r7KqECjfvIAFs9YquvUhJ9ArQy4zsujoeDZi6V4oLB9zdXRSMQ/Um57s4wma
czqdFc5OK2yEh8CnHJoRFfDceC/oqteEJ7K4AJjaqOLrHNt7f3LV6lydgJHDMuU49FG+5IJfc9RA
WwDEnZQVweEq+gBNvGowR4ExLMx7w8iZ/S+C4TpdgUKaXU2x+Qf7WGKQwG5w4xR+e1uhDtjmOBB3
onYWJbQY/mPcRgJRZc+ly/Yr+NOIln9H8zs72swAnQ70xopPPZ3Nupmfq10mRVfU83FuxsrdD1Gb
nXRLuKdjSJWC65XtmRkTC8GNPzsPfq+ptq6wihuTpAE/JLzE+FKbx/98Pt8WXRksL0NZeVT03t3R
bjYCCsbCSN0RhrO5xTJSw3WNZ9xH7gU6sXx0vkofpilVG95u7eFNfa0Q42F+A4A/kjOeGain4FPr
OwyNbl2VljXceX26qekR8FUSdYn96F4yDZpEPNnV4BvDAMfhCWI2H1IjJ11vACoaqxrXOfZm6+sP
iOdfEdKVwCSwZbPMXN92v1S3UO1ctFCXSVcHXKxKdzk+uS7M4qhdwpxMVE7xJwLHXcGXuoQ3smLK
9h4IdIBSnpqiJQWR3pBA7ipfC+cvipb3dNhDw306qk9AjhW169I3q4sQedKth/QzfUJp9NsniM7x
DEYO3VyeD4s4DKC42by1FKuJs9wpecvFyCOLq24O7RChJFV7WbWwQCVUyY0KuyEcnIXLbWsU6Mf2
ahFjWm+zLhe7gnZBXUNxMCaqvQKFNbJYsfNnQz0y1UMOxstZ/mppDOs1QRo7atqgH6295Ov/b3M7
akg+QuzReYFOAU6tvx9QwNuZ2uGge8TeWJEdzZUDHpfE9Gitmd45q5W5CrXeTMHlml0teUBr7nOe
HHh57qVHe444EWovOf4i99PdK1ajki+2eBPPKszFSTr5eeUX+tAA701bu80iHzMa13BefIjkAuP1
aByxC1FhJlYZWQfHvpOSi58PdQaUgyqkJTa9VIGYvfA1qnjVRNc+GIGCJ3WWnXTDZxnTYRxyGVwy
yLAz/Um6uAWly64FAt178GNQQxxMezfpa1yJG5esnXsIuEZ5IWsO3JfJG1hYYbc7rT2jOPuw/2UR
3Nz270DuuzWRCrbNofzj5/0gAFdFR9kNiDTtK+OumdtEBuWp7KSedYV2ILUPYJm/itbNrrKk10Bc
U+i7V4UBD086CSKMWdP8l4LyQUSKujgT6s08FeOIXaXP3RwU5BqbgztV5blO1XHVDRPNS8SyErX0
84ZhfWSEpAaAFbUgnnJBrUUao7naHliw7nB89W3LifhvmwyjQBuQLuBmsCRKMRjULAo7f9eAbs7l
YN0t1vXloHPDPY38n2qyXfGYtW9m0X/GN5u8lUNzdy//wbShO3/cTKVKULtdhtuNUEfculj/NJlK
9qthURvPsp6svB8IlBYg8QGu57gmwxDOb5zjH0wf89+kshiiX85g5ngykR4xae8dJ98UQ/UynbYe
DqpMpva+mylheRvKeKI5N2riV6jS3GjuRjrDxjL63Sg7RUQy3rbKpb8D/V+R5MvA90soEQdk9b8f
cuf8Ls8QvUt6GD8TQ1uFOIGnSu4sfn/L+3Tyxvj1XPPef24YLv/Ee5gd7I499QQa0Pxiz/DmMKTL
qnAzbrb8BVC9GVmzCbiClhTcs2OQg9Aiy6FL8k7Tv3uU+3VxRd2Tj7qBXK4dTrxB93l38cw/dOmL
znXlSGf71s0DudF58B6e+wF6WBjZpj3tIHJmKi71tyP6hMQyrwkELiFQP85BcoEHIkgedubkBqqc
K6v0OTYrc+1H07fA1/JKPoKUkzFIq+gESeFEq7xw9oujGClAR5RkYJ7bl+Dk5Js68Ld+3W+futy/
zLnxrnDtQD0xpbTsuTtYT1kc/klvEZf+GtiVbj85E88j3zPjwUqwkU3eURjWj6X1iQFYI/aSzamI
vcLR47Azej1kLSulBfnoMP8L2IaNq3Xdyz8GuuRef8QjCpQRcrY4Ifz2EtDp5FZ3biv3RG1eI9mB
fhe0LSZB+vN3zrl9owxhVFAeoJa9Hr41Ha+Ic+jL0EXL2WbBGohrZRPI8D7GgPNfWvERPNZ7H4Rv
mxRZlXH+3z/i16jye0+zSpnx/Jy9XTg8t/PthpVoTNISAiCl0rTCQvatRxgKW1CyTEPPANWUgUDF
pZqbcyoUXihzdW8hoyBMcxpv8jVdhoGc0tlfmXrk+eNh/NfL3L8kMYMeRtFuR75rzeqGtVCvqnmr
Gbs0wcvhvtEz5vMuxajySDzVZHOHyoROsAY7ToZ9FHxmDNjhZT6hvP5MoPvyUqQjAebYutwlERoM
YaHXTuJDWrtE7Is1+Nf9tQ3NhjpsQtph/J6nF+xIFC4Wz0lNZNLvyQVNEnI25YYlJuCIcdHhrloT
lzqPYDaejhpkjVHI8AEUgfKguxzbaTYfT5HQwRSWc3pU8f3b6PhqoyKQwAHIBiIuleVNeMYRmF6a
oYgNQRxCOtYqe7i4afeweLs5DAEWXkOnDufTyLit43X9kCuOqyOW/FL+IXo+9iY+0gNwigHTvUzM
RiTOPUpOwRSVydJKDDsjIHBmXdpAwJTQHnjoG6GwpTUBvMedv9c03UH9ZpoA0atmJ/Za4wiAtgEc
H16gNMLMM8MuzlXcuZbH4ACEhlAtblrir37+EmnRu2y19N+L4BzEnzkQkf/0FXZ7HIvs4sDB3e7C
5sZLq3mLujUmDf0+xGVWFxFzrcrKuVHk9Dt7pP1IQpRFVjpnF335NHk8G2TzPgLJFq12+w7yxSVr
cvHPRQffRAQJy3G/Igj4XCRRNGJCNH/jaqS2PKzDd0bg9eN8x+4zOQEYzxfHWjb2TvXxaM2ABP6Y
d7vw1YywQEbN6qr0GsiU9NxiiUo3YKmnq4hmnAJFo2jS6BHIMgFJxUUi/MkZ9pc2pQSQGvpGycY4
9iQNwu2/1muE1nZdTlalWY7GWajrODRc7CBlFrVEnPbIdRLwVqqQbfII6p6watdbcP6+P9teYjGy
n2Uh3Mn9sZsXs3GE3WGCn8EdmqFfq5k990ojwrwAD9cRM1pHkou245uNziuCHLK2VMsYVHV9iseK
/Er91ePLMUufWAO6JoTwYXdEnv9Gj76TOpOQbWW0OkFNJn7Ap3YT9xxR4qpMW49GKpxlBDjYVoIq
2CdQJh/pi4tFFCVfMrXncTHPY/oMu2b322WqCU9f4iu/d8nUymnZJKCca6FtXgy6E6wwlmUNWwMA
2VXKeextnLAmiZTFenAIg+f2gEZ4wtaFU1x4BHYDPUtabnnsEOQa94WcNxPLaI/hfagbrpYhz9aa
3PJVHuCUq30NrbkpCgxSjqvSjNCFTGRQUmOgj+plygOtNukV5ejOy3ta1ZG8+BQmWE5R7ZIrnmki
EpD1WMOGwa49xAGxOj529VEBaQ7VeRd3rq4f3VsG3fFJiSCXlH4lhsnRGyx9NzBoNvILdUNcWi1Z
YJNwNxVKdD9p8ElEzPsQ+Vv9d4RnpCDTz+eYvWJTFDEK+/RFzRxXuecyGHizqLiLX135okUjfqqo
KC/KxrXNudzE/VODd/85FBIn3umDdjvNz7VrRp26CKoS+WrCH7LxKpM2QfdMeXVnFipa163iRom5
LiMjqebLxRLNGky4XDJOvZsUNhWW1ys9KRvmRh8Bwlbji/rWRCuxgSl4Y0Ugs4f5mEDfjzE3sKQD
fqV0bslgapYAL3MccuqB7Mf2v1uUnWFSEAu05vCj3kE6IPH0g8jI9YJFEYwSb03LvTCR2oc0/1Tx
GBk+4yzBeThUGT+SVMQ1gwvnYcoMKEO970Bglt++yBq7SZ6dIiJ6O3auAgkGIVB0glomoSqkd1NH
7yqVaLJKrK+pfdD94btLv3FuhsAdB85GG/W0/+rDMhlUF6WFHxhuHSgCIr8b5Teowaf/eI5s5jag
082746En9VAMegAr9UD+LW02IGl+hLNRR0RHCPzF0Zk/ZIXTJzevbwptjHDcWEgEsBF/KI329c2b
PQkubf0RtM80hPiVIIlXftIu2xqPIg4Az6zCrrqXsuPWaRISihcq+N0JoEGOnxpsJybFoFV2ca3q
4EtTn8DpTn3Y11ceI1PwxCD1720u/XTheyKKwaR0rXrNLvs6PMjsh/AtgAub9f6Yix5zC5qQKu+j
YDCXaUuyNtJYYhHTSJrJG38YLYdLlSkeLg+HxsSi9T2AtkqCLZkab91lTMPZlHzuB/sNmzxyfOdF
CxnZXmDIEfz7ItyQjBVXPuyfAuDuYmyHh5vZHp24RLjTfYQKFfyR6c9nHYLIKstMjS3HbqGrjN+l
JhwaMi6LagEGUg6jh73nreMT+4eaG5D4o+/kwDyvtGdKsVcOv8kWbw/AUB+NaECkas+Qwm0ULK0G
WpewScOTfecyocBfFNDo9ISzgTPkZ8dmM1bBXGJ/c1ovWCAlZcgRY2dA5r0mxkgYQU/FdSl3B5w9
rGpocond34EicYXV1PF8Q47jtPMmD8b7OSoLhc3u1Nv7he6TGX4tNMovSKdkq8ncllRwASfO+M+K
F0psVOQl78mxUb8UwXa4SLsFRfclqymmwAbg/h2rIO3xcBXnRHl1zaIFIsDng7lWjGYB1daptwtr
l5O4qq3f3g38o/o6QHXaa//pz+FTwzXrA9hL3qbfnp+BegKJtx6Tj3f59In76ASCpp/Wjqh+Ir7h
gtOjRfI7e5uF9avJ//2JSEBGxhBzZK/UlGDtt4V/7OWmEnOsfYSNXcd2RIS8llNNaqDNEEXeLtmv
8VpSV7dS4kGA/5y+4MC6bsdSNfuWo12Roeg9itK4C+yUA3/p89FxuoZcwnMMwQquOvn8zjCJTeil
Bj00acGWO7Wnv6FlyfsOGqYouTCcXQX2KdcGT4WmvWfBNZ79Pg/sDpALOi+DjVi7wnpwQfD+Ep3h
dn6ReAiZLiITepp5lAs6jFiKSHitNJhAmf1gEd5pL/6YOfA4Xo7RWShgkxPrdU4WnLh+4KNGyA2l
YCRC404JQ2mfRRHQJvd1Sqhi07KE9y6yuAyHWMAdC9c0umuBqM3/LD55u6FfNQQ2fgoFOM5miTt9
j82YeNxPA+EVeglZm6giVA1e/R20cU1RsVGRjMaDORGkfFb1Nn4Khu3oC9iQGqmwJRCbP7AQrLKr
YC+GVOpljBEyjoRs7gpHR7+TyFn+fjgcK2bwcjE91I84ft/vr1uOZPjPpbUNBWOw/BKutbglMPX5
Y33EqMzWC8akehzAHYhuGQ4TdmTVBvukn4SW5DL3W/TuA39cesdD+1D3NxfcHkVNi7xDHe5nywZD
dS/aDqfJ1MkxBaCjNNH+UlNv2SKIPmpdvS3pBPBV3tE9TCyOGAkY8pphed1KA2bd+2FfjO6GzQaM
l0fcxxHIczVd6sI9HbAiSB5Vu7oMgrRlSu8Fz/Mdy98JZYvlrkhxzzipCNZ2JvEMjaxIHriTnS9c
PAVjiAM1gR5TVAWs+CBei4VHgMDRuLOiJJBUBTXL0+ilslW/gfenzPHZYJFW2UV0tioi8cVEg88g
Nb1JSA8D6TUOL2BkjcgImd+hqp7rQetaR6IWF86XvSqcfTfH6bb9pyOS4ytI3qSKpkdo1E1sfCHW
NasmP33qjTds5npUSUy/lr54EDyawvER1jOsmAoLhqJTclk++spwkmzQls8E42PJbPasf2uVA4Ak
OVH+qRjFTv+ch4gMoKQ0tvDoTa5lysKvIe9s9DiqTY9nuSlGHGSdThY3YjQ90oe/TcgCDVadL55O
jWmTW5AMyYqcBqscgFet8vIZOJQR+g3X/CYnTqkqe/LkbRv0Gr3OER3gnj0T98f5vFWbcOK/9okk
FzCFzUIY/N/WYUR656fnycVobN5/BeFpftDiIJnrsBlm8L7VR0O2iBCCzGYaHXaWj8AfG9o9Z0bY
WGMEmRv1tKYzK0KRGC2tvzg+OjypPeWVzSxCHpcCE3NbNDsRRS3ainGkKctnsxvczGot6fwtd6i1
APyxrCHU1yXVqOkI8O0pzAkvprfaXhoQmKZNtlK8u6/0B1Y5+/YP0FkaDVnKeN0dZKhBEX2d8QkR
evHeQ3Qo+nY4jKchJ4LMjQaZXIaD5QYARKwBQhz/9QU7XlFJh+VnUNu3w3VMCPTkgA3Hcx1ap4W7
D1Gj+K/xUwXlqvaLX+UtoWleyV9VnS9ktaaTCdpoNBT+qjia3/yYr7F9CPchGCSg2T11gH3OjtDJ
enWgOOXw0mjHvjj/mBjPYRPe1+y8UQoGOo7lNkOXI2Z8S02VC2cLj4VY3WdAHIIsfUsEQhBg5j/o
m9gRUrkqzgoUcr0tsr3qOMCYSPodJtw65usxtpVal2kzlMzy5X4GcKUe2dizuYQGY43krWDbeGwY
K7mlXCv9lFMWHMukSWgOpP6fQPE7XWlXzkhBi+BZTOsljEXHy1XzASPvJlHuCbyyUv/j9Ij873NY
Vt4qN+VWrawjx2i7nVmiaV48xmClDsQha83QD8pkchvUF4ByFC5n9I5YRj49xZ5KSom8ljhZ7UaW
iRAungCKuxK9WKkjBu+QvbJsXka8ZGt8Jd9K/9EQGdQfLeYurWIOnVReXPyl0KGkt2szGRH55140
E4ih5sica/jNCIobBgtkyagcRGZl3qOU7XNSc/AKyNP1c3v4zgSL+YUlyrd7WTmukizBY2AmJzq6
t9kLwXelcnlL6P69ym8utNASXGDruJ1sw4hFPBMuVlGNycNYpr/ykIAp7hoDSKA+IWrGJf6i9hu0
+qGFAURuMIRi04rx80oO73ymaHSlRj+sNE5Ls4rg1rTJDkw3oq1w4RfJwgEAVw9EJTVWFE4Ye5e0
/iBwH3qy97cQ0dl8GxPcIv0BhFif0qjkcVE+XMBxk1/UZ8jLR61VQFBZcnOX1jOT9CitSo3HXhPV
DxFKAYXJ/DLg6PE7O1RX10qs2h28SE05yHGB90RnGD7cPrAIZSYsw6EUvKaUtMv3jwz0WI28kKNH
gYJv+mpr6lB1OwA7TlhwRZNopa0gfbCCCEZ2b8l3aGe4jTJyukRDldBgi4fWCpbHTP5PiZmRy/Pf
pJUVL+Kdeicl7diiQX0g7YAQQCyUNv9w5GdjbXIHM80d8dJR+rcHxU4HmXqmqebpIvYVxpJXM+0a
kWTZpLZanwtbdtHeHN9G74n/EE0MCJIvoUBgXNOis+bjYEq0+mpMcBtB4s4cr6xulJE9BK97KYID
HvJjQlZhH8pBXfIjdN4UDxxzS7xrId7abajVJ2IT96z7IX+wBlsOUdFKnx5sPEnkpy1g3c2zzV+A
rFTEjW/0/gxrmhYOsXDHaIodF3SV0h/sqYAoaGjWpemZPUwn1609ya+ELqxKS1ngtTVs79LoKK8R
s3HytjEf+mI5Dvn0ap1mb4IR2K2aqb9oc+UXacf9w7/jSEzj32ey7wf3iLiILrxMUXCymW9wYXw2
4QsCmfSSVoBvxaHpyWIe430DmPhxndWIIyqNNQBF4s/3f0o4PnQN9oPGkW8d/e1JIX2TRwvqO0Os
g6PCJkCEIVjA85Y18wBl2uwvXKtxY4HW9vs6ce1OdGDnNzSdmrc4/wZs6TKsXqsls+cs5RlJCQo9
8iQafLUdJhLmW7tWSH4BxuREzN9PAvmRsF3ewARRXIs04f83dLjfDEL1NSRD5Kg77/HLk2cGka7A
hJt0dQuWW5O7Pp/DbGbKFgDbmK3gLHLJxnGlBiQ9y/zPqgE44pOoKlJp6njFWq6EzPx/J1/YqOlm
hBeD1Nsy1SA0aUQdYtLRKdEI4R/5nkyZk63B0np7b9OBHZXY03JjPI96/N545743rJNwxDR6ReBa
E8QLFdVnklhEEeTcM6T5g2YbSk82FUylny3TOyTo59s1wXPFuac899x3OGs8KMUerRrUFinu8QG9
xoFWH5Q20j/MH6nLSeWdjM68DtIZEP0W0JteAFUxvvYCAohhwzTf+r8rznZ9cKcxWkAmgVAQmurV
9WT3UuaeKkNpB2Ybd/FtwRjJ4H7cpUm+BOw//A4xzalM38VQ2LclOsJsEOUF1745VYipQK3KHkgM
gKo4yEUhXX7fUsdyhoREFOLuxsP+HqqKAIReYVfpKdR87gs0EuBtsmzp5CZA/4LDOrFZ0jFZ36QW
Cd3OvSJDgn82xZxCZtiBJTulFtYjuo2pLIIoBKhSFBLKkLKNWpeN3OFIrZFN3tF7xGKW/ez8pE71
pqTvgqs++/P+vn8DWUXUynQpV3P0nPDXFbUxjTtDEX+Pg5jlj6OqEURJ5vX4x5AR618yFsijYSNE
hHUKYJFvhSwOxJBKzryozQnn286d/G3vrE4gMG0UvugP47HNSRBp7nh3T5d0emu8BciKD8MPjM7T
U1falTB0z96fWl4ULHpXHRUsw6cI2MIq/gCekd7s7DLSK5za0gC9JGzbYrTY9zh7CWBMewjCYt9K
hHhv3ozRFjyxVgG+PkdclXmqhcwx/V2zdsKz7CwrZdCVx6EfCXqKyR7fUd6MbLlkpaNsZxld8nGj
25LoVItgVD01wkhCVMtAzTQ3yN797gvDNKX6J9ZkMr11wh40AXLQvXjHeX1p7mndq7ICDHEeGU1J
8OgCNTi7Cb/XuYjCQNiYjaH2SwIEw8mKkcbi+C5Q6Y9yzpi17mLAh3Ie+ItKTdl+XbRXCMhg/Tv1
TVr+QAVELnDE/PLnum6cog0kaZTzyQLmlR63c6DT9aniTiXCGewd9rhZ+qz6MdORSF6KT17GdylS
XMwtspFW5ug4tyuKIe9IlaFWm6B3DCcCz80ZVtx3tetfIm5tjBxwu5cnXfs6OKCxpdklIItsZ1OF
N33cA20jeHOaaPXRYB5FhX1DerPIs4kzDbQOZgKkUWtvy3AUp+X+96YGC3YZfw2C2Fighk0sksMr
/CSo2/WGpJahKReF/23wf711xHkBUdEgpj6pnSJOqqlkLO7aPH01WdqdZPH045oW9hqzbSoDR73I
haky032kFk6i+Sbbdib9wMnazpREinNPwKzYZMqLzG8IvZ8INqIY55Kv9UQQ7liFSyVC+sFpmrrP
BWkaZdKx9IAwh0N+pO2GkDwCm/YA9mhWUSowkt0pa0WuDE+uHPAm97tVoETXIqGypSUHlRo1Njfb
Rfjq9BcXWU9W3Bhkc70clgKWE9VNgY6ubx3yBqEjWJ4W27SMLDfn8CS9HIg/EXe0i8czL2rVLA8n
IVilt80Il38YdNWyaxs/1JbbrG4eQUqVbs0tEgH1uBjITXHi/DNDFO1STb3N6iU4UcmaURttr4u+
26PN2QLonH6U4YNqhE/N7qCA7c16nyjQ1TOr3JkHI5HLDEPhH/DgVQDOxlbCpXg/MxQKfBgnvVwH
ZAFU1Sg5JyOLoK1hWn32ZCWwkfLJF5EchwGNZkCOu/0nxgG7oGesmEkRVo7hPPHuh3hua/2yU8BB
LC3qOtBuioJjNBcq4LWdGgi7FFo40btqPyJ47LysvgEQmtimZhNj2/N1jaKhkpRXjOBIF9iCY0Uf
7bahwwwh0HiXAlveufnxe/zb3ugMGa6giFZXJcirzxHYNVnVxTkITbNNpTjCJWnpUiB3y54A6yHI
MVE1ynWQh8Wb/MWpIUqNDlBrRwHf4l3wkaHRF/oYLLn8BtFg7c75KPAvmQwMBTo32GGHPUIz8Imn
izOneZahBspfLXg0ZW+TG0Q37ZlXMK412O5h8yg9PlvhVj4iPeCpdOxS5DRchM8A5ATUZELmR2k2
ftw29ufwtB5hQ09AmqloaKZUjd6E2pHgfRbkhkryWXfBXFYdrINmxpKB4Ih/kHQv8FqEuGqco2LB
c7SqPnnWOg///A1fT+MLtkzkQa0bL0M5vXPisOHT/78uVS39V432FC0AHDl6Docks8WgRDiRpF8j
jp1Mrm2jbGtnGGTFRnPmtpJMilxBWnVMdNtpBAY6FfDk/MFQ//Q1uqsR7gCyFi9oMqCoyN5k8e7C
LS/V6U8EBrANxvEU0qzbFU/p7M2ugeXTf2SiaqIiOqNFvns1c4PIyXALvg15FrYTLYK+v6OPLMqn
OggHWtQVBhSPsomPVmE3c3J6UqJa8bB2GHC5LtncMP31R0k5Ql6gyBydUf8fm04DMbsUhJRe7NvL
0UaiJhgLG863nXbTVEyR9JNiBOSSPOqceZqiSf4ZM9in4cq0bctc1F4foLhSoFOhT8bsC+OfCDWR
sM8vMTx6JMciA6kxMWgSGjj9g4zkWxxO3LvJ6oUk0PsvJcHwPw25WokXKlY6vZKM8ynwl8SdJxpz
Ccg5Gm2A8bG1gnDUEMMnc7W/+m6Fr/BWaIQXAM2Q9ywMlA2Jv4lxu8h9UjCQNW73wDwCGWODCrre
XGpvcabEbGKchBH8zNHfCNtwtqu2PLsVmNEshXqbM8/RnuBJJY/cJpEcjyKn2ifbeb3c0U4MGiYP
q+Mp6ssPjF1ufu5ESYS1SnYPVfjPqB/ZL5UY2cSYpdzg8I2OwHMpJBAbEAJylUw/DCrgaIlpFUDP
XyIV1edkm3ieLTlAXGzTpR88TMWVBnR9EGQ3a8zhnM+YbxH6f1cFgvPQYjqMmclvg8LiZGMC7HDi
yZund+Kqz9gr0mFVGRNWZFvZeIFXdmHIOdAqTtKXQ+hIo0zCe/5d+kW/KV33sjtksJJZzO4LJpSV
rHe9lxmJckdUaVG+1/sH/oezBvklh0aOP4hzKM1yBX1AR4XHMuDcf5Xi/YyyMMwSDIuyToHqzgL/
bMZe/YEU/XBXbSTKHAuASw5hjROsa3HPO1jWpFWRghRCp2zeucuLXdpum15syzWGlhKURtgRGFKN
RYlQ6t7TQOk8qvjgP4lY+aPN4Ibhcn9R6j2/difVf9gLD0JGOyGGTR11YXlOSSx0CcasJfDU0ToT
oAcB85VkWDN75MoW4TLOrpV+qN1tA0kFEdZVYVNgtTvBrXyieOH1BLn5Wxb12CdB1S7KZEMAcdwj
cypCASdcD4Voo0Dsw+hrkT138+pvTPmRs1ndPamuwxuC3Q7aW8tt1RmkPI0Q5TZ9JC0jVNBPndM0
tek9MJlu6BbaUbUgTSILMRDiYJak8th9dIdcVpuGl/PVAMJZDzZE4nyEH9Ek88ttTQIuqHP6FAlh
OcEN8QkleAwhA0Sdo2TOle1F+e7IeNyFM1NFko8qp/G+/JltbIrs2zgcUnwMCwqUU2LOaYQaEX4R
33CpUSw14StawYAqnh/Irt+fNLXjbOrd1OiGK5rp6F0YrfJlZQgNK4sJ4eY0t5EbZIx3MWziAdyt
H5Z5xf5m/wSArILWFp8UMrZSce5yzK519rUxgou0NaGOtgM7FY5IlS2JR2gLEC/zI+l4z5+I4okc
RZBOzYOlCpCQgd7J6fMP0XZnXtkVmuvDyfoNbEbhC324a3w/4tD5DPFXBLx8IekGLbi1oE1wSnX2
BJ6/PvfUPyLzaZW/rfQupi9B3KSXakvUbApTltl4QGdjhUTY1cn42COe7DK0EG0f79YdXAxPG5Be
3dE3LicHAtIYHdzuHh1WdpEWqDE3KnygYzeMQjrV8xxhi5drXrFepJozDflrmNaFePk7V5yV3+3e
oGoPswK/jJfEI6dvV0Ce9R4hMLgBYPDO15YO0MBus1+qHgQlIETUoZ0J2isyGLzsXAhshlGi0EY2
33L5F4EwbSdJFt2zDYzEZyu4wTfq7a0jmeQUlaGGQfzpn8sBcy5UCoGIE6I0u43HJuZu6pMvx7nf
wbr88/bCw4eR9i72sZk1lwLR4GrZSRbRPP7H2rZVR4Wgl2fRRLAq79tMe02o++UDh4E2pHLn1OhY
4/bTnnyyEZ1oL39YliX7zBJPK7VcmU8+12GkOjX+UMS+PRFVDUtf4alVA7x8ZtP+yPOlk1Yz4l3X
exfmqF7XwQTSTlTBL2uHdtdchmgmX3N0k0AZNe3X7dmBDVTO/XS3ytgsFvMCIwdNR2/QrTW7YnCk
3muaP6OtV5bzWZSbuP8yJzkOOgOB1T1SlXWqEpiYeKH0COMhZqbjdhUUyJPCQQVpIa7O/sUBe6oF
tC6UnGNj4Dy99B2kjP1xacKH4mCeV4CZ/xDjqczEDjrvBBJSK3SLoHFqaBDaJmok9PDxqecGX7Yd
eiSfEHGN/OXnLdyqN3reWxD3Po7Sd2vsQSDhe1KVTpCjs+FYe8+93WVq5HZLv7Q4zubfTQL9YgwB
SNuTgPUj46p/koboiRB6woYh32dhbQMzyEF559wXdAYa5kuxZxjoubbMfOUYd9eS2XSYzuRm+oqE
ib5vvZfZOd2vxqp6Lw5wwNTf2EyUdmkRMuwy6P0nWYFj+r0Qu3EuIVJtdygrjxuiTbELNqF/6p5t
wNm9At5nT0Mm7c+Ul/ydOeTf6xgwW48KkmP/yPHdAFSLGaasPKh6HwB+Hj4PG/QdRco2XuxyEl7+
iJayc7LyyzGZKt0OFe6ujo73bLcTvqJmij3KvXQK/lxD2UcNln0h0OICPiupLu9JSTBM5/U50H3r
K7iqML1kOzUUHmz3HcuuEaBB8fa9XonjgHDko1etCMTj1yAmnN+EZpfQ2qolqEQrWSPAaxX0WvbE
sI9FIxazJ2aleECAMeKvBidvYnEjHz1JDKtNt+AKtruY3kNgHKYYqLgpXky4yelxQ1W3gl2YVKb9
77u2WxcyV5LbA7xi0i/A8aMcAsrCiIc3+lcenUgvPQqLFpfzkvctEJo18FXebZedwLnHp83dRwet
YnWus2V+I5Rp94I5EoSZLGuy8Bjf+NhiofIWm4iYNi5kH0Vm6yFRxqHiT1ucLCOyT04FCY9vVd34
bKx2Cj4++yRO4Z+XwqOUgQ/fatdo3KMjSDZCBqWgWf+1lvPVf0myV8AWNXEILzba7RPacg93boQl
hy5O/DY/rxFQ5tsptoK7uzTA0kyrQYTnWuBj/pL2FfT1n7tzq6lpE03NmbpARxHDv2WuoyZlhza2
uls+qjuzd9skLF+zS1NxfpSF4dHXHmv06EPe9T62FGA7mEJ+B2Uhq5R1jMXhhKK4jLVkV2xtj6s1
Xb4fOAnVyQF5oXE39gQr6VhjcoInQ6ubW8swOo75uJSNrX/o+cpuP8O3jbBqNrgOp26mDPMNnWOv
wee1RqXo1XDxD78VYza1xQ/MH9oySaMbe2Ob8ejusIX1tLhyPGbyo4ar8XJlUxkIoExGASAG/APJ
y+adX/mKxxLNb9HmddtdqRq5safoj0wAaQMElhbKAu2LooqsXntz/MPdEhjICko+j0udjFBJIxcF
i4qlH4NV/HFCbx+weCQXEDXIQnxIY1ox+HFVm33J6MyLt1B6duxTMuCxwGkkhSLaOk3AgnM7WsT3
cyqKeSDAmSOcm6xpLMnWX5BvyBTxHh4joCTAsag/YKJYLN67Yy4tHBRPbaDtSkkn6MFnytzd8usn
bIT4mgxkTC2JYt0LisfGMEPpZo09RqtbEDSJWFBwR9omz7dp4qFTwFlF2hQGWRKKoksjQ4OCHc26
OwO0DrslCJWH/cO1TQg4TTdP1vvOIbN8TdFPlzPNzupMTDKZasv6VhOZSvH+jv3de2hJ37860Au6
4/WRoKJSTMe0aJeS0BJGQulCPP55U3fKNpW/H9qllZDZQUF2hw8x3DNRq3iWOgD9DyIxvDzhrvfE
nPfQ7y3J2pmLrKTymCRVjE5zEdb96P7GFvW1G12896z3UOn95JUJSMRx53ikMj/aMNTXuneb5kTj
AuT2gAQ9RoDN9m27z/q5mqXc+Msa36suhnLWZNB1tzzWc8UzRpNhTzBeLIe5JOV8ds0ryGYKpPbR
1gd1qiX4JgA8vK/xVVOlCyak2xdjHGZQ+VPJdzvC/DU/8bKxtCF7EX6/ZwMHPTRJQwmrf+5I4hGx
nOAndCrjphaCU7N05W3Uc0/82feMJkDY1jA7ibiyGkazF9dXIapqmBDyWvJC4Ck2YB7+osEWlhGk
AV2QXdDiyqjY3MNVieh+7rOOWGK5Hx0wpYBQbZvEnmWpVHt2PQRw1S1WODZTGkpwBTpwzk0XT9AB
3senEMOW8mWkNhsiovBV2LTXIhofFlpKJ4s4thOw+S/Kj5qtao970FmvUWMx/oKi9kOO1maGqkhh
V5Bngl0kWfBxOHKB01SLybtgBF3XtVW+iYRgvTE+jAzqrEpKT3LrnQbREhclxzNK+3pKKVer20ro
uze4VJKEVv0v6QtJGTgV+ZJFCCFpu0bQu4zfMFFx9tLWz+HK0LN7BPK+sf5e3b0hkJThNUHc5haN
RFrLB06+f7XGJHrozmE5h+1M1X+YlSQww/MWEAP8LHjGkDomPnQ3lW3puHwiv09+1dZlLe3Lnidq
Fvq3XulutGEiqwPoUl40uTj/gmRHV4jpZCTayVXo2wFj3tKPZTugWa41kRhFJv707s7WVs7J9mx5
Q+KcBoET+/F6HpQ5JTeOkaWhb+JOeLY/kjnSFHf/HhdBSHzGWZ6wLm2UpoklGHi7UrtN/2ySyOIK
jhEuRgWWDysWTtkNi4OgXb5hzyAGTorG+KBEXEXIu7zF068jVf3hq+8E5o6Bzj84JM38+SiH7W0T
Y2DcYQTKJtc2chmwLsQ9sE0IG28dvmDLJc+VsthdftmoR6gS6RflGUX9Xf9nomCPud7+ULSJp9JT
aBQu39A7uBufMud2zU8CUD/CN5hsHeaLVeea2UXaWlvDMuPbkHsrZ7WSS4fqRjFyREVUQEEB+HMq
FPRZIAAxvUTDupoosY2NHbysedxVuHgjt0AGB1gOKx0MD5nntoN94YvTgeq7P5ofnwnUUQJr36dq
mGy+ssOFAnikMMdHsmD9vVuJ6Os23xByKPr30v4LhX/7w5/LeYVHdkD+sx6xbmSFdjsc9Q8nNvV5
N71GTxv1vBU8/RcMbjkeE87SQw92rGaBpkRIhUzkzXCa4sMeeLflNuEtEpZ4c3fvouCGlj3f/R+D
XbeFXO/NHQwmL6ZnDSUmqEdqDDbd71bq4EJvO2M9D/lrU70jacuUUSEeyU01z6tklNZmIZtsqFWW
f3+YNtnx9ubDk6XzVYm4s0JMX7yLjW3U/vvzVWUJLs4HKP5L7UZu/Y7TDVNj+PG90w+/fLB9+wK4
+L0pWK4OSthIAnKnzpyG8NwjamvtMle5n8OyYllNhOBnZpzNlZDrwL7SfwH/NVWdA7zkNH5DceNi
YFGarNkgHn9MFC2bK0747gjtvB/+Vo5lu4XIH6x9PK8whG5NFds+sYDVAj4l8rEKHh9nfaswsT1+
pnwraF7X6UfTQP7tzDdVAlfRV/AYY0ocxcz/TZJZh0vjlZ9d7qPwJSnkjb1gr+hA8u28aPSunHHL
ZnDfmXGtcnE66zYAbg3JRwYUG4K+rygds4AheqW6mTpOwkPuuIvJlnnUVZHUjeyDkrAhb86lSUwJ
wH0o39RvaWgj+zvqZC9y4gDucalGVvnIsM2navAsRVR2IWu3ND5XZn63tkeRrTAKjpZxycXxNBto
/P+0cDLfjAvO0hwx/8DIt6vkMZPRdqxMo+W7met2YxlJ+w+beJAwiVlNwLLKOVwwy6UKdreK9Nrh
AOdcNpUGb9MsrcK52pYKzqcCgJlPdZQJIoiJyjJXkjS8WOe18exWhI9YubSE5ipHriZZjiiNxvC4
m++AMAguh+sYKLHOEZRA01TU2C+sNuZ/3KHkYBSuhDQTKJxtLkpnfXfz0fIe/XkEcxKox3OvQ9Ai
kznHOffh/q0LIInwbiT95oYCWwQjo9d50FmzzbbL0sz9McPvvYFHxXdDG2BWKY2g+x1xF9qipiF2
vqNpW3TKspmcycQnkVQQL4WirinHeg2DL0TH5rIKFJ5SMUWaeRQukEi3ZymcERZ19qpAPFr4E6BT
SdUUmbhEErR0qQ+Y7AhMMv8njrFC3A6UrzvbG4MfuEwpcKkPz3SArqFxFHoCBeVAPcH7CLUc6rmf
lKXkSPPb1C55mnV0++PUhJMmhyvfsE5pe1+iH/3WPfF7pcTSq/OHjE5Kr5fbXHeG5Z6rh58IYIsB
tkigjsMMxx3Rk66Zl3Gs0nlM1gFIO4/LB/ndi5gvIIgGWsG+rY5CjCZnQiPfkn0gQ3RppcaxA2pF
0y/N9rM65zmK9hDBnhDx2M5dn9tlvm4wRbKjlek/jGMjdzUQWO8jUoWKzPV1ik/5JsTJSw6eRgIk
6GXYMXPI9x5FRtKl4zagNvW081c/UWziVx6CAJzhiQNARGAxYwCXqg+mTI5dVi7JgL0Do0SuDouk
5v3ockh1jLdyGHogoPBhSni7g06Y1bs2ApCIBnn5JpeT21GaQEsRRyDEvxgWHghj1HwQyi98aJOd
tsNvIkUr4zS9ts/nc3qWj3QQ217RO8sM1Ys/U6f8eMMHKA2SVEofexVhVx+CFvLbigoxB9ADt1gk
06tEKi31kTCB0oZzhveZOlqts0Te5wObXfgN6+1ILUn01c9ba1GlkvUJNggGluheevvzTBLMRBZz
TJTIzld1tIM9OJ50owb5dt3DLZJ/pgytbftKaUtwOaF/ur3G5b/qZmdkn0VenUOgCWCkZGXwtYyI
Ffdip+MFA4JUydtDFv44hXjEvZBW5Cwx4975d68ozRslHtEd0mDUclLsUNAwVoewcyXEBpgWfykb
HueNmKLdwWmlv/JdqaZXkupCxK9zLz1lwD+LP9ObG8v9G6hVsnCXJ8VSnpl21S3zGLDgnJFKFcd8
DZBSCEdIh5Zd3ZdEh3H862Riw2ggt5DwA5VHvOb+UpyrsBBbWeaobQouVft6EFAi8AxJg2JPeLrb
pAEmC3cXmwZ5a6dkE4heGatwdRbdss577R2QPDiYWXqGVREeDEWTldE23VFV8lH+g8m5QT1CYF+I
TVjAQtr1U5QRAj+C9zWlawgv1u1HEgvvn0da1tpFMlaVp1KnSHfHhvnXO6rJZKLspwzAoRfilE/1
UfYUaeVTUKfqNdqPBACUDid/U1FTqHCLKeYdjL9Ykc26mzWbQtkqXuAtS7O4XlOBioScAhLIAcP4
pmpPqR4QR0di7rvTgnwGPy1XgfaZOdq96T4MWWNfvBz6sqztRUZKT2Hc6TQWpXlTm5Qs/GVWLZ1N
nUO234UvkkDnBx9DgV4RQo7vo/B2zHg+0XqcVTc+G59nL+YGPIgB5vaMGVGUVMdTtz3ZxaIdLkNv
qwA/mhcIRcqP3rO1PiqmV1SE0cK9Z5kKsQxTJua6cXtJ9/hteeltNueApr+bh1LDm573CwA+sXKP
r1jCblbxrRziagqhVxB/5PuwsE8YDCa9hAvUk2wn20VjFZzgfgJRK3vBdXEGiUeqFClTyviU8HZS
iYIQl2N3qw7lErmjx+6SHx5mJZLRO1YQR5g94ve4BAg7zJoNSOPsPUeQY6kywyHhb5Znrr4wh2ul
4Ig4KYZwZpJcROH+2JxwLtSNRORCNcBeknPPrNK4puNWA1Oqv1L/QrUOU0q43kAwFBMUFgs0Tg3g
iXzgJfL29BG3o11h9YRmNlCuXdj0b/m9AWw4n0wuoFsKGCvJmYkAvvx+tn6N/nBvapipEOumjHkt
0qFPAetkN4bDlqCW/UVSaQDgXrzHrbrr0zY1w1Ia/noZyB9WJ/luyUbLgfcnfX8r4Pv3i9gmQLA0
RGMGRUtTajz6f7d2Yx7ocYWsYgIwTjSelyrjkqs8mFcFspQH0RgZztuOqFpTGe/RG/OrsKdE1CEQ
+a2aCLxQSMK8oI3ABvjGNX7cZhpBkJ+d8/WMhnHJFvARHTgMBAQHERg1WAQSeGK4Q3R2ZGbOGYiW
LgcuPeXBrBracmGZZhoaIeh5A6oQKgJScGOQwt01BivKmsOU+uphrElFOhd+3R1Qb+0TkrDOozGq
XsE/5fgyYOkOrA57Sbv5FWdErSF1lgHp7WKOpNcBFhf2s+QfnTwCx/DMETMqVd1sPHv70KV8q1Kd
YLEV6zIyIa7KBm9XDPYvybFtGT9XkHeR+OvYp/KCZh57BXQUMZJfhyRHDEnRGMR0pjGqdgyIGOah
3joAj1Gvkuc0YU71w+65o9U6twplf8snn1CAi7t72YbPV/OhSjyg04Y0U/sFJ4fxe33f7e7hxJBj
QHGiq0KkYjwOI9vpCeITFAvSLFPcxVoSuT8RItmMbqmwqdYLhZeWhrLBfmugRVNXSe3q++mYd/a+
mK94c10cHiTFEeTKhimZeXpfVClUTskKAjldeVUkYL6FT9sn1XQnQyjSjZz0dZFuf/sYpZ3j4WJ3
RHNiSiOJDzCM32Q9mkFM9zLL7S7SlMa75xWQhAExaXwA6W6ycFCUZXj4D1KJkusHxc8VjsXQ97W2
pe7LSjY70MXoa88pWOC0NW4DkihYfSta9yAFskBy27gQX+hvV3fFaasPUpZrXIfdsjWprPDpedzS
EjZyY9VfZnnlCoDGv7K0emapRk/VdpiIvr7N5yKReU40w+xhkq1FX2Ub79poOe5WwJnd0kt26cpY
HlW4B1yuCjD9q6TM+mOXFNBmDGAcU2y5NZ4NyUXZRggH/4kPMLo2rKVFkl+GqUhrqbSTwrJQohD+
ULk3pdzszOHQ5Uk/Rd2CZ4Yr3WMoAjsHUWBfoph37jNPymsEGSLs3W0KPDL3XVA6DbIuv7hRECXM
emyj/On0T5C2Bmg3m9Tsspcwd4CRI1Ybpa9S/LwgDWy5Ce4wh1YfTDLvmfgTvXigGPZdmWFw5KvV
nV9BzCvmFZ0wMhyGpz7DP4WNrfR7OoTkfXD7v+8ttdTkhReikgPTnrXPCmtBokpvakFw9rlu7WoO
dyNUaO6drS8XnDtzIsvr7E6sbe5QXz7y2w1/xWmUMyGVmYr2/xxMYUOLL103Tdhtfk6rNtDb/G7v
z7MZ7Ut3bhQtM9rgbX6UdLw+p7kBV7HNstSpMJNT1RbMitYrDy5Fbl+kRPE9s7alTzViVzec4IwE
uYY4dKhzKP0cmngJgLtktq21prxJCW2bYg7eGDejv8zgRo8lpQbvt0MjUelEYwAZ/PsgCn8YAK9I
Uj9sfU5XrJGinfUal5Yw30/TJvaKf9C7w47MZVZlkVLkTCxFhjE/JYgGCLGMer945rQfoRoql6HU
KpfhtaExggyRLscTY+y+NQq6S9aO8fjwrdMvGU1R1WS1e2yCOBGKhWUlZhhHJZf4uMZ8P1wwz81t
HwysL/BEFEItaQBXa7Xg3bFn/CdouYL9fn7+TPnSvjO3F9C43hD2K9IJXRQRGFxa/WFan5rrqZUk
d6Y3iFQk+l8ZIRj+NSqMBwWSQgKjzs66IG9hAcHpEEDBZyYCIPyraCG7FERBb29IpM/N05nX13MF
hd6cYJj9xT8/NbTwJeq9Vs3Wsw4TIMkfSfDegxQb9mq+t/ER7KztFsHdLNAsOP2Fj+yxOAFGxVGb
hBSovx7/Zuqr5hWEus0g81jLx7l6WsKI6lkoWM3dMnsi8XysfYlhd88tjoOf6/w6zfxbNADJ7eyR
YDOnsf6j+zq5l33uox8fFnB4ow3J08a3RnPOA530vp/u72SQe+R2NNMAxZE+vbl8EynjhFe0IIDf
o+I7M9ixkVyegW39ioWWgADEn70lxL78Pddc4P7YfSLqhdlJ+YH8rB7QygsOtwAb3I0Cwt+bHrpE
urja2Opj89hINFyI6hhn5N/9bIJYFyz36oOvFxH8yx7qoOR+PDyEvZzStfIEYZOfePf83FCWZZE6
C2udnTorMQUfEE4sdU6NPiM1PdVjNR7ghm/koaLuoYx/upL7z1Lm10tkqmn1zXgdHJFY4OOWbGCf
Nutm9WWBGZZ720Uzd/I9ZxFGh6y8A1bDmsx3+imkkKUpDcYz5bWOkVGclSsyhCj/R92UmpXMPn60
/JffaF/Fg7ATQQM7KaZZV/QGX7LSrCnnZ5leKru3/5Hx6angsJ9XLyF/ME6Yh6k1XYwfKLvOoR24
203Bcpo2DkI2VvkDXBfCfOeO+1YexC4Q3Nte+n0rgvmodwIZQkNnCRzBDMKGG9YQRPFPsnE3ZdBe
oA5FVaNU19s29nGmNcgkX5xWP+vLg+uv/PiNO+/hxOpFEbecU5Cmbzo3PhIN7S0/tOkEXcfNerpU
1ovHw5vArVJ7EG91m/DB99/8Et93fzG/UhUqfpJVoowtyuifDa5x7MNP5g87h7bhcRSz6dsoe67i
XEuK5t2opQ6VCJHnrwEW1W9N4Yf1ZotgecM+1MWyieeeiH/kuN1jTva5BvAWAfQzCFBz0q+RR16D
/gBl1DRj+fPfv5v5lpF4OCiTRJMDAUuJY/o0RdfP6uzimErGAgg0iDH77qXRBBeNAX45eq0p88gH
n4Sc0UPpiR/fRMqnLVgU1Q6XxW8Edx36v2TT5TCpf1RDK8uuMem2PGCR1n6p998S1LuQA6ZXdoAU
iTU3c9AQ9I1IA157oMX+mS+oxkO365EC+QAVWSGpAS+it0g5SJLkgpf5qC8mSYU8aXqngHIynv57
8Wc99lfBJIJxTv6ThxL8WKsBzeKVuIxVOX2b+yem1H/hD/6GnB4KM5+HQFbUL/W4vhqLELLompo2
wdjrHdTss7OcrHtLOVCXgKZ0pXdxsVcvTLsXohxDyfugHqMmy5sP4tcqSAaYaLq8Y24QE1aRLaiC
Jg0oG1osLvAtSEUDxJWklyXsC97lGCN/gHtXLn7k+BoFcMMHtIYjlWwoPsWirlwH14CfAZktRZxK
Ccp1EzjYby6tdsH8lXiAkJcTUFjM8QGV36pev+Kb7YrjD6vfoJMRfyQNj+SQvOT160xNB6QwDgkU
vkzvg3Y1b5jDrT4RoGjHYNTP/UPGr00G/nwc8eZebjlGGtFc5fiYHIfIJ6R/g1JI8qXwzAgUx5gH
yR758xasBez79jcyrhw0I1Ay57lQBm+XY5vKLI05Y4NCb6a6B7oIJ0P2DRC+Xi2eAZIk+3D8nWSa
a3c06lIQDDcsav1IHgAvjZF5jKJaouCbWQP0zkKnlD+w8DhlYtLREpMeGVJuIVAwDFNDDmUYCKzu
ohbxR5xgnO43xlrA3e35MMAPAO0tpBvfIaIiTL1+uIUuzAX8LjTYVWA6S4E2s9kJ/x3K1ooyuPdY
00Nn5DfRJgHqvK9KIyk4U4Q96rnxTHP7sF6aClyKLL3hNjF0GtbIVjTfjx4xBV0Y4ZkHU2GIWY6O
HY6lypJhcW/hbEXtNF6/RhOsQbV5bQuCgqnoWAVkzwJW5QXgy+aWMyBlZNRxd+Ey+YLOVV2CfUl0
SjRJDBXfbOTNoHSZPNVCSaPpe5Lrlae/znHlAC9JoBpM31nno/527BtDOHrt/04a2jzXwnQkAw4s
BpukuYxSAd75DQ5xnoY293bX55W0Y+T0fVEi2kFKUEmPaKaRZl6zVTMohXe324iuuuyCJgpDXtZJ
L42iwsQCxFNi9Vw3UlkQPTFNxFhD8SJQFEV+Hszihv1+HuftfNWmV+8FDOENyax91jiompYLP2Jh
H4Wpj8lLlw52BuMafPu0fCx8gIfDvmKkE5ylgVPAexsTKkPqXmFiyLWKOrv3fWvITuNjqXQIDgWZ
x88x+u2y3H81FOq85Ya2ssK/lCO3wFp/L8GJF3bpFDty1OB7paqT4Mo0AmXtj7ivEocQWLJxgAPH
fkJ1tZWgvJl2DAo47vcUGFTP82mtdz+UdYgg4ekso8bHGshWm4IGhLt0pKx44dWgILG9KIWxCrVx
3L227vci0W10JKOs/YdxHvLKjFO0VrsOHWDImj1g4JY0/3ZQPaCzg41bwj7BXDVTiT+gYHkYJrpR
qup9H2hJcvmPt3srAPMCtYcR5HW7KlN7dzsxd1VtYJyL4P2BGqVXtMznc/7Ttju3OLqPOLAWVwwS
SDwKL7QL5ETMPXLCmCgw9tFkRR8Kht16msGbk2GGFzoxDgi9CGFJ5wTz8kaxO64LVqA3DzHZK6RD
e4ddE8Jjz4r7Y+pYRuY1e3jk/uDbab5/UbRvLxEeToi29+nZT/q2sl3jVVxzFm3JiMHSBdfjwn8m
Qjlykts5qTPvqdOS1SHopi8rHpW3z4kJUNZXApJCzSwXOvcjx5gfcm7ANtpsMfmknRpQqiGcUfCJ
PMhDNJhMhzHfqcP0Wv72k8smnyvYyk+OGs5DDcwH0BirP3qK9W+4kWk3w5ZL1nrbHqqjShwc/yM1
X90Nmzt8gdJJ6S+Y5tjJSYm1cEn4Jxk0Xt4DBYWvjWPscqBMw6la4O5qt9jR8siqUiQ5HP8QO9yn
Sev/K9bjPSg2jRsbLhJGDdhG01IA6sZvQ5wDbYPaiRzprP2tE/FAX0Nur1+/Cl9K761x6O9GjZGg
kNj9fSZNE5sgOLc2yLjRODrvpp0na9qKb7g3Fy7N/q7q7q2Dl1oeLPzX8CsAf56SLs11oCdByi1x
s1BkqJZW4tkGQaamD0FgiErfI30EqzQF+apCN9xLKw1p6xBuh2GPeSeRg2ZmFnaHUVdKjijXdMqQ
UtQNNavMSADfy0nKQ8gOhSWaCef7VOWD+JEMLWUEA6QKZPVbVqnSX4VCSrQ9nZnzvmoRwDP2GrhD
djzE5If8QDgoSrQfLtOknl2xUacwl67WkpUrH4ab1UbOymYmFIqU8gjGcDlBYZRj8KEPNNdZ8DqD
KnsBWRYIWnlp9Tt32ty1nlkhQunv68fOGUTEaANjPlpAz8g2q26WD1mBD8G2nbkfXr/GngwNFdbI
ZlFr1zki4FimWE3sIiaUm++cPVsaZI6gDC0UofmYYfqmLucwbNQ29nZa3/N2cL0KbV9Jv3l7v9WR
uWod+9IdPMYeCL5bZyWsNCceFtXjpcWAU4T2rPBpyzBbq7FUcThShETny1sLp7t8C2Nfi3WDsRR/
/g+8KEy92QVSiPvtFOZedp2bCF8o4X/DBSiu9fDqYyYHILkc56ahNbhED08vcbpMxOigw+ZS4d6s
xdFT3V/1YB4lzYYPLn5jyTPUfN3No3K6IosqqhR3dBg2V8XPa79Iv8j75shxLU9jfH94U0KhSxnw
dEQQMFx7spUIeLunOpo8OGj7hWFpCG+mXJ3cTav0Chvh+0AXYLHqvZ8+4aMJNoN4QKe2xl3Mp4vo
H8dPTCfXITIDT5qb+l+wWYVV3IdjwLP1jUT/ubSM4/20qDFLsTc/LKRh4WD/SMSA0243OHW6HdXX
SbOJ5MI4JNWx4sHtE3UmNbTNmddI8vTSBN3Qf/m4d5e//Pu/kMNsCk4lkpyjDJDdFBPGy2zZ/QGK
RK0gjfHpWpwa1WD4S+UnHVyExTKuqvIvi1XrFqvJe8BfWCGehiV+NiOamywa8BaKnjpObheSx64b
1ansPTOa84ysC2FzjCptBIwG/T5zSMjwWiukWXW2MsJWPYNAgDnIRft6QWQpBmN4TWi9LkWnIRxY
HXWL8r49iB+Jly6B/w7/vA6B09JNxGi+g0sA5Uk0snpOCOV+38nI8Q8YWfv7UVfrrjtBXNBu22Wf
/71Rr0ycJIpCAv5k7ky3UY2WrDH/k18LuHkVzuYZCpgEdaU0ECkdIO+Pf817jCvKzfbd5+qTqTzC
OgOg0nMHZ5xJgaOgir2KJHp+BRYvj4GivskXBMi1gvW7Mhj8Blj94Wod5m702effKDMf+FlE+bYV
vBBjaiJum9b+t+4uNJwkpjmUf3QWvK9eN2ehSFQI1At4zGWgEbfCUvcTBVCy+B8mar7AgMEd8Sio
+hClPDQu56tgv7Cohov4AJ31hDz9cd7l7bdBYswTUJ+qUYpaW9VHXA/EjwVoxXSsAAe6B45LKAcO
heyepRqZDyCIa+1Z3QyrU0Iy5m8PK8/r7mt3N0ZC/WtoJROmQ7NfLeGQ2dmdcFWHrP/xIg+zbJho
9HJXWmDOjfZMtA8uKXy6bXD0yqUNvrbLAA0F5c3kh8/PSzObSsrxZbw1ywvBCq2jRVW/ivQlk9fj
LJfeLxOmis/Az5D92iEdLzkkm8v5uLLjSQrqgxBXUw8OJKcFfvYnxWzQeFPcMH94a8UJTXRe9bhq
4Kf2s5IPXjHkWZ27QDzuODV0HYqJ/0DtENi7zlcv7RMDxVo6jIdXwHI1C3a+sPfHba5jVwPbGJG7
a4aN+k31B9ESszA+IbSLV3SkwD3UqIjpWFSNSjX8H9Frtdhcp4lfwByJRccc67rQeMEkhdcxDwas
iGh/Ih1V2IKGrdBtbgJKmzgaBVp/terTRHsGKMhtDD3drT4by7NNvJ3xij/MjJqQNSwyL22wvsLP
AYBFgUn27rhMbLod0f9UtsAx/y8asm37xwxNCLqHXqwjdFtnFEkAHdGqjtNXYlEdn8yL3w1ctupf
DsvdvwFa1oVsXFJAZgwYx1L/306sWfqEHnYZnRHVOSY0yefO9vC/XtvwykEWdnlRXJwUQAKJzMT5
bt7NziHEu5q8F9prmwV/Epv+HT1i60O49eXC7IlH60pbIxSgfmn0pFB7msusI1pAOuNLHpPXA/X/
9XP+Y8UK+9kVxItWeEzGPWng7JwnLmqPa0kw+DkBrbMCrYFVpThSOfWIkoJ86B6ecXleGrwpCay0
JkUdADwsmxLShB74tcWcS5cj37TTMNPYlUXX4/tQm2hO9RTQzFy4QP1lpGh2R0M1cLdjyxfvNoIj
+1vBZ2L5S+f0zdCF2AKcn84iT9r3K192nKduQtJo7kwWk/DlX8EVQGjl5lpgyTr1Zzp6LdA9HWMO
CzbJBhAEZmP8NbyiM2cPGJcR6WNsA+6dkwHpNHnD/4HCkbejbFExfuH/o4KPlGDbxjos3kYIkqnU
smCFPeuUGMjLie40AjyVbBrVvT639sfR5Pt43ooT2cpyQX2vlPARqgeMAhhIDl5OTgPIL676B+qJ
eLda3/Npyvzzr27HFHk+FmkSay/B2AATCoQOdz3IZ3vHLgCerIil8RTzILg/xn7ef0Ow7KXTXIZE
okoi42F1SkFEZeo3fzoHgjz4pI4hxh2V0Xzwn5Ut97J0kI/x6tOul+gkIqaLJUMV0wYhAwo+LtbN
yRKNAQd2nMFWi9gF08dBuVdOjh/oWDaBMC+9Lua+PWwYIdDFQgmvuqBF8ec5R6flvG1J4VCVLr1E
CQbmbWBTc6xfv7c31eWfVDpUTI+uFDwjJbUSpJkgXZvX3etOjGAQfcnCABkpFJObOU9jfQ+1hzWh
WHhAN8blWuHwsbCC3VR77QcNuL4OG1L/7cOnnCBDsSRdEemwTGw0urdknrhu4UFWW73VpMSa43EG
vGo4iRkNVutF9H2IVka34xuSV8bh4qGBI7OmyhZKLqDnZ8RLtIPVs3QHYytorSIfcdhPMOcesO9V
Otx3Cm8DE0LtHvkZc5zKU49mr+qQ64TVXkzXv5MXBWyCCI+wj2ljAQD9QL5zFex2hHscnZWECaSp
nB5185Lg+5r8A0gJVZFsBvlML1OBLWEBuItTrgTTD2n73RrTcf8vlqaBtT/hbCD2IK4VQ6/xuXyH
rb9In74ihGb2ckb6qmnV4t8civqEGuaIEuT3oSScdNknnGcSkpPjR7xo6m8Jw2CQTw6uyMomBiSv
OTVcTOloceo6iyAP7QfHIp0/RDL4qLw6HvPL2OcArR0sg81eluD5lDpbtqhXt0gvWIfKSLvT9hgf
mfNUcxp7NdH5MgUjkX1hJFO4ujA3wptry9h/hVmlRhOnD5detJmqa0kbQpE2ND7W23eApdpwcQws
UCTg/7MaLkIFPY8j+J079K7wk7ZkuRo4GLjTncHB1vE5v/w3/PmTRLg8MaGL2N31zi2+cjOHm7Zu
RKBR02wMqgS2cxTwIbL1d/sN7I/HoKg0eTarOUQM5EQ1aN3fRoWdxjXoC7vTY2DgsWBs+jbjYwMp
vQlKXHjgNp6LSUirv6hf4zjDjfXgVRPX/ClvjpVcjXTifVMTO+nYRrASSOLZCpAmlNQbSSclPtfy
Nr1tohI6c8VwUAPQviATc/peoOdAq0T9yfrz/tNVcaDYlSazSQDWCOF2Q1QH4SqYSdCzRBUb9B+H
1MnPYVIX+48o8KORNFnwZ0RWgDES81kBgE7myteaz7+l8AgkN/XTflZCRgdUznp8Hn8Hb/TvDSZZ
U42j2JN8/QP06Iccg+//60RT8fpDTKpBQsr5B3bAOx5Fq+piDLUgpF3UlheARW8j9g/dIqcjHyDh
OTvpYtAqVv082L5nmduQFmuOIFBkaomw95ln1kpDhduG8HzOmgJpCEklFO1gWXWimN3CeuQkLweu
56cDwoCPKC511Mk1+hpICftcBhuyCR83ZSWjlQuLsvv14hLYRG8AWFHrQq6jWxG20iSw03xb5lMG
cr2bHtXbpVK3z7k21j/gIGYypiC996FywKSbp0gXf3/30K5Yv6t6ne+UHO/2mvz6LzJTH0zJS6Ku
d8RD/YPtmb8P+Oe5FP8iULsASm5Ck7npJF173oS/eXw8f1Hm0ibMSPv+cTTs6rpnVQs8x/DcweMP
sesBbGI6AEFd0tkdKrMDkvnRdJ21zXK7JujH1kdB+PAggaTuI8O39HTApV97/tCawnyRXvrZeVb1
k8Qc/2xjaoP3NWyqn2Z/jIpXK83s0q8L/WVb7MRhsBP5wlnmBqB5Ro/1i37yzHTG+hosxoMc76Po
CE+3IrVV3e0KJc0QIlacM8jwBSUyTkc1OsN52Ne0ytt+lYPFMh/OdYZu65skgzjEXWd8mGvOFN7Z
lXJPmZnpDZYCdF1iXxqulSuZJfavrSTC5hfYHAFliIKqOIbv/ewHZhXOI1m58Z8tp15vhpi5rfN0
LuMYCkpQS2KNAnQkVYHDrCATi2lOMGNv+UL7UUKpS7ziuSjoLTR94KvuxNS6KHxiSmBltL1mddpz
xvdhcs4SNH8AqwO8PyDJZJjq/Zf7mSDoEWlT0A3+q0oUfcwBjxpzExhelJmDGO+pxHixyRAlAC+4
9vlmgCoSBeRxl2HPHdOg4WvtNs/CmhB/UhfpS2uPVp7KrZ1SAyzaI7EmmKNkN/qBaxuEd/BfzIEE
eTrm65ild6goNObh/aSzokKZ0ejDjkrFyBXrStcjTDFA/g2X/FYCbRgZMJfyAA3l21pwC05SyVpM
KWf/FXfRl1r4SdLP1GigK95MfKgWtJ3CAS5J0pOJajBR9Ohe7IBPr/WW4QXJRkt0eX37hpwASLPZ
S3Uu4wcSH0Uh1pZU04od/S/i3clb1Nxp+pfuw8FHFk91/H1yGaxhWupwA1AXNkL8PD4unljFbTyc
HJAGhN4z4nwMLK7bVSiN0CIfkHQmcxzAlhaa2at0CNvFC8eU8IMhLhJwwMBKyMnKcN22WW1AQed7
uouKClpSWGEyUZbQ1PaVKyLmmtQ79X6oDAhZdkyCS2SD5QqiHdycWlltYS8RvwdkN0U2Ry1znwMK
773uCgtoCa3V93SCDhi0BKNBZ87sPmtXa5fQWMeBv4njFuVt/3i9LY7DfPq6AtBI2ceAfa7dZCVO
UuBul1EKWB0x+tBVXqg7rNmV0BVo4klSLY5BgIJgae7tdBOIwjtl/rGJ4Xix5/6iFmjTAbyNzwBR
eZvX0SCAXrtN/GOS1BUmB3SOzdvTi9oqI9glWwWU3yepi4RanUam/ixZsvdswtsNv88wVVB7p/fz
oYp6Qj2OvKHIf0ZUS2MNGUiDD3eKcJbAGi8a7uPgwSa7vg5vy97OzzbbFEJ9L3t6MKmpyU2wbywB
T9gqwre1OTP3G+Zl3E1EuGGdZ8lX+Ru0h1RGVX3DeKRi/D7+hT1qDsYRhsv+pXMwzmR60vhrfoIU
82lgK5U6R+IY+O48FHISANxXPtL5bqF2FiopZvZPrDK4NhViOWhnXeGUhQhYckixVhYeHLi8QiYf
tV0XMQzsn0cWrwE+bCtRFf56wqmXegqsFOM46deRMH914F9WU+5gd1a8BderGUYHAfsdGSgW5zmi
w4iB1RD1kvAakqtcnUpzK2gBGRIXErQPYr4sH30F2Q7gXmTJ4Q5xymvu7jJGQwpm54th6MWVJYXJ
m+uWS2gu7Gcdi8lLDAI3NmucCub4ohIpZQhge3xEJNSFi5oOgIT/X6nBpck4P5+UPwSQEWbfANwq
iBJ/tcnWQaJL4c912PNP/D5HAzgOE0lPkyaMiya2cgwEW/whFbfABVne4KgHpBkqygh44mhn5skM
SCq6tJuAemo99XGLWN8PAo4wHW5Va9GNjtyPTU3iaEzK+MTcYI0HmdHce7BKvTsKfF+m7Ryxm8rV
w5vbwQMC55fRN9Mc5v2IhCO7XaOaklT5SfjNaVMv7ogR6kbEYJav7FwAXCBidw19uZbLt/tuLYDN
FpuDqYlZ2V73uE2EWhNn9BOvvAwvuB6FfVgjZEhCgp5Pq4d0+5I5xeQK9s19AtNgfhui3ep3TqXB
X8bXxp0QhN2MxWzLPjF/FpOVbKFZmDttAAiP1jqrCuj5RvPdnpqZOR3KOa2XskEg8N0f38HkdQpI
WCcOFXlddSiKu/0jvW3O/uhWW9nMg4QkzwmkxeStJjn6Eq4Ui03kFpQvyqoMum/ytrmNOvHOIX4G
uX7C0yfusyrJA6fGffA++of36+gg3Jiw3LeYLt+HngjQvzxCAwZ6v00LdnCtNrBZWp+2N+4GcvRX
5ewux269cJF4SmKMbsMdyKByuToRm2IrzB67oqzKhOMigEnNBLLeAwjIeLr5cazX9h3HqHcMR/yi
4Qh6o+BDFijAhBopsz6yDgFe7hmStgtyX97V/dAE7Uh/uQrd5gDF/wpMhrrdcTZYuxPhLVoFj8KS
UEQolQ9VjDgviVBok6M19hFrvM54kWdnQo0vaEovySMPCN5LknkeDFaMMUgNXyUdIKF70OEIsZ22
cT+/j3QunmN64RNPnyaogMTZf+JI2OyZLNIYw4mh+j0FRrGkwMiN3pVeCbRa/FaVqf9+BHaL1Yr2
auRh0xtr/izX7YMnFn8h3kZQT9+YKW1Bhi5iIRqBiJJY71zV4CjAnWYHcZm78lI0UL0O9diIauPq
6MVv/e1O4/AhAEdFHUfa1C3ZeMY3va/7fCKRcw4eJEQg9NfSkdkwhDMqzRGg+GU5r5tAAeqAaCg1
hqmStlPHW1xZdCyeGSiD8bF/jRz4v/WPSt2GYpFBQVku9+36Kdxx33sd4SvDM7m2oHY8Nizm2dx4
5XZurTuQ629/cK+G40aUftB/NBN8r4YZ0K3/h2oFDWWUyhshQSYlILRd8dwOAHTWPtpEqmxEUS/m
r1ZkVKtjho3e+vyA5unzqVlTmcQf12NF8WI8o/NGsDxxliC5EN2XIEmBneS4xPzYKWn0bWOQzs8U
EZZYVJ1JYOT4RFY3BJk4NDEC8xW9HjeDV4IiipP0VIiyS0UCQ8NR+WnS+M2RPPfGQsx+nLXIR7wO
IIeNqKXdTz+AQmRQiRJ2php6RITQczmM7iDz9jDV+tSMveTJ401vodXSJoj1kqGBRFVdqf3ufYSp
xv7vP4+pWqDqxAebZrFxWGmzvSDmXGBLcq8j5eBy0C/Uz1bObloeKt5qji6b29PtwfFuuiPj/1Md
qvDFJjbM2ehcrRascHFSnI6mlHB5NVEWZ+lPLqU338T1Z40CHdHoNlK8Tp4TPXhPf1sHmjecKjId
mY0zMx9hW3fWgo65tpo18kqAWSpFBFiAN9Y7FjQzZbkQJcG94QQNO7PgGC4rEt4/SvViUxTxsCM7
cW6c/tKnO9sVvpIPG9DDf/wra2yMSH+7v4O5XSEFQSOV6uC2ofJyd41M7NiZZuW4tmyfHQcs5qLx
zcPhjn2i3yhnxlnDyMvumpVosyL9d5oWIHUsWDEsB3Jpg8HktYGENCu51rinXIMG8SJPdULUuUuu
5VdcBB/IGtUyZLYwL4IFEVX6x//lCm9ZSGXaFFAf2iDuM4+mRMnD3gqAAtqBsHDgzgIRjyhKevu8
TwsNxAEyDpviiw5+vt51rcslsUz90Fq7saxje61yBzcnrBbpdsXgn0rl/4ptW8UkIn63oszUJDk3
TAd4EOhYrylmv3ruu5Ni18nlSCjGq99Mxa3iv/IoDw2YWPFo2+v27lPgYrdvdKgNkELKSDa4fFTK
h3lydhn3PeZoenyyxb1Ymw+MFL95aQMoGbOvvZjN4cMh5yaT7JsaTiYMxsG3OkkB3hROpcXInjVx
H3xbkTk1LvdAwyT0ZOVqXl8bUKnBDw28GMBKMcUfF3ZobU6LWKcyUrVH0ZEOPx61mNY6sC8kXp6s
zjmaZT/dTeXDdqDvyiyR/ng0IFf3uH7KHxPQSiuDhcKhGfNsJ0BaOcnsL9jqBf4zfyNu89gRF7p5
+wbqoELZxnkb/4e0gcTnDK/gGf8PGI/NTHu3pf2O5VXbEQ3o5guxWj5zSVPOcIYQoPfkVydAwjw4
iaV9mKNi7KUw7on/1yaNaoqNuBRCcE+UwFv+JYxG5a5S/UM5Z3z4MmpwfbzjGi/XB0jmBx/Av+ZO
nY4jWiz3Ri5QY4wpwvM7gqdAAuCs6irovuZ6ETBocTvxWYAMLwvnVI3MVVaEAfG4mhh2dq7uo0cc
LvYBvBlCmrK+mbHcfHkZ/9j3aozZo9NPGdIMkLWsIDlf1NZQBJZ4e6yIdYRQsleGRSPclyp9FGXC
+yh11rAKPpMEAcCUDmUtxgt7Z7BqbQhB/oWlp5x2sblaHR5i7Yldms4WHSTesl4grcxiXbIA+yCm
0IMQniU4cxPu+2Lecnglvo/FQ03P2ReVAJHyaqc5Upri7xOyP/OqGrECgG/zert6goYr14iuzcpt
IiLKRUOPT0cx+9g25Djo/aFTFbnksH9VX8dt4QZG9pBIasKfXQiG/Vvq7+pNRKIIbEkdE+u8rijL
qAp7o4xd5A2mPFaUaTmnTbhgG+r5RjtBt39V7T9jhcabdAp2S3W3+DitSaVpXx5F1SVuia1PBvT4
40MxdEL/h1H9vuz6dMTXEDnfO5XWEsERsfQvY54vGA4Ma9xafDiCUExngR9e9k4I7r/JRx7UREXH
aD/HKWXunVZfo8NwBh4BdEJz9ubte141MgGEeDU8QOodySmVaN0TxAIPVX4YmwQSDDLBp1XCFQbl
jUMfWeAs+4ZDptIhA4NGCjZOmGCKRul/YjP/t4XRdP5dSabqMLx2H/l/63ZS9BtkpzP/yQ/c6teh
vzfUhCPMdUCHzJzuVrszVNoRmQzc5RQJoHwc5e36Eu6mUT23C7sYL8yBhozzTYERUqwU6McAG10c
a3FuUsWkIltAWVH8puE+gM3TdGXOMD+aNj3qseCzHpzq5WhqrbeZmVSJWd7j9LOjZ3xwdMNefHPS
1kk6Re0Zu9gfXf9Kq3uFBLD4cAmm2hZI1y2yGa/8chh1JJf6tf3+EGcF3MGmnzBV3DeEa4t+zMQz
ezn/V9QXiUxl7+C/8aYOuuUvJzXXcFzhlXaJOuxVe1NqxRsMfkEO50dIj4pm3t26P3hK/5P5Xk6A
opkbVH7iHrf6GF773tEU6G29j41PSXLnGfhqh/YJ3t5j+eadWhHXKAB4F283Fbzi2Z1FqFvMTvvr
10RPJcNwfUO9QI54fYJX7jRSZ8esG0lHdUlnqfkbmla9nFMxuyy81FcC5FzjdAu0OL7ZtawWC8En
tbgVhVFgZAwWioX/bohPVgPWZPLx7G1mjRsaYMR8ABRiqh3WlYx0HGAjy0jcBzIG/ouAwe+o91gi
iPcEMJa4QaIW+MjTPFEUwqBiuX5bwzLKZ5N0jGW5LdH+A/qSACS7BvY3VHDpvQOP3l1VPTXMH0vh
n17te6xLLTUo2yZ89jxN3kg/umLGvvj2XFq/WO8jXBcbyChphpFGNd1gQEZhkdbZBk6rl5o2I5Kb
/aq51gFCxuFtY7r4axkHcbI+Ol3Z4CyEgyY6OQMJZTxRKyTdClKQUkI/vW9ry/i70TSPi7BED8J9
rUmN2MMWhhNdAwfbsaD/UImfxhxzlioHJkjPz3n7AwOUtdPCrqeWFQDLWNhMVXCdNLDD6setqDZF
H7tFAQ7Tct/mIURdI4NE+TvXZw334Qk3CZfWUwQ19DZBCdoCVT7AeBucaUcmRAq1zj+WNj6aN2qk
J0GSUMTWNhHFB8Or79nya8thTQmvZozs5WVw0hu3B8CSU/LzqtOgBJOlYYmMKZqIYr9IJo9FJacI
wV88oZENrXqDZazaxWp6H5S0jEySsfF2WnI6NGUTbTz5NjUnruUrtdxzy/sloZ8OtlEZXU4R324G
SLsRCWsnvi9MssCRZ85ZS+hEtFeqGsMHL/sb700zVkaINojT0jfZFM0pGd0dn4hyuRBU5TbBkPkT
NaiW4/ILnGfdC6nyXL2dy4vcv7qhZvV9IcWzEbc8Div3mgOyjPXuJtuYs5H7N3GxsWE9v7be113R
9yg2cpb6tlM3nUd1NI71VDLFwwABge64/t8CD3C4GjaQuqiqqL7FYxR/1V+fRF41p5rBBuosKfmi
9MJHGpEAZGbUDrir/K5tbd9P/xTh+SJo2hdoW1W0wr7u7YgeRHfFN5H5Y/Gy4X6+tXVZ+2BNhcO5
zh+swblC5ty/aPP7HITSY4Q6FZ/R1a7m2pyM02NGvfsUD8zcXhPuubMvHnMWet/RVKyeLfSztV0r
ACoQtH9gJzS/L6SinXBDkXbZLG6oTG9OJZGfIyIKB78G0kgGZpvDCHXfLxCy3F3dwcewi3ZZvxMa
CEHT5WrCy8piyzglPemRW+LpcMjxqtsyGnrExhB+AO2+Pu4ZtTEdQxQU5dPkFzSeFLRxWiF/Y13/
A4MAHasYEKc9ne+SELFPxm+2Yi6PggpBeqpbu/0oltPBZ+BoDekpVeRxZHb+Tb0KM6ylcmHCVNb4
k4nbw9no5SkIE+rOrubuULa5wzS7mZF3yszyKBcsAM2asVqUJuaowt9cq6YgoorXd16i8ZweiE4V
tqlvghu9bjG8M7OpJf8pIflITUhA3Bo0Ush7jfvE05a+Hwgaw+yycSy4KCbxxEfOdgx0cuuvqrCE
TVdXn81Kszqeo9tDOfjRNNtiyCcPJxrZAHkE524oV26vuHgbel8uLlTUs5rrrh4QAzYDTZzRALr6
rXF84T+T/fxBnBx52z3KgyOGrSgWAOrkPdTPtbM2OEii6Y5l4W2KaPNPb3XVxZJ3UWlfTmJjeUG/
qTzsNc9qSaANQe/x0N5wifjwinNns5H6G+M3EcmoaIk8dgpiUtipY0RNrOg+X4wxGEigE9NmEMsm
pL7s2vNhkJjABrM72TuRhae/SSDxiFL+mxsksUBHfzK4wecZ/hDI+ULUs0RWTJO8xAHD8c23w5WC
hFRHIbpFAOdbYH0MI2/a8cdXv7Ys1l2JRu/R+lbQhyftBzQraz3p1MvjrLNUH03OAjW/inzxhTxq
2f9g+b9h+X1ZTbm0sgpMNPuMJ8kpK/r7xXbo8th/h8Xzdm0115xlLyrcB0O28D1ReczFiWXcqc9I
TWyGCnlu/3tZQEsOPfqQrbhlEQGHKieoXZ8tPDS4/2K0QufENHPTvkhuY/9nksPMRIXpkvZdClRP
+kO0j5MJ5izfXAx6a6d/Yy6o3plomH2okez+IWHfdBWVqDIsSl29Ph0GPJvAlpp6N98dVBQ7aU0u
nSjALPVYeM+VZhZ4ZwcYvLQeVP2JfWnhm+KLfSZJi2yCePFldnwZhevAHptRpbb7mPzJIhRdTJ8q
o5JOJrrtYA6XxP+1u+Ha1e6C2twD8fSJEXxPSeIpLzvYhNg73Q68kwf+6FsKSTDNQl8ctD4q9baX
B3V+apVcAL4kRgi0lns135pJBxvqtgo9h4rXPtRN57SrBdBzBHWu1xCkxUQLy8cFNwjAtg5xPmMi
jzkFhOzn1uyf8JsVVoN0dX1oG/hWzFc2bcpeue/bCU2W26mKwi6GuuH6VeTeXNwd8esV2BY1F6LT
gsUom/9OWFNEMrh43ek3iIhmwA3q7JDKxYRhXf+XjTGjTVY47y34ZF4QmWKmzgabbunEbSf1RVGr
cxcWdEJQiVT77l5a/lrdTOVQdoihvfX5LxrETei991NJdOUhWCxt7vJOqMmu5RiBtkwga8rXswAC
dAzAzHhSXD+ZlvqkA0smoJBz2gInlI5635Dlrn1hvyfBJH1DmKC/llmjwOz17ng0d9XE+Sn3OHfR
w+KoET0Hh+JDYqfqFQERbVM/5lxNZ1TBBlX542VzS0OEyKYGSwaDokH7EEaazkbLQsx0pWWgTlwF
g+4TRAl+cwHAWZQhOWzO/w2y+H9/3vprxyNp/QkCPDSPvrdmwEuRnRpYmGUfcv9edxbEKqtFUmL4
axElYi8B/8CG5y4hRAhvFplkAPI74C60qpIFSGfIg0S7h6Svk7ZWzo6ZiFfABcnvlNshXUt3sua+
9o6ydogZK5ZiFk5n1iJtvZpaNMcs8iQh46ZGptFI4tIqSHMUcD+WermY/+EV0OGv7I7cFWJzuWNx
U5TC3BUwdxLqdv+FFrzVyblGIhJmeB31A0xMFipPqUzB5BdjrqKaIDzipkH1HaUwKn4Qay7cgvmT
eoYYO7dgemh/tAqCjUeLfmW5l9lTRFRrXZgOe2PxmY6N7ppiBkyEBJAl/XN+kEFcDuE4FdHPclT+
/LkdYs4tsTJwjE7kWrcTP/btgl0mo9wai75/PvK6STDUpOFMIMGFLfvIarShQVLnd6JSbHFVpP1A
JaRBKFKlUOuh9twcmpnyCgoG2Kc7bAFVOb9vD9N/ivhsGiW1Rt1cBIvegaavA/VkBqTRgqb5RaRK
/HFTMAhzn7+WLMFUQMxjbvsD64n4qmwCRf/SfPnAzC8LAFUtNBA+YHtd2re+2bifqiEGWI8YItIM
ApQgVQQLm1ICdl1OBWl9+3L1WP3iXwvY2fCQYcH+2I/MhjY+1xTZSzqoinkuym3+SqMXAqzzbo94
QedbQ1x0lFvUwoBc4GqPDBPpk+FTq3nFeH8mvPTy6lHnjzUnNI/lH3c15hmZK6/MSKjrvpNO6xBu
PgaYRpvEI8mkYcx6ZKexzjKAW74lruIb5CxhRVuFPPfpE/NLXWfNbudilnTrlsS8jOl4RLeH3UDB
f/TSCnDgzkeAYOqawfcdH0Gae2kx8oo1t8ZVVVb4Vk9EcnzYmm85Jfc0bRZNi/HoUFOsjk11Arnc
16jXEFgR1LHLPC0nS38tqIWoteBG+HNFNNm6YfvQ15yh0+fXNZOPHp6ct+sHpdLDp6PYKm206wRe
tWC1Ea2CJD4few/nH6KOov8GZgFwZ7E6ebTnT16VpXi+VZH6XJ2XdDItbjRP/YPeTTGd2tJEEMpa
cdgxiRkjlvjCsWE/1FXYFh2/Zn8iEhsCEwEWoIeDoVOwAdJhvkw7LCUUQCwfYFiixKW9yFeFc77s
varOPt7qhIDHUupZBhLeQ4NeVxiV1JFFbWNUP1vINGFYsaqs7H4Rswtg4u60Ed8U5HbCIOkwgLBl
0akAdnIt8S0thZy1zMKo6KJ9X5FEQKfjlpWlBRTdMp5osI+SJwKcioURnEq/JL+YgCk2LjouzJ4q
lFFQ5vNjZHjQogv0Yn+yjNjXUc7bB//Jrdi4NsNJWgYbV03GgWHCqMlP/viE2RNy20iYDMmfJO8X
E1df9BnvnhAzersd+XdQGq+i6OHr2n02hYuSPdmTI0KykcgzNMJnE01ok+1zhKqRv/7C9qQ6SxW6
6DB3b/pGY5feOVE9ZxcywlwNSTd1e+nGcAfBTIXXPYOy0XC3zBqnR2bxDJVM6f25qmyDd+2nmLUn
Q4tGRmSr5vFLsZd2fxAqMEoKitjEs3O8xi2Y3GWOTFAi1wLEC/8Qyd8U1F6X5Ispf/K8uz1GUfJF
gpgGeyMDhIXCSu1m3JXF31t0WkJAXmNBeOQtwFrBmPpyJqck1kQzaBl+svoGpcYlSoDNojJChEDC
20lZVGgHKZEE5tH1lL4LufeSvfRvZv7jdtOMk5wh2h9yFDWtiTpdICE5UCNapKLOXLgv9CrMj5fx
nNMe0PHSzN3eRcFTArEfRZC84iUw6WAVv0ZXif04j3h2msQpJtYXtf0r0h0uwpg0+eiUNG5C+Otw
jZVtjosVnRW/0mJ2CDdNkKcszBKlnZ3pvBu4x/4//GnWXamxw8dnJORGnMOWcAIc64QfBjmUa2Xw
JPqYcC2ZWYUCE+r2hIhMAEIOc+eQGpDFNJTdVdzjMuopqtkYA+cwAnquuhJ+HO+exIyqKjWnfmkz
qCGt7eXLnuaJWwH0I1zLrb/tMu2W15EIcgm8oJA4SnUXoQeqpO8+NAceSUjnNE2i3rZxztIQvIbK
ImKCP41JAT4mWAnHOpIldOs4n96OVuwHGQbayS0f8gfLvHbgjlo4CKALxrH1JuPBtFGW63CYQ5kL
oQlquKYn2lZfhvI72b5ddEBx5bB/ZfATtI72cOz+ZoSEzVC8saGq9Ky5d4Py7+4e+ihHvhuK66QZ
FBQ1wxo+KKisaEyh/RKqmzDqqkN3zYKcIKFzmGUupBvK8Gdku9oQZu1Ec+Q3xMzaGfoQErYI25JE
Acte/tCv0vwr75o27VlAn7FRBJ7NM3EgvCjhRI5pt+TlYDL5rX8ctIJIXTdFHPHJ0j6SyZT4zlBV
ZCaLfdk9rt3mH+feAxnD/VQsen7JhDU5E+mLsYQh6kb0FqbcdbPqpq5SV0XbN7VPZuHymYl3dZZT
yCpEchXOzZBsS0DeEVpqxBQwR0P9TrnlTlBH4jT89Qe0t6PTW4Gk5dAmx1tMSvYgkMsCA1ZwU4De
8wzMcNjcI3uzKag57nWJO7eQnH7CnosWNGOKQJ21P+kLwcoR+VqmRq1RFvHqDj1xWWZD8tQMvctF
JWZWEXCpP2Qmv09rQHB0OTSVkDyWOk+O6CvReGzPKG/tuaHAYsMgzeSFlAgitdOXulVyMvjcTsjJ
ARSCNJXUiAmvsdenHs59OS6gpsnJM9TuadEsPk0nslMYcBi+HWfne76awC1/pmG0pCXOVWjH3ifN
HQSqyoOumpnH1//e01OraiILLt2XA20/R9CDcPSNyiJWKFgTJNDOUSEobg4mLU/Wer5TpcdoCGQR
Zii3Fp+rH9Z5DuBz0Pi9Zob/qlnoYWrkTAPBwf/BG8lOJhcDwbZE8IcIswxyb0vZeFQ6xbun5Pxw
egXOQ9q3JAPKJdrHtJnyWdYj7uxhI03uyL0k2QzuPgE8zQyACb1PJk6XaUF5v2FrNUNlrFJ5Iw5J
+a1vIGJh9YrJYsSBAQofMKtUjJyAmcpC1fW5rfngshb1dPKBfj06gVGSpn+WVKRhCxfrEpOtEA7q
zxaxTk3k8QdcxQ9m7HqcZ6MQqcRLxji25DukoYKec7eVOOwSgrEtMdO8Sjm74aNqYY3Z5pHd4L8Y
5I9/R4P6HLjavZ7b6lg4RIxuUXHk4H2MeuP546v3P0VG3AFynV3NAsJ33DR1Tb+RM3LKADBypXwi
S8BkS7AHkWxByyBfpoqMgJGkaqwPgOX+XHmCWnEc9PsJuhX+HSroUICCpWVXayjy6EV/FhEJOtJk
sdnErQ6pl8i68o5QeSW2+V3G0pF2QqGLvYKvPuD36gQlBkWbe6DgaLiQEfSg86kBgkjyfJBcemXz
nsUBmK1nBhD6LdvOfSJ488IVaf43JryTDph+4rnyXcxdO00qVzBlFKzu9NTkuC6P0V9qBmWsx+Eb
i0SlW2JpGsUbQruhzHeyO0vdm9KVbtBH6vJuQ5kVQhvgW0L+9wIRr15kRrNVcbwaJgA9fqNwNIzE
E7XPLIGjmx29pt0QT9Q1teYK4oGBEx/ZGyVDwYbXgZzuV6q+R/9+/bHqeGa5R8zPdbiIY5Zs/BrC
dI7iFJdeHOD2fgoiAzMtzoe25eTJy3/SBNa2JLgW6/B60DLyFh5vMYz3I3KJzy87ppK1SQqi+csB
WcvbdvZp0KZ8SxgsWDhPA0xcL9YHKCOon4GGawiorU/3w/XGwl1Mf2JdPx59lfx43Rb2sJtreN/t
Vt9sWdQRrJ5TYEcu4hFQY96DYJNhzrmePHidqz4HtTwXnGOo9syHmkDzfcW+IX9XC9sTIAxTz6lF
DcAuFS1H06/KIeoXhjBhmev9zVHyFUO9COKXcRMYHLbCUXNxcpP51pYZu6em9dT8Pqgq9JnpdhFw
EVvCKbzB2ZMRowHLswb3B+3/WDR7mP72zXHHWV0lGHGxOTLGQFTEh7PwWC4Exayi3kW+lrjrk2pj
NXOx25hQ/AqoRmLLx/OpwvZeyWVYJ0F7uHMUGxiM6K3DnbGonjqlWuELBiuTy0/618N8GPsZFT7w
J6xXSqi0kbi/B+t+M1Sk/aTaALDqh+51Vt+dwsIaD0wtCv3010F3juU2SRMmCLeG2+0Qrq2dfyqy
FaW/hLa6q8yKmI7lVOnxZFGVBGBeUKx2AQdqKl6EGAUsuAp7JV2tCZ9Zx2YAAl4mt2zrjwI+9Z0+
bxx/p5H99uqgr+Njl95usjEIDMXWe4DUDnANUyjFKmD6MWSgo/8iXRL0jiv+aT/oO8kI6cGVUu2V
4zVrnkeCGYC3ECLcovhUoNrzprql/afgnD7LCyWZwYT3sz9bTvmRHbjpsDwlwL77pW153ZrK9Tox
HS8+GEXDVChEn1EQ9TWH0W5hT+UQZzeR5XTDrkuTxw/SzCgjnjO7j6Vu06O0TU70H/j74Y8yT9e9
jtW6IwkptIvAVpRnaCQP3byrfOXsIkQhQH/lo9B/xolwoorYlWt0SXVns7i3mdbZd5tUBZw9pmq3
1rrRxF6c7D8zdCv8P0lmfXr/FVhrskECOABQ2b8g0aHXtpz7FuEjSjcnSbLdAcUUvuW3s4Dam/Hq
jOHMOrAs20sZXZrAf5H4ezSzXAmk4DuRuC6evy5o6bXlhNgrSHvaNKUAuDyJ8wP8OWAWdwO0J5YU
k4I7Lgpq4AequyRHXUgfIIUMXcqEADkxNSG30/wBz2ddfzLw60Rett9WUYnmAng+URZ65b5usu2e
t+JGX+AIZQJB+OLbObmWJRcTC9LWZvcaSAqj+Kh8eciqFaSlAo/0WCMw+dALIjimy9DJLFisIic3
5LrbFdLdDKykoM2xisYf97g86iIZv3zKsPREnervTZ+Z1MinJ4680wDMbb7TqlwVcGorF3dhE5JQ
aoqrrrJWT2E27a2ILUYbaSU6FjHyUF0cBymEsBBpHNLFRR9OUV6RVsZG0w4bRUWkzHmiW58cOudm
g/ezL3r5NLSv7PelgnMl8UtAO6pANGVeKsmmbUohRvGNShPT43M7YE6pM7Ak3vROlYNBPvt2MohX
2T4ap7zJf22C67H7VWYHgN3x2YHY2qE2cL6v8O3hni4xgug8G5EJ8scx3fAfcMipUF86aqEoVvl5
XxlM155sbx5FauLwrRRjdqvWYcPBChFKMvo6NIsyAOrTE00/cQ5ok+lRPyhA11CrI2kwH3Kyp5k4
8t2CAGnxay9A/iDNOwcMAq1tlmrWNhPS3WYtis+QTF+7nM7dMGUZReOMpySe+Xv2wfq0FdFlImEI
h2fJgk/YfROwlBkxrSf5AUzyxmNBEyq0dOsA1c9zHU9PcbV1r2dJGGdygY2WUxPz/VWFrL6Q++/n
WEz8wSCdi/lyWhJZUgg4l94FFm6c++hdfTF8QwZfvF1an3kjMUbywdJ4W06hSYLMMvYfjILWOiyw
aqcDOUJGUE4cof3UA4cNqckVVkTx8k0BmB36mQsHaCQFXrAt0jPtRiatpeD2x/d7Qw7vvuDTg+FY
CIYFP2RcJ5gFQ2R6GvsNSTl5EytOQ+BhFukUhwcUMMku2o7mTyQvetioMYzA4hb4AxiHC98UuxYl
cVGg+tgUaHKTFh2aSh5k8XBapII3lK8S3aobCfS06ecViLG1TV8Ju+5bwt2TsX/3whicIC5/ue0J
mYh6AisJcknBgBMR70tpM15YMcUQITi3NdYBfA3TCXkUQw7owEMZ5v6ZcREFSpXyA/ODCk3UzMKb
EhIeFkeuYDKtoxApV+9IedV1JlTDbcPm9jBy4EeOgyJiYMiF/aQpw29zbECWjsF/XYcyAcy61Qgh
UkGSmnfN1O/f8dulnQ3oAVIa5CxZvYvqR5jPZPrNQ+np+aIRWmQ5NuQT0g7dfWRTfe+ume8tF63m
z9vFpvWhyWDsrGEJoROLik+TMdBiZUUUjMXO1C+Bmm2B6MEIveHmwCTMJK8fQgHp2qCljKcyVGSE
oCu5nLZABnWTGSFF+rsCQtBiTmtGiVZ+iwHgm6f2ekcmzBXZ2CVPqpjt5MhGcdKF6j9yqbLXCo+x
ZUHsl4snCX4qTF0BToxgmb3uG8gFA3JejPYr4KPCpFImxFrPZjS64R1NMYys4EYFdIyrI7hfFqUj
rWvk83OpAvAKZHZ24iTKz84Rbk/nTPnA+sNj9nay3GxqC3spzWxNGJTWirUy+FtelYn7SvKOOv7L
cjcCgmn3TmIjpVLtXWM70Y+N/hO5uzS6H5BRKRbSv5VXrFhTc4bNW9sMJsJG3wWV6SpjyeRWr2OM
fCoJqu9ouPlS+/coNbQ0gUQnASHOdewRMPnSqxnOZmQkvfBHZf0zElNwp5/72wHkXOZbUNNiy4ct
YXh02Q5mDSkqe24nxYZUjDZT2HrjXe8GDbnEViiIF88rf6K1CMAvEeI9geUeK9ktWNDchk2SvlTR
4/lmqS4j1ugXVBpa0dcHfcpT2bI2tYug46aU4XXcrLBRrGStmnAperH4WoDT5IajbEQCYVzvkYDh
7lbM3qoEW2UKJYHGbOCUQ0Ft7TLluNZKli81oSqGCv+sMadSbMVj+in0tSiF3pgIy9m7Dzo+Jdj7
mFTRK7K/N0EpfWagod9c//HpozjagJoQU49hGELMGTeI9SrFtU+T8w/zwcKgWbH0IPlGJPiKaGeK
d+9JD7cftistHk7W0CW7PnNRkCMeArnu5qHJ5b3/Hfd8ZCwtvKk4uy+codBU97GCgievTRhu+J90
gY4gGGEKVuJnNTkn8sebiiWAy0xPz286ePSfkvx75CQnW5XHOAmbFYkxP2aqijXA93H7aN7PyB4+
bhVBuftp/P+6Os9GSz59V7EMTccfeS+9soapqjRveUO7hqJIlxa9RwWxTpo2qYgKo4V6B0Iu9e6c
10z+QjmE9G+V1R5dUC38zkC4QpYy8Oi8id0LfdACLWOthkceM/uVdMstPmNFIQGy4dO4Xq/+N2eB
8LBVvDuwNgFtT3N39tJONRu3jgEMJ2lvmgqzbJELkAOJrqCh0EcJDnLdqAwpX6hjiAiGqJS0aRQx
QsBDgPdemaiXcrLICgKuBAnYiTT4t20BlujOmxDaNzEjnJHq/tq6Tzjt0AX0BPvrbXkL3dS1zt0R
9VmLEn5zNshcd9whcCdEblAuAacE4ovmzX2c3+guddN6M4vTwyjsI182cHp9KueD8Rf9Ua2/eFXP
SyYBPqPFfCi8BtUw2yMf7I+GyqJNTN17+27AnXXyit0tkYb4xNiDQd3nA1FW/56qp404meh7QFEs
+OTErPIlN9c9/D0Q27HNlIEdR8vD9MHCxOOXNISFA8KZZ+WJ2V97CeNwZSMNGhTn5iziTMoxdI48
9PSuUTkWjiC/gmof+VhiiZlINqoQdhsIV0DfzrDgOId9MGU2QfWljRufbCIvYiwfTS3pnzvIctjW
I2MBVB8/OnJxg776F/zL7PfrTXKnbDCcGrqzCYm4Qn6AL0jpMbOwqDaN09HKhIrVbVpA9s5Vkyjq
vGVKh2ie52pjbQ3mDGQMAeaRev/nI026K2cIO2AyAyswqlgjPfnOVefQx9UCCicvIbEptwKmgRSH
fmkMdZFgvR+aFym0/0euvZqdUYoQFoQCJ2MWZ++TvjmgBsbowsy2zHFyzjU+RDywa36lpUUhVXU7
k+ae8R4BzzgcfrDAEJX/W3qwH/G6Z10deYghHr69zB0sRqvxMwFOy5dXGNbb8EqCm/18GqvMFGMu
UZiXkNCaET5Fi3v21GWN2c8tmAHga4zmt317J8Ik2CWuWKD/Xb0mU9FRULqE2Tlc4Y391wzG4bUv
BL1MCHvdDCP3hY8tJ03b1TqvFljXzoGhtf3yEM1JUMGfd5jedtnI+3PI/ssKWCsIDDEMsv/vD1Be
QDDQb9Q2P3yHMmZLSR7e5n7bM97eIKdlRjWr2atuGi7wnOZZ9VAIrFTMCe1jscUMyqTIG1XmBGqB
DoVd7yhWCrVkw/o+oSVF0uV/B+61plPLNTh0HgV56MzxHyeKuD1LLzPe0fqTbS9EuBulDwCRCpDj
X7jOxxg01QxSWZdI6VA55V8GKBItQhYB/TIRUSSCwi9AbLuh5ikWUN+xQDrc55+dq6TQ76EHDmQn
5tEvoGmxiqMGum6oE43xmpgyIOffsaQQJ7Ap5P4RGrpmxY4MtpOYNubs3CfYoedHr1joco8Vj8cn
0VKJOuBTK8L8yhpdKohuL2ln2UjPcJh1yfQHzkvZmxDYIpww4UVDKwTMjgw5+YLUNtdbxrdphWO4
mK4c0Kp4OXFc/5DjUQCDkqNMzG2Uq3O9H8bJ0kw06BsYiuHDMcMb6Aa6o1E19HWtiN+xJRiqRgsZ
Cm9qHOhoe5rRdX+FBjdVE3gOuFpK05Scn49dYZYmN8zdZyV0w5ObVODf8jSYLGtNZvSLPcXNYE3o
FuEgYmhulUTXGfFeEF1qvOTaFuESGc3KC7AH2pIQ2i4mfHzm9rXT/k7a2RfYDtZzvHF/5gGG2av6
ol0LhGD9CQ+c9SPxtNTECFvwg5NWilgh0Wr51p3Fygl/CzuNA/9kfub9qfFl7M0gXei7W658uXZ+
v6tkvS1ixvxWaEvRAz0uJ0o2NCd1IHLXaedew6kzumgZzzEkjrKMwVw3Z3xyIw/NUTUNWtGLk92I
QwR6J2AYAFWHcfQArJyFyKfZnpf7yDJgGXnTqEfKIFbn8bdR88oXqVpgCVjlebejgutkY2jtuWMA
jNyixb5czgetLH8yQlqPvlaqIlfeo+arHSR0tiNapm26yQ1AbtAk/92UN2Tz0X75fS9pSAjX3Oip
xSbxcRywD7sBLI4sllK7oY9z2SxGv012KHm5JVvc1WDUJwaxflVuF5JnNEZb0Zj7a1J8+yiejZtD
aze12OqGDt9jrZGWW2SKpjzT32XRc6eAOHoPDzj5zJndTGnW2pI35WqK9sJtpICHmCqVecNGCILd
XJRTiNZl457X+fIo3lDtWcBtmP7df70W6mlE8f01s9qLwfB0CzXghyZiV7inaEH+lsjn3OcM3tPZ
VraMFbxpwAxMWkrntFcmYhgK+zuhMjmuZOhuH+cf5ibJpncHY77GKEgvqNCiE1cgKJlQ+RnDykTV
uRs4EaSD90iji05D8cmPwX7tIrC2VpqHZs55+CDuxMoZvVwfwD0GkrUmzS8dfNQpp9mincShPfG8
XTkdxtIO98nvtuxrVoVX/g1IJWGvmc5n7nCv6reYFdQsHjLwD86TCC7iuE6I6dIt+3ySWdx0Ka0e
5zQ1Ks2MCn9Eq4PHB/hAYFePH3DOrxB/FAmG4o82grc+DtaOV672MO4PBfefr86ikVe0T3OytP/p
sPJa7IFB4VLmOt/Q5IpLo/GnRJf8zrSbNKYTzCwKFNV++zOZRfxjtZznga3mOlHZDTArFlhBleKg
3VxiSpqzLVXErVy+IZGFR+Ya35LG873o03gDy9BTW1WQmxzFLeRU6jSkj6V8Tfw374M8lgunYF22
KRcwW9aEK3y02YM0MOlpYD422KDrIrHsHRXcTFwmMQW3Xa3qEUR52VZQm63UN377YfQbRG8OlcFL
GAGdmL0/QuTWseqvaL0C8jNSJUIOIA+iN8rcHRLefHCjuI0Qmm+ZUGKen4xf1cfuM8Xy9nyiUTiQ
TqFQIW/kNh1FetorIrnH//U9FK9G1K48r3jO56RxCqvWi7Wv3XZkrp0Z7AJrBYzfLdCqqcSg23qx
KBv75MU50mOcoR3l/F+8TAvI//Vt8V7rMHOFeC8Kh17E2PjodcvsgDyWEO41BjHcInL3zeoYyf/s
0dEUunY+32x2VOez9qQ3ajaEu2hKHiCdl+5MDUTw1KjVLEYxWYjkCjAI2AqNt9IB1dCgQOSjZaK9
FmrvOWgoKqv9s/WQ7Qs3UPTx7dd6N+1d0MiVF9r8trtZ85y2RavIDJrA9gf7gr3ichTqW3UBx/n4
Bg2KKLzd4o+1EI1+WG6qKe1yq8OW6QKoK2xEqYh4+LhTSkaRH8vx/jjFXKmR9pq8Jg8Y4J/q+5CW
dRcAictrAWEGhhBsJRorW0ISoiMua+Fn3BbAs6phnO1RLl89oet5DzN943RUI7Js4++XddIRXuMq
c900C1nH4TgeEdQYEAtjTDtcJ3WJd9LFgKvLKf9Kr0v/PagpAeUQVrqkUvmEz1z9ql5s0OB8Gye4
pjNLxUZR8o6qQ4aLMSak8Ai9/6KU+PR0mWXxL8iCXGn2QOH9v9cMWjvFHYZ1Dk7B1ryhoQ5Qkesa
/4xdlxpHxuHiQBqZ96KxSvgXGJKu6cYAn7SiW71Ch1+IwtE98Z560TouUPA9lnBebeEpKm/fJGss
ZqN+HFPJ1Uva0n4evoVNwUPc6GkKbNMSyci2cafE0UZ8KzkDINxPkqY1v7+karvnZpcCxbMWwX85
vnK1Xdo2zUyCboN8PelxiPWsIx7HvIqjDyPIibkrAEWM5bNoByPA3osQzGX9e3pcwVJncE06r1kp
mfcnskndt0btsR9rXx1RqjJuMWzFCt/NpHXXw16vgtqet8uBS2LM2pCZBVgLkPz/+CfVzrP3rlH9
r4qP4qz02WYXmItYwNHQRBKlphzWhH7Wrh52AFCKjl0gFBViSlDBXsOlxiopVB1EBnUMKmkvOYX6
WEWhJVmUtQp5Wt06sXlbMO5sMFMgFJgWgluXVYTsF/sH+XD3yo3AgOaxVp7C5MTUsAcyx9CsRZ4c
eQ+hUb/tzFBqIPiW2u0AhvAfTE4ZrNQOQ1PSlcZ47M+Y6wx9yR2WeavEYUDE2sn97gDp3RFcrY1j
7+JMU6a7gg1ODXgtepN9e+TZEwHZ4YH73JhiZRYerpjMRtZm4sf8scpCOH9jAL4rmElsa65/AtFZ
w+TtFJiEMrzq1Qlp4TBQq0ask8HKIr3oeeKcRx6I6nP30hUclJsObwIgF7xq3ChDrKrNCpOkUnjs
yyO+BCmPZ8n5weoEm3noIok++mK7ABrF7HOMEjnf1VDIhIyb3ZuGiRPYqeUYHQ7Xye+pYFcQSVFW
XPXdhy2bSKw1fjQh4+sdO19oLy3LgGdr71qy6xzDKtC8TJVTN0r2drWSvBHddb/NKvIYGXlV401Q
Urh0WTvXTFyvZlD/oDJxexUGwLYJ3nnLC/4UeRo9g3bpk+iOy67B+iIrwggEU0bNPf/VGZanEd3x
lfHji8XI4wdQPatPwxkcv4XYnsFI2CA5ZXqBwvI7SqB7d6awcwnpltPc2KZaBzM415mMHKvc5N21
8jugKUfnTc8xtvcbjW6ZusRseQ8yeBbQlF0QTk4g7mAoOePH8pUtjLhR9+gnXKz8GcafzXU3PZ49
mkZ5DWt3jRUrl90EuOIPXoHR1hjyyzN63XFy3Rva8oQqh8I0oTGwTVxH5p4mv3wuxsZLFjx3zfHj
Ake3B4VEr7x+/exIq+D3EryoftkV6zBvll1TmjuS5aIoMfK2wC3Elo5VgR6qywLZwbi3Z0vJOpnG
W7Et/+pAXZaIa3oEA+LUrhCly6sS2dFEUMu8+NnMrbqAASdEhD3l413AJ4YR3iFpzEnty8PIvjAK
U7f9vMwmDXVHKR8bUMLkC0Df+eksEuj/W1UU/2eQOj73SOnXX0dQUGfIBFX47e5ae36n8WWn/WBW
psgjZ8Ix3oGxjulQ924sBPQmjLwtaFDr0nA6lHVqXHPbRU6hjUEDIOmZbUvVA5mP0SgpMv2EGnHD
7oxKaBJJ6O41F/nCMVJOrIZnbXQngQdiufkPk1Z07AW9wD2/18WKNogZLNFIJqiqnX2Kx71dvLxu
MJ7gyTlGTi9iH+zGompf6YTTzXePTp2BakQmgKZe4ZIoeYydq0VKLgqNqkPjeygp+98FfnwYDOwO
0SUPll7hUtIY//edy8F+zmFDkO2Yj6JFuN49BKJU7CbAfcXmRu85PJ7+h0ncOVFTntXTmh0EOLB2
24abXw9ZH0woAGYzXNsC7ynG6+OYPrqjwumSHn0YIW9wrJlm8bsFfCxqnlhcbuzM1VOGUDxoyMo7
bqOFxiezpt0FO7krPtPq4sZ1q77Ssy+OYRPypzrGy6XV8JOvlZofzycnLYzv9ONH9LvOeNJ+JMUu
3x2W05OxJuAWdJnOsLuBQUQWyYH80hn1+DUBzspa88abndCFZDkyvStjdifwE6oiMw2cyEvS8XAn
iIonhRrOmFhlB607wOoPhI+yane7yFmJ3jDn1ugLDA0qmUCBeAoxfw+qXoC0w8SGEaDoNqXFx6Su
QUJQdC+IJK7WrVjpVruvhgOiOLW/slv9XaygZhlwcIiU5TRgiHvrepPa/A/SEnGonwUe4VJpSOYI
BUw3OeQ+bP+kWRUqMTT+NL23fkYhn9hkoI9EFQvi9qdwG3xuOLQCLenEJotIBeD90WeXKSbRidz9
3Z7PMUn3pMed+9i2kH5Sx3cAboaBjfHU3lkGeSTP/emGXZUOMU4A5h3wbkXyLZogwlzn1fmuSTCZ
Ap8aFxMS+AipWtuhxxxa8ABBXP6kSJjN6JngD93rP51X/M8+SnPPxJr0JZqGkezOa0R/d1PVVnoI
9c6O+TPra0Bn+Me31cjw0e+2Ev55gjJQEhvwnoi8Iv6/4l+gzgZYxIM1r5jlsHbLRDEr+LqkAcHk
Co+7D6o/jMZ8WRP/ZiyrUEqLLFxFrM/FdnJdOhXEuNLCTGm99uLkHM+yPh3rZN7zcsDA91a8r8/z
8GCob6V/oaT0CligfS8df/3fK74+ZJ21rjUAgsIduo5lPRsj97lxW+LGGNDCinf/in6ualy//sbF
SM3eoJhJpWNIL23BCIFyFYQQTyZ/rD8wambQ+fHgcdJHLcGBTtFq+PFgb4YiHs/eQgNkAMkTxV5A
gXivzAvnUxJUpF6gvqS/F6Fsvakds1jRzPQSIqK4Rrmae/2k4K7bylq2qiUHmuMpD5jkh1lL0f3t
Fa/L+JIzMnavEUnxDSPGqOF/Er6bDuEye5OJTEX4K4oZZx0syyQAKtCU0H7sHS3d1B4vc6xo0kst
03xyWqZwSdlFr0xVZ5173K/WujattCuUf0TpDxcIv12+TppkpYku+7Gg6KNLK4zjhJbLGZqAoXa9
50wo1czJxA/OgdLyK/uEgZniq4kmg1PPEeEG2tM87L+PRJHzKQyoLwfUXvqbt5XBn34Oxg2afZOs
1+SSTie6/4h0s8PhsCyJeGmKZOmZIA/TbcFV45mLl9Zk5ExH0ISCkyaT4lXGwO0UZZm0UPTLzcI6
Khi1CAGXbipHcy7QyckwcZaEazuBa9MKUyPGDpUKxjAOArqjVviysCPQ19JTCqKFUztntr3bgs4l
YBGh2dNZqw7+XSTHJjAq2hhirp7/Jqp6wQC7osp+W1dc16lIRNoKZYCj46Dx0ZSPkCVf3ivY7WW3
E13h5usYCm8XmUVQ1gx3O13QuPj9y8o0QFCygCKns18vmoyy+QMP9BrFy558bUdOVAWs+QfOCW/S
FOFMVFz6GeCVwpSyw+ue4g/9ru/V+KyzdxNB0LfCaDFyPEcXZl/iUhDDN+SSFB7TR30h4ONYQyZq
SymOyAxa+bqmxp5bABTlj896wvtCOfY8SDQIs8NvEWl/kZq+dUL7GrcNzR2e2A3yL+yb7D/ugRaY
QQu+aR4lcOAXpxJADLPVdxlHcl/aP3FKlv4oR8T+pRSxUhU60qzrO5sTAIN8t6cyKGg0tBfLIrXC
50MKs0oiEja3L2uKezltbY+4m8/4WABjHJMRGfZsiCHbXhjA25bxexKK+sHnKVciTwUtZFMTaIRM
w+5NvDnZgKWUjXnXKYY8r2jPmASgaoiFeV6Euyj/r3Hl2CwjB484R9NXA6m64RMvwiTSvyqansb2
jngBhQKaIDzr5lZLxyW/uVvrtE2X9Zl1uIwGk1DCogf9YZZKFx0eRtxLoi2H3oBdlZboxlosOnDj
ZsATeeuIrYT7/JYc0UFEaNVR1Zy1JgBl2qPVv/Pyrki2O6+gKU//Y++TkJvWWtbnFS9SLjutv1Bt
+sy7/U00Y5lMjOhxku39F+c0SY0F1HW2RtXD9TGuqF019hf3hdYBYa9Pqquem+yxpMaPm2NwEUWK
TBNdHdZ98q8Z2dDy4XFZ9UxuM04uQ7WxOu8t+LJo0i1yTvSlZyZkf9sagsxBel1G0DozfCftA+/t
Ht0qC1itcph9vV18zu0lNdKhZhBxgeQ/ozYJFxv7AwzZVyw9/iuXFCRohxaIAUUiP7Gi7wSHw0Yr
w2vR7IWlzC6YMZdu7eDGRIDegQmYcXut/Fp1+wTSvypR6oZPt2zTvvIyN4oG55aIkr1wZ1znBPl9
A2gXLGm6cAsWuLX1E7CCFw0yLcNeLqlHZ78in5zQTrdhWwpRYJqXNaUYwm7wBA7cad9AbwwlA9Te
YI48IPB5WRBpZXO5z2hlxXBOX2WxcepENxZzwuqUg3CPAxXXNuuzCZo5HyS2ftBFC8DDeaRljUAt
r3VNqFaUEV+k5IFB71qe6H235tvs2xaYRuvLIQGy9qHKbX1HoVMs/+QKdqVCivCBDWmJ9m+5S3a5
BpaVT/0HP6Dt+Tv/mYgoRe6aIij+b3ePEVjkqfMMSOT40UG2VVYUsOv3fKo6SvQjxQ/z1VqZT7xG
oPNZFxRpMrZIqNPPzWY6EZeWVX0u4SVUrwSKitQ/qz9xgAYXdQtRtAaol85iGStPmIvqWbiVVhVE
tN/2XtMbo6bvUm1F5xYaH6DsMEXyWS1VAlltb9RgsuMN+CN/bJ1afMpsMrGZ2a8WUqBN4SLBOrJx
ot1SWPzlIEntruZeXUcYhNBSQnUeBvo23Ot96HscKUAqcYSy4y488VlBKP6q1V4wP90HMythPg9z
rH+8H+Swdho2W3fVp9gaYpVoz1tKb2hYa9NFJAIuvWh4MrwDYf7KnWvkee/433WMCSqDE88Q8mIA
FmkHL9uUEgkwqQ7nDXF3gM8jri/8RBbP6V+z95Ht/1GPu3uAUBEDUejCJOxIynGrxvPne9B7+Bj+
8SBiNkaLplx8pdGOACClZ10185p5wqOnwSuB9J2AWpSTSf4yy4FfEKrEu/yQGz6a+SWzqvAL+zYp
Yq50PXpND95voIaw0OpvIpZCA2pW+O1+dpeER2NI2UtFa175n3kUhbm8RP9GNd6T4Xsk7nRvPdYU
zMvO/t4EHvRL8XiM4NGZ83Ot336sxpJIsWhP+otuTJqYzScoz0knPYMv06hcf5A4s6Zk6Q1sFYRQ
Zo0RhCTBet8+NnK7DUOx1c5fMt/2h0yimrpa77f1FPys8RBcKW2EbvFdkvnaUPfnqtW7o0zcrMuv
AITmxW1gKoi/n3SGBWSY49V4NFCdNMKAK57wwrkHON/zxg5wiGm+/qjEMyISvwrw1fXs3qZuuPr4
GJq/3qP6TEpFsh/k+FnkTA/S9jpus7ckPKZ5OJfyPCR4no/RzkeI5r5RuinEzRkZkRurYQf2Oomp
/QacflM5Ss605FXah5HX6OMnZ9E6oC4rB+SH9wbatLJbsX9qfpBFsGBNosdn1xfExtd9CcwC/Eu9
TuHzZJzH9pRM39MXesyLKx3TpiTf7hiwNbqDUiyAJh80PBcaBNDldhTebqIxTPV1durI1VzoaYk+
vq8kDmTrBFMEOPzGz8dEcZxfDi9cdyt/qhKwjDHd4UOGMrtwroUfUf99R9q94V9DQrjnf8MREhPc
MGZ+mQtD4DH/m69iU5aJAGZ1qMMw7noSVpTYCXBM+Gt0LOeg6C4ZOAEZgbydEL6HiCZ01ey20qeu
di0QqJllTvt4EVBbF9+ECPerjNToVp/HEgM6MoER65HDwVGuwD7WwLfAPeA8J5Y99UK56x3YWIxn
HnLaOrcQQbVyVyOdwX7D/+ooq0uY1IHQ+IFW+6O+IFpv+zcIEsqxX7VkMThaLSBov7MHDPTm+erE
mqJkU/QtEzE1qaV0TMOa8D6L5DjUFIbjbOzRDJ1Ok7cxAfrOUuh71MiyitydvMFXpCk3+xYpe5lQ
0k5QlB1GaNcDewQr+XQ+tsHAT7/dC2TL9e/tStQElEYdaO3I8cgrXv01Y52zWCv/a/q9jDbNMNfA
SkRGafA7CfTrDAAFDCmfHdlNP5t6up0m1/K0Be/JO/EB5myfOGlLBLdjUY/+0UUbxO0EJqS07qkC
cakkRZ8DI8y/rRVg4bYGI2F61OcfWTAxvUA0AJR41N3OY5JknvxvLO++6KK26b/xYFSER0loQnLJ
9IFqKB13IsjPwWt8rQXbVLNb8cJ8/XU1Lc6uGh6h+aW3F/Oa97VQe8tX+ie5fCUuQMQWsFzTWShI
7fflFSiSKZtT1RAjPh9LOFpVASeb59xPzdJjerfvtDSNpsnn7UV9pM5woVGWOkufJDy1RSmn7TsQ
fWf/w8EcOvVUR+zcoUqFANaCGPzouSSooeXwrTOOdgaPBOO2vw+RGHhe60r/ecKe+mVhDzLTS6zw
aj8suz4OeLTst6LpoW2YT/nZyCCsu7mdeQ4dcFPvMaosqCDYXYHrrHme7v0bg9GIb+wJ2437z4GU
nk1VlerttB8t+daJzjcA4jFzqp8qEsbYffQwpN0+9MrsQBrMheV0vxPEk4rjvAWMUBk+ee6tT9di
vZNGGY9+nH7R65WEo1TqSAcH1A6Y3iBA/N9XDxIGqNTrUAPY9cSvEx0Q23Q9PLdAn/TjdzhARCkc
GmyUh7CjYKEQOgUpe/iWbGHrL0OE8UFHhotsQDWP/AuIjB5XMTeJorkqPUftiWD1cWPA4cx0O9Vo
2v4G8VyTdiXrgRvbB8BjhdyX1mfeL8zNM6qUSCFidEDUPZzx8f8uKnCMD3gnj4K3KIVaOgXn+/ho
Ve03yOKRWWEc5Cyh0PNVkAg4rXHxtCSkw+sYZTmWXUWFySfg/qaOm7pjJVqMRqQPibUxxatR5rH7
fAYRepKqVILjCuSC1KWZDlWJlvr597jN/gtKfzFlMIGhQV2wJm2LZOrlIVyw8QX7zmFYACaKxLkd
S3W+2WDKsHm1oyQhSkfkghX9fTQglNvpFlLsd0QUe3aBTf4W/vHJecEBn8Kn9J5VPxfRLiFgWrno
PU+SH5X7pbKK6O8yiBu1fyW2VrNKK4BnznD75+T+jY47Ofc4T1D4CuVzCX/HdPwVtURcGc1p6tA1
VlFDKjX/Q1P94lgj0D8qtkh7KKoBqQo1Cw+nCgZnfcq/eEdf5tUbE1yPZf0RMWEKTVOiLYr2ch5h
gq82L0hAzdGSIc5tIREkff6speAyKwUX+wgYEfS3f8O/y25J4M5FhZnmX14NyRqmnzbkax+uPKaJ
yH0p9IiXLU6NUGt0UN8/g837br7S0dFi38JbnujVD+5mXUAt0KQ6UA00+iqiZWpnuFBpxlYWVJDn
jHhl5EZjp63PrnXvMkBYn7FP4Qft2ii8OkggIzBpHqXADUOUMJ2VMkiCU0aaBlkcfnQSh0heeqyb
t5d9EyAtxP3CrcuZUgZOj6mqev2a5yS0OSyt2jtIQaYIK1iSNfliWSZsMWsG2rQX0A0nt+E3l6Ua
vMmFwkiiceoYloQCMadXgRzVLiQBS0yjDEoEdEIoZBD69+ikKolOcs7ZvafjCnzfv2/r60hxIzBF
EwyolrPsNz4VIGyLpHrwBtJItb/jwaNsUO4x5lCOqRN9GuTgEf1kwDjJMSOE6KppksINQBV8tUmG
xJ9Ez0ys0h8mmtKh7vmLR3yhSPKmnSzxlcrJqeuXY7gpFo1Gsek7+hjfQ+3PHcr0kZFCH1IYMMli
fm02C1atNXzziEWMeN2cHNV/KyGAfjPuYRA2Iic0gIXxYZL3+YOc46CGlwv/YQhxZII+tfJ8yHqa
BzKxvRuFRuS5la6viElftn7eHz0qynel21F0Siy0Aaqj4/Yi26+N9WdB6D2FT2w5UIQT8+LumJgC
nY2WCCjBYDf9LgssPdRmaKTj3T6lXLZldygIZjKNOuDGeeGEYsszRzsKZKl+ysG28i6s4f8NCZNa
66MmtQFRGyh82+HnlarAjEXCRi+EtZfY5Yr5ULErNXCmg5faEEXiNCuzo2K8YlNIuquNdINeJwWE
ZJ3x5jNO9ef08Ei1u3t3iexIZzER0pK2jqYUXAWuQkPhnxFr4MMuiO6YZmH+5CfPIwuhZXIDvCsY
82H01PrhTE6tq+UIokTFOfllu1U5gdJAl2UHcX6yrzj+GTIiiDUunyLjWURan2eLFKBKwHk0IJtU
0QrHQnrplw565n8ldDjZuA7e99ArODUcb91K+a1frIrktex9ykYQ2Y9ItfRPVhgEjvXq99XLqxUf
aVvJLreelmrfViE6Kx1wWiBWpLe6bYJqWxCmuFQUdOx5Wa7CQQxmqG6oCt0YpluEP0u4Q1LarFKK
fQ5kyIjhqSNo1nvJVAWKGGSgqBD+nffJccjLgsbBu+RoA2YbMwRQ5fez+itVnBWw3i4OOEuGVJxD
ms9/6488du23Qknu83VcrYPOid/CG0Jc+WWqoSFBCVbiIakRCi9n0HUmmbFrURCqG+JjSU71g9b4
NsBwqiMjhE74nf5C0LZw9y+mMuGuzsl8nXX/Jw6SdlgJ2fAZWGd2O9+5ZP8JMSQj1OQMMqSfJouT
AEF/s90uwQnAw0+7mZ7yk2G63CfA/8wSZr52173rUeLz83x0FTmSYllgjFLF/e7K5/rwk3CYhgwL
YGiloO+30BTeq6wptXg6er+9MtHWuJ3FKewkx6CPRSrzXgLIhQ+N+Qx8a6LBRCodJjmcbE0UNYdZ
Z5aRa1SGKZVkb4iT9s0o1F199sbAr0vFDWFB3TmL5ZciQFQSL6RjhA7f0XPRyB5GrpSk/Ag5BwMH
qlkPG3OC3eKvWh2U6d6K6IxZCBrXven6JCtUCmr0U/L1P6T93aSqPXuJPmBXyysgqje1MzkZSu1/
1pamJKHp5aNqTrNiRwWi4+/KRp1b84vPzaeVdE0pGOsae8Xp0VWPWRZNjyZ0q0D7hLYpyi45ctgI
t3jvik8ndKy7ywdGgZnLqvxXIcfbBRP+Jwrn90H/VwD4WikkQsUhDiKkIfEP/h4usJWp7a1TVzbJ
FwCKQMcAhdI7TWdrAKEy9A6VQC5tKvugYCv2ZkYK3iKVF41UgYRY4QDR9fbkrrMYGCsQnyhMdHlo
fqZJ3XEl0spvTfgklIOKf4x7EasJoLaIwyRa35DaqtG/n7AuYD8RGOJ90PUVlFrLHhWUHMELluxh
G2+6j41VBVwFQVOdM8EXxaHYQqlFwIWllXh5SsB8OkXT/i0riIV8GDcIc06mJxhYnNmRxjt00/ob
cHlfHxO3ZwlPXGmR+k3IF784WNHVCQiErCH0br6P/aiFKeNpkwWSA+D5f/MWMe9lSYB/XwEvCcGx
DfpSA8ZUNchnnUQIT02nd0DjHfNLISPmdiOuSa/92fDkqYjuINT0nrTOy/55syf2U1CsLU7/4Bjb
xpn9Y6EFDIXANFG1fV2+2d7W6r8xGxvD4RtkJRWT3bCsBTKlrCcypyTiSEUVayziAaNRCj1n/ekz
QYtcPvdGbE7vDd3yQcFeBc7njpblCLLDH58jFROf098wjUoHt3hcQEAF4K7skc21lb93XH/FqIk4
gq8pb0vmfjFmeOuo+lBimsRJS89ztv7X8PWEeooO+hWapVkD0OqCOHtgJG6gJo7g4ql+pEjCoxWY
gj1bYJtYkyJcTdbZg6d/86Cz0bWuJN07Fh+qEEU0hUv3SYM0ldikDUGyTO6mS6mepAOyLKGjjAUj
FPHpmZahV37KRaoT3EZAeym5BB3aZFo8zQ+i31+/R8sRYL/Hd9onEOUV+2yCqacsYL6zYEtcp85l
jYBzfT9XRPGcSUklLCbNvxZgAg7wjs0fRa7d4Ni7L5FHC8+eFXFP/8lC4gy9eZRXbFSu9bj+xblA
QknpCQD6phhMhYrsXoFzFwVfMmuKKfHrvD0sYKzfYMCBrqIQUaVxKIzQTIfhVp6KEZtLBzqponp6
/24RG+AGqbs7oGITaI/AHdMiK2TSJkxO+MvqLdmV2PSgYVOtkwCJlMkZvr3EIHKwCcVEyeRFOn4U
laS1vwNeqPRxtyDsrusNe7gE7MKGceYdkmvWlge0xF/ExweGLkb8ft9jqChZdVvqbNmoFJ1MRUaU
xBmvNxdgbLLQRN77cRsVifCrEe8qQxzNOfFmHDJk9QwF9nfk2HNVfiVpn0aoV/4sH1zLmBBJDfaT
OLOMWwlutNZtGptPzNd+lqz5LsIywQPIPOgUAuqVmgGqlz3e/eGkEBWGaiIZ7DtScqxHPt36Eb9t
xWJFz9bK3fv07ZPUanrLY1QmQwHCwxjKJkSh7ymjMdkzpvKQbFB1WYCamnbr3oeUc08D94ylgw1f
pKe9fhco8tTOZwfiEgQwEusRr+rKfqoQsH/OopA26/6KQZ1lkT58RgANx2AbLsVYtn0PTmd02bQI
50vpJ+3SS3tcP18FLkPofSOwPQR6RLw+nq8/QhqBag5UvbhWVqZ56homJLPNeNJTOXPs3Hl/Zplv
vFqOqNBvrHeS7wjzC952xiPekKesgB+yFMzjDvPKKsmoTXbkJ2rYuaL/J35KXGnW7+rKTMSZGcnI
cK79oRERQ46NWWaJv5XyX+PbM4Zjx0L+UrLqJb4xu/peBl+XxhdPV0B1d/375rkPW7SwbB/3pw6z
t830toOJBYR98sO+gstSOR2DlHGnheGFl5Bie+TUAgK0dpRf0m1XKZg8zW1U6rbAbY4NWNjHCNfU
dsvfT4vX4S/xCkL11tYtyksTTDoN7hG7RjmCZPp/muHbs3t80FdbACd34XfAntfcwJ+QCgoravr+
KftjgELXkHA31QqqMQo2EZ26VDRHSCIcLDkikpQ03GAr1SouLsDo9KtOAlekwlwLPJ0QYsoYCUSp
T2VRRNCXwow+QRIbuAI/2+L08nykY/NsEy/8NSA7w6r4SHi0qYOYTt5EY+q4ljXmCD7QhWR5oB52
9bPdD1rNoec20E7xqQP9mPOqZcA5cbOX9W3JMkOdiBjetDLjSq/qI1SnZ94IUeeaoeED93YDgOCh
xpSa+cRaOdGblnbV41kdQ9l3eMBkXMJPvQdGTSmE+GNllcFSUOa4CKcxcYTnJaa0QOwJlBWKYqc1
DlBPbRzxqIO7moJjFgvZJSqfSWINBxfKMxdbaKpUu5EIHXCvkep796reZ7oMfv35HJ77/Rhw1O0z
1snEALJ2pUW41Iys7DkUC4J2ms18UL64e7VBF2dOsbp2IYpWPN0EPOqELTnx1t2lCo429SHyYeMS
EF0N6nKKnQ1Zu2Na5zhjANMpWYwy0VUp63PNbHwyBC7B1EDbS6efxTcK+LFt5lENssy1iG+W9lh9
zTGy1pY15IBoStlZm4/MCtOXASOT+RjxzDBGV5XkAhElzgQ+m4qCR1CUWcJh/K/0KVHDHpm6QFe1
m9W4bIAMY2NMXT2/fuDseCX/gu3e5/+/bf5LVKkJ4iAXFfneWx1WJDCfPyUDPArxq6FWrCaCNKrD
wFfs3Pk0sJkxO0XonPas6CzXn5FT+zZayQgxpbcTwv0fxiIh4VhY2xVp3jyeVdIvPfw7AuWSfgfy
zocT3lGmbDaXrpDTn0EpF5fZ0k6MisaPSQVW0lCi2ifcVFiCH6VqDI3LTnM0cYALU5oSKY2HWpVg
ANwYj4c+HoZyakId1XFKWpY5RGmAI77x2ZpEh8uq4BdAnQxIMxNX+jWmw/ZQeNHdv7nqLdCUl4E+
B+97tqu4+vjrpXnOEWJSPL0QeVdovn1nVkRA7lKE2MQOm4BIuCI1yyb5zhzkTF1aKHypAcH9C1+q
BEPO5bmtWOgPRf/W7tUz21AXHOk93+kDgwgJRl9TqORwOisxyvUZRiYXJEQMhSEUtzv6HWl4dsB+
amBaBN98oTzGmsJ6GH9kb1yQzrHKyGkvavGUI2Gi0wEFAYffZ4CIHH+z7g6+bWsQm8EsWc+4GhpJ
IG56zSQd0xN388GB6o2l3EssHKp4WEEGTNdCdSG9fcvuiEaryEXhZtRTnvmHoxpPwanV/z3rLap7
uKpFvk2UhOud8b0JGXGRgiJnFnqecj23yyNXLVqpkE9SxStxCtzbgih7OHtpfOBVEG/i7nMu4mfJ
t38Zy0lMFonpHwHTgVT7N4upbvy9uyOpiK/qTSrsTkdT/kp2giOD6lGY95Y5/W2hVLZ8DxYRTYL/
XzeUVxJuNmjM+GtApJHwbGvaakyrXL1xwPQp1zHGJ/FieTpAohNDQfCQQVYhHeTGH5/Arxw0nTog
4tQA8b18+3aptrJ2XKZQCK/4l8W4tjlhAS/JmUGtR+HrNcmyClnEVYah4JH8Q6twt3BSrPwRNXbk
X0HEYukWyh4ho1TOVP9AAkO6M7eTd2f3jbFXIb9qTmw/rxi+sZKtJXeShh9YEiq1Hb/CsJmYt0PO
eNGU2k6wSi4JgxMtHvoIHy+msTTEy7LJ1NfurTAtGLHrEjaZ2/YNgWwznUxPdfKZZydtvUnMF/ht
2/kG1mgAddxrJoz0vjY/qm1DbpPPi05GNPgBDYVgSv1eUOZtrGwlx9qhHNJjFYyTPpoerR/0f09U
RtD9J22eqt04D2ZMwNFCmKJwnvoNciflFPzevqu/3DFSZL1YZ5rotTZWVIUyTiXfHz3od3BqYm0h
hoYrk1SHiBYQCUQrCT7TkoD5GksnRNivJjGI/Z2NeahtkJHLKwYcqcgI0FfTIffTWPXJaaSc+dpN
nOQjuUsUs516bCDBPX+6GQATdfBptUxOq37ZFYTseyv6Bvsr4+t9568Ja6/YkJ0mZnBGrM/Zyo5J
9axt7fbx1puDrbrjWVRkXNvXVymmsYacWqSsHdfz/w9vB1oF3atlhpsAa29KX/QQ7EHQwfDY+DH6
cYc7nGXqIMyu1NZtJkR9jjxoq2fSw46AMjb+Dc3aaRyVxhtDTpG6g3phQVJs5K6lsYoviVKjSW7b
4fNpyn4Hfa+Klqmcum+el4LWSux/0hasfAauLCYdxD5FU/jawXOhxQJqTvKc4TUSRHYfSEaibhk9
ZyLp70WqaAUH3LDK7Qfog4Ub4lilgAFXHAp2dW2Ap64vTnYOGsu3Zq0RhVUJWVQWQqu9xXECvDYU
tPT0j7aC51pzPfDaHt36elmqce4hwwm9Z6go8FdFG5bQh82Fc536GKxr70VJ+21cWYH+JId7q7Mj
YclrxXqiDnnqpI+/0ps1a+1TTJTwdFjWzgrYICye1NncUn3S+50nyWjgDa8AzofaslIfSRZ854qD
ly3pL90KmZb41xC5s1dwtXJLci6f1nziwduOOqeXMptsGfpI6U7vG/Cr19n+qq2Q9X5ltva3fe8N
0Qvtyx76OvZ2GheSBExpHp+dEfuNrTnG2JXR40wvgudP7zkhCdkvqSifZUFFh0SLYTcEXQcvApN+
xBbYHt4A1ihA+Qux7qy447I5CPZ5y7mYSgoe609VAgl7WVGb742ifkPQqEaNhFZSEkNyIR0x1M5l
e/W858qykkhkl38Gwb55pKpGZE0doiNXr90ew2tpZeNY85bHLpNysFyFmmFLrOJgKMCmKt+Q7f+2
IZx/8/2zQHvbJOIhuMXg5PDos6Mzn+QZJ9r8YsQsc5U5uL0Uh0YHWx+IAk9lDovkZf1INyprTOgL
DIXQPNj5Q4rvTrBbpVTehoXwSO9WVmb/1NjgE1AhUYaGoPilEfcUO33tKHzxOXH74VcblZQfDNsM
bcxIZLbwJO9mS6iavgq6WSYNqPm64fkeaknLu61pkCCLdubwwgMVjrKzLxUrVClPbtNe5AoqE0rz
zXnKwQVFQY3GRlUvFcUnuHBKSm/zkJLI3MXGL52h93H9LdzBPBXWYoD6/qWFAOZTpV3lerCAfpXa
93wasXEc/SZX2GWI49Ylh1Y+R2269sbL6OHc0tnJmJSMxoUsprT7RS/hfGYSLd62rqTEefzkMooa
ggRL7a6UPCTI8AAfE7tGsq2rLycZJqzV59jajaaWx0LPw2gi9JAIfD5833+NQHrBjHjRVNqQ4+uV
Iqxw0Eyvh4rXStbNaLQsd4akSoja5ehY8YkrQCci8hjoTMN2IZfvL8bytVyt7sExqce2AiYDK0dh
c0YgC2bChXJXW4P+COnYo4bOwKymg35zXPjOeQrgau6pUxO/CkmJ0yYUUef7rpSNqvAUEPrswQOX
SApEZpsHy8KnVcjhynu6wgTK9+n52AwUwYwF604eywxorswDW434Zug3Og55wUUNb+9Z8jjp055/
SVUIwIBeVRVYp0tof11KSD4TkCiJbO+e2SyRy3T4t6o5gOD779975EdkMB6JNjkFJ/6tdSTdmEFF
Qj3Jt67l/LwVrtDq9gahR3NZeC8QEW8sT5yDv+dRlucgGHYw3EQkUeBEgRxHn/0bZaW6hSyXPIM7
3S4BMa69vOMUxLyVtbNhKXy0kiXhdzTHZnkj0zDnfSKjtRGwrBqD+QcbkEYjWlPOrm4UqbiYaHbt
L+kQCqpenx7na2IOOw3ZjVuhBCvpNDCeftaQLvwxzG59ktHvSO607jxPGAclhOqXDmr6xcrPMfza
/Yeswg9YKtktLGWH18+67c2TBm5q/bpqlGopYi2xZH+zJe9bxS+qzYjTQh4f/S6GQXcVoWJIgMdu
Mf16TstrxPXvlwxG/xjw6HCxFfDSvVn4mj8yBFYUliBY6qf5myOGsmDvpXPNUAFhuXa8eE0Kk/in
2maadd2E0aN9AxDMWU84GlvuUXAObGlvtstOsQJUiUkP5gb50st0RkRFpSQhUY/QEh9Z5ai45WfU
8KvWrNC5sHVT9i3YGtOAL9r+LNlT5eVSNp+4UpR1oQdtLkTadqNiNn/QXCJxvWfhAjrNFdPcTVBE
VknmfqgZD4A1LIf+QNnpwqPHoeRwrq/mL3cuylGNz7GkmeXJpBzf1eUWc34TVjuptKjgOMYusK7K
2wAv92rTWWlyS6dYPI6dEBfOWOO820zubCWqxCJMl7uAV7tlrjEXc2hejtDQo4H9m1PLBiUKPgm5
m5eoC8fWE1zi21Ql6LjyKvZnVLGjdfHAQIJjz/U9zHj82GsO5TqNhKm6rqmTMxUdYGVrrmTjyC1b
NZVPyyhbbxnZURjIcTRImrvC3RYipKrS1jB+lNgyHXMUcynJEe+kqXcc5/GSgvwlFjhcBf8GS9sI
2f+YKZipoS0uCoucocGqYABweW8nwzgsLI79sVRNIQwHVWttzpF3MYZbgLGfPqe2AGavQhJx1JcL
ms4o51UvS6gU94KyweRWeYKG1PT4v9RG7wJpakq/Pylx4Au2yb6FlUHHuwCAdIDn8V+D3V8j/Ezf
WPOmqrPY/Omodxtp+brNPc9SI3XjmgtYM4vCHBjEFGWrhQf3ZQ1HNofP5X/Xa6+q182x81GZUWEM
rYa7TlyPLiHdZrZX79fPXEMPm+h0HFmujFqOl+I5YrIVvDjlTxa4W6ZHgWJFdE69I43vjJHOtXbB
aC3xX+rLdTOtykjQNNABpq80mu67CPeqa1IsWVctpgkuvN7F1TTZfoon+0HzZgTQdz3cy0XTP9gJ
Q7dWKewSbCOTwB5Jj15W/89l5r1iTc1dz9k+Jyhc2JjZHJU1QXO2L4sC/2ywK9D1eQYyPFwqKtxQ
V+ftRv0VYkR6QXvrs3UzDkExvZysNm4e64rd3/kefxlnx2PMUx6DTDqyuiYQ5TK1Zb6dan7WthY4
lfk/74qda/64RAd4T8fsy5ToQyYFTl3LI+NFTUW9pBIncpzWSUnCWv3cPv/hDNYFJuoFcEjaudwS
6VYFBfVy5l5OYmRAltXF8l4Q55U73LnpLAQ5AE1wzSTFlkbV3YzIF++Ts6qnbLXvjp/TjbFrt5OR
26GJf7BxiYpjj04gPBzXZCtDv4mFSTARPzwi5bGjqYTsH69cwouXt57iAPMZ2b73RV5ReYq7a0QL
D5Hmgh7D+0pNko0k8nqxYSP/Lbbad/HloZgEsMJd+zhCvuUOZdqtyP9k+ulih/hKmD1NdNxP9vzb
vGZYcRyteT6Ap4Qp7xY1NL0gfo2HKJEIy/s4dGqqV4VwhU/tV/3JHShYMHObme2+3oRWtUxO7bYT
fuk0xz+xFqporDEhGwcHEDWTIMUVHk8+KsxYQaGCpH+YdkYNB1H8aoA/tszqEXyoeKqIXRFtTcXZ
iFvvBvICP+nbV+7Mkm99WzRZHG5ADDQD/1g43ctTFKaFs0bg7E7BiPOMWxJP0O/mL00mwnUL467j
k3HUeBqohB1oi9miqxyYOa+xo8ixXVmFY5ZOxAS0fU41yvncd7UTrhuiQ1e5OF1DpWgDK8I/yujK
GD0aua+42KN8qcG+JODyMywDEY8oQdOtlxWraIor8W8jLc8HWlGlWI8aN+VE0M1VwamFZmbRucLC
0b3tCc6z/BQEMXDjztSOIAHgXOZcPyPcbVHrYI2dIVUSjZRJj90qf3EwZFYGcBoYa4d9a8TiGqja
amkODZzTxIUH8JdhUTd85iSi0XGhPEhOmaozbAIzHvuAJLbZ/6Dy8E/8YPlG3J2Sv10hckONgEAU
DurPSYZRySD7znh/9Rd8Cu8f4oSDwaUW3F6LUQ5gsLLNNairYg9TIeLJpNIVZrV6aj/40nc5g7t7
7C5wxI/PAn1YeGzENbTGH9rb5FrqY9/FnLPD20sgyoihVcq7gJ/M1H90A6YNwB25Z+tIktV/+rLB
iNXo8gguBEzwnufXoapUkcDJPaU2YS9YzonCHQzOXUx+DAnHLxb0guKgS5SxmbCQniEOP1QQBawe
B8JIcqL7QQ7IxR+9VFYG00JJKnh71+h1XIkA2NRtU050FgH31kJBiKRnn1YjzEUczzJ9Igu5HREi
m3kHlCHvCVFVyMttKLzT2vcPS+U9weaYpHzXTC112ixBXWxYNmA3bp3+bYuZZTJ+Co45sdkTSLU+
hdj67zQEwf29W+UaxwHk46xAr1vlNN3wqRH60imuicxai0z4C4HSQduVaemsOMs+A5swgv0jJ9F1
Ewr1PNxK9oc9SOKlZZlFBZ1sEdtpQP6wi2orlXd2CsvuMbY1BVgCgAsMY7LSBfzZG4MOVuWwBrDJ
HBm6QVGsf7hOfCiU646hfZO4j6KqrhiTwDOhec/5c6wuBF4CUf4nMgZYYmC9fuV7YsbJqRjPcIGr
pi6ViMpfcVJYkNmlXpMEWhzCwE59EKYKudQe5Q8O1T2ZJA5ojGU3LA9ISFm9XUMGdv9Y+6zFsEAv
rwkAVc9hbbWubHJ9nF3PjT6L4URCM1SvFMapvHjIo1EGXZiZWKVe0vzxqEqJhEuEXtmSe/53bCfe
4m4lvpjP4Wh2pEKW9e5O97RLRKlr2Z1tWfu4sOUVbgops/cLbc9RU5H3uXnctBHA5sXtrt5YaPXt
LgeNe+H9ASYSxshtf9vDWKWsLuOrRWbL0gocN5U6fRuKkfCE3JlU3j3xRjdfscozMbHaCB0EnD5x
3seCq3o6wMOh6bT9gi/W5i546UlzC+IXTHfAhQf7H5x/LoN/0zc7s3cxSSsEKlYNXJTJ+Spxs9D2
QALgQ6dwUO3qysO4pOdeUUo54s411bRDEAEO01oM/vEQyNWNAmP9YOCCgakuj3MUvfSb74hXCqAV
X1NqlkY8jH1xpg8R3n2pmfJcXKuztIvWfyduXEQwDRJtwl1thnlP7aOk5b9sdb+vknE9f04dJLRy
ePpIkInJk0ikXHYQF0UfqHZ39OLC0cS+fK+iv26DZJE/LQRqU+4QXI04YyX1qzpgXUeA7u6GNHDB
Jfs7EFgqxJcrmCelrVbf9LWy4jjhC6ZgnYPhMNBFisbv/naJ2POePADvJhEMSmJ01YZ0Wto+YZzS
TpetdBVb7vWr2PvQbheEgrlSoI2Cg1bTtbzRTw/mwm6Qx4FNRnyCaTHUDu4legabTkg//RST+9Uc
SOB5X5Nqwvt6aA1q/gdkLwiK9XiR1QPAlE75GSxmD3Yq19Hkahk5EqMOuSCC5pFxQDr5f1oWess1
FnFQh3ItBeCVV6HeswSoY7BpvU/gWaW/Ogr9gAnadfv9yEWxXINbJVqigclOnMDkvGjI/I6/E41j
Og6u5PfDPRCF3ibvxbdr1a7uBrzID4fRPeG104ycq88zaZO59Il5IDPlgIJg7pLDGDUKrSjG5k8C
6ikNdwylzHCZG/0R1H6eTAXRSLYsD0u/+vglfg2N2lxGBvb9fwqo/PxMvytDj5mqSkL42RxcAkQx
SU9Y2sCSVj0bziMJkpT2zkvJu1+NROv0uwUhR4jEs/cGtDssLb6EfAXb9iX87+lZnov1PqZLEbvw
HklN/NVneMD7mvJth0OmdxtX5WUo+LcXCKvGGk7UaKDFUtJdkBbpp1LvNE2PNDlicuLq7NOhW1gh
iwPhz/i0NUiX9DBtkzkSKXZfiC3pky3KizrtWeYaJDUkwanwntb+mBR5a/FbUg2gy3KUFj16kHZ7
nAd0VMItL2o9XNZgfpaQoxYWnUNGSv+U5r4UGN2dlChj4rxjDHntk+nMG8FW30HqjpfO/SwzjGrC
WjL4OjuYnjxZHA4kx1TlrV1fEieSLP8HYnqcbdttJnXGfOX5pWLw+jTNZc6tp+wsBpLirMHM78Qs
6L92CWeyPoHOpH2X8XQ4c6h+aOcn/JW94xg7Ytu/QmeJnXqXwxfC7joI6F+ftOHYOf/cHb4Lchpw
HE83p49naLih58KfEG1RoFJUgNw3H7Beb2a5BAsyI+B1LXqYGlcBrenmvYiJEOLxo4dX2hcAgMTs
sIvgHLVwEXSmfhZMYLHJf5pWottL84dRh3oX+j1xsoh0p58tVZs9KXLtJx6rkwQ+5Dl7lenL++GL
4Z7w0DdAXhSc4OL/QplRLKqpXWggG5Oru6HpTBBictpcj4LggPj3jagCqCYid4cjKjUz+FZuZJeN
wn141aGzDiOAI7Bk5+0BjGq7NXnRAI2R+Nf/GBTbMiHczdBSPEYt/IL9jC16AToEJsmDhla9qJHs
TzDy7dNoZ8+gkjxgO/gP2WaCzV4BAlOZI5Rxmv/Z/howrq3v9L1sihCq9bCTAho5wsWUVYTVcv9X
1a7CWJvFBzPOwCm9w4ulxE4bjjPdRh2A6hjH/Fzv6Q21vQuXv5rOBZE5HdxH77hYSVW7C9+hO0Dc
g6i8+LtR9WyX4x7zgUKcZsfHImBASuri0yyix0l+lJd6vrnGTjQSshJHdGlXPvpMo+IRHWT1imQJ
grdhKslFBzxJzYham9ceBzNW+h+GlD4tBlgK5zWeMPqigLFPEgQJQka42NoVstzFb7QQh0ryPgYj
VW+0NNY7QjPsjQC3Q1mPkek+vUS/6+XgzMNN9HwdNRfuI0qNe6IO8cE1QvSMyT2CS/5Qh2vTKkMr
moQx+BOfsT/Cy/E8ithVOD4SBYIaEZAZmqCzBh5uf0kY/DbrSVZTJsWy1Z3aepXXgROmcwJCPhEe
f0qvtzyhCUfrI+X9dbi135RzH9e4Hsy90jtbUeUbZOZUsfJgsWvzfL57u8nTtEenTX/kz67TmhOF
Ja2Xx9zejDskeu0kNZDUJqzNz3PAWZ6zv9Uu56UkNUjkGw4HbiX6AbBsjJ2q21MAzvgrWSE2f+OQ
j/ouIFrfVBnw45W3o2Y4lh1RRxSyNHJ4l39d7Z/nkj/qlDux1mT7vB0+zpa+PnpYGhFqP+LNvcNc
3L8qcrp5FtPU9yGXtZVINXknH0GsI//3FvbayDfVyh4u4Naeds4cLSw1m8BYNKe6y9TJDsSuMriC
cUthCLrgpV6iLBaTRJq/896CnrSsa8bo++MNUqgHJqyvYP2ICzXnSuyg2LcwUMAc+UxEHY7Yutk7
MCeB8FSIypq7KymoCoWrq5WH/wp5uKednn78ZeSObkbIUYy548antu1A/rUzgN/qWXout8EeRyow
AycEGzMERLtt5BTFjt6QAjK3be3Xvp4Fr/K+Ph8ANxcrwSTDT4vzSiZA05AgzQk7Y7iZNKOa245w
/eQ/D39kl9a4fClxHYITjDYt34kXahODZ+1WZC26g5yaVDGWfQqvZkOubAJhafRiegOP3O4YIkUJ
lbHCHIpr8T0uABo+hBLGIdf5W2qB8iExfvw+f2jBM2GHwqndy5e87OowVfAlw2gF1OtT2LEVP5lw
zWgznzTxOFry8SdoBEEbAZQAKVD1dtk5vPMy9z4uz79CO6VBhTR6NgQvwBzGmprYQXx5NVXsKGKn
vpKQ37zhmHcUqt9n0607c+nvF10lAXObzNWovDURivwHaofSErVp617ANikiwqzao/zTsnK4CkwB
D6G2Akv+YArAP7kMJVIyLw+F4mGQRoMtyG05NN3nc3E80YvOqzRw5VOQiZkK97IkcGK1OYhNK9K9
Dh79FTTUhkeF1i8Yvho4EHUXQUTexeeRgTpiwougYXwcJiHSBiL0T09NqRBa0LPokKeTUxNoyoFs
1wBiFdrNhR38fjlaEvq1F0wuNxUD2+1W9GmhvrsEqa1LI8u4YV1N1EarjqSviS5bv0tQcwJnEQhK
18pM+l4NEGHI8dLT7ZsxEG4Zo6WblSMrCvkRrDKygUIgHZNlszE00k3mvAbTCk2KcGwCngj/ohp/
Zs5xm9T87d4/ORQhBj1oh1XheCuroX+uaPp06awjb101FsekWEpOHc39LMQE54/Vwo62z71kxEkZ
XrdWy/5i+ReDJwUmJkAx3fqvEY5eRXYILrQwy20GcwFG83klTuOWh1aM8KQvJMEgzccKUS09GpY6
609J/YiQnjb0ER/Qc+9Cfg/xHgORHAEMCzYt9qdS1nDOnMCTUzTBfWuyyIaF9hmoilxW9++XkhZf
/WJIgpd93c5K6oAHqVZZNLbK+hK69BlIyAIyWq1tO/5pMG64lAldfKaXdaXse8QCiaDrF/Wass9V
KYqr3ua/jrKV10xFyiWxQ+ZIJiIuypaMgWYY4qOZc7jBG6b7kp6Knc2R+USR1DZFYb6KK0/GxfRy
kDGBnOPIERiutqd/laZbpeeCw3lQ2sRF/l6Mb6VhYK+1grPIUjuUw5zP5PSkF1nvBjwPdXl0xdGh
uXRPSEKjb+qbvgNeuCZO2t//kmoINVCYdr3juzBt1qSaV+2CtMuLb7imBjTdVgPAvCJlVVGpB38M
iXgTZH7RVV59VS+9lZ4GgalvtlfF9siV/XlV43az2QpNktweuIOWeSE1TidbtFnDqXLIVUxqm259
wwfP60dbMfKvpfLZUw4OpVYF1+Q86PAEw02T0MsbxwZGRY47rxep0s2x/QpBlW5wLTr1gA2n61RM
3LGdlqdtenKWkmuaUrqub8w/QCL33eGpcNAZB6i4pn0C3IF40oPpnBeC8GbpDpVQI+oLSE/0Pusq
giY/SRFKfFH1KqZbuHxtzy4fNjc/LGttydG/QkbedFioVyze7nYpCQTFPrfrPVTo2k8SsHCkZDjW
Pr9Mre/mj4njDQXft5JiigYwf/v/VeWLAZmVh6KcenjlqtWUZwKbvdHN65GUkBKLQvqLErfxZFYf
T747jOfMrHMr/Dk+JjgYUx1+1mWcfVlZFrwcs5tWEiOp1LUC8ZaGKJzZwb+Qu7YKurSVrzoX7oGS
NEV+0T2vZh9BnhItv4JlBqVti+x6OKcAF1iKWCOFAuhuy1xHWjnr5sGTntVc7gLUGZIEQU7WKize
fveBb1hd1SgeSkSCHXtlX4xoZ8xv5WwjFUK8Bc+wVySmIkcObMx/4wvNUJPoekmEHHZzJw4Gm0a7
09QmSYM3iuZF9wBvs74ip30/Juri/d3MNKJ86CX+idNENJkNlSHMx+EwnHJMLd2r9lVCZpFzCL2h
3DpQhjM2oLa9fQzr7QZy1bjcAvf0h+Ok5tyOa0jv8LwH3atTotjamcYeKDNFVMtuJZ81cWPGo2e5
R7Dh9aL5pddwScLqMq1o+omvfTOK4eMQqaZZffjQHySTsreZwy8xp1/BGrSo2682wejWERirOuzk
xsenuC3GnqFioEcRNkKHZMZ9IHfZAb5eQ023jF3W3guqjJ4JwIsIE0nY455vJ59wNQR9T+JxQxW7
wAYcwzFo9UIEO6FTVtS1YtsZHlDz0WNrJeR15zqLtFrUBYVF/c+wOKV211CAKy0oVvhAsw8UbPWs
AxTs1x9KtWHPzM/CwUJ7tfbWyX18PcNpP06kY64QHQn/BGTfEW2N1gaz6ieUidJHUM3+R49/OfVu
PnEl0F2kmyTzjDiB1SmPoNXJi4hZkmsDYmhSoRMwkRQQ053t9Qy/+j2LUjAwGzGpS7/kdFlWZSsg
0B3nhxW8w0pMyPWPxi0aJsVQAiT/TOPNFtko2nPrZoI2bbFV3NMn7xvy8N24rXY5yGFQkIams6Bx
Egw9giFgC41DiXfjXK2OIB/R8YtCB4XMrYxy5JTuJbWe/kyjQMKdFsZZ3G3TjvLGiE6N7qdLEqFY
2Qx3k2+OFBjV8ukViv+0i6MP9wWDqzRVwfSYNugSKTpXjgHtJ6Xd0jxTDeEGN2r0GU/Ngof8ri7A
LrK/QlB4not9+bNBbvBnn1GFSUD7Jurr+xaO/a3zjcIiddu7CynX7OHWBhmBDcYQzfeE76bUAhZr
UefsGMnYXispICV0/MAWeHvmyQ5qJjiCFOVM3wAY4O1hjKqzU46IEhKSOx2DfICwcKmIbc5HB423
o0qy7w92aqMwd0Gszq92QA61ZqFqoZdkf/sfCPKBUonmZ+9YtDPVd4zxSEzJaV1ufEdvDIsT8sxc
bAH+QqnioFPdZMjM35wA4EHoowVw0g6vZFaj64oLwf5OaYljgGA7a30fNBGbohN/hmgtNbGo4AyJ
JV44pY/CB8etQ+a88wauX+Nd3DsL2xCS04BqWgg5ZijKklWhjy5xNrp/fXkEfwvXr+nP/Bf3aXGO
V3ePBot/DPEM8is4r/bAK19QSrSN+ePOuADFfVlEajVjaFPEYg2dNI+ebtQZT2UZIBnbO/JFbUNr
0ia64FUt4zYL2sC9WXhhEf9ZKBoqNgsU8Zmbwa/YRPcPbasEiAFdtM1dODCwKblcSecnmf57Nhp0
dM4Faq5RdoUtoO21pP92+l+ul+gcerqf5JyoQNZtNP5FpyqXRgwPIdRJa+MrgLq2/gprMR/A7JNs
0m7k5ZmJAllQnzlJx2YAdpO05eyESQQVjcuDGlmrsA0qjVywG4JJD0nbS3fcesozfywyFmMUC7Yl
mQGBO1lRe98pd99366juiSJuTz5OJYMrVi3EJN7L0trJS/p0AwNp8HRijlzd/q6gC/nLeDyLVtK5
mEu7iokOahbTiiked6ednqD5ek665hGhpLvVHSeHiYm8G60kMHqc2LlgettsXxOFJoFyI+2LFTKe
j19DQs7OjO8wjhCH5AVmLmyjnaBbyH5lwbTbKemfS0qPrTrHVd+6wMdmhtg1KYpLdKI5LgzNBWya
B1VhWAddeIEzx+jH/lzAtWigYeyf7BgRCehkDtfXKWvnTnBw0c24VXrwG/lbzHqKqrPQDJ9xjxGJ
2V2FJRQrr2IINVsOKr5t1iPtjd9cgbaZyDsxJygkOsqDz/8b5AIs4c1mlFf1lgjhD+QK9l4FxOvn
FSs5HRv8dZyZ5IUYeiscsP795T1T705rTh2blHQAyoK2cmW0E8S1uJJN31BTt1rxoZzfQSQ5jcQy
LoL/ALt98pLzFroZofZrVUbQJxL2xYnB94+C3llkh6JE41Tj1o6bjzJrCBFrrDfCdlLibBBj54JH
+G63gvfWiMQ4X851rnjqrsab2esNAQhF0REflQ4p3juu/+6F45uNMa7HfGuV/I5KA84A/KloBHXH
0OAPe1q21F8hSOo5WgmRNWc2g58lSyxS6YkbdiFeqe0YmSsXcVg4tpM1ZRZLAliApzZR1d121XSp
2ekGk7DeNOQPaRuPPuS64cwrpjdfk16rZPP3SyrxsYZT+sbKpiUsb/3Vyi3HlCF3dWd5CXc2W5s7
tnySKVKA3YEwwnVYuJDbhjTM5yO1ftVgFDN7l717lIc7UnDLeU/1ohq5jZnGQHWqLp6BpksltdYh
q5mdJ3nYUQERuWzpF3qki77uUZouYWyaKznc+yNknLAxEMd1kcA7KtcrAuFejB2g2lYH+m6c/zkN
qFYuixjlm8n48KOchh3WDYQUBqy18YIHSk3X9R8oqvbThP/33/40767DTaMnO7PWbYixW2/cQS18
EJWJdMpLx7ejAVwgkBdPa2+U+hrVj93JwYH5RKEDbjykowjpMySWxdvBDpJrTYFsSJVHIUWGxbto
N9+blt5PfIEthnW7tlyEhHi9fHxrCpvE+yGH/RWMTJOOmRllAAd+y+2aqRxs99d344m1tU7GaC0P
AOP/FfQK9W422xZewibZeVHoUG43PMhjjbyZOB7c+sDGheAlsysP354RXTfi8ISfME2rGfQzdqpa
IgbgBnApy+mV9mlJSGMQL1ul0XHcrfV031bYIiAATJMlBtQp12EO7rRXqHlNasqKVnbSFfXfjseP
8MrjrgrfNiFlv96FUbSwMZQGwkqWz7BfnHIvO/jv6YF6KKzzXG/jyNlGKvOlEsU6n21zwUrbTSdh
qaQiQrtMvDVrqluBea3axjJJPs0cpwT8RKN+LO1t8NPIMcsGETZm2X7+VqlsEAgq/Zax44F3xJtO
5oQ3439EPPPce3rilIXTlQSDI6yGCrqefxje0ktPFX9o3BaEjWWdQ6X1kxAkYnB4w21pz6XuCOT9
BG8kUqqxk4dZR1Zy/nzJdmjowK8nxGwhXxTxTFXwlm/z5DbZrYtq6e5cc/X3A5auhILv7xHjVAPc
emzhlOtYXiz89Dmf62ZYoNsdFxynCIASpzxpor1MzEHfmcq0W3PFApk3iIjq1B3fEdDXA9Wre239
awtpMoisP5jcgGd1sm+gjkqEYkjnUInar2mWN1WNPVDpcEctbxz9KXOxX48wfFg2pRwwQMijrklD
LaOcG0JdR9sGaKSJgdQw45DiWUsPADmwmPtxGWDB6pmPWAHjQgYNwxw2Fwg06NeJlSKxJwcMnuZM
9Ah2NsL27rhVunYauFmgx1nRhwqOFYPMvcYRW90OZW1aVfaQ7e0MCTJ9JNkpnyVDGHuLDcoVeyeB
zX8D8B9Qf1iPKxH2Dl1PJ0HEGuunfMpjEzn6wrzEiEaaR0pazMJ18tOpjDe9eU3BStsW7yNj4o26
5mRttDaD8cvwW5fc9DkA/xRXHhBxNOJQzpg+i1Fd2kmhvpjakiOP93o7jDSDq+HDA49UkhSkUlkT
qrgUXJGDIQ3VZ4VuEIt5tRbIhuzCfsldzUlmhqiMoKT23nqRDvsSP//Zlp/7qK2sfqgcVEawe8PC
LhVQskbGiIkaG7OwfxToRhEW1rCUwh4GEmKFjUjGlKOiD1JS4P7GTln0dBIW7qFqgtf2g08hbhkI
yF9W6gRZNOr4XrSqcnu2chp3GuKH6eBMg/jSppNsTo045w8xg0aRgGzD3PM+cpI1Kg0LAyCuUQoQ
B5GSbfUvNA0EVgOrdtAItCvXWoA9t+brm3UPhkEFsJjlYihnwRqnvzCq/s8hPLQHNg4tvXKLSwbz
uoh63WLj4Uhkv7TMU0OVO1NN3qrgUC3UsjufG0X1TLlifpfo+XsWMRLe/mvpTgv7YaeZZU9Ur8gb
waDhG1BnHq/H8URipmUQeq3T5bWi4XngLF9PKChRCfiP/Pb0g8qW48XeUrYJw6Z7HccwFvcE+MgJ
soGZMqftosUYVVzAA/hf9FTnk2klTjwe4vGmgFGllC6piDNa86KTDDH1/mG/rWHA91an5tbzVEnJ
Hz0Qe95suMc8vex4BeoyMzsKgI2yxUbomaxLwP2uk1+b53qcTM95IJljBL5qvxcBLkY9jPdT2GaR
WhB/y95PoyoDtjFcObQJkFwOqwj0Ej6DYkQkzhBp3G4828nvmnHP5u030wnV5TcY12kYLJoeCfqu
ubWKf/CITVg0pniiMf08BJuAXpuPF1O6/5sAF1a53H/uZlVzeHVM6ElLwoF6PBbT2KPBQBEVi6W/
K7o9vzYzBItAiXFMHVB3t/4akUlzCif4qNFVZ7n4wM/ze/prX93OUozQ/symLzZTMMRb2t2DKOfu
9VaZUYAqwdxVqxS2ary3vSH1miXsESqFf7CWtIcnIG2ASWtndwLIql8KbclAp1El3DHPGq5AX9+J
il9wUHMITlptoQLWceJMekgJVaK/AjWTbIEn+TEdgJiEfbRewyP3EqBZIPxEKRFql1mTbczfesuc
KiT6pJAtlsCijkfYaVPHTUv+BbYFfhX0SD4B8VVWOlCfstZk4ulS8iXNCVybnBNWdz+hofQpwP2N
3i/YV2MRC05ptRCRwQjESUc/45Ws2MZVxQdficMHBqnGryYOssHzATDnjE8N1PpRuDr8RjBNNJaz
F8sB9j3fPX7dWQJ7FhXVb4T8eCgk4HZQ662C/TFrA9JVtvXMANFBpjK8ZKRksvW30Std3vakFAM7
U/STLC0xB1ZdebRjnazh+LWm2VdBIR9GDDzPNnliAD9r4MyKGGRluH6rz0i/FORc4ihldQLT1if+
n3beMvBaWc+Ir0Fl2RChnmK9IcQNzAA7s2engS08qPRv4UL5wRvMqOtMzh4/cdv62kY8Ii4NG7N9
SoRIk/5Qx1I745772BzcqfOdt+SwNZ+fNGIDTtVDBoZeqyGThzstVjCld1XGBx6JcU8rMI8KG0C8
3jTDg78V+ZB+qTbKcl8wwxngqAEvwkyQ01xfppy1oKKkiFNb6Du5o88w1q73DH7iAr5sDED96mjC
joZEWRAKqShdc+rzExpS2PVNL/MZ316k+Nox3+92fmhgX6BiEHLsUpytiZP0MnhpdGpqYB77iydG
eUeB575duBOScwBPYls7CKUsuqBK97atJV2e1EDPVcr5sJigCnauN28si4gbTQM8hUozVs9xGHC8
29+SbTztxopW3ItFjvvvlxqUCC4v5tyhhoQQYc+OAxQ+evFbgdd3QuY0gYcNH644F+j1Rmnu18MD
6pfVxYv/6gCpie94q3S/T3++MKgCS0sHuf3jProFdnRUJpDCO3CmGxWjnS6Prw22IlVuuhPPx/1z
VRwMAoos2ACXcDaD+g9gzG1YYeG9MvbAI2duoI1DU7/PMA7fr+dIqK2F35/cCYjzQoNnrWvZ8CaF
FrA2pDv5rluD13Nq93U4sOLlAHMYnYfhvXXNrGjgwMTNF9u2uUbULlxQ+GXNrpu3Hpt35TCnJ+ce
/NoEGhL3wE3dBVPbBYnVpypWL4Xife3IOrKJmMTR6Om5EZGNLzlC84cuKik4JxnG95IEt1/kfBk/
NNo1AJtlP0tx1V/RdZqQll4L2HUmbk2siWlZ9h2okx++3zMyZXRLbXP1EsTAtOdYXiNitAEuYv/o
d8NuZJISF0refX7sCBOAuj12lyNa1RM3g3CAYepCvuAwKq60xC8Legyf2klfQTiZVSBaqUw8DwxB
y9Vu9qqPIfz9skXQnQhgMhMyeWwdOVhUi9NuXloQFv2Qh+/siZJyqrge/siOL+xfNZ0l5UcTcYet
1iOohyZT+fs3yr6v35k/J4ry5Cmap9+nUzR5YX+ynIrQo1mYZixDwg1jfXcemQ62amnHqqzHRI64
6okycPzIyKLYu7+2jhXK+G/A/VQzvkppl8A8Yg7+Y3weIPxUrCLu7uz+9Y50AaFw5ah5B6dvPFMO
RCFdt8Hlgd/YCUEYPhWV5SOVkdwL376jNi7oZxaZcLd0QEmVtTsLQWbfpgAWKDQdPYcTh3EQQvzl
ac6SQ1NSJwuGujx85vzKkJ3AVZNWUYtoSfI2Y8bsPGvXnHgcnDxKA748pyxkDiAze53TD49nb2Cu
XID7Bo8FKJJ3U9Z5GuTpHcuzP/jQiTJx9SmXqr2vg6nBH6vMbJL7/IZ6i1JMYfmtbkd+WLVzrB14
MVjylGGiMZWKWjwYPKBgxAYzmV2KPkcSjaIz7HdSKrl9A8O6/BMyqvwEC/acoZnZCioyGU5tQUuV
6LZcskvQHqzV0UGYb6W48wf14FsJE6gHD2hswQIE64sH2MO4fjTpcAmRfZfjsKnj9nrtazIEGg3Z
Uz/YdNVWB69+Cl7LND1F9OgBS/WWbOywPXOqvplqs2axLXhfa7uiOWYxatVgs5iKG+5CQ4KO8ZZ6
LpJ0gQeSjtyQSq4fJVEe+MFcxnTP/zTc3jtwwsFV92hyBLHYqHi8LNveKowgIhymz/U7w5n0hXvn
QbX33Qsf0NcByndIoAklKtUp4kPY4EwkjiLLIRk2V3pqcg4DScOItia9pi1kjo0REH6SRFUwyys0
h8C1FEPcij+oAMWqeXEaT9fw1umF32InrUfVjlCNGKT8kMMdnhNuvzQVKKuPqXF8avA6vR27lv3Y
Ba8tLN6s2TbtouRVt4juAyuRkccY6IxeD32XVlR2Dba6K7Lh1dR5xDZwYwky8JzbVPZPbLWosBur
SlBM331DkaXtKXyqyKlRoKK2QPYwKuDf0J+ANpw6ZNPhFqM8nyhdvjO/wcGB+Bzu8ti0P6SfKSl9
OuiRK8lSqkbeFNO4H//YC63Ef1sVEO7pAJ3JEEE3w/mn3W6+uH05hyef7nBcnfOq5CEA2S2BRoYB
VBRW25XgC/nztEV1/MZStMNIVCY8C1H4O3MMw8uedZ8Cra4wbQyf2hbWAMSUhH5A1No8LLQxqfDJ
KRlGPGGSSNh4XuAwb6U3nhJC/PHkVpgCDLIVf+XMfZZObA0byl558EHSuiNqS7ruQFJCBh+GdE5u
zMeX6yeBdjNicVnvP1+YJW2Zt5vHYB3q6KFwm8wCBQrqHbnEusJzmban97gt0ouZLo/KLi3g/RcN
XTPYij3PM1X/yBi681yB9gXg3P4I+3/WDwkRwyFkco3FQknzKx/OnIn3Ugnda2jJ7VnP8hZG0PBF
onPJXMVCgezTmjXQi+Qu/96uDe0F6WVLgjQ/ZyHEiDQEbikMttTtRzI6eVVg9Ivi/qLK6JTk0vWT
Fl4AmuRQtVjEMqYU/daLZVA+HNBIN7uiJtEOc6LFJMkUO97OBwwCF6yJN6ZvTYlUg2d5PagAxq0T
tkkDirQLvGRIZ6iKiVHvA8N1IDl+l8vyEy4oXE0hydPNTlXk6V4/kELdYh/21cQQIoRVUsnmKj5e
H3F7Bzuo5D0yEQmaaOIMTnG8NRLEjTxEzlO4aqRoA+2eo16diCsV+vYvcj3QmhS71zGLqHHQpwJT
hPlKb6TKCUX30XF5HH5apMF3QW/gEEaQXeBfCSjnqcPIEn2l8eYSjiCZILQUTHIELfg/GoRbd6rc
TvGywQnuJIthz00zcPB/DsQDvXSeJqWERa5bH44wk2s81Hs87sHmDgwszFbH+qf12yju9jaFo80y
WGLWSB+I3D6xmo1kHlXJPtxaY+OO4A9LST3HAN2Jzu6gQO7PvZ65bqnPEnU3mLh/WnU9bwp63myE
OyPz6LjavfV39acv9U646yxWmXJeu0DL1Q3nMAQ9A9+tSGgXtw2QmNQunFqNRe3nWB1E08aUAAVV
ZnPKgBODzfvpB5x1pO567yqhjTtP/6IdTUA3winrxTMxQHRaippuubsTLoVxgZgKXElQQROoHKoe
aAYQm7Hb27QLhu8tf8ac4mwXOtgpNTjXWRNQ6GqSM+DnavJsVwOXacuYL4RtnsxDt7B19SVeV0wn
NPMcFMnHogE4l6HqEPI5CSKh7/gG3Jf41WYnzmbJfeboHuLE1S/VhlwOutlrGVdpv03fq9k7OrRT
6QWnI5lFWDaW2dLMbhipqMJqaK85Xhanw4U6pGM1ekaSbAmbZENoDBByT/4eQFzmE745sAtuik5x
BZrHGNF1LpB6sB8lCIag7c/jQ7PoeNf3yVcNhvDoB8lxwgfvnpDMly824s7LhC2qaggVvjX0awq+
fYsAN1QQvbg5xIo2rewqkPhrVEAntOmunxPlTjasr0Rc5sL2cIOpQWdWVP/twZ80jVux2LC8MMZx
skeNsg304JzIqlUJYaU9QOFhdb4zzK0QOkh9ehvcgju15T1W7jNy7BAETqWffTDwu634b7TwmdI4
0+qQeWB8sAATT1/1hKNJZ5hR9Jvi4C6WragdfBosiG6RIC4PogWI7gxXpagJz/bgMRwmLANnIpfz
QUJWBxpOWD2PC1JACA8bbb7eY6oUUYe1KS4pKY20cz/2gV102BYCfxVx6XXG8LA7aPpUqhCfWG+M
inrP4j3TXEy4F5eI7yXQyIUQGxfM8XGCxVnJW8FxEqhVVpqXWxPMGBzRBIqVrMZbQlT9xs3KA2iG
ONkVh8ohL039LRdQFu6PLb18xlUbEch7CbIeH1t5+P+K44Fo6DclhXrX2rGOFm6FKcZN5WujfqPf
9ycro/S2ctCatH0Z43dOlkn3ScsrntMPkzVdHBnP6ynWjT6p/8jnLCOuWdGGwIGhnQ1tNTuDepTl
dfXHW3UeOcVGBWPgkXlYTp/u6npIQpbvKUp/dgFWvgE5o+vHl1yUIWvIFKpUzWsOextRHBPeA30t
NiRi4rsd7LxEZvxi6YTmkxqnaOWAhe3PEceeodio+5PDJ+rIsg0H2YK+oyoyAph+12V9O3SkkAgW
cTfFrxINFU6LGsyYq06nFOsCbjwIw4tYYV/Uc/vXY86UqZr6/Wp6Vl4p3LsCSneYDbhTJESiVsBE
+RFWDnbYhtwxGzp27qSy50/wKpPmqBfAsakYPhIUA00BL4LjyYkE+62roD44ZN47TiDn6nLDFpuG
Wq0YxRL7LRKvYzRAncZtKdIm5Mbt0SdhOuuX7PcuykD7A8h2J2lozM1Em7SZCriufXLattjerCxr
/0DXNe+xoRRuGSzBbl1EW0ItD5jmILNvhYfCXDq52KOYkKdtQumbdiNNCgjF8zVWo37w4FYTH6UM
ZJiltrSkqeKsU/ThLRDFfli+BHoCr1dPWwTZHEDStUx8j/tcsoqMWkldVLIMmV4j+0Cppee6KvmA
eUhxgD25dXUGLGchhRUZP31mavAbYD/c/AfdtosIu5QzXA8rhUrNeyWtLEIRC7e5sLFvtUPd9dwh
aVTve3WiYrg7R2hPZai1YhtC3uDk+LR5OIqed4oISjNR8mtdegNaE7PM6CnnvOQDqgJAVoSONzZm
KnerYL3xeVSG+cDb0aCEDKmJ93C+eEkJ8X6EMV+GdOOlfwatGZaW7gA807ViIqnXsgvNX4QDkdFa
s+CLec4mOHM2MWOYEh9vN5kr6TPACxIILV9Ekv/oW718NCwEwMsKgorAZxk9YhACilmqYBS242/J
/M1stSoGM9jK20QPBzddpuPG9NYsFAKRx/Ae/00EGCuNdAS2E61J+i7IOU6SyE6+QO/CPhfC5lBB
HA9NB8iSNBv4LdTTrdQJ81kzuTSkaRGJJmZr2KZVzO51mmHMc/kkLHMRRgsChNB5ww1A1R1gEbIt
lbPt60OMfoFZW9dluoz9S9yvnwFMrmW7SnI+2L/SBImE4+16lnHurnpTEp6Ir+ZJyB9ZA25UQSJq
fzcu6tN7QWwDn16vOgX61IFCqcjGzVG5M9RVkL4127nBEBYqFVvfvH1X1TcBClLjYXZYLST5DJkf
4qKhFW/GQH2BCOsm/d0cn/Bvn0zdnX4vgQliBXi94IHU0+JvVcv+oOZisHRS+naAdXYMviFJSEnH
MCMJk7XtkMwQBx4zjksmhsU0IODbqkwZQ3vIhOTCKNSI6KLDZPPAlUS5t9jt7rrDBCGAtAGXgkhf
QXIjg66Qru6HJN8BTI08qPHi5XX2dm87cIBUyTfot6tWLplQMJ5CeBmaVdVcOltwSxJVaWbJGjum
i5Kp+x3J0X9T4bKuHdt6tL3nvmF2CKx6Tr4jkVpwgBwudISSkRp32UEk/JponltJwzHzFU7GvvVC
nTTASS/rPf5AnZMxjjPVIdaOgFVj9Ck2Tlbi8IZN1INuE5tNLv42Ox/AN42o1BWp2GSnHoEur9Vx
zmG9ojp1/kIQR/r7Uv5AcuT+7mBZ37U10DHy0sGsGdkBdCUnyXXTQfywe1qnFEF7h/HK70D9pwYc
rSTQSQ939wlt280xKyiMODASrPJu4dSK2Je83TzB58xpZ/sCvs8JBP4UBqiART3MMYYvPFxrHO7N
F3JkkzKymYCt0YlAfkZ0TvwyRDBQXJkLJN8JfRa9efTQ/1KhEh+73uVH6Uvy+MFG1GrUCgAU4641
GKSB2k/BAWyf44UV4U/avDtJcEs+tl0wMux0U5JFAjoLWbfCxH6WhMmX4oLLTzyypl0sX5FLhedW
u+mPGyJdLAK/TP4oNlG24v+j96n/Ivi6ysQ/sMW4kHElWJbAwRVgQ8mkBAfyHT0nUJbxE7pfjE6e
SiZO1BBkdlqfjn7J5G6XQa7zsBFVuv2YoOn7f4iN3BMkdgND1axKE9j7uwmxnChrK/1oBKlT5CNM
8+xoN5vouuzz3AMwzPzPcqOLspWe12x1y2P9mayNUdP/LsJIvk/OevVMAWWK+jeXPbhxSQ8z77Iq
73gx5zL1Df91u6uBUDAx2hUilV+UJkJlMumrWQi+Ds+w9g19pYj/9Ud2uJcK0cxH7GJxxwFOmEOw
zf3h4LyX0j0uvaRDaC6+2QJsL5brg6sCGyl71ptXpLt2TArj9V6PCyy5zcAl5pA82yNTp7bL6QRF
BalZsbr3UxchiEInzZtFYDfu9y7WLYuVonve/kwiAeIifiP7RNipkCHhp7FSmQHH5wNnBcnsFf9a
3E7lbrc7zLaMpMCGDxBVmZhmbF1TcIB6BeEJM/JyieJdqhShetDNxyU3b3qVlLRSElLQ3IrsyaKc
zYx2ERMVILpfeDjO78loRp7JiuMGmE257bZDpEc/pdYcBXKwvbPF8Fz1Rv/kvR3JVus3CV8km/IC
h3TKo8Zhp0x3DVxwzyae3zPRTdMmTeqMrkCRCrIjcRz47QOiJck+rKve9euAZoxgTU/uMHptJ1g7
RaJ/HOck9px5GT5hqmosSojLUjgt9w4gk3zfxVypG4ATD2BFUFpKYGGlGbDJcsFXG2b4G1lZLc/m
I+IAcszhO6QfytJuL7t5hxDUbfSamBoyx63xB7a/JX9KvzoIOVodTtwteVQdeIdWNQvBw3dgKUIp
RoJjRTpWOvEjxrDbIQX3zexZpCMsRYvRcuZ3gK27KAMxUqzqSZiwYSYgM5qPwH6YBcW4dbt9ot5Z
hmEJtVIZ8KVt0IjYmLwHAJaLZ/KCEH8HIMWdtZwWT/HmaxvKMn9MdzeGV3zuWGgvXWP2Uk4L+5HH
CmpqoKXJFfMCn4esJiUNI+8bFyKheT0/7L+Gj2teleu1FtMncyv4QL+WvZfFOEw5fKQf+ko7zw2z
NzJzdwu6uhDFC8aIkI9qiuwZwz+l7cD9unerDQ3iw8UoJ3RyPUYs5fRJVm+J4TEqElCuSBNrLn5b
4U23O/oKlO6VuehnzCO3KsUQ78Sm4NF1WSvx3GMSq/uKVZc0F+PXVdA4fexR/4T5s/rod7vDbOgs
drvW7n6bDYhl+2z/iWcGLDiHADoewaZ/l1mgTeQw9XNkF9xgQYJePXh/Amni7gU/Ej7rp4M5bp+1
OStJ3JLO/Hc9Wi0MXhQqVLfgL/gmeZ4ojQfxAkTV6BOThREmb5GAAPW3/tEeKfa/WNpO21DeTm+L
Vxeh5eqnS9My3zGvUCkB0sQ2CAQCPxj7Yy8QSpFzhP/JyFKXgteDhNhIxhrHxfIGN7mAJ51I0oad
3srbSvOOuSidaxiTX3E4UqHjayX2M5+K1ftw3iPkzveGWodNekslakO9jsITwKgqf1QKIa4Mtc5Q
iwaelOY7IkPl/fsYTo8Em3dX8Z7bjJPGTSFOoiOLP5XVSu4AhL3VQSwzlHPsmqwXA/NctWmtyUrR
/8DgwVuse5F29w9hGPkv8r9vLPmZpQ4FSAT1XffY2nPixojwvAwvpZr+w6oDt5BTqRCNwALhW04C
LJvtQUZKE8tN+5CPdP1O5wRI8c/ee5IMYWcS8ltioLjLlG1J5Fhg5JL8im3hAbJdIsUBOGR40y8p
Pj8WIcp+YcdPz440L7ZXLD5RShcmhMhrbw1bU4b9RGom8Lv9DC9J/8N4tprDO692TflWH2MmH5jV
3izSEuQ6kKExFTJTyK/rBBLLQjJf1pccjUA0ZErO2BPUOXGbrizYKGW2ULa33RM4IyWdPi/5ZX6r
lTbh7CRbHK5kQgTSUML1ysY9ylRk5XwSKqDaUjD3KzgqGjgMhbYgn2nPvKaBffK292wVnHBwChnu
vx44eJazd3juTycB4HtdI8pc279HVN0iKAiYjOGwm0yGstSVL1mycACjCYuKw2HV81eIKfCNA74B
NnYB9Q36V1acwpolyb9y+HRuE0ZoHt6l2qLXutfsVz+4+036aYcgzXUxBCbPMRTmk3jJzijNViVx
vs8AEsu7uyBHmRowkf6rz09sfwb6bX4U+l5vpZDZzpfwXQMwUl+ZPmIK7D0RephDiZThTmeN0LIi
XTKAh8oKpB9HQ2uVwNy492kFyumqnUCYanz4pUvhyEyNxRJVUXHqt3B58JD2VG7ob7/RKoer6L9Y
wR6w7VgImplXVbhAWIXiCsslM8KVlUONNAkjqgHijeIMOqgmndryjibbaI607gLOeKWpA2yORRU7
cyJc4++jl1ERQHViaepIPlvQGt4RtRn4GNmJKcNCKHynEO69bV0/pR/9QUrRUC6P7XkFYNq85839
szLw0foNTEyGazXvO4/YA57J4pAzfFLWuXZKXrNjMtHc/8HRiFEcRUbmqRojH99nh4d8DCSLXEWl
AvrH9wixVYkF+UVm9zFu90mdQ/lhA72ymvSnje16L9OuS64/TDr/+34RPQTSF6mptuYosQp3NaiE
9cQAayDztz+RYSDIuC5nnw9Ax0fl1gFZB07Lyo1t0B9ESU9LSLFSyoXnt1o2MiqBSsh8+XO7oInd
5Is/wAOWvoCa4+kZEcCMw+DKyl2SemE/rIpOchKMExmdHXHCGXXVTm3z1o4Ne6iyn5wnphNeFe2U
QhV5JOwRn/O30ch+OKNw+GrecMt5tLzORbqPdGVKjOk/m30viCAg2mgP8CgU2rXgrXH8a1NpDOrt
EhITBEKVc/v31icoZEp8I4dVOISvgCf3nRg9RjFelqjKalNXgGkrBq1AMNlq6SZhQLZ0AMG/4IEP
f2N78tx9A+70rqN6q6CLtqjDV5N218RBnYLn+45NE61vEFwSWgRLtWvdtNS7KgZKlncqAI3gt/pI
KNrPuIIG1TMmXljhN+mvxFS8W2aJmPrglMhaVRBQtZgGSInTt2TEjS5s2ubHAngT61zKipKvRW43
y/Y0Kmt5YcEKfrZ1iE0a9xy6kXaqmwr+W6gaw6OqYhFx50BEVPL47Okj/KjPVjCQfNiZ9ttj57eN
PigyOWwg4n3oSW7+PR0v5H8wX60NyUz690H0NgTZYTIJS7tzp0KCUr7OKMJQrDbS4tmzm4wTxjLu
LJVLa/rWH+3Qm5e38Q7c5fCq/6ce2xn/MxUM6qdpuhZPbR6dBj7JAjBNcZBuzaOXH+ZtbARvpe/R
IPRk6cFUCUXr8Z9DRJ7NAOsCyt8EwiWl9XyEy+eMjQqswj1T8X/4SKVlhiWi+Zb/LQQu8hW+3IJk
BZq86X9pGPLIqreFGH/9k9Rm9GahGx6FogbcBdN6ZTWXfEIHFY+k51QZKRZZFepoAqBGdpwsA17L
wIXbMLukt4GFWoeYHiGcr30Fdj+blMbPUB7c6YC5pmYVBsqa55H/gpnvSFansmaP6SsOB2SanBao
J9swIAJgCiKnFaP+TS4llsK5teWEa06LHOqN2Bs4hEE4Wn9Ip44ZgxO3IK5bS6mUgFiZEelGKa7I
Yt/t+7vWuxoAIilQLe1QM6I6Ame/YCulUq7AAspbPoPlynWsfRTbCj+jdMXljFDUibLnzUVQmogM
w11371HAjpVhueJqvU/mjREOXo3X992qkbzAieaALBHT8b/udrT+kzU61u2+Wjv9AKOsCiwpSnib
APYSGkh2yhpNz+flgh/t4SBcwSHgGwu3+bWnKziXIGJseNYSiaDq3Z+WaKoxwGTEWdZ5i1eExJ9e
M2uY2qbpD3IhNIyTcnY/yOvrW6soIeLIj5r0yiDpvosSPPvJQja9Tdnd6iyvuU75/aZNz9fh9/Ke
pcAGaeXvZNB5IqMoNhuuwrdHa2e/jA9rEZJA9QhxMI/DPK1MxuMscGRrlz0DGxVYEJM41f1Qwidg
l5mO1Ah+U2ZaB+bQ4yI0JGxsiIWAD5XwFhA7F35Eg8jLwt26nYSbHZd70a7j/Tji+22JwKuXRTBw
BzRMtyfGGOz0dE6S2odMhbyv4Z5BvYb0Q+m+jDMquwF1m217AN4cgvB0SntZupg5BjiTa/ZnIWGj
bhGPBXPTCsEtR6TralO7KPr39VPecSEhK0GZ3irjcS4WhMTMMfaOCtiCo36RnRdDsJwV/08nA4DK
2RaqZgDEqOKWHl8PuI5HRkiONR7Twh+ASlxte5Vq+QjNNboKHhWtdW7rQgz/JBDKiU6RY5MwowbK
ehAAPI/GJNPqgg4L4X7S3yDDdlnQL9fUzltErU6aZiVKvdu0qsUgm6/Jz7oL/nG1GXVcvAIA47gk
QSroWtUy9Pmc0K5LzvcRQS5MBBmMrHHDC24IJqOPX9IQrDvoiSARnQ0LunqGKoGlUJUFJr06zGyk
Xoea+AgFcwWGwap/6129UoXvCCa0JGr/fFdf3TGrEc6zv1yDzo92rVfk/c4rGSxdMPce26ToVc7t
6jSGgewpo5p+nunFdUr9v6AzpP4xFNU4fUYqj+OWGIB2ZmITLVxYPGKfKrBRInEvh/ASmycxk26x
q12MiBPJBTcNlrBWTWcTehBCpe0QGWkryWt5jKs78ap++uD8Dq7kZVhSh0eSC3J3axIApJt1YZwF
0dOy+8TCRcPNHHVdWS2JWqm5VYjiVgB8FdYS84F3lbmf5nbWhPoAb793+izFkDBnWYoiILyThmtz
jYuBcGOllEX+gF4smaGJ/+l5bq6oK/mlmBeRL7mmsfCOgiVE+tGKdPswyOVoVBrQeKv3EYvmb1JV
aAPFxdo461/YY3fVCQogpOR7icTuaq9141oTR+0ogrVUjIVFY+8jk5LNl9aQBkguvMf09QS51PnC
SZKdzOL+0f9tb7YdgV3febxf7rulyGX4MuXbB7/WiXSalrAZ7YmIVO43hyRWgxLtojlv3aMKN8iy
LiiM9hQC0fs9VhmZJ+A1ABAwTMIFu5ybaa2+nRuvQPWboDLYS0iDNnXeFV10U3cXy4Pys9tcDdJi
jGL1ktIf5OmYQjWeLol62g7gR6iB2htRM/i+mvVKGA0MA4NUW4e3j1969mFkbEOY1IfIXtMsXSkm
6AAtgiP4mGO3E4opdC74BRjGoNrRZ1J4Ia90paXJuCD6JuThP50eYibfruUPjbVKphrjgM1PUu/b
pnopaD8FQLpv6vr7ztzPiNGkqVLrOXODRPpCjBC/K3o5bfygjXp4tjskm/c3HuNlvhrx71Ixdtga
SKlCbAOGLlN5OWpmbuzq32LxjvhbmGJHkGMdsIGoHpQCp27wI6ow63dM8Of02fdvKr9nVKMtcPGD
1dpywHgNMWd0IAA1hm8uqXQi5vqyw/te5Sz87l6eCRVHouYR3TnlaWIhfd05mhXVIRXY4wiC/z1i
pSsMlNlrVFXk+lhsHUtmPsXpVmwF+TJ5Q5bhATN/mlqYSfKtQBfgEZIkypkReyFOlEzPpZQsUv5S
GpPWrz8iqlb+Ab7ieqEQ11OxpKvHDwPfqxQ3z+Teei8sxVWzP2Wi+NW75NQ7iafGXjKNOFmJ3FYi
U1offKPHzEWFFoFj44KXd24q1BHcRNR8JQAgJvjE0siTuoXypBsMHC/j4DN3qh2bg3ukgr1gjvcg
r/OP/b6Xuw/E3j7s+L1mpPmGOcJJ/Ap+UsJalh+JQ1x7YLQzdjA6pmXsTr3NMDe9qm6Lz7De46ex
PKu04bAuGKQvA/Kjz5u7aMt9e5wvuooE80Py7BueCaTrKYmbkEoEEtX7UghsghNCRH0g66KaTESn
xycHt8b+/PPjv3lC+8iZLCDiuBfyh8CpVBZ/2742OpBUQj/mHNwzZ2HnoLwqSi2NSpnnBeT8bz8w
fukgxd0BZMQiDMceWd2U480yP53LaNDBrOnLIezdcxQrGbcswvuer+v7RDZQNuVbTRSWBwRsmJu3
u7qbLjbGzfUrqAHmgSMii+QyvIHROCJhT5IwvO3AMxGaWB+9X4oMAFlV+L8XjEGwmrt0UilmHsZe
gmHplhoRcFV6TO8k8Ue8k5O/t2XbI+5DXLhQr3/mDuE8/n79xJNGcvA4WUO4X4w6qTcVm366kXFI
DixD5zkKYQMZxICVYrfXmNLfRw1tDjjx14BL9lpXFQO53af0HmTV/8SxzvRqdbHKXm64/u+z4eFn
oH/fO3oGjXNFCCWWjxg2VXXKciKQVUqg12tbAxPb3OJ49R6ds1QFG+YfJEwsehkQR7ghfbmvVSLo
OpuNcMfzhS0rOQaG9/2OP2BsfGUiWyB4m4hA8vlHDj1zuXapDl7TWCvjMNTEkO3jjIm2TIE8xoxW
vjxKGYvn+Ar8RA8kn0OmTxUQH03b1vTrKRIMvRX1jHBrj3SyAcmw2Az7nUKNyJ+q7yf2CprFl1Qi
KHFonDVIXK9iTJUjZDqtcNF9fN4WocI5hMaEX+KhN0sTciaFjUxNlytOvo9qqAIZVDt09f7qkJae
6hUFY5SmM1KomtEyKdxrF6jFi9Xp/RuUpOvUuqM172MonPq98Q/VyiTQlSyD+ev2CIU17Xji+Eqf
5SFRBAltVHhJ9jk4EvItmUntcz8MG3LrJX2PwoW5Nr4si3pEoeQBXhzYRkL2wLn/3I/DEyhvskB1
JUxZa7XvXe4EvIzWQiC3paMEGGgwgIB3hJ7IcHGJj35szNMCdekAwNysE8QzZMgaBA7Yws9Hd+Xb
dIrBHy3yOtJJf5j7FFaP7lNLQUlYmSiL7iFvTHZvXrj6d27M8GcmUtJaIDOEBhEXx3rDFCfi8chs
ZLF21lDgts+E3UQdCG9iN6kPctT4oMyetgVr8cNrTDrBXPwhzjVdOEawpUfXWC9hWvkDeQRdCKOU
OQJFdbBKQLeuFS4J2bNTPQfjkweEWOsL80jkvwHuKouSNzecqDJ+8SN4IDCF1f1wQcif6UP8lx3e
WcPtw3rWn91GH6dUyaJ5ayPO+eXBt6kWW1kfka4z09+LurgfdGlv1rpWiztU3281ffxgNNsRnVsC
gBYmgLEWYzRp0L2X9gpwiah5GMawbT5CmIX5CuoQCnoUgYsiloJdEPNrZfwNBDWVxml5HX0/awRL
uC4RlghUtVZDq0aHFHPm7frRGRsWF6tWnFBwuZhc8vpm49yDqEAMfKdVpqVTwr87N+hGCv1z4MpQ
mg8qCCOJKRlmkCEvQI2BaL+cMi6FN1yytTFQjM00CwLPRTIqAI/Jtfh4dcaQJWJh+qtQGibUxkdi
x781lDqB+0Z3ngsM0jQGdu0Gy1VYticZVSCDbzbJ5dVhUeHvHCl2Aq7U8EvEMYVNIzeTS0qq+nnc
RO8zwjcG+syExuh6ls16bzNvLeG4qGu13727AMjiv9vQ5c+95VFGk+QIXLiyCgGFuTB5d4mKEVpW
rzUNYbtxn8WBad7DcU17BlYsLdDdWMP5HHGeTBeJ3TVZwz8bScq4krBaKrNCgdzEHFQ5DJK9op+t
FUBoXI1/PNex1E2z9t35UvF6/EPnQRvm65weK3P8oSQesl8WjRbbZRzaYSEOAIfOYzJDrO/N8os4
pIxmpDt32vK3SC6Zd5w9OaOus4IBkC8/Hi7KkASypAEjbROTOGO24STrntRvp2fEixGv1WT/o/be
fkVuVx8CMcXntA9XJZpKqvLu3n4aBy23OUKjTL/A9WpegDr1c3ejdqg2ifGMtIPhSgbhy5frxfVp
QEEXvFpkQFDIdhVjZ4AWdFoooF1BVVL1Zg/rcnfbt0+B45a4bpUhhHRS+eaIiFD+D/jeNfipf6az
vJACXCBK4rmJ+TTK91OCaz/dxgFvPQlVQhuucweUQUB3qbNrLVWu5PzC31RlTSd0v/WatHBzbRO5
z1LKS5bjQIhaLNJjZjdmXVC3hTg16ONlXg2MnN+ul+ntFbavnQGRy/5TZHkgkEYBDkIOhMviYZQn
HVdNuKTX7YdXvdXkgxHE9EK9FGs9LXG5HVu58XTwNa42MfZHdyV2QTUg9ClREWUYh9m9mFUuFRiX
SoYedMm4QTOL6W7hcKXBTLlPgmWgvsgfgxk0FoABTWFXtx2swdIlMPsOuYin6+YMO0aXzdOedtmv
C59Jjip4fo2pPT/FZvEcPqDNcoWfNJRmOyu1zqi1u+dwSJpJiknqLm/wwwLRPcWVCesQ5f69Jgsb
ivw7VnrYOdEDBOPRFEZVaSaVT4UvKeiLuw/ND4KcbSBBP0UQeOrCJvkRp5BlZ4umfqLn36arTeUA
wk4vDPurFQ/eCwoLiFoASAUAy4+z/F5lyXgMaVoVueiYsnhsocE4hpxmSDoHyIJRpAdJJf0QGtqq
WKN58cFifLcZgb1Dh89uPXYin1OIy9Ft3VBHhSTIuzQz2TstSn/VkevuXcTz6pmCyc/7XzUo1P28
CAua9cPkL9XFKGDGXsO0l0QSmZOwZPeC/JuMhYGiz4rb0NvIplAAni6iftM1vu1ZBgrBv7b1F9gR
hJn73dZX01Tw6qK9mE57VPyA1TlV/MHNmWGs3aRRmYvRkPNLKYX2cCwD96VGM59IgRk3wNNpE4dG
MtkcjHmb8j8utFN9HKkg8m+CW98wzbDapSxnXCUt2NsnaQSOIA3R6mSMxQTc38mfwwGrTkX0S69f
9Y5lmJBhEYeu0lWezv6AAUtjNhAbrcSCbQO3l9V1DN95Z5wp/h0QV/xAZ0rkh3rKBTUZqiR8knID
bJ8H4ypy1MlinXyS2XOsXptkXiSCAOdRxC1K61PT+Uqhw1PD57iijT2GdMBhgbXa7eVDJPVosUs5
KzPot5rBmrkDiQ9xv4LZ+Pgpr4yJX9uMHQqdLwQNosHZ8XHGC4/rckyUCMvRgUfcNnmG46wwXD9n
vf5icO0kg3fkbZVrTG50TjB/OFDFuHahlnrchPeyVjXG0bABCxTrlN57sQYC2xJB7XUaNq/hn5oE
O6mq715l9g3X2urQIZiIzaTM93yZFMR7BBSAIPlkKWKl/B3FzKYZ5PaJod4Nc84i/qmP01P5G7zO
ApJDeExZUfZLhLKEJ7odGzfhB/hvPjyPnqYdkH19Q5ssGWnuEd2iuCHJLWkbodMrRo8I+KFsFwa+
6nGxbtJYvJz/5ZMTSe9WEXhwqg6GDPkDHnIwVG8u89mh9PnRHGHCBrQA8jYb36Rn3gEjBirA5LA7
4kzqqbdE9iPbGppPxf8bjUSoS09+ghMgS75JIkApr63v41WjdRMr+y2f3E7q/0sDItwniWDY0PVt
IHVtBKQLHafB4sEnUUJzRTZqmiV1eSWaIzPMvm8IH7c6IVwlfvk2nWhf1rR7GseCHXS+bLnxIo/S
fdD2qEy+bUf2CmedxOjuR5iRIYhzYl4JhJ3zEDoDoaK0mUsf7j9GorYSL5j4K9fLQbVAF727aEYd
6ClRk5IFmACBWoQBkz26h4vNbEB0m+/HcSRpEot3bWQSkgMXYa0YUXSRytdsgyvlp1BmBU5o1nGy
rW0+LkAG3fjXpzkcXbB6WzHykL54x7WptbY9tfAO9sTkpTIEbLbARQ1MhuhGKw08wR7TppFVt4zm
eAdiOn1Nxxr7WhD+MBhsmgUnR49HIBSV5Ap2qcoktNNGHeLepTzhaYA/1SSUt5Hd5DmuTUROyfJk
H1C02cxJEEIwam+SJaT+DOtSi/iNE0z5d4oR8FqTuwfcjs57lLK2XyAGmoL4L3sde5QHTu6T1Xgi
goTxP9YIJpSgDWLACLp0cUAAF9/RJgB92QtR40hH88MqStzMB14yId0OgtIvqrfhmIPVw8FewCY3
wLhCrGYQLOuJxLT+Gv7hPxOBZT9ggG3FvfFTH3PD5GzTx6G5CQySc/0+q6y47TFbApMPRROOEN7r
fXQBmjkErMBUMYOK0KfOVW94aTZF2gsUhdQEt44fHMbWmsR5u3/i9BjOLlQ5kBR+19S6lEVORPvW
yXtRriJT+DiltGPvgzhjnxUnMES2edhjovD6ggdSMpVHfG66FtvgdWS8WSOJrBjNQkiU2hb2las2
F6AJBDTA490MO5F+K6BMcM3QJAWK3H6uBsweyFg0x6rrJL6teUg9eNGAvztZumdlonry1e08hQST
3PXernbXsyoA/flWGwMWtDtym5EVbZUkpxoJmuZY+0ZqgRRmeTyjyOd7v4QtzSTQ/RT/abPBo94F
/WWtQUAcr71KaUc8rBBDWJhU4Z6WY6RsWKF0RHLbBBDQs9e+X2XZNEWcxAswSxx9JDQ1dNUGESD0
3mepXvS+dXoWAMIojpfKoyvJ5mgl2xE+6vrhZ57Yqv7jZJYtVMzvuhqozf4TMlxLyKj0cIE6L/Si
5CDUbA/h+HDLwsaMTMDtpokSX2zTeGoH/BhVOrYuEX7OM9iSqB2zD/jAqYwtXCWGS2jR5jaF6jVS
2VYrSn/QjOV8GrubdYa4/1ToaHFHv4wv1/jZWPxwuF4L5SSR4qPI4LY0ks9kykGR60P4GMpT8Iyd
h8GX+kfMAixeXco3CUdIhyTPF0QIg4CdQCpgxwrHkVrFeKSIqYBrMjPuJbnboGorkZ0O1tZT109I
Z805bBQw11/5hQpte0T2pRjfpl5i4m5RVC0PEs8hfDq1RvU/N9sNhqVNuHb3LUuLpV88wyHBY2+4
JLPra7EHk/FfG5N72Sl6UAzb1wLen6mQ4gLrgtRb3EobK8tSE9XwcOO4n7fFOO/hPItAapyWvrlv
fruVVbxwg34E3IhvMCE3JDHSbVPc3yKWybS797vbwhUux47YvW0UipkUVC4RnzDi360NV7a2noQ+
klcPUcNVwAukznXaaDgwxZ+sJLrlwR4t0wPSipVF9pv2oEuG0FwUk3NAms1dg0JbD2xQfEmOzyrf
8u8CxdI6r6VxlC9hE0QH+ZmsYZc+yRhNM6knFFIz9GfMPMdLIE4MCAnF4JWBHzSq5f1cLlatAe03
/4+SPGlxQ0Jkqxz2cILNimG0gdhBoopoOWcq2rqPzjDspMejCl/V6HFvLCD1FWNAvi1idN4gIjhy
m4xC8787ZUimvtVCguCaENj2wcLCRl9vJrJG7kXYGFpY8tnG2SfpR2xkbOUA1vlv/cDC5W7Pli9r
3JwR7qeJat1EudIsTzfkZwVS8EhwyzLBBrbCZQvbSXN74rGTy/MwmSFR85zVVuzLqsryyvlGX0Jl
nulWxc4TOJ15B1r8iaxiXnxNMAdchgkjlFiUhBwKWqo9GImJNZyr3OVhBBrNONotnOtVyX4VNtdo
IW2A7z48cv9xMbStZMgLyZKrCLnHU861JO3Q/q1WjQAZJZ9qpnGV0IFM47Ri/n49oq1gse8FkHsi
zi9UgSC5rcIeRpNun1Bfh0GYXa9x9X/fg1T4UMrKTdD/4Mu3Tl9aCSxBvch+ZdxIXWgavwEem7z2
MhUJ5pRqRjACRfCS7MVXYtHpOvmMBsJNgvdaEoWRjtGoTptVUeLjl2DAgXeQ2Z3XBKNIDN7FYsJ/
8Mz6L0JmlBMcZ48FuG1PVP/guhhOhyOipQ/oLub/Axr2TWtGj/ymwKCyXIdxoxMokYqJX9P5uN6Y
7BOH0ngqOtokL+pHxwe7JIdeIovbVLVrwLl8tpwffbpMciD/xkZQ3UylVZDF/D4JK/JyZ+bmFOh9
6d/eFmucIJFsm50KvnpLQH3R38fn3mtCGA8dTn2EdbJohpKbt8njWpz9MwS7Yniz5O0pajjD2wCk
ppmWIJv2KjqHh4XBvdP2o0bDHLNfZZwt2O7KbQW+aO78ujD+Loj8Nz94MfPHZhXmt9IMj5O9HGjy
C8Ox9fwLUWhnmbzLyM+vy+90mhVUNAQPrD9uf5/rJeMoEatrj/+9455/MUuksO2JGaCsK3TZZ/tL
3jMvXdYzwQrNx/D2iKHYJdmUOzpEWvEUMVbAJxfJ7LI9EihaMBYQ2OQVkWM5flgckrc7PxFjAkKM
u3mBUur8TpGEjSLPpcKlTN1RWhwdq8KdvuXRw2tbzsgClyKyUxEhmeCaWgVqQP35QwGs/fzoHtLU
uDucwO7GY9VrulDDsIK7HLsXV8ucH2PaGdAyO1a9NukwrwygJ4KzNFjDrVscNOLZLfxPbhIEgdSZ
cYUpCaVKROQxj2vOYTxiLeT5pqcZyc2brh6JHB1nKp2pFi0xn2Fs+mvU2XDKbxoyFUScwswYhSW+
IE/HsGcB/GlXdkXMVSBw8s7fS1UFTDL3mZfviuKA6Txa//DWOE5Y7D2T2Zh0/cQGdVAvRKst2+Tr
1qCIuWyKS7WR6NXotgUDBBqeO9QNKL7pKcT8RmUHTi7NnrrDeVzUMEu27ax2Fp9mtmBHDtUZ1a5v
Ry6jdwSxNMHVFZOIRTFri7RWy5hek0nitfgzx6UATq+aGcY6ROx6dMbUtwFWNBxnSWjTD3GSEKNt
iRGr6H6BmYCX6T0HswYdWbzwpDSVFRtEfx4FaZd1mF2cnvw/o2MGtN84TOVnFTaXUxks3hd950eX
L3sod+Gl4hanDhvTNHwiP7Wj6IPU042Y3PwnTP98KzmRmbU300+kApuda1a+gjRNUKSwI2OwhhQg
qN+NYcE+GQN1WitqGR7VTF8nAYGwKjMpPNKxAzKw4pFKfgOLaZwJ9q+qMnEG7nEtekNP1nfqxaKM
+NiItgEYVvdPyG7F8xCe2MvfRwuIMyrPPACUNLdYJ8e4EAZy8EAbqYsnvfmfJZkiNiVCgSZr+nOf
DgKE4+qdrBbsMVHwoIMh8E0D3yEwmV4wjsD3XEGiGvBcLFF+h88hXCAkn9BwS7ohOo0XyhLa/X/w
dg+m00BbMDwpl+3K6UHCNk0RyypkIlHbMaB/Sv7YZXbYKXwT9J5MkTPug2lBAFOJA+uTerYgTfQ8
y8NFzVHLWExYu2elSmBpTdZkYseSfxOyd2+H3BzpXVyK1i6LS9KzJ/ImSiHVQxALFz8BBCy7tAsm
OnY9IY0TW/3v43380jyXonpZ5Y08aH80XIlcgFoaW7lkuxY8vvGGuKvhrXJ7s9B9zFlBW/5r5v+Q
MHLjD9EL8D19lqqKQHUQ+dGOOhUK7gdwYYxBRV2dqGiMPJ84PxwiLSq7HElG0Uzn/5IQ+b6PT72H
yiOJsqGvm3lnExFo9+ur/Q8WC6IZ2v0TJXdNWaiGVBZQp7o0bnK6lLFUPptFUVhlvoTbfCMpcX9C
8ZWQaWyxrc8wUwYKcRLg2HJRyWh3x9HI4l7WMD7JaUUVcWNp4XZ+Ev7eL1lJBpYXFCfJpimkfmhu
FUfOwL4hasSEepPIyYZJv79Ty7sLxXygqm5SxSKNtqMDZAptIRBlwRvX0HqK7wj+6PFrSjJFTHN8
IKeT4yHjQ6g8x9q8qmbtjMuSpusf7VOOapCFdndcS95l6R0Q0/eYaPh2ZVq1qxMKlWPXrGUKrsId
ICjm81pSIqPMIcn2eo7xXihuZm4Q7Ee39uTZKq1nWzl1uuS59euJFUywR/KEWlthiAn1Hpvfw2G5
3k1JBqZYMS/Fw0uHMykD1eN+e1y9ByfhavWk6Xd1AXMSyZrd8Nzp8LxlsJU+dG29eRkHGsmFykXv
hWwTJHpKmXhzZ8yDwu2Q2F2SQhu0rvoHPNofhTb09a1iGDlOSyqzegVVz0fmMLmwabd3JqOgtqu1
FJ1rToEP1VR5h01xgPOOIQycFWKaLiweNnYkVAWmche+dEPQGc+WRNsAUq02yPCGd0PdkXb7J2Wy
kzsvLq+k1nlv0zI3DMEyvZgw5u/r4ND5kEipClXajqFOL3ywXKda0bf1GXIKRN3zBq39t18UosP5
z8jal4cVnxiIjUspp4u9UgkBk1Apzlx/MLPQzWgAoUSiS5CXzJR2/k+GyHU7RwshhQ2evYKZmz2/
WISdg50csEV0Kj5MULIP/QpJ+lEj8ylaRD7dXQ9LTL6yiZQ6FPTRVsYQIOGN+QSn+twimHPvTfOJ
n9CcHpOBguc020w7ZzWzhxqLfMfhmIAqrc9tPS0lITEEstJ+lEzDBGzHtV9UKQdYCgydaok9aHsG
KDCE/9Mab4Lir8UdPzVMhpbHBNUntMScM06Fhzy00eLh+HNFzumk5/JFlUhU0ntmkJYsJrkcTdue
g7QSoA1cbNp4GS7ejdLm/lh85SbdzPdEyIZqM3wnEFXJSSP/QrP7uVAAbge9guWQ/06p258csJQa
b32isg33b5IE2Yq8tQi/jV89VHQFG+Wbr8j3tLZzRiCnOyKhyHNyKYDxT6YS6okPjgZSsiBi7REg
Mc3YZL2MRUMy+Ju3zGbiit5Uw9r2C8cWcsEgBVKf8bdQymKQ5Q4aERWY5nJzfwguxPT8xtfVtgCw
XBwYp0r4iGjr1F+m4GksuhTgejd7SBP/6cTazcZtZ3DQ8U9O584LdkZKrlEl1XwQ0flDzJ7Q54KD
AL68+UZT8kPrJSUDRIkqXheVxbvv4Z8skHm4k6Ts6JTwlLqYCqAzIkclZ4OC5x8ndMaTh0svMrZ1
ZLWOkcRfqknlsWWvnp/k3Pk0rGpdoJNdgqnDQC5/Y3T+GnAaRbLl0wfKH8snqoeLIy0KfMCJbHyg
4BtxS0m4bTN0/aj637OoySYnldX1XcZQGSdAM1f/CtPQoDCGXTG3hjlAM5SdFJ/Tw1aYOj1hSSAn
wh4ys7bs8LDWAmn98QIYuu69fnO1xlpJD/dNvhdnwJ3Yq/YQJ0DTJRnAslebfIIgkx76gUgAFluG
bsfmdLBDc1B14AENUM7kWTli7p5rxwjJ6mPVDSgWbrpT2pGjanuvv1fTq/1qsSI3UHjCu8O1ubeG
A7X6NfU/So+Gis/mqh6gV0iSOe4F84ZyP3NyO7KjJEYI4ozXC0k9+nPONceYw2hdlzefMJcxUSen
GO8xBZ2qAniWJywBR3rPLx3f24Iqd46svfvRD8qU03O/7Z2mXPvFA30IK7lVnoyT4VBJRdg7/LV5
mtR04rn2/xHXzbjvrNjIejoQJeN7HRRn9Z6x2oMdOjglpDsqF1HSBbss1iyP8ZtXACZuGF2DAQfI
EAss2E6T61NalAL9Ja3y03PHfaLF+4EQwhTB63di+lTxwa3cuwL4i3Hl/vruUmg9S11JS2u1rpxJ
dGzufEbAJkMFTpfIAl98KWFjCXFuJ20U72J0hc/CQLYHGYXnnA5zxDwgcu+IZrGSNeekWkVcJrm1
djB3YltClC/N4iovVFG3KrEMmyfJKn6NOjehKLif1gBXpnyy3DIOzxIxvnjIQODZbAhJmeHNiTwf
q5Ubi6BgJcIjY2QgZigTMUv9XRJjgSmErR2vZbyT714zT/hbkm9iQdxilOdcGyTXqA1te2UBf+bC
Udytfpb1SxfsXk5lovmDdoeW1Oo5QDBdm8Zm5HIOds996iF55bVDY5SIj3cR7PTQb63Sa82YH93v
1IiGZ+vgCEn/2VIphE6vGG9is/hFIGIs39jCQZa7hUU4YYQmDfpVpttf2nsODgsO/YXhutfwl/kE
P5z58VvndU49mABSl88z4CFcNTJiRhZICEiDngxaQsnJc8WnQy9DcIA32ISZXhtMqB7gRLw+VJQm
qHrh51glxhIS5+pfISOtYJbqVm5pA47Jic+AbDl5IzmDAULXJ1f+1bQ1qAs8UyRKHQincer+424u
lWt7jk+fHNES6+dq/9NNeLAOQat8vqy90mQwwO59foLw75fwUlaw2OHCEmFKXJnr7HUrT6KPWD+k
Z9YwtJ+2eTIxMzv2fzwHLiR47wCginic3QmayTxg1ldNvkWq21tj50IbYd0SkQNxUpNx2iIhphJA
kd/IaGiI33nPI3K3qxnjFYWhDvNiglL2NYk/6KF6fMDshBGihZtolBl/O4PqdseKtO/be9rZkcZC
hT52Ct/fadbIayhacUbIOJOmcgaRZ6bC1VGsy8WOW27JGo7efFQrj7PTDIrIOcvlyvp2TYCHz4We
MyaMiWiS6w3NyetoRwHZ6g3g+Aqcejk85F0ArfJtSmJCJWsf//oNz+jtAFXZcAAgLvT09La0zD9g
l+bYIrQjzcD9up89fAQAnk0cXJmLncOKqgaVDr5l7+2xUUrdz63SmZ43HlrN1sa1i+wVxmMnc8iW
RjxGltYhvZakRUrhaIGi8xepHczRpG93sDRdkmaJhVm42OjR3xRR6d32vOTUxCqv0xCxgKLbJ3VG
vWEoYMuKzP4RvBvSG95yndXtyDEdXGMZo7Xo2OnsHq4fHqP2I+sSZBEzU5CCbpUxuY/17/5EHueD
tlIoCyywE2eMXBAiYmDtgJdRyYFyjwj9dXE//HIytC0MG5Hrb3wzphCqLsS50X/WqC/fxdJuK4nZ
vUyTgwRoIkUrFWyBE5xPQmb6qqTlmlU3tjr34gjZgGDeDM9L5ZozFY5LYopTU2B9LTw8sQoDCmqN
RjccVQ/pbXwtI724HYsGT6K4j1VAGGM9CVmYoqNZsRv20oULg3eUmj2wbm6Vy74d3o5yhck/j8ht
BVtlx6LRzBt371Z7l+3g3tCocyfrxJnEgHG3D9N02XoE5jsGcdhcNdjWOAcAASkbQ4PGhUK2Sr/E
ZecP+EkBHjUMiC8RXOqAKofN60S+hXIlageQXCkPmyhXNdxHuX3Ys3POicKruhXRUVioq7Yfk5/f
v3eJxJVzixVcAPC3zzFKE/nlSvrthxf/ykj7chK2PSEqHxDmFYDWa5DhKQA7meZiFXg6s1JT0MBG
Q1PE8W4wLakGStoVz0Yi4uxrMGnfgb+ITPDyL3AMl5zFojqEbvDyejRlAFdQfO4V4XUkqY+ohBTV
p1dm2ywyNMuIuk3RmI9Nic8H5+z6l2JQOAre191Ij0ahH+Q9VsC4BKrbUP8AjgXoUw2kMQ5Zd+Tx
8dTD1RAPm9C6h/74LYXiZ7NtELxnx+g2LlwtXycFPncNbvzSaksaRynrnwtJKXatf/mYpd4urLIR
vGUgdlzMpKKuKJn0CSlewS4av/6u1PWSzVQfOZBc8w373/NkNP4Mnx4KSAqSZgBXK3ik+u16wC0T
XU2ivcpd1oD9BS93Ls8VFjD8XtOb2kOVryFDK1qXWhQrdKhIg46EXqRCB92WtzLFtJou/9swaNOd
ctpCuVna9dCHpYSc35ol2ABIsGDY23KdQBy2yHERccFuw3hVmort2HcCmGSBt2WAt+X4dCRWWy++
h8H1mVdgaEpMNrLDVrcPxVeiTYHg+g1FuoSMrOLaxsIdJj6iVBc4nRRGG4IlzKpzj6XinryL2+Bw
twA+BB1OUquxtPDYFUC+THF6PO2mwHnkXq1tzlTUT79V8rzzYR4YLW1ljvwIVlZJPDDaHnL2JTgI
BnEMMOZ5TDQ4kMOTsoW/2k2+xCtfROw2KTEyWHcqqPdi+OKlESPFKMDE3jzauCWeOIUdD2G/9Fj2
qXhSP7zG5m5TMG4KHUySXXJVUO7Kdc2tnCDVRTbbO0Gm8OhVuXz+51ypuxLe4aZzLn+6hSJAGgt7
CCoj6OyawC7Z7FfLjh4U2cP7ceqohfhSDNK0522jbNdSSE6D6M4yOb7gz0Z76C9vUeO+BQOtmD6X
QDTtQfnpjONQVMfqBsrQfMN1fdpsoy8PJ8qNd6G4PVSnZw64VuwlvVC4mEKfERiYMXhda/sWG+LS
YBGgg6WDVQqfNfOOyej3jrHEsEcXKi6ZCCt2lSDW/pVnrKunEvppAWYnl1SPrPppb2HBKxAdd7Tq
faptx92JESrwg/dILRMwTwx6snMgZEhhf2TmVvXU/BeGFh8oIPjQyy2HoPgluhoeBOGeuKnkc4Ck
5NglO378Y/9F15McEM4T5G/fv90+vUSIrv42G1B61Ri1bWOSe/kWKkVpk9+BCbLqizH5xxuUz1ry
ingFPD0JLAE7laRmoUGwnB4vdjVLqa5orepAGx/GQpPfgLmHwWcGhmzzL8cXQyjVkWcwSO0xtb9R
T4DTc1kKD/OyXNQ1WeefbevFbhaPftLQ44GX558gI+Hx6uTsHGiHEzxlIslnVd6nSNzJzHhf/0xk
qxLjO7zzb8koadi/eCFaOgmPYlFxCs8ykX0z1QZO3dzSN/E7J5zv9b1GHnM9B//KfMHwhMNx61uY
TknYYNp2mj7YZ1FdBPowDVBhnvUXFFDw9uAFHpG6oDOtQqEcQ3ms4e1KcXxlEiFZU4p84+OWe0QC
PbTpA4C41iQsQK8aA1qnfdxaCR3wk+DAi9iz8PT+uaKJ05+GECJdf3IOVxQcI8QqNb535qWlk9qr
Z/C7zCq37VemYR2UTRHwUekDle80YHletqXPKWOMotoTKZs7bWc3LPciQcNOCXgIuhhn5/wJ66K5
bYEMZ1l0YHx30lZ7aJKKxggKf1zhtUVq6IH6qOa7RrijLRkvl0r5Zo7IsBtBdGPM+o6rGBpCwha7
EigiZHU7aXaXjRinyls7mBQCWWvqc6XpkYFJrLHT3WUeEd1GT9rT5dvLRl+fQeUFVL7tLdZHepw0
wWb7EuHUoJUDdOl0XcpH+KeZufxjTEQvTdQV6mrYcmlwmH0nuuWo4fEW4LGJtZ8aZcLItV9WoUIY
5ktrUFpfJmS+/zjjIVGQat0HMFCzH/9+81xpj+I6EbFYKKvu06AAqvDmy0AXV4StiYOn1eq4tmVu
/BfADtMo3R0QLRCR4zGgdKhnnzppN0bEYtGr9WbhMyst9wIKblfXH+osWRB3zV9zZrQQOKp1L9d1
uTgbHW1FQu97/WB7IBeqJ8KnNvWJYW4L6ZdTZLTkac60gV2wkGaI5Yi6DkEisizhGHRY2EpNz6T/
rhNT6ylljJH/c+/dWruL9CD4RmIKbnCFGfQbK2u0bZOZ2TDsfLtRJRshyw9geFS1H/vtyDn3XViG
iVryioHL5hy8XumAOdE1euYz43XFnfgHIDHe1oWvBdTnBZriks8l6IpwMaQ5RD5ine3a7c5Ip3YC
tLjhtt9cHPYCPRdCXdvWiZ6oG4cUQp0qktGKFhbKvoJOZ8lKXkmeKmTKeDnBJaoxw33O/qtP7z6q
hwAh8oJIbkoyl7fOX0685ASQDWSj3Mte2qS8iP+0SpgQMGglVm4GP5r+6LUClu92T+YdjrxUv/Ae
YG6rnwsTVRPwS8QSHc+fTnCgV9IH9bDZEZH9sSk/EhQkmCiZaUFQ04SAHIRhTcGKLxVjmQ9sQw/2
Mhqemvz+bNyHsavBnjr2uaI4vq0UjFGRn1tbWWVHVSYCmzpzOheKFd9E0/YOibqHefNGQv3Swvnj
MN7Ht8PwcHUQL/oXmoZ05Z81L+wOS8KMhEHBBztwtb1vdslv8PuZUw8ICWvVdRihNIHq/luyra7i
lo9mJtLxiIE7SxJE32pYVRmHGBWlfw7l0rnh1ywMaW2k2y3VA9WvHSDH077WL3/dDllHXVznrzlU
oeur6YWJAKVVvLAvRwetECLP9YwjPl30fkse4lBH/W933wxPEMVbyeg1kbrTp5oefaoxdiQZ4o0c
Yj5YdOq3tNi3B6VBdbmjMfl3qxil8T7lh1y6PTNK1SqVCbl3/eA0w/jlynDZO14pP+Y0uDSf+RGg
8+giFa6IxdiivbNhvSMTAD1/DuETyZs8k3E3xIVObVWeoXwRX9HVZAH+WTVghJCtoZb0uhKSO0gL
PA9CUwpbagh7QxiRRbNapeLqypM+3Zavo/NEdgj/NY8XChJMTjB0GK9G0hsx5pXw/r+wY+PbtWCc
5PLHQgwBKsS3qwgVxQq3mZULfmlOr1AHH5KVTy/mM16ThA8v78JXwlz5CBEXN/ESfHsN5f0ZlK/C
CtulCTMM9UBKVlpOEdQPp1PMmuigjwYfxSPyTa0SpZ9qHygbnYcsg+YSB2jvXyw9v5EWln9TEiIs
tZw2zuaGax7FR1mNteEMucC0GWNAWJ3fVsjcs8B6CIee1O82VT770RGrXhTkZwJrcrUPKJCnkzij
1klg1XyfK+xH2VBJBnoEKDY/6D3i42VybdztAhw25HTEXIosJUcPll4IbTvwQXkJwZmQjp8e4a00
oTtbclfF1ETsylGz/rFWdETmI07tPHL12RpwP8QSuBhMNBXqu0301AvOgj9H6BXf0s0P1LuRuwvS
LrWhpZPL3V8FAuuEdSIn/I5z8wGDdLgc3yDdeXGsRInXqAdphiAXwVqi+/iZZbYrC6iZiOcdkS70
KdUs/r8jQQGqvN3F/FKVcECIfmmcTpsXeTuUgCzcEi3c4LBEyPrZA+wp46TmiBnONth18MgJYS3H
sp05wELc4wpcLjlZtu4gfiv8AV3kX2E9w91Rh/lT0lJWX7YXkd+R8qVRRbCrN3QkhQFqrviXvIZW
ZoYSAATyL8+r91v6K6GvnnV5UGzEmLDO1AlvcTyVThOvNMw09NKBJCjPpuPhxGIYwPM2fj/Bnl6x
Liylpac76JZZfl22l2IVt24e+621nTb4/8tXPPv+qITh0tm8ujuQ720aKKBxis8iKjyJUVS+vZvp
K7ozpKNOYzh976wRX7gLUPOgBrgzFJdKChOlPfbwufJoAQzIk42YoQRxtSjnmFChFiwSch3vFJhr
DLttFpPKs/VZlnMiIgajyMArVlaK46BJ8Zc3CShN336nyGIigmYKPUVFQ0ppfVwDCx3NocY0Yevk
fJFWt0VM10kSmiHrNVaK1GsN1Np1s165rgseH2H82A9PH0EmNB/HrADBseGTJu9JUYqAbuoWa6dX
p7fbGiPa1fnzr04Q0FcshyV/601waBYRK0VlSa7OMK7BSP02vHO/ppcaSPiI5SuQ4zLFO2iK6ED3
UisSWgotvFer5NRtKRDnJMtDI4auTIO/ItZC1m4RXJWiSN9LZmIM3VMbZC0RY9/gEMQTv521Ay61
d73PyayVTelJOhFut1mFLJ4NuhXOHbKKvDqUTXJBeAG9VDqxxMHEihMSdnSdZ9Ecv/1rzy1VWVZu
4jlcQYLZwEC8MHr6BUPF84cVWO7RFFxJ7jTZEssIL56yVfod0QWYbQysoraEHSQ4mRcu4rEaF0FG
4Gspu1boFyrGHplQaxt/Vf1E2V0igYOlTxubYUwmmzwzrFVvTgoxNiZplonhUFHhlUBm72r8Q/XB
wXOgiJxpwvT8ZJxAK6+DTigBH0tg4Ap3TYQa8PQQxwMmIJ3PZK+ThjXREr9X2NzzvisclA8kkhp8
fXZH6t5+HDNV1ywPTqbwpiB+hQUlUPlP06qF0fn83Nd+C6fnnQQ/RFJJwAxdRtx6rXqOQcId6O4Z
197sVOv3AKvamH2qh8I+mqsvNuX7mNWRQVOwifl5P5hQihma84scWSWIqx3vkUDJxfu8hSJPgomS
b6T6BXL0Hv/pzSUrsBlMoiDkhUjllebo3A2o+U/VQV/0s6IJuKpY2KzS/csMQbHMreHIoaGIP+9E
0Ye2TFyko/jDqbrxmjamacKw7wm3cWjx53qpd0OKgUryXSCbwcEW8OWhmP3uHTwU0ziCse2dIQ8O
4kssj0EWWdCc9zIOT/rpmpmgfC2l8UT1p4kOxmElsq5OpOXAEj8GVYq7RDILqkKvryia/529AHVd
HeG+g8kWPOMnCg5eeTnxKYqPu1H2S8uDPI3I6TwvhnHVMaNfija358rfHjSNRc9ZgLoWhn5aoph9
H2elFcY8O7wYyS61d3V09IraPpjnNnbaQjolPFgK39jonsg4KHt+NBKTQ7wlrdnrPNZLbi+RnKth
QV0KBcQF3jTJHuRRjUm6QhpOOhaz9C45Y72TQzCMsB44ymFNLrB5Q/W5jJ73ldLgdA4pQcWRz0Fx
w+0MxfE2SnHg4PEVJmznJdQsKVQ5tYj1eNW30S9STEKsv4om3BYajI8T/pYxqOT3FI8I0de5LGW6
H6O0237tG1UZOhNKoS/afxmg+vg5z4o07ZXbb/Og0dyijru7LfyrodQM8yV//6q6T0gT403LunHY
mkgHbDRpBTQLtBJsRRQHF4FMs7f4jWztmOfydXvOTkO7Wi8Mej5XDb1gsF53quc1FuBwN/JGD4hO
8XQyWvNtxl0RLZv/t/N52sitb9vK9HA/Rf57dhpprPHYX06nFgxpdutUokegn6UDTHl6aD3Cb64z
Ex7UgBwFWETkI6c7tBP2akT9CSl/p/6KtcpPJYz7hmmS8AYH6D4cnE9TlCDtOSPMMiYkUpjeLnwi
XDuFJB9l+ofJhwvPDA28m8pgjBp6O1Mc32c00Ckm0bDg6wvy2MXgcGDsI41LMpMBUFydZAqru6gT
jQBGFTmrh7dd8Yy8W+Djz7xOqNdmIes2lo23EzdiXjSjWxbHWutkBcyBYyybVWGNOmltN4zTNz/9
wlIWwV8H2YHun6pPX7JzxRDwEgofTkqjA8/dEBt+sqNu6Vzadi74xoxY22BV8+ke6TfbS2rLqdFN
3qiSsarV50dqB+bfOT2C4ygMguhnojyGr9jkO+W0bBEHWsiWr1kCXq/Ca+zpg+J/R1yzLDJeHaRN
peWPWrXzbQdTf/soD5uA3MOkf0DplbnG/o1BNhkwsPR09So77JGkeNu4jv+cY+ioCM59XwjuzGSa
FC/z0R/CR/dWwbcCp5UXsjabmPjaDfPHKnfj5BX9bIX7cFRjdX9J/5ERtyUESYXhHWL4JFGGO/o1
bghYeiFVJK3VoaUfbvilLdaBuGESro35QUMb9jvgvS0PtM96rkOrhYBf4YRa1XMHnu1IGMJmHfGU
VcICAZ7nMVJtiyEEj/1SHetUrP+2gb+wI1XWEHKDrK/SImLPhQIP0i3WKbYekmqb0PIRAhmEfm5/
G3dzZG7hs9cyftOqq+/OnYYiptkO2uHITb5BY9i6uTNiZeyuIPVfXd7CUj021CnRDRCB/gaNk71T
QgfcrvYxNzrFQO46xV2j9l3Gg571Ks13vouxcgOc0xFa7HElpr5T2DElb/hRX8h4HZEeDpC7mrok
ezI2s6KhgP3kajNdiqXPV9Rtg5WXuLKMvtMLLwpkZjJUQtiFv0rCN36o9/nf4qWjLitLUG2AVz8m
s8UkMMf6ukA7S6EPeQKMOOuyHDewAHl+gTUIPk3NgmFs7lyOmZ8KO7nRBVp2goGnOW3ksnQUu6by
ECQBrdZ6L2tnu4JELfjIfusVhWi8m1VpiecfQUWdpDcgsGCfUFsva87kKRsBdZFaqRxOWhXO+571
/EGE2D8YLnsepxsWjsoXi3VrbdmenkwvygakxtixZt23Ku2Mq1qyA1wTn08ZmRBh+LyW/wC9SoWD
lffv+VxN0nLqJPTgrRy/IZHnlbVmFcT+4q0xXLOBzPc7+zVXEaHVG56L/3FnM4ge3SHtinXDzcXW
cHWOtShK6Yh15VpcqIXlfqJPtLpQbTtYvNyL9O1r6tcdTWjj4ioFVgfiioCGZC1HrPs3uz+SWrSq
q4ZxAg+FEBjXtc5BNSYtdzWkaoUBtrw0yecv0zdLwlRT4gFirUtxjodWE3pxmt6/wL4VHiFeCqre
j5oY/r/Sj3EWov8AmQEoxAkimFZ5Npgx/Kf3VVJe/O/8SmFYdAg+BNQDRo7PCr33VKMnq2nIoeFN
zmc0tYWTJ15pP4lpIPL2gYvlt0PWEPD8m5hbJEvkVQUkahz1eff0PdZjGodsQuLW9yItPJkYX1+X
upsEJKVNyM0hKxZEnk7lr0rHiks2KhBOKgMcTVaLBIRA6IZRrFMwKdbpq8XR8ebhkUGeag+RIqJ8
SW2675cwlU6ai9Yo3xHGF0wCr134RCDxgpcBdUyhcfXPC91pBU+RnP/2ejJSRhVrelBw6XjamKwm
HVNf6g1rT6PJtMEKy5Bp8B4Msg39508ROr2AP6dGoa71ErVa+70PLH+9mn+5EHXNI2/0+adjIlOO
PQzSz5DNgbOx+kpiyEyB4WUCL2g2yPky6TKfCH/p4UQ+9VJ+aOttlPXuVfLYXxoKqYRaX9fNDTll
ryar3YdV5pi6wqD6Cafl3JT7io05avBdeuwtvfIFLo2HTt/1hRjlymoaRNaln5HemeA96vE5ys06
Of2rfvog9lMmLjy+K48I8KViSkFA53WfviZIMy9jbl4OPvIwWH6+xQ8VdaJBqtqV0T2piosjRGYm
ovf5BBp6ICSc0FlHX7QB+VsSYs6RgJXrFg5vqNyrVj2modLDqGVK+CFOhU1yWsRbPlEnyyLqBNni
FLOcjjfgfmVMHmwzfzufuZh0ZNcIMH0Ls6oKZX5JgkSRVzQ1wrPNVUSLmrQPkZyIC8Z18BdUYxQz
DGOGG39168bb7wB/xh0sR4kh37R4bRT14WVnyESCWUsTq93xA2b5RBKrLdePrgnNrj8GnqqJXShN
gR64pFvsuO51nE+nOW8zLrw3GjZ5j1PaTmWg4yOHWOTioTRtzVd8A9V/lKEJlj4/+qRGOlftacdU
JKlyopOMTJy9MqjJwAh742O6nCqXmiicmXL/0+mCFOm9QSqwzNH8U/T8ULEReqhgT+lZDotZ3/w5
aUDmPOak42Z4cAhh1yEyrrMIpdwhS6V2J3UZofS0XC71Yn4GtlqYBAyfzax85AgB41ovvR3F20G5
5Bqyhqkr2FMX2w5/jTIMcjg9JgoL7yOeHb2PGtNoSSR/LSqpkci5W5DwVunGfoX1hFPYQ9DG8IJ0
FdU5iqBEn5hmdMUue/U7WEvxJqJVzR0BfJsnNciGj9qsNKqFpCxgCNwZ+kwhbpKPsx8bdfR3dK4G
uOuYplODhF+m3cHCcv96LcOc2uYPmMyN5CKJtue57Qi4UJqjF2xmVJ49G4mY9kH0z9wKoFj3ToVF
lOk5/C5uggsuD4H/zvwwO0/Fd2mizGr7fXmjLs5n1ClqCaJV/I4i79asjdeR8rUFxyHTGjHJv1uq
YB9bVDewYnBkvkc6QturbyJ6eG1N2CLPzrVS/KVjzitmf1SZmZS6Y7g2C69OL3TP49XW2H/zHqOX
sXo6MRtigg1keXKxQbtMckqdYkQ0h9PO3YY9bqw0nRgMBf67ta7J/TITbt8AEdTFQhrQdaOf+H6O
3yrx2VijFmJW8iLMevbnRkNNteyCykRBVByc/cgrGzASpuOtpNQSASx3M3EVTfedzV9N6l1RXut0
W89IBbqsSAbZTLQOW4Uazu3oKAqthso8ilmcJgBSdFw7RmHBcPWKkdVjex/8LXQbOV7Mc3wkfwC6
55BZ4gim8b+Y17dx5RAY9Ppn5ZX1xbBPBe/Nmt4HqrU7MUKGS0PSM3XaHeUdyZMUVnI9x1YZhut8
+a0FTcOPSI5gdaNFDCG4VpMnkPcmM4DuOCzF0z6usTiOGBuqOnW10agsnkSZxX16TeTKgOxeQLwb
ADGfE081X8cvl+PKd16jKs7Iy8OuYbkO51dvAOo16UyCMzotkgxwhZruR00KVTv57PiAhOadoXHD
8EDv2G1J0hnwBil4z1zUGz2uY2Azpa3QKprHMpvLP7BkHoRoc5ol4z249LaBnL1xwVv+IJvTESwM
LKrHqTOC0WcEphNdErIzTR39qdkTWHPOPAn3yjxjL3hMs7iG3N2+GfB4nZmQrSIShS7J4EeEaP4L
GPsDxFexKUcU6ZgMlo/+i9v9lo7totau4vN8mPMhAAf3tBQhTrFijditVVXh1bqmzA+gm3hFNLbp
0sqBQnUgHaauQMoZHzNtYlmw91vbFwzBhGzjKgMVihde6FLYWtO0f2Jl1mQggw6fM1dBIJFL1Iq8
3UiXgh1O0tjRDRBWggWyuqvSVV6OEBgimmDxux5ZNlICsC4GjNtryQvgzg04HZfd+lXtpr9uKOWv
f84v3zMx/UsjZJpEyve4x/TKcl22li0m9izYpccM7xsU6+MoCHgFR5RkRGoqqszJEUc71oBYdZDj
lw5VO+zR2Clj119yvirgGqVnZsrJckeYjCIx8SNkWUaZcyUZZR5604lxTYVqOGTeDoYR4JMUgUS+
d/RgDAiSlZqtWBb4I8FZsjxsMXoxBXj/CGpBz/TOvsxU/793X5UCvLOBW1XW7EcFzZyk3lLo3wY1
wPbkBwpP/s5mWcgLfc0hAp4uznaE8ixVths5K3x1I8pNW8XvGI7yEqfE19VcuCFNtJ5G0ST+D5vo
L+Dfz2PJ6ZSHcL7HDQcjTz9DQSQDT8vlgILw7OEnfANqg564R7GvWTDHOT13A3JVx2SGiDcvYZZm
ntMbjTZ1Ocrs0YBqm1aMmMvJpadEnmYorM0/OoMbymnRv4jExWvRd5wj53eI/plkrSagPFFZ+oqn
inFEF+6tL5gT3rBUwiQwJlnQfvFesUBmmvlDhZ+4n+v3qgimSmFF0eOLCJXDpP8NgNPllBPUoEmJ
hIuk5T988rzlAlAkcJd5JZz8Nt+g6UgbVfh1cyhEjHv0+HH5gAQ7ePb3q2uz+h0gEuWr4jx6RUxt
dcOF4fbaRHokOSE+6Jagw1ldAzn2bKPT4b6yaeawjW4tzTco/wSjK4gCOjgDUmNJEYEGPVXhI0GA
Q427Nu3pBKycoSEQ6yv6G/2N27DW6USsvXAVP/3JwNgNE8nZrsXatJOyKMZrlZvHwL1Xw9o9RgNn
Q8tamsl84k8xAJqNcxPyhBOS0prUIy8qJI0RjIIWtZ/EOM/24Me2SyTbTb9BQDur0U0Hjm/wchDN
6tCKY98fAzWvvVe5XwsQdAhsmiTi6FiHCLxPBLTIEJ5/es312n2z4PsPuWHtVwt5jsY76DswTjUw
E2BIf699R59z6El+L/w/2UE2hOVYwsY+PLu8jON1OPvE7e1dKAvPcaShQEkhv3EJY6V0OJDuzfGb
6p2y/CKLAAejSm1yj9cJV6djhb1pEhs4sLUoackg0kO7v62bkeymnl4wtCOMEJp4h7tgyqZsTQ8j
o7rnn9HBrBHaHl6UcoSl32EnLoOkMVwDHPvgbsi5Aw6kubdVprtgAee0CHGwHAUK1EseR8OIvOR5
1KCDr/gJhFEeaimMGL1XTH+zw/AlUB75qcJb48nWyg0OnOnPQ8vsuzC/BNPGJipGpi82AKcvaA3E
iAcqdKrCLL2paqjNkAQ7WiQCmE4Fc2X8ve/d8ox9f6XDySOvODdYsRe7Zc1UG1sDoudRZz7z62L2
lAm1Qo6vfKjt8vXSsi/u5S4DdtkuaIyUiViVjOIFYXaLqZHO9lK28f3fXMs8ecitgdI3J69r7H9N
ghh+3XsRcmIF708a6/+hC+R1lykt2QvXE+mNM7xTVq6ZfIRb/cRz9q/9lriZv0GaUYljN0SmgUPc
Sqxj1jgb63YJx8Pe1724WxNH/PBkkjDKISOD62X1OmS6FkpSK5Do1VIpx4wlhvelRph4LN/L2xur
WKbXSPxArEqKuXZR9U0LEejnr/td+Q7ugSbZosjN8F8DSgelJ6VaAiuZsULUJTHrufC2EXpCYtq5
S6yJ6CTqhzqiHyvTBc4BqfvfqCZfP0Xn2a5frPmNH48WyitDLALdR6iRIchtgLCth0KPuzFFTDYi
dOFbNpWs66kWiC46U0oDDiasLUiF+T/D8ktmWXT8KFBF2jnOiQCo/YSrbtTkEYJrSDtbVdKLnuzH
gp5tcjVLf0sQvGc7H0N7LOBb+rgJapYVQcoDi7YGNvevt2DXCy7ErEJMf0To6dCwpAPOlNsPyqu/
mbvD77MSHzkBFcYuI8uMCLV3omvBcvEnjliIAwXScKK2yxwPs4uHkVrDMXT+IcsRkMTbLyhx1FaV
Uf5aw2t4D12fyuOJTi5bKbBHvpPAbV79WxedIqmcTUsUzYCpiKt8iV9ixeZDNS251KUOR5IBxU2P
XxI6ADW7yUUMar1JomFwxtRFr6iH6TBs/cYsNaduRbp+jAwGd81W2VJn1smOlkHIqhhqlect2vzq
JGqb96Pz5f2J9FbCntOPPWket/SuvjE3ysmMZd5K9Z81INK/gk7dMaPAMc0XF6EprCHz3SrvhaXG
xCDP6lZoF+wpavJQhXTdnBTZcvgdEfmJdgLOGXCXPnc24rRZZ0Io7Jxue/Nj93rFzc/3mXM76Yar
SdWBxsyaD5hnWP+89dHXUVTeBJUfscHd1c/529s3u53ygAXgz2LKpyQNgE83lwpQMossmeVEDVld
BeHpMXdPuY3azyey1pMrRHlJy+LglYyvUmLwpg4U8d/uOQOpqOSHDIYdPMCfN/SXO3Bf35nQyfGV
reAkyoO01MiF7JD98bAWelkRK2xu44g8ACOlogAqP9uTNAvZvdGJxi6WqKns5ZNzFil/UCeElh05
THEokWQfO7ZRcV+dGwpH4yctISrQhEShjr8SWk7p9FQl9er4c05h4KlyHgS8MR2U8mu4Oj3IGMwm
GngvLerhS9FkTQvsIEzb8zxYcD87CIN6JSgyALY0Y3AO/h9OS77Si4HWxEwb+7ziKgw3LbG8y/eN
bIQjaoOuLGYzJaf2sOczWnejiZDukdJSqSIZDXuJAvsbK5eVWg/1QY0+xD2KhzvvfD4TB53SGpo/
o0dxdO/B6Vd+V2nbiwuTFphj8JYHZ2DiHFzaEggh/5OZbJ+N881qCi4uUSBUEZgnn4XTG1yJLQNe
vYlmH+MZaNV93/7M6vV/rZJPlofBwe+hveYyW9u16P3fKN3qTIaPXfSOOzk13ooNBS5w3hiWgDX8
tUvegvzXs3R9AZdESeUz1qLKFTsJeFQZakPh0pp2qy66WNiMCILf9SNuNBh5ZUE21iFRRY6nEuFZ
TvyxPjR/2peCP8FFksp+vTDKwVod0rCbO/cGXzsq+laVbI4UCVfDqEb/4CRBSDE3L5ToygHRx5LA
q7OmjfGtTamToNzt+gAImnBu4GocD2vfRLuaz6yAXP0mzvLOwR5G3A68Kcj+W9ulwzlAKCE7QnSk
dhRaHo5wQdBSQfpccIf9o+gwf8qJKSBYU0Ds6rROY2PAUELIkJeni7MN1z2wKe4BKR6ic3L3sJdI
c/KzJkVXAxlHMbKhkYyPSGEwfhJp6256YTWm44jZ8pq8icFYW4B4M+rrAHQEA+htchpHinJ+4GO9
klb4fkGdyY8KQtHOc/TvvIaJ/eWAfltmLBMvDgbc6w7rLcEsoZ1xzYLzf6A1JYjG35Tw49MdFFzT
Rvz/M7Ep+ankAxEqwtKlV6G9HTgDpixFVWj6tUS/dZ9xnNY9y+ilQWPwZge/24HbieMeln7VuaHZ
eQ59HBdaqCcAQIivh3uc64D5534zJPMqVFeD1sk+CK41EnqH4lTETYe6EWIrI9uJE+ukt6f2rdXK
dJZSO9J4ALfpj//+QnkQDqo5i1LtM8ANmNxKWU/lFciH/pjIMLFuRwfD9oWSGv7ufXfJj5G99KYW
MH1Y+8IKuuWHx/m5gh8qF/fef3WNcIjhgfa33vjbvxh73cD4S6sKb9yBIVgAPBwQJTaY09I+7Ge/
bPIHBov/ZYZLPGESgpETTu+VAE6L7nda9aGnK9lAnn8tH18L0G8IA2OzDarw/k8fT17VsrP6XcjS
NzC4q+TQaJXBsCysnHYoZH+UzmGuwXe21L8CbHox7Hh4Tgh1+dxhBJsC2rf+EozJUl68JnTwMKyj
oO/wd4NGEtY5rCXGngqcxlzIOOjTf+/GENmgRs16upQ3jBDdHHQJd67gdV0G20VESZh3mIFBzKmZ
lKzEaIy5K4/z3e3eT8+JLF7bmQHcQIknUUvNFvfW1xc6S43nQ1SL32MTWDVRm+SMK2H/hPbBS6CJ
bhbK1PMK3Hfx8hLUHB/1yeZBTKmeEbMrrffEmZ6YqjFWKq8NXxkP1vGdl4Vf0fIHutYNJnW8xEsv
DGTopKlwH9p5gafmPUCYngGM4AomNQaG4KqY4H+tdph9rqjSBkwJzWjhjJL4PsLEXKvmHd/oVP3q
+imbOTXYZZq6yZSRdB2Hz4j0j2sdohUQMIgXPD/sgkM5IGi+0ow5JwkDzRqQa9ZPPAwT/ISys8jT
2TLQk3tOhvYI/KvSQp0ZYlG5owqYO5KAoZUit0V3JDy5EQVlMSH5SX7Hg7Q8tFS1gZM/fu7TeK8k
NvT1PwPYIe6KEH0Ab/DcPKYxfSBjCrttdl1abPcveud4JF3O9MxcmPRuo6E6ZHvydGNGAqqgcfI4
/w8NAIshUrrXsMA0F1KQsB0Rj0EzwCaP8F88Km/OEeZL2cBD6ZEd9Nro4p4JfQIGrk687Tw4afLv
m1z1lUdKxE2ZOWCpaWFT687P8Y4hhYhVPNEVqu8JPvE7WbE7rxyl0FnDgMAXTQPiI5BsNavv2oyg
5rUjK6bpfgTXHvYVLlzw1BzVvoH5K5Z3TEK814nhHTYp5UMkxXejRV2uKEmvBYuXLbNUQeNRDOva
cLbRx+sBEFOUAL+Dj9z/Apr2pZvOrGADRx3BWr0EFvo2yBfKpbnTLqHnI53c2tqNui0tVceDNHuG
Jy6dpE1RN7TsWbZcXW61vh+s6EItXhtJ1CtvJnwXXeLr6om/RF2uN5Gfj76w7uRr17EalosHKloI
FkCGUBlGjohO9fkdBKqB7P+3vncdquDOnnaNkSDONSuLrrXEYZlXHpG67WgZ9xP69bUDlaKetDFr
QYJajiGaY/1HoKRdKk5BYNrBtUmJEwiOaGOxeoLeuQyU1TqtjywjiZ0tcGDYwi9F66Qy9UE7QUPw
VfZOaziGt20z2RcobbZKdRY1S8fU89DL+EHOe8F4rNks6PrEywcXAaj+JSe4NkXwzSQ82AndI/f9
DCdlw6Ij7etOalovPGj7HsDaf4KPuO4gemuQuEkUSr8bG2hl4LN371thHlh8V/g5vYIJzSn3p3a2
yyshofBhBbv1/nFKWFDDg9V0eHTAKJziZ90VSltxjn3BlCX7jRaBsm3yepkvsMZtG/5I7wI9ViZk
qUwWQHudHkAuAVd5BjiroXDJ2NFHo6zUJ0l+Jr7CK29RcvDYoxNppVE+FqFkotEevb3zFpCwcnFS
5wAAUbr8cNJcma4j/yuUlMeczlNeuIR5SKW4TzHftEgN++D+0Cj57iBYoMwmCSEdKUNRJqLE3uac
7EcLXaQjaE1xAVmeJxhaGC4Td+ax5LOhLkM05NONXGmoIDRv6BvCTCeaaFhdbWYNjfbNEDyO5ri8
NuDPe4Z7X5dNmOuIgVvGtpIPyfusO96l1yau6wG/LNxbNgVFh+lsDSFeX4DqsWzcHhFnRuRHGhDy
ASSAon/U/s6ycgbEcjhCvaKLFyTH4jr3WTzH8P1UezN0FDsdSe+xCn8uvUC97g5n9X9BKjMOcmYV
yvPV9Yt1w3lWp5k+XJo9uYl2C+bur59y242kRpOOGhbdfPJb5J5tBN19Ei290CKPDGycBAdgsGbd
C7Gh4EhAn1EEece6jamde22g5VFVKMGbHiOugfjeVu0flZTA4CS8hnaTUourrmNOSLZx59kkmO6f
YpO1IpAaQktn59Lh5zZyOe3aKx36U1msHRcUIJjHAzyaUjzsXa7X97BJ0jBpPhFBEd2lACRfkolo
gYurnE5na+7o7QctwOEtNrvgAYybTKZ/wklyQT5llgIPzEklEzEQ4936ycbSUZ2dsuhx4fTGeiJT
Imp8+0Xs+v+AjiI6BNQsHI1zZMJTXD5qWNcsTAJrMdZhM//EehnJ7b4k8v8QuoIVTrryadNnkNUB
vOWpWAEpDEsMgY5LcALjH+esgCUIL0LyDZ0G10kPVG+Dqzg0AVsxlK1zgDTfhJtx35AO/s2XxwxM
hj/2whsyXRC8GcTuJFoRgYVQIUdMIFWb/Y8yFEDJfJqloCN4Np4PToXMv4AwkufTkrolp2OFEL9h
T9w2ZbDBVDoSAapJmV96k4snl3UZkJBqxCku2MkXAnF4e6qnb/f6itveaAColZchBB8xTFSB3NoC
350Z7F+x/mkdIGIgwHYs60T/238NxPL0VCTnGXGeUV5AAgOH7pUN4h0p/RSn4PbdtNeGrVRBZI5N
aEDVmTK1m1m/tQQdR5BFK52aLCDWi4vz6eFBBTlIhv2oKc0T68vZqNckGd55Ll1HsXFbLqie3IEf
R8bfpcAQW6DArydHkptT+uqKLw7t5TlK3dCW487coW0HtbPsn4yYJFfsgYdD4d5I31rWN5vb9rER
+C6uS3AMjuSX0pu6sKQ8cTQSPR2nERlLSOoVIM3AnrHxo/OE5rXdR/PNHQtZ6ppXjZNvCu+cWfmh
cu1EQIvqcQFDAXmaZaRp2tXsfPGjRWpfKs/lVPdJYW3xMDB268RQiLvvwPEri9R5HumWIRe4/HmS
KdVAbmXO9AnlGE1GN7jVMBoQtbucc9Wym2pLDvo5FzngJhI1VlDsbMXbjt9B1fmUIEHcVKNWdfKv
sFrVjsf50RmCKkM+IYkjvPd8tEWdbxqvZjIOGJtKwyJlPQtCX3/5vdqnriHndsTR/GEo0yzdUiw/
DBgYhqsL4J1t+2F+TpwwHvRABT+By6vWJIxWIfYGNjRjjC9zCHuxHt5dMta9Bm7NM+UkWq6gUy/A
t49JUMfw8qozYrNI7acADvyjjbfhABCqmh0niVIOnlbzYIrGAK+uIcLSf5eSWhntF5w6LzAGxs4h
tS0Ztq/8iKaNnXqoGdmKstEeKbFABugFOVhaUOUsxxG1ar198YbrES0AN4jkWaXVKDW7ylNF1r93
G+RZmOFhlm/FeqeFRiV0XxK9acSItri6V710SrOcKzqSv5ukJGdTVs63KGhk4gUs/7vRBxY8M80r
AFbztcHau5eNbPHgQhFNCElA220btYOcRb425LBAKFzXbnQ02XQQ3RkgnOfqDnoEsAj76c2BiyXH
5M13Gbv5fa1RNHAlmJYKiVsXMwWMdxOt9483nV1oGAz+M1Zhv0adXBYc0nAN5/51q0uXsJdpaKQ9
gnvtsz8hX6hElCYb+3nwg9O8zmIDrZwfId3hlzoFWaHEiEF9zsH+mPoaoil/XSVCTeG9MGPO2DN0
8HSelmRo+54Dm970fWbmjTCxpie/GCaBdHdRkybh9106fezZXx1uGQTFg6oWB7fGMWLdZrJdw40u
H1XzA1hwbmzysca2X72SBmHi3/7RxiRkY5YZKkmy2VjCbfiJhF3DUZXDuVj8BvhnlmgAbNwNtrLb
CbGmrZR9IVCs7mGaNJW439iD8+kO960vb3mdnof293swTD1MWoEexpFw6xL4S553yFtwyarBcyVj
JctaHDx6qWA5Epbhg8kKaZqv68pT84Ehw49YyVuZ4f5Ux7pXfF/CaN/gIlSEI6QP65wuHV3E7FCR
+Z6POOPkYCU0quv0lITFiHUWtY3jQxeZs4uy+wpEO1uwULxeBBlQIphZu4dxtdwimiY+PUzxpJPl
5G/UUBkEW/4xGfeYKRklIh9HhT/9TpsnAkATSxH0vSWgozBD7wl1JLq/IPRgRz79ftp5gJXGqN7f
iYhJ7pdXye0wXMmtMq2HouAL8WqfAI3FFOx6PmmNaC4oBmbkl+ABbCa+r+DiBmVgvChv2S9rEiWd
mswkwzzafYPScD8Tkr+fQ+go9pF0DqO17z9IJqDzrGol4y892hnQhtn7uo8jOa6hpy3FKiKCJgir
X7Yz6qYRHWRT3tn/seqzKSAfAJB8Z0THBb6otx4Wp08u7oqOAPCAkPi8yA3btXdGN4cvfuf0/ani
kXaP3WHCRVkGy5f8IesrhTWHkaZeCYukDNxxI0NptwKsH7EagoJfdNPH8Sb22DsPOBWnhMYK5z2Z
5JiMXm4pAq7Rd/pwFLdmuDqj1UY5SP6rd6RTJinAO4CmeWTzLZD6nP7y6Yi2il/DufnfG/p3cqmj
FYnPjj4FszRkLBuNbqDYHCbTSR3Qf4kcIR4fU0rdJivHqEXK6VBAeBDD7tmGoMWz7lw12Bl0piLc
LsHYWtT5lb5ZMQ/5e0XEm2Pjlgojhv8PMo4R6C51PuuImwKmAqjGn2DrRu+occuhBI0KOYC5tOVE
utAHgTFcisIgj6iQ49ShxHjy1Jue/h9uEh/beWvfO11UkVqjf1AJzJMHC/lZlfwZ0sUBDIE0JsNd
n+YgMor2iAFWonm9gdBEFOh669ZKtjFzEclpM534IypSLFv1DSu3Kez50pGyuLli03z7tGaNjigD
j6K+pGE33SnAcYV2l26Gp7S5DmE9bTDpz/josIAv8WHuORoFOrHC1QKthLeft2LLKeVQq6UUGHD2
3/3bQIG52FkecLhcgYw+3yFmVODhDT/wviXf7xYPLiW3mXjbvOZL3u8ovok+78B3xV/nS2X32pz5
b3ITUwPEiDfLKGxGSowDVa5lzCxyeWhf+ruTLedt4crWpp2OyRHCXQtQdLmAqDAg+CsecPTNSlfy
JucPgoIF0RZtmyGfyLb74cas0FMs9JN0hL+ROlGsk0R/LlLkKdO/E7Yf7or0yKABYMF3TbNnWftG
vWzzBNpZ8ypyH3UdU1xwV9ajhOz+h+EftDXCFmt/SQtmSPcPQvX2vUg3GX7dvfFp4+TNdYjFTLJO
g/2hg+GrBtm+SCEyPTAwuymfZ2fT49ARYmSnwBO3s+eULfL8eRVvHzi5XXWU2EYbj8k6JLMCZfl0
RHxhCeanPK2XIhkylQFjYUg0YLIy2qqQu/TPGsmDk6hWXgUqpKILCTdx5vpRjhW+rJFm64o8ImHz
S4FawHhlAC3GjKWxc0aqB5CwrHpQkcDLmUEXSHDR7FnyAZXIKMMNOp69R+bH6hexh8VbbzaARxIa
sbdefCFSIxCoC8E73mww+YgM4ND23gElo3dFd0DcgmAfDIq7Y5MQ3LmLmGvwSvMKQ8RJ5Qnxk2BJ
3X12MCyOZy4y1sRun8sOYTk3GSuIzmCteXV/FLDboBgGjBlSRirKVO//kkOKLcan5iAQuqMQqHi1
Nn3x2Dvwk15Q4uCxomjfSdT1Ivh5ZEqOfiIe59xKtZZzZ5JR1Ogm6CVvtS8seia+UsGflV9hm7/y
odlZVWKotaw1BzZNOrMGPtlzUse3FFOCXQRlBBzhBIzZ7MuzDv0TqgMT0+3D31YOlyCfxkEhsaia
qWLwlXZdfPcAecGoCFMfN5v3PQ140weR9Jk+MtHEisQ07glCdOEDHZKlzRP92lRTkiJs/sVL0Dtr
M5ZMaWb5Sj0vLdFWQU9JZjfcg9hPWa/+nJOB3sTNyeTxJdR1ObO7PUmJzZVGpe17ifTcJfmZkjzQ
885in6ybsp/sG0xmOqSWcWSgkmYnxb5dnOA9oXPEu9SKIZhAVHqOEJNEsF5XNe5tuFjDjY6Zpz8g
f/48y0cgzmRIi59klOwaiV74BPem20EyCUqpA/Dfa1RGuqZ/1gFL2TSeiZ+cthasHtnaiJ8/7lba
9VC6VB+0vjVAjmCmigyBPwXoBNqYDWEIzW6wR8QXPFGmvHrMJargBLu4rGMzXhT1gxdH8QLlCloe
sdLVyLWZ/ciUjcJP2B+kKsDG7TYubuGEj3Y+lmTFwgiwnMONXnhJ/Q3eRTbSaQLDWQFIdS43zp3/
hrRdtjNwS1gWgYMptWSfPOZwYU91TIv5qagOLTcdCOV1kKWoXxYRXS17T/Z3PXLo8VUi9hiLpese
XiZM3ObdEGq9MfsYJY5DKynV2bJ1WKGsWgwi/IGHGsd0KJEMlHDC6EgmEyOlTidFAdGHAdGPsGqb
lejut8rorvS83vF0uAXF11pz51Ha87wCP5fTxb5ZtyWxfkkHS4ql3tsykCKmVVnvNEgLJ9qv9JcJ
/RJy9LDAlKy/Hz885tAoEoEX2YCK7hFSyy7EpwXBrtH8O2JrJ/ZdDe3Lcy2h4vtYEwVDcH6V6Pjr
0qF8HSPaecZvlIOTP5VwniPT87DpKWT44ZrMJzWizPg/avYD+lRaaf7G0DTag3DFz3E1VzaDxFKi
Qn1BgpBMYvCbzIvhH3eirw/fcfj8LwQYdjzksEz/B3Jwm3E+MzLOg1AsiV4WX1z1L61B1KxsLskL
/uaaqXsJWbFmXOhm/8P5rSJOO4zZqciOJzMZdfUyCDDtPOGX+RK3fydNeduIo486NwC53cI/1x/B
Yj36fbSiJ4YGG6tVsSpeq8vU4XY268bbNmZOdDXV1iinKzafDbfCMYW6ddV9I5QVtsKU2FBekb1G
XBbtyj0iUFuhBCkEJXQWUyXNruVoUFPFvSRllbLUqwE04Y+F6wtdYvI3bj/wuCHNBSrXBRlbQ3va
zLH/VKm3KJ0Q6rGdo/jTKJ603b1u1Dmyz4yrDlmItFv3OO79h8SiatTbkZrBJh0se4M8i54aPyGi
ImYCde81vXw3p5BQbAECRtDjttSDjl6w/tzpoTSCsXEl3uDzcCUMmproQUKvjzBdpV4ONTSbv2ou
wFWz5ahUi+TwjJKf8B2rkkoH0H0NB2j8dVIsQu1WQTM2K4nGKlO1gwk8STo5pHzR/mKfar8gt9bt
XUxadMWeb9R83IkPo3Bo2OmOABHZLaF55IfrbiHUEzrWLMPyM4TUriFNMZz7DZGVTdGsFjCW7RAb
goVbwoJTCgKUxMcK8mWv0/8/YOqYivdpbfqTKSw/WxK/6JxUrZWTG4injHvA0Zn5Ir7c/hv7GAS8
v6pc7mY+1sd/FvddRw3Ro9DZWzz8Xj3F1GNAH98aNBVch5MSBXQ1TBFSg9mcM5jAOzuFuuDxPMju
uGjY5cd3wZnBc6EuPpbAbhBk4zZoaTp/C3hphRgI/7UUOr5dcHh/dKpkIDHb4UpAAEBQwImcuxF0
Mma0VK3odKaEYuCC7aAcxL9t8vHyJBchdzD0M1OXd5/rswYG/8/4IdrfGNSkYLxQC0uqvJvisnMU
GcZjUTM54+dJKifMCJe9RX2Nj0vrT2T5JMWPlK7OnszCI75K7Vo+KW7pZNHG12YLjqDfKB20m9DZ
+6K/i5383D5xTo0wrrJdWadqUpHE9kaUYOO9LWw3WWCSIQTIw1NNPSkrGs2IwAvxLhyWU+44CJ9o
Yt4oQ6gsOlli7+sZdRCatqk/5PSNnbxdyw0ax8BRjNKVLXRUuNg809yFCuQs0/udivZT7r6eTTCF
L6MTmPhqbIyn5hYQG5wCI7WndH4fSF1I0YQ3XuCtc2oC2blov25TXmvM63W04MRfDOqh6Bv9Mp51
eRW2vC7yBk6yFtKwArSf73MFptbbEfHL778hiPRtmOgyqfM76/8noPmQ8uY10B6iPN/hmPXWmpJH
GicsgdZddkJUxnZ9dOxh/0KMCpZJiZ4nTAu2SNdfUik7+GRf+jgAFs7btzGMNcpt90r1EWkE5WPW
W0Fj4aOhK8/EpPg7ROYob0oyBVm9q6/vc2ma8qGEsN6enTwylyA2eS9NWLZZxYe7TyvmaHmF2YEl
kOdy28zqoovaLZHWSkkQ/hPUzBB0WNdvTxJipjLGIbKzjGuw6uHe0DYztfHAxfRokDXEIWtH2rQ6
URdFcKhj8Q2ZFSoLEaOY81Z3wjopjKpT7aXXSxHbE6rIGraqibgToyrcmGG0PUM64oXHaYKVSrR9
pNYlxgMOwCzwIiuxBxR6U2Xb80NSheu2bNP8t0sd89DzA6Yyw3lDPOy1uGDjBoEHqtHGeLClcGRr
thtK9G5aRRniRsRW+S3WISp0IHCzq+jfiVXxktsFW5GC+RkKwTXWpiEr9mPi2ebPDh+7h1u1+HS2
Hx4HJgPV85tsZg26oAzMIU1OaYqArg/wSliC+bMzp+tY7OC5myfJTJs2ZElfK5J4N4vKZm4iI6nQ
pjG1mZ6SvJeO142JJbRYHvaSSbpYBwjQTExabCF6QebFeuBJLYdS9uU86kbkOxds1qCpoZdQ3Id2
A1G++a8d3Us64Y7j1g99cFapTiwr/TgqlK01SmfUxQv51M9CwLD98F4iCpr/lpRvHg+bRAS7dzkB
OJ/Afgyybs050RaaLBaHWIzElJsXQAmjegYJEqgPEkVTXt/O70MD3M+7ikNlAVRb1oS3GUQ7P7Tm
l7BNC9ENjKZMk2/CLyOp9HnS0KeIkHjJolwXUGeJHjj3bg6Yh1dcIG0eDprbLieQgp2Z0slK+2wL
AxrEE/FMkA9TQ+LLSe0zsBFO1qfNxxX6EjNdmha66Lqhvd0UqlLgtZOp7nFeSJLlK1hvBh2KA9nj
S/DrX3S83y/Q4uqALq5jBUNzoGaveH/aebvkPZUKD+x9HJS5XXRbSi9x0yF5E/k5vr2u2Bla/QrF
cTnzzBF1MVoOgTg0F+797yjXsGfd4IpVMFZhH56Pr6368uQdvKvm4A+CwC25tJT/KgSdjPRUit8A
5byHHAAaRZkbdJrLfq0FUUB6aDmYRh2KKO6lO1s8U8v5QA0ccsgFHb1Fl3yJwJnbKfeC2PHS/vgB
4Dwok/ApEJmWpMhzpMQWUQWAWaad2OoiqWLv1AGMTo7CZi+RzTjn7il+BMQ0MhLMjZX/r4NZVroA
p/WGEMXztjXvvwHOeV6SzGxucN7ow4hjXD1Niocpyp7p3WlEzpoQvaTYKTXZjOiJCJSUhAa12pNZ
tzbG6lqiAZKdH9ZbBRBl5ORm9B72nEEAgzdZLGBi2DVoBJKPid3eYDsobMrsRuXg2rWEDcgpNfc0
/ESZ0sq9oEVEp6hODOjxrhaEFMllCJs4FK3owPmTWgcnFp6iUun5bYA4pG9dFu2bP+lXtp1vA8Cp
cLlIrphHquuS4cZ/JQUTRlbzPe8jv3Pm1sowFogSNA9y5He2ihvLOXnZIaDSfX7WsxEIyvgC5IZo
kNahKANVcdwUyCYi5v3jobOs6RiaYYYK9QMw8SpYgT3ppcF5dILUBAkMruTlhxPYMv1VudG7fuZ+
TpRqZRhutqEil2fAGEzebHI7VmgDlgYJ3uQCT7m8Y8wQYVC6mEwwKWzr+svEUIuInV2RlBt/crRN
j+fUXcfh9YmR1M00RfIGN12MafXdSSuHhjLG6GhK+7/HGMQVOHc2PMqVxJGF5OELD/O3kyjOnCHy
k4boTjeqx42m9A/CwL1d06Ww4xLUF9X4xsNm3MPTQufTlhKlJ+8Ql/0PQrW2dmn2otSb2aMnB0f8
QnNT2MHO0t5vKwF6CNeUDiOdk2J3f3BkIEewvtfOJLLseFQan6g3vGl1v80/S/eqYndPq00rth33
I1VDQkcxMcmgA9MjqPjpFimTsrcZvWgG6B3UHA0hMlfP2ISsDwd7niJTGujwLRtOiCCuN+qt3fUn
i40Zn4hNl67spj0F1zGLE6ZXml/HjH3T5WcPDL1Lr42tEeS8xZXICxqCE828KkKQjDxzqalGDp4n
slumTFKOZ/MGxNl9ZoOpGD8XQUunOUXymXPs+71+x8pLcN+fTI+NOKi0m4vOBJ6MCIjUcqedFkSE
KpgpZhUjRaDi7faqOIMk0ZtReq7j1dDiJ6/50hWiu/rw+tdE5Q84aQ//YfIuJDdQ0D3q934EWBJ5
LauXyCp8KdInu9m4tAV2kFQSjJlaUj8meIewEPgW+ETzLBwWD63xAE+yr5k9eGPE/6+IH4VnCZYf
PMScx8uCrwU/6I50b0kG3JcIY5x+ByHG3x6+siNfIt8RR3xJL4eSxI/UIq+XwGM7YOMBkR3SPq1k
/SBiKZHxCgyp76/lgiq+xxIRjjDSNzumnzU6ObdqHw6oyP8EQxG37rargaIn5IqI7Hp4wJB8x2P/
b6UdvHw+tArqKBInzoYJgRRP8dFYNZVM/BAQJTPp4jvxbMJlofwYiOsYnHeJMg2gLpFxVzPNK/7X
0M9f5jRFnTRWZx1qQ4EW2FGkUFjaCUCJ28hWVQ3fULk28qSEm/jY3iUR/eWpimC/n53j/azmfqJo
JSPbV8KbryJb/76Hy+vrtTOM4a0lk1mW23dRo2dek8syzPFF1c25xULzInR8x4BJrcQIbgUUfl0J
b4bcIAHw/nObLwCXemiOv/nqt6vRCUw6Q331+SARA6G6/tAnX5kACxALftV+D6vjLsiJPBtnffZU
owlmZvlta6mQtHz4PWHog1AinsWHh28UUaBFLsbF6Dv37uuAHS+evRwV6Qx54pFKwpjqKCeePZH8
M1nwnpnOVxWasuO24ZXhD1ty6VVNBd2ZhJqXXfRCBZzHdoMDLYTr/lhDKtDmJGaBOkO0/30s2kwI
n9G5KQvFlXgJJoz1aDEwmUVtmEkT6SaxSfGP3uU0dhSKilVJ9bMa+FDgFbKxGLZJB6gYU2K21JML
TB6UuXf0S7PGSFiWBPkNP3bgCbGMpuKjYZjTNVaZzjMREJhYR5a7odXXY4qRr5b1rNG1kzIAopVT
Y4BJG/SQ0BZe7412mCenGjqGQCCv6y5OWSmdvUb/LnvtUFRk9uFpfORd3TomppJefQq6MjAJEIm1
vycy3LoydW5DtasvcwJ/b0YXCGqsTWKm/+DM/oCEOwFDx6wq0nt6JoQwGa/Z/l8UMUKlvy7LEgzB
tm1wOhEIrRLtNnQrj6/HhKRuVQM18M5eiGpmkUbm5GV28P4R1FOb3vPPkASGeSDolknMds97KxYB
Cg5Sq32qRv2FnBlh33PIVFAoe3BaZ76F189qfWbMJQc43gayrzF2PMqTTqV0R/t1u6AyarjOEW/m
9rVFStqtmFNlRivgupO12BY54abLHlF5l4eXWxCb1G92bsKBrHFwhkoyeTJ/SX2CtA/K5V0FIhNw
A+zuwhdQtXY7BwP/vjd0VCXF36QkLHDAkRcSy8NLpiGT2gojQpyi4kHO1aT8s4EBrTHBC+PbnDhM
n6ZEZDY1orjswanoiDo/wRS8w+LAybBngLqQbI3rVpf6bcPo0uHDgn/nV9G8w7Wff8MrYbVsitJI
MPvsWrJwodw9a3EpzdtVUf2pd4EdfL8RWsRS1WIb3GSuOfiAwm3F8OXChNtIvIujTFgBtUpqqros
BgI03H1AObkN/PaMj/NouDuKvrDJKtP1rYfzie1KCZYUth94/U346p2Gy3GuDIb5a9dsqdeoj+gx
6V1yCaaWuSZnwQj4v7lOOsaA1hMUif/udCBKtxBiR6n+HY4bZ4pnKgEr4xnDNuwbGzWWsPtAljzJ
IA+hrH2Sm9o1P0yPnrpO/2mMf1Rp1usf7H0XgjpQhwVRorQnqUaF8zPNtpDdWPc1x5vGRbXnsBji
xMk8KhG8UjJM9CKrwt7njrz9uScBkLw9oQ/17zMoBOHK9JBN1HFS6cGgutpBtRxSoxSWEuvu6wzE
7vXQsQLC9lxvExUEzblqWuiAim0XcgnrTEp5L2an8TU1wo5mnGPGC3HNRaTjB6iyCw3lgJ/byGjA
ll/kLbKPGEhbkTtHRuy4anXooQq2XqKOVCJti+tPfLIj7QKnBTaPmkOSk7UX28/PXsskcpWCG1/T
ZGcLLynixgV2ycejwO68VCrYAXKVgqh7OGGECr+rsuSDftTkY8IlIigh4o9LNyNsWTUFpvmvsD4y
8xCKLN4XbeThBOliKh7htF83Fd8nN5RGuitJOz88Iu1AqI1BeGgkmu0he3cHk2JJBCJcJ0AgAfPs
9wOUFpfbbniPHf0mJ5q3TaHjnOrmfcB6PEWNu9nkedn87EXfirOPMa0ZXqWOnnLIN8iTJ+cNwzg+
WWsN9JMCQjo+8i0103DNhR/HwSIozUQOroXl+qs/hJVO1ilz9B29cfVqUE3bGz3vu/VZS/83eAx7
qJjfc+RnCYhSs/f60yCaGY278XpG+zoiAQUXpVpUfTKc2SddzSPkr18uSkx8xQ2tzOFpSNFbe38+
B7yoVG9PbbJa2j/njJgBaem+wMCsjwqjSS6d54fpT7nSYPiNSxaV9aQa588XlQ3u7PQxkBld6pJj
+LmF9IQKOIEVagUfIy3out+yhXqGsoIaZmxIyYiR+CDo1wksdW9yAG8I4FWRBWlfMPfbMV00ifyP
N+31cLWsUaUs3/zUNpTuwMg9MqzyDWpo2tdKQpms7rOnHi+jV2sqsN2ZzWULlXbe0Nxz+vDSKXQY
UTWYCrwbNrFRhr0DybnWR8i6e6AxNKfMeEKE179qRKElJmhZJiKspbQzmIpiTFUDSoURGwdlf625
7ncdil5oE4N1VP3k3Ep9RNiuXCKLqTadVyKaQ+jGShsPJbmMFefxVp51ACwKF7WaMzZklFyJeMLe
rrMxWIoKdIQdz3ADSUg+2D4Z9wRsmdX/g4lZdwsQR7/JRwIaU4+d9XnYk8ZZoi3gS+AhMBJpBwMj
vL17usWxWbgt4ro7s5RKh2KvvBDg6xpNXYJLj9AL754a8jk7+JFFGI+k6UlrcwX+2tULtB8XISk6
LY1oCiUnL4iFO5ea12X4baRi7D1HHB82F+5ZHVo965+/gfeiCKCc9a3OqkZYwBqe9F87A88dAsCG
owtn/xZgKnkqaFaPblNbSZBKFpx8H/FLnzh856nMNEcVy3/Z+SnZUgMsKs6rM6FTwGw+nsXDjWHT
aTI/OnowYUmvp7DGZ46c6T8gzGjij3UoSTwZSuRXXZqezZ450bXXA84QIqayILaNI8Ljd0lornG+
XmyLuiA+iUNFw81yojm/6dOyBG3pkVyiq0ICwnjf3wQ1EoPE8NwV/xFvtfmI68vd1jpcNVu4ZqiE
xVZx/T+BO8Pdf714Y41Z8jrrZAZs1MVpIkMuz5zoilVrzdMvZp2fGXYroCwYXUscu1anPuzTWsVQ
aRM78nngOwZr6M44vscZ6uIJboQkVd2WwF3A2UREttaXpxLKUzKh4Se69avQY0xySzr3gYG0bw65
kBjXuQgvZYBt9Uv2MRf/lBeTnroxY2+IlLW+TVcEaqEZ6QpJvgbskTUvB+kZNZnYB+V3pVC9idbv
LjGlbUxHUVno6nFXOS0DftH1rpFOcuyMkiSGo7wDIp2fK64+WWbmAQLYOlOEBx1j+9jZSKKnKIKx
fiJO1F6pi28+xU4Ee1OKZvjDHxWe3+ntY1ab6CS57qmbJbEGiJoBGbTqGHK0s+5FeAi+jB0eMw3z
enSTkXrk0herwSVXhdECeNUYXk07irfYQ0F7E2mPRHahaULAKhDvve1kVMu1XLUdYXmB6zfjs1up
2dqr8arcyCA3Jjv5P+CSXkGqLWM90/EXo+c2ELAEm7XT9mtVRkI0Wqu/FebP/c+f93lyzSowUikS
xXEDiZfgS0f8nrtzxU05yydiPuJ+ctaX3NTVZpeeOM4a8TzpeLJbM8c0Wv3gHt8xgl6gAV5dPlQP
L42ouw3bfX1jULtqzGdhL6Jpj9LSbtl1eSjjyO9l1zi4qtDv7sX352F/3guBeZrXade1vgIAQqSM
lAgCamzoVKgpMDf6HlyTt3soFrd+21EA41CL4rJbWc7sRwCsAgd/z0mx3xVClHoSwyYDlC+P9ecP
rpCYQKa8C7TxX3u+wDyePBb+Nq1CeU4Gios9/or17LWKGX3/pWXCKFOJrCXD8ZCrjtkYXlDdaHzR
227c8XvzsfRPBgodUK8tZY/gPvhCDfDaUXQ90fLsx1JlET+LsbDnafeBnZBIC3/VIx8c4dtBYemo
EPpHGYwZ0jW7QEVQhSedyoBac7A/7ynxPyanQRM7K+R5Bj2fPx/vPZI5vKP1X4/nylLnz5sxia7s
Az8eqzV/B8KIRIMn2hDU2F06Ii+gPiKlPEWpfyqzEAS/nDAv7fFS9ZL/ylVG1/Uk+lbvXuE7YmFb
0ogO61cjA+iimObOTlZevXD0aYyiuULmu1U7JbvVtO5c2RdG2Xlq3ji5qo2l72qU80DUETSLpFpa
nwneXe+AoGedn7wi9i2asINQ8Hrq+2mzAK00SgsL3+wnv8D2QRvEkbOTnTH1ZX8zq52lNjWlDUCM
gG8kvTRkf+Ucf5TyuUTL5wOtI1M28i1eLO9cHpIvdftiup6rlmdbDINg96cQCRGbFt9xrb96YbvZ
iafewKol/ZayBbvOmQfa/RujF0PnUjvtyHvvEO6g+5/7QpCItsQt0O+4Kix/UMrgYijXtkLCA+UL
fC/dD9b5ad1HeGDZULv6nln6k+Pjf5X219vmcXb1QlYxmxaTjhwOD+b+IVYl3vMOdNCQCgspOxQ3
5tyjuopqg+p3X4NiPyDKe/rc4bIt/xI8R2gTBi1TcGqbqNwfhni2lDexDNyxYByr+H0e0qsMwkwN
rbcg3KKrVTcVEl9FFmG8QeFKU1EuhcXXgxkMIC9fKK5Isk0f6+bQMmHcFUtWW1ETG8X/eIq6+77x
zviCHthCp7wi2eJo5eFqeHVXBMXS1oyEWrUNDnGuCqzhS6eEAsOSJzo7FUlNOsXYKTSvorZbSRhb
Iu1pFMaKhP/ZFZzt+m6pYNs86W2Ne9BoDhAIq6BHTJX+1j3cX4Fxrr4F/iIBH3QnClQrO6Tv3Pre
jSmi4ZsvjCaEAfIQWTPETst+xBWh13OY9Eel3JMTErTH6QLyqATV6knDH1MdxfHRRqAwtM7gBeyP
k7FyTsea/EHEfNGRtQ8Qg3ywGRfy8Cs/Wz5sYD/E+nw2OA9ibvMsqedlPf92uFPwFLjA3GiiVsK8
0KNplInE3b657S0KSMTxf95hAcn/L0JUY2xioPx2Pbm/E6+IrR5NYBWuPiucQV5e9qdhaLteFJhB
eV/nXDCuRv30xJZjHdSsrY3p3hKGZJUki8ZM0yN/U3AJxd9iRAsG6LRzyo9Kpxxs6BElQcIJwhlE
OTnfQ6CwwRscIIRUI4ewznWbRF5HrOJkvMrI0pCW+jf4zt4CPOWANsIuRYixOLiwZtqMVVZnOD/o
+9b2io1G91Td312kLmYfHuxC4RzuKfgMiCOpiM8F4fCDgggtRXwS3CMUYfgElOI9UfVOFfqNiMzw
QyA8gLRlI5Nw9CFM8m8opWlkRhMBW4nBoSvwTzQ4AEGFxusd9b7PEpb/jmXAULxLproo4eL7pc9s
PUNtPFGc8YYl6zZtWBdcagFNHqg/ip7qva7/XSoAwHHXfAWlcFGXBnCqHZAPau/bQy91TrzB055q
DolRPvbT1TVxOIVeKgzPfs8kgAJ2IIUsKK584AqRUj8o9vWRbBTdYDPt++VPgNFg62E1RweqpEmn
YKHvakglCH902mi6IyAjctv1y3Euwx2ZdYz0nuhB8gdAasM/h0yci+6VuA3yG+3wXcZ1usgkZ+1Q
dYutuQV7EGm7HOlZNpuH60mSEPvNChvaHbIHz64fjroa/4bPiSBy4XERJSptxlu+3lHqz0eYdI7b
8kXXocQzTcGiGLnunCGMHJWtMbh4EYx3LfiStjtSkkLlDx6kQ2N6gkCvTIjqiikeBh2cq+o9yy7R
WdSTP/ar0rwJfNkIynqH++KjAUNcqqiilLbuO5p/2HBa9u7TTDS8GEzRd7+TVjMLJumGAvO/bbOs
e8O9xhWgPJSRS6GmQB6NRMe9ihjBTHeR2gVT29TQtXX7APCE2jltUwBgIL/KfZFSIf5SenOrmuNH
LmCVZddYcBgjZ9k2hc4IQBWAAMFjLVsdievn67Uy9M7mCs5SziMSu6C8JuA9T44ltU4Z0QsjxQFN
smiYthWnvFWEkvJ9FuNKwOKXGQMPJ3omyZb1GkUQzh7Qw83hacATk260Sk3GD9phuwIGCfSzgoJ5
Ig5P7WvlPSHeXnxgM2usFOyb+CA3F5u9EOdm/VwO6A6Enl+fLRJbZmTWyH/XREYzGWY2lJw6ieu6
4xE3ttvRDhtU73zSzvusQW9+Yb6eQekqzDP2yKU/gT0EEUURTmM/y5u/v8fhcg3gGE/dJVVpBS1/
DwQg/IsB2MGnMQLCdmUhS4n71hfcvo6eq1aELD3iMhxlA5MfitHO8W7eEifWC//JUQojtxuYAb9K
EfWAx3CF9vjIcolP0SGPxtksQYMeYxN7ujXy/CZuizi8T3MmRcscx+QMe4Mg4PQ74LKBuIej3TJo
N6OrDngEODp70bVXhthaX4BNm6PzvOyk1MqZ+k8DfpFZCMYP2P8Jkk28qRRZLPd5GwRExttquDoz
U21s7Khp6/T/fuFZXN3svSy+5ofOwiNouAXfceeR6SuSW9a9nsVjEf7UJ0kMJFYy1V8OnH+GwIYp
nL4vgQK8F4Cq1d3E3KhuhgqHaM8Y5Sl0GbAppsNM2br4UjVPBmPCNvy9DQWllJcOTi+fSe59E78R
xS03UmvwsWKNdqTDpiJ1zKhDMrFO6SaPmWpl2S8LIqW46krMAjJINi3UyK0vxxOuPE8ICT/rWKUN
0bdXxtHD9Ys6z7ix1HmkEKAyPxbjRxY5HunVZnMu3MYC2gIb/N1j47Z7qlwOnGjQ9i9IZq7EqDQS
iZhS/vKpP+97qT6V+Yzhna077KXGyyvqrXbRSvMknQFJM5IonhkjBmtWZ6wD7FCnOf5imKL3CK3z
aD1NHiVAgYoG9f0j8gy7O9x52wSv31mOGMKPNfI8JfTuHwNZ8+B3WdtxGi8mMXqtcQtUUFUzKYEN
TOetMoQFWI0AuyG/jvXJomb/fDxMjyDmxe7Pr0VxE6TA2vaumqKcii5du2boS5hi+9z1/4gSycWz
DjOf3u2NdT2KTblEJzVHPBcSg6dm6sof7l4SMhxERrtUWs3Mt3xO4hrmrSkdOOniDMKCHMl+n8oS
hOI9jeN8MEaD2ajESjp3Fioh8gWXBANuYSqL1xmEYzCiUshfKKQEcuQYnmangBCals5+EHNjQIRQ
CWDiocglrl1Cwme+3g+v0nQObLGmU3P/YYzAQ/Wux+omU0+y/ojHq+zJYAAQxdDJh2OvTrWbmwTZ
vjrGcFop+x7VOGHMfoZqSW9iUMYFpOXaoqaNDvMU7dNxso0C1XAJVRq0d+SjyoD+vJnnGDdTT7//
k/GlL+5SRQqqp0M8Ps+F59gW8mj7iaumRfHNTbM0y5TvFQBL/YGVpLEidzFC9q8QLIEgBuZxefrE
h1EQXcxwCRTqriIuDpRlWz0+ju+WQpqNWBe+q/q9x4Zn9omljTt81ReEShbzTyOYQoRR7MY8P4P0
4maJrJngAQrhoehVh2Fr2U+m2aH6oi2Pl9m0EZyXeEkxFTgcm7AOQXjdadbf+y67GyhqgIkLApAs
qCg+MORX6Lff2dodYZmy3AdAC1UhQRjdHnAyQuon2b0nzLVGClYVB/7gdwrw5Sgxw6sn5oqn/yKB
nx8nZchgtlqgUt9xvEgA7h7hpSZCKec1jFcPg9mjeaDipRLWM9iaz+c+DjyOZFgp5xH6bvtos6OS
xKJIaDntyL0tlDPoZRZmz295Fx0jUVsnmPqjk9Dyh34CwohkAsC+4CIqVA6UQA52fS9saDAY0mL1
2u47YWkb0ONh0eCoGJvaJTuEPwvm/3dCHhrcyX/DxN8FUW3CLwidFjST/MrMWrQOGWtP47lI2RmK
thzklNveEkeKIp077rm6x/gxQu4pzvEl8nvX/hU0ljDkVrqP1exkQGwh3skUUsUJZIaG+eKm56TP
72oSV1RuhRpEn25T3eZKnDXL/A+KC38HQJ4FDasfN4RK45LxtcL1nqfInzekKZXe8bF6RN7TqSDI
wiGjUtj0r776zUijKErEOiLTLmrbRJB7rvP/3ocLcmwClljbX280mk91Eu7yByIeSn0sPU2QZooF
EssryCx3SP1Zn//0AwjfBEO9vGsDhgccGGgbUH0nFr6PCC4JWw4t2eS2A/0jAjpK3Gt+2EWIEwdy
FxjaqmoHq0Jd+SFpwfHj2sJHzBYpoTUlhdXdw/F5tmt0ijlSwhO7Y+OI++vzn65J6+EpowJvmXRZ
soET3VSKvDxC6fKNntAJ8BxeVh0+LviUK0qjvfINhNVPAP6FT6NUNcscIW8HL4LOf96ta1DlbKXH
MhtgLNEdKPgl8Fp3p4ZDnmB61/vbNCU6jtakMk3mb75tzMw2cPfAO3BENBVtBh8bAQ4DfwrxMBwA
/nRGwtyoLL/sKBtuehlPj2Hikep605saRq8tftMcRyNFKRvfGJ215dVws7l6udLyejoaZon0/r2r
KY9NkLnyAQYPuyD55VbZPQrcnf7m7yqZNyB84+hUDGke6AQ9K5w1odeH0TRoQ3+ZeqYi/NRaHkxa
F7QLZqDgJNPtNgs+b8XVm97S9g9TtUj4ONMSdSHoxA7m6uAnLtHxn9YcD9js6DhFUobi9UTWuOaQ
o9tXl0AnLTH/wmT0fQfxIaYRg0mpBcmhj/v+WH84nraNDSAFqhN7af9I2VDggSit331IA7kXxNRE
zVBPx4LZt3VoDv4QcnL91IfjhSfavLTBpud3GbJjuHWPvr0WSwV/U4WXhsxBIk8+hqcehwD8UlWj
YiZMVU3Afph9uAMK0EAqVAVZiC9uRlT4DIgexbL3w6eOcfQLvHGP0gqBfy4JIIrs1LfuRlnZa8W+
8la2NTnIGvqwj111opgRUhT6g9V799hcB11qi/su/pZSbCQFHLXlEkU+eF35hCzYWKr9mfiqG7Uq
t7aEqc/GnEV//xlAbWvA1sMxQPsyvFo+eQ5xckKcCOXCYHwi1Lu84u6uAM/3wGFF/seVgVrZnmgd
c2h1lVTTJKtzYH7WMq9mtEqz3BuWEG0RsBSxRVkMni/q9L3c9zqBgBA48O3OHU8pyuk2w8Z2axS4
Fw6qBvTuReApjGkzuBOeLkL7LstdRXWG6fBRU2w86ylR1RFZAHUknBvqjT+NpTNOeWfeyiQC/hr3
WygrVemwOHMsdGxy1j6DYKVtJ06JpBVv1ODY6KhZf/7AOen814KN7N2EAURpySgd3CAivOPyGsRO
UwAXr36SBzNWYXRd2RNJxd00wwbxLOpJBr6plaeaTxF3/5WjZkQz7nUXf7L86idQ6A61pJs8NHBa
tYo8DrHml6dP6vPeXUeMUpWj1C8uom/L6owK6cKKV7+YmlC/4I3/u1UocQLNJFzZ4zHRCXm8V01I
/gVaZNF7p0PI0r0SxfDC/adMZzny37wcynOhRAdezwa/I4r5zUVoA+VgJ+ERKlv/poZJhW6G/zxH
ufuxnDOVyI7rmpvjrXEBE8cIeQyi/aaLyUVI7QqOXYz3CyJeb7pMg8RLTo96XSRvuFhfXDzuqoBt
ZBSYCyLXsTj8c8oXxHDbPd5tP0lfcqOEC0Qw/ca12wexuKOd0DnBpAuLvWjEJlE6M2HnKRvD21fO
CtfvdcwV02ud2ZucppXI0tvMpjlUJzfw3rYCS+bDhu8khUj1kc66CBJkmKIWB0jqBV+T9kUzB9p8
vwewPg81BiXztVX13UHWY8smfX5jXdtu9lY0TUXXlTvTRYdkC9kLu4eWyzyGhZC2f6eWiZErONqi
2nfgJvpUxYVoxpcpj5a+d0mrpt4xE4n1NmbcPZEcNlCJnvvzn/pKTWjbxSvtHkw4y4/xQVLXN66J
lVErCTHdQwGK8IafGDBsd3gay0gaOWOn5AQFn9F22GiOJaOSlNbBxvAQoxJB1EUfHT6CDZXoWGvf
o7WClpa6MseHldjTQJdBaAvuIw3K0N8qW8eBIcy4miXqOJxYL/fs32m2/Rv2PdjdGf0fE5tDWZFA
9df7ChF8A65ETlfqJGt0/k6BXCUWgXETMcds3t7kK/PxLQu9gsZJkrU2zF32WajbkqJVrTz365yz
YuR/kNlhXouAhF26dhajBkgnYJ812MvigHkLLuw6HaPuajpgLBgHlYZpKlEcsqU7GDsvMd+EC/fB
r4BTYJqYeU2VZTLqLBrmTOyV0cuCieMr6RHKH/IrcYiGgyDEXkK/LlXO6+8GylWoNMUI7VkP349F
g/Hv+H9vDaH0hqiBHsj3zaSFYb49VKIB4nbeKfZEOa3Z4sHbY0J1F9yDrJyM+g4IdT9UVJ5SuEaY
KRPw+SovrGqCBgjF2I3Dh/O7BRK7GMMMlKfKnNThNqskoWEzQxQELpz5sK+1U4QQl+I7GTXz4GWw
sDg6dbJNpdQMTXAnl0SF5o/ci1HDiIWXfAFltM7Re+38B69lbG5IyboJ/dBVVITc7+z+g6svEows
dyaZknwTbudDdqOsm3ZhITkN7WFFHFaQeIpP3lxS7CBh+7Skrz9ZTeKdI4lxyVfeEYQl5RtkUtHE
heYbU/6r9uAfbWStJ5cdZpVgh5qUXNs5/k90T5nMRSWNnHLokJqkFrU0xVmQ9q+UE6WOyPwX+1gM
J2f64szqCav5YOF14Hk3ffPQZvAUY5R5YHwS6MOttPc8JwWvA6cIubIy3wBwEdQ4TB1I8QBqaGme
eKiGiZnYgrFrtp+QDkUirsSZjJiqOqZgb4kbtzUgM3EIcR2hSsZMcpGSmlxYbTR0jB6KtYKgqjJM
FnUK8+pid414PfRPgQfv2S9OJghVUlqLARorSnABjHVCy7xJ05dCeJBZ+qT0K0RBoBlThR9e2xlT
tZZGhj9rMeDb7LWMVtHzvx9XGIyF0aUVfRuIrHSkEwK2McB+pVbrN/IorXhbiDJq87ku22erIrDb
c3UA9QhL4pg4e0Ql68SEabY1SKC79uu+XsIbEvlTfkhVE3QU1MpJ/3uysBh+oO6sMD2MxT0Q3E17
7mOiR6nMyZkCi7EupCtNY4qMMyMGz0XhS/bQgYBrSBeeoeNYbv6JwtDossoHLg0GaP1vBFo9xdpx
pr6e/SBG1EYo7Np9v+Ca65VeB2sw6nnn8S5Spe1sOaNnUCxkJrUQtD2wShAGSV7aG9ElZLTiKwvN
/t9etffL4Ol6IMgNtxsl/HJMo5H6cWquB6xAEFvkv/9sgPFU/cElB5t9Zk1lWNuI5iKB4eehyMir
iKXeCgeptxeOAQMwzlSxR0p0AhQFT85bMQ9bjWfFMOPXtwJvLW63+vt8eCwX61umyFJguYhbIYj7
D5GozG/VEUHjdkz2e8nhBc2Q3Ugokj4T0coEaJ090H8V3C2beXfMJTj8wLomj7OdAIFYhKvnkdFL
LLw0zQo8PltMZBALLYmeqWuaAH/NXxcYCmRUl1p9KokkE5+mgoYAfzckjPlv87L1tqzca65JY2+3
QpVS4Lc8wwvtQZu5F/d0SW/Enhv5pYXCvDqNtxfpKOmKBH5CreoONU6Qu12p1iCrK2QPxKeQoCME
PBIxjq50ihNRsMJCXVXszqggRP2+3SdHVdoC2gzaTV1GapDM28k5/ha0niS9xtPC3YWy710n4bU9
L1TaQS3thFBok0SM8kKYzHR1mQObRD6wxowWthl0NnJTtSx3Wwq2dkk5UL4h+xLZ+vdUMBhu5F6i
OgJ2N2kOWuJy8MyIGYA3cmxx9jdqTvNx4thUA8ZbZOXVLWtKHHwUsk45O53IdlJewUey2impqkEA
pDNokkw+EsQkoQXx3fSPGcc0fwIQ1AML2ZF1HTulRozHKaFGQb5xDMtbEI7XV9+Ui/5pUrUplBMc
rSFKYHbd3Vel41V633/vACAFv3g+/xY67xe5l+UWEtnSW6od62+8tv3V8h63QMPeqAMMfbXq8rmM
6RkWpYiJVqAhQzR+Vl9oHgL5L8DGLqqWH9BDUKK84PV1wMYzmffofeMBuQhc/bLpavwHrUoI9zDe
2C+cMPrAYsZen0eus1kRSPlgb/8w9F6CnZ06s+6WWS/2Y2TrshZDQKdOEQQuvsUtMr3lCv10FVYG
S2/keLeHD/DvxmkIqVg+Bnzc33Ssc4tCkh++Tj6WGQB3iJL5PfoJ3XB18wjqiUk6eDdNf8APZOCL
QkzH7/H/iZ8yjUj6vRInQ/fxwuzBcbpbKo4qR8Kp5F41QyE5VVzgp+02pwQ2OjSpXTynCebtqcl+
f+k9frr1jqcA4EPIzKeW2Xf0XlvbHwPmhwxwdlBr2lhIb+XGWzGYEBoge0Cmq8UXSJFFzisFGanL
MANVSbhFAnvdRx+YdnnJq56yQ9FC4QdA1jiOlC51gjDIpBJYbT3WFvPXkl+C3eOo8GtiaDD5Js8G
+MiL2HzKygrhfQCtUn/um+h4kguNfurx77CgCTm51Ff8wFCTSbJiX2C1jQCscmHklB7rPpHk2e+5
mvQ6sz90uX5L9NVnFALxozZlmBz05eLFSMVqoWgzGgOBMe8s2gphZnmxZWqw9g0wXK2bYspkcGi8
ZR8vQc2b7xhm/oknAUqoA3u5igczByK7fJEjLyQiuHeBwVxH87GFclaVuN7TdQyqBr4b0+w6Lr7d
ZkNOwQrCpVhSt3aJFhPU/E6/384mvYp15UjPy/BYUWAEXVFjJ7m6acQk4lkfwF96A5IrHfggJ9uC
PqOWbzc/FOKPBTCaA9/hUNdH1hZ5L31wHb3/7VE50gSSZCWSOuFa3PGl/ITQCZWjt5pNx7Xmfu+W
KeIzWaR7S6TeNMRra+QPhNLPhT1e19wl13c/7++wT3vOG4cYne3j+lp6CZlhJUAATweIMFdd/Gza
U2mKcuTDyipkDYHYfuylOjSvA4ILsVyJmxEJR6hW6NOle4OS9APV2Evd0o4mVQOBYfyFH0Y424HZ
l+qhWKSCqtcnLPWRikqXa0zJYKHhsTmhZ2OUb94nKCVvvGYmwIWo/6Nzh5wafWTvkWDKINDvMsZK
AyiHuiZXnchY4w9ot5PcexWzBJeW7kl/MSqz6gDUn3dcJAMCyh9k6Ai3dnXkyUIfvZL4W6ZDc6r0
JpKr85LFZO6Cf0fwXgVU9z7XvVFYQSSr77J22XPBQuToQOFu86MOs6+Jsu4tk7B7BxgOP6uZt9l3
pEdzGBpmD9DtrL1fOtOFtKD+QWMRgy94R3pE39BvY8TmOkvsgsqos91NdeQBfYhEp38Vb/yrRTJC
e2XFd7vTXFKR7CV2HfEoDgviQhmEi0F5MdHXl1rxUovBw2Qx2K0ME2uy3smXUKOt5WjXEpwrATme
PSebrWSgVW6GpkTGqH+fqZfU3egVLZMan6ILny7pqiBoofUyXS6eq+HtnmKdWNDKrfuZwXXkNDiN
CzOGsbgwe9W9us54rTwyp/qfjDKm0qPdEj+PQg0sdTP9it8q3dJore1PB/xI/QrgypE6i9+hLqf/
Fabe2J3ehMSImr4kIBBuuojzJSIhOrUF4sY7qvLbxWetgWgWWspqlYs28HIxtWatN+IHDTl8yfRe
T8Aco35TwVk9C5YchdC83I+DkUX9kl77r62wUDx5LID+tJhcOCnxhuBFykxWniEiqDJiLpDHUCHT
v3h8dhUmIJyQgAJixrRux0EF1/7DQBfP1k4s2DJwFqk9w6DLCVCy3BTJp/+9QFkd5mDpKSy6rXxn
8tVXEdqfyRo7QyUFZxcS4NSGi6mD8W424MB+oJ1oN0s4diTYtCQhOXH8HFOYJhIeAAiDDSFg9XJL
oU8sjCHZxRG5m2FVs31B1MhR0fR+U5A7kDcmETmhM9TQTexVuJDKLNm+aTReYNpCFM1xA8Sujnpr
I1Y3P8CzgyifNdJgHeuCmlvzUCe0f/aIwuINKKNUA6CoLc9TuNggySKqzK7Oxk1ofzHqdDoG5fnK
PT8XPFi/adN9ckGpIOjpDD2W5nEzhRTzT4fBgdzHV+VLNpzWjkjQpnbybK0xFxtRjEWoXDJhBQMc
gJIIsJVhbnQkebhFFufh9VLgeMGDHJIJrOprZqls02X+OIcwxE7dXNH5zVvZKksyTcNkaA9Jmtqn
TWvTH1CA0SFQzZzxGOhh3YE8Fj0mxXc/uTUbvuhtvRr8VcLEUFu7hTQ+K/Y+FVVOOhnMJtftlkFc
XyweSh9akklXzszNxTyOpiYvFgBCeaQ33gJVt6IdKK3sVtmteOWfngE5nqr0qo+AiItmTQOcyAe2
XZsolOKmAfOAb6Qpj3whMkavXcRHvwx9d9tY98GK6xzYhfiKejUysJGpKwBy10cW0L2DfjHs3qri
x7z1ldnmOLhCtRh4FyqXW7BF3b2PdWVkGp81SXQvKqyBSD2Pjj4eAOXqT0kUNz8t/effmcYeanXC
F4r/71BzaRhjJgabVGW6I6nf8TRm+QbNSgoexf8aXEpj5rEPEl/cYs8Ay7prvH59Y8ks/Q9vBUEg
iuyjonJhI5TMk4TgUdQ4G9RztfW5cRowOP9nm4BpxOouYNsQEIjZ80CryD1Wt1dkI1PuzF0kF37y
LIYKa/LZ/hsF8SGgm/QkRwXY4ltxAIyVoSxDaGfPvguqk4CUKRvlOoOlpnWtQUa2lCMr3MwtRdw8
T8Zf7TycqGBz5HrNdnTAjlb7PjqTmTCvdm3LUSMY4HuP4CzZWcMCM5MVa+5tHBN/i6+8SJoYl01b
Z0zSuwxSHODAySWs5E3IUjn96hfc1Z9nCfWDdHUcJXUN0jaNhRz82f4yYS7Z7Ai0cQDFJwwn+K2w
z12sA1NCwEgn9XAOJWcNsVKeNuofdZ6fgDmSAU83eWv+/07zwGpj0oFtkGqw3c971RZtiaH/iHt9
f+CDYIp+/YKuE0sZse2zKVrk5jpM9es4FkfiaHR8/zABAqXSHxfaVL3aNCFXyPgdT/hcXzF3yb1h
uL3MX59253Cooi4FXADjFCIGUtcICfRi4cAJoXMraja6QZkN2UdO6Fy4cXAS15oFMIPdLMcYv2ap
i5DyrI6tEBhDVkJukhjv7qI2oENJUCVEq6wlvIGwrXHGEeqC2/oESs7Xf2zyCHWdlm9u0cbogJLF
cHg3gnq2EP8O0AZ2w3LiF0NdqPu4Lm570Pp6Sril3WWkYlakCnZGD87XokTU6MzNytqoFz88X3uA
R7wyguSmFM907CB53TTNJJ9ZL4N0tpdAAIre5ltXdBk8f4nFhcyZt1RnUs5z9StQ34yebAU4r8x0
8iIxcjhb15ta8EZf2l2uhf8qcAo5dLLpLzWhAkSA3Xp6Wvj7LdHeXc5sUYOgWCz7IMdLNGZQwaIe
JSViKnpLaFe0UeO2teKcKxPPafvPULJyla7PWaj+bP9eBqUh8gSw3RTJd3hNEbwI54bcqrDE4PC6
Y46a5zp0KXXk6ZXGFY2VdpnIG2IKuhsUjEWE/uHUtIY1tKpWuLYnw+UsXpKeAkpexUp9x7QmT6yj
X7PF4w1xY07oXo3Gi/rXd4VqHnjZb+UHv+OjPxPccagXyZVmXtXFzzBIEG2ugP8ylyaM926UT1ju
7WvK454z
`protect end_protected

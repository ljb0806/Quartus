-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LE9bjWwidRX3b1R+q9V6VwSK1JaAUch4Nd8UALxHOzhQgZYEpxNzvxO1LWZtUses2yErFUpQdQHh
mMYWKzzEQVXeEdrTPHMLfYg2RKXCAcv6uHPoFrbX9PJsOorh5o+X8VCBchn1dwK9zYyNeBmzxiLP
sIctHck/f7mKK5lfSmhpvJhoTCOL6zAnTlu6Sk1k99JWryISvmZMEt0AawvPYcpqlfkMOYofoA2o
uDD8o/+dQt42vBLjIYhlRphF03Yx4/w1zOQ9o3yORn1+NbsdSteJqocsdT/qqr5BOP/zVmw5G11t
7EZBPWBUHFM9AYh8Xp5+C+GjaaxuE9jZ4D9WgQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 102384)
`protect data_block
7SXugP66+U3PBNbvnSr141a4IVU6b63WmYeyBk19TZp0mMYpzvrLNpSfU6n6HMuLykbvifwPXzPc
UAxIZy/wxX9ALm/OXai+kiWJhLmJZFf7kRYnEvXUjQyH5+ZlmtoQ/JeCZro1yAnvvJdaUAQmN7e6
CZ/0geSUSxqfSAP06tgL8d5wjd6u246KJaeD49RST4a0rQPIcF767BlKL9QDB6Z5LFtLDdChuKoZ
rqwcFzM1aNZTe16Vtwb+/12cJb9SMbYhZyiYxffWt7Qvvs7B8G7rm5ckkcwqQHCb1tiShu+ykdUJ
Qn6BOIrct4oWA5nbB0LQx7QpcZ7u6tRs4d/iE/Uixkb5zSGGJFUEjtRMsCZSHVpOq2HXZ17PI+/+
hmpnDXLB+H8OW4qpsf3HA/tfXvZSbc3PCpu+6rA8O7NZTu24/SS95BwfuLaK0IrbKv43c1K2EbKz
jU4OObOIVj0OIspWoQVTLWttQp4E6VaB07SXWsxXQeAQMaLN7Az3mjrdj754he45Xs8XB8Wufjht
iurS7BWMboX3B3bwG7oqgDhV1QF4m26TmSkY1amCJnTd9pdivs+BQZ0fwiBWy5LigPOXJx4rMa52
FDrbHbzrqrpgtn9/XZ4ofca7/rehpcjTUcQgOMbbFYKqZZdPKCxmYoooc6nc4PB5o8sP3ln37WW2
cvzzOQk7Gvyp8+eonKwh0bk4HdceEyJ1pH0ifFN2/sKjwE6ad7CzxAsUS1lY/XJhdrIUciyoASb9
zgopc9kz5NSzKjwTpFYo1/rJQB+64hW3RGg7Bi4JEeQCX/rFYghThvU7hqOcI3/7Jk+XepOz4lI3
utzEvBoTr2LMB8dnoelQ/A9pFgMSLcafzuhuVKTvwex8qHytVCka/DK+DEcFr/0nFLqfqXKIGfmZ
XNFYHUFJMmXWNou8JjbAqlPHKlwWO4CTb0q6DYdpDpeIDEgObA/lI7/kYg+cDXp+lufPkOTBnEwA
FN289xmsYCmo7lp+Gp/wx85Uef74lRTIl87VgIOYb5NKiBnMPMJ0K5pbWTlNRqlNrJNkFXyosv1O
wy5a56nNI/VOjQLBLP5v3ACKJjrk//sGhva1qAf2VN9/4o4fGcO0AkpbRLhC5LOxCweUjbMCgMiO
2hjiWfSaYxiEh2/XnlIYslUyN5TRnJ4fejNgBqEhEsVomOljlq14aU5ECQD2E2mOKB1XKcaubdap
5y7HQXSaOIKGRZizIsgsqd7VpXGFoQfmVz9pekq25t88kbBq7rDR28xghS8cxJwiTrFnkDRHXWQE
EWp/bPVymQJzzu+Phm06cOvF46KOXLr3hUnykqWGEKzJNjvw7+/SQaUVuY0qs33HR9Z3e4EPT4fR
+diJDw2TxE+1GM2dFBaBkLzr8WJ7ZNrT30jBCB9NVBVGJsKDhPMVDl203PzOxQf7UAdJ/1j/YxHO
av9IGL/YRinD52iTPEcWwhlB+OAhLr1qvb+51eqxyehHbmuDiI9Sx37t8ZQsZS5Bj9MUapS4R4Ft
poGEoBZfE5dRy1rO9biaFQ6hjCbe5cLZYthuvq102JqvZApdEN47mUlPCOs7EOZc/98BI6+mRfB0
zEsInYYU8eSpMXBc9bv6WmKQ7rUjQ1daMKzdcD3czajEv7LiCFesuXk0MR201GKmzC9PyxHHM/QB
3nDTqxbQNUvVOEaNBGd6pdaIh+dKQP3tLimAoQraqqMxNKMBZ2zaDUOyVe+L6AGMnO4sH//raMRC
naZLuVo6lFmK05nF+VGDmUR9ZrS87DmqEx+oaVg3DI/j7M6VnEjrXqCryu2YzcCg0F/x1s88Vh/N
lR3FGtvrpzd3dPG/XJ/nmunFjLSNmDo4S4ANbvzwqdafPaEi2vfoUTBnX1R7LILjFRQ9oMy73qfk
01YfWXIdA+h3yaOyprrNcZkpS48OPr5OS5YfjTyeOrZ07Od4AshPctqw8QvP4YnLcVOw6owvRS0G
EIftXwvunHGo1bU2Ug6lyudqGfpTatdD6UBecqXPX6soS1kov6jG2lsLnh1mr5XnxXNT3US6+DLi
l8UD/TmmhxSkgTrYMSXpFb8ShMq1WJzVV9ViINBcvL6bDv8QHfAatpLgLDzWDMpPW/OYq18Utr52
2hOpmVYM5dDzf9uYyfQP8Z8oE1W1g+6PTRT8w2s3Bvnp8VT9r8Hd0bIgbtPuRDODi8oPb+dho0vE
W5L+tqfFfO0OgKYPnD2SizTFUELNsbNkckPzawvdgstgMauc3UZXoH05CU0Eo2lSOfT+40XovNvf
wHMWwk1GPR8Z54Q7nbKZqqbPcsMKg66+zaBz2TbRpRL0OV6MeA8Zym8WQutERRxNr3DQTle5erXF
BhB2zWkeZO0oltsoNroefAoLRW+Y0wojJaYeZKcgT+7zGXxwKCEv+0a78BlcDa5C5iYvFZdUO6P1
AhkEpUxgKBehancXbmZAy5Oo8ZB8RZJd7N8aApd6mXRyzakaClQEKP7rs85Lx7MA4yo6+Eg3sESq
Z/Ryof2I+PsWHlAyV/otXc/Xxi+ERANaweULxuWOfPTaJsjTNs10eZcKoMVHS8CS+Vp0IT3nPpbr
Q43DrseYe47oDR5DYINZ3zjl8V0jcXo0/IP9jt4LWjZWU2UKQQng+4gyiNU3u2YNFRtNCn3WFGsy
cjhMFl+TbF/hm1H7HbwUW+5fCqPGPxXB6qq0Ik/nLt9uRgs2DcJcrprFqVC2rQdXdtDpsul75jkY
55WRRNbhBbFVkAkq/HAADFwOkHKDCTeET0F7NLR9Ul/zsnPYuT7oWmPat28kiB5Yek9fxZX1NB1f
31K/lKO+t1Qwe1Im8S0nxmxqSp2AmIG9D/WmvlHuBJavpYdVMaq9IZJCJL+JZG4l01976ktwuxLV
Wgd+BnEKQzE5PEuA2viKiR2oNeBRQ3iGUWAwUBq14QiofOAG5fAtkz1w51LH4V0wosfsegnY8kkg
ydDs3bL0KGNBRrxN54r8L+U8fxjOeOa1PMfY/Y/Lj4U3xg0xWQeko0ZpRG17PKScWsUEflRyNW8g
id/y2qHK4KqdyCvx31jCeVkgWmyAJGIB3UtD/wPx5tNb9ilAu3PFuaO/RBwo/ALtEXyLEm7CPsgl
F6KC/GaXg2pR94227f/T8txvoJQ3OlSPIhipUICoJoLcL9/eC1qu/icI/00rhYl76EN5dZSnD64V
e7tna7B11SZYoE6v9KQCKzyvcRJz4A5y+pKiSHlkRqz3F5gavTWe85pG/RXAE7tN/qG5o62j9Gmz
5UcYqHJJsFAHeNoe5MNNsQ4BmaMwNuzwfPYfz4kZU+dnup/fv5BR4RLxVWO61yxagN6pC1cA5lmg
+9avuQncV75Ef3WeKJEuojDYpH3n/v3Rw/WImhX7zYz653ZoOZhqgoiBkO/6IZYrpxzA5B4axzj8
by1CqEiXk+3FlfzCN4s9FMyaQBIw0Nhhqd+i6P8t76QGDNVeig/nXETCx5qKzEFJAg9av5wuxH5B
e8a5DFMGdW4rY6nla96FrJD2rG4s6CBh3cuIh51U/26tiSJ5dLh1JgIsIHOnDcHx8bnbNOFk1kM+
/CIolCt2zvhvf6rOhVfOcvMz8QPLw/G1fvERk59B/jPfZGJWbUlA4oKJNbbyYZ/A/WkDOHBdwy9K
/0cKgcufXSHl+2BRbLpJQy9z05cgrkqVKSnJtQe9POnuVuo4mNDfj89O3gcfaKl6FYQWJICHYjWN
seqNen7N+bd3TX6fEChZon5nEMPPbu4qpi1soa9jno4bLeZHpq/jm60V3ImFwPVTvG+JT4QHasm/
jr3qrHTdscon4lI/zu/MHUanFg4rxWKaccAku834R8ku/0RWqE/76QPrn9iZt0VH97FJ41vg8pMb
HAIe1GwWyUuIOMZzFaym9yHblppeMDtvKxIVin9m3YEimz8dLmnWqJbXYIrxUktchOPs6Ti+uCH6
gISMnIO++SrllLhIvVI91gbPURyvusfSclKJLcB0Afa6ZMgPFzD8OQdQ6WboP826YhB3bU+heINS
0AxYCL4eVJXoJMRVrpU74M0jcbx8ss2apek7BgitPO7YSMQpjlZWVIiXx9LZ2sd9nlqF5LssrL5v
FYvkElP6rzho9Du5SgExXl3LIXL9CX9Iv+CTpR9I5uIbA6i5U/H4Nnw5FJjtmv6oS7ZOnWfuqS46
ln4byU4cxB28813QSRXRii6E6Mtq4742mfUeMYk2bN8PPM6WnjdAZuun4EeQVTQcJ1u/+VxTlxU0
DGeTjiGvs3dK4QVQKlPCZMwiklFT6typ80AJ3D48ioTrEJ5tIERKa8RzhbVVySrib0g95DbWOP6G
h28kWDeZBnXMf/AOEH1/AO5W6tSD/F0nqAcJmhZHQXOyDSWudmyfgoRmq5VsMo4SmrPbq1okeTTX
8/IqeM2UOScM8DsUPc6XRHV2pjqFfnFVbIRk5IqSegDJvn+GmGunHVSAQNHrWI7ipW1BPtFgti/2
pQcl6a4oUdQCjyZNtjXG0x1Z/GMEA7ddtH6FnORLHGiT4JqQug05j6hN6OhBYQNcVwlFSaLkpTsA
U6NDUqIirGij/B2mx4h+oY7JiGX8YHsJxVIInXnM7SkckK3WPFkwhmFmW1sBey2gMCBSoLAMZgL+
+nUlc5z0pgLECt/fKr1qwU99CPvRXJJAldskpa33e99mh4edNb55JFUALDNWH2QECFSu1nqieIyY
K6TzmgGqhy5+kjBBTLit+goWHQyVaiT3hxHgrX4UwB2tXqo3Fkz2dzT8Z2hFr25DG8NrXkWkh/X8
JxwhWgAYqaEYtxBY5e0yKWZUn9rMG5nhIXtGZ9ZCfYbE/FR0JAJABY0Nwaf5hMgt8YPg2xwiAb1G
khsMZ2cUIAQbBg7wOmKV0cQM+K/ThHrvZkAum170MWRjJGwZA639uIXC2Cvy5WVILVad+vV6f27X
+PtMmk2uMt+CpIEDfbMw71e5DXcOAeFVOfaZCuhsMWSUN8SDZjzXNYA8l92ojrrEGvBqzTigafPQ
YxsMz5D1yUFis3F21hbL/Vzb3T9HGgPS5RMEOmwRX1MKRQM1KkwerOMVUhRB/C9FJTTNneCklQrL
2OwwZ4J/PxVWUFH6oufqY0phe66wLh6mHebVIi1qgkWuZW19q2EcHrstgWI25kG2l+BrwFKj9yJ7
kSizLLU5kdw3S1dL+Kvn8yOouvF7qhFm/rqfZmvFEUhaT2Vhm8g0eEuUuFVJEppoabFosfYlnUh9
s1GGGVBGbRduxI9dOKnH67YHI0MfyYJ3ImdtXMsyR9D2HeclTd6ae3WhEgSGxZwJn0mXUBLYK1kA
DiGaBcroLkCW1s+l+CK2uUe4nb4mtlHTZ9bpYysLbP6lmFexZEvZtO3Pnie85kdzGwWdFSy3PoTS
oeeT+5O6hVef+1u9JgL4pS1YpddqifenIfV2XwJJ4fjry25tsOc5leLFz3QgEQb/cZNvvNnK1VcS
ygi7JiJDjUEGvY/Ua6Ub5KAWelCuOuDAy/TB3SI3qL58Mgya6uYP+grYdkSRlGFFrfW+aK6URqjo
kZxozexfqcu++4ZTmSt2GNGgER3PJTeEtkL+Qo55lCWCzNTiCm3To6IzOH+HR4ro+Vjlsv3T+Ev+
FHRvTkbqiZovxkNsaTZNlBnFPMEiU1PC5WLlnCVI6+Paprk++pVu69FBxQgSXmQB1UIyI378NUsw
hSsXXudjECX1MnJ3jltLlcQ2sqJm642o83Qj3badeHWml4mKq+TXGcc9OydoTs1FaAGuU8rpN3XB
sNskVS/UfusT/CBfkspLnXQ05WAa0C9ThE0P1nuYSi/1gvLZc2JrRnorhJjPYBQWCdLOF0lMsTrB
kp234Uoo+NJ0MawWPwScnWvT+9Efsnad1fGUzXVNVJx17SR4gxvIanOBEJ8okDlTXz+Jy8qmLOOp
qecJwOyGpZJ78Xe6vur+6bFxKYCoVBQUWtKI3lu41toQW6S8ILDbnoWCTM9kxXvcFLGoTJBFg2g7
s5q0onlw8d2ca/F5OcfxwHBqQBt0sJQQCR/eIRaZQwvW0dF4IM/SmywPCD3GyKD6UryCzizT96Iu
4JRtlfeoMhSWwjQiuRjToC2fpicoS6yibEeUWgMrNIDvx6TvhNBklNYrzd5xMrvSm5K/hLZdq3WT
vdtrohHdte7mAwHkpyJtE6KiBEa9149i9bdATpqx/CZa6rGK98XwpehtlAtQ2TLAHruzWSY4Aao7
KhPQ4RV5IV+nRk7OmFD5ftIBkCJ0c91lDic2BiWhiCFuYU+ngI5JPeqrJh9mW1cbMpg++kDVrDxD
4haKhVvQeSButpe20L4KCFhRw2fWOexMTGdo1p6L6qYXP6S3P51Aejc5GhnOaTmD9N+LAkpsoP8L
XfFsNDxLnBPsKbRoVUv8ix5HZvTnGQcXKe7mkzv1GeDxu9CloLU4XF2fq5CT296VwbiCAVx7khFK
gtoxD22D9HUZ6ZbiqQBQIHx6qxDetlzGGI050UwkkHIjENEw02i6z71Dv988r/OkEZRT7T4mrQN8
e9tu5V42J484/0mUmbcgliAo7x/b4T41C6RaDayfCR5EGnrU/q2/yN1pVpMho5g+z5vg3mplHcKQ
TPTmURsus/HDB4xxic9Xx7ETr8PkBlI6IpGixlxfNGibFqgH00fQK8lqUgR3Rm58yu8zddpNcNB0
p1IeUZ+9BxFxWqMkJDIOSIpdQZvg+AwdNEZRv6Geahm+iJLRYqT/v6XGh+D7YzhGJT6UbJQjI7Wg
sNVEKLwsEhbo+kLqtpCo+2VZMcILymWa0uA3QsoC5tAy9XsEg8/fr1UiwLb+qJJP4vl1DjvbgMe4
ZzJDpBLX/dZE8ug1jWlSgs2PiD5j2b3Ehh9LMV8iSpEPmUjaIDfTilRomKiTm2nLrcdH5H2alWTj
ThddYSYjdJQyNuA3RqNX8O6Xjc2/yQiqozVj1hKhZHLPFkmsEBMAAENd1cSZEWhc7d3201Nyduvr
gwukHlPqQb36SXWxAsWZSBa7uvdPX/xKBvTTUzZB8PRWnVcwh1GeXesRlmFF799jxD9dEk1PR0BL
UpMJmB4XJeLMhps+XepbFqz0HSXnnbfCKnvEu8vVh162ZDFvJlldz5FjdUVWMnh9H9WG4LKRF7FW
sDxKfISZYbaht4jUzgtw4o2vGD3goFgwR4bHGttbIGILUk71F+huIQyz65xDacyNMc33tznLS08L
W81pZOLqV4UVoAoAIcHtUBuN1SHzvQIjYSoyGCD/kZ/rGC2aGdQYP9Lji37s1sQdbPR6IyEM3A8G
yfgjqQEgaO7i2Q09Oe2asR8bguH0n+KH3ijzUgfwm9kOM3oz2HUmS5gSMlHg57KMSg3rptGostfq
aclzJxxn4723kx01Kd4vGW46GtqPItkp8ftuXRn1BSN9ymcdUZLaPUzr3C7W5u0Sm5LQyQz0YsLS
CKvb4GpV/opLok9CxsBCRWvwJwyy/d2ocVi0XEN5YN0XChiVErakZOHrBAJTNFiuhJzcnz/NGwqa
L1F8P2+yor3sW/MxKShKLJIBg2geWyEImqL3AkBfWybkdSqAuPmZFq+/29Nwb9w6Ynvg/geB/I7K
HVo6d5bC8NG+PcErWiM+gsjy+saDuAmJ5ztssEGAaohBhEkpGsu0tTriHkIBd+I57ZQe7CdGA4vd
j31RDBq+gmC2csrFqFgJkhrkyW3A+2+ajxNMYIYxkijILVWcUr8t7aa+29VCFWyC02KOadnRNDWY
s5zFv3JU1xOVwgUutKLl0lSVX0WF/4NJsTfLk9pjOjNZT3LoPhie3OzAgF99uCYt3Cq12KbEd1CN
263SSrHRimGEi8PCfaPGMotvtE+ChM5DwgmEfhNMFrFMxl5+Fm0ydXaz2wVAEy6olGcxgB8TD1oZ
fQ/nPIdY+fDra4/hEvWx9TkJonQ9epN++NKCfW3cqzmyl7l++tu8BlII8G7SKzgin4emtGCT3NCn
EHPdi8hB0tPiaNmfnE9RZxWX8bkukplyg61cJ/mFcEXR6PqVrUwZ9SiFOHPAonk6Fdk9E9H2ssuC
autWhT1J+KeE1lVrulCQwkLuV37XvHjyjbwxaJfBWWWDEy1WnRqRWz7NA5/eliUnVeXxSQrG3Ncu
onFZ7eY34luZkSvyDtXBFMiOb3n4wEeiJejnRgRsie79FIdX9uuPmD3ozTwuc5zIBsmF618SKvPR
dcpA//UdZiDD7+/xs0i+WbUax8KXzsHL+Wp0VzFTYLJVk/8r7QGfvVscqCBhcxUieXvBRaZWtVGk
Y53kxGaJAt21RHdrT3eegSjevTkmUJzx+u5wwad4SR6ZVpw2oVg9NuLr4ZqiGYH3tGphtaOfjsGM
iQLXJmSjWLjIB3z7sJFRgih3cNPesS2chFM77m1cbWIQO2zyrsqRu+Sfox0wQTR0lB4s9oerRMHN
ydkWDds2zm6Iwahbr3F1L27lOHnYVRmhnvEwrIq8HNftEuFqOsdopwYnM3EIIP5QYrsiUcb7MjAU
LECL+HSQGop0j5QaH1v2iKGfDtP6qyZoAyfp3wKOEdIm0U/GuR7cV35/7U3qm4BVnBnTnq3EccSp
bT6LvpVzRI3W3+qeHqdbCPMimrFCz4RFYEjdgJtDVrRw5DCNJfTE88c8q0qVKH6XxlMrFNdHVLwQ
7RegCjgYCa7DXX+LI3kZfp0++8Zw9/HvonArnNpzPAxG8XDb6L3oLE/1qaL+jVaN1ug77AxRgh09
5yUPnIVLkUaPoI28WwOS7jMFW675F337jlE5jjByN+92m6W5fsdywf/Olb7PqAloQzHEiXDQCeug
uU79HQyQXpWBvFc/KSP5XoK99jrFRObsl+mlpxIn1U6C/Gm4ng/z1QZkRUrz3+7GRTglINdCapfM
t9xH4cO8sYo5/tlOLEBaXgKLoz6V4TOxV3hiVo2mEuZrPFIHFk6YiaNns9+KnUY8OFw8i1HF2uAo
rbjqjONswg6TtQCCWb5ymPiMt3LPJbREKRH7mTPbkOO31HXhCzwI2xJORDHUXch+a1uTDW6H15Wq
zhFV8Wk8t0oaoZOImO0Sg0zY+M06/bfp43HDmll2TmxzeDLOYE7l4XBarNxJ3dz4PnpxCdmF3Nv6
LHFfPynHPuXQcwz+dZLc9H9SmpJNwaiGgA0Vig7JeWNE72l/fSM1g3K8TnHbEKXE3Y+zE0l0YLOO
g+aYbFYCT8gOFinj30fJ/TH2GdNUhNNsWy//9fDHVej5WFQYnaaNrdcNrwkxrQ9lFJZBF7k9nCLi
alAujItIeNFaVIjotidOvlh01KIyGyKXGADRBUb7vaDsurbAKgeCWGxFHp3+Ca+nYoiO43ApuiC3
JM9ocA5HmUka//91IpIB/7UJg+e6OMgYjzrux//u76BQFeQjzNfzALxpcS5dDUlkyS5k4DAva7nH
Oygn/WyCpR858HTzeomPlXQlUyHWWMB2qG4l63UPHslzP9TeK3xgMJHysUB9lDi4idaxv+cuVvhN
/9/lA1clz4teUvSau/hGsZtDBjCJADtCFkYECG0dtGRkyvyUkyZh1MCtgWCS9iGB+cBjxT4rjSs0
s85dgefR3/ed8Mx/b7hzcDFGOLod/jC8w6oSZihnjQgWSLfi3HoShOxTW/2oGwtRRmJQFsQ35icd
Bhkz/pOlo1Oa048aluB6pAnTqO/GkO5vMYQrprJ9PKSAf16KwvD5Ua4LO5kw7nQLpa4xmeA4nE7d
UGjA/hF8s1iGI0ea8r8Effvvh1u9uAPloYkR4LHw0fLuobyXig6mANeLIhIMt0eahSSTKVa6tYgL
vefqDRep5lHWIlAogIuID782caLSDr+5t9+lZ4sU/PeUQoZcB1/9W0OM1AIKtnD6xUZv2/orQz2n
G0x7P/L2RN6vA6pfj+if3yNOrHCYLW9eFBr6AuTnVvbIO3MX2o/OQGOTg+srzXN20ynFeTcBs+Jj
VIgbpEFHvP7ijAWI+utZxBV1cUiyMzU2W5DQLMsr6lYklpAaKs2Vxn7pxyDf6RL/l0Wh+V/txPir
PVD+TPYf4zeVyVD0f6Y/Zr9Ndg+NxS9OoXxF6RiNV/eB06JLI+pYgZh86/cnFXuj1aDORY4E1X/o
eDFc3egVfI1DLry6LJbsXHf3ZkJ7HXA1M13raKTtk4L/sOHJa5iVA4J5I++ThF/H6OZdq2oW/cVH
zEuNzwdAZ4QdvC3qUUwcwu58jIYtUXeYPKqmCXPzEZQcMA7miHkiXiLJn6na17fOovoYOf5wINgh
5nTagHVZJfyQbUgi3qcBINw1t3usMi/V5YKG2uoJSQZlVm91XsBndoXE/6cJKAU3sjcd8n3O5KdR
U2W/SeMfUE02pF++3yLhHzGNXaH2gErNmmjDBBXTkZPJIrV3WC+wJ58LKHGGec9s1oAzhyi28iZ5
+g+dgrx2CDM0OiLTkD0OqVtxe94NtpVTHwyNR8uq04oW5mgIzsaMkEIFBdQve9TA9i8sCrRmI3mF
8pc87e7MLfP4y66srFGDlFpns4+0QvF3ZZlBW8o+PUXBqAnTieHGFaan4ZVnGxV6dKyChTEYMgbl
6q6w3V4btr56xNXucQ0noRkykgiIbDXm4qS480g8WdwVzjBSRH+vN8OumG5ihGLpf/q3OzAfoGoQ
ZPXeoDgOgVMaZTUT1kvD4ZXTWUa+TJHtv3/PWZvY6MpFr2E2idNc5tDm2ELQXdfu8yFt3P1UBr4b
0kgIGBl78B4bfu6RmMxxbQ13A6evTFxkFuGtsRXgEs4suLx9I/wggGDAnea9llFb31oqR5U1GidY
V5Qd4MGNWKKsdz/9/gogiX1Fq8OAhafBdtq4YiTEZqimgFH4blfSHZf14PIJFEfLd8TNTNRZMZt/
vIQinF55ykNER5gT+qGDZ0XXsy4kbK/lBKlU0EEXkZnTz7CdP5fmABThtU3S4wX5zxsgRvHRsYPO
8xThTbbZcnUkgwvDki0GhTKkNA7EudouMMKKpJweI/20DOXRwqllAh2HW/9rvHWWl1ZD4+vSH9rk
dCVjPRC6XRRxnNKzaR3CtQjmezFl+eBrHijR++chPgRypqrsgGXT2/Pr9l0uKGFmM8nXzDm7u7wK
XiXxal+t9ZYWsHU3OaWFid4MtNmAbFJmwK1DX1XaJ3Y9G2XS2akVBPatOmamS8mb1dRma84s66b+
fXZ/C/+gRxl5ZnHwOjKIPDTrropg/5MewM70wusqHXJ9T83oeEmWUWt6L1oYAR3URF1PJCNeiBGu
xc1m9/QFQxRVaVbomGUF03VQHyxxpuETX1GWmWmNn/IC4n04xmSLwQRGhPbIBr3YbOp6tlIqumIn
MNTroOi6HQpJ6TGpUBfTzkFrugpOA78NNzQduQO0ZMNMeEtlusaVGU+qrYEqGtRVxUo0wYf9xnFn
vskRP2i8mjkNgkb5S3sO9MyCAfQ0CDwhQLw5sqKPvqAjm/Mw43LCibWJ2Nnn7FBc+hG1yGerKNBP
34DAjdu7izKeGaoyByWuf+BWjkTUC9zdq4N6jz0Gm5ZhUcRPabbGyIF3N7eeufJKdIDuzhRycv9k
QfkDxyym4M99yKa1jndxg+AD2MLO9/PyGH0TE7qe1rbcrTHHgnyr61aXjkMGB0f5z0aHYmOhX8wh
ME3gcAfvAaCviwYdJp63mlERQZp/9E2wJ1RdeI4zCy4TxYGl8e+IK928hcJAUi1U7aEgkBifGtYx
caotRxliZvJOtW4zo0nXP3r7wDyfm6arRnX/jZGtUqNpdtDUptlBew/w3MRYZOUntu5tFkvEd8Ub
z2ivEKQxsXVcwatnGPEDNszd10q41Kc//zb9QLPvLiWTXSGo4oOKNxLmIJKP/DgB7P9qYo7M6yjp
7avlPm1byPU7hb0ypQsOD9/4H3SOGP5eab4G5DJP5LGyDxUH2ZSBCWfmLcm/B9nSRoaj1zWxWj9F
uNCanZ4XPBLoW9YpMLW0Mm6P+a0cs5v4oFIVAg6cLj71+uUmIk9QKnEhJbi9mMBVlEHkeZaBInId
HhnOxMoh35wzKuY8Z82dtbAS1TGSC6Ra68TazI6eMbyci/j/8Rigp7W526TfBxhSdNua8ZKhb+f0
aiKPyIKsvN7Ca9sJgOBAYyhD4MmZUsgZR71vhc5Fyhb36IYILqV1IykSfHh4hFh1Cge/tLJzycVK
jvoY8Ywo2lC7uVapXjdzpf8coK2giJ9jJ28MKgyjVYfwah8Fp/mAZL3hDHGccrFY5hGMNdvsczJ/
CdFb1/nq5VMjDTpfy7LfO2fS53hM0dRggqEZks00Eiv9PFo7A+ugRGBtKoN/Z/pWPGk23+oLw1Oo
neUUU+6+wq0UP+bxPcyqat4n0RUQsQoZTNu+61vGN7rMBW2YIPiSRtzmCU28D6ewaonfGIPyNZFK
GfxAcNi0cgypworouVVvzKXtlG9f5cP1Uz5bm/QHVdOtmIbaHIpXTMY5789NEe3yqiJlJgmQUqcx
79MRq250ejhzM1ABhG1jMlVpDAmysw3f7Oj+6JdUw5kUR4dhGFyzhd4wDX9Dk7mzaK2za1vCJ/Ov
OeiN/CmkpXUQoubhp6xP6hPEv4Lfttp0p8NDXK0GkKl0bx2XAMjoQtFbU3Vt506uMrcBacDixUhy
kWKAyEjSZa3KfDk/xPVL1Mdmj6rFe+N6aAeHbQQ2BR+9icdzFUkGcEx3STS8FS0+vVx7snE7PXM/
T2/j7gY57PQGKgxgb7i6gdGGecHw2iPv1r4lUlpIbAQnngmyEOBMxnfr0l8otPrad0M474gzFIx9
+l0IyBfGfGIOSzQ8B72J/iYarUBmXf2h4/Wkte1JIIes52f42u8nZCg4Kme1p4cX2Vd8Vlll5vdU
sB9v8NEjxyZGCNi6Pur0OgbB6fDPNlbroI6bDst8v+09pU0CuuRvZ1RnPuWvxHyCsODMHu06+sRj
vIqo4w0Ih+ChKm9S5cZJIr+gtp21fZl6YCRha2JJiejT6rmX9dmQkV4YZ5FxJM49dkVsL+Lqpqt0
VB4cdGSsR6v3ek/ZnVjKTiQmP/J/08bur+0GMqcIFVZcBEE0Q+N0WYPrIaTzMH1jo7qgETBaPza8
EhPDN6n0RCSGTvbzM7cDTYokns0CnHCShqnqluk1VCJVDi1P8GqqYkrubXXA3q6rV83g6H0LYScQ
8Eb487WBrkm6+kW3xw9H9ehd6z4VTO2QFTi3i0sZAGdDDffavkIdW6QQ8qkoUyeEFzvQoXuCTuXc
743eAnjGOY6uEJJ4Ac7r5kagXXprB+zzK25TukOpzGF00a1oGn9JvRHyWZTyAbKALyb7tOLdQeuf
Eyhm1mrW7cRaobGp+CEfe5tZ5vbcglKR1prc0diZswbwjmANPT1ZR0eoyGjpAudA8wYzQgu3cQ/C
Hi20dQN2mILvMtCfwW5XpY9/CMYaC63NMXTgA9XqA436C8Dj6uShnneQNjWxE18oXIYp9HuMgDy5
J1gt/3V1nvdybNtkbneRp3dtmRxdHfTTUgZRy+7Zlx5pX71FJuIED478NdoYG8/SseQ5DFsmR1w4
+tUmMRybKLTWSqp9HgOWpmcYxf5Qvps/GZ1b1RJFjLZT7vseRRYzDiA4bOULXX2cVQsZAaBAbUUW
DDEEoRsHAXawxdZK/Odan1eBgKmrKFtm5Q36J4CIjenFyD4IIZLpZ7HZgs1HOzcqvqmsIr9RmVOz
TlL0tJkARwtyL0f2V9BgCq1UWSyCwv07KB3xmSRZqZxV4mEmPb2MJdKb1pZuAQCfGkVgu6RD7LSe
Shvq4L5ZVDoB6Iy+HhqdXO50deiRF2Lh7YtIzK8T+UfBih3oyYeG6G9HlW8y7agr6jrY3RjC9Qa0
c+W8jcpCj6tWilqiFnx6mNtm/UcaqPeo9AUQh+OXb2/UZ0Q/S4Ax+lhlz37/NGeXNjOAZv5PiYch
t7SZ8KJiiRyHa8eB9O18eQjzGVdraSWLhXFgsBVm6AvkWR2AukCbPo1fpiF9Sy6uSCyJUHAdzrAk
sOfe2yCg2oa1EH4HvfDAzQPYrNJw9VSfSBre5oEbU7pG/6VqHfb8cfOLvb6/dkC89R78MA3gL6lh
wTBZquTeWXvDnYPH4uVynCtrwpfX1yOIvz9T+JusX1lbjAb8cZDTwGlk9QFA0VYewn9t3hF8W76P
fsAcg3z+nbDPF/W7SrzlNJvcz1Rj9xKfspant3ldCBo4WrlJcfkSigQSEFHFtpyKDfqX7uno5BW2
PfsTRdAin4BwNr2OFMCDoyo1kJfDQw1/iuWkB2yCCrjQc/5Xpl0FpwrFgi6tG8Lo5p3shcBfz663
eLOWv1ulS5+PSLasZYH7FY4AM1YSXQspdEW4jfBYiUpB6XZypXR30Ro6nWCkF+zunR8GndzCwHn+
flZYHbPfVbiHiquFcpDvDTZko3GvesoYCrlHxqKaHIDw/QFCjTnDb0D5dY/ECRba5fpS3Stavoh2
zQ7HWUaA7Y02L8u9RjHr4VDY+r/BaxTu/cm/RFuriZloEAtCQzUth+xF12II+6vH7vdAcay8rzV5
3to1Jo8yfFunHq8zzDYois+zS/rnrlqe40d/2cBf97pPAJV9M8FNtIK3zIHXwGkXUQz+R01B2E2i
a/3VyR+pUTklQiRg0IAIvA9t6UUBl82Oe6tx0BPYuod5UZ0i+hTCFh/QAs5Hv4JmTkoOlspzZjKu
CaEJjVOJ4DwAHb8NZHgbA4l0OAzbW7IhHfSxmGdtUZlBnrO7Mh9bZh1njTXqY4dgMNBpjXzEqfTZ
P/HGFEMWZpXjA7B6aUgXknFKc7yUGN2LeV/HlxJl6r4YV/c6rfRCTFN7zHLAWpy9Ctvihs37xO09
VAIIQvZ7IiZH68+KYhxVTB5puuBDCBkIDGXpzncsvENF6VFe7iZzVXADU7z04GnqtjbCi7C/a+Oj
PD1zefSxouSE3IyfPV3F7zRmj6319ejikSkzhcRYl9DSLZq8UfioqipauFb3eL8dGAWAgcIzuJur
NrdLEEG+zbE/ViE2GeJYhBtldhRfxXTwIXIVO+wDF/DevxPU832QWkkQKZyf2Z+COj1FJL+4Hqd3
Mjw8C4DhNeUEBeXDo0xVCsNYzFe4m/uA1Ybvp7OjMHb7N9GInb1FOEJMhWkhyWBvIO6QmkTjSeXR
z51xSj4QDYr9PlIouLyvnrLIOgXs6GMj02iWcVvcOKF2IUgv9udaDHfvDPItsOL8nAmv8X1lgF3r
agGKawJtROU4zwaDjTWR19B2xJX1KzI8ZANtTwkuIud5IyqAZCBhXLcAM+fX81PpxYgW6/KCyh9Z
IHvY32Qxbpr87cULb65rUUE7OSLGusfU5Onj7YJXx2n0vC7hzqC+UeLKbgEiiRYldsEAJQBCgvFj
fCf6wRBzRbofpNp9oh9XuLf6zXME7RK8OhcPg4lrv+AFhDCHV15q/79CgwSnlJ694LUR9rU2+RRt
MJVPMet85kHBO+hM6QCtXOWe+KUiz5qlJnsdgi0rAtMsYfHxVldqNW2GzpcDTEnNkAiS57RB3VLn
DOcn0urDzezLTftokygGgkS7YF9qRS1O0Zjgwk7FXf2cZrPQ9qou1KfcInBJu1AZQrDk6iwbrUWq
gaNyewQ0lx6c2VLKYru6VB+drM8B2gRy9aE1TcG4M06BzSMshWn+xCfzu4eK+ZTiBK3fjlRuLolz
DmypF0tAtNIXe0AGKR08dfHgXwTE1wB85Yt3X1Ogn43iqUNfAc4lJx2AuulXMEPgv9e906ZfdEBF
4O3oq1J8f9O6+rC0lFfc3KCkONelLnceCfSUOjkwIsil/0d/7KI66zMP1rufnQbyGxURyJBlErWf
pY9V49h9L1M8ORMlCSt6ryVspk0WmORrVGCVyT1c+4wMcQdoXZMQLTjKs2zX1xKPUXF0ik0bPSst
gZnA+GQAIDxr94R0EIcNmq39TgUVn6HCrNsYQvev1fIGVwRohWESpKA1t4YZeFbxzpUUD5yHFlpv
mtdpuW5m0fjiOtc9y3kG2ImFUXVWdJsce/ij2q2VdIt54J7k+fp31cJ+f7dYzT1A3mOvuep7FTbU
HjQuN2NLNk4LpxHgOvKWhaQnsJ2QsZ+axbno1TIERGpYglmEgVSu7XwRi9zjadbEJtVp6MinQB3o
aCgRdQETrFhDCWRoOo0mFvUv02CnfkCgfV1cX3FXp/dwn9ZHY90N0wdGw5Z/YbCFTezNHXfIgPfv
VxQiEtTY8QJuHUy5J8XaOC+Z00DRAaSUIihL3e29eT2jdPytRe8r6GT456ms7umrwmnAh+MJMxYn
kWdl3Zbve4id9Jki/VPkrW6HN7gJ0LrgAFC6dhszPOVk9hzYCj4Y3tUnxx/2YZAwsngfo/nFBXja
UUNcq9tZDeJzw/stc9d72P4mA0VluWptXiNtFeS1eoP5/ECu1/9CUYEN5CPpwJ97WN6EqKEKBQMt
zaET8boq4iH7N8N7nvG99gSktGRgOqnw4qdgNOwS4MF+FSmUgnIKI8QPKjkvk5yXd2hDFZ/fgyxr
jPOFTpSW/KcSgQzK0AkEzADI7m5N1JW7oYJF+qMkryoyq3yZ20ik6dxvsZ/ZX8cZ0ZDpPPy2MIGe
GdRdtdgCVO9h5E/tV/HTfXJB4pniXHvkMQ/4TFzjaVYoViLhE3OGnVPRO+atSwYY2ofcaUb6sh4+
mIKp5qBoLhWPSafh/Ty95UL7WcW8jdLL7Pqza8glBrVtRBFA8TB3VjbGGLIZCGUNh9kXrTcp5Jx8
294YhYLIx9BAKMCGLAy/5EIjkHkY1ySJVO6HcKEDXajxpa0tUfErPsEFznsew+9Qm97WDAIb9whT
3QDoLzk1xhxt5af1JKlhU6pEulvLf2vtSiPlneKeptRBF9z1JOgmujUPNSzzJhCbpJxo7UgxyFUb
WLLt3rGNX0wf8KHjw1Mp9BsjnqkwNySea+asdcCW6L01XgU9H9TJUgsBSvn7mr0pLT3+bA9Gyyh9
8jWeSX6gu2bG42h+QZrXxW2hHIG5IZPtriLcL0WTpuKizyF0RBv6BmwydspOegTNkBI+wkNJmn5e
5kgq6rCrtlApz9pmADTbclkqRg8ZhiRptQquETyZ/xiWs7aownQeD0Xmsomd3AayTxufCYmcaiuL
Wmn19xTrMLYvpFVe5vy36Aw2uFTl67dqrVuelwSBM3LGfSAUcCoIA5ZFoXSj63KoGyKrJ0g31w/0
pphRpUM1e+CX4ovF0+hQrJJyC9Cx08kiDh1GAXTYbPNivWVdZftxzszba8qpQGQ6nirSeGkpvAcX
NImQpWzV8JaKFfKMmOHzRmbVBXF2JoyZA8hZzMzQ/UzNqzLcnqiaDB5lVDJKDGqIkI6E8g3QYsoW
NPO0cCIJ9DAncst1jP0sT0Ddv8kEo/4nliYerx3XpG37b0dxZUnyIT1pb17B1hV40xdS3K2k/h1X
9nVj1rK9i8yOc7fsiOgvZ7UIlvBiuzItgf+3G1prXL+r9SU/qc3w9eq28lBsXLWKVB+73gCGIS8o
FdQYOUorLulLJU/+P2VhxsaI1LaRXTSGuo8zIMXG281/b/d0xDzKXR6DYO/S61jHiHmbFCXuKRbn
aRJ4xMjy7hNaZpWY37BBwOGhhhRFhcQLI/dqv0XHevap/sfZSPfeIfHKNii3mPJh3ZAMM3tNGCAC
vukRRb8dSO0P+ipxiLe3/BHzbeM5KEDeiizMcVZmzt40zppk8NgKzD9qp9NtxxEk89v2X1CYcKbK
SSOsnJsYCeiw6ckZZr3Sm+Zn4Rk+Li51kV5sKAcUXGSdA1LRIoq0naa1124YWVc1YQYQUa+bbYHR
yVEkq0lJkqu4BKClCJVIjYrDsIKfXtBlJdm8VFRrrtNUkWDcxBbdLwLWQrKYr/yGM4fW4I9u59Vn
8BfvBU8gJd/F76s6qBkUIFXUuFGvZJehU81tx5G4m/OsP8vWn35A/IZ9Q+9EJL9Gy/azXUu+Yzre
F1Rx60pfRXsVHJs1CabrlmET93IhVHk6O+PLgMtoeVsvXr3bLIphpWh7t1D979Saj7fZzEjgVRn2
k/RHq0dlWlx9n27I6HJ0SIWA36g1d6LAxVYCJn9KIh3MtGphQM7igD5uTNOx5r3vIcst93/HNDXY
JYnQLws+JAQfuTAChKNWiMBJ8lsfD3H08S+9L774vDC5lu+ZPEmePLuhH5QuI7Z4riDIiKCEPNr0
oTR9U47DIzLiBPdzeKzQuiivIR7mNEK9K4PxpGGPmOno4OAhT14Ou0ypAOyHHJyAwaCJDaNJLFyx
YS0y7DW/SmC7hNsC69Gwmo/0a21lxwUjpSvTe+tDYFNtCT4/S315PIWyVsn2LjVBHSYxTLrPFpnt
lgWR8yIfF+meRvC79m1uGKZ+turi4l96pADWDZLelIQUsZt1SoONjtD/WpQRD/TJpKXhmNTVlVMJ
40zvHuCIBgFB3tqV+IXlCYOHCxjAB9hmj2OLjGoMJ2raFQcMqbLR7IA4ANaPELCtIJjCbUI8aKN9
ZSytQ/9quCm2y8cXIgidAWNczP6mfVzcgKORa0lzlBHjra6KJIpIrJdSy7khy37isOj/8HsK9pJt
OKETJW+xyliFcvEmFOf6wyHNFeVyvF3skuWwV8ko80uE33CyfGMkv5E+a0UMpaYDJgftiGYEQvHf
pxVQaQJ+wDQfy5qe+kvYP1EOLJslDF2CF6dRHW1a5HFYANet/HjGdTGFxO7zFnJ7GkqlkFWH58YZ
GLwI5IVxUvRPguUI+3KaqsXaWj53aK8U8ZqG4oCDqMZDRTj1Wn7b9Dx2amUvLiikj2HRwCjJGf5V
bOicjQV7OjPFuqT7lkaqRSapW8J31IGMygsS0wa4X+15pLOtRIxUINjt/azv3mN6mYJAL44mjaxb
gX5v7Ws8/0p+lcoPKulc/ti7NjAKlJvmIGXbJBazaLgLmdmUeEaTwEz6A55Wng6C+8gtwzm5iM0i
ujZIHMnpTyEPXsoPbrWd8QGtVlsuh6SH9htU+hv3aglgywbzXdnlkZxgNv6jaE6erCdvLOVOMuP5
uR8jYAjnrPGNuFfXeZJJfQxxymunQb8hTs686Mx2Tj0P3dmQqo/89J99hAiUZvQHr1TPLNKEK6Ce
KslsS8IiOByil2jm/WPSYG3bYd3HtjjShhGuY+A810V+u5rT0fHpXpYn64sdYtGtKw+hapM+VoBn
u+BkjWvrbScSioUZJPb6NTZ7dB6Zs85xW2gUpKZGBDVyeFZbYfzq/keDsEzu3xc6f6lPsh/pVPXh
AqwfFIjabzx8/T7OxwVGFv5v22vuFoltABw3jcr1reB8ZSreVivLqwABQHkV4JZNwnAJh0Y+2Uhz
E1svIBSOjYbVXf2/4k0BsK+6Ta9motJ5ZgUttFw8N39CBUQ6Lrwt4kjdGYwzQCnX9JutHcD8jEJe
jTdVrtl+wAfvS8TQdafTW+eLG7z7hLyA/v5pcUte7Qw1pjrIgWH55FXY4gsTRCbN/rIzCztVtuVN
mH4DDzIPgb94EoHAhgTwpYmdPSLNKHpmh6WsNlbCmFbMk1E22FWFUPPgi0xiG45QOB+z09LwgjZ7
HAPM5UDTp+4CyCsNC1/UzAxP7n1XH9gBbVx9TAXSGSCBZElCxePnRVHvsrKOXvpRdfTIwUW5n4dS
dgxRRoMZlbFNp9txXLHHe/Q3kTtah9bfbCaXpYbu6nqJmVbzuK8vMUJfrOToorkcEYFQDiDfmE5I
9a/et4ptUh/nbN1V9sShH+toShxG2/bpsFCwwinrKfx1s74aAY3PtsODtdX80hIbyptTx4a6of73
7Gf2PtrTdyvwQJreUER+qMtGqg0C3sFs0EKMtsRw/f66ostbJYi/ikf/P5Q5s5s8m41GIu9Tnlbb
eAETqN44ZYVZmt/KIFBKHXbHKU4ZKgHr5qCsEmp5W2NhNPYa1hoLLW3iyXqmdVbMrqLzymFYe5L2
psRr/872ahtSZyZzjz9Z6V+/m518k/7fFlspzAHTdk8XxqGebVhw6ZjD4elGjV2n+FfZuJ5EcpfM
L6kDEedMZ+gz3JBe5WRH4CuirE7USqIfcftXLSDrIv8Rp2zzODpOdXID3kH2kgJ1OtxkuJpC2Bz1
YReEuZ8t4GFs7Y5b2bpAWDV/MQ6Zq8YXQnTwXaTS8oT69RK+flYyjSEvuh62axn5GoTUm1dAn5wj
3lHg7zFqaFVFeInaCAKOXShlpjGsDPy9aO+m6kZAEUImS4vrqk407lTMymQNoq4zgeJHBgneURfo
/jB9BFtNPx8lZsqL6iTuFqM3GtT2WXFQS+Qi5QP2wdmHk/wg5Mtq4xI8ZL9AYRdxLvaWQnx1lX5k
/qHK9qznqVuAJ6YQro8Mg1cgKZLIb6b/6VoL1c47aqmDbPy1rdlM+ROWnusF8wLjwAojQFTD3bOw
lI/r2ZGVliRIUJN0z/r7Rj867iDX9Ls/MtOnwC7R/Us/A1FOk/2HwayBeEmApmaQvD+FWOLfQhCu
maKawkYHKoBA8qNoqx615+l+IkjIrp7g0nqh5FR7ZUpMIvgkeJxx4DZC6yw9fvF2KPp78QTrjajS
TUhSNr+PZ3eUKQrVRJbbI/1bNcaMkMheTUxYU6DOomS6xuwBmagJNzVmDOAKwi04DXBtZIiqNK7Z
A+nG4K7xQ0WZ+8SuaGuTquSSFZ5WKaTrohYm6s4tRK0V2RRxlHbIknIy8A1dTJ70976bTYs3+9Xe
sxAMdrKXAT9or7I0+0YHl3I5UhHZgKOfphGwTQgXWQW4RkR9C3jOjBqIAIopMq8yBslevZQceCg5
Ux9W+DMSB4nl4j9SiZZELlUeIHC5RkQvkpoaSYzlp7yFx0CrwQrZPBOz77cmFJf3PoGRC/Ex0+jP
v2iHUXr7dVzD48GPKVKfL7DXXowV6WGPQHAJ/D4FDdMXKd8LKPQs4PINEqEe/Pfj3O5a6IIoQTQh
WwFc5NHDDXuB5Gx1CEn9ewfJNhU3SBPykP2y82dtv5WImrUmzJ4PEOoxwfcOMLrq73JpXyYGWGkg
ttEqW/jR5DL6rdiZ9dU5xG0VJdgrmhtc6ci6nz3yM0ZJA/VDoZPio19vDOYHYKDeYrznC1hQ4hig
URPZd5NlQ4Vjf1tbd0v7tDO/a3gmziFiW1dvpi2jUakKALFqqAhOdDG1uY8HSZQbS78sWe6DB6Hr
xZXHHaV+CucOTTXvCiwH/4F3loP7xFfy/1PybzkhPLuCGfO3dnqZzl9czIGx+pXGJyVGKUxq2wpJ
w/g1ZLleIITHJydZu4B0boBm3yJBAojFZQ5MCW8CI1RG8Nhj6ULzhb8Wf3StZISQBkq0Y5WM9gOe
jCxfER6nG1/Eb2T65bytr+4MQEgxVXqF/Q3JkvCrzMrwIrgUQFLr+oKiS9JNRQUMGAunNk/pm1f+
LLF0nN4El3taQwN3QKFFwjiz1kfUYXhC+oBaMsR8GSeIqJfMX87two00eC4YLOMDTRzwXASjD4ot
vuDJjzj29UqtNzId14kldNMigNTMTsFu5Kbryx9YDGh76idAHxquYFxiXxWrlH48kBl4qthvrpgI
ncePqkpcHOASGk6qni6Ivw0UdkM5D4qvMpWFhr3FWmHRpO0h5vWf4PvTnnROimD7B/VvYN/N7pvy
yWk7oa63ncbxy8srhw+Y36dUVxtYCRrvuIsiD+qQ/YulRj2bgJnhjiAvD+K4QaJJ5AEFTMwpm0Mg
7+mS2oCxNLDccQeT++iSXAS5+PqO0nR26WpiA75EIrwfWDiMvrAmK56HaoLEF5T50Tv9QV9KIxBA
Ss9tPIGRbUAivU5xjlAWuwtkDaVvACKJjNzN14DWrhOvHR1aGMVZ17ZjhIE8p6L4f/NFIYta1oeA
EC/+fDs0PdVbYoH7RKp43/7KtmMCaI03+x6swkO4KoA5+qhToc8pR0FjuAwyqDUzLZxE/6pB0Lpn
55XFlg495W8UvFWW8XRyNbzPlcdYwONecasFNN4lPcKXikwHEK3bdOjoFT3fEwtjHAV9S21m1dAG
t+5JdPMqQO6lNyGlSxPUuA9CKX4Rqo2QC/hM4JydR6sodVyz2pajJjtLxBf5iyPYLiP1Jy0HYQ9t
FLpWDH7UiHSnvRE4eAFC7rm4WcCbkCj2bjtenFBAZYGTmAnmb1de7bhCxwdaTugV0OMikUTuy5bj
33OjcxD1KJzXMQmGQG1m9miyPF/eWVMOMlk2QPwtHEd2zFVd6WQSMPAJFqyj5+gEBWYZmUpkYPxQ
EsII/Sph7k9PR6nN3LGN7EPPKvE7s7NEF8XV8UH3QNTeDBpN402JmhQ3EgaEFv48L8pM4mbKP7xF
X/Nu6aAs0I07usIFP8q7RpHz4k6t7nuPTUM+koXfWU0chV3meXuViLhoQfIzu1jaCHSQJbNgu9rh
Q7fMzVeQ0mFVj/923dh8OrAqMmD3VJw3lERrdUHjae4z0kA2U/2r99RHoN6daG9Z1kK+6qdeuRfd
Ly6+wY1kltn1Bh5cKqw4AScEFLfq6aD5YMqwlaG0xjm3IwlSsk74ZCgax4DvEzT/cB/0ZdNHKSma
dYLH4SIXYsNbRpmSP6GWzz2m9w4DOZiD1aGnbtTi0pgtSKsDeU1fhBsK4pVcMqbmUztXyHAaG0KS
WBol+8lpnHBVmPUlRXUo7RkF/bQ/WXfy6UFkc961mYuopUkVuifjeNsVoH5FeuFsUWY0yzKlqK+5
sLj+/9QjanrvrHYEWUUp+u0rtvTWHX9dfIXFnxMaPW9Qg+2OxbGAuvYZNlt19/9dsfHiMHdtrStW
x8zVPBFZCHaYjPPlwz9UHhWMSACjuKQY/F0Y9BuYgdgZK1rRQeQ6eVDmyWhhSm+KRpz4j7HARecT
BJ9e6o3Q+wnlpeCUOK7BAoFyX4pccSvuWufxvPzJ1cb4SuNSpElLMGPXyiIZjy4XuUXpm0MlbzLH
IQi2+PkBIgt4pVOL7jcI3TaLPbbIWr1mbPHIct18mkJvWkr8OGhm50P/B8O2WXKfiB94bgztjj0I
4iCYlbZcAVMITB6Enmx/1m7UhLNvNWTYcZ8g5HbqejF3waVInD533e0+5o4IT/u50avOLXLX0EDs
7PtfVAIAexM7dkFKdVb0PkgM/dq0di0GYTlLddqBEPHIY4JdFgVusqHkoZlgdF7BZdLVEeZ419/P
oN+QmNPQIg2p0mLjcDbOWQkyLTW/vBn8b5+Myzu8YIJIcRs961b+wbVQW2swA0LWwQBDaZYumBss
j+Sx4caIPO1JiHXqRuEG7KJVewIl5aXm8LwXOFDgtIIcnUdrWmofr0CF8ROzVZv+LVT1kIPe//8l
sen+t4FaHotZMNcnMNHF4TeDvBo2c9w5qEoaqgqDbAkDOd01OzWi1U2HPdm1j83D5aeCw3riVSLj
UyGgugW8RE7qTpgIrajEWh518+1HF1N9jvFW/3Rym5IShWI9PVaQRnOduate0S50Qm6I92On+sAb
NCHevjTF8kv3vZwrIV8oM7YmDreAfcqtOg+a8sNlpwL4Le40/esD5NS7U67QQ3xtG/RRdCohx7Xy
EFR2WT0wymGtnH1wwVsnExywGWgBkVM7x1kRvzUXGlEoMM6N8sUKM8QqiFKjvL31UXReYlClShFd
obUavxRxJOQaZLu/TRUgw7S1n2f68if+b/YqawsJ5+dLLFOMw2KM5W/Fb5e3bBSm8vUy9vIq6rd2
BfyOo/EWz4iVdXwfIES2S/V81mSyTOhM1t9BMKpmBlgNv8UFcLo6VmhX1JTYZNB/RfpxY0J/YGOq
1NQj4x2ye6T9/PtTguNlfASfuMIaS4rV/6OTOYt5yZkwJekvqNBYFQFoBZUnErf6s0oLYmcGwtHv
i5qHoAEqXIbTnqwCikkuyoh8PGGOG2T5GHCAu3L4i5JF+HUPZCQvMtYN1XNoRjWj1OSLdnrheN4z
ThC8srhJ5CXc1hOSZaVUK+wMIzX8hj8k7cVB+8AHjhfE/PnS4klHPA/w6mXpF5TWBjqAWC3hFsFV
55DXkPrTE7oR77FPSCeAyqFk18/iLAZCvB9xLFe5JDf59mj5AqinztmI0JJm+CpLhfcrcpx9h9gH
IrgMFa2tOQmzeZWalX5nmoCUAqOmVve7okQguxQRxOnaJTcNx4rujkI10/bm0bmao8Hn3qxa+YfZ
jIBGyx9fZCzvaUufqsLwIoJoEpS4vnLMDEyivWJ3DzbckDlAd6YT8JaEtFKE7OLHFQHOKMxZERBg
sM3Sr3kIdEoc96EtbjjV1vC32HxkQyo05U8iRWa4l3WEWyUCUUyT9IjLcYQnF+Vw4ZV07HU/8Muw
Jjl3KSNF1eL2IPPwkCwUYQ3pf5suNDKr2/uIQxz4qcLXDHlfYDLZrb9CeainOW+3rCiroAvIMGxL
fUi3YEY7swoxZZA2TU5OHG/XV1X78hs9eKHfZCETS5RPFNKYasq55WZ72wx+6PGMb3upfcnFMJ4c
MEV3wiwa8twduUY0yChhEDPV74Hz3mcnkqQ7J53uKle1f92yPxwDSmIAjd6vxdAbQciqid46QQad
I2KG7zDRkq9aO9LLVGv0/YJSWjGT64C2H6W6jbV7k5H3PNVeQxlinHOXP9X0kltcY3H14OxJi7uX
9+h1rGARnmFYYc7XhZzdl8UtsGbWDc9krjH0hAErHnbvviE5timuA8kxdUoPZnzCTi7wHwwj1x7I
ZXfQ+t1tXXx+CIgPieLWBrLCTqsCuW8J80ohZhJrjXGC/V5eJtKXCPfGBb0dPpScaZL2PwkiwMNg
TMLZid66ZeCuwvwVM18dGKjCIoDnA7vZFCzw1WsObE4qTfoI/nyB25h23pppi/lFZxu5Fnuijuea
V7bi4/O9Tvn1Bi62NZNpZvmS7h+gYrWUxQg2SZg1RDdDMm/cnr+2FwE8E67znk5xkwMezKB6FTuS
eOcWcCfSwIhaRYEUE44rJvHtbq9aLVWmHPfucrA9ekfq5/7jJWtYtBE+/wyfrCSR4nJk5Gl/6nHh
7Gh327M7VsJdvw26Md0asLiUDxMN2SUm86/sQGgqE4swx5sdLZKnHH166zF6LUyCLSf5Y1rMjdjp
tU0aRdnK63zuNd4rTEVj6OgwpU3+aXB/WiLkhuOyYC7KgPfEBZPoYXt9SW+g54wG9BDBxO2D9+kL
j/iJ7aWQegW6qQQxEtt//Jnk6KPwzm1TLFMhgmcGROR2+8Ndyikcd+me1csqlItbZ2RiFj/DwzoX
lhfCNdVjX0jP4ySOAEnQWylOzjXxfVxxIIYEFyrZBAJtItAhj4/yXNv54gJezaUNqRtHjanFvz69
BFkLJPpVSp6LfX9nDow9wz4VqDepfo7ziDxyj4PAbBrvFdEQVZdJ0Okh8g0AQQ9uuvZHkEuKN6vd
OuswzWXfWsZ4Q2gXOdAAqSzyOxCQIZNdT0CU5mh37WoAWkFD2rZbrxmxRbF7RQOiyT7ykeOu5DGb
vs/TLyXTNuU583n+qsGCduIOXit6SKlyOzArCN4n9omhby7rI0RghYXi8RuE+uKoSJ5ah1wr+CXa
u7AA+WQR8xyRSpZCIihGrLH7OZLLl+RBeJboi4cW1V6yFvtjQ/jNK3egYu+WhH+qZN18yPy6ILi4
N6pv4k79pqo2G4e051QwWSTWkCYHWaYlKvBGN49Eg41OfPRQ1kc2FPL4+/e5Sg6o4rQMWcd3aS6l
wy3jkeBYBmPR/HvXdccMDD6N8z3bU0zUHcY7xUe0zqgO3ehfOJRFZWZ+oGtf+Mtvvk+F4N+zn9S1
33vZ4mbROyETTN/J/N71CHqhNgXEDAjfzA7uBvuc/M7tQpsZZvblPJmZFzhBK9KEvRKDHyU/Owxn
1GJRefWVEXBVGG9eFKKssPLPnHV8TeV9EFKPbG/k0Rw3B8L7E+NBygwKM3YWVFgQW7LS1elvRFoj
pLljx6Umjm0RKszfOnlV/tDK10DU07lasKmsAuUg/pkDaSOdDVDWnaU2O6pXAskfzfXUDmaNdpPg
bl3JguQO1o7eyZWzI3zFR7FonTK6n2zzo4LThr0Qmfo/1Rrk3X4uMHL6MR+/FCXhyd3ruVwUoD8e
AH1Np0I2hKW1ZJVnaQ6qS0GdjhxHgx4/k6NONXh44+LY+Ky8ZcmkNWhDhZ8iw+kp8tZ97qmPU3xd
RPekf8GjVgFKvfGtLmrpETAY2vn6LS2A6b8KhSjsPCoVFhOfhqi/KwnlD7WUKgntD8NXrZDMFIKx
kOKoNo9LRkJ5taxnh2uWcdVwiYEHUfoVHGgQwjjnE6Z163048fe5nNhX2dUGw/s2RE+CUW9fl/+2
cLLPraNqjK8Dh17djChPnRDzgTRyjy848j566ldSFbM7ymEjD1BuN1QeRi/C7mzrSIUHM2TgQ6kf
ebUkfo1zaK5KMvhTUPx46Bp7/4R4p0+vD2D2Yv9VJlikipp0p6c2EV7wqVQGaX0cnLFd7WqWJfmi
cvFRGm1E0ukGBLs4GlHKHOiciakCeZaATV1Oudbb9Hovd2N9uwW1zkOz7tfg2eYU2dPdYCB5gcLj
U3PzVZcNmJS80m0s5K0TvmEds3iGwW3KTpGZaz51FbYP8EvnhQ4E8U26wyf/EsrHet3Sb3Wzy4rF
TAVt2ZcCpwZELFlfHSGU81K8kk73pFjcm8CjQ6zMAvfq3rlsESVT19Bh7Vk8lSwdZp3/qL7hfZPd
TF6nflpid9XaB8A6H43/V5CmE8mFkal9Wx2EgickVww0W3S3djn7rwb+f4tYuvcLYG6bDHxgHbUs
2MnkYtcgbKOBuzuMpZmGAKMtvwgNYlsqEM6OY2Uupz42Rj+jHMYRuTem/y9X+//pqO3HslWi72Hz
gcBFypGuHyR94rKdGYCyDfs8cw0YulN97Z97HYxrw6ogn5RMhcfR1qjty4zjHQA5yfklRPVUGwCN
FzD2n3MbFJmFVdaOyqeLhxtFTlPDBlv4H5SZKnc2TziMuqthavcPuK5Xk6VIXS47PR8cisexZcFh
a4SoRk743a94CerxGaw77UwpLRwYQKLgSIcebGOOYNRufkiLHrX9A7lIie1wLKXYlU73HYKSxO38
9FDMe89g/Hziz4GpfUWPc9GS/0/ZgYuA+7dDXsun3D10naxISPmGZrPgdedwWufUmTr1gcpVsFAA
TSCTmQ2jSzHHohjkaWW4rgxu+YgO72sEtaY36whyLyWg/bWOH8lvkkgBs/N1mkAAOg5hGnwICr13
xcAp6nS18oa+xqR0VYUxzytcbYzzyF+lGdhzqWQXx6O5l6SSrO/MqXiorpCX2SC0UPAmXyCK8On9
XlisbIcStY31C0W+D3viWIxBj2KhLliQvGxqWto5OBjG/Qzc2Aspantjavwy2hi2pJXZ+HPQtymF
t/LN7CdcmtWkrGeprTSDeGJr3iI1H407VhOZOje7tmPBfWhrQKh6gu0qosoGBDwz4fLW1PjUZUsJ
oQ3w7XEgZ3GiJ4iVoXhdONeh3MYhaa91kjlOj4CtZZlGSeZ7I7vq3/ADSwq3fbbXEiOrwyJVC9QI
OtdaPZ4Uwu06fTmHKtq00EecB9zUbweZRg81Oddw0k9lmtPTa4GMSejHsl9CSzENUj0SnGr3OeBB
vXcRwrG8k/q/7lV1iKBhqoaom3VzufPo7QPGLcuq2ahvUWzZtSXODDd7FEIT+Wdvqxa6sutIOLES
kvTlc4qXGC0hCNT8HLnIX8xO/NlDj70ly9RIkihJPPaoENgAm+yKO6i+b7mCzhPnAiCVaZwxnVCO
TAPWKzjSgqLTEdPF40GiMhn+ajjJevgUmOsGugxseXkRZ/9cwjI5BITaxFknqncOqzYignac5vZ9
yWaN2pivZ6zozLHqUz41m76J8lhFrgb/C/++YW0Yh4zGODVt8Y/4gM1TZQJ3RAQUhTb2uqU/7gW9
5KQTtmMhLwL3akh1J1X8oeufNCILfuWZqhy29oevBvW336QSdPLqP3z9Hb7j5Nm+JW2F6Of2mEMm
MiQ9ApomaBN+bkJiTSoval9vuBfsTYdjNSVhxAlaHN4c78AioRYPhaG1nniqWH+7+vvH7nsls/PH
/6JLovsLdHhyD/c6VsslcmL7/ovckqF0SvRYX6sUaYXKUQ94YrO9YbstI13+Hvm4sABk887/AfDQ
3YSQmpA/RVQTqcqVoyXCB+ttbrHOrkgNjiBVAgbKSLuhGkW/2sEdv8X3QD/3zpsMr78+t/WGfgx5
TYnZUtnKWG/5mkKlsR01h4hXg68b3sryd5LpZyPxmn7gHQq5hsAj6bQOuTZKCrMjC1hcOOoIIOur
rsbwfySryyh5wBZizg3DKfdhHbiimMCtrlN5KHaZEY5/4jyVsIeqiDzpC55HSwaNPfHafPa/LPbc
XJW3Un/V4mGaeWuR5u0qEr620IWZ/Q+zuI/Tchiqyp+alT/sakMuDhEQnM0YvCbfKX3xDixIbIoC
LW/HidaaTj+Z8SYZRixEXGJj7VLqJHQ4nijPtfMLa+Nm/r0GRysdtMS5OEaQogC46baREdLfaBx3
9sIlDU8VYdd4uCm+AV/qISrqXK6EQFy+wSoo/Ks3mF8CATBginhAOMRjjE47nIkZcdVpWQvl2wu4
6Ce7eTDR51d7+F6vXdxXIxi6FznO26W+6BnEa6NHsoghO403k77Yyf1Kr9UNQJZLwWeKbGCbkzaY
zDvju+JdrY/JOxw+lxVvP2eudHmBRXMnKwRyiruC9e3IQrolznV34Mq2kms6AVGqp0CyagZdJynH
aBepZwhsUImfXXapxOlLU/OHqBK4lGULZjOaDlffhDWjKA6ZKrlDO0gzS3Mt6FlYmcmYL+7rb/NU
wgK3Rk0dCf8HyLpYrHJCJf2OtnTsuvvVlMXxGjzufR6joazJHs8xKTW6jT5GCevH5J4TlnVH3lkA
jLdrDK+5Xbh1JTEZHvIJUb/yG7e++haMC1f0Bqov494re/Hgnp5qT58cgweMwC+kHhJBS907cIXA
anOgQitybF7qD2FLny7ymJMEVAl02S6c/VwAEKrYzrIfRWe4X7vWi6eXl3lJLQ081tZCjKxxo1jA
86rTdyUpVgnCgJC9MJLYcCRvgb8lW5wVDBQ+P9GjBIBJlj/Ah4QirFmm1yG+SbaaFpC548EoRMkP
5yg3VMXypVIPJNQKgb8Sl4qxlpkldLJyY/k2XljxzpRJglPcZa+RpFw3L7qTGwYXD2/+oHRlDZep
liExq+0jtrpu8wtzqZkVwrQYrpZS6IJAGQ5bq+T5xgKf3QL7heXXdhtmCDeSOwmIGamGVr3Q5ng/
eTXBo177P17Dn3E9F70u91SovakiRtpjn4KPATnbRvNgUV1MZrHrRi5UvkxpXCRufo2FjEkRVM0u
fU/JVZbnxfzir75HftEibj1jYXNpLRkROAt7Yr9Y/GCjdqLYE5Pqqv5jyHKL926T7qICnAdfNeAL
62NEUJ6370qDZaopyQ1CiNwTCP6lvouyBi8dg+MwFoYrAds2/by0+KOiOpoq7ZwZRCeBsprg0bq/
1HcphDzLIh+8Dt2LDiTi/e8jcjsfc0n5QKpZztGms12sXkPadfEc/Ltetz3YIQRNhS13wduNXhb7
d48IzhwYuoIGzd7ajIQkz3xnVBjWgeMYqHlQXiO+mH8jxkpGoqa3hBZvesI5tYIWsfqrqAPOLvPJ
ivn+byUrs9QHk0/EGIPuXwigM3m7X+LAhqjScFxML7ssCqucReJeoUE3xlGoPn3i3v02BDpjneT6
bQsLAAOih4VgYaBCuuKYQ/tF6BvMbKTVF3yjmDsaTA/fR1ok4IHLM8UFqsXmk8H76mPQ54M3c5FV
A8HLaAfOYefvmouXSMz5TLC8j4C8pmsz6jMXUtAqzHC83feRBNBZPotmsYgxZC40nvz8v9E4LVt0
mHOCaXP+JfhEx6E1+ZVJZq16qY79DpAf9B0ibZxa9smO3ys+p/I4b8Za7d9jWwf3VlNhSQIzNfrP
HfWDmmcDvQQAMxYiakx/Fn3oYpzMHaxfHmIakuZNJkuUxIBob7R2TfArxuCf+l+4Bx7jRWBQgIHL
njbKdAb6lb/D+rMnUXDBaOyPQdxlkGrFs+Q5WZ5DJTKB8YW0mwNfwAGZ1xvXankzVvxNlVR02p1Y
tqQ1PZ/fVAY77TOyLUyKSXaQigg3ZFPH3YWN4s45VwZ1ANSO8/O7nKMevEClo70IOmM7LJfuRDix
wDWR0ZL9AezsfLKozze3N4/YDh8V5It8Oe0NDBBOH4aJDmdtL6E9uNGgpgA0kHmXY/Bum6StZzVh
xhhnMXRG/QOiOlbf08qPMiNt9YcggS6dDw0R0FU9qk07jzsL1P0zSnKlJwBB9ci1K4CO3Q57RAlT
YsVNdjjMrmkPdFqE7TwIklEZkwoHeJEfBJoCay2WFeC1VUMEnQ4/O9W9K5MXJEuHY79Ze6vJYu/t
KIABl8KDBP4VmDw5/sNP0ZqI2lZ6HqQ1HtkCkJjUgq3uI6kBrwG01g5k2fT3nYlrgMrMLgQPzxVL
KB7Dc+jlVJ12Apv7xE14uMlDz60TB+pJG9jpk/z7swpdwOohzO3tjWHoQBEgaNcAh0dHpTd9xsIC
76zj2R/hQwdtbMd5zO7m26G9a4VM2yU1YhOz1VRjzH3B/26PZ4+7srgnVVQcEcCbvZkCqyl0jdJF
hKb2ZXQW6GDMsxpEPzXbPgMtUnKvzDUI42sWQOtJWfZJq0vHS9hZFRM6RFe/VmMsqnaqWOMuHUIZ
Tk+ovGPsf/AP3qKTqdHCRV32JSjCJyQ4GsnvNJmtzxSyLpBpetHuXTVFj/ZnzpYXYc2wGF9htRMe
eSGRgPIoqZb34aRhqfWqYx8sFqRYALbRVzlOlMU8CJJnKNA0twi1EHPXKnBSZLgR8NygRH3mJ/y/
errO+HKclh3UwtJs9RTf2AenGftzWQJfC/SMuwoYaypCXuaqiiBSDGIQQ2joiNdaRy6iTqEwv/hd
fDZCMEElmPMxnsDeqZZ/nvwX/xDKFjuwT8rG1ank2T1UeqKjsXWr3Y7c8gCfwryr9C7yAOmKHTrZ
qp0HNn3hRE74eaKtHhmmt8K/xnVSxSnLjGOtcNrHnCrz3r5vWX5BMtfsMKYrIrj0Dow4nWDDojiV
XIB6xhG7enJ6j9sbhI4hj8gSFFgH1WJq9HSlrNlkmNvwcPB1JolEZkVHBkrvne5C1pMTZa7SzQ8H
fWgdh9YxRElFZxksHcnYyAV4XxTlMksJAzFje51+HIuDcuRSzdbz5vyWAjn2pGDJoFZ5SvyV5KCm
In6Vb9CqL24UBsTRV1FWFy2VFWkx7XPyVm3PaQnPV3M4+uVyq10PhBe5O7GiD3/5GxBWZiEl10Dg
oWgFx1JsK8ZYmQ4Zwm6GSCOsVrIUgjMInXSt+u25H7YeGslClgnG3316VM5fbxiPKWAZfyiF/1WL
cRt5gLBfpvi5kK39xqHXatZFkIWY4vGGZHzewT0ooAqOpwDBn8tXxCDquBvTQfPvKDJU8DEJJdt0
M9qW1LawBpS2/lAi4AhG10W/Poni4JHjZb1CGkFm8fcavgz+J137IF3u/z4ezKrr00MCl+9HFbb5
NkByzaobswiyY3FsqWhj4K0OVbeDWQERgDsUjPJ7SzTHKPkX+NJ1AVaQYEwY7fDna4wh1AMWPzeX
1UetWHToa0FOw2KMx0x7XpRZ/OdwRmPL6n5Mw5i1WiY/HqRMI3bsUQ5La1OpyVLo8kCdm74Y6Zz+
YV27toN+7EkXgP2Tbf/rr/3Z89AhIv4iGUDn6MIonJevGdlT80U+nf1+Wr1S93vbd3fCiseo8u2M
VclzI1ZF1gg6Xkzn44Cq60zhE0rLe3yKeK9z4EObsQLQofMkkyhXPfKU1BLklNZyePpU3/7PMSRm
qddR99rOWq6x/xYUtiT6/mojQBZ0NFbUCVdCqTq+lAOS3Ds5hSjvk5bETUw7HlHWUYaRbkG3zJ8w
03vDx90BH5R2nJRMzWC4Q60V/fcvVPzUGQste2I9xNTUPkpSe80R6Y3ydF1mtz9FrcHvyGctiXFz
F6Zml7Ozhm//wOOmyTwEhjvh784au3M+CdAEKjfWqrbpQhnQb0uFlpT1NJEE84w7Vi3+RC9PTxIw
M26HH+HJN/6vHBZpnPcIfqqJGMEY29y6QfAOqwV9MnN8XIWGJYDgVhrP2kMej26yd1QWX7sJrPWT
6B1WowjGS1Hv2UHZtbS2jjpP2RFODyWZ5JWzuiW2vXmg5e33fTlDwFgVfG3YFCg+q/WL4gcT2o9T
5l21YIwk84GMRbjiZSbfQoce6jPI8E9AvrpUeOahrJ5DH+AJqgVB5Rde7AaexF/ws39Ep3hH5tOv
FmXseZjHElBHQwQ7nbs1DqeS5auhsxMmvWp0CedPz+VLmG+pR0j1m7hZfGUHyrOFgGr3dRH91P1t
DTTf+XC7o0fjgdU+d9/cBbVnmWVGqaEzOrrz+M62wOUJ+E3NF8+MjBZJ3adPwCi8ZbH8V5bffMZK
PMvPGEnlVoQoKoPU9zYMLTA1fH3KN1nxBdlFFzf5TX+dUS4FQUSi9L31suQM0usnqD7E6ALnwG1g
TJi/IZ27obF2S5MczE1rPkatZ+3H0YRBFjqlA2QxpV4wNTb++3HCpaXIqunbHGSVCKuTD25JZ+4N
31fO4ivA3Ev9xXQYzxBEul9TZfOAceC1N0btDsENte6yQdprzoAVYOKFT0ZYVayKikg2P8B/X9tb
BcKU+HtqtPcplZT59bojqAT5w145chqmzC+GGztQxh+2x0tLdo7q2/tOcu9r89fXdOrnrVEZ4jdE
YQ2D4r0QnCuCkrIFqc3hYK2oa27HpT10ZIDHCa3PCcZ8qnBER3VLv/9KQlObPPDi9KZH3Gq1fOb3
NysPUS3GV7OvzJ38xYxPTFfXbdno6qwmEZZOPBf2eANWzggwVpkSAqU67pEwd24MBJc5SXR7ARz6
Z/elc4Wri8WtcauYtIh8/JWTRuG2GZEaYT9c/nnUD8Ez6+Q1YFfgSezxXhuWdDjDLfNjNSSo1m/x
OyFmUkVTRmfu8mo7OqgK1LBnJLfdYP+RIjVSVxyQoaUVYjgGDSaK9GuAptHALqlwlCFZ4mbDtVyK
ZBD9lAWiUpRHl1l5NZAr8cHcGqsZ3EeXrq2Kk/rBTbkm5OLxwyfjUVJtfLgZtqjyIyEg0tajDime
nRY8R4XcppHIGigaplJMUVbngIo3TDvmHWj2TpuNnsQMOXLdCMFazoz+V7lyzQyVSTcOS3trRn32
sdv3YZmflC05Q61cUeTTk38vcB0jtDo5Pzx0JkXo4G9VPIYfGwfNttBXopdCOhmLHJINdiZkr5sa
/fmgSazEwAJsysuF4ELJc1J5Ep5L5z3TIUo/szOQ1xAxfGIGB2RHYGi1Jc6vV+9yDTVV+HV5EmmM
YxlXn0tYyCohnrEOc/2Z9thwWVah3tyDuC0yIsb1DYargDAiY/B/BMoR9FX5XzT3YRwWEiCbKxm7
zndVIkvdiSmK1+4gSfEeir2kQz1GdXp2EzknfHJ9C8sXjUQaIHxhODwVCZKxKt5MAyuP1Cj2Ryq9
PmYqynh5Nx4HzsiJ711gaKjpQqEEZbOe87MHOUIhFlxzW/uysmGqDfvjDWoUI2knZHksG9HFMD+Z
y6BCEJrnZcwGo/9L/l2H9xXm/55wfOtrZhUchwGETpDhRuKoM7xB5MR8zaAYGktEzRfgv4wY5wlu
kiSvWhA3STef7Ybd+FCbzowNh4M629biFihEJJR63oKFzQy+7E5iqMd8zMyBW0C7mLBjaJDteK+p
cjnBxtwvYxm1QSH1OgXepJ6bbDOx3Fh+QRmVozNkOKq5QYTjg3YlxVSMAE27dTzW/7YpWIkdBo46
v0Ggf8SHC/vb0qXtLNILztshYg+P1F/UWz9+hm0txdQoe2NojL5UI79D4jiWEn9WFRQulXsp2XE7
78LQUy1UHksZQ9wiutsqGUX65+QlzEgFqkJpzkgcgNh4N32TqXLe37EZrYi6eWWvxocGK+2BzGw3
YW6MPQMNMN7qLIGrj7UhEiTi+KqHwfwufJ8kOmOFNKrL0BOUKlC3acuqWxkWkpWISH4UKnLYxMvb
ZvIMZ6SAnEDvHa04d5uKAd0nis9kVUNBXTcdnrEc+ABiUnGJvFy12VXY4UWmXwtgoce0BwMKErvm
T8MOL3PQ6gmuc1Khgi0h5Bf31Or7aidUfjzVpnVDpuGVwGR1ecLacGjaKvohSokiM9j6ze/cuexq
KD9PdGizINDDqqlbgWaIgC60uwAcMMJuWAHL0cU6WtXfDqBwUPEbkensasDADkuKSghwChv+YZvw
oV0Xbi9nqqKeVcc9wSeeoAxPUqOuWgAkYnYpuZk7SVppdOxOhezZXSvtnzsikT4PFFnoejCCEilK
VPUTv2w8CPe1/vUrBJw+Zin5ImI0XKz+G8pncv9Sl9Lf1e0Ik5w3bc2252i+ODH9b2st9xy3OLcy
5GwzZICTCyvvpNd6wK2gofGtb9uVvaVY6Im7gMS86RVg1pKXalojiv7Hk0HhP3/dWuXtw2cYeF81
JL7CxI3w0heUxZqiwuSjzJX5ssEbyqPOhAEaXBEjntkLAvkCwGwu9jztZjbjdtOO6o4OX1CJiVdu
fUmiUowZiEBKDLc7TP+mXXOXfqP6Pm+gpxRNJykSbMci8MQ9KZKFWKVAJtxuzHIaP3n/UZ7K4iO0
MLL22S/WpzCF5MZS2EgVhQ8oBf/Qo29g7T2sUysWt2mJue00DxxNybiQ/GoVhe3xON9oEQrEPbwX
N6xvwDvapYzFzUiAyDIcY9I/oxL9a7fR2qmSpnVdoWCfKa8fJ9IeQxQPHmBinsvJucBQJpkv1VqG
aNXZ14ZP9nwDzz73tzRoPOdVHWTyOaSlugygMc2/WdFfSQWbX3Rva34fX6sW7I9Gr5kRgk/iIoqC
Lq8TYnLUFR1eOSZrj3PVja+dLiDKIrENl8Vec+7ND6EUQOxtflyX+DiZheDaHyCSf6R88geLHwCT
q5jOLR8actZ4uxH1mc3D5J4y7Nxu6TpKIhi0Q17fKZhzBzPsrIPqfbGNrcvCvCnpmGg5B+mpU5IU
ZSQKkRhZok5DhrKgyJnGMTTTmQu5k/D8dS0vBkVQfl5pam82hKeuaI5S3oQHjjZHR+ZTbJ+X7wjB
XqCHW+syzFNZn+g6nSoy22jN5qACXw4qJIVH5anthV8quxf8Gx0tKDBV3V+i6ZA7svslvmUzDr3+
ARwYLhMLu8PRoC2Mvx6Ey/1aQ16NJaYzAhYKLz1ZPcOGC3DIPf0JfGPtYBwOsrpVDeo8iOk/o5Fd
aLsmIO9pAgoijcM9Dcb6fuHGPew2IuaWB57rNMdnolodfnwFZ4VCD1JvJL22z+ZeXdhi25WIvjci
1j/JvY+mJ79V1mZ7TVae3PPcPWW2O8kR6hpNwzsy/1QRCUBJ/069zCC/n3dQVdqzf07pZt+e/Fnc
GNukXhmp7rDk3TS2ofT5qS8CFDZxTKc4uSngSo27qEmqR6/kpH1GtbyUZm4faH33tl5rA1Ma3Qwg
S1z17Yp2DGbF+eiYIqancLS6CfjLyB/OyZ12zZOJiuF8yNPdE+h/L6tuQ87O67/LXa/ND/a4bfOR
6rbEKdzKhvv0918VcVGQXwEvkfV2vrf9H+U/bUoeuSmPVEkdaFi5ViWJ9mGtxRj48AjPqRvlSNSq
AoB91iIitxexkA9MdAxJGtMUWKMvvTNhk6eQXWPIaf7seHu8HxLFAlk9rai2HbEjotaoGKTxFh1+
V7yMqtKrTgNmLiEKj6tQ8Ucr/rFwl6gPxmtEdhtRnr+RHB5uKcY0JAI7r5fvZ2x0z/qLWiRskwX+
tKGQrBw7BiAmVOPWEKovGOTLS2V+hxWIIlZOQ8w9McEbErqG8UQ0KuzUl/mk8oCbbNtKtrHDBCXE
VtVSkhrkmXCbibsHjmwujWx4f19uRF67OUEYIqeqhXdQ0ZmzqNvpAG3CVcDKnKxecW3rJTBAg33z
eaZP6cjKMwmDvXnQejLqAzC7tz7IF6ZYkW/UdvfJ70Me/7vKQfiGRSKBvbvQd/IhajBCK0T1qM59
U6vfarpHIc0pfTAmyrRmtpZDfWfhhGdWQKKfajymYj2opmGJWY2BRmGViuG5IlImEW94STpoY+Zl
pZRKzm/7jnm0QaEdhAk3s42CIjO2ylqrgTbHH4hxBwoANy5e5x6Ogr/c+pe+iBkufjAXiZgmGmMu
7cE37JIg+sY8HcmlbTAeCz6UcAjp3xb5RU75yTJWWvbSwBeIZXygeQ7G64cNi6b73063cUSkX5fG
HjgI2ujuHKrwKyYewLaAc/CsHhyHDobJRjo3aq70RwZmSBhvBADDUiBZck3mA4aPmqjkgZeBEPhs
7VUJjXAwYEB2DVgEcgi4EjdzEGm6Rmm56r7D/fuzaPGwY6A2YpXncW1mPIe0sEmdJywgXY519ZR7
+spC3Hh56dR+wtqOszYa87PW5ii6FzuLFSJ86k18/LIqv4h4uZ3j2gG6ZabfQqEPN9e8AleLMiD5
pzh9dZVhe+IAmYRRaqVGN59M/7oHmasjigNN3NRjkKC43+yel7TB041OrIDyNbgY7sgC/hkwkCnY
Ku0I/rCRUiK4awS3H+/T7Lvmo3CVKcArUefbaj4/NN3ZpCpDAxCZhOoQSqlS7eA8MmlJy8DfI+rc
DWKocQvsyA3GAIRpsZbcgf1pvxjQIWWmuYDm6Try1xbJ7MpEEr+eD+ZSZZX4A6VnYZ4RD79qaxkm
ef6Vn7/46VwqZ3pDX32i/AeGApHE13lfMceOJFd55H42hOt3dwE9SU9qrhHOss9oYSSYaiMwR2+Q
MYAsSYnqOtDDF4dc4f8fTswnPpdxHT9+KYKwqqjIs34yZSCFgeOm9DWL5NKFnYsOXpj2px9+XSaq
4OlqlpKgNCG+cOJDSgI9M8K9/DNDCOCYpg5IGyslljlDwk0ounkCmSja96+b4wImonc7/4me0Zhy
zbmRUnOeeY0XxqfiRiqa3grzKn6YOKXBOUxadZ3xlBA5oNV1aV/rcG1paHWvjAeXg/LdCpvoXZvZ
S/IAnTqw4On1o7AWqDr9UNJLyQs+EY6S+UkyjzvuNRMRGeBQjUUBZy84WetaBx9ewed2dgWu6MJU
xL8rfi8hfLDnFtOPD7Hf0SSUgKn0mhzFXWhs0AiOzRAKsBvJINjQGvTX8uVahcbZCMl97cSpr1L9
tZ4ykHZW0yNDcHrcc4wjUr1/94sxQzj3Y5366NzLvhUJXB9ltFBZBrFfdhMtcYlrZvJ0BcZ7x8MK
o9i93xGdBi01vPLEp0qPTPht6ql8YLfk+ZaACr9bA+KC71hTcKFC9VJOblFDKUAIQ+ebqzD9bMv6
VZBxvgm1OWFCnN4ob68edl5NKbvZeXuKAajalk4lhfUABi9ts8WsXSPMJOmhhwEyZ2NAuPS8rqsU
eE2DWddZBxzmUPmTyZz1V61NlvUlatqzmeBwEIIXqEAKo79M9It0qcxC/Gm3f0dTj8V9teUcYHp1
fL2a7sweuMCiC6Zu/4UNYpmfUveFTAzDL3mQz6FFHdtUpf+x8zz9MOoLSHAl5XG21cU8qpd54BHW
q2/pbRnYtGJcQZUUSVhrNUO3OePbA9ixRtF5SJyyIqKVTp9UpcEvh8O851hiVrkL+GzFfg7w4zeG
IkDRtZlOSP0qo4evMNBk7tu/u+ZiBTAaM+jy4CTi7bolQHA8LXZGE/88vrnIfNoTaqLaSxWBuUuv
qdPVIgFC1coDV2AEk2Sc55+zns/5NtsHjvo547S6EO+tG+TsfDVFhmE8An+dPD5Y8EciAiXzPhUT
l7kHX70ehKSXMfG5dnCv++yQoUDPGHUYP+ou5lfOsrcyasQKgZgJjwvpIMdZccls2S6r7M1a3HTV
55rPPZZRlIccVBefdldMJFpg+/FGGMAraYXTQKO4/b5/nGcZh+hVg5iOSchTJ1VltWSq4kxKn46E
fTPLpHZo8lilYFoDH2eo/6Mcr8rPi/7+8VSlP6fqSheRAsGUiWAqmQFTmi61moQWrRgxYXTEiQz3
FeIUyyBBUMoGF2xIOIHKSzVToYfxOF7dRjcEwxXWsxzVqclFmN4PcNMKAtkUjUGB00Wg0lxq/sNS
PKuyxwmWDGhdcwgcND3x9BlwTv/IlJU0oJmdCYOAscTeF+PteWRv02hKWn40+SBLNVbL+4NgYdG/
sRzijb1MqjtR0Ed3FqGcS/ytdG1Jhb1l47H/jMoU7CkXXNX1cmgrQfEYmIXHlPYsDMSy1C3lDYIf
PzEhGNodvy97uh/Z7fRshxuJjYOWrE7guDykSlk64Otw1y3Cg4RmHwEVwLhdS6fl+8WTARuyXhMn
oqAQdfIFxB+lZl6R4T7L+SNWr64NBghgF/oYC0wk7YPwSuDwa0mOc+RDoMsLC39vNVgNETNNw/sP
QLkRktOHrSFDLK5rtVIAonNYNnkLUsEZ6IbcPnzdkkE/8YddaSm6LtxCN6y0icUYabjV5LoSyblv
3Ma9uvjm0CYbWkIjC1BasusaZa/C4vfEVEjNa5YiF6NiReIv2S4fxXEwiyG/V5GV+GKMz4Tq+LCk
QTQjJAuZmpwBfbr+urjSG+H5soCAhi6A8MKYyW0coD5jNnNWBpLN9KC/1N6A8R+oGvjJRs23/Rt0
/8PeUsqBu20Bkbf+4Xzsdn0+ooqonUGUJINjSZqHvdFmIfcFBOJta3h3GR0p1/fn6oat66ylPj1I
J5FOZybphg4Nkr8lrqkXMIWjtFZr2e8CNOebnxQlUvG+prm4sfHVds98JVPHd6zWQ/y0SRgGI8bl
KhS8hNdWyE1rZ2s8L71lgB5VNTZ6QqqvuAv4M6l0bttPSjWqP4BvIlwBDbijfRCspXOP97gAHMkM
CYEIyOurTpjUmN6pYeZNEkulInSqsKwYuibqW2xivyXUDLVAIxmj45pL2lIzNbfpSGxKkJHsgZS7
zv8yLxLBjwhMTKIavF3BiLsq7x9w6PCRF7J+U6MLx+n7J83BDXiIEWaPqySlqncAC4JGdB5WZ/IR
yda9aMyLRHrILWwQXjZ6WtPGaPURGfI8uVqVuzjoPdBBHjL9gWrpoovoBZsFiQEUtHsztpGUPLrQ
03KjxEabofpwbWV6bN4w+nurMyuGXfZqpt52xstbc6IwrkczAMGpHZdkXJEWIS1k9EZMqJChvTeg
Q6QSy14PQUlkIjn6Cl6aYv5/y20yYMfIO+z9M3y+DJo5qnBUlL9Ilnf3D83XRfFP9XqcRGcA5b/Q
LMeBt1rLnZy8boRAB7yzd8ow+kdc2KKn+hz2Jm7zTcuqZZAAwQlyMWybhKK1SQiori3b6lkgbrz7
0gvxHtzVLengq9wkpuK7xfG1hlWv9ztlJjVK1to85qe4t2VUUCugV5h3Op+2iDsEEY2l6GxLX767
057KmoVUwPa37ieobSYOWFIfY2OnXs6bGpqHMYLbSJLxkhm72N1e0nRBLB0zVFpo2W/2VqdM7LzU
kaaPZm7JsYf7nkRmqAjJj3DEccjs97qoIbnYpZ/d3T/+704JW+2dZl6Jw3N9HERV0DWA18kEt2CF
I3YzTilaoyDY8fIEZZ+ycTUQm6dzS/BIZABdbIPNus1HJnW7XGTB7OqZ1Hj4eNuYMyejIUpNfJE4
wyw79NORkbSq2wLSvkQfQ8KamHum1k78eyxh214KzhXJBd1lp1UjuXUYhbf17QokKtIECbU3pe7L
dddghN+QPeb4QRpe2GxuvbTsNH1tSBqOM0L0lvTa2tEEZxiki8BbhM4ZabB6ApfL9qGpP4KltSBH
jbkkN43x51PuCKuzvVUjneILvkJ3EY8IEmV8b7g87CnnM4yhKmDl3Dk91yOm4/lkqEPuPiZET7Y1
LSMsrUqaOzJtjRWuprZKnyIDTQjnS7uHuCnvuww6UVHfngeGUGhOYLg2H/3cLN+FUpE5tcCnpELf
gySrBYf+BhHhCwOEMhgMaf0LFMNq7lD5R/AUBCmzAT6HlMO4jKFTEGNFLtD0K4hGy2h5aVVVczTB
nL+b+u74fiDGybaaOGbCeZgQzpOqnNh0w9tjcrVv4xgN7fAcN5fns7QI8Jnrp1aumi7v1psBj4cN
Vnhu92KUHM9BbDIU1Kxmc+fOSmoNZ5Onnkm74pLWZI1Lh4W3j+G7UIcENcmJFWgcN2Donr1GB+nm
hVYTFl/lhNjyFO8Yz6csrDOhubWpfguJgMjkfAnwH/LmW5WnnRlbIkf/mCRHDayY0M2NxHL0Ti4c
QjB7IJAZitdak1qnpa+K361IQZNzZqTCN7WseWYa+ci5ukOk5m5EuExseBwrj4XEUQN1BlLFrVlM
jljoLzvSPXUbNfjfjvNxLwnOchl2sgzPJSeB0t66xbFp0FnF6kSaB5bXzgTEnoQ2qDq08GHP6Bfk
n5YtOkpWFfk/fdiK+TK4m4k3KjC/LNqX6bKzsHEYYq5g3efE6rdgPaSsdxtRi0sv8u+BBvtRBzjj
J7kpfIXiExZ3lPk/6CVbMqn+DAzhn7wI/2/CgUQ77rUKnxrXwcRMHD4pR0+9rDSZhrT6J6Tihu7D
StrS3ZiABwEPwCOgiHyOzPRhYZ3aGNA13p3zkxPWD1ntoI6fj0kjzpHAqxwrqHFuWuHfj3XUnUfH
zAocdwHyau69LQLkPIXCozlSfEXEDR/pc+ID17wVHOzmJS82pmvhgfCsJFGtQtCIgk2GJET9lO1u
7YDxIYab8Lxu1dMfssX0qvokle4gVcGwqhpBWgqghzpW4RsPxT1jshSDTziv/QqB83soGTcxHlwo
TrxWphC3RwbUCVbR8tS6C+6/PPNZqIHuNlZqitdfP0wJF7YXxeNdv+esznaa62DrZCmiuecyNbR4
n7uU0r5R/0a1Jjvz1kuPR1w4q7blVwYbk2s5IjA7Wkj+sPCpBXoj6EZ81YHbJeccevfKq+UmRDDE
5HhPadd8aGZpc1WCUQ0vgKcQaScE0Ph8ouCxYUsygfmMhT9bLAd7I39R3OZelaxQDGubfg/wq+xC
wp+hzVqPvOcocRh2pM3/ojOeyCdCSbC3cZjh3PYGrqBEXhEz8ZBwiPoQDxzpAxLWVM/8GDaBInaO
iUco0gGClThxrjtbe5Hvfolj6qALXPEU9P9ie9PLzFav9nYp0Qcc9Q8ELZygdkyQOVvzqSCAIS1M
zqGDGLipWGY1nYXJeAgoMdjJ9tIEAennO6NeuMQd4pz9C0XJ2Vkv23da0Pmgt3Jxh+ZoJ0RcXSef
21O8Ve3XjxEAc0IChDOJqTNKcRD8TSyZwVZJrw3EI3GeHSUrjbyJaFtaLBtO30EnD+dF9KZ7oAsV
cjP8vq/Ef3HKu5zuiShu37RInmlGGkU9JgmDbxQMOAduLu4iwRDEfUSDBOfiVgZFmDV3dS7ssmoD
BT6ZNGWkJ5KDZUift10wtjUU51prkcM1XgPNnSO6Txx5B9ehxUaCDutBxe99N5JvuU+0IylvOQDw
AqYEGvMp3SA7H9G7ir9NB1pB0LOKBqZcXrUrul7oRqMNEifxO5AVTMTYdSf19qErZUb1EZQ5VHjM
2xeOPdKSSavcyOWRT0fqxnkMBoU8dzSnk/LHlIdKL1fdp3s3g87i1MKCgtmK8w72C92GCKxEWJuq
/iN1bzznvtPUvXqdOUVmqeUGSPpT7ETey8pOcc7dYlm5XGV/KSo8nMmxa4wczAJoHMhouhPVRfPU
chnKO+CElcGbM52QsK4px5aC1PAKY8nEEtosP1TmbEaiQiDr5azfBOR9ubXY3GMn3bZyLewNHYS0
aaUGR0HHQGQBvU8tb+hW7faHAqiQwu/ypbH0VTkoGapwa93VItqs56zaTVQhMVydF9e7X5pJ5SQ8
s96ZLX+1dYnRqdqgjoxcwWiHrEU3DzJEN5lsNKo22ilq/bQXlSv898BE9eE99QiVQhAmp78Jg2yn
x49hzUiOBgj2LVsCWO1msrGSpBSbuJ6IZF7hsKbYptflsZd99kBnKxclK/j69ZNW5eWD3zVfcVr4
//GGgTcPSxou3lp98PdCTy40mFUnuwbLgGHU++uRcDow+7COrCT4X10+esWgtD7c9SkG2sHpCrPA
jRkhFcpmJigSmdGptwO4A1onUOZX4jOwDKfyTUzt07IHJG3O73OUa1fO8wszbF9MSkZ5qC6ketrD
foWYXZ7m2jcrPMYdbqlO7DHph+9RHAy5kbJYNtr1cJXi8DUETE9GYgAxVzA5XESiGjNWhXvDwE9p
VvvrKMBG3nf4YtrPoB+KuUsaKf/Sa1xkRH/rMCxc4fKGV6tIZZZM5pfotmLgnrBQJUG648gcYTVa
ZWkcuWKh60uOwbopbLfYVjdw8Gi+N5kEQMVjoHA1cygKam+Hfxh3xG5Mdsw+nvEK/VCu0urhWJGb
W8+y6G5RaBDgS+fI+jaKVMhqabrjZohxyAt6SmGV2Q6E7djMR9H3UyIHpfAXdgdTTsqy9VI9P8t6
5eJo5tFu04KeSyHA9dA05JEWSyF524ZDF53mbNnFSVo9s2EY/UtxFNlu3tiJ2aqKGSdP6Eed63uc
1bmqd2BvMRPYkDqfZPnLjtsJPXZ+A6N/5ARcsVTntpH3X8pFNQqkPPprGeV3Wv/9fyXhi6x5Rohx
VJCGBgRTJuU9ECCmft+izkEkCcsNROql0oHxAdUg1NxePio4LdUWvlRaLbE39I4RdY9TTDo8BpVq
39ONisTAcabfczGBnBG0MnY8RRmxPZWi9fKyObda+v8I/lNzUWi/BMyEKSR2J2/ELuVLr90K3/+h
W2pL8nAvo9Lh2ENHLdo5PNqzn4GD+3mBqCeegW6qUhiGAvbhV9c0d0aYUwOBhV2OgA09FbcE1oWl
DKbLJ+icKx1gQMD2EqBgXfnux3jpbRK/J9bZ6WPPmJziot5/KT7CPFHdlG7eToTZ8sjZQmIc8bUT
Rmv92PgV6wbLHR+12CXU4K6LTfiv2qTepuUsRtYyxAxbRMYV+/vUYh39Xw+U7SHt8g9XB4UQSkpu
P2ZtGnNdhdfB40Ow8ep7JfFj56/l+X7eLhlwU/4ExG+oFOZY9Cx7smSrSIp/aSs1A7WY/m/l618O
cbbexXBmWw44ocM0s0rVjHCOGHBY57oheJfwN1qrZXPmLAX3ZDpaA2vlojvwTJ3j0nTLeiqNpxU7
W6uZuTbu/duE/jmvDGDj4KiXlF3W2o7XVgeDuZ/esa6uu5coubMxC4Z7EArr2KFMHb+WLJMmHeZ7
5wwM/ivEWvxAwEK7/yYZM4AGPbdPI8QWnxKWmaL1io/6Z4EpsKMJVTaWxoWMfz9nu0Dyoof4v93f
IkPz7u2gn52Y0xDvQW20b87xSNwqtE1oGBCPP8nbHtUNBfsRyiAoSAFSWiRe/FeChn4oOjCDJ0m3
AEHebB6SB3sf/bIukAD/B9INspUgFRdJ8Q0HI6zhe07wIVcBMY6aTVFDQkrlrmo1DBObAYV2UUp1
hJs4BVO2AArb243cmRZ8EEDqI5gwbcWJd/qxk1kwzGr1RTjMdwS7dWnmu3NxmV51uTEi6lBOhCL6
hcO4up7B34w0d43TagwujoB1OkXwiF+LGhMNw4Wa41K8ydHLU/fraVjARfyBFIo1tFbcm74WAS1L
b32UKdhbY+DxPRzxB71Mj+FZP2gGRw/h+RMPqQPCJ740WT26jUdXGl9L9wcNs0Gx5J4u60TSwgBB
qI/PkTRW044Yt00llHNLNsYjmGVYOEbQ0BFkGMMqhJ/iuPhO5jv5MMv7bh7tKkMjZ0eg2ejBvT7B
I1hAeTp9vLRuJlaewu61uKtqV/VwLuorY3e4oQzh21zTg83oeAo2ng5ElSXTpfeflOEy6zluQBiD
BMx5yIisu72v4ROrz9/C2K1vKOMDcrGiRnaAwRqBXEPMFCBESPddtU12HKINZLRyij+vOZmSCBWa
5a3RqpFLSFYWXNueitKAbX1NUcwtdN7RHugqFpKO4q+YW7oGs1BvTOQKjVdDCDpZe7w8PG9rVCXD
Zol1l/HyEWeIBZVSUUfOfJqwG+hYwwdXfFJBq5vnEv6s+V8NHjt4MaIU179RTDwt0+o4y18/FoEp
bLd0TBx/MKlYn/tboVjVURlGHoWAR6rbZUX+vz4b669aAQWLpxRGjzqn4+4QlSgi9vqYKPfBueiP
Nln8kOE5po+LZh7goNaxNkQG3p0OfFayxvhnrFjeVqJlA3j2qk0FIXW7ApBQETU05SipnkMF+LBv
Pu41CoZek72TMt19uZ6bs7mPP4Xz0xsMzNdXphq+HFX8ChOMtOApG+6PVA37kV5Fbaego7asJC/T
O/uP0Fz00pSXbsgE1vG2bNqCeHwC6Qwpq+mja0EpVU4B+t/OVNJ0LcA39aG4AHtaNqjzOYTAUtIf
w1gpDKUKO6OWEfKuD+vUMO0SHd5NTNN0mfLhc7OZv34sWigBhpQc5CX9Pn4rl59fKwkB+FnvqJsn
OYglhQHsidhFQBDU67rcjRJcZyQyAVqWvtc+7hZNXsm5/mieUB53RWhsXR7oDboBCaSPylBSkLdT
isvWPoro8uwFHF51pu0TyavmnLKZoPhZinOSm0CQ6Xigko5UnVqvXYTGU/mLrgrvKIWJ4fTHkb5T
ZivpwMObDmAh/hQjD/qpxM8Y5Pm/AKcJXR/V7PkHwEpV54Qbhle4ieFvvPTwctPtr8AozJUfHist
9FxdvBaZQT85TURxwH+h9n25GxksZbg7GvcZiMj4OOk/KBV2lFoI8LUHRhMb2+Ru4xK/PCw1LO1D
uX6sK6fvIm/RcXIXYuP1SZmR2HaDc4cHlGT1NXRh6IH/BrkGyAhbcApoNkJf/O6y1ziKDoMCeBeE
gDP8uvOZln2SOH4YvqGoEj+nuuZswKwMWJJPDiLy5022B/HraEHrDeU91YD59cGillImdg87YWvu
QJMYJJLnTqrp1x09R94r72bfn4udOaBSqZx7Orl4dylstJb0BojBp4eJOxQ5prbXMvYm7Tr8zhz0
tLwGDEzxHmTqghz2IwQ7jsC0sfNqgEXdNvupkijqfK72JM+2GkdnlwhoLZGZSimXGn10dLt/AwF6
R5kc0g2p5Jz82X/VDbVPBt8ftYbvGjEC+yHy5nj+OoXWyj7yrisS4+bDV2yeGYaweV9j0iz8I+yR
G1BivFTehxELvIX5E6dPqHTfsRGugxnXK3CqGl2t/KSPpX48U7XKWJ6/ZRxeFiIR4mUywTet8jFx
WeLyw4GaYudk3Isn5AmUpOPKZF2nqbyUHuF7Cca8dmPYecuakIvv+zh+lZ/qqjdYGOBl7M+GKsxu
r/XW1O/f/p1WUsx5K1TDOCfpw+F8T7SNQa33SPskbDv8oaof1l70jtcolTkuolKyrLoU/Og6UAUh
eXsT98HgNCrrlxeyma/oWt2EKy0BT8ia0VHaaivHwfRfbma4BYCCl1359oD4NETrrs+cES8H89hc
jUPtwda01fgpMMccr4Z7Eg+dMR2xfc5cLbgGlNTFxNAVpl0gFwCMi0WNB+TQSAkSj3EPl3Ism6Lz
Hx2pcgELc3aEqrDZNKhr0yfbujEcZq25f7qhy52t0poLnbIkOrl/F74Gk39xRuMiO4mWAmvK+cqW
AfVC/4fFPzRYnoL1pYqgR5HMVv+pIoR+AeUCTsxs0LecvJBC5234Jpyt02RNtYddKKC61aXC3hhK
OPNuR+xvcXxoPICC1sPRRiSVsPJieNVfunZcn02XpZ/7BZaiVjlx8TR4wfJUr79jBfjE6tOec9L2
zLoHxzpsexfJXjRIRQhQAiumGCxZWriuLGrlbEZymmMFAx/UPsFqGDmV36N1A36sOAJMf9cPfeBU
OuOVAtYfUogvDuVlimuGVncZu7XsD75SbWCH4DeovCxfEMB8fehiII9/rbNxbxkO4TfeMGL4clt5
fDlNgJKM8OPovjKcf3EJKwMUBYQef3b3b5kaBpUrvnC66qtnmth/vxiEqWnO40X9P2DnkywX1FGD
yHTrbubt30tsEGz+J2czFpPCOtEG/+TxVFQe+6fz9IW92cQvOnMdBKzKethXqdKNvVJh8PPJ0ALc
vW5zvMdurncnQ0nqx8sjEunAOva01SvOtRLjlJVeQQyt6yw3maD3SGuHPvX9hv3fq4vnc6LrfHAt
JzmHIVPPvtmKM/mg47EVICmAR94jSF2RQ3yO9Baq0GxPkBjERNS0OmzIvr9j2xh0bGcDWE3kl8sr
5oy7xnuv2PZX8aQMMIHe/rnnixUrRkH2DOAS8rJyfb43dIofikK+PsuvdCZ0Kq9cwFOc8h53gtNw
EQwW5JRXdeIzPiMeot/zTj/BoGQ2xvlJD0hpWwO4x0qMGcFvYUcpIIWpfq93Q9+0UdaoRUgjmiNP
imdScXeIpUTX+7fspAJNbI2QFiAdKk2GbI/wwRRsvPlWCFRxv7xETU421eOs6ikT1/+EIURwYcsY
3Zo1p8fsv+hTfkvOtpNOI+vv5WqUHGorfzrGZ5HSCnSlxOJnft84038bJqIyed3SoGkv9f9NeS4z
GMJdUBRUmYQcMIoOgPBuhmvZgJhsg6cGI0BFvuPbdEh1xFBEOt4ZJcFqA7WW8GROLSB6aIVHUvD/
+Lqr8OYXJfpVB2Hwry7yBBf8g7MlAs0ztg1UC4lo1WjmIh+OvDC72GAU980jsprvO4h3oTIQjwgt
S8S3rHagqckGqZJPQAf8x2p1zxU900Y3a8xp36oRRY44eUFA4UX9yNHPhGIy5NNMgw1BPZgqRQG5
u510wK0xsB+Njh6gcswz+kw9YzdXrFT21dvT05TmMHHoHvdUUPPpDzHTUXLzo6n7Z3AH9uL6MuaY
dQzKm3p/jy1/OSH5vmGgjphF2COFjo62kfZE0KVIby+zr4QjF625148bZW6gcqhykzTw8T/SMaTX
lzkbqYKb8fMu+PP3ssiX4TJfQDOIE6ugiYb3+3jlabUa2q8IcJSl8KqBeGeeaBtPlwtF1W1K1cPl
b8j5qb1WMRHRPj7R41L8J83/xa3HhLnhBXBu8v5kIczdLrzrMDXXFcf5HPLxVacOybJeiiz/YowM
Z/gfmDKm4YUDSbFgmqOX1+n+MgGsUP7l9j4P/Dm/EN4HMLwwWWzyCrTsYVulYuLmEM6t7CkYGHYb
vX3ldFUZQx/pqun5S8y3Xpz3tUewq4if0lEa9UGlGy478nzpvQplDXLQNJGLNgeNwpcyths3AZj1
wnpyMHsTLyLgxjK3HTALspBPRL+LBhdKzaI8yLoVmhgOwj9SObx7INoB6PMMCNvX9sHosbiA4B7z
KWiYdofENo5Y759WMWgobZDDRh0TKfy3E1EBs/5Qb8vBXp0L6kHOqn1gaj3yxGZNfSwY+1DuNXPU
e0FaHIfmCUYVPvgKjMKy9C3Z1KYKLsNbmXFSAaeDpTE4muNO+TjlIJWnMlV2RA26VWiclCvQSN+N
4VpjW9VmizBB9ITHIdsOEEbSp3/mOWlHofG7W4qzwuzNmhseRnQAGeCsj94ogh8hRcn3fmOgIYEj
O6eFylDW/ooeqOfzrNoOrrUZGWawLklTdJ2x/L8avMLED6cwD1ZCq2HE8HcH4OVKr+sqHNTyB+wM
VV4NoKMgDuRo/oD4/U9ByA3d8pzP/XRe2z1uzcc4/WoPhIDPnhnm72w5dkzuBpxUd7g8SRznPg1M
anlFz6hdW4NdBHh7QcjVr7Mi2grA0EC6dpOuij8EnOKKZY3cg3HECliFcd8M1mpG7GYxWigX/SOw
UG6xtQ1CkShCu2j0qcEcQBavaV6HOQaq9mIoLFZgyelIIvL+QkaaW4dtTjY1TjukjDX3t8olgdO9
5nabMmkewsqx7Bgy4S6khZ+d2MvwBCoN/SHNHgPexYQ9OlCPtSWFjm00NyUssdGS6c/yi1o3kvJR
7Xl+pin9QeCPpOrzrY60LitkZqeoLzJqiFnvUQBF6EpTpdWE/+J5sMCJSVJMjCPGdVABczlkyFLN
w+ZQ5eGXwcihitGzAzXIKt0zV/sRCApvaRRJS/ySTLf1cBtDp4ae6ddI0Jxf2DnLndjGnUk5vXwl
Ybp3PoN/oCsgOviVuOI5E2RwXJPAbGv8VM4tDRKNtnrKLCK2yCrQRj/86DdC6jhdV6gFCOtqId2D
iVfz66U5cdGXoRPK95A5xnLlcLmUXs29lzDn9cpaGKDC4sUe4tiOeNg2Xb4x6WPRs8ZO/gXakeNi
gq4YzgxZG+RuHegeARMyUSqX+of0khqcDbMJihEUtP8rFxJC9kcaLr+G3QIUo8Pz10RySVXwjHmW
J5O7m5sJxBBt7PLmKYeBInEpIhiqMD7mboUBcXWlpNHEBVWfxkqHHFA8sqNamsmDGUNw8xKAVTgU
NKGruQ453QEyme65kyAMcEDkqfJzGXj9FKBNofRx8wSUu446L2tqfhTtl8Swp92s28M8KsWzkGD8
4IiSMQtgi01ZyIk9hGQML01CbQJ3csA2oAhBfvasUJG30SBSLbhmjJm4RoScLSymzS7U+u0yedGL
bc2tCTvaqxAW5kXd8QAzTPDIxb3dke1K8E/xMMS8s1XjBWT0stNzXviau/Lrxs/o8PMxIi5RXjpu
lDW2WG/YSPmknD3Xu5pGqakyedeNJdnh9/HxsPHSIqful85EqzJcFwRElm9geeicE7PY2zbT2LYc
hViXAGa6Cu1oGDBgec0mqFa1/Twkkf7DPyl48KA5/pVxEvymjiHiT6wKCe816blG25pTHJnJrj4J
ejD1Kqae3vj0DW2c0GIC91iCVR73Tf52yOGU5UDHPa757BG7T1ImWa+nJXIWN5847SsQc2yhTMvU
PPsJXzrhdfJEYK073CpB9PUyfNx+i30XSF0JwPt+zahZalO6G8pmAIS656DMI7ceejKGpgRSgSXp
EHGmpvUAxOIpgbanXVvOvHvM52hElACJT813ArRc9RNdIbqPgGZ1u16ESQZ57Hq2ICHvQZm3LLzO
Goy0vKEyC/FAJvbA0kAUff1w4Rm6//H7aQ78/dfCTXWYTgsyEqrZ5YmP19r7Ee5iHEXHOmow+L5X
aefi/F8f63H9uViXq2PFxwfRg8utaQFwLLWaDriQoI5xCrIwYK4RBAA/z7DgPt8ADTAJ++3LPDLy
CKLId+f0R7wadU2aim9yrh/UPckiQwyRIC0EWOfzKJtZR7CKK10Xy7oEKWnILUlsdQBlf5Cg7GGC
54HDijI4n5RJJofZ3fV14GA1VLd1U2BTBgjeaNi5upFaws8isomB4N9OG+0+kw9zMgipIBkh5Qix
DXKNN0I8yoM23Eul6/KOhkeLfBw7WCNi/wl2vd6aTqoAn3dYfRMWw6HcS85yct5DTXWeJV6aLvn4
AAsg3a6Q/C1S+14MudtK2BujlliFd4aKO0VR+Rm0lsTv0wSQUwl8s+uoMQZp5oatlR7x8e9fNnXJ
wPtDLtRdCZm9koNjS8NtGSxgmSnp+p88SVwZENaG+3qTYQIi/cLWeEaGZ00y2poIfhAiboPr24ep
XZ1bg+ElCEktEEX8xVHYG8b/pSc8m5fB1eu/zA963J0WODFrkqAlsonEWHsLe8ji40hWai0X+5Lw
vgP6u/GtP/+JkvAmhzMpbU/sA88PwqBbcFjo0CQ31XCCdSY+7u257+C1fSLb9Y5pv+OBFJGNkrl3
8zZSWP0+DJbjSuajpsAiSbjfIWJhKrxmz0bJPUOfYpTIbu3wqPKXZdOaSnYTM9g31rzqj3OK/BeR
PIsGRfJrvsGaEMUqJHs1auFrlv8eOFD6KkmMzKSGJEKa/jW+sL+b7k5zziCSCY9rHyQNU2XqgeLf
oaANlYxjDxoEPaovt/oANYOFHDYbZ3Q1y4ittn90hbdfaglKvvJWIMMUAk0IidcDxQ7fHX+NumpV
eQdgLOmkET3o4X7LGpCdIXNBen693nGJPRDjhyF2AYE/33/55q9K2AImr0ciBb2P6VGjRNglRt08
3i9pFGmj1J4eQVZJ4E6SgEHBHDH328dV903yrUW6qd4pytV3/XwJ3U7eq2EybNOY7iZns8/mWhdO
EOYDx++06FzCPDb6zyfjprsLCE871Id0p6RIhbkcyqMk6lQClozZGvXvw8LJf3xCg22tf17FY2pZ
4Zswc0NwesARqw6SG8thPR8zsC3/JkqTsIM8InIfhHsm6iS4A0S6mhviP7CoHocQdduoE/fnNcl1
41WeHw/GAzrvEnKSymkQ+3tI+Bg44THuZ38n7WimWl1EXdKN66fMs1aC1rDSj8hNuKCCYoFfexqw
tlhdCtwf293pHMK83nqgxdvyPnanJXWSfWedZIIg68Il5qzGmUBad/e85pXLrgIDIB6Km9cHoI1F
wmQD06hYtEwKEwI7IXz1XHhVvhMhYX+SXdUAj0mfYZxlvnLqOp0TsYRKe2v/LPzZ6Orrmrl1IUW9
MFvMmk/tafDbFDqsneRYJp2WLmBBvV+ngee1ARk800DLWZFYTuryh+S1rBmriOJKSSe2iMwZ9mbq
5h9XSrnpDw755REE3z1089XVJeMn74khSBoUddMDCTkl0gqlpVV8UdTq7DE9Hmsd5P77ynuAwL22
7GQSHRtjXUOPg8kjJRYnSRrJMlsgybqlULCJG9s5k3t1sZSUabCBXugnsT1D77xbj1u/v18iCW11
5HPEowuwErlUnODmdU0cBzh/DUZUwlPIug0i0nf+POibNE43ENKl7EUBJL/KtDCqcXd2kTXmf1TS
NWjFixY132bU7ttOiqi5XP5DTCzlLk3363nZoVhRmR1RDplaPT2m/YVS/mQ85KzdjP988OXZi2jt
hJnne5MIpyQc/aBZubbRAWAWv3Vy+eSuo1eq8QxnekEE1X9DWPaVohRqOEjAYpVU+QuvHjMbz0Ox
9CobUEQlX0Q4Bvvuxcmpk43lCTsKpBBtD+oTlG2BsJFgDD3KGyvg9nWtgyIp/jwTKtFr3DkjCu3Z
1whFCQrgbIboHUBtWwNJLs2goubs1obzUANEm432mt2h8t/UTSceF98F/li17rJSwQChesu28ZMR
QkDJR/3DTpfegn+ui+d/2ynOp5IPJ4E+xJXFTTKbRwozFTCbqdPpfHztAWgu7lSITrzn/Xb3fSJf
+OKf1Ep7KJ9blfHUU3sSdXo5W0KX7EuvUzsTrOZf2B3Ils5pCJ26S04U1yD542tpmCSt6wJh9ahn
dR+/KG4PmXCpi/+sbvCSlE1g5JBxeVr1TPPzIUHzrWwYA4yul4kCvTwvIHKSGGlOgZ9bm3Fs85Jj
uHV4Q61pY25fisKrZXxWNO6Qq0AJ7dg+EVxS6gamZ9fQc/MWsN2quwRABdYTUi7EFnmZq62mqsxz
1MvjspEyU6PigRh5nOMyE0F4iyCdTgqSHz5Pvj0pHTYXkm2ref/WUnRCJzABuVnUHdqtVfXinCxd
AXdBkNG5/DKkjGnBgl6G6PAwca3B4kPN46TIoE2eJGz9ALKfoz8MyWx2KAypwouvG++JXbb7he40
rNC6qt5Zb0ZVH7FbsROZAhW7KhYh/yrB3b9XKVsZ1afCBWc1v/SfwAP0ptajW2kM8XGROCEUjXpI
qqMsyM5mAq6/sPu/bpvhkLnu/06LlISpHtkDOjQ+08fvrCXkvwFfN0C5eKgU88PHw6ZyxDMWOFvi
SV94rI3R6mk32l5PUPBPLXuXXhGSMHGMjxrirvnOtFWxjbh9Ffns9W5gYXeirg/f5VSb07rZKJJt
FWK630dzXzuj3UMYPXOPu/gAMncZyBgAGozoQlpvHU3w6dL+71MXPpz6TVBlxxS40UG8pAt6HECS
HI3gbLFVOMX1i/Wp2fqoFzPxq3zl+OptmQ+KNWiiT/DL7ItgdpHmzx/4op/xOWQ4+4g4v7xb+aF3
KYoTlZjiPyo/ITiSBFEEFh5AleJh9RUiV+yPGi8pFvGYqNNKbpgL3bBgfQ4JUO3QzzmmOExmFC+q
2/LddoI3vLcGz5flZxHE9AXo3ij3SPgm2GmaLmEgVL7ztShOPRV3uypWgaDbJ+RqNxGLq99+FoTX
wai0Pyyrw1+biVUcY22U/l8sm1KfQLVNMHqpXzsxqOTA7syY4aifjXVHE6gEf3UZ3W7jeWmXMbdY
gFPLPSOV/yjrWlH98q2BmpN6pH5++wtMWFlJopetCYhJkbxFiv6SQVPW/eYT3F3FurqAIPAQdWXY
6/8+5sSZM7/SsiwQcp1SF4ij0MN067EQYC188hsAdfVXs2zmt32sfs/Cwt3RzqZ6OEkhf1ooZnPm
WCb/TmhsZiLQCrPqbMS9HufLFIziaW7B2eC6hOlxaFmaXulMFghWfj6OlPRbje/vi6YrZ+dTNP8u
deXnsUD+VGa9mcv22zM1icPUCST9LCI8PLC2a+Em3Zw++W4bTepYQn4OG4nKhu+sU5Pm1EpwUaXo
05y98SycNgaTWJ81jvyUUyViP4CTYK2+3iupNWpeFd8UF7aX0pCQuCa8VFVJPpIVRn4MTSBHb5kX
3/+n95fj62lrjAUY/l29mV6YJr+4nZhQUxHNOcVysuHCCF4Bf94cdknffWmL8iPtONyNGlzTxOBI
x31RziQLBFhXEaP2gs9cP2g0FOSj4zAlBreSQB4KXjUYOm0a8NzqKSoxnp6fMoAiqo2CzTWBWXNE
Ty8K9rHG8wPeKwaCHos51635J5LJlZ4ukHFZXPP9zI8isQM7ydtjT80VMZHB3RSt5PssfZZmEjrS
nwYFSqt3fThn5FydGpctTes05UrL8E5opDnpsvV5morxtIj2W6kFil7xN+NbfKa/yydWPwtMtELS
xwxQVO5myBYDX+v+v0Bchq+QH5MByC6ezebN61rq3bNW3d6PmMbOvtHvFjKE+5iQJI7BQ7y1T9zk
qomRsZTwAxDlX95EUdZWnRzHem6AaIhOJ0gs5SXNR4p7CzNa/09jOvCn7cvzWg/dPC+yvtWPmCfN
WOIcRIW8+a5Hia156kElWAqhtY1StQaksWihqnSYq001MHDVkd36+d91Ou9jx0qHjgbNoyMkrGvv
F5fRmLV7OfY2nTbP65XdPsxW2cVqrcfUHWxDaTeEf7WaKFiv3gcmzIiS9EcKsIRXaZEsoz7cdGQH
ARhwIqXJSyfZmyU1bXt45TZfzSmbQIA3pZZFzB+JpRU1MoxC6Ak7N3dsXQS/ALD3G5rZ+dLWo9PS
yWzAhe7DBPq/gM+AefWdrHVDaUykJDRMAgNSFZEIbVf+dDrAQFMTjPdwM56R9dQ9uozXEBx1i29d
7VXjpeP2Rl3QD6syGq3SUWCMCbSlJnrakF60AHxbvkwc6ENd3bkCE2nmXB8SEpM4k+kWiPe0TalX
DfGKVKE3/3w0f26DyD0bZcCWcEU8J5hhiys1FwUyZSP+bArsfdH7q3+Ddc+9smlVEbvPwKZNlyXZ
ovRTvIbrIqvpPJBQbTpAcNEykfr54Gpl7holxj1zVrMcU7GX1EAr5rCouaeFD9eR2PnPRcJczrLp
oGYFlhftF/VMnnQETeeX4tyJeiwvx9DBApEJEIL3a5QalmrsRv16ylq4Se7nPa50KGLbZaMSwiCh
kOyMGs012hIwR1QuMbphJBmAzKHv2d7F7fw+Zhbb89hNfDvYWCmCbYhAw0ypcrGjMC4mLqn0qEg2
mgf2UlE3SZOh+I/tGikHa7gjh3O6Hm1fVwiSoTZD/3i92eXjXMuTIUL07VxjSZTmkzjTmd/BdYLY
Kns97sdtWAeu8Qy1vyLDDBSYXzYTi3PyA6WQQmphqPv7JJH5YUqG8qlP+gM+x5PLK6sNlBKliMYC
SQAyJX4K3FhEUpmmNag8MghK5s6j+Vdgawofrzo8dxfsJSXeBMMcH7ON0PiP0rBl3WroXPVbjmOf
gCkNp7Ax5pU83xXRrYQTxVg80iS2Nslvdo9lSVflmHh25mpzpXRUxWqx5gfznyXSO8QuzXM84A51
2wIbXoH42L/07FnbcyqaS+VFuLmpqu/QbIWXIDxliQcfRy6TJaF4YJEPPr+39vw0cVqSfIGvgrg0
8fd67rDEOCgOZ9Sop7lc8DjIuvgqQHqAIAImymCe/85IEIzqBO/Dxmv0rPGFFjpwwTBuYg+O9YzB
MfwEHcvQlmwJP/K/2sXfekgq+0zK92VgcZqOM6vZes0uh12jjqp4sMZbGUVJbwjoNa8TWiVpriNt
7EGJQ7dZyKZNNVVIw2CnnyUZ/WR4xsbhSFdQ4j3Fnz6wX/FlTtbk97zKHdP83Q9wUkOlKacz+LXG
3S451xUXt6Ek8BVO8MKwxBlRgxqjneKQdzERyJdJ0lDQe8SeAdoqy0BVldnZQkjYMX64UcvNqYzn
Z0jghaumsZczuKUTkPOYB7TYzBbE3iLI1Yn+QiXwTCIjF8HirZweqDE3v6gHUcYTFQxXrnBC9dsx
XjciF/P9/OXV3RrWIrhD5ldy+yOipgKRVWp5HQq85O9Ygyy9MlcleQGUPzDvfwtGc82UpaSNmi8J
fvs6P1foFF/iPpItToSn23EED4ra0aM2vEPgYhvKGndT0tARu0EYNgmlNo3/C6J2WpbtQVQoy0ZS
PubNQoL9u2xQTa2fP9kIj6lgGgqR4sRghnLgLnkhoa/3Hxs28k4Vy568UodXZTxnFyQ4JMSZZvpC
8Ps8fndxoUOtO9UYhNmWLhls/AM/gdvkRIQ3EKttqIkcdIj+qldwO9BJSgi5z4SJ5BStD6FN3fiL
ertNfND5iKEYdztqh5OigRE4AkpF+aD+pIBPaBvp1WS0NFGC1Ybq1eJyofNULn+hSxkaI3mnHMWn
oCi3kdvXZ827b6siV6JyHp/hOP/LZGJ2MEQfJMtoF/+styRTU0eCdxlotToPzdFMuDl3bnEGedKK
/fl9yu7OK5E0AOBW5aBm0FiTOe5hHwl8Txbb0PTS5uGCKvAlYyvG6SGMl30c9u8nv1WXZEk101Ve
20rqzd7lQOhsC5JFW/sKVWZkuvfuxh6r+qOe/MPX3+srkgjW1FwQjWQm7hBKmni4hzdkGgDFmuq0
EoO3lp9ZabL19VWg8nWU7TJGAevf11F6NCpFwUlfcJyjEsw1/3FCvUsPZ9XjSqg/USJj4Ty303av
c9vlh8ZxPv3Uxme8SQ7voIo5wNbP8QfGJdYrWidnVSFwqFM5qIer3IrMyLWdyX1kYFavQQJo/jU4
hlH0u1pLpUdsDFGZStE7SoPZxflxvCm+l/tbm22zZgWD+BuCEZJYfQh4BAtRQch8hNt9DMfC/M5z
KV/67uKO6IyICjWlSfGpVRMCacCPiAB6FGKkJ2MkV7w7RZzUGKtCO8GSicbkWTDuW33rKxwqd/UG
NYAsPHHsLxhw4EraBvmgkg6uvqpVzdkI1Y0kpUCA7fEHrWW0sqFbInLUBO/igW7TmbmV+YJH81lL
+BWtcYRPz2KLWocCbdWV91qr9Cc7je00Azfutb2fWmr6OJtHhZbC9jzahIKMD2/HGAADKE4GMjoh
71Jpc6GWFO3JoruA3rFXnS/NEp/yfPOpkzgP3PTy0GLOEgk2n+h3hvITHTmnau+rTfsvSpg0tgRB
2LET0yjcXeS8c1HqgJU0mT4DCnB7rlgF0gufaKGzTV5qH+mqcOXwA7waCN2fIUc5gGN79AbEIu5q
4MW/v1ftMHDTGPMkzJusCHwUDTP8QeP7kKxmDt02GAtBq+LNq/fScKJvh894tLpH5hkdI87nt5cx
15BYap0uiS6Pc5mREvyJeonaFiZSiJihgGSQxhVfmQk1Mh0WlRW3sMhD6uzOZMtDWhDpJvlFt/Kt
4uNmGkoEIyqZiYNkCBhFd6AlnJ8e7kHFU9jmnZdMYxujT+R6yv8MIp7cdcwQjzbjjgNZCp/lxyqX
R1RgbYds/t6o5JNk3elDTtYKu6sEHkBuU+SGYCt4fgOYALv+pKxvipERwcPjvqYoU009id8ppnNU
/dwfGCVph5xVkXsDIm9fVR/Qbc+DZt2dY7gxFq60SdJHs+I4km6IzF7B0GVSKKkqRmoLrSrmEbxa
jbERFqmB3MOQeWeBAJ1i79O5q46Tp5hM4VPqFpgjlLHfyn2okXY/dBaPx2CZOp9Ky+UBqn9voLXP
U0OjWMmu/glx4dVW2KvQDyYnqDHeLMz+vA3bl941GE2eoFGA4EU2kUncrYqSqFit/qaL1J6xm4U4
LxgmeXvL/x0c0q9/rt/bYGIDRZAa5BMjlGB1nBs7mZ2lrfdUU84cg/mdxYtUOjDmCm+TsLSdENoZ
sqYQVcDBxqrimTe4r6jpg6xmNMkJJ0qh6J6HwK2L4+cxV9IJrtVHOmsEherXoBbs8DQ4IfXvsnfj
n82a2y0aSxI6XL3jHSh36kjN31TmxGqIIW/HNkwym0JpZxd248kjGQHLPxpO+lvNTukwI4nlhys9
Davq4tb7SXiIQTqppFwn95r3nXhulL+JoU45LbLEC9rT1SZpV+BzfYoIJbHQGwlUBvNbQKDwbtF4
u8EcYCvy27/MmaIUtp/RJlZHi+iJ3P1MGGStrRuFq8rYBi1dTovK7Xwv5KTW3INfaXtBGvxZtvRR
A5Mb8rrXErYrNLAAItOB/gNOYT9V8CSKZmyMWqhHnpZl/tWtYQFUovSxz9u0rdw6Xgk6RTz6WVRZ
9n8pAJMpRyrGsF5A6jqzC+Qrss31VBKsDTHCRmMRE4gkRJ1WHAskoFr0ahUoTDwSjQrkY25pjCZf
S8EHYehzW33FQevCF2Faoojb2UCFdiE4PjEWipAioYbzSP4QDE+hFThIsDfk/EUAcHT1n8l7QIQ0
LO/ikGZ/Q3pX15ij0jPgu/LiS+gbUHYXdmEjYGF8JXltKD6yeztJvRlrNHsTsEU+hoY8WWEPQ6NX
hovjL4jHvfhA08W6Em8wPlKROg+2/a5sRaZPO2TJdK5ao7Gmluiye45UNxXCD0G1K2v0+jDWryrY
ieFqhzkRxg4PrhMwKHRXcAY+1H4y1lJE3OORCt8PVY50zMen9FDJFc1ZYH9BKt061JA+uXS3U7au
XDXlYMXaFMoAx2BnznEaEoS79pvkQ3YcQYVY/t/6oofpq49GkBT185i4Ni8XS2grCitw6NbQ0jhn
96cLESacxmbzj0TYQNQpL8paluJJJPS3d73K+DDKQFXRr55FIvA6Qi+1eEJIGmxQkumM5ccD93mw
I8nTJC58Wr1m/8KOnI/tQqfdHBlyqh8tjscXpWoKgmrhZ3VSDc/TKzQWnCDZaw9xK8sgbz/ku+n4
Ofj3F2hDFGwgXO1tfxcqIVhzMHCgWnyeEc8l/L2lcppdtUFu+Nwf5Oe3or41nQxREl2T2HXsDjrn
JVcxANqPf3jssUsX41kLhaTMY1FDODtzjm999+EWnoyw1EAXNcXejPLb4pyMgzkW5uVKU0rJnowH
2s2kbjhIDN1bx9vWAwQInHmddJLbJnByeKP5WkWufZy7zPSYtGnRRI0ozzLGPG6PQsHN4b6ZogGb
Z9JBPkoK+ikde/fjLDs4gre7yx56Me50lC8HnEgC9R34dG9EZdlk/vxe5+6v3FMbrDn3Rvd/z2n6
XVSqHXXt/IliFWwh46HbMdtNtt32+qyU25GEzsas9b7xUrmNFHWwZtBVF8tWH+MOHCoiRhvRaCZj
Kwi6agK8kZVGdW4nmTXm35u0oW2OZup+0eOrkvi8/ic7WGS6JEKZoaEktGhk4+ifWQ6Du1T+QBKH
PyPSWqXFu33vEPfDqilCe+66q/65Vk6SGEj3fIllIcVAeSTzFedKBa+6kMpxkJ1HXgGRDWwMaghM
D8hfMD7N0lzACSn2m7w35fRP8rjCQZVho6yaSGt8qswg24OHgMgASvIk67otNDyber92sp9ieikf
6i8adBUJllgV+VlFXGcq4IWy8taqBjWnpCOStSUEzPU4dPNFyH0AErI3+MsjtilXho0W5pPzSZhU
FqKKpy96OoGiru/9H8gAmVPJV4pRv2HG5hpWqKRw97deLmyyu+wjAaoh5ZCWP2HktMs0ZRlk2I0R
GlJAj5+QrxunekJdCUGoyray8MqjbcGGkzEzVubI+cHIbKKNWOZr9/1YqnhWFBEM2Z3r0DlC/fSX
5rGGdfv+ltzhEht/sBYgs43K7BsCL238zUms1kP4sg6SXk54OwtfkFz543QBGKeNX+QMCTOvJ8vV
1ZId4AZ4v8szXWkAVFPnuoMikqGGYF8ffaLCDjXBryDZFvzDAuseLTLcUGrfiYE7PYkWqncppIM7
DBbd0jonQnFd09yIiHMlHoU2xRIYhGjkraU04bzFCIEJORJRAJaqFfrH4RuU9Jgx8QdrF7Wp8+lQ
L/SfAtO2hfeOHVxme9PwHXpSU6GIwh00gUe4LHzJl8484Q2Fj48b1A3WDuGl+gt7s9ccNoOBDfHS
5PX9WS+TU9VojUws+Gg/j1AGdFz4IYUw406kiijlICkPv4DX2PJP4I4LVIu+jXr6Jea6l6jQNjXl
CDprQu0xL3NTV0sAWbisxp86CUcTQL1gOaD+SeTc9w7ydwyKpftzpKO+UKV4bt4HezGd9SFCevml
e0Q5FXa9R6ysqr6n/X/9x11dnNhANKnEwyBzFdTeenGwKWGiLAPWfU4hy4krYddY/+wJcUs3Omzi
04wJBz6GnHsuOlvl9i8wWZUJrj6udtbp/Mkp2ibD62hW6pRjKB/K7LU3z004YQAzPPTrS2/Af0uT
QW7gYbNj4BYLMNV7zM2kRY8Ll2BTgPIP/GM1rL8bhdDRNkP3uFEB7wkYVtxVf360zDF7TtZTWWD2
Tgx2gcT4VQF/NpeUVOBOm4ZRdgSszTOFBH2WukxN2LO3vGe2Kpf1jbj7dY6VMMg6NhRwC6LtWkA+
Mqp7X8XTeqvZHTDQzGDItJPA1oR+bCLx3LzW1rgpm+3ZRIe/oDamvCq55XUVIFYnSpD8WUlWjM/K
MlcqPek6vzTDR9eq6j+w2ZvOOfakddcujZ+ZSBOkgAIpjsS5USkRDLz1yC4TIQFSXPUil/gLlH7B
9KLIyVJVzBomIy6qaKcCkAtpYzaUcqQvT3EN8bwxV3uOrDC/rmFirDxEoeOX2B/vzs/KIdxkHDLA
lHbw0gmJYt1roFEopTVUXHezHs2q4CI/UH6S6NQDkl/tt153gPI6WMuB9Jn+FZZKu88rKDPxO3R+
ghB3vWRrajx1ei/VFg1mhXK/B8XOA9IPcg6MQfX7CcTVG9Q6ZxQ7lq1fe58bhbuzIiW8/DM+DpaX
32ql+D7kCIFMcQnqlUZSTEa/tL3t+cFQ9xEAhUEhuW24icWnmRKDzt/zKPoTKpi2r2yTb76yzAwu
5krr5RYkIS3zqLp6fjUeCLMOAt8h8Y8AgKoJWA//pFawCLS/JnVXrvETv48H7cicH/EEE/233zlu
dVU+ntRGrIL+OjczkFC3KVeoTiGaX7U0RU17OoQ0jkE0sF8sYPBSlp65cKT8pFbPRO/a+sWdzrF1
hBYDpojL6vTLodVUW4j1DMKUkPGrdkislmgXUk+nkmuWLTRSpyxE4TqP7hOcGfSXpXDhgstWR882
YSmvxk7AOZg/z0XA+6rjH7oTwRYhi2hvXYIvfsUdUOd7/jcembl62pul1/ft3LbA4VL8XIJ4zoV7
crzPmSOqIFY4qxR2WmUPef4iTKtAg50mgWWCupvCKxJkn+DN/+edrfp+9xQSoxLZH8hsyuIq4BOw
HHrvjx/22JdiUdcXVlUP51TqXfmasc188VWZTUjS6xxrGlbdjUopkmVSAWrmVA+ghS2iQCnApwON
OV902cOfV/p9cA81NAzhrS5qhsmjBWO3naa/zmf4E67A6JGEKIvPxjpawqhP2RID6qtZqQpH20XB
FUHC2SGLVQnKvuJQVOJ9U1psLFv7zrmgh0g+/GtZC6F0XA1T3eRkqmHNwfneKtnjSw6SfdhTuxBy
XDhE5zIiKYHlKOr+uLjk85+CWDoPQlO0xhcBTv+qK6OaEMgexGiGrAj91/W+tzKWOEHtBfLIUO8s
mvMsp6dsD+Fk8iVhUp9Km8rsohCwh+qheJp9Z/3+KGWSknZPm8jvvItmxV9CI47CokzQHPu7ByN4
PSEDOZ2cgu3ZimcygFbPQETBRXqNxFrp1ZjhsUl32BVYEDcHGz55D6p5Y9Iyu/OtCVDGWpTSxQAZ
0VGsgAHN4ethUeKLwFyngSnn6ebUxmfexu/GYHwzfTykH3dCVw5qpjjpFwKqkC036lDit88WRvxL
OOdXAIOxVd1xV9jP6UKCEx7i2zV+OCqRwIruAGITXO8cBQzj1Ka2NDSYWDPlCCyBnX4ShojkL9lK
2Zr3TOXjlewQWXWnyIylrq8w+pS5RfPZ8vfuqEkYdnRZL+fqkm7rojr4sWYLffJzH2ZaamGB30fC
EGmsY6RrA2HmIXrY1bdd0841AYBc/4txlJNJZ/DRl91H8E8Gpl7As/TIU274jLtMAaYzlhWh1DB5
V4XABtGZD4DpJQ1yOxU99VhH4O5k2fX/4jtiktTr9QSE8uZDAWvGdtpBBdjJhe6a0MeOfJk9vLtA
f0eDhPP9d4o1rSGNTRXj60f00ommQtkFz2xVYLGSemwIg6hmuL2DfYEf+/j6MJfso+KGUKgYeZGW
4dNYz8PNObgj/TKYoXQgyv+8oDuZfz1soCFC1Tw7DNrqMBf33Y64UyGbTRfCBHgBNbnOQKWN95k4
Mrtkx5+lkUZILGfCaQzHn4u1w56mk5InOQTZe5LKRLIg14i73TTSxKGakjffF3i0pIElZvcQnT5/
Uu6qimD7cIg0isXerKWyJ614V+6p/qBapjWgtGpWzlOyh4mcSx2ME4kgiYOLJIgpVyK2hWxAx9Hz
HNE1UnxhkxO8vg/ZB8UlT6jUEVqQZbjFR9jhilx/Ww/Ew6ZupiBQ7YOR2DC0L4qy2d9haWjqGRbc
5rRb60v6RsGGi1OGLgzYALqAYgcd++iqyQ9bQiXQ+npxIEq6M/+UjcCtc3ydlqO+7x/KgMHV1qcF
wymwtN/1mvm8hGfVf6ZtZ60RWBPxhRpMuhyFvsLQSMZF9e5hYdIQ3O3ZRl7T0EZRKtZH4sypXDqN
lFgRr8R95XeXAUa9Jc+0G80+hJyIfOVy1xar2v+ArPqfBWjLjK+hhv8z1kurbjw8mLRhGrWbEjSE
MEVM+uG/Ms5zZxyXatvdgrUOQtbSk+QihWSVQTC4rmLTRW4Llmf9PZ1Z8nw17jUVUw2wcXVkbEBD
23fcs++L0XZ6Nck9LfPqYeosOHWOY4IboRLkxtSCG5zJOvxQuBcil++9AUqUVNxJpObQWQ/bF043
t3xiO4+BEa76c2lOmm89hpjsVoiq3+JQ5CnK4vtJxCZ8PHQrxfyhcg2glz3wBAR6CzdKhGVHhqlg
v/ZAaqYQoNH36ty9pu/oRa9peEgiaRw+oqdK+/WhCK1LAKZ/M4EaRdsjPmjsxPOXNY/dvi3uyLgD
NzZuloy6hRemsvYICzlB1cQHIwZ1VoIJBpHhD9run+qK/yGxK1oiE5K/ahz4yMwS7Q0Ac1dk1XMM
YXvQctnAdWEs9t7tsTBGZlw3DcDD0MEQLJHzWaUXq46Ze7kmdoQNOTJLdBV3aBrWQAqb3KGjRQkp
CyNYz0GfC5S6r3fAQgSrVaw+ewTtL9aHpodnao1kYAx8NmO7xyxiBXtsLFVqyhxhl+lrgMuQzEWQ
8dtUJZcasBdIFpXwjpGULtZnICBaaZIH8wGHTWZIRcAgOgj9NzSKRhqbcpN6IhG8SJI3ZKGaV6Gn
muYTu6VD2HPC2DvYa1ICZ/zgvc8MkdZW4/xxXqXa9BtXjgFIhhnmd5nCYCrKHWFKGFSzyRKDjUp6
qOSSJ0ld4mnkUkbIm+XCOoTRDj201R7t4JXBT/OJchqu2C6HaYauAJfdMCL8oe+V6pn86U95mLJS
KDJwYAI7hqXjMs3IBzZ5yLjyIDMyhzCwO0Yt5eQ/SFmTRtuHGVTU3I32/8OnovsVzPtZoY7VK70J
0j3JEPUmuqivK+LEsQVXfJCgNfxBj7T/IiCjGQ6znjVDSHnuIlVWnuvplWeoHuGvGEVJF+1yT0RB
IcPeyLfCyfk5erJWAD4GWiRvmZwJ+vF9D1KorIaRX0kMqnVT0JOcKrKQhhghi/+DPwHTmJ7nI2hV
AVGVG220/H8oYjNLEG6lMT0OKNcNlF4Nz9AePgl+3fCKF2Icpdr7viVLYbAM3hnOjmDjCSqRv3I0
S7cLklp8KI/deKww8liSh/GTE/bhujph4pJmu3eChLzhM8sXx/kbEbSt9Zwo4toHgH0OpKCDH6zU
QEccPqpyd/L6BDFNK/KyWETcuOujlb7mDxq0tLzLlG9EHA/DOkKvYBeDsVX8nx4pPR3ieYY5mqsW
aOsHZDIUSi8wCkMDKzbOptunvGQ5JdgK+jUW4Nc5HJSek9Tw5dV4bIDpqySbrYPDTN5j9JiXzriT
+cKYIeX43au2TbwBnvpDcCMP+X8OygsRbqQbnYf+gZmJdflH8QmHVSNhQQD3aEOqPwMcyGSt2SjH
gOUYHxj4iOqwSzJKglzwlVfBMMTY24oJEQH0Wj2omGuEQunuYizpNvcqEj/gmU2rAlbCG5Om2yaw
sA0KrJGDFgOe02H8dj3ARNF3qa2L60cQR4/AwooKeJ3UkRBWTAYNEIbiESz/9zlzK34yF/cibnYw
FqFhpM+aDNkH3nnfEfxcxx4RI7AufUdXFJmCiQ63B8A/tZvxeMeDZImDiXu1nnXOpmzoYwUi1MLA
bZuvtOFMnj8ER3bkrgZOb2bI7TC0OmjAjPlKRWqQjBGh0VfmfvhCeTpbwAJBR1It7WLc3NYvrRXq
Y5rwdmHCWG5rrKmazS6PWE6WedcJxeD1uoiKHwJCc7A1iyGTXit1VUZOx2wbFcZiFADIaTp7mWOe
3XQPMEabR2qcZXRHd9Wa/v2YMbm/5RdGZENV/Up+BxEPae5HFvsvrOO8zgO3+ZSkepyStmLT5NVn
kgP8E4FWKV/FvavPQJSQgSQqm3Jtf5HNS0WGxRbhb/yPZJHxRAIIELDyjHfUYRy1GrOO0CsH268/
wVsTVbNvYV8feD4ogG49a2am9i5GvIRJPlMwHwoncFWbJaRztJ8GEBzrllwsrc54k2fB/tcr4sPz
jJVBNjpIAo+Cr4wLVMh3JMUkqHZlMbRpAYTkByocWPaSORDwJKg+lkeGEZRUAwpEkqaL6O5+8fFe
rH5sIFBYP2MCAil2vmzZryfR3Hhpx2NdmHgM9YEy8rCnBQbsdYGi0muayRNkjeFzunfGTKwmL+md
qNMpPG8GyyX5Rcfttom+r9/GXxEtdJCHL60kFynygcqc64QyBug1jO2EPqPnIL1IH/vAIgYV4xyf
Y7YdyPAZz9hXwJd9Z/Mb3AcF5GcChAHr0EqlS7FUcejnYeTHcgjEyjSQuES4MnKk9kaI1FAhEHxD
oWyROQI6WV+xRu26IOxBWhdmAoqQsnQHYiV+OB9xhIiiBOvxeQ/JPy/tKfX7Q6LrSWb6IOa1PcTC
6TIC5S/d1pgDtVej2g9nboL2K1QJ6VcKG58P8Zo/+tVFinW2k3NNEGRa+5fiKD/kfaIFZbZ5zfm3
qNCDWFL15TQ7UlT6KI2MCQBzxJSyrnn4seOkoi2r5iIE7nSlPY4JdKGft1HCBzIc0iyVJoFX/Bhw
zDeqlkx+ufU5yZkuSzKXN09VKq1LT6xsWee0+b2YJFXfq5pRx/ZTAaH1qw+HrJmPK3yyScCVT3yU
stXIR+XdEJdQv4MX/ZvK+rc514+LmL5b8maW09BypeDF34p7k7SmsREBtevuAafIKDo/0/v9Yaau
2KRF1ugw1OBlhovc4mFzOBs3evlNo0qOhg3IDd9x0P+6oZPv1ysVU4NOJE3yPp9abUWORzvVHw9o
XGqDLSiC6SEFvAueBmt5CqiMpu4HAwMeUCJGA9nrRHpgcQXw9zUHINZKUW+vmSw2iPzgY1Tk5QhO
EK1i74CK1FlsnWtOkq78eQYcQd4x0NLvk3TyYjWyINvluVIJG4+vSP7KQY0G/YjBUAz0Sc9aZu/s
3WRHUfYEcGAvMXXYLZHOcUIqiYFGw10pCcLChTWocNX3tdVzkpYiTzZgdiaImpRXdhV3fh+v28BO
s1/YV3ajjUQOmpfrRlyNMBwR7NG8oHKfb2QEP7Qpv0sRhN6c4VdXXCFNkAjnBOkdR2hZGz+aH9ZG
wz/5v2O8umrc5q37fLzImcRrypwZRGonNrWUboC0F15ySTVXl5HIPRJiXILhb9TngXbH0WTlEqJR
FPVo0jDFhbQz1NC3mSkYvVUOOHEbULrG8PTlsM6e+tx5/GuQGnA/Z8rNXiMlogaOAvvu054Bm2WC
zScjB8Hi+Mg89iEVHGykO8t2xF5hFZRVllsHc+pZkeG/4BnU6BT4mkx1Er10fPE/NCBRI8+EeVhM
1PSAhdoBe+JZNET+K3390yZhJwgs8rj3Swf6L2dR6eFO3A79G05oFyA+F5FjU/S1tA5wTwv9Mb/L
6ssweR6qh8gv5HdmOErpYFQZj0sXDNmvBkFa8jA2aUgyxK1VCWsCVqniqhjglyzCcrj4SDOSt9Jp
h5YvsBjsSTkCPGR4oFF7X/KsPWNjhRfuTI8pV1PfC8rmhSrTzsLlQhfCfSjKB9CMjhg7GwcupJUX
2Yyv4i44F2bPq3+v1bnt1oUPfXCNv8mIOxLEoJS5yCkUbfCVAVlAq/C8LCOpUXZOVlAWvcoa8Y42
xfyvAHb59iy3wFg60n4DMdr/9J6CZG0reztsng3peMp/TMR4+oUyZgfxCmgqbCLK0rCNU7hYop08
6qtI+EEZ0F37jOuQ/+MesFFpCcvURqURgYtVAz9byPRPYQt/j2TY/A1i6JtQr76HzI3Zt9yYamLE
FdiuVYdU5pRmKNQNrUhB1bzjHzN5GAzhNIiMKZl1pti/p6gjyjqAwu6P9t7KC/ATVXRGl/SOYhzm
v1nf10M8Qa+As7BWmTClXvMD4rKHXrIDzGyjS2zemvC6zR1eWMfhXZDMfbjEnLoVTvSS2NJU7Y5A
dOD6KhD9f6wvd6+Oq/xVlvqW84P1mkTU72IVYwYTnPyRyD4JrTAYXZ+601FclepFQ1fgcFMv7SP/
THx9gY1CEMVoX9PCFEYpupPm60bgWaYu8d7VePBGW5lRqmYKnu8aj2tKzYOYXvlRPzeXppfS0Kl6
t0ZYovonjqU3erIoOaDjyOotQQiwxcY1jFePgIsrJ/5tPNV6/dt06t+Av6+m3+zNijCBhHeotOp2
hweHGQCiJAcipT8TTEtm7huj7CpJFcnY2ZxWXqX39PQDSsyHXKGbeEcJxJ999xXBMr7IQ0iDtBsN
tcGcTNcz916MevKzOHZEHndI5gzxrYpj+lYBOICUbcIxZnJWOvgh5Ylj6b33dT8yvUBDa1dRyOQ+
e9LvA5uBzvQfifN3RoTVw7qssQaPU+f4PiaaZj7OFmfS5YPDVi0Yam1lWs9aCxs/40LyQnadyQan
jdjbbXKMBBZl6EzobBzgZWq/LI5I+sEjGqPEgFgjAUONAvE0IuH/EwI/d5s0kvxhnuCMPmsqERce
S3Ys/eoRoiEonCvmb9952a3nFaKGUu7279Hv6T9/wG4f4id3CE7Td2z2YPmk4eq6w/6Ms0+MdAMB
tPuBEDlpP8hxqWj7cpnrk2T6sfvDbUWD/tQ3XuxSp01dzgeMNGpLSS4MWtNyM7WYymrqY6GYjRst
yFXSWKYEQ0g41kJWdoJyxDdoMxysV9qDJSz35dhD+YwTONA43Llk4KywCTtwDxgS0gxPGfSSKRO3
SMiIz0ju+ktdOMYgN8fQJ0abUUAmievGy0v918rO5Z7ArM9T/AuBdnSiIDW19S3egkPOgblgz4E9
nPpRnbv4fiGeMmFylLBGkKBKhenbHaaMv1mCp09wYFTl45Dd6OLL81IZzGg+taXq/Uo80zLUh+cF
C8LdQcbBpcxjLVw4w7FzHiRRoEJALQTzT98Rc91jIFUpyD/KX95qBZP2TYRdf4cFixJqtwiHo5Co
C5V4jg49lnLXCfkHjGofOf4f+X/y9NrwTb8ZOLSxwtj13AV7pZdJ8FbmXERJDPuWyLtOh+lEJHk9
h9/qGqyoyWuBXEViHSsRYpjKKK7tsus++kTry4t3jXNboCE47JgCrxeOLqLGCcBCelRR0LuzLeiO
vHH7fADsVdm/gTdP2qTYYLnMhGCC1mOf00E4I5sk/nYiOJCJ75kwlCIgiGUAKZyVonSfjLSL4drf
CY+aH7QSovInULZ62knk8yXCXcK8dDZ1X0KoZJ1oNifvzZbnXtJGf4JDxFSFtvmYRp4fllLvvuCN
tWB3R530nT6qyj3v3oOKHNfWtrYcCJP0mKhIKEZDt5MdSlRh5CJfAe+uvB5sxMqv5OBOlAhRTvLC
/Qxy3/PCuFTFXF7pWA4Con1Kj5llX9z62MSJyD4q5fgv2CZC9TXzRDSgIAxS18FtY5IIgNK8DU1E
JXcKo8KpVLHiP5J961axIGotjhmBB9RFyCxgZ6lvXFsCJhU03COMtdNwdaE8iJnR0agRr9UQXtdX
EMfSluIcQuIcO0sKK2IqFoX6IBpJKkqfXvnAIzMBmnKVZb2sac/tc07p1thCZPzZCpUI9UwpZn5a
rM8J8YcWjnAj7uf9yRSVf5vXnUpdKw/AZb3YKMVYdI5AZgv4fWr1bY4KoNTGOb3IjJa3p4MvMOrL
MCe7lEcehDQoIZcJBKEngCqnReCWQeXe1S0tWV8dL2QGpYW4JD6auA+2oIdck+Tu42J1WJ0fZjKq
ss9Psan1T4L44VRaPVEFKg0rQzE/IqkewtIdSKXgoyThjf+pt0yl0YD/hRXdYDKbQLUAshs/zut5
gWiLXhoyplTkoFh3M0vWnzS5lX0PDoGHUPAwqmT55uypnHM3su1hDSRLTkJqDNUBeXxrtUGu6tZ4
/+lAp5OQCu6/ydyerang0akAfO3cZI3iGihAdTXRP+7QPucaaaiodHYwa163aIDRIyH4Jiufc+cs
H2STnJ2MqPwnK9UOd/qmCLe2Z7Bw9sNozGsjj8obohtRX8MXZ+AAm0GuGH4jS5JmpdgpQ8D9LJIR
JaAmpPJI6xlBMXJcrIF6/xyDil93OAQRbxf83NSLSbP/uOAdvlLQSjrs3SSI1wrJ5OADe+9Am3Ty
61xljoFeNR8hk3eUkm4bMInPpoR+MzhaftyXjCfsJAgvV5sRM3bflWWcZeJQKWd65MeuV+Irzues
tyirMkuufsOg+whkbvIWRpbm9L/mF2sNeJ0vPkY9oEKhadsi6W5TlCX9YSg00Hzxp/D1Y9bNdM3s
gaemhGn945Jxexhrxyn4hSYU+2czDlIRuLr1EGwI927qQwVqaDzvtZFrpp/gHoZWSVhqyNlCVQ3S
XVDaVo8okmwJd5+Hefkq1SADYTc3yrKRBEHDUS9iX++Bj0B82ZHjE4A11mMdxJ/NgTDRGwaSDGTP
bfSRYoWynfUWb2K6KWz/iw08v1NITlz7lxsXkQXqI+rumBSAo1JviQrASvj0Tr0WMIT/ipPnooQU
JBrblB0nUrFXfWTpPRIDJjFSv8CCy5JnTM2RUQ6eI1krrlWFoliVweYK/MgpRLnwtUuUfPPLw6Dx
kscs0vve1gL6FTAACmRxIVTlyAFiYoCjgcD23roeedCH3j5rn1MXlsY1ArBn6NgAZ0Fwi7odvrsq
rt3T0yN15CfNMfiZm1XXq3IEHttKgKjSU7Ho1G4cdYaYnzIdAUjwEL9GKxzsf00FlFYgMPHPWJ3M
GT3Rqe1C5F6ORbtJndIEw7QLK0SjEz8aqF0y0c3q496Wt0UgN3uJnaVCCn0+fPAY+llZveL4k+uB
9kgk8LIISftFAAYcFdRPoXmxQkSPOb4ZGo9GulVmvSfNDbK3opEFu8vu5Kt8wnr1Ju9N+90e4b36
510n+vBfhkzOHSezwoJ3KS8RlORCNavbbKZMJdiZBgfR+tYmB5oYJ28WWwiTr5zTOnOz7QNU23vW
nxTMPP6MvglGaELlnsuN/uqwDXrPPJQi1swA3nBCB9EeroS+64Rtm/5vShgUuLGa/mXDmolpy81l
bBA15iS/Wg08P4B8IPYtUSM1pE0VBPTAojkZ9ykn0jwIb1VLAlF3kVKnZ0gARTsgURkylDHxDPFr
YqemMOLzSevWJo9a13UeSyjEYvhmCBDk9HtSTP8CbicpjseDIxyyyY/uaxmei7V3oQ4/O0Pm64K0
5hlp0cPuJixMrpfe4Hg6Ia6ypEVLDYdqEa5JwkVgvTf9aeHvQSpMNjLMuhIYR0dEYOAvxgihYAti
qzTnn7nN9+7FtcYbc5ZicXwC3fC85WkiIQyPg7S1EkbLv6JezziiytJeRqFUx7XftWAAsOWj70Hc
WbqNwn0sPMMNfbQbVGfqtGgYcqJ/PnYIZ5kZsLLpPMwyDZFFSbYN9D36JHAmlqifkCTgPTFylw3+
pOrevnE3O83mBNIEJDtdaBMjWm6RT7SEhdJswhdPLugzRbRXGOqDJLOe2gL7riRihNIL9EOVe7tU
EMqsE2SBiv83DdUuCH6I6YDTeCgSbRS18fO5jkhNytEJS9W8uCSwHpKVHHJukxym6En3GN4ctZ4Z
p+lyjPgVy2CesY7wPo293LqP0bwefGqk+LjrsUcFQBDWJdjVO6in0OBsaUTmDW9jYnUUf9izDhwA
xvft/9J1CAtietUNXE2ZYFmq3Gkd8yPoG0uyJYBFZynXIwZu6HONiGkmgLzCRPsB5zESZrgvb5rx
Z1mpx3t0ovOxl1xGAjOwS6USUY1kJSG/7NqZ5+lXRLRW/UQ9MxVI261knrysKdXf5gyvw9iif2VG
y/ms6TrYBWhpFTyxZmIBDKswz90jxukNIsyMiBnMeGpzQNdijEbFslFRCoGriL9Rv3L2B4SiTWFE
GDjyNNVcP17A0pzlIyxNu9TLdAjLke1som/cBMJN1aHTDEuuU0LqCCg2VIxAprn43PijAE/b4r/E
nh1BmP8YqIfoocWFAKD7BtFYlz6nh/xit49gzOGXL4pW7plG9mGP7AKiQmkLflXC4LXxYjawq1bN
QCLB9GhiLfgyk9PTNk2Vu6+PAEK76HULIIG8XnjBQjjcIrv/lszjzz5LmzL4E3GVJdF3RJmv+gxD
mGqjd87NlZJuj/trpweJM8x8NW2NKQuRQFNLa3Jgrmd9nNPZn0wHD/qchfoyQf08F4BkN4DSHz2A
MjdCHee6ortQQyaRpDnnD2rhA4U8Oz+XBHJ5bTPxsnvox2N6Y2jLdueZtOX9b8FTkktTRyrUaOaD
4Qa6tugy9j5dgtaiPD0sCVUF6QsGsmbqIiBe9qWwNGtaxGaGngiiAV1JCXaYHmfMeEN8ioOQXkP8
sgAHDbXvFGb76F2nWY5wYFug93tg2XAUQHzPz943dDtl+PgLE7O40rdQd13LBwKSBENgb5r1a1HB
ux+DxbmHkXToaQEGAk6nCugXZUdpoh0VcJIEUOKvidu7hp1spbVTpYbWDHh3yrOnlPpyRGWpPKfu
qB1gFEpPwkFd2SJNDZaauL+qgjpZ0DbE5VQ5WEB0moCoL/p1S6KFPoyuBtItLIOo51cQ36XB6kfb
Jff4p+aDYm9bvO4KCCHnTJt7zolYoHh4jHCRqz4fMO2KHpFydaVtn21oHLS7StqfgzE0ePHcc2VN
/YQvwTSpwqMM3wF1juuxrVAt20ieOVWacTFgX3xhau9Scx0VjAj+GIS7Lw6uenI4Sa8a5gO+iJ7h
XxpVfWeAUXwNlDooF0vlbNOqKPPGN7sXMP5rHw5Yb499wjVwy1aGqXNL6jLHWpHiHBlKsz3gUUQR
Ozi3gyuVT+KInQQGiqfWaWdQ1T1IgES+7VqYjE4IkXv1SgmCFM6p9Q12pRMxZnPDS0l8C2GY4ERn
szHlEChvmJpz5qzcWcHJyHf5Y1Y/pUat7PoXKM5bH6qxm9dnnxrdNYk6ICzN6ILHIIVLPdlP1g1h
3wkRVnbDWGK1qJla8i/qenCJdFUA/RgdLI0rF7Uxc9Oj1gVImP0wjVncfD+9YiTXtMNGzK26rBro
rlqtWInV7Ro8rdr5JtI5vkyOGfFus8m775iYIqc1pFgYJd5pn4ksRf6rbVxhgURm3nr+EX+TCpEd
XcpdgsQe4TwcBfLU3UjTUBpQ3y58S9cV9GQoqlAmbOf+9BSLv+d2oxX1jDSfgOIQTX9JNUafrG4D
IKkBVmlHAR2yeVf/mHP2wIljIu3S2N09Xfjh50PTh1tjRevN04zmuecL61+l014tCUvD9HBnU6nw
6UyzyQ8xGd/mmwRNPRWfbkFNmomj9uXQqnFc3nXLh1ggvXhs7dWMK9cb+jNHcgIwia+VQqvLH3s/
qxthgHoqrUHIIhwV6cH/f4OISZQq2iUjMSfhs3sIvi8WJXwK2yJqLWV48r/OHUXdgWFj64755Kw9
jVYK8WpVXFdHlFzckSi1M7JZlhf36Q/kHT3YsFJIX/X0oxLlSWItoFU1I+J6/NWRbzO+nPkUj8Cu
hjONjkL8HW9cfmHzwO4gnpELvjCXYPYHRj4dl2CNgwJcvfiDdwSI7Y88w47UKA7smoZ66M4UX6kB
sqx1XVUlo6EsJQbfSFExyK5d9slJlKzVWwnCm96jZDxZuEVWxSSUZba64kK2asjPQM0c55O0P00C
q9rGiTOWwO4ulixZ54b701uLxb7hr/YJl9wFJB5IVIrDERoH6G99LmzMAh+eyXl4sIA59njdyrUF
O/GI93Ef1hNELNU+3sMNEuWpLI/UzqH/4IuSQim5mxnncV1GQRiVgh8aOVfTWsBZyLMOjYVyB/Kf
vjHbA0mCA0TIdmIsyIro5X2+zT5q9sHzcw3wj+vbwcpQ+g86CnthlSvdjqGX08pkMq1B+9Qj03BL
ehLGEFIwotptUhXSetndIeZyNHJ6OibE7TByp01mlNxi42jOizXd842zPRTcfxFYkBP3nb0YMhIE
rPrO+J6f3sBDWML5ts55a4L+pqUcYbflPclRwIGkeYUZN+iJKIKblPNzUEd83hWXq4D3ZDDkI2nf
3PmIxUWTSes+oO/Gq9JAavWPWn+T7say+AamQWWt/bL7D3xmpMXHvPbUAKUNt4BhyKRJa9cWTPSz
k4jQ8q0aOPC4WgCiH65v55IMyXCfeD/byZ+B3NLfmdFnpTvvGFIZLE5MPt2JPtQsKZ2XAiwSBA80
Rug8IFhKUYH8cwek7Ad3Z100Eh1ZjiwlycyL3bjIudxscJreyxoCHUjgAbakemrpkobNyG9oRw4D
SvEiBvcje43Jy5283de6s9VgeVr52HB+7WTm+t9THLGSbka/C6ImzRVeQ4XAHP7Wu+5WAiaOnRM6
wgx2APULSShtFNP3NaWhOLp6MfqruwcO2OMZzerp5BXmqYf8TF/EmwfmXOfBnCFzTfKEa4SuWWAz
xFal7V9s/gIr3VPlCByIgpzYYvPuwEx57poO6vMlWTS6dCZUbFpFPC6SMrol+5Fa0kjGt38OvJix
OS2NVHVAwQ/ft5J9ecMBY4ub8jJvqeqtr9ecikNgySRn3PzQ94XPDg9hd9jWyGvN9UqpDlTMBB0X
XO4muZSJFXJeOlQ8a9vo7d5zZmEkcM8CNNQLuPYkYmA1+MIc1i0OVOSudBl/w5siUGONqrfa2Q7W
dbvfz9UJfk2nTmk+oVO52TbduvSP0VhdJfUVo5UB7FqIb9Tzs54Teg3xcSQHv/Bvf+zbX03OlEnm
P435ysBjiivA2qP0bWc/xM5Z9avK1XyHeJqYOCnTvK0lmsKv7mJX7jMhTT+bBToc1xhXGF70PPF/
i+SX9JFYQ//AVPF39vE2EqxvHtB2hZNNSE4ixFWDLFQNRzt4A2nuHWsa/q7+WeoKRUyOw0jL4teX
wl190arek6VjKoCMe2H7Wv5ZyyoZAByCvho/Z0OXGF08BsiG/kXHH4DangKtyZJjHKBzu4YterxW
em6bhCSQMOXE+9uIUC9tKumpjBhmCCNA7/2KMFmSDSe3FmhWgVbpdn15YYcBrMRyO9aCMCjyYI5z
R1TqbMSSxBaPj4GLZ8bww/e0MUl4PtGBplfDryVUGP5guwICZLfh30G10tg/iGWJkwD/wD1E0Vvp
qmOLX7bB7sDaMAunZX/0egG9TAsAwVuA5IzYIF6Vd3NGg5fJnB9ytHEILrEI9Lf08U0BK1YjdAI0
P5YbegecIpqOZszgdmXN+HeQidWu+ItfNPaiBsKLJPgpojAypzRvJIaB9QAQnXrz3na3VllKWpxi
aP1gHZmjUE/bO3NzO7RKgVdmyqcDhQCK9TPVX0sJqRTnCgAPxYhpFC6C+1cmXIDdGNJngVmnGE5X
pFO8RXF93hbQv+bWQTRq89LAWpix6EtErygYrAs4dn9WBPcOPKKRPU1mjA3YgN/VD605UaUCrk1C
k45tqpy5oIdQp05LXyHrPdzqYpqgLeQXpzgTnzLTPbOItLN0wUBRJh6QUVMEkNbSZhlTB1c8rQhK
PaGYnUOWp2/0yaBzrYYZ4R7B+3dSazDObYMMWSYH+r+aBbIWaCpB8iRyVanKHATf1uUq6+cPRVF0
PFpIzN6LcgAoph3Qqdz44Sdr/BMvOoRc2C6xEBpWGzCzXPYKhs3gEYWRSp//zV3g465AJPuQHRYS
wz4JD1kcMhQuxAt/vSs1G04qkea3TI3RiN7bjLYYXBRj6yASKB8HDi+3iabBVtvI06xyFuRfAFWv
U8FsKqjXsw1LWlUlx6OurPm95O543Bo2cOCAF5ypaWLIgw9SzCIHfhe9ne++D9ftqkzR5aOrOMVy
SqHe4mM4lX1tWCYf6464yrtOZYgeeTGA9cqaFOuqXSKvrhaCp1/xheVghveru7uhWfOeJ5Q6f4KN
WHeGTc2cpF5cI78VcGBUpQpsQ81m7Q1iDQWI/TrzFaqHllic3b/sLcCZfotDFH4i6GSBwT68Qzi8
KvZ6fI6CojqU1SkgkBFXhR1AkJDzXYdAmSCzaFXhhHLq+kukoup66n91qm1/mbLsQrjphsq3GYK9
fsPbTevzzI93U/EsmNZyMNsxPCcbYEeXYyrinMW3se9USDwiSz9D9IDMsg3j0+X5fI7CnGOIwdIV
nXIQo2kAdTv95FVlt5BIHLsfChUeQf4sz3/Q1de1wgpV05pzav6BSXx5tpZvVsPC8hBHiFQeUHB+
Ctp6Hs5Ph/q5Wyt2VkUqJ16/EJaiCI7g0NIOzOeRv8DhnU+zPF+Ex0QTeNxySki6uKXArwSK+rsd
IrUnZ16pA0B9jHu/KIm62eE3sgOX79HtjHJ0/5UOyidznuON3D6e1O3Syuti3ntokwOY/TllunXJ
yC5B3Zq9do67ORBqp3kGNOm8WL6t7ApWQKLHh2dTV3uYvzttKmjGxxe87SA2rNNJd9gYgaYeEQhw
KOBLzMhf1tB1mpJjJHWBpOpnxbTXnS9EqNR1BZm32UYobsiFPD6FemL9P5I1LX6YvH0zZQrKjFRY
EJD2+XIzkgbBhb9sljhsCzG8QBZoQRiiXSKIHrjmmnl28Dk5zxrfoJhqI9Wttgr1aREZTwlk32ed
QR8gKPMwKvtxm4aK7ZxIpIb+tzvMIwSOafs6PKJpdF+t9nkjxIf2KVdOlSDLzW7UxhvVA65NMn5U
5Cy1FGuZ2sgxdK27oeBwfTdNVP/L8KEyfIJw5pYJcRFABA1C0Eudcv3I0CC252aIS5k7eaizEX3M
I7+dGgtEht++LdfrmkKGur2SHuMVf3PCiXtgw5J0NzQOjZcSJwrmD2LrLYOh7IToMopnr4ZOSKk4
FmO1ND2D0cmeNM63bfNaBRuiNe6H324LPcX+40OQEAfqzt9u3mamAA2TUwbw764J8nmNT/iBbNqV
NK01J07taQhMWdBAtwsNfGQa5PLNtPvgLmieKRhQOAV5/6IZNpIwdCWzbm34AtZWcfQPiU+tyD2m
j7f6C2KMTG5OSiLS5qPQXzzgPCFDUjdJm0+qdWEi2MVY65VTqapzf/pP7OTg5BhrNa9wb0sVEbYS
EFZjZxSk+n5CpKQnMwML9P+8728WXqN59+gD3Rf3rKzJYoGDZpVo4G5k0eDY7qTRKDiKHm00t6kl
qgGESvSSlEU8T+fry41bQAN0C5Kha4KZ6Jqz1uE1gdMEj9xnpymu/HCGuQyjtQhoe7TjKUrscKsJ
SoTP2DjyotbnydXG0JCbHubBduzRPttLlnBiDHCtgUWBZVQisRzGESKYffsNDtgGCxjOrmyNs2RP
7DaXLqZC7B8bNTNYKWkcmj23kx9KtLGH0R/goN7VR2FFrgayjLx9zU5+0JirLZVey0/d1nLlfqf8
7bYxp1eSrXehVqGi/oIk3iYEzPRVToyUXrV7qydz7TbrA/2ylTIINARqF/laqQCZ6Z02tl+8GrbY
bOFzKQEJGwFVnqIqLTu76FAEsbCUxYpQ6oFSWEhKTfRF2Y0bF0b1Guvj8uQv0Q4NBduqNkg6C/VP
oAJlz9sEtbAhQT/u7tfRGkBlQQ/m5BJ0PoMA6Lw0weN0gLC8os9b1nAXAVrM09iuhFwzLogMe1Pb
jO4Gf9PxpVc/8p3vtwwGeLBSXIEQz/qERQjopM2tWhKrfgo9PRLWut6IvBFNY3TPf0wlEeUR9h3N
2Asje2iXofNXaSGZKJAkDbF9Bn8lTe4NwRSIfsdi8SV1tuG1EfcTQdTbpl9mOUdSdQO1N/i6Mw7d
LHLufo0beK0MZuff64xXrJemRbMI36FJeoGltZ2uVtaBlIyAlB2hYwaBZBoyUhWuH7CrP03ykHx/
T+aQzZxCPjjVd1/WKjQgoO6LP7r+3dnnNDz5dNEV3tcNVNqOnL7lqRtXOW+7BshD4xGlumQvTCXR
qqzhg0hL79aAIbOEYcBMyaZspHa4PwAS4dPYmKdFPTMh3ULTtgk9rAPmM7AavfcwVcTazJNHitWs
PFgL4DAIHpBXwddnKgrcXRpq+R51B/Kc12LNs+tCpbPVRh+6enIAUaWyHiGMcMtQ5kyFS8C6Tie0
VrPnhJ6O6I40lNFMcCN/L60n5kEn6/WSxLvxRrvaYZGJF0IIiYzhn3ixy/xdaj1b1TvgpSlI8sD5
jUgDKKDtVjFJe1zYwlcuAoQwHhuGGxmHC4GXmmZk4ZphP1UJNuSTVpbMqLAIPcn4aUOTrvMhvkSl
0XOXqjf4qWGIKRvEnxjpMFMWZbGMlEvYP5/QK4HMAUEArPA84HCRLSDPl+tPvWTnX6oL12jtTgUG
2eKpLC1miV8Lb/fpx4JwnPxctQXAydAKZoEmxoBf7Md3dMBBTQipTzNCoGCqDkCMKYGSPMSNssvs
fkA4AEHujzMPohWraUGqM4awt6mwtulgHwtefg9Czvu5aUOHvQRcKZ3+mH7GcokdfKAkuTvqd38M
tZUShh8M0MHYZcl9Wm4GJB0OTgQyM+3pySx2NIh+3aPUrhh51Hw+M+mtYFUS/AcEVxYaO8pStLwP
rSl4K+6PkH3wwg4vraIMvn6FQcu32KozRR1gEQG7lC+/qnOfmQHJBMpTFPvx4HEa2lEBDOWhdAV4
zJFhR6reQfQHTz82U3Nt3SGZdtnTFXiqz3qCXX5FRkFkez77LiJb320pNSPj2KXUSbCwheA1ZNT9
FmL3DGuqyj3knJFOykpiknu0zehIT2Olf4U9q/o9Sw2WJ3YBOy02DpCF7oM5Uz6SR00+GSGYNtWn
1P6uVu3HW/Lglf/ZQ7nsnNyciKG2jYq3BL3205o9XRPBMubGABRg3lsNaQyn6aY7A9CjU+OPo1yA
V3j6Udf72oAlsB/RyC12gTtcGsrno0h4IFk5z5v2YLSwp/j5TYdDEdWf1yzISFn/AC1JwWw58tvG
ic+xWZ8CjyZVq6scehsR1Br1RQ6J2F93E9zYGI5NiPPVVgQdFtH8dTD8FoyCmwTWkm61+WrfNTBf
CcqNmcolbiGvUt+ZIxFC9s9akzJQWN2ZaR8RK5JbFV8OpH8mz71+aYTkgIZNPm3kOLIuFcnMppe3
yR793BpCaWgmzCldL4h+8M9aBbcJEPI+qceugBjH1eBiKPZlMUN0HhgHg0nx7nriI21spfJWTzRg
TCM8Y2x4H5ZfDoJuPG6rM0hhzuQ+gjFUOKz+IaSrdIWIPWIj19vgIHHnvfYYejBp2OP6aq5hh7Ia
mMTz9oGE7Q6k8q7LXL9x8qFgpBCi2vorDCUVFY58nCKgl5QW7d/+A3VoqwCtsRWTTCBk4RxlFRDt
eRifWs5wpdcOmVSb1J+00qXsTpEjjwlcWk5LF2Nc1xOA87DWWG53EIUDR6B7PcM7wrwvB0vH4ikf
g/OUSANANazn9JInPuwYfE4TZWMG92hEGwFsljHN4OvTjjsppgd4MXgHoxvsI/Aj7Ladf87hXD1P
df500rd8C5Wl1GVPx4ifQl0z4Tyd3Gp7PGzIEf/uu9HbxZyQjVf+20Yx2ZamMmLnUMrQfVykgwc0
DDtitj2cTMdGHWiQYvPdCjphqMrPbmtGoRkoyvMA+JGQKQxkgdpZqRZdYSDo0spMC1RFe28DNA8X
wMJXiN2PDv94+QsxVzkHdVpeEgtwIKx6Vd3Kgle8bCSYLS7kmnR7rZzoGw1VPtjxOBXoctl4xoJs
AiHEcnnyI99BIlSQEkNh19MpCsTZkQv9WtHy/Uk4GkmLGOAU50JOPlAu5hlZNA1A2MZJNN2/vTef
xhXytQdRYUI+dB5kFrSpnsKOekybYotoykj0wo+zVLX+JP+tU4kHT4bxmt/1FGYjVPzZzNaRNy5+
ZENR/Nm/FanwtuF5jD1RARveyzbgveaIhW4s/2cWKCc6vuDMuKUYNEER9n4IYBdZUQayHG/szlkK
9uJjUFVDXuMMEzlb4pFoBaSffX3tqPr4e4bYiL8yEsTbjGxIPOihnMCgyisxLQZCOHTm26fE9rUd
PBRATBiJY1eJ1VdyrN4Jc9PPyM7bGAGXqBtPz8JX9/vxq/M6dSfuImiHbGwilxDjPPe6+S9488/J
Zq1C0ErhEFIlIVx4KXgdSQviCGUlIX5L7Zml3uYNiwQ2v/clg42XiCKJinolcWG4RKqHXnQt2R+O
hEXSHeug0eCvjQsBti7cDzar46xtBegIzLvOU/MTfewYW2eU+sUohVAY/DZwZa58rD1aEzIW9Oip
Fr/i7gbWpQ9ozQM2o4GIHsPNtli6oBVZLiS84pKVi4aRNk5PFeubCwL3Ev0bK65ZkPWbEgUMpZLh
SYPFUSaFcIW/fFmJ16WKQS+sOWCYE7qPPBqAlP4kHQLvO6i8Ijh1ZiML92kpEX4gTIcaWVje59jO
/Tzz0+WLp7Sa53/h3d9/zgXkpSwQsdvmZf7Ya9CMoVppRh+23sPjgxgm4G7CJgCWf0CiVX+dxsZp
MlGgUD9RAsGtV+gkPX7oInNV86pJmgY9HzajlEFFx01AC6vzBj3imrgpfUE9ahNHzVNouaeeRAyS
xuVcV16NbOlAomBm2G0RzhZLMuyH3XAs+/2b6WfW6JYIfmoMsKGlO+QIcTTLWqim7DYl7Ux0brGY
slGXWfZbzZ8bHUUloSDcrcpOjXAjR6YH9Np87xnpjj/ASTbR5cKrbCgHIYIh7/jT09GOsS7I05pg
5uotpoMpkKSUppDM7NKPBT49V+VLI4R4RYSCWqbvD9AvgiX2LgwjJAzRTsHVivaaLaPZ7gdvG+Lu
Xt4n+hGxT7Fpx71N6w9QgUksrp93gre0yka5pR4pJUDOO23f5P262Yloarb4wjDgFhXMBP4BkNRm
yMYZaayVWdEqwrffUWfER0TfDbQ/tT+fnWsKXek+d/jpQi2wBAzevUZprSleqcMQfkWy88nBiWqx
T2NXTAsoqeZU3rFH2Mrd4txdJnRmyawHHJcz3USPEu4ISWwcmNMmhhegpEs0xkFjLbIEELFBvmWX
EL0BNlyJyam3hN9Hj7DLdh3K/Fp5Pdm/DV09dZEbpxV+ZMVS6ouxZ0XWl9rAYYQMqmZ8uI6ccPYx
c9jNCHG1sQCczLx0WCKs0ebrMIqfjqLuwj7oY1nPd1y2uhGi0LBTBnISpuqnEZeVwwRab5vFoTpw
0WbGDXZ0C34OmQvKQh+OzsEKhD4gLhyegV/seLzp/YKZ5SEyb3tTjCnYRyXTc8e5AB1cl+CqUuIP
x7aYKiEhqTlVx9pHD1ImXtl/VuT7arW2B35UCLYs9ugKdtTt0pjkp1TmnnNNYcB2h6RvvmOEUW92
APxcRvjyu4sHNSxn5vlLbFYHJ0nKHEAHl+SjPOk997reAmzGwfLPpFvDQnSqBJ85KDOuMMpqZ9Fa
Q+k8K5XOhrcL6li2PYIOTyrd8h7pQRnQPo/DIN8tERMRaDBlXvGEv8CO0DsgMKSeXypHHrCiIa91
AdG5oHG/BZkDTkaBe2OLdkoVBUBd7wTshgAKH0m28BglB4v7QiTm2a4paSOtVRU2bkIzhkTr1mdu
7P/NKYX3j1ZZOmHt2tUQqeqUV8UaJLHjlNHdOeTrgkDpSBYrMrBOutxgCLvrnOArHT5Ti6EabSLn
VOf7Z7/EfBvYv4OWi4GZCL0Hp78z8H0GYSYwEZxd8ilanwJ41lCXvFMOBxfCOP91xqQi6UNI9nmh
ERXE3jqPFAXuSAlyIyylqo6nIHZvIYRISnoZk976TSjxCtCgDq6+octNbhBK2QN/Qg5yHKGNatFM
N/rp1wsetxnBwR/beNk0l4JQqjOkeUPXd9j/EdLMy68ACu8t8s8jAUnm5LBdHUBnSs/bmvMcA3H9
5wr0IaiTvy+JNnPmoZhn9wt2SqP4Uj5MeCutd9r0/F2gpXH7W6VoL5rdM3+z0nySTEet5EsOnxGx
HcPKozHBeWdK7JuYfQC4mqTsAeUTWAn/jINtxclN2ThAACe98kAlKNgB79elA9+H25QVal6g+8YO
7F0KO3xselT7uW02hWcquGUAPRH6Ofo5AiVW5YuZWnls3tNqRSlugjTWDyE16mDpGMXiJK0OaVsA
zuaFWsSeIj4HFzX+epaFZ2uwTR50YUc7POGjeZR2euHMQ95BKwy5PqLJ/IKQJUYPc3lxi6CdDkbB
UREEf1E2+9P0cIzyuSV8zdrXur6/MznNjA49ZEIlMSYdVJ95mPCg7m5JvG3B1TVuVAnif5qoEMOt
AaDIrBYj0G7d1FHC0RNJdPg8S7KkdSD8jacXe+MgEJijl6T+0r9KLWMee6GmFMXmrPuGzXtAEOvx
96kjQu620vCr3F74rHvyMdRbhOh/R9Nw7oPrsbeRW8pFkYLq+oAQiCu4F9BJu8ALo7ZzBx40s/e1
ELCHOEQIYonE7BL/pqnYNYhLSH/FGdI7q3KtWm07E5O4uf6cGWaG672J+es84T/YC0JNT5666Wp0
etEggU2lb6ROq4D6M9Lb6PixyQCFdX4beU6Fy+tU7TsjVjgHufiSaFiQbtS859YSfpUMtT3DE0kd
/NxwfgrO2dZ7sUmoovuMA7bmmakvmso4P4PSM1XEfdMtvpc5G02ZPg9iRIYk3jd8xx28e52rwZxj
67/GZHA6CgjzgW+MhGTz9J+KF1BSA2k6sFugu+A6MgyfUehKTiCEcM14H3DsEK4vpxMzwoW5ZnWe
nnFkRPUoRP/N+qBP4sw9Sv/H2vuW7pWSBi1ty/VjuyLA4pCx34J4IVuZqDPqMwkYB/RaYhpw198U
TVDL9dHzBfBdQ2yDCNYUE6BLMupvKb6X1x7EZej87WP4zDg3FUEOWIWVeNQJZZYa2NcYEaNQ3zES
3AZ3kYodrdeWuh9o227X+9Ey6xKez8Ib/isFLG/tRuYPLfsNMtWb4mUZKuye2GWWGyekW8ATRUfc
lc7If6xh0MkTRQid0QGH6XOkrQD7VFF1ly8CAVf41Xi8KfPLbI1vYOEGMnennsFW+KNKYAQ1wvKz
/bK/jD5mVlN7CCYGx8Uudsw+DEYnrWdAIkCIEvgiH2WrhPHvFoJUiu3+ULfJ0HdExxgmLnFeq+WL
ko5REDiB3OolwltK0NTvrezzT2OI7XLG32gR93lVWloME8000EY6bQL+IbwCjoVMQqL3DVwQfo8a
LAGli4gQ8JOR/lqFrmGN9pXJqx7btGltzHwMKyYa7+YKlDwh8RrAV0yOafPEaBai+wrF/gwPev+d
AsWLilTzV188d9xWlvdLuQB6lX4qHnoDfn8Hjbk6bls5xc3SA3m9pQRZkE8j1N52mq9VYmlBtox3
31z4M0nyNnf7EhNU96xNxsyroFJNz6Sci1mZILRqOFmfXEZxrWOT7QGqY2lbKQ48Z5pm9kyqtL+9
9LRg3kz4sZPWdNqE4K/vT85CxOZc2W+sNjsHpZ+W1KIr1Y+7tTo5T4Av2BV4Qemz6ucZsDRwZXnP
yXxVpxCx2/Q7KCvkP+MjD9gVrVNUGbWNi1cpHqTmCENHadomAn3F+iexVXGwDe1ISN2MIFqA279d
f27+W1BhzR5jhvDRXe48uc7dwrnNLEJ2pgUNcxG/AYys0pB986X3naYKK4jQAJnnDriBkleyanTA
rWtcKXacVCQ/isTTAzr9qqkG+S3Lh7a4YR2aND+t4L/k6fzQ7aV6FTf+psLZM1LV9t6TpBKPiG6Z
yTBqHmoXpg5XR9uKymW8gfP6AU11edD0e8z/OJgJGPfK/m8QTkMNdaVuiZf1buoRRrKBCy/9fU9w
1u1Sk6SsH0Nj0Uu7y4WokcKKnVBSXBkluMXI8hNV+ipsTF61PyieUuxv933GXjhxLAoYOJg4goYs
EE8gqr92XSWtOnZSYWmo+Nz4gv4W+ghr1B/DZy3++hwNZR8sjVY0ezI1WpbACJacFt14lNI5QHei
y/2BBwwcRPKpXkv+3xg2IToWbm9OR34Mhg/CJIuYjlZPEwEHR3uX945dsE3ECHNmADSlIWOsPtGu
sXaQQrCCIRHxsPSSDOZ+uTp6aW/B2KH+6Q5A23r8PpkwR/eKvNZFuM9jJev/45VI6UM2guF5QTxf
fKqvl7lF1d1Sj7pdYqochs5lAb3dST/wInI3pCbT0dGMPB2uCMKD6jxCoiQXNIBoojiImYTiyl09
KpxKsJ+eAHNEbrUX+eWPLpmvLTi2vaHi5y0UQVmBlomyWzbElxkRguVjuQt4cvJSKsvtsRC+2zFj
2K+o2wNep6OP1cmMNaEfBbZSYGwZJCu6vM5EaB1LxSJ1ghhP6UxU6rA8gkhYqkJaWC9Hd7Ijkx3a
Yk8CSg+V4M0KCJfvPrLo274dtfzF5uuXGjapQI7ujv4sgQduHCbmQNmYPQSQC5q5Aae/Ksv6pfx3
GhMTJKpTRqCC7gj/D1aK91pgaxgrip20fKKPpXjVheNWeCGoK9omwzBUJ3QPJms4AaReYs2TKlVA
zmuAqKYkZGXBkKEqndeZ0pcbqX0HnMeaqiqFE3O1oGIhq13ug3BOb3QUtre9p5Wk3LM2A5dQNpIC
xV3NoCGBalumIKCttyEqYKV7lbNY1WGtwlL1yvqaOj/pv1azbY6mtyyu+l4cPDdHs2APcTk3NJFL
SlH8HU28UAri4uaNfuB8OvQHfl8aeWGjihutqAsOVlm6ZMI06tRqjfbpleVt3LdE206VUbiIy4X4
9T5cKx1T3IMHxKAR1n0zWVIDvkFmUdNI8rs3MQlX4To4GcThdtMRnQUIO/oeh3AlTHwyd0suip77
TiI9uQ+mIE55HBL8KKRFKxzcc83xfc7BwK8pAGUB8ShBffOd/EKS5ENN/OiNBZlvwYbJ0qxgjFrl
wbx1M33rqelXPkhXboL/Irxqtj7jzIETPg7ECXVldf76QUKwkF5SO0ywX+4sMDUhtvtx99QhYg9K
EvSjRdh5vbTuQqdT5siBjastU0A5F8QQKBNhHENddX54/heKW6+JoC8xtjlxrPiBUIgywy/BRRCR
cmcB9P1QzOsvjQLAOzZapC5exl3TGTFbgSMAdMyL9tB1v1L0RZ0/IqhYFPuWv2MIZIBB3icC2t2m
8iC4f0fyH0xyMG784hlumAnjxCBKaBv27YfWbtTIFoOIvHwV0RSgaKZ0FZsbloEgDSpGKJMedCIh
V+c4nBeqSiFaClmwW9sokO5YZlhgWQ5r5pws+DwZJKVwQYcc+g+xK9McLWknvQ3fjHtlEv6/y8ks
DGM2KXgnyssHYc1G9zG1ZKVk733+SYPSBXSPGQPsCgDC3m72flN2WV0cKqgBYZpWvlhG3Eh4DjrN
GQM37qz3f5v/pMlNCkErvODnK6pzAkN6POZavBQvnTqboMItC1DuCDatVBu2BJ0FZE0NHGwJ+MIe
/5a8BOTr37EJyEDRANW98k/77CyBtTaK54syoG/Mjm2S0AJt5/9MBAAIcKLdp9GQ0TsGcnlWTvHC
RYTCzqNFRD3r23KISaElx0Zkbzr2I0+rszyZbwlIlTpRyeIlbKLJMNvUNp1wVCElWJsQmodgLSYt
3jw+57zjItBJ172nlPFW1AdsJ0zWzP5gDM7xRX5kodyAyYYrRMuN1Si06KJB8B2qPwl8K2Lq2Awr
7r2V8IDNA27pCyX2rDYwlKBRVFPb/8YFDhmNzbDGHQv2RcT0dU0IUupy98+IkGo1sEE/Kyufqe+t
TLOR7Qo/ietAm78n7vZcjreKu90KqsCh9vd38qBnNHhmNZVFEGiGzRu0Cly0iosPEwFf0k2U2gcY
+aziDsGkm0p6OSVo01sR2ioTAPlTvQJXrjXzy9bxj+hukO9yRTejRr8ZeGfHi2xFoCguyMm4uBjK
KmxEu/ObecBMbX1HLqCoIPrHkJtCzi6iJfwTp+n38n+DkVTm8nlJYfm3KTa8zgX1o7KIjUk4f8zq
jgkWRkFK6khxCmb02GJY1MzDs5cG+slbBpy3qpIgbmIdnVX0+wv+8RFWzXrSnkzNqV+2ccFn3JyB
Ac77eGDnZd/sgBWbO2/76MXyFtEwSwA730O7Jy0cBurvM3w3MGijqsA4Xqz6bXQCSdsO9SUe8N5c
QmOydYBUPgjmjhXpYQFMlBR5Qbgu3vtCtgcpmRNr+c7Ey2IZpFmrfuUImVq/1fuQZ6oEWh4npr4X
3oklEzkIfHE2mbDcyrySKEaTLZnSLzn65QoLX/nu0DbmeYd0RIDASUJjCL6fmn3inCj9sqme2pyh
lS+O8W3XTwiWrJGGnbl7jOeNZVLPw/7tTeP8L+HEdkytRDSSfutpkAb76LHjACHRN1mnpIAreed3
xcThF9kzTP+VmNaygywXjwDyz/KYxZUgkDYPl7Jh02MFxysofQF9R7dGY4RUXI7pE5qMngTFM743
wGap2uooK6UI+qWaZWoPJzKWqGT4nb4YYFhze/8bSl/neM2TaLtvfPg9nhb95cXMZKzKKxBTkkCk
tf2x+mNO1nVcJ9L/5fJr10ZfhXGdo5IdLhJ/LRExSDc6A4e7CvB1ZFQqpNsrxRn4s1J7k28IJGtQ
vuvtl4XKVmHKx3LTj0KQ+8Jmt2dOX2J0KNWWkdzOEjQ0NidJgOaLkwnwdw/ums3+IRR1kI9q6X1p
jxaW/xAfZBjTvZ2wUdrZ9ZiNpVaUOsFhPF8ePWJsi6CFpWzewFqmwrlN+SratcG3ECVJhiZ7E+vL
LwaJ1lBHt+Qri64EAl0sY37umGNRP4EfP8qjwRkwX4ui//2A9cH4GdGH0hpuNyrP1MkuLiakRJT4
VmpMRyxJLVSixGLwX8NdlV2XQXiibl7HNbfrvTe2FQ7SHZ6cAmBJsU61oleAkAQ77q6s/xxa+z6s
9yDBz6i0Db5uckgA4fz8MrFTsnKeglE7Sq0WbKiu2HCmBSiIjdm3BvbM8jal1T9Dh3XZgH+3OIdp
6oqlrTukgZvM9oiDyAJ04sY050f5VDopgEp3KE2HBKB621On7YMS0tA4lG15x6vYcInXfEz8P3LW
cackgcISbgImMPqKLpGcc3hyetbgNXlND4jUhzK9jugykpOADfN6ulQzDSMTPQfuLDY+TYcMTx1d
CLo9O6fdSW49BGnQf+gV2IPa4ooSfR6di70c9IjndSWSp22mcjzKp1XAXbijH4nqikn1B4Tlfnqo
1/W9yJ4AJ66MDmvmNtpRWCoLnAqXDMzUuAkADzheA9H+6QwAumXOkT33evUhpiq5+JkdY30FO5w6
uj7SWf4oyZorKkt5J7XHfo8QOF31LVGASW5Iu+cDsapkmhKijG9vXRLp5rw9ezUSYKzrO74/+J0h
C/+zDvFlkWgLWRonl9bm6FR+bRBVx7l4njsppBvJPGosTGCHaFg7U10ShiVwxTRWeS6zW9OtGQ2f
saktjpNs57u5rEMkDhEoeBPBAoVHXH7502StF/MVGhSt/7PJMU+b0TIC8IRlaCar2d5fFxNxRcX2
4GejQQipKXx+WcJyf92cKp2bPGaaxsSGJDhdNedv0MfeuWfyM2A5dov/p+1oIS0G54ZggAH6damn
cbeWzxuklB/I6guzy7S8H8haoHo0y3/SCA5DdM4Fr//vVsME2UsxPSOdd8ToS6vQHu+5y/nLmR6V
bCxdZ04Kk3XYVJ1zBkhQvV2bbBzCTNcdNKpWLgiom8aeWkxwLlDq6GfvZ9OiEjs7KL+IPJsAQWRq
D38wisY03yTbGUMKXRWXay0kuaU1q8w77Go0yia2xeON1dUUYwBS9G/+6kWKn+XvOqG5tQ7dLICT
NfiOLKUp3khdkvaI0Z3riZxKR15CHeM/p/9stu3ZekBCfUrD97GZLCqrS+sfdNxNSsOod24nO/s4
8ry3vMRwG8Mdzx872E2qPWa1H9nWCsx4q/CSV8sqM2Nmi55JcCE0qwXc8Fqr1GzVDhQ/Co4RcgjF
QgZiu+X6kHf6w99+qGTAGbfK7jF4BZRXUKmkW7bdhtqXPiSrbGIiRGN0He2qIA/QDbSoY7YEW64x
q5OG+R9J6hypHqItyALjr/+mrT4wNDs1YZeV+aoUOus7ryhGJRo3qKDT+4utP9ysbfgruvZ4IhlT
lTZl6benwCxVvfaHsw60RJSXVG6gZiatTbq33Gk3sXtGKeRhHNHzCK+HiKLK/UpTAp2oh70ctPYY
0ThJznKZ8ozzphAkDfI0X9qk2YvM68OTxWw6w3Z2e7gKlVZZ2HORtRc8qPiz3Ii8483Rp1OmJw41
39/K8HP4XLI8fbLMqMSEZptbV4GsJYZyGCjOr7r47h6e5GlBQtpsVNkx4NNkYi3ezpVrkGg9lBPW
hXvqptwaSUtIknDJqODkW8lgsjpUVlU2hy2qp9mh/M7FRPaK2N0kHq3SFayjmy6qN+HmvlaLPe/G
KgDgRnVEBqDS+CXaLUY/Qh2o60BahMWYFg83a03IiSgClK3KqZ2kppEEn3Bs1JXWsUdnVv/J5Lvt
4O+21N8sfEaq5GGLqR5p9cb1hBIjrfJvj2hCN5/HicmulPL9Vh7iF3XOar5vjNgFMzZGLZuN//mk
U2JTITNqGYPLGGEqEdNrCE1nRngcZ3N61KuKYPc0ZfIDHRSxweBbgoBMy5xRjf6iCMEosYr3cPWS
G9U+JpOjRsiNLxZWwO8BpKZP9+ratsTKeJJH1rpowp5jFIC60/YIunQWf3l6FclMCxORHPja0WwV
ypdUDO7hFcnqFtcODviCNT7EstQ4UfdyF9ZmYrKiiy23u0zWEs9S+gUGqwOHrMH7Jwp9rReX2L94
zDmMJbVHDte9Mo0yGK0x+yKUkc1K5iKGBVQLgEglG8E4wDhFtOChiuIJRqJI9bV/ExYrEewsiq59
deEcjv1oM7+/W+KMzAVFSA63zsh69rcYVr6mYXBxB8DUS6IpLiWsaNfxFXZHKVJ07uH4xF3FESTj
uvXV8dbYSh2eKKDVxEDt/EYSEtV4u3qJbnWDFPdUQu3TPHa3Cc1CVZ0/0R8AjyK+F3wB3iIVWYie
5v+YNQ2QJOH7s8l91kEWKdAbhyKSJPDJSzDlPLF2WPcwKdCtSskE+nneGljYDIXSrsu6hUPNgbfB
MJUoJBi+I1Ngco9qc5vF/mGeN/47dBLuaBA755zz1bY1ZBi+3lzqJLt/uMas0Imww6QxH9AbV+P7
Kd6hxXl4nYzpmn5vORHzdOoSFo26c/I5TrIsfVUQd/rR45FBC7rhpoXNzshDrIHKyYdYFNQZhOn3
HC17y2YbicjrC0zBnIIQ0vZWI70tEfJqEIYonBupWjl+Rl4C96orCo4+QTU8gPtjrHNSVRv06GKh
B61AB4HB1scIfDBRUi453HPRMXXisyYkaVK7eV5hnFyLQZNLkqRagkATGQP8Lclt5mKO74zvmvGG
dEau63ARL9EqJ+bSmRlSjKOMV2wm34N84WcT4rZALqldmq2fRdU1JRJP6a8mmgrpX9F6UWxlFiy4
bOCO8PtolrKVUeq7M/XyXL/gd9TOF06/OfrNahFwhx1nzLh/OciMNHsH1+U79up3htndan9EkQ67
nvbLSeAhicPp5npJsDVkpVEvRt2zeLnObWMI7lrohPXIJsVq7YS4AfCNNozzwT6CwZ+Y+MkWBZPn
4zNvHgjulaweuh5SIrsLBgaLyWIS3CHFNyvLlKpXVIidnnqUWfPMhMRPCKbzF82cdE0RHlGn1xnB
gHDqShVrqf1cPBJ18leYFs6O4bIdHFNlM/WmFBQsTLJ2WfmPAvw4+x76M/s4AopkOOdErEUiuVgi
soxy4wyXEi2bVUUxTMml0WhmOtInErSjgzW1axC3LA0/ARSKM75TGNnAgsqK9nzM/EkxLPlQe/2u
9oBZBe7nxgqWti/44e69BcbLeIC7Eyh93xV6MqWtZgo7jrfQxK0vPmcOAzsMlmPXfwttS47ttk4y
4wogJiwld6uumM4dI2sd0PBoc/dJ9XtenMdtgFPdScqflV8kZjNC9gU6gkxCzghGZsBcJ225gBRL
69+sB6tb91efcR/k9wEB8v2vIQ0Vh1cmY/6fFHlHy4YS6X4glBeubWuHq5rX3HxQRzL69BRZwJKb
52I7xctR5nARpK5WMt9yPZnKaTkiIY5SnFdM/uiYZCnLoXO6iZO8lt+qKS2Ubd8CCTJKlxGLSEIk
zrtFL/3NuBTbzFnWvXlqVxMfJCuHUfJ6E+hWFiWW1FUN2Q9nxNDw78B8OyXh3GJc0yECo57ISBFh
xpj/0z2plFLKf2FC/GrvakHBI5Y1beNC2YF+Ig8TecogT43LLUX7w1/sr6iiF/cJaU6jD+Ebw/m7
s4xZbvIN6frVPlPjeemfXT9jM794Az+JeQWtXtAgfrlWTpJSzGTi4hdE/ymA7QZcsco/6DaHyIBV
0g4hIBSxwTH6rrWm50PIsdE9b8mRxC9RNd3PAEgN5rdpOrDaVaPD8PqzZjg93IyqPBgmE6EUZ2Zd
8yLrZZtMhXoxT1HWlFDwFOLtXJSuhUhzWkCBeuqEP6IeeoeEaTF7cxPQcJnlcmchhpOP6TBfmreI
fZLaeyVugvKfDrro7mmqa7GsKdHbo3fTup5V6KXwDrxpEpaESZzAClPMTUzkENgT0euLZKW5sWkk
/l98qk53MlcDp1bucBa9zE8BC2Mnd5lvSS6Dc2D0hmQEz1ctY2WuoTokLgO8LBRUNc6KEz6cVT37
9KNIU0beqiDYggiZLZ/wEr23t9PwilS2cZsyF5DCoIf05my5E35qzK7VxAzVsFW21e23stOrimQA
pdY+7BTokR1sl8rtZrUDGfeO20tT7HjFXUWDNDaX+F0X8k8lvCCw2wtd9Xw6ShM+qhgSQW1Ak+U8
9rd+A2xPKIwKXleKLempcwx4ThwgfJCheoa2efMEJGjJECFsYKfP47jGmuuOW3xThwisjsRtTcvA
XxkYVo/6eilqV2ybrVd+HsPqqDiYTEYFhAdaCSJP6NLjoNRxvlKFdQa9XHiqyKj6jeLoEDw6ShL2
HQ/ErllbTic7U0BZEVjPYfAUPpFEinViveLTOGpWmxmTvKoyzV4J5Tz3dmORjdkxWBH2+3kY/s/3
7rKB6qvsdrQgayZOTYERt49y5IKl5B5gTT++++h/x49ZQmvZmA7Y18mCxb25Mk2lN2KPU7hpQQcT
QYaP7QVvhwnEKHTxvEIj9AGrlwkTIJsiBe30WxdQhU9pmhcwHkuTxLmVyq/SvUeST/b48IaK186D
rh7VqxCeasiz7cFd7EA/VFxa+DfoPDO1IuEKIaC+f9KAy1jKT6OauQmucRxV2tZeshvWBXTOaMgR
GDMGjk+zcMPHSOcjOxO2ok37VD95Y35hF6jdVZ/JnGUVX9+Xij35+H4jis9i/DuLpzbyIK9fxZdj
7iuW3nNyYyXn8qI3WSINJ4H9iLA1lIK5jWX1XNm6Iv7Adx0Q1GKkCDRYgJ4b4/dE9zYHuD//cR53
Qo/SNSV5Q/OBD7KOsngaM1z0uq8AwjaKA4sDhdvxqHYjZ3ur1gzisMFnJMqNHkjx1aq1ckQE4omY
+K32unAOjvA370wK7dG8kfdhdqO2sTYgcsBYm+zwFI0lug9/KjLGLkeCILoY9PppfEkbb2EO0GNH
ia5Yw8bCjRNb1mzxA/VBkgBVN1QHAqgYrv7764o3wbFHaz9Zp9OzO1FVDUfRrp+YzX8U9xzMRUhK
Ub4bo3emRyHTfldjhx7pjmT9ZXsJWT6BTeacvsfhroL3KebjWmpo/9gjA1UAf4P2jUSYs1pr//my
4WSx9Ct5Q1OUaa/umWE23hRY1q+BJ1Pye3kEcOW7ALppoA4aMVR4dTBnSSa/DaywyrbEP4xZ/TQZ
GMkiVspFgabQXRS1XVjR9MIZjOxgA+SeP/LIfAd1WLdc6dmF+zrST0uB/2+cHAHeeTl6OABfpmgy
o/rPqYXav+UPvmMsRNxM7vyvFXeHjmMklZw9SBvop2iyPQr60LMSOeYDMksfyi0EXthD3MkQxNXK
BaAxDeNUtZGAp4oS9rKGy4inIsyk8sHNsY7iUec5p8zPh31O3AGYle6rg5Riwzc3QkCgBFRcySnC
U4N/IClg0ZXhkHwk8VqQsathPP8OXJRFvTOuDo1mL3j4Siivlo+uBP8MjOSWNV+2SRhbpNQYN7KS
m/SZuidCPc8C6XVoGMgdea42+JShuGiEXjipSP0Eyr5nNurZAfkODnKS11Isx/3aZvcUnGPagiYv
DoW89HbaNPN6RyCjQxRxIURJ3czAzYIY7qjU36J5/SSAOKd7EHRkjDHD39EqOhDVGs2IEN9YiIRZ
0eag9hETmGAN8m0550UkLJBxCk3ZqYlXwjuDCHfTkr6+ySkg3GckbmK6y4Zb83LDv0dttZPYzppF
q6FRlFoS5EhjDz1lNay2ZpGZUjfD+PXthC3q3VDbtFVu5fh6h4OeSlWh+oHfFWatIY68SgtCl886
KY7Q7vXpCQz12xaBRAW/3hngkFIMm+o7Eu5J/UM8dbkRWo9V8kpJkn+HvbogUupxe2zt+UvZsyRq
ajLfDnhTO1g9baOCtPmzpIToi3wcaZafiwC3pTMccNe2W4PuY/nr37Y2wW9UT9DEvMs+Hc+HVIL4
lcsROlbnApe+1MMBFJWXxzCQoHJtNtP05IaGbcDbpcfBVM/4TambzqasTQs0PrkBgUpgEc0UlD9A
Ph/xlTuJ5pJlEni3bimROcvbYlyqhRbliZ75elpChBAEshe3zUICrErqDLOW9B/CMYHqXh47LHtS
aAO9uVOpFNTSejxRmCQg0ZRL8u5jA6MqzdzjYjdRN7DfkiPcDuUwW3De2bwDSyh52eKQaWW3gXY1
OuJOas0Su9YE8yLZ8FwyAMpKw422s0QB9CNpsw5Kw70i9mz2fJ14KpaNijuRD6lEpk0Ymiz4kZk9
jwFYpEW23lI1Fzhw/Eqy3t6WlhUrKpaFhQ2W/6PZpXOSJeR6MEaevVuC6ViQy5jWdrpG4iWh4rO8
K1cStjtOw68BZCg5LrFr3kuUt30yss+/OeJdIh1LhpLcESmX8Dwemfy/106kJpkHK/0HbHwQY7gv
OXyjNC8WKCdiqjjenxSc06btIQau5jE4S2KpVkYz4pEXrdYIeBtLqzFHxHG6cJMi/NlJBHo+1i1O
mXp6IGN/zJLQ0P9M8ln0EC56XNPdF3kYeJoCXc8Ai3kVQhWlkwX/WMotNoOxrU9W2/A4ONBKcV6z
ENORECthKujlY04ZDbzvRyif3UcUk3cUIy53dwzal70SmAnNQU7MirW9AkjLkxj/FTUiRmdFp3Yz
ImcRqDsxUOriy+kgmDxe+74ExICHtpkh8rYqSb3kE37/k4aKQY3kedrShulfCOaS9bbIuwdvyiRd
Jwb/IT7T2ZkHN7Ifud8fYq2KEiUrDOEg8iqJX7O488ZaVNJ+eImk632oe2hcRJxLNESXWDhbEyWM
UomBYrXAiLdl5+HNY6vX4GM9weN4OB1Fz4xu5tIJwLuUjfTiSYUR0DQUZO89HoAp2j35FD8Wqt79
Q36860rmHdYuMt5w1KIpBzR78VqbTZzXhIvFIZecsjyzAvEsDLJPFLDkx53wTI196NnJRid76qfW
3Uzk+cPMct61lNELq8gU1ffwVuzdUz3x5w7gEjeK9TT38tpGF7NMwRHlTjCYUiPCr2MxfEeJ12hg
9NGt4HbZixtrS24SCzJDLROVfWVM2ElwWMeUglR9G1mXfawkjhbMgI6I824T1cHu47Twmtu8VC+x
Ppzhy+qbB6PwMlNavEQ0vWTggORfaWEYc+aF1MH1Jog/3lAfM2J4osC6ZGLa4Q5/+fsYZvkRE/rA
O3DbxyNrajiepNItE+mLKBM/gaWjZkb4AhmvVmW7JdVfaRmIalqLBvM1wrgTdPaPYEs6wnws4+RJ
zWeJrjoz7wQBAsihQNMwFr13yW2zuDPnoOzyprxRXYc/rf6siWO0wwUWL7HZfpNwvVInsQ40B72H
35+3MBIf8MyM1qzQE4CwA6ZW6LZRF5vztaFcp7LxQ5wcOq6e++ectTGE8/elax/NqyvXEAUrETP6
S15RbkoSgE0PMMco2c+agt4UFgstVn39qJrsJfqPZZ3X/bc7n2DxzbAscxJWr0Sbex0/4UPMHHTY
7vjWFcs7J3dTGd9nVmNe0vR38jvi31162tLOnKWCkPUD9ugq0NX9El8RcKpj4G1b0ORvrQLAOvY3
/AS4/2zWlwAWalWkmILDhQQh7ESJsEwNhFTqnnf5DYCt60Eoo5wsi7qKztepaEviteO5YEjC/0bJ
7pO7fExBMb08Mx2CqTXDF+j92/KCDieENuQKGq9V9nClEkmTfigLJKC1S2NNW1TnbRlC3uamNUPp
4HMkgASkAS8TKWYPAh65F5Am1A9VwhmV3715CISXyFIRI/RVQbNK73HKyE08n7IE2wEbP/9EDvt/
iOzrRs3JKjfV22PsGVUbos47Xsv+wjpUiQxa3Tp6vttsfGot/9sekwwQ+pVUwgUtvI9dULW0GRiz
Xs3m1xhYJp+qoAiFBVuxXwi730od5RSsGn/6tM35rnV5KGcpl04c9apmnao93WQscdU7it61CwUk
oj2TEQ4SfIXMZueQ5HkEl7qufNeRJ72WcCem9A0KaqnVq61vJoW7I8781MjJpEVZOHrVZ+ppjuUq
ZNqJxcHlnsDmnkDKVkZknmcbbIJwQenHGDyE04SKtN9SfqI9Tz7iaLzCS/Gmaye1+TKIKpaH8Y4q
t+VI96inoCCEX2xpTQgnJqPNBUCBrL3O4Xjv4gwgi+Y9+FwMSTadXBnVu4vU0R1mG0bqoojdvYzl
7ZKiUjOxcks2gdY0DK8kI+8+YlZpKKrX2YIKuhEFmr3jCJhtE4zVM3sJmnyDpL5l7tFaIjp2FXuI
edgpaBvMZerdY1oLaWTsNDYxdFs8xqbWhX+sfWdyNu7wKpyjk4Ek6/KoPjNWjH8v38yCtw2JjpqC
vGjH/fZdwmXKCwzXPxf7SEf8lKtl7NZKgAw9dzFvWWGXbIAVePvSMUw4ekT4Cp6seS60NZFe91IV
QqCU7HGRAnE/XKfSu5y8rjdvYcRSd/u9+VbMEtY3tLfvws8TsKKxuic53LOneWfk7yXBRqB69tBS
WUMVAxGsHjQw0GlMh4zEsNWBTMCNTt0LFz+J75ONTLNdDWxlhi9064qc/hGERrljBsQ1sRR/BqcU
UMmrnIeu43hGDKJwWRpi/BqA350/DqW2ao8XFnBW88P0PYgZCXf22RukBfDi2qEGf/whfBwF7yh1
of1u4KbwGXw2LY5fPqrieARjBWoR3GYuHyV+1LqBi1PZ0MfpTG0NGOShRv16C+3C2kgnrO35suiv
haGSiduSzv2jp1QaamBoKqZVlaLoANEp0bBIN4V9XvCaz5lbO3tXTijBULUXl07WkWC9wOyC/iHO
Z09UDhRULeF47ZE3d4XWT8kdVVSwhNUnkbsQiulW1gwsBNQOOqL3e3uP5a+WPT4ynXZ0VaBfDVVG
bOGyxwEK3/+Xdv+LDN/OeTYp1D/VrUztvLaRf7BLwYCx5Qot+29jLWj1jw5j+v+2yMLBGTPaRC58
1nC6xMOiQYpcCddoQ7S5ZZHHEmGTOKZEiwfKZ0P9p65Hb+EOMkhpUqPEA5RtGxYKqlA4Pu4YnfAe
4YQTR9B8bqMBvO6FssJwAYDB1MpoiVrKtfinbpUqCYTzVbtkYe7v0a2zbS6zzLs5tv3+bKceEMk2
u92gRTwcYt4dr6LbOt9hEFkZwxHnl272ZuK/DhFapsIH+bQVYVb0AY3GP6AyshF1cju4BThFVMx7
Hf4hF03Ndxy5xgcGyhUhw4P+E86zSH3F08G2dgxlI4VtaUBZIETqoRh9M8uwW5fRk/7eF7ih40zS
9uFox0JMy3VPsTfNPuLsTOanVkS/0PuzIikjUEwT1iRTe6T9Z8WaD32NUyTdeuIxwzcCDOz2mUQY
eyEjwvBbnvYcFJ862BVhHUjdG6PtMptt4Jl23trsjok2Rqv10nf6aEUgz3b7K+0J4Kx7y+HfTFRU
HI2v06RVxzrYm9rfBEFeyvyigTOt4/NA5x5gnW+JhLmzCev0XcysQrupi0Rr5EQ+2UJCIq0Vvenj
zUXdq/Hm1SLzeX8wZTB6T45M8Q6tQ/IfAEvq0cyuvaIYU9fdDoN7c/Jw2f0Nh+eNmSPDKGkzSkTE
7FLDoot6VqBQ6WRmSP4Hehba578MiYC1oVygc2oaav3cGFOgcPE2yqDdZ7M+EXFtHgjAW3cSBROt
gfrg4qWAzzXzSxmGUbo6PhLaT7nRsWWyx4CcvhQFimNYTnJkIBImcM1Ry7MnNM51YLOUCAPOThW6
8O0kF9qgmacMnzWNrFwkIlguS8moD4K9Cep55qOeUMTu0TtyCKQypCiWEDRjBrrm/aLaSwzoql4o
iImgewQpRrVKQokGvwY6LVwu/9hOilBp7Uo/2l5Qhd73l+QVguq12Qftt/GMI1REO+q1bAoOqfiC
1FhqvLpgLQG5Vq+mDoIlSHSofK5JLOKgIL6PweTq5nRtYQvDudQpevfHzjyzqaRX5BqMCrVw0a6P
YGuERleCSxQdgo3kn17Dhtp8K8nha8uRPkVrHIZjL7ypDmeZpbMlbgwsRhgGo8YvcSHJpWadfikC
3XuoPvfWTe7de7+jli1DghQr28w2tX3pp/vy6eDN8sYIrm9AqjUCRLo2rV9Gd9opF25+5wjMUBla
0zWZJAsFn85BRh69aRZFo+mElQpU3fIUMeHSy3gtydwZU/296XSe9C+x+EhnSNUR8ql9t0TJs4gl
6DgPjcPb4GIUSpX/MJ3HiFKDK/1z62AZN2rFLovyj8jOV9LYWhULZDOK0TBxtff1uW72uOe8fX5l
7aAb/B387Dg0eUkxxsc3cFCtY9Vf8r5qUfi+gsSRIlA9de/6e5z3yASqeBlkZsKsyzuW/4en3k0r
A2/fUlDY5aOGP0nlzOTGbutwF43fvqeO1AVB7uKecLQ/j98d+NizrZmqYlI9vBT03x+tltqA/dnE
VW31BJJOOiZHPQuE6UuP0W+OjZoZcLI/kwp0w/pWprhd0ozUnGefT62xUchZ2MPSYvr/HUVhpLng
s/vrNAMD8Y/LjqcGC57s4gxZBz8zmVx4GBsHp6PWgAM/Tt5wpGe2yabhXoz3tc+4hwmVqXlD8Hdu
sP/ha5Qs5UTaskrVtlE2HYLayh7iWe0Ocgv9PpHVA1P6wEQYAAAQHc80UQWYttuxCabDFS5CXZMB
0nhKabadZLcoyslnbExdEcmGM/b83ScUHGuTrLiMlvq2HoEssWpTqrcjFKDV2D8b4SplfN1OTEvP
DS6yddpOpFoCi2feD8uZbZfdEpBKqMCgooCZWw1isyYTKZoW813+C3GUNv8LIjOBm57+ysvcUqs7
hFmOBgRVIR5JZc17sTZSuHjp1t2DHX1gwoCRhDHgqrGYpXD1QUNb0qwXrqZeITQKdfD0HS72rXTi
755lN0SXpj6L0SCUSgQvBK+AVek5XxYMqVlUwKaV9rwd9DS/0Ea5p4l1HSqAPdFU6GPSGhr7LLfP
wtUR1/NOc+XXS0ygNQ5MhyNJ/npaF55ivI3s+CR8/GIiNvT1nJWqVMfuzDFNe6nw+BCbOMyBk5QB
rLlq5dyc07xfmy0COr0tINVfT9+tBqcK8oiBiq0p8FHR8cWRJRzXuNzFAVemKJejNzqM0M5Rdn2E
tyFwerT3wawlVl5UkParDf5ptS99+JUZPUGGnqOPkv3JnK5JDmP9zUHB316hYH6ZIyYnfgE7X22M
Fdv2sYg8TygzWf9UB260B2cmbrkgw0h4C4EOnGcMpyB1IEEqgKpZsDuHF1iwXaY71+E9NzMS/i5b
cPoUaMz9BasO/HdGuEn02Sy9Qy4LbqMopSKMAfMgcarA3qgJmvRT8iOw5ed52Fdhs/Kl1gF7xSNf
v8CTB/LOOkNcieR/7vPF7MCB5hpQzyYCE+NEqAb6xdfsG/khUiXx7kdQj4VmOjM6WAYtuEcH8ZUo
AycLjZzX/5QZnDAYNZpgSX30Tw5WXK5y1Ugn7coq10fuB0lvhMc+Ji/SK+elB4LHi6XoYgD3ewNK
NpdxdgSI+zfCRoSiDaliC6htgYuNfeXcJ3+rrskwuO7OJF3Oh+na3DuuPMk3LZckZ17ZGlSeAith
E/oX2ZIkHfMZiwDqJefF2EnjgM5WFps88dhc4AIdbAFAjDRnzG6hZWm5VJ+gPpvBqigFWhcPUrmr
h/Tneinq7HvjFqWU0YhY+hjXx5pcZnwKVO5aOHvGkYgbADatQIfWTI7/3Ho1UmKhmuDlIzDDVQMw
fIUfN3tJn+ecl1BYifMKWZxlx+zUZtltIApTMsF6enHcKQL4jKAj/d/gYnsdbvOzEckoO46uBdkW
PZ78OQYuV7ZaKndoS0yaDwm6cTGvfvPDMLJuyskK5+ib9DllqqZXtCa9YJv0ntHo+QWg1dGN7BL5
KhbQFgnXOw0SDVJgc1f3L33TxY5d/akPPmuSjnVrrxXlj133VuUmUvZvCiwfZERNLZsUtUJVtYRR
YeyK4AFnHoSHlbZ7VzUrumRx9Z8cXCk1+Pw4CzNfhNaA8wG5Kq2Ds4LiSL4QRXhXeMUCDHmYXr4P
QcjLkxt0RASw6zwNaeSmYPiBWex17Sm0reCQrGMGItuti3KL0m3YURdT7gwYdmNUcklfpgMaCnIt
WTKUjQcI2RCmGckOHY4vIahdQhb1pZtduXzuoInbzTatzlsMmxxZCXQfC62ECdok4BNyKQP0Xfkm
nsEoiO2RZu51CCpogzp2avbnyBwCOlPa0TVNBaqnm9kmMtzCOoiqs56WnwdLVmIeY5CO+Jm3Fakb
lj8hhEAD6A4hvFieA5UVDRg/YzylTFV1T6GCdqIp1wc6VXHJ5NhGL6jebK4WGtIX0PAVooKu2Qw7
JhflrfLSSU5xL5B3jqEi8KRmXwkgzxVkJ+MmzkvPQlLUSlkr3ZFJpi/rKNaUHtWoChmDKs1hDQcA
Hh28vxTGz0UCuiLNEAQNC2rd+qobQN0TA7Gok0QZ6iwIoyO2y9yUd7TY3xLiy003S9dQqdRwHiCd
z5ZrYDKWJrzjN2+9Ih0OQB+0R/tmXN21tE5PfnZugeTTPL1loWwef3qGwBtghaVAmCp4y5Z8ZVzm
k/P1Dv9vGi8IAeOfTVuG8HSOzBEhZRxDBS1NXwqzMa15UlHZu4i5itlBLdmiPozrnNBg46qihN51
STiztuQKQfm3Ow1FbgwTXeer4PEgfCI8r+CH+cvOUNJvYz+OfaFawrW8wXS4KUnPSYvXH4U27xbc
3W57eutYgZjhWY1CQemrhknfEZxEFTSoZjVksgct0Tq7KUS4hlAzebgoXyfe4xggEGl9W8MBIrsl
83u+E7KyIzQrggpnumlSZpKUzavKsQelg3OMExmcIIK3WoMFS/FAxjG9jQ8Yc87QiK3OMiquE4Fd
xxb9l1ICXScTYS6fdQQxv4l9aC7/kGM7CAlWf5SYNsRJwNvpcYBX/Lvlw0I6gV5VUEaz/PsN0nND
KGUf6K/cWDw+I2bYW7haEEydxT4msjfiZH3ehBzVi/t547gkRan7PXyIdbm9e/pkZiIhLYm+sMIi
+dsdv4GiUWe95tDqIMHsIqFFO68FOuCaQYF5a8mTAcR7R++Ya55cufVRUAxrFc8HbCBmpPNJdisu
F2rWGgFWwjjQD3TJHLrtKFh21qQz/PyuTA1YK7VECqRZMPMrWHIAgaI/MPihTX3+azihgrkF+hiA
dq6863QhOEB9kdWXFx4PAYYRfph4pfnriDylrmkfRnABIPpSD0FmkQU5TvMS8WZr0uczbR1UZF/H
Qj1FczlOfAm0CQhtVjYFjrpO5Ya2KtxOV6RqSxP9l5QmlkdOdBE2QVoEY0Hedvv3Il+naX4PPE2d
3/Ykyl8fSH1+NsGheqxCxtxG8hol1skemBOmV0qnBXeeEr26B1mcOfp9qf5prcbkb9WrXUxKmSF0
GOMvOA9X1YYOdfkAY87Vh6dSlrD0PBhPdPtHlb10qHUTAJz2JB8VSRSQt6McVzNEy6LGEQvSQ91x
2mEPIPDxM2aKYu+fo7ddXQ7KdMEN1/d5brEWSGeJIproLT15aaCSWTMJYfPBhPcJrOsfhQNnxjwf
QBCemaSF1sPtaWLp4G3ZmPA5CHZgL6Ww9KHpmWHCYMIeqbGz5njWZkn8QCGbjZpvE5cuVF5BEs8I
Xl2UgwDFGf1orcaRLyHvfhMksmCDl5iogyzCEH8N12AKX0U3OPH/GWNOMoGagPALzUGIDjkhCb/P
SoByNQv9y0p0NWIFoZ422XAjpayaF3U2/YcZKfLtfO5GaDDqpfH0HWUuadg39VFSn9BO3lk7IXTa
Dv9+INsCxnhTCKy1g6XTfToLn1F57L+/GTGLUThvTRiOgkkGY7OVqouvzGpvizpnq8HEzRMYFDef
e6XMhZ4SUmBdWxjWRdtYFPkvA23oGNfqaA2ygGRcQPwQGml7Ajny6jVDROae1/NEmUo78O4xnuk7
LPrICxFfWUt+e0aX8ujr7OUWp4rC95vOlbSrCc0/w6oDLHcngjAXZYROsYKy4LAMBhaSdni6Xt8P
1rPt3yvrrNwY8F2237LE82szQqOFEJI+uE0bEI2DaS4FnWgJBxvm/XHrt+SHHwdRDwEULK1nsTKU
cLhqK8dAy6mPoIYBtfErY6Ruyg/xt8qNc/WLSb6ZuLuuJnlBpzj0nPZf11I/1cJtFxCuv2WZupjs
u2xrMJVAz7RTsHDnrtq7qFngTRqtz3MYDQB6c6zLuWc60q/4Bs7pTqWeiuLXNEBhZyo4cfrDNV3s
HCUzXRMwhudp2q9tSIj9ljPtWvVpi0eWfPv1GKTTZYGkTxd3PsNt09o4i5UsrhQujxahQwDaANR9
CMbfIjPui4I+y3buC3f/Wef8wEVf0bNsytLep/8s/ROrG5cyXnLpy0RdLYq6oHl2Vq6pyC3J9zNv
o14yqoMF6YW95KXxvbo0TJ28gpSGTgdob6E8ERTYl6ExNRtuHrC6pdPAuc0DeeGyLB/T9pFmMJ30
9gYqHPJyDpHv9xxzGuqSxQtJIU2Ic8v6pmGQROudXydlDnL0JOUU40yWYMM6t/HLdMiuY2Co6oln
LiGSfhDOQ6PK7RZ6BkLIa5lNWAqLVNlQ9v/fbi9OgOaJapqrhXbZByE7Oq8nd4ZsKO2dZVCErjCU
B2/fTCB0KKaSFEozePmMKm/Pl1PrBv14cpuclpXpHHyiQZhL/D0Q6lkC/5QBFVQ3ZH+Z/BRNFWmz
A1JALa5Vz1X0WgjFbFPsRyYBK8WkyjaCKE9f3+r6u7b94S1IEkfOcPR+o1L+nQYSE6HtwQKAfVKF
FTcscuA17EOPFa6Hn1GpAO0tGPUmdshckWoMDG2wyGqE/1B+fLUB8ASrAsJmvUCB4debF+A6GAvP
/d1qNgjXMVVUJINOapst7IgZRl2n0wXYIYPMhk1CtqIADO6NbuclB6/0udtU81O4zA8bsFjFLT3V
DdPdbCjjxvnKdooa0Wr4NP/5g6+h5Ute0uMfYXj23ehNSqKoLQFqVvAezAiKubHw8LYSagQg5L7E
RhXApUOrKU/DyFpCXCCxKju6122QUR/JorfmHDJu+xulQmAHxznGlyqAAFEKI5hO4LLDdrElE9bK
28vktcp7sx7t0NewPer9AlU+UnD3RtzIcuq0dmIZ7K0E7DLe94XSUblbS2rulAi7bcLoGmsTVjj7
ekqjkTHQqvPO+I/GqP1hjvOQIjeJjHsIpOR5kicjjNiEsdCfztFu9DZ15h4y8axibmKmdiNjsKna
QxIIXHICsDlZTRS6zuHf61wA+YLAdRbdGWab/RCMFnU+xoeD5ZpaLXb/MFF7ggKSeXAhTZk5Yl2K
Xwwaqbm66zJH7YHTt++xFzR8nKCdcrGjPWPu8JRlusbwaJnL1oSgk3OwFbB9Y6hlI9yxBZV/CKNO
j4h1nUxZ925eXfOmEO60JkR3MhhzcjDYsTpWQ6f0ASbCbXf5ZThGFtVk7GGSG/ocrg691CSMi9bd
IUB6b1OSb+tnNoAkQ8NsO3uE3A60BwHYFM7LzB/Ph1+jrLtrUVymo0ArwS+7qJu2aj6Z+c9ysF35
aCI8Kgj7gsZ/ggrFT9e3XyigJObMhu1eyxwx6AFs6zhPN6sVG4zoEmzke/WxL1Qg4XHmr8FZP2qA
iXo3Utlq29Np9duZIMsaaCGjOqm2aAfktGqWq/gpdv6QB3i7WSKpK1LgE3PA54UEPm4gjc+0P5Az
RzmybEUYXPaZAVQJzINSQphx+NV006GGuWC/Ly2ZXeIlMJq1NfJq/74i92t/ym9UgEm0/f4o6lzn
strJKwQ8FSQ1AWifasNWAUjMBlwYGjFnlMdeCyEOgiWwQSXhaf3T0imnrJwkJLF2asiMmvX/ePUY
GsvNqHzXvQnFvQh5GHZGffub/OLwHOOhXfJkDHJqDdXLSP7lH2nRfcLr4hB3qqL6bPDjDHATmu2s
ZTTiSdxRy2LK6A31sA7gJoZcBd9nI0PKRWNt24TqXo1x9xA3s1SgXaRq6Oc+qsQNrIUORWKgltnv
tU2e760NTV73KhIfnEz6d21EAJBvIGNe2Eaea7fAiIkV4PmN2ivwzaz3zvG3iK2LAr8guYa+oi5U
Klo6TsMQ4CQHm7ot7lotp1URO/beFTES6tfnPRJKmSdVocaSAg331m2veKw+BauUHRld54HUBOqk
TqYmqB6ZSfmFfZwA6Vu6Ep4dgb6M+/Ey3wy1x9mkWYcV088Ip7Zpg/RflO4WM8svB6HUp6FDCDXV
HcvR0kFdZ42rwSbMWHDYRW590qXGYoi3VCRop7qQpX1dThrnwImhU/KcwozpfW354czs8hpzu9UB
OO5NY17luBZFhD0gMaW1OQlyfK1SyKtrHL4683tYIL6fWsyzbXLAJokpsjGNYVc+tRqMlrrL06aF
lJ+R8tlhRIBAW3vGYbANbbJOJCesa1tiX3z+GOZCioYo/7TeItwzh87K6ouMbLLskKq2mO0WoHgq
DSUNNsqX4uj3nz/61czZMnAUT/0yl1Ak/mKM2VDDgOJOqdrG44iuebAwy3TSpEXMauUcLS3SzAtn
9iCzjFmI6Z/mI9gZJ3KYTtO11R/986F2HR0eTjTwql7vdLbbgm5vpp3JmiW8HrBqzshJcl3d9EDc
ma5/WXJDdhKNHOV13nKZynwqDUh/PYDIPqIACVpWRWUhQKVXGjSZMNcy8bEd0c7g0r4bhX+jsXwO
8COTve9hBKwlTF/kNGsDTZmzXf/Wyzs35T3VD2DBOrZs/i8PstGe9cYo7OEVsF7AyBztktx8Ym+L
3vR779cbXbDo8BuP8NS4VeYOcb/dMHmhydVAn5WCHZcOTUfhzr+aOK5oJsKBfjlC7xeg//NvCuYI
cf6oAkDqHsXHM0xUdFeUJQuowuRfuEQlHgE9M4mB2DiPXdI8i9+0PKispACXvlPqy7YkIZqfrHh9
7z11BWDOxWreGmuqE3fPnWs/yJpScgvF9WHC1mjNJgCmrwOYO1NT/D45Nk/98o5jLwpk8fovQp95
MqmJMl5uNw3TlluuW7ZEo/UvaDUnTeZ1E+cV0oEw7rDXDdPgMD1dSkd1IGMEo7eo7QUyh5ccCvBB
NC7Q4YQ/IZ1mw9P5eoTq5oV8P4luJh1sAYOic0tQXx7cM6ReVtLdGyRJpbodWQFHOm5MkgA8K8Cq
ANtS/HpEFKqU+dt41J+h3d4LQ1rJGuevbMiiRd6+Kcq652hkyWHsdap0qj2knncugEbeKOI6eGUq
MAha/SiDe+Cs0Svb3XBsmtf5tWcWIt4mCa4pFsXJSLT53jXNHmlrTDwqXvr6cQsAGlVZYJ9a05Np
BoLBz96HCW3En18/q1XCnqN+UEZlJ7x7s/HfzHdJ8O3NFE5HHTNZXrFrhfzP2TIlCCvgH1tHlOCU
YGkSrEZps0fXpcKi/1g9aPIyaT3k5QyqF7sqbnCXpHhDuEpv4KvfgdcjxXGvuwJYG3o/KmeINQq8
d2QfrD8EjNbrUzML8ZdBhoxfDJDB6qvNeEQKg2Xtq+nU/BmaiBfV4wbB9Y6rgsnm1sNjSM+3Ijyb
NeYwvQTk3CMpbHxfSmk8bi8R0Do9MQV3Iu8W8zEWWWZZBWAISrxc6nrPcmqsWeNAi2HV6lV2GMnN
LFjuPpsI3bldSkTHDTwwV3bklW4HthfzI6s9K3l4/IGZckTHxE1f8XK6PQB7KhN9JSJUaG1VxgmX
h/SpRe9+JHh9nOLEw0LvncDw25onmx1N32NdfM7XVPj8C1kzQ0TnR4MfZSVmozrp5YevcQkuhHzA
+RQT2tRR7hV1Ik0+2s0n/THX7TQAYc7s6nmJbUmbzi+uPA35kaPXnCa3e02yfrvnhoa70aMBOmva
r0c4DLGYakhzWkPx6q+rfF01d1/iU4gmvI/OkMWRD8GPKOkg9dJuON0m+TispGwq2+Nc1lsHBfSN
R6KDla0qJ5dSI2J+m80i02UpmI/xcFejzcuPYkK2rmsXYzcNlNx1E+2DzJ/HPxpCZNRvpiIpWfGQ
dDYwJYygeH8ajOvt9u2cQV3wlW+nCt+HC2QY+mai2PrxiFzrvZWquRt4rpjUj3+87C3a2sJP+xzZ
xy6H2axDB9JzOgygiYaeXtjBRmo+LsKb33FguD24N2cRygbxa20I+7jFMsoRHhPMNacETVFEF2Uh
qgCyzvAyjRD2DPphN9CBk9jyDU0MdJxeGvaBtON0kV9P8eSe8yh+39LQ9DnO07ueMUPS5Fy3EdFs
z9+EgfpNvIti1CBX7aws0SZp59xjYltJDULdbBMqUUPhZ/PjbBHPge2rMauyfq60ovmLtBR+1d5C
X88LZWhk/JRsrb7QBx0spBKBeU/gvE2BH2e+oPkyhw9xTIvd76s5xM1aD6HQZ6V8k0nmj9CmSjr/
HjtdcOC1pkU1aekAxxkKijb8g6SYrMUT1yMuvTDvqmFtZK8GeLC4c5zS13YXKTt0iGtaXFUz/+HN
m1uubCEq+qUyyAyv2L2ni9tKfCpXSpnZKVguh/F9pHebvdBVLSFOGgHAgUZ2/3uklKyiEDDxk0La
tGVRkpif+bIXWJTtLf7077uTF+X9W0t8OZsrsCSmV62q0280G0VYSwJjzNornYvyBpIek5CKNmVn
aT+6LsrgcnBO31LNajNriY3WZl9aoYsTP1j3tU769TU4S8Smfujr85xEY2CtyaFcudZIo9QkiiUp
9quro5Q5zPlp0KXG/agbZN6+zlGKYEU/nJ0pKeFkqP4zz18bv/xdJ9HugjuKpaFa4NiXOFNMhuPj
QOGrpOzbnHUhVcRoTjS5TNpv/E++Rf0e9O7PNt0gr/W0swC29noj2V0KLzA6vQyuheL0/BeUjwPK
vhQ/byVZcU67zdOp539hMbAIeguahjDV8GitWprOEN7TN8+jyTq/ffrxVJKm1wNM6GQNcfl+yUJv
YNdKd90DzVYBhbE0SLUrbsyH4yC6jFVx0ruHoAb1rkoLkULs8BUKqMAjcmCIrxwa6VKs3v8cOdNU
fcZyD2BysCNplU1xerJ/7bMYTi0FmQAtCR4OsW6/da7pneYsxEMmZ9vAonooYRkGwCWLWpKYsupE
3nwIU6/exywT5Jv8kMzNxLRBaCftZw8qW0tHIfBvsWIpIaLwGDNSuZsLCn7+tMBGYuxEzFYQQe6U
FVPWqRWvez7xCtXDio7yMdB47hTD2JJZPuzVEhbZTrgnbShCJ6pQDLBJI1i8HMxEZ68ru06DVSxw
k1Ic7GhsDDLffVX/cUav87aMO/sH32RfVrBRpX7HheKo3YV+LwM889S+RmWx9lrjOlLnLzqmLOxn
RSrJMI5T4oPTTbeZakFBZQPqCFfACE+AiUKMx9MKENUaAibW8bEvJ0G7z36R1uO0RKhsvyK4VLVy
b+OG0dfMc9QLXyVBnSWAalPT37gjbwoweYiDzus34HwOedHn3Mj+AUdzwtvEac+GeZAm7019kMY1
oq/dLZiTOzLeYoGsMCvtXSBy3og/KxqA9m7D1GJc/8y8y16Txmtfa0v07ABiZ8qYdRl9vMR1yoUz
qG2t12nT0pmvzWii6BxnmHM0FVAmE4aiSmQR2ieb2BpDWemAzSPLcpJn4WfjxJePmUi3qhyhECAI
KKiuCR8zV5X1BpaLid1bXEmd8sC1UwvSj7gw2jl7HpfPq+S/oNohz5hjEdnw9qsEAAuKxP1pDlgQ
C/Bah/koaQvng8UZ+6WfNezTiu56KwQT+1sl1hNYJTBV2erg2l7m8W1yHNf10LY21GJCHObKjzQb
ftIfd+fnU0kjr8z00vSvByvf6TIV9tChqHbgxITwS0eJfd4v4pWxhfciz0oLp4yVsajp2hZvG7Bl
ck//zlrQSDPhLZr72wpKajTMfU8P71t/RrF/9ZCr8m0jMouXMpAJN4aQNr0wOcBPbYA2ectuRq1R
B39N9vgtFanBeQnC8YDQXvOvpQCkDTm2EPfYEhJeAxO6FHVJKhZOAzBBDi2QzWcSmZcaTBwvgzjT
cAIxgPdDllZnh7gPK1twMWi0fCmzpnv9Q5YEmYJNjJC/OCJYcBpkYA0yTKztXooyRN9JGg1py/QF
jC6cLCPOKJrLNdTqmnb2ho45WmC7uSqf7Y0JVrM1Wwifjcj+YJ3wp+ZRlu8TLJ0827cvKJ6AeojS
7kS5PpSRDnSFD+zvkJJilhLEyRDty3iF4XEQMNQ8LNHmCOcK4CgGvd3Y6X/sDupj4RvjzsZyI1f2
TWkgvW2svVntjbt1p/88JoMrbbeWQ7ecZqHN/r5rz8E1owH5fNgphtvgSSDSXE2DKUZG9w/32zC5
vhxtYmHajQTszT5emOr7qEWJogVdriC5jYPFz8kXV7aKmD62GlLgm3J/pd+6c+Oe4alINr46Ai89
lR9B5xNG6yHyrrZKHJR/h+JsOWcr9DeYZN2tCxR2YSAYIVwMff7vDL3dsBSigvEatNMYtvHAoy+9
SofY6p7yCslOdpnuft24W+FppZon85pXjWszda6qE6V+X3ZauCl+1LZ1rlfWYyeIaz8F+C0daOG5
7PVGGCNSwyfzNg8S2WkHpuqHXM56PsLD979dhICGwPP01j8ePrpH8Zi7XxOwMolVqJhcMCmv/Icc
D+KxHBkxlKrtCfdHzinye12TvPJ23PAfU54ZTUUa1qH4kltLq/hmWdGmoXG5x9UEIVMBGmExJW+8
DhU/LjmU+nCz8dk2hRh9IaQQCSCAa98V69hzY11uuCe1FI61rn0L1ZWJQQPbRjZ496k7RsrlWe5k
EhXnUsvgUiFIlLD7Tpi48NvyFW2bbL/SExhov+spUGtLmg2+55VGcHXryPUNBhsF6fQqEMVffRkG
LXEdqQGUfVAxcZ7bsHWCZwAJJN9ttBMdUakPYw6n8+aZcSeGUOHEvdAvkT1mJqOKc604LpDf/xzL
pj8MQw/fWgmJ+LTL/zovQBzM7dlu2+jH6D9ymzor3Nf4a13XUPjN6GJVCJjlO49TbHLo0LssYOMB
33dO4kSLc1Lg7VDncB93vkLKNoIkzFPmIuflxzWg3H/TwvMwVr2SlSWmxmeZ0JaIQsl13yBUAVNE
jpACsZixe5HeXQSDORtbzNJkLLvbS0teOKT5fl2YGQhGUY6K7QpgXSHl3NyUUnOIFJ64mkgt1o5z
xglZWR3AGCWBva9ycdlFxGf+WqX6x4894K6e+S92irbelcRFxg2MsL1OwExS7wt+xwA1IqY6BZhW
xrg56EYTjxXjjSy09LxGg9rCvY69YVME2+JloLvFowWwjqtfzmjqK6nTFlhJORr2nLFtn1xt8G3A
Hv2JGfEI6QzP3vCimGQ8nBOAZ2rHRSVLpK16Nwcqz8brFedShqJP9NS/NOTUh9y4H4n3rwk0BtrU
ZmHRpmBeBBpB4nwv6msgppZrJbUzjwWdxFJD6/y5ZsHVpdzSiemf60Td1kloPVaV4TWvVykdhBmA
q4v0bzVyBsBCLbdVdwIbVn4kEiAYTZi7Jr4bQJ9OnLoQX/weHdp0ccaYd38M1xSyEJZId1SUuEV6
3+tUUxUx7scpBwMYrU1oh+JD+2hvx91VvkhA1R1himfg3aXU3PZBzSwOnzTtWHvDBHhJfIMV6eoT
++kzBx7gCLVC3za+Q7V9QVPKcH3bDwlOoHLzBYkyox6oz0YQuD52gzAXnb75KwYk/7jHjyohx5JT
PW1T9bvEKHCKHyawLMEd0v8Y4BbzpawnWWynOQj1hkJdksEPgiFe+MDxsZ7ookcZUUBuPIhZ+zwc
9fZ0blx0kxBibXoY8qEwSSe5oYsPldQnmIJTpZBkDl4tMTUxWGzBSU+pmyub0JsHEM76fOolfIuP
dhs/VEAkVgdKI1f8EFwM5R2osJHylUCT4h09JwQKYDt+fbrUzxa/W5uLsKadOhRQ+kdZAhdCALcy
pyzdiHU5YmTVMg81ZkzvKuIei58hJ3GcEtIwB1XqDF5KYfNnWAWuRRrA7Sb9GtISZlQFt2R06PFR
4X2HZt/goaFiietHHl9+Nen0vIuQeYRxLhFfGHeDJdvxoCNSUFn2YfERN57FRs7OAo512D0yKJT3
e9wYTP5ok9jgFHikQsN+o+Jx/ig/TuXBikDoDlgmhRO05leWV+hboemdE+kk37ZcEuGTd0z4kC0N
vEMPoK2uZ3BpbhYMxNOpPj43s9WCcs8+kSz7h7Q2E8CHw8Prx9Whw4izJNPObewoOvTbaD7RRs7a
/yWfJMyidwfU8Y7nFbMpElVQzIsGGwi3MfJSUuTD+dXhNC/8UBL+AW3prZdrTCflVskLcHzcLPiC
iq9VnZQKM6URyuzVWGwsHLSglLLTpjf4AwLxg/GfRVbniMlRjilcty+YTZ0sEgIKjSfDiokBo8aD
jMMrtsNNCNL4nFo+nqguExoRIvzZH/vK8SzFFNgcvW8Uc7C6+Zh7V7xyifUDexkSsAvHYLAOf968
X9dBNJIbtTTpAAXRrBFK6VcGYWhEFOprqI2KMeKe8G/oLs6m3+N7N+FK8SEzbIJIzcyCWher/KsH
LCbqEHC8zClmV6jCe37YZtWBVh/MowJH2nAdhwHvTeHVvYhuUMsX+WDbipSJM2KkHb5AY6Lpvkh/
Ci0f+UvIW4nr3E7dYbsIHkmq/2KQ6C+EEX8r+pcm6P1fiWKT8mi5xQ72CgoVwlhkU3zhjK7RyRo/
KJCldA+sTZtRs9zMUKbwFxEhi4/keRXdsJ73JAZO2GL4m+7Ep2AdTqsz2kajJ7xTnVkEC6ZoJK1O
B3RIvBhznPX88Tl6J0B0vf8Vi9Y16ER6CAGM1kEerO9lgX2tMlwAUaK+X88Q2LXgODuhfs8L6NzL
wOSeYC42IlAesFu8Z/z0cdvyQQP7y1DxQkDb4LYgpqMpRF+fD5Ai5HOJ1Sph/gM58zb9i+XxHNOR
ZZ5D7/6evKXio16cBTpzwIcEUyxKiSfL8nBTrQjfcAgOdylNf58ILenW9vdnEnUNz6Rsn9Mcd7GP
jDWem6oV/2lLLjheSVTluq1N/ZeZw6WNlmiKRtEa0xahsZbnlyoutpFbYCWN2eL6+s0/yAzNRJlj
Uvr3+1sMVpqehWVCW9D+zc/juI/s4cUhTUTJphJYq+lqMOMlS9ogILnmpwl9HkP3wVizJCULkVvA
30B2wXGmyxgWvb7XHkDyvyBp8Ho5kGknHgm1and8yYqzqO9Ff3WPJG1qFpyY0+s0PVC4UNoj/CNQ
cxjy/g89DiJyttrF7QKBKQJE3+X13OPoxJCH8xLGZvjKRBSwxdz9Eg6UDsbdhEf4GzOUI8+ObSlE
reT9QHENLqxTro43xmdD97Rmm5PywuaDktIatOUDUkcTBH51xWNVTkivyI0pjFilzVVlHF4PU8R1
uP53EH8LF3AFR/+soXfcqyASOhUTnFy+D3A2VRll5cztIEJCJcprn8QI+rmkwtCODCDWFggkzJys
OmYHtXMvnfXNcssZZDLkjtWPWya1E3UEYY0Qa4AKDZtQkTWYXWtabyV2vXqaxkb+AyuGGJY7DAUO
or2dNwg5XgC0kyvVP7Ump04JX8aQZwlbTzAH5Cyi2pIrIIvPVcSCFrBgNnFZ8VfnlCseHLhiKIiG
QMRw8nL0QJaZXE9+YTGMefkBSZ+/hTFSP6SsI5aXyDGFnKF7nPQSlEN2br7d2dTABWR7/uKucRzp
uRWDFSyDtC/kbVlimE3LrmHOfTKBWnvCBu1HK+dQ4FI2eFNtELdmxMJXVAKshG8ESRFfgqaFsdyW
9KiScoXH36OLmAxNquVQvABmLh8Kb/i2REeH7+zucmHopcxjwmrGbPvjAWdapWqh7nvzg3VPD1wI
bBXKYQJejyqrQiESiBAdkebS4vx+ybEV/RO4rH3bDU4G7oz+W91R68j6/FthB7NNJDjyxqhQHqDd
GRUYMHO84Jxto70sDGzAsmyqUt+jW1QtdYFFnUUNN1/RwMprXkNO8CRhNxZH6wqG4n7tQYQ1Y3vj
VFvWffotyc/5rHhCWBelT9cV5FDO3Pf/+sHGY+DwKh7j7Y14oIWIh7FmE/QY1YoIwv2ivwTTkJMM
iFsk3QNSvHhYYiwSYVmB/Y3tvNLS0VzSKZf2VVot0OcJcys/DqiTRWHtaJvHp64DMT+FtTZpfYFm
Eexnl5MyWC35y8zaJDlyLZo7VcaPFzQmJNFxGvqN9wBl1DYNMT1LuLC+euoiD6qyfazbOX06uats
5EAlk5w7YYHigvyRByeegkzZUQFcbGxmch6Kfop/pNF0vzMxnnBYN6muVhaqZTd4e1GUG8d8lqHQ
pkaMrbMISiu+1IoIOoy1oKyBVkmO1WperaoKeJK6qNlIR/xn6Yg0K626TMWiaXaJZ4e7PDhTcx9M
N7VTx8qeWPFqjGce4GyVDTA50bwLgXgKrsL6m6nKxbMghgfzSIebmEdFGbs2kdcRJqGuiQFzLl3x
9ETyp+c0B20l3HMOPPbHfTX4XwATje+l4hM8wlT7LplMxUi83b7ZbRDYHU1sY2+iv5Qd3YZoy+Fu
m/Azz1Y/R6DlIyVbV6YW0+MXBqFBsTbDtfQWtD8V0JdrQqNVj0VBJzAkAUrW899YL34DX3Ry9R+A
bNHWOvF2Fo15NiKjYzx6tekjawc6Zh4pOphpELgk6IumbxGDBaZFvuVHjdSAZ+mM5sHc3TL8FE+G
5U3bpSAR3gS736DBfVCDK1u2eQwIcU2MXlIFBD9rFvj2y1xgD+EzGyfuvuI7fGKXyLWe+Z5/UvMA
mtBdcZPCRbLsuXAW9pVG8cOLp/YpIUUmVoXoA1/hWH9A6B482QR+n7ERIY7D3cJ8rWpUzgW5+YqV
sHxcyiDfadQIUlugY76JeY9t71kegnzfhOZMerpLxyvLVneNpGU9iNLEzhrTkpiv2+OGWVvugziz
POYHXIAtcBWn8DhZQEpYe8zpZWuxg290kU/zW8wUI2B9bBqrHg4q/X+Sh3gl8qXPY6do8cVGwlKj
dGBhaKyGUib4FNG72fwGL0q1+s+g8myslhP98cuROPwBHjQvBUC8/MD4gHeS3f+CvF0uNzIpOnxE
+GsrIen14+1fcn2B3JmmuekQ0xq3yXrxlViWUDvn/YRkS9yD2WV+TUpfnqGa1Oyg2sgAob2T7Yv8
kpA+D2eNCbelLNbgaoUObrXTlL6l3hE95saD69XrgCk96js6uMsxmskKWZWjxSj9y/yVJiMytqd4
KP5LXJlJUn7G7qNI2b25e3vHQnTH+vO7QD8A0w4eMiBYCg6NqU8rKihnOadw/mshIxWVjss99+NM
grYge5EShFifKYTCrcYvfaFL8xyStWcMmrmhNdLJQC8oNuRZGu4mwvdUAoIbp8UUJsmuV/pkI2s/
EPDYpPPlDD+UknAjnMXJoXGz3Lpx8giAKPo1VGL5l6pC0jiJiSGjtiU8xeRbyS2GS95Dju7XxGwR
2M/t4qdyLty1jkRFiEZdxEU1auq/MnXYhPZ76X5hqfargs/tWbxPu7jAdU0XAQ+tF+UelFauiKQW
wnki6ZGZcNaqCNf4qBGcWxleRppJdBQbMqPXIuM3zLSqPPVbUOIT7lb2wChsVuCWqmbcbANwbgsT
l4jP4avalisSLa1rgP3IoSg+z4rRMXOV9YcmH2KOVZbPI+KAJprIgRmi6/eEjwQWWAq9COyWLcCV
KnjaEgyJ+y3u/mtoajWc/p8534kplpLwvncu/JccHMzpAEviqQUFz84siu4K9qpxRgSZhw0FT6uY
/59T4zEKMRINuzB8KCSmD4m+QKh/HazkgonQGHttEhLEdDSmzA0MqMs0qO7juJ/gG3/dNQ7nJGih
dXpbvh7keVutN7yaTusKPo7egDSXb1tc4jH1k1HP0yIsJ6r/+kHtkh3p/ClH/ggrKzJMa8vtBprh
kjHVEbMlML3pqo+q3wIbgT5/mZkA/mHIJYBhIChTrArZkB58nmW9VTb+fzz5plw2QaRQDIrEGFTM
CJzdd7BQ8QFeJpzWAsyUI6dVMDYZt2JlHrUy92rBONOhPdbuZNAbIusGJnIbavCryYqVkksn281B
N2JBU/u+mKbDutmfiaAQ5xw9Scm5H2F97NDnFECvwmI4EEmcZxB5LoLFGDCxkyhGVC55J7EC0ZfJ
LuT1vfMOYcOmkoMbCQYplsvOF7vPQQjBrd/NdYxg5PNJ5DXJSRn7r+aieXFFhGGM0IutFDq75HoP
Z9ghunNpVJLbi1QBwsT0AmCy6xn/322uf38HuvMI1E2KTUijHTKlfiHVl9ka8juNpF/9eQLlc7sA
GqtAsvc1v3Q2/M0CSowVmLce6GjNElZbRqQq63uGZp8fXuMZM2hcg0NfWYcHJzP7aA+hqBL1orFm
vFjzYCXQYbiwluCSZl+qNS9M8R2aULCdqBAEUCtnqwfCs8FtrM7iyYkzg+Fk4idrorknVlJJirRE
efr+3IARbWpMbxBYzithgACVL9qe4BQP5DilkDFsvPcazFAL9urYFxwPTQkxoLFVuSfKYvyZFL1f
TC5UOof3CezElYeAwNK/TtpbWexJ01ZxxbwrEpau/9TuW3FhJQ53dw/dWQ6eVAb+WLYi+zoFiIRR
0nZkI7Bs1tRr2cBKqjx8S3RQ7YT1uVva8g5fnMZENsFBPBPiaxjFFREKiSylOFgAf2Tdy5w8TZVY
f6uzOHnbWTTWIO8oDa6kInqKxgf5fyzJz4ke5ZtdFLo+lNZvmCahzehTgXA9tsNXU5zyvG6c5otH
o7dHMXOVfSsxixHsh++2fqT3K7wTPCfptMo/gU6+I2CUzPqLWnNn+taiGxvXNsETVFvRy+L1l+Dp
5C/dBTeJ3aDzgwNxAT6y8dx3mKrqJJBv/k9Jp/7z/8Rn8Q7xtNf6EYM95u7UtM2wgUBnV1m1AQcD
1uVeu1TdS54Lf9IbjBEtI4ZU99owCziaGZnv/BsYwq9kYbMJUiyW+qltnSlR05gX+iOORW2iq+6/
uAzfnNGhCwktgAXz89Dzp0JqcbA1BCydfDUhVdB5je8BbRbQ4ISVH48sH9bq4Pni1uthBdayQYG4
Rf22Gt+oNVKFojdK5XDgtyJPQBSVqqgpiH/3Ivi7sn8p/Z3SNwcYi7egoDrpXQWE64dGr4s7oB4z
ads3DD59wECvDM264sUC8cTWeIdujNnx9c0S69YIZAmb1TbXbOjFMiKTyMwgpOxHXxIfD7U7yxeB
aH/dOdUIQFq6DWsbtFLhTCET5Sb9Y9qtyeecAJ5318490kD11UoRfqPM2TF7zU78xUiSA2rLG5VZ
TbVtLJT3g8SMu8abOoQ+wIhBnT8qL7F2x0y3Mn8vnPrXADkOB9p0phG70BCd1N1hjjt1E0oz51JA
DlwWCOOvS1UGwnwrh0YXnmA4qcH/YQZS/C+YcU+K9jn9RAFpgH+s8zTkzjtZYzUPZf9LomrGixFh
hrR+54ImciqZFCw9rR3w4Med7Y9Rfea+MYOPfZ8G4r6QAEfujqAYJ5VzpplDoXc49Lo8/Y9+Ap81
JX5twFei5mmpUxOGVWjL4ipeT9d/OGtQa9jfrr6I8cIl5tcm439dDcWESmLAmqneOYG1tFrKxX/b
pL+MVEi0qblkCKiGMy/Z4J9kKkUnVkSK7Q/gyVrabgbqczq3AmT0SvQbpkR76dZFZxufabrk5q8t
uKOUibJqWc6qMQ+SnSHrsYW6H4lAOUuzztZLd09QXeVUJWNxofomQInD5CUM5WfD8jWPhfIjzWWY
uC38qU0Ml5jwm+yY+6cpkiP9+nu/MtwmI4wYEgR5wvisj8MQJXqouibz4251fouY4pT6dBnLTwU6
bzSQALYBkQyPsd/94hLBmcGUMRQ3AzPWmSW8lPP6vNsuFAuImJ7OAbcWCXTgkSlHgS8JT5Ncq8IT
F5oxB7aK8bO9rRNFfe6ThJsNoqgor3SIhYpJffDxsFrnQq9cOT1dRirxF76ean1jBhv9HxCU9g1/
9Aslc8G+4D+cMer53tEKaGvUALjdXCyRPag/PLLDTs6cuoTgCFwdCcBvJKqbjK0vHLooEERaqzDI
oCMGMWsQVDsCuKsHhPeCgZPTdnLtyyW9kfKQpD8Ox8UdfnGkQw27ULCWf4zzSAh4r/+F9vj89ONp
P60u5A824XNIEMUQAEcoTrtIQN+wb4xXaTeGbjVBYNHJC7bn4zjuIcvajJuHQ3TXpqhNGcACecUh
0Wq5+xwZ4cKs8UCoUxzCgDdBDiBNAEomFOwcmb4bsXazTYduWtoq2TIKOO2eTYidIgkBACkNA3Fd
G7bTolVRmHeu8G4RIt0ow+/iDKlL7Hf0Nj4pknc4ZW5T1bEvQ5xE3d6oMWHqNUmGWLqTcbqObWP2
hG9d5GsnZ3mVk3slcS6MpZCjtgUCWAfZc/+FYtlxC9nmcekNTZTNoiQ3OBfBb1FBWO0KxHUKYr2g
YvUXPlr+5kg4gjQeRzuP+rPVnYExYGLvhxhh4Md8uBdoh6yoi6meQkjUcPC0sAhrRVnL8hsq8yG9
qvlxjIacNWacc87lQT/ao6CrQGLb6RqJKPbH+BkiONYpcJ+KOHOBoELtAu9kNAk2WJmLgW06U+mj
eS3H0RjaiXtmwNoGb651ghTAMGU3th/hfUv3FvAkiIQfUTR77XHqlXlR7ArmOjAXOwCUZPNIb41w
OfKULn7JS9O4ggAUTxgONkCIMd+oTnEdd22OYrH6PFstj1OWrDZP5W6twKsHEKkUyA4CFsClqLBD
ImtmgQr++sP1dXaPGRRVHJsB/7m+FWZL8M7mYeot+lDZHzwpWgjN/RJtrQI0zgXUYveahlCGfvBJ
En6xLzR486aOhL2FqlXZouwbV9h5aBMgbBPQfQ/cTGytOrmnaWF0+fPGEoQ2qC/lAktxXPa8aPDH
V83IAbCdr3cGQxCYK+a2QZvo6UWWnBwfOpchNsxcHoSeKG7uUjnXbDmMY4K81HFVLNdeedgDaDOD
It/T22DB1l40GVjlJ47KKgrYHPeUe8HYwRVgKt6jUOy9IHuPjkj5Qk9/Jc41RQoW/ggBFNX4wGK6
6qr5Anf0YUESwEu5OExMQBO7Va2I9iMrNhsmNQaJRZQwFy56SRWhngHyXVszUYiXzbEkn3y1Y7aP
1pPqnbnp9MF1eXDcDrJcpxvlhKW6vJmma+KzyGoF9iAWdVx8Har8vxnJ/RHikcV+Onogfh/pMMj7
YLNJtKX0TPLNjXBqNeO6EQIjLGZkm4hScoTcYWYs51CvwPPxLYTPmOSBuD+VBT6j6BtyhaifeUzz
M3tpdl65pGThuHBfI33VT7COysaSLZU7hsRw2KE1JeNJDw+Xw4Zug5KDoOopvSji/ZZ8dVzbcVJM
cyQz8Y2KJiFVrc7Pt6EeFurP8ICX5NnHfn/xNgvQpENgeBOmOfxbgrk0WaCLQwkdAqCV/g49axxq
OIgLeZhUatD8liieMWkOFkezwro294rDfcFYRMKoh0H5POEFYeMbecUx2ss+D+BwaeFCq30nE2IV
bvUMYOcMTM8RunRvUCjG0uopsnC7EA2OLUReJ+hTphn/W96PiAFo2Zuj4cJWDd+NZYJ64eaT81Jn
EFTvZ8zms/wJ+UA1RTat2/LUhzjNMaiNSABRo2vJNpOf0ufBxR5XP4Fa8KyToGzyTcy5l8FYEv0w
jHwqUvlmwAupgJyYzXcMMW9ZVlmyJ1lL3EMW8XFcejQGBAoryz3klm7i+fVlJBs6ce/YQaPEXK2l
dRwyv1VIUpXWQea2Lkyizwi0JUeOu7Ew/Nsh4jt5nuGOOzjZfKu0d3kKdYPmdP/4wqFT8+w8Os7G
XPCSmvd6MufxHuv/oXAFxkQEp4FoURnFQFORi5XjwJvOYT2l4HLdlCSyGwN5l9jmVYNNnPBJrztI
Qyg1CoaRThRrsB5MhOtd6mZRVVoxAorZ+ysAVHBv7VWCzQcbabf5KXDGOmYb7AmwyRGKMBB4Ew7v
FXVNC5qK/5oGLmYF4F/ZjX0rWDUq7qgPevvEU2XDdvKldY83RxrT34uwRzWW2vIXmk+n72tX4QDb
EpLEGX1wx6Ege3pIxWK2YyeaNn9bHJM5ylAGSXtd9Cju7iwOcBxFtepspgbNGHhRsHUjPlD+QYu/
45MFxPUkzC2uHQlJ68J07AQj9DGUaxuV87yqjhUFWfQGKK2TFbbb2waseKV4JyTtY3iDy/EreN8N
Nm9IR8SCUM14lZdWBOMregaQ0AWy1FfCc7oTLvgs7ec+ljlydHDJc+scuvzx8Z4D3d2NBMyJrald
YeZMIqcROYU7TW0QSepfOke2O/4vMZF7/HTBZ0+BGhrwCeBQGLPTq7aNCckcgeazndHMT8U8uZT2
/M0a9JWbHk+5lvSXYV4nIPEcuvlrg9RHgReTy6tAvP92i9Zwph8xdqeu6MBvxgT/cOK1PNss3pdu
ZeDTjnmJH+OAnNGrhDm6FDGsNGJtdDnbHGtiHMJFhWUNSwTHZoGsKhyuRtuM3u6DMBmboYa97IxY
hz6zxlMPfQfc43+TXdF/LBAUUDB8mdA9h0AmwzR8OgB97mH5DX3HsKPJXBceVfKXZdZMtPbMU55K
lJfvDmG4mH05zsbY194LfqYDdpWr/8fBQ5Mr2qHVJoQRyD8x7YdAvN+RWXMGDLdUDLhO82OlVIK+
ISxsQGKXiUFVc76VraIdvBKzvkWzYYcY0Bz5DzMId6GHNNNePeyrzWbCv5YyeLB5lsaPxxHf1o+n
CA7tXmdx66hPSNeyF5OV3WMRicmf7WJ4tkete9DUEVuSW7CbISOAjpwsSULn2pwee+uu5sxQ4kEI
uhF4TFonpoVC824pKfekTN9ZJQjO9ZO75RndGakqe/quINrcJbg7SXAMVZqj1wYJPvy7CsaV+I0H
2tkIY1cLj3+Ax3DqSiGcjkAFvivZ4L1R244wTPnJoWjq3pMi1TI5TRzL44WVbV0f/JeKwaIIlT0U
0ahuB89TQymBjNhdy1oTa6aJDmoJxkcl3kxW8h1kWZ4naQFs2uIclCxcRAnWg03fv4agi/2MOCcK
E1y4ur8ZnTa/ehTNUqD7ABPrh3TlidFdtszp2gj7OrPRex77WqefqI8+XwCmKKQHwQCLtWXNt/EK
xA+9byqEohXaYgtXJY+LEHk/jOwDmhmqv5yGykqLGn9+dXOBRh0RoCu4eOmwGhU2pB20MoJX763M
fCwx5Bj+KD3p0bWYS0LOcpM2DfOXj5lXghSP5I65OukHVkR4OIc60opapRS6G4onYX608h7nPyB1
Itxldn/1+hmVR8BFTEg7OnXn1vWNiuc/7xa6ErZyHU395HewoAa8LQlXxgWJIeJ+dGLz+8fi6clJ
lV0oTEHqdaqhIQNyIgdoFtgFNkuZLMUBUBQSUD/Rr4Wh2H9/uVc37TpdflijtBNfsjOS9LpWwv+C
reWsDoKzFinOq0zPm7XwoT32B0zR2ZZ4IchHe8OwWpbWLCe9tXIuBqQxgvCBgaNQ8p9Xp2Zxk7IE
JX39G5z5nxa8JZDpO3nljQVKR/e6EDzzdCl1AfyRMsYJ9UphUE0aUn9yE7BFIGxfvz3iXedLZMjv
R4fM6y0DOzP4EDhSSjmJ7oHuIIQslu3yWqHACyPooVqyM/XMZhrkfFWlX/VgOfGUuXCn1OAVIH8n
siqA+eXwXWYDsWS00r9ZFP2Sg0z/USis3VOi8lrRtlt60pVjoDA8fq22CZY4MZ+Z6k1KEvaGLTb3
BSDgog5R9TWoNd5CEQ9f5FKeUBH7TANfVQh8/3sx3716c89du84uU/+/am0IyNxuAFq5BSIQEw13
F/aoOguXfAdUj6X+QkprSsWb2C1wc1F933sqwrVIshVN8PYBu+xtZDBAmUlSg6xuesN4J7XCYwRy
ywPe2V2/L18oHynZVWagJ3gFVgJnZHsYFWuhyXfmcgu8i23v+Rv+zpbl+1lZN3yzLdXh+7SAaSRt
SOYBpnLDaZZB2LB7CznGH2J/+q/1j23YLnXh4j2pSqRPAC/97kjJnib/EooMMGezq3d10BTCX1xN
5huzPWRFaI3tCmpr4IFd9eykkGMYVaCdAydVQjYU8h/FB7Rou5OWwuFh5pSHkzv2+FOgFA2kIUJB
j7/yn3ZVv1xZ0T17k35TSDOHDn2E1WPCBZvLLh8SPDOSugLZF9Xnf4I8X52cO+WuTXiGxy8SoeLz
9568GABC9k/6ziDr6/eXWLrjUhZpNgXmjAvJzbY+z0Qyglw3pW+g4S+0N6t1UIpt20fta66FuI1K
q9nhgHJrsvBtzfEwklvZSk9BtARE2Ll/0+gobZRnnKdS1WG8sC2f/aheny2gazYzHcxpNHC7+Asm
6e+o+oT6vm2awmcywiDtJuqnPywbTyr04ab9ywzSpz6ud2dl2M4vzVaimD578nIgQ6aECgIG2Rli
zROHAQwQH9sSBI89goQA2ujP88HQKVtBYMAP8yExnxliQd8nidKNcNKSA+qPNrNYq8jsmqCwAVn7
r69pqsZLt90ZpkF/dRh6Yn55va3afP1GAMBAaQNlP+UzZ1YPkAaT1F30G4etNdRlGs7SvcoGkuXf
FZc1+6bE6BrQPWpdfkFcdSoULhpvEVlCPD/z8UXt41vRpdcO5Kg7bi+PhR2l9Sc3ri78pExm5bA6
2yAi45mfZvuvfcypwtvYhBmpQMXoWNaARPmr08tL6Y234WFPCtV3sTgwr8E+nfDEBIaHZ7aMzdr9
Qx1v3ZHqPAnlwy4L0gvgbbHrU1Q9DabwtUvVWWc49EToUx2cUs07mO5mXKIWdFcfyGH34C1GDz6x
PApIcC7zqXRI/WVzieSs5XDKgslZuxhZjQ+360cO4SKPdaG6rTnkcX9xrgZ6R5VigTktM/upLb18
zu+UQ1S5ceV5J8OGS7zUi8NPVvHnbWfBufB3YtUfrtrzb3wPD/TkWo7bq2WxViMF71A8cG9Zge+j
KucsCdmT3z+bs3bqo+NGGZeB3EfHPM/4SPKWfKI4Dp20RUAPHqllf7oTRs9Hn906TJ3h3+E5+bA/
A2E4luEoKSkvrRQItEuzPeA0BuRilwe3XnqVt2f9tZzm5F9AT+N3eSjOBNsQNv3/pHNdhO0P7lBv
ZcuRieV12mv2RddZIHtgPEJTN2SX6ZxKh8Spa2JbFU5FfXDmzsW9acG/UP3XjnzIUbary+MRyAZt
ZYyuGscLKlojTXQSVyp2Ypfq9eRZkrbBSMOha1X6uWIh8nYf56N9AMRTPPW/VfXvCV3dCicF2A5e
SdwcMQURBEeTC2oqcj4VucYZeG1BXT+7lALgHm8LKNTrKIYdqk3mx/hVMhpCU3/0h6at0dd3v9gn
cYfzPDybygJ2GRbiSrtxzya3ruzdzOJu2sUOXlSIvo+wgABt4ld80RGNTFjj3FK37QJaSix3Tpe2
zbr07ufpAi2WuGwO/7qbvV5asXoZ2anvJ8OdyfXYI05G9cdfNdRJnoHHvEBMAFznttQ4BXLrci32
Jey9e5MQ9MFUp8iW9eyxq/3VT+RbhElWzZm5uuN+EXQzWFaxprmdiPMlTVeNl8ylSA9Rl960Ll/L
GNZyKMkZFkuSSBdp4NX/9X0CkJhDvzRRx9R1/Uwle7Dxrk/Db1QNnZyvmzc90zfZllKlJRGNCSvP
gCCLcy60e8M7lJ4Lv72OXsuSnsiHPf6JZTVGQg02RklBNll+WZlhWO4MukO2Jzfg+DMx5chE2h2i
yAH6/H6uISJIw0GiOFKh8RIvi+HIm+KAejMpuxIlarOHuWbBB3Orn9ENs1gRssHrH4lHq1tZFXV2
PAwLujQXdLhrJBD4Iv2Bpk5U/FsQMJfbCDISujd012pHNORpZPXOQWCeFiyLNP9rFcmSPoS63jt/
NkNSw6Ns7BZc4vFjv0pp2G29hGjhV2shzXzI2K0uO64/AkHiHToBtfu/D3n32Zy5AofbaynPp1Ew
N6Phzxr4UmeM60nrnFhk7CjkqiDjMZWa/HavGs4/tqkK8AYgldZUA1yB7786Vt7EZfyaWZ+b0uKu
jIGOEdwES6Bbhj5QdmVTZgtatyu0HjZcxY6yKvkEag/cCZe0d5tvJQkI+LRc4/j1N+UVonVM3MaC
g7AVrcTIYkKDh92MMS0AJ4x4VAt4JNSNes0doHfUhFPn4bVbcAH788BUB8AZJ8JPdDjiRoOc8O9l
GJtQCMV+qpHAWXQosUbArRVgy8FNoX7kCzkVhuAAguWrwa+yhECiX/y58Y0NflO04br79AmiSnA0
yAo++A4wLtTPHM2JhW48gY0MqCoytRAKamOGdTwPEZv8a0Jkk7L0Ve+RjDXFTb2m7aDfnsllL1o8
xrmVBFCD/Yu0bX9gc76zsQOTQEIJ0/6am0Gc2tDN6JM3+x5MmWMv0EuteVIdYsgZgSHHvWtP4+k7
SB2YIrX2+PpABX2JpbambzMUmq6yKc4cI1Zc0S+stVn5ddZWm70PVw0tPnqLU3q7fogU11sz+LNC
ON0+WgUO7GyWjsZNrSwUXRQEMgRRdWt3MZ4UO25Vvoyal5rCGHQ+FNdhWqT/MUte6yHxAO4mjugC
Q6ioS//s5fWSPf8MO3ymPqWwfqrEMqwxJNY6bQON831RYyMUkDhqqu62kFIfuWhWozcbfxOwsMZG
rgCQyMnw8Ilfs6uF0sqvH4J02Qcgqj9qH7NggwkQ3HbndppFh5PXczL/ZKD3jli2gFNN1jeVUv24
QvUGbYeRmmUsLwKvjsoqNV+k7wnn4kbIMiRxWYhEHxHf5uVebGHwEU1tRqqGwE428vSXfkhqi77z
scjsMhvuKhxZnm6yVFzsidOl/0wor6aDvHXHHLZEQIqYS1BdRHgDYc7DmBCTjZ9dTWKxnMXLmKjD
389AIhsHb0rZCkoiWRWy+PBb+x2DPjtmu7+0ltYla5pQVTfGDEPu6fKyPS2XPs6pSRCKTrMPg+W4
DOO3T9lSNmXcDMhJZ3bTQeesaDLG9DApkIm9yZX0s/EbEEUTGivj2DDbeuS+Jf2mxZcBh6J4CcOO
rODmvwpPzLKvH1C7b9Yqs5OvWS4wjMClU8Qd5Jb0H482l8hyTLnR5UWbWedXTBxqCUETQCHS3tdI
XZmvzPLU5ymeHFQ7MRaT58H6wqifqI8iGQ1jj20asBfkSGZzofYo/awZFzEkCXtbLRrSW++AGfe4
RTqCiHVkpK6F6IhNjEXImItvJTHV+H16zspSQLew17CKJjs0uU80aKwumqqQp3YtVUJMWlfClahX
BXQIuXyGHkGM5fCpC5bTcMH6FjjeIlXUFiCW9H+xjwgSGcKEVr7YPNT5qe1EZdria4Ha3tk0A92G
a44UJt9VdF3kvCZYSibTB9XkfmzAEun/7UgfZ5P66Z2uIqPj/2n2+h0ZOIsM7qCAqUfnuEk7cIXy
Oyk9sYwN7XMdr2gPrZ0WNLy29/bNLhC7pjM+rGrxKUbCAJLl8vypc94aPl4PdRkauk+pgIzBvYQh
UWhxlCQJonl0Yy9LN6PnA1qIjFQ6UwNr6xh4kAoquGxhFuJqPUi5Si0zmkZV+sEiJc3zfzKtWdx6
1rgA703AG5Aoe5HdNOAZJFgw8fwGn8kr9To1EqdvsVLW0EL1v4cPGC0RWMsAx01XD3u0kaw3N/MV
F4WxTc6ibZbGNH1hBDboYrRUxh4J2gH9hwSZ1sfcU71cNMmk53zwPplApog4z11SvXKH/fCefAzM
Z6IffEA4l4osaNwk+MNR0h8gCvtmmBEBdcEcB3TuqiFrJUom58hlHEBvDp6JSZp23Dp5eQechpv+
0XdZ2vPZxF++q3jLs8C5rzoLkJgiWb3Erhh/Di73x+86XuFU+wxf2fJfGdZ3LkEgUBt0JQ4iusiV
kxJCQjZ4pP++7JTs2iUM+hLvwvVZ6yrNOwuhlSvx7pZjGYCGxmrdSfC6/DPBXHYyVn2J3Scs74+T
9gzq1b6uMasyCf9XAysS/CczBiKm27uuQasXsUKuL3iqaiRNy0CZbQ24avfmmxtrVSF7Qq3V3CRw
DLQ8pRdpp9hJyPugMTKIgOAMJAIZgNKPjJv677SMk6fIdh5L1ZX5X+Ogw9tL/v00OncHqFisV9x7
3pf/ITsRTpa7XLWyGQV7Mdqqgih50O6fuZcLa5+i63IKZnZ44AS7KGmX0JiOConR3V/Ecw/QLeem
2sbDZ6twr8vbEaOvCGxhsnByIost3mVJGX83JnpE9bPdNAtFtKvMih7jEB0APHIBdzxcNmfWhrLV
lNF1xs32QzqhpfUIRLb4DpZG7xl/KxOK8wEYD9OGfiTVDw4sGHqRQiVysLAeBTtx6AR2t7G6S00b
E3rXnqgskIhfEzdgPtKrlpc2VBB1yQOFBxgK95YJDbPS9EAL4CbV8kAehyalnMGY2wolJlSv9t2x
CmurNfxhq0yMlD74N5O3yZ/FXH4kuzSiTy5c60Fxfgr5ql5SAJimyh/VDyUtMyDq9DAWCkoLpDpi
z8Oj4m0chB3x+qsux6mmF1nQfDkGbF6+LkBwExAT/qCpqr90NHjjQPhUqBvlio/v5nyxPllSRd1K
yBLEU/IV1oOX3+t++5oCQJMq9em/ZskwyIkgKqAF3lH4qnuZmtvwAVIu3BT4elHo41H7oUW+R9XY
GdJEj7+OYJzyI9TQhyBlCykeiKErUEAzHpA8VXwBpCRiRtangGFDX5FRUoKchPsOTIdCMNYjsC9e
KXujtfa/i//2AqEyS+ymM6uoSbE57LZXykgJ12xx8NmvBO1vyf9eZwihksT/cMOR8b/2SOHk2SPk
jGqKdpz0lq4z41klG/UYd9RTOXfgBwlq0ZCAARdTFVyjnmw40DYkEuSEP4ls9+hU/YlGfGt3cmkN
uyWAGjbiXYptbosCqaT3yn+87yknGs/XCmoC8Q6jZG4c77vSvXJWvovnwIX2UYYG6h92bcU85wLS
PZkv1pOQ6xaQsGedACPVtu6EbBmkqqD/++KEc5DweIVe2eHfaT6CfP972GC34mhf+fZtCFTEjaQ4
ECmSO9nBaO5bZHYpXjmmnc5fSwVXUblci9uBRUJ7RvdxXwZJsdewmWc1HHNXrh2ABmaja7BwUW33
jwJ+qi50s7rILl4tKK37NXNibZL6DPIDCDrFCUGE/5PeMCN5LmfXAGAhf5KFodfF+9ZlrK4Uk912
QxDSYK3lxHw620uThMsSISTHtUtZvpbuiSe+U6cqvhcemkjCH4+8eZKFF9SHLVdJjHuvkQgWFTgs
8UOfnWXOH2hAwaWv6OELG5Oe+Stg0RsQMpHJRWDmZCkz2/WUZM6D394QCzwS+6j7khfZKGWT0Et3
FmUh1l8I6/GeBC6yNofJz1j7DBORhRS0FfMxoTo3akrhebKc9aCzqTCxcEOCf9yB3dvBiXBxPx2V
MyviCteIAMQZnKU/mL/di05Gkcu0k2izTT+kPNXlcVwi5+OEFJQDka9NrL6bEkY9LdJczShK5jNf
0W54ianHCeFJ59RowxhPyfBOxdkxPxxYreFNL4m6gCeA/F9PlG3h6yVO4s8bCmZM+6iHjVoVTekn
lrPO0S8txiytlhj8GZAV9ILlxbVoe10OPPqrC0ynks1nr+Vm1K2CFAcgArS89Sp/IAW/Ibw4sM9J
aJlaFJ3YTRX7QJUbwADrRqcmhNNEFh6d1MOmRW9F4p1xxWQT6GFGXLELNc309S+WV3OK5RJdQVCh
WsFga3BvvUwRS3blE40Czx1MwS+318HjtRPhauNuJbUVhVfUUzvePX9DK5hphw8rd9ktdu5t8NLM
HU7rgGX6nSvZ/2bAzDfoY5HAuUzhNn9ZEzGQPWgsxprhMtAFcwykWgPB3TWL97hhzDX3zXXjOsgM
dTiUAwpshlL4uUC2xBsQt3gXg5dbRxrb3+EC5QBtDnveXG3JRNyQ/qCQEPRKewd6j4lH/y2lTF4k
t+Z3mQ+8+CNcAmujHexkHjoxeaG3ZW5ZWW/KDOTbgLVIc/J+W+NM1/Q/61A50x0AOGUsYqjm0eI6
DR3Wx2/eJk4Qv5YxscwVWm5DvwltFz/TX0GIh/H6tagZfCi7ipMWnqLBGtz5ZjcQNTKl42aUkQEG
SYCC54dec9mnjaWcS9E2BwGPBxTVeBIp9y/fuwQu3uMwffLLP3xhXHccIJo5A5f4Elns2IXmxwUT
dqeAG38T2vzKcvJXXi5UrQC/quTWcvY4XZdT9iKqOmcaVyR0q9js9vt2fcCNPdsZ1MNuc4HTU4JK
TWt8ef8rUGZqqmNji3YV0HD4LgkN5RcEjdV53drPXFxdLC/jEx6KW1L+zw0L1qG/RX20gStX25a4
xIRfjz9gHEd+myxtKJtfEA3wgjelNiMKrGlWgqigejar3vjdrHRTD+LoSWzlSnWlTiq1Lrvi8y/z
L0BPJvjBkRvZIpY42/ii8fxRA1j/oZUAVn5DOneG8lkMCYWDZbhcmMaoQK8K1GQ4bVFHqtq1+EvL
m1rcwWTVEuEKR2aRHlPmAHeqAm8jfCtYrXhJvsgYe85iTTE58XVuAdgadWHhTAcPYuh3oydcbTGq
WRn/05E4fhLuPp3Iu1SPfP357DafEqqmar62VZZU0iV8rcpxyOWcDJbKhvhQZMB5kKUP6obSyPBU
BYocRrqGDl5pZEGksYJTCaISopaHKs5N0c6EDY0Ta7I+y5797ozJcDnbghDx95nLKIEAC4iDR5L4
u+WW3tZE3AOIGgQO641tHIDIpvydKs1P8xTVyhlql+BaRJQhB8oDFlJs5u2UPJ2yr9+aiidhaC04
AMyHo/1HeX/OYFWWoiLMnDqG/eeLTkvk5SMH8tic/twnLstH5NHt8xm0yH99p3fQJak94wbc3DA3
1oSMVq5TMkgUfockLFg+YnUuSlPlT5X1QhRE3e82ZSHz1bF88qu7a/w5rQqL7VGp15ta/TAQAgtS
FPg31GBRXG5uWTC8yDopB8LJvq1vO+jrUTbTuLkNrehib/H5qRIGrltNJLQGsDGuTDMON/0at5ut
PS5lHGvYyXp2wR38j2mYDWSIW4ba44Bcx9Jp2WjYcd/mlH7fZah96kvqRZtY0x9NI7tqkTu2FUxE
W3tZvgJZjbJayA+Al83ANWP3hUlQ+P7fmKML/IMPHElYyjUaPS9jQ/qquu2jo8s7mHHBh3TNhWGf
cJEV9gmpDgPZAqQ+E5oGKjidmtGzVdAed5K66cQG2njUd9IABG+APMHaj1G+17IcQ8dA/4OCDxq1
yTyeSpJOtzsw9iNsocV0jBj7VbqjBB0XAFK7Aq6Y16ppq2nigj5F6tH/nU0LLoFQtEtX/A18M8Vz
WQO7+TJkIOX5o9a2Bb8RpO/qcdxHEpUX2cO3n4Y59K/SvcJejRndfUBq9ku4BvbpwGqYRtxFXYzP
mnDLl7q3GbjFsU2C/+haPzZBOlpjxs0fcEuV+U0wdpFiewqe4rR8g+jv8UuksB8P9l4IUCN3yKG4
6QZ7gTdYeCVpJLLMNhUzTOTA1Lwe2xqt30jUFXXdchkUwuS8IiOASmTVCYzi/sxN+F5EEXnNbBGc
ajTbugRoioYS7SealOS+26TuYU2ytF7FoMFMBamA9qlH80pqgPu8b7nrK0cYUYwOw5ZBBDZPk9g1
gqJeh0ZaXVBNU0x/bswLFopXqfPpEYnQELIENOax7wYpYdCyA8T8qAS4MohU5tyMCaajCQ52Sr5I
WPUZboLF1upLGoRpu+QwFCLeZ9N5i0ngSNBZQZdb3Jv1htV2RUCl4bVGnNwiq16NgLcNr4Xp55Kr
FUVkl6QM+w3edqAuu3MRQCVuQVmJ7r02FMXnpJO1Fh8BrY3zs7mY1cG0ykSTAfNf1JCIZ21SEUaI
mmcZ4opsF6A2m95MXz0z7gmKnaabsuFr5EQnUlF1NGromZ9hTJt+YEmUd1ljTmrJRQaVj+UgH7Z7
eavjxA1o2kqM26c7r297vDy4Jhh8u8CMa14K7psowrcfCIfPwQHYzpD5laKzwzm0GMDxsAvyzed3
pIbfx3gd8M4ny4ApaDrgoieb88ZS/AoffgCeQCfskqQATt3wUWf+IBM1qLpaBbnPQB2cYP39oVYD
SORqBPcS6c7AiNqosa3zuktBYxaqehofO7u/4vXXWba3Qb3Fl6h37xEqaj927QIRAocWnG3iDxs2
F2ddUTt3RxqSeR8EJEtgoq/9nacS0JvnL1ebgUC5ps7JQccSnOTUOanOYb2XhvIOHPjkB0B2lJe9
mlwiNo7+3yJoWizouWPQzqDPLVhobrlFy8138pZex67Yj8sq7glH+8nlWtuefIa0dCeR1TEiLXlO
1tgVxrIdIoQ4EzaCwZE4pECLU74ZremQXtOxDO5rXUZ0Ic7oHF82XOw1to993VjDHesUCVJJ2o+7
cAmYPSdri95RfyKBHzHteaQDgSjhOZ3Bwc/CIlLFL+QrcF1gOZKigMbB5oaSN6Xnkv4mVEKiRsxm
tkabwmTzP0s+rTHsSqK2pt2APw/fCPYrskrDwjT22pCogD+hmlsuPNlkFJobitPUpRsiiTpTAPZt
bHhw7WEy1JoOcRsutqnawcX9gSU5rVV4WxWaLuKZJgPllUz5BaCEk2uUrWbWx6P69qpfmAyF56cj
fLe5YOzpViVo/BRe4BL4v6Yis6HzxsaNwylayUA0oHIOc+DlpIUKS/y3R3yd5Dd5UJnKHf/TKkqM
Elh0iX4zDuSG0zgafJ3JJ87FkqO0bs3YG7OLF88Y5gvhOmtveCRgBWqMGjICz8zfh+FPNuybLGzl
UF34JE1zZOclo79nq1qz7YR5a3evz427YmqSiT/Q0/AAfy+ihPRqQ6A/DKqTuCwXkiq386Q8Rgm0
cL1NXp2oF7F54MTYjRHEVs/ksxs7lUdijVlDoDjeyJtBtbKle8oJJUfqd6sKOsMtapwEnQPkNYR6
hh9uyUitpifycCuoBtQnwFXSaPbGd52AA2SW0LfB58NuFDeW2E9xejgysz1YSjrdgVPXD9zpGSkH
xR2FeGRXeAv7YzLIttrTllJDIAUrrbuW0/U3a1ibNQHfFlTh3sRI1ofPTaX19dzLm9IWjcOf4ogZ
CstoJ8FSc8UAv/OlD/Rqrr1UvWJEQwe6Q1iu7Hu1fjwYQLyM395+YXWZdXOCPdE9sMM8IVwInM8E
NKmqp56wjYjQa+0lU4FFKEL7zqs5oCmenHq7JHb88Zz7j3LvvqnKuq4ZSNl4bng8pT+q5nypbznc
LzprjX2nFzO6SZyqbu4ER4fY5p4WXJ+0wt4nBoJaRntArKWwceoHOwr0VSCdmFYsUdJzygqudaem
7AsNg+NewLbxnrFrncLFRUIAGA3WDTWu/0bnZGDMOW/n4SWlh6MgwAIfph7F2+CYX3AAnHweVMnJ
Jdtf/jw7eaNiV256TLwq8Eu0H0BekNYGAlsA/XUByo/VUyZob8KrdbCAnAMwNx3bqtz1sfoafBlI
Xb+sfhFNueoaXLYWFlb76LgkKul1ErYL3cLFm1dv8pqAhCywFjr3qW+nGgjHEda59g7bzGPCovFq
cGrisiX4fu4P4ZYVvMBj6jn79RCRwIkXrfFpTTIotpSpfrJ6ztOpg6ujoO+NVYdSkVJRZYdPjR48
3aZzQKc+JpMV2U399fm5HX075/5QErVCCUHhLPz7h/qmOl2/pohYqK7l38jq2THjq4uq7sfnpmv1
lf8iTAKqRmf+UXJQ3cgkYXjs+Owup33ItNiAG4cux6HdlUxXiRniUTICbXFIb25kqiFOJD9aMsjU
p335qGARzU6brqSszwbawHWHdn9MW8Ae44dYUhoZsN3+jMx7YePOTS3imMpwpwO16zn1+/C24A2L
A2o0RzVYSDKvlwUS4Mzz1Ui4NTp35tnWZTqmr5SuKIYe39s4XIQ4kdF8GAs9ojUk0hBAaeuWb0H4
GYMr2Z8EiYqLXwKGnD9s6oj9nT9u2QradtUADgxvh+6APet9c1ESVMFdY5RFelOtBPyiymTe+oQ0
fp96aY1pGXgn+rAYD3vT+CVLNKxdoANaLR3eIlvXETiAxx4sSzkbmhvYd9d1PVZhB/EH8o9RcXui
eQOJYDxSJcYmRzPWJBEuL/WjtCiI0jyRMepxkAG1bzMpyvlmUKRh5QL1Rt+UbnufQ5sMHlUEQ4uE
HTUbf/PL9s/ZwtLJgzhheRvW74h8DqR3ZjUsKRXh82y0iw7ezJXN8nZmMAY3NwYUNYQBPOVoxyf/
P6dADIgG2vg/uNiTIpHeS0LrKl5NpJwWJvfdq6C009nqru3RHXyRzQBL84m0kaKjbJOmB2JXeo/0
1jGWOUa+71cG2ZhhJ/u8ROzQJuahOcT8u3QmH1Au+eP09z3XpFDghrlr7aoL0JDK069Ys1eok772
DAMfEWLYylifUBva/edPq1ZqPEig2ofo87a5Znwft7YelJRenFsjxc+8foPBLLZ1I0Z99RE6izpV
Se0Vf1wL3oOwsqFlZCn/PXgQnEIHIXDNmVBc8SfcYRwjtuC8vWzx3+FRGAeJGqSJd9quYrhT5Vka
nWXpt9Ph7tzlGAZnIlAdkAjD5JFJwqb7hniliJ+QpF7HSdLBwLUquBmSxcnPKd4AN9RWUmTNyQxk
FwNJD/AIItQQln0jdlou85oThVJAo0QYsuQ6vu3Ql28ZbVwVGQCs9S4VbWbaD08xMXydkVaUoTou
M/9J6TyP3vQhSARW7n8LwH/YtHybfIcmmi/lLEpQy/tdg1fHePwiXh9r7xmOiVr0q9Fid0L50sqg
TlOTj+NcHdpmIKSEghrV0XbPsjdWfzWyoj1GqMt7wHwNLlSyyTuBmv9U5XnrmRgJ1+sG0ggfN5+G
oMv24VKfqdEWfY1y06hN5KY7RrcSXoDeNiU4m4Lz3D4arjkshD9lF0ZZtkvJoRlBMt2+t+8CjpyL
jHqLl2eWfv/WVt6kFVYqprsftZY2o7qdUedb/ROVb/XyGbb90m7TzFfTczbNDiB6aRQASW4iHMpj
4mZI2efHFepwad2yTusOyFfrE4ILqJuuuuHE9T3sOcfU1aMeFmzYmEQGQrMVh1PAUlSzdwmoaY/L
4vYFDy79J55Ajx7ohB/4CzTrURrvC0ODGDtrn6jGYHJNxuITKl7tIJwHubBF0ep4zwx+XXZRX/nl
G/eahFrpqnTCjh/I45ND3Vl4WruJXL5Aw/daWRSgpwBT0WMBq6ZeHIm22qN/Ae6rITjAahRPTjS6
1YIy3AGrBRT1yL1Y2trAphRcPf131T5xNg2U5OcB1A21z3PsiPTcheR27/3ogAuwHl3EgPEA8I+h
rNdunBey0EwTvZR83fiC1Kxxny+qniBe5EWznblCZDSavRtFeTuZI0CZIoqTguoZHY2jfiGyt+0e
l3Plob4tio1+1agOLgug7XRYnjnFGvJqDPq6lZYL/dafuRXEWr6b88tOlssPOD6Ym6RvvEbncogC
wXvv9D1rP4OYonZKyHDwk9Blv5AKwvsq9+4FgNzzZgh1mQcO8YIkKc4umK963pqDerfY/PGmOYNC
L5FSxRN/2GyuuGB82ZETaUW7dWrYNytMbL4zY75fve+dJQltuCYw7ZQDYCk1PBFEWFcnSz86k+ja
ikYZn6kwSQ+QpuHZllMiou5F9/6/j+0fSzLGUeTsptb8SEwxvGtEqLvOWxYox78kgiU4yTd/advW
G810pcIxkX3gc1OZwWZvedJ/QyGYx/W1qRYI/eIEMDrcHOQ7/dWgKRnzmQIqjV1GI+OMV1MP0lVc
VLOwYTpiQPQ93cvV0N+iKBqmlnpGAw2l3YmLIi2CAUNMflfzvDI9FsnmbU0FXzdeKTtNiO3zzU8k
JKVkVASBxH58MXXjFTVuo6CbOztp9LRawA/0SAAO5LTIgtVwkyRZQfcE/JyA4po/7lZXr77e4zUn
O4cXsTAfIWQEJEZvCxaMdakAZVHZhRbDuRK89/SlylYIT7yNx8jhkNnv9TMmNH6ArezcwgWorqsu
s0lcV4KKLx1IkoKzJcdbQni4UkbTdNpvutifpU6i1Ceg73cn1sFdKqHKoRt404DVe0rU/m0XBjoU
VPAp5SV5ReYnXAO8Jt+fAy1SJeLe3XlbyAuhgTxJI2adLcA9SKWiIKLVu2W9BBXyVTDQbfE+FRrP
4Hjz0/XlZOT2/1FABcdgzAW7On10IU3iz0Wf36TQmiWKOmxDA6BzlSps1zBvj34WZpDl7d6SbehK
0w1GCfJSst/tS3zcTWpKHGcmRqCN0akDsoYz6tBsuyGinqWQ4th9N1k3cFhrrQr3J7MR8mSUQu8N
Vxv7kZrqhumImNP3edM0RyqzpmVgAL8364X5FTFkT3z1CiwyCDy7xf+KphP3NC2rqSykNAeCfEvn
wLC2kO/pmZLe1KcVa8388UbfT9Jf3D+dmfRcPe1yId8v0VJwsiJWUdsEjMELMMp2JY3z2e2EXGWT
0odAb+kyIs+6/GO3+bzYcbl7y0nlofDx4chPMBbyfjVEVdRxaFSdLAJvF64F/blmZVsMt32bxl4B
9VMa/Kqa5zliRZOz776SntjG8QRRWyyBncq6QbRmrMLK1zzzwlVnuQHi91BpX2UBB9u1ZohKSGPM
qlVFBX2iNm4nvEkwjTMEg1p5SBgikBz0cjb7kZOAxob31xaAFQUSo97uoeJ2+/bnslCBqhASFa+o
MBYO4u3bYJh98b6nGRChNi3xEl7hyC3r+WVcKea3HNi7Z1uSODrka0Y5SEJ0ENMlj9wV7DhzJ8pq
1yAvbCa4GiHLjERojxLpjApWtQLwR2O0b+/l5+pf5dGK2MAe9t8NXak3oLtrwsRuZU0SKtw05lrh
NLTRmhqcvgLYADvOflHkFn7Mb0m/zEhfRbSW6BcvEmuYJIOdex9XAk8jV7wI+rdnWW5pIbFkMp8b
4mH7tFyl0fk972Q3vqFWcBTnc/BeUqP2X0yREH7mq4bpEpBeQEUI1+HX1RX7/uFA4IH5yS82vaOw
p4o/wWAnwMIhAI8KJLoqaODCivS5134MAxfiZsCRCwFM/mRNBIMlJlWDAh/VTDV58tIzby4qHze9
EhTdXlI2FDyid6ob/sLEZRJE3Zuh4cu6yrR33ozQbmG9N1h4Hganrl1I/H/+Dfqsn5EQEqe7Sw5k
12gnu3WEbSwnq8gfFGmYraEbuiZKO/2mOI0urnQZLjQ5LG8h3HBmr0TX+Pl6YPX1TmnrjxBxuH8Z
s0/1JFaYsgsIkRDE4rEfMCAHVfIsZJakVB3gHRcyitxLenA8a8lp/8DkpJoNmzEiV3S3Ip7nihuR
s+CQtLI/uUNKeTEcNjUUOKQUO+Jse96k5d+65gTc4rYXaXFZ/AoyhgRilv5XxPtAuO/1O1RszLHq
07/BDE5zasayVcXYtoLtnjUKgFZkZLG/mIoUo8uTfepIW3INEH/mIwFmwNIa2h4SXDFgEgm29Wkn
2dkN2fcFJ8zIAlQhYzFWaGQEdlLHzv1L55hVEpSYDzMPWrGAizntHBg3T2Vvy2uBSI22Btsd0QTa
bCk+yOtJPbytiVLVYt1sJBc8JH/S7CezhVFP2WfpQKf/ZYQa8wYXHXYKLi9XwapeLSQ1UdfHwC8I
je+93yKPd1r1+bZ/5ZIy8OZrqDg2ovC7ZG7LCx14ME8n/4fxpTPpbtdsPwVhxRn5KE43xktYA73c
mFtgsYdgdg6p5sgdeG5SR1WaZnQY6xF2k71U8ve26TVMfTZwESxpjHCNE1TgWfRzgfYyjRD7ffZJ
x0gm9vUS0vfE/LSyUmCnu6e607fBs5HdvulK+DuMdU0PmgKFiMRnA+MbvLXPggEtL65NWmUphhSe
n8kHU5lYCKR12Av6K00toquSHDeK2LZN3mbS0FOn5qfkBqeB4iMDn6EFTWsl/LnyNRfYi0KadpMp
16WNpnkfLGgwbh9pJ9yexAS33CSK4BScGhZQ0EhqOZT5OXr7pTGSSAd4xL/y6J4mnqNMp7XN9qBW
hCrx8gyEOys9drIQZB5YlYLHgHE6ytrn+Cn8QXpDyUs4+XBoVGwWgGoq3LCbWBduwFoJi0uHxhdW
8OoGO5LvXOLmI9lVTryKbjQ31d11l4J92NU1sh4ES0y19nWdUiInUk8JUJmOf/3af/fF7Dum4vle
Cv4MZ4EDYI3fYxerXfwuzW14m7V3W8SJsJJ7hdQOOb76mXTJZMHMS056dihpQhSxsTiuRiSW8SGs
UKnq3M8gb1obiC/ZBxqVez54x1g/YOHZMEniUjwA/s3Rf/hKqC8+HGpU0Wwa/l5shaZs+W5p3osi
L10FFBNWZLTgBKW3lskgv3etwX2q+2zAOvuyKLUdCLK9uqxrL8zu3btNLQEb8mGJRH+3f+ndd8nR
PoCMGPIwlcAbBM+HmD+LoTsZiyIu3bLMF4ddOE73UAogOqz4uf4MDEI3sV1gZ3fVmA8hMbSXz6Oh
bBvfzAiVzcy0L9/WrAd+4+EgMHF+P0+X7OrkS5XUNmkknzoecvkq/jALafH8Vmp/qMjHtZujn3Df
p51iuTPb4srIQRs5rnY5rGO9AalCnfaGjd6getAexWFfWQYF+6HihH3KWm7w/0VYkJD1bcQXhL2o
TdL/wH7jYAtg1KeVuWTVeOynvRTBBxVSefXZ/IW4FF6P31zqh2Y+ncq6HlZo24O4WmpYsa2mbXR8
Mf2QpCyj2sJwna4QegjNubyW0N5NahA1BjGWK+NOBXP2//EN3Rmnv4/vP8NWfnN4AR6b6YZcbPzV
7iQKbeYfSLe1KaIeWeRxkcV78pzwm896NttTZWgIQsEaooYQdzhBRIN8pYmR4zum6BjwSY8kqy1g
+VBOQbFEmpP+6h0MlKBo7gX7kEKS6+iRyNZZkua2f/9q+t0zNTwQs6FWvinzIYcGmoZ2TC4Ra3P4
LRxm9WUJwntntDFXsMPpYYZwb5IH5PPlvf5uCOBGYUTXhkCw494mzrs2SVJTN1Pzni+ZDhdPmte4
jhKjYk3IF3PaglBmb8Qjo6Ugmsd71DMf6suTGEO4wEpvO8Pn7Tg1vp5nOBaKWoaBpkwtCwDPLt+T
Ysrx3pBe5r/AJCbDnthHdVf31xj/b248Oi+LNp/vadrHY4ZoNeHYXE5Z9GNlzDikpZHdAOjWZSE/
vouWXnKDsaHWMJUzaF3ETkc0Me9iovrLNVpgZKMiN5sjKB46MUoiT170cMQwzyC4nc3Uw+8sv+O+
fhFnAM95Gf7dLFtZJoixvFfDptGlFoRcprJ8kykg+zMGzd/SxZG1wFydwHobaqsAkJprR0KxSNV7
NG1y87fXprNaLpwsi7HmWzdRgewNaduxSnn4yPR6ngqipYUnXLXAbRk7WyXDoR0N4ChE9gKQ6xaw
Ax6Z96fB7OuWG5hwM45LRiqattUzK0hHaKFLePeAbN7Ac0uj2brRXfbmUFmPPmAfdgBlKWKJxpOP
rJjpB49SXfnPkWfcEBST8blxH4Zwsw8w13NsqdlHB9XDKzm/l4ydnqtAXEdtlLCpdE/ZHUwKZ6pL
q0eOJGu8hFYTtXYZo7atJtvj5LuBdLsA289UY1jLCkgW0VaxX0wnJ/sTZgQG0p+qCMsLYP3VYpFQ
oXpDNiCFAcTwwG4sZClvKeXyMpuGoA+p1ya286F1aQ3pHXG8cS14mplkeiPm+YsFkupL93IZLhdS
1CRpklbWEeb9knVJv+CnP3Jj/jPjNk3XTqkyHmzob6rgInWCZwN4j40lfcFBvlUC0ly0BDqL0qQc
bR8n8wXdgiAVtGBFZ5CXHTVEdnSQRqgqwsM/a58D6qUORAEMZv79Xn+W3KHWzSmZm9GoZ2lBxXV8
uBs7gcu/TklxMgmzqrKXPPQ71lR0SRB6tUChET1ziYLe9v4QBoB51251qHMa0fGFzwBl/hXi9POE
ug2VxblIo4TfA6wtxHDR4335ydr4m6cFBnmRHW5Dn+q2F4lmkShcjnBiY9eiSYszz4ghmv05pwpp
UhQZFflP4RABChDFmwSViM3ZnT91gSqAhzKdaVFK8RQSDBCGmemjLXu1O/0rdrJDhpv65mkNztRo
wKrH6XKZtYcbNuzgBaj6Eb08HKfoeW/odpFjbHqCiAFnfllx19LWYJ4lrREuBUjBvP1SrYDPQ8Ud
S7EPlpdq8jJJvyW+2nwn7Xlhc3Yr2wJKBKccnZiWZKXmNK9EwNe0XDIQUrfidGi+s0dJ9TaZNAn0
42xiKFBobbsz1J343xEg0aZf2fok01SUep8/8JRYgIFReT1jzWRgfaa5n05hDZIODObbSKLVl11u
8nMG5lphEzH59l3Qlq/qKIkZXV2cAawVJIB49k65KoUibkOrU9jN03wuhGtA5z+Di+4cs9PATdl+
qqEEPu1iuCG3t3A+yfG6ZpPzBulJ+Xs4a0IysD40UPXaMJzBJtPI1cYltsSeT6G6Bj/qblcXRxQg
0yaMIZl8qYfgGlHull+o2ObPjp8XNC6siqMKHNyFlLP8KuoX8VtSS7xLsd/e9wt4H4WNVu9ROjeM
LNHXM2VNalQ052edld7fS2gEJAnPf6+/uALlHGMmJ8z4l2DYxMclf0DjsPShIGqJo/hbOL6zYC6f
zZwJWD/8UYNZlWSByko4pRRvIaqsjD/xKzEELGdSyyDUcQphFOE6aYyDcakAuW8Le6FDuNUmHNnQ
qkWyis90z+ai5RZFgJc4OzwueYDTqQHPzqo+idOvpEM8Ye3dpnXUHcbODdzrE++zPuQJ5ls5SlHv
ObzWQHjBIPsfKIsOCfRvtaTmTyHqHHPId8o1ucSuoHmEmNb+JpzglEULtSg2CqLgtTyai/Jsyhns
fBZtuKZF37Ch8y42+6ic8OjZjWo0WM3nLdA8eXRKVlKA2lcgHn8dxUZvBoSZ7dbmvhE/pd/L9tID
zmMGEBVXorJ9uPWgMdn1yrIBZ1SE3zSF2AFsrRXE6GLZ4L3TsiA54CwIpROPZtcn/9y6lBhbK2SY
jJfwBPNI8kHhIiwDQE3XHWAZycOEP9ZuA4qc6HSP7/mvSP1cjeih7HpGD63uFxbcuU76qJDIB41a
lc6Zx0euSs94H45pMGLw3+2XaGizPLYAXK/o0/FiMIhFT+Xw51tDKcCIvws+xAhf9lfYHTRt3vHE
zAwUI/quZ3mSKzEqb6umtwQF/9CfP8NbY0JkQc8EBqm88AjKDqFVla0HEa5KoTI21lr4b/hUDXPA
yZI6GsPHWIZJPmRm2PpNTyKJ5Wt1HhbylWIeRKemEk156qk4a7BXrsfAu7sETK8MQsSqNQ/LuHwy
k3AuWSwT4IZuJjRGZXmn0XbUQBiSl/iegbrXhAKFOvSgZQ9k6afXX+M4V/CehZl4ugmCvo4hzYuw
oKW8SXmSznNURsuclznITnQ6KAygTsPNkv9sy3c7vzQHF9/1PvZwXwlO3EdeTXaKx9RCX55TFziS
vxx1vjRW/X/7S9S4TMIHMSy4LOmX/+g0rLYrRTARqEfzHKRNmWLLacElIKQXQiK2+AGj0e7CnumG
i+K0g9IfePEXjyQuPuI/ukfdkEtjwk05gKWBXp/ueiYKg9bE6AzhgfWFJ2vZb4pyYB+f2Jg/9nfU
p9Fdf6k6wcLkTvHcfY4h26fFMnNId3bVgpMaHPhZeb/pdcYLZ1VGekVwuZqfXYwI74dNNaLFAdUG
dmokOG5cCo6CLhhyC+1BD+m3xF42FXlQiXweOaMR1nZhpBYyftyY6DpCf4MwcVJklTpx0Lec2mi6
Nzq1G2R0hkuCrga4cNA4XbyvT7mgKM9I1mU2Y3PML5DnBCf+HInzOkKotNstMp1MSr8bRq0WvRDx
oBsSChZ9rNJNft5WhGRk2wsRC3shkTeBdh/brR6qHxwZOMZem2RTwffPVMph95I9eP91P3wieUtU
7U6P7SUs0wqYqxSxTRx1Tfp12/NwhY/aYqxqX2v0L+QNtnuq+3QsX2g+QIg2gz0a15TgwGap4s4h
3l12NcLecjftSNdOAkEQ0ToCy+rU7pbw1C8GrIl8Y0+Ld44u64O0Gml6DrGa/DCJ2P4D+yXD+4Tu
1DFCYkuHCcqzsfCynRJhXMC/YKegnbqHXhLfrrdLkzP5NcsxqPk0/s2GVQ2SL/0KIYzyJ7y70ufl
ca/bRqgsgpMp+ibA+gJ05ODFkZaLW0pMIhrG0uIg+J3y/UnBki4dJ8Pk4Ys1ACU5anDtAwjAfj+y
VAlCoAPJ4v01g8Ra00S2MLR3DXHL4cQgCK7qBWlxtd6XQv3F9q9HH4QLB6NjpCwDIT0AAExP8L3E
D7ySnlyj5Ba4jqEwKyS8aUBtlwqmS6cLqC2PTD+kloaLyzb5p7NI6G2DXeSRuP85CsQvYaFTJQRo
idBctDg438arKoBAgslN59VFL3gA0+ZJ41Vr40aYTo49tly+TjRTR7wlE7uMqHeZsrQ0wFNKNdbk
6uW139QWOTUMqmBqzcSM6TkcjKMoMCMkpfIbQdYJJBO2QJb136JAdYT4hWAvhNDOnp67FD9vFXMo
lu5eKnC56WEIH0uNkVGL44Fyw2MVzkisWemclIqouc5H9t+cIv/80ZS7f63yhj3AlSC3jbsS8Ryl
7aHmHqqAFuWt1sFj1DQ97bmywCpxu1LoL54AdYW95D3YD/Krl5gQary+EMWZoADwuLWx3XGQ8HCn
UvJSvCbJS1SY+buR7KjMR2HsGqiUT01tT4YqsvhcTWNGEr6bR7J35glBSR028bMrK0nw/JJm1V52
wT4TRn9Tq4XEL3IaLr3h+2es/BQ4m/tEDGYuGts5hfI+7wVPu1rlTeps7KcaCRqAqdV9ROlH8b1T
NKH9OYLSCplUe54FLOZNXGI9nMjO8KawagJTLWGmkkQFuZTJ6MYE3cP8JFY9v4jtZDeP90aHtfjW
whSdgcpicbT6Se+6c/nyCgb9zfCtxccvP0QT9BG0RrgI8nmNI8OR24RjHXOC7u5uwu5AbFDlHdrr
BkDAUEb6lD/zddD3CEQ2VlYu0yHiaAbp60eTO+obUbHvEd27iUZV3i+Wv3rxUGW0xftLvMdTek/6
fDeYHCVScgxvVJddmgqIkOCsGR0Zkj/tCBgP4/n9tLp2OVls3D36zsYeYo5aBymxMyejuit+SEWd
T4gRTpSjTV8PlHOCeJQ7gpDPZZ5YutSRCDox4HfYija9sayoZ+cI42ccrj8ta1BWGR2d21+Z3mHr
CvPgpkxTfyN2V1EZk1I2WfL7NevLtcYHh3c53y1PCDxoZsuXsRRsAnwceWsVqFCs0unhXcHhZBJj
wHx9ldK99MzHOMHo9Eep35PDd2gNyKDznPX+v2LCITsdIyfy5lFSDruK9QwZ+ixe7mSRce+kZApH
GfYInLJN5fs/dTO9b7NjsRTZzSH7vIlsQ9hYTgpw95ZND77sHLHt87mwyqL9ygJZt2uD9TfKykLv
k3Uj/xymmJb3xad6DdIJeGjCzGA2BkpKE5WrIxW7MgjZnuAYoPVyBGMnaTZ7+iefDN1UyEeb57tN
TK+LzwCCU0fIOURpiAbIRf1lPex614ve/YwxMzuk8Blim4nG4obqAFL/+FxqrKUXiUH+0DlTDpkM
m9RZfBwyowwJndw9JB/xc0AKfc6lvW1bvfHmI0cOdbO7XQKa2e4LPgVDNQAJ8pIx8MLb0h7POqDT
Fw4G8e5MMS6wCoBMbOk/UaqNmmO5Iqm29P6Uvm9ye4xV/vvS5uloyKCj+7+c1jIm9cn2G5IxLNLF
UUeQ4OSWoYn9UNkHd3pgaG5ib/XvAmoQEOMTsuuRmTc6XC7vKsN17DwaW1+awLfvvQ0jUnEkE6zd
QR8xpBMw4MiHJgRUg8/1bP1IDmRgl5bwS9qxZXn36TJRFfdR3jbefa0FLDeACOz08IBtAvtLAJGx
Rc14mE5YEeL4l4pA+litJ2hlF8cDppSXGeY8OL0GKvCAhWQ10nZ8x6qedDNwCd08NSsQ/JM230zI
ZeTL0UY6rZmgiaPzIH2AeUesSWFImqRNjxLUqqtSObnixJHCZIo7IBYV0cV4UfXawp4+bq8zhfzc
XTT6hAj3LMSOL7/g2N2A9m74NPJqz9Vp9hK64lhAlF6KWHHziQrN2KboOP9GKJA2gjJ3kmpPH4Tr
P0osspSGSOsIGju7tikaE/c4twmmcveGbmmBB1mLgzsmTqzJX0c6bY+46/q9rGLsvMLQNOOp3YTo
joSxU0EyReDxFDhGlJwunPlZC1MKzy6T+Gjv3+o7VAfUZNdDb+WGrdQnPqsGIcMz5ROnZnlpBr/t
2X5gAuiky+P7OHoK+oK4AMg0bFotXJKRdjTp4S2rxOMvzrlcp2oiWC7W1CxtO9PCTKZnYG015ygJ
2GVnez4ZDg2ZgkXWMtwjAOztUBnYL+Ct7f0dAr8IiLO29Dpm0R89LwRSBffU567vQXNIcJQYbksr
KfTO/pAgORU6WKRh4SYqdAU5C7jYiEFreMvebrtFJCUXKj73LIRNkhvn83p3BLhioPBkwES6eOTc
QnMZRHndlCXkkwpcFYO7MYe1KAsF5nta4cDv+aXzOm6fhRe6ls4qz2nYsG2pSkRQR/Qco9wPeRnz
TmLZ68yUOO/eHtMXNiDa9HcH0FHWnbBHIx3wEQcI6gIUZ6PUpEtk8fSAJB6WlHhIVVnX/M8fCaRP
OwtwSEEs8lTUTqPPYFU0YI8f00zqXDwy7Cm52ROiHzohuym9zguNzS4c5S7AWgNAVPkN4MJr+xCk
ZQ0Hxox/Qu7lQdY8jtKBpVEN6fDMXpaJlbflXVIK7ulzPmBVRasKDUWCJtRP5kkVIQF7K1GqHYXG
XHzNeSX3tgA925dM07z5vrFsvUp7hoDwllZ7BdgNj+sQVGpSzyLdC9mf5tHL/HXl/xm+mMQQleLK
Hu11x9t9kYQmO9XJOf2C8ioXr5WZhzGzqVG2cXDYHMSn3SGZfduhPV+VFyvr4a5J6tdfjButcIz5
k1nAl6nvBPmBaNxPZZNF1rxdcBWnvSOw5b3U9pqy+HlQousNDW/RO6O2/houjLofmSuPRlV1VGEW
Ie+hKbkYtGt2mw0k2z0R8gaNP+j+kDCgwh2IeINtnSBUthL4dFD7coSMksT42Bfw8rweIi2Rbt2L
tEgBwoAMcFbpmC2YErUtP3DUzmGdfyWFul4oa8+BIKk0ktyzEEY8e/hRgsMXYiZDYp3oOQchF/pa
Kg1eBAT7Le20VefZ51UukM4CapPDKBjF9qzBRvMvtyvD1M2NsKQgB7C4BzRiXRETpehStai0mRRK
/Fkyc7vOOZ5kOHmiXTuXHZH8TI9Dwk30dyh1ReIsNCnNThUHfCF/PSXrD/zBG7pT8hnCJPVizk3n
ntCDIqOajk4w9gFQUeHxHm6VXOWrl2fyJPl9UJqUc8F20arJLb28JI75Eg6f3lkY7IzcxILxCA9j
DO9e4pvB/QLnG7VmK9zmIHl2G6fIeuhG0311nm7VhA2PicDpPo/YlScA3+5PNW6id+3C/P7LtWlp
90ROtupwSZThHGjQ+Rf7OY8u0p7D4ahK8EsKpeN+gwyBvU0Wq81J1De++MxR4fJSdxrXcw3lFcGL
v8lvV6psBbigPQ4KY64tDiGFXXUfOa13bUOHhyCsBkDTRhJQv60vAJpgV3InJvDX+1GkeY6BTdrg
F6dqHpUor4fhWgBFkQXcigPrhE7xMIyXcCCOhIRpZwfa+hV0rrlomINeDsbvmnZIJoDBx0l4lwOo
D5o9rEd4dlTJGbIkJ+Dw2TT9EznUdWI3SEPe548LKZ0Z+jeEFhcwobBoU12DHfu0Zle/0yJnQ7Sj
aAUXln0bGbNiDrWY
`protect end_protected

-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NHZ7OTFJ2nLlWz6LcZb/7CIFRKwP9WYIHXBr/HT92WDdHPeLhPK4G6jZGu8Kw3ZlTkrO5uNtqS8L
GbzYqFuwb9eTiio5SDMupdv6L/ZIA9t5R8Kf30uNgZuxGROOx5/Q7xjSdVl0U93v0W4GOiIi6jNQ
FPhMO9bLbCmQfk2J200ETezEES28Rz5L25CmkSv1lREpaD7ud/0iQESWqijzfTsPL3xXCv3StzLW
j0r/SwKthz/PrGrtsBLD7RirDM5ytAnwxEquvm4LTYLJ7uZlImwqvTqi4BFT5Kdgb24Lk3R+fizD
f8K7lfVXAe1BXNnOkzU3gLlgHmVZ+jR/XlTSvA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 71328)
`protect data_block
jTIbdAJycChI2YBuupHRKlNdf7lE7LxKs9eUr1saXiRoPVTpnDPC6ZRnBw/EO1p0Ebar6AVedPQW
DF8PkacsnAl0UoO7LxTMa4zpIezlV6X3QQmGXXTzHrdFSPyecQyhi2AE+mdvL/0be7zeaGgM4sgP
HDt4bNDERPz96SJILiaBPG4ZlG0I2ca0aSBd97lU5EzG6nXowZ3BCLa27O4k17MoM9fPbYsZd5ZP
mLoLpS/dp7jAfPcXlSnmbF2C/pJTDR1NWERd1v5E3LdlAPFIWtZGmxrZOhQW6Fis17NhosBdneph
90elVhKfsBsps8PNhLNr88gik1N0bSLbq8LldDXFSJ8AlPMMe+kfMZbqa7ggfd0Qdv5tNC/jf3H7
XctO7sl52B0Sgh7QNOq4EDuIULcDXCks1VVls52TnAIRE1FhMHtk4xxLpSTtsSxj+Ej5k99yUNU3
kSWrrnbeizOVfOo+Jw5vmttPFnjZg+AgKYwd1mDnMoSnka3F0+FDQWIElToULoX/cikTMExr4bUQ
fEB7CIQQGgRRCehJ8sA0HIVzP1KQ2J9bFLCqwq7vexDDmNTHp3qRqQyzKTucezJ+rdGi/2Xz9YpD
u20QyNviX5KhpUalT+8d8kfkG5LT5SbgRhEU6+8zD+ODfqjToTbzNHInMy9YDLJRmWCzgjPNb/xv
MiS2Ug99T5j8/p/torFIG6jtMNkWmOo5Z6pD4yHnLKY3WGWOfoZXQvBpS34JyW3HCKmU26L9xWAV
rorNTF52ndPgcFcImUM4tGrMG+ZTk360e07EmEhKh19AziQB5EjAs0vYYaokXj4voQNZVoEP556m
jK3ygdAENSa602JJFAUsL63Sz56H9jUunbo61M4XoFyHd66pV7Wz+J3jTOTWSNjmgTINqiOjidJb
OI8OXX2SxWo2gf5pY+EPrqyKJttWzcGkB+QQatcz0jwGzsby4k+upj0b8ykntFcrFiEUbJjnqtV8
KKDAKfrhXGufo4oNsT+ODFF2StNOaTlaXYAxLbZ7yM/T18TCBipohKPvjIVNBgNIUdxWabZRs+7j
eQA1shocJA8g4aKt4jq3IRAzJuEKph1vAwRcyiqQVybTJCvCQwmad3fYsv3PP8ZQIYPU3G/Lnu2F
kOzJGn0W6CCjbcAKVHycWd3p8UZb0XqqAY3SKGy1JOxChxFr2h9rwCwof9SUZTR1Q8Zsxhy9SMp4
ltQ2ugzWUhk4ySol2NC77Z28SnLUa9z4oqx1LPOBRTVvzJV5oczLrer8Vu94wvIyYyt7gr0lOpVQ
KXSJD3LNvdnh92VF+OsIifL5Q336zjNwXSYPvCoI3zmIRDmQjJQuf17LkZygvUj9aCp/3eMLO6Ht
2x+ChkbRouA00yH8yOVwqmswXM6G6sitD0A73kOcw6yayYgGUackIZeXoHoRpIpDofev6B1Zkj5E
Z30vKGP+jYoL53oQtoCthX7zbdWu2zl7OrwwIdaqExZC6H19ZzvXAQBGpCFEv9B8Xax1YHjdO6dk
eLNRXj1CB9amO26cT1sPxqKbJca+VuB2IvVQyPuOXQC9pSANV6U7J+MJkL7ijtb1U2j8+1/bM8j9
IqkNuSER5Pr13SpO6hQL+3wknJobAMbyoiXMyoh32r1A7vF1WFDkiMaa/0smyaDldClJ0dNlSgPR
QwAnQl0SODGM5U748dkkhPY6sm3kcySdKrfL/P0/uwFVjB1IhrVhX+L0LKQj2pObvpAQ+FMcm7sN
43EDbTLIGxRwuUiB96gg1/vC2eMgJJv1/9w7QKQHrl+TNqWdwDQrPSOImgZnX6G9NtOYc7HMvn6v
4bRh9MVYGFP/IsujRbVO7ulfdTCZbDxZwGr3Fomkxki2bVZ6Frhr/I6EDF+I8I4s5NezXZ6OZHP7
9xS4QFs4V5uk5g9ml2QtaVNaPCyajfm+aYhltGZNXwEGZQHGJMbrI4O4mF/gREDQxm6QwGal+Qs7
vxSyeoBMOPN79nnC/4xcJJkdNzHjoGgoQJvjdb7DD060TfkAG4kyDgO2tfkXyGMD1tlIQNYjXtep
yKxEOCQoRcOdxYGVlUtfJRfpLKoY+XmUmP2eKmwJes08mwtSQjpRsGKmMBoQsRIKsnZkSAp7loSQ
e8E632ZxIacIZjFkC/X1En+45CL7kl0sqhGEQIHIK6Et9mtgoUb3/7O6DHhgO5iTtpkVvov+oIi6
q+KYxpqcM9Vwvwwwoq3YV8FZVxYr9qVmyEEgwKGVlgBYr9w+1RWQZOQKCxoviGx8GSr3d74aOFUB
C9vNez0b9f78azpLgpmBLWelJTNnyi3UsYnqCcNAUNJZWHS35vT7AxzWZc3I0GpguJHGlw0rICTx
nQlOE0HgBe6IT1WM4Zq74vLo127aagjPas5RFj3F26wOqOROfx3yKMH77NAhfOa8f1r//kD4kWVT
jLogHqhlEUoEUehJHnPQ3aF4518JHPAVA9txdaoM8ST4e/hIUKl/lcpT8kFeOdkMM4teVCPU1Pb/
wB6Ssf7LoInZNCsPPApdvq5WS6zhBpw/QZOTPDgBsTx0t9o+OUhGEw88zRAvU/qgg/vkS/O31J1B
ILo0ssr7ilg46m9k0PyiPPg7sHzI0v+PGU/K0f5j+zO/6jOq6u3lbpmwGdU7reA6VuQOf596ek1J
MsYweuX7CmqHIy5DphfJN8JlXZ9Oajq2UnNF4A64u1mH8du/q5SCCBvJtwmW48L0eObn2F0LVMeK
TZTgesZr6bjy9G3n4feWIVpx15RwwnZ/bnGcl/86KjkIZwO+dyi1RTRTuB5UCt0g9oqlUWt8uWV6
McOP6g/NZtKkvTot24sa11sitXY/QV9nWkgfk72Z3FHaLX5WQarJrMUCFVIQOAn1cWeA+FFe3UYl
V4BagA2irmHTA7/c3JT6SJdHokx6LDVTzQxvWmAz4fsMGAravgOQ0s/nVW/neFPFJ8qiQYo3CD/D
fw1r3h0OATYnc0WeSJf0fjZiHpgLISR2wD4T5TPyWIVlABthTSjLP7Tsvx4h4dDBb536He+jLjyV
9eqgCbraZr6Oa/x0qRhkdegmjVYDmncHXqCSF36uTxew5QCxS5CzvzNA3JqoypnTNG/wPtzoDnQf
5OUpQniF81BOko7d9u+pptkqaTkNcvkM1zj3c0l9Hl9PlR1ixACJIT5nL2phbEiNdPBnSketlJrE
i4txFwQeMoKAbhmrcZor4Zu3F1lzecsIAvTM/l+LcmnQ90mNlqj2BLYyr91uO0MFIr//IgLBFB/2
5BZLfEkmyhfGfDydIHVVZq0bfjhjMooYHg1rodAgLYVjdvXJEPupfBcaE8JW8AuUFW5Az9jVFnAn
9RR5JET2Y3rIFbFb/aZDv5c4BU4VRUVlaAexUem6PCEJJJX0lfG6iYq6YBkIYcydWZm0JOIoYOl/
LNfhjFYrDRATdxLhH26Tyg3irXnZOHC7kyXb0XPVe9QaIj0os9Zn7sHjeV8HxC0BfdWDb/Y5LOhX
ZDnxQW02Uo90bf1BmRdhO2Ad6kOMyD6NvK8m2/fSTVemg3bojszo+EsZiRzMzFpvsc1GZIzNnPUF
784kXRAGmrH5KNQu0oG4US/p1eyU5MH6GVwLmvCgZy98Sv3j4tEzXf6xTxQvoH9P83NK1N5uFYQp
OjhLWCYoDQwITVNHlqnyEIaEp3yhGyDMTb+y+v7jk64m/PzsPN/8azdeQo1dPRgCAmgqBegZLalo
OlFHY0RKfJ/Jkx6qxU2umPE6LXmdFkjT0hcH59A++xyoCl772mNxDs1ttBclsvZJT478oANcdB5S
DBf+lVYOHCQvhw440cbn4mKRy1LGfn5758ZOdSexJhGHyIMSLfsGUeTR6q98pKmivLsFONHNQhPg
o7LyTdOUJfFfM2Hw3RPxQOiYYUZl8hcm1RD4flvvuxk3FMp1ejsTvvzkudhaOG2PL7n3nJypE+Ry
m2aaEhGq+eNEN4SWiMkiI7ML3tCHRW25tRzTRM7AemcTei60/8CCBvUOi7b1ID3VkssJipUzMYO4
j1AaNpHaWAyYezGa6CIdSf3hOtSK02gkv1t0C4HbtmDAST5wE7Qq8yFTfadpntwzyAG42CrraRCW
pmQQSdje/csXngOPiYY6VhzJl8MwvWtwrTk47blJhKDnavU9KYRrsklSXfJ/+V91Hgn8EV4st7sy
bBikOWdmGdPFwnWXq5QEYZm12g0c4BMKQ+ycvRO6Ba+8d3zeTZ9M/nqZxo6WPVWVMrdrr3zRgALg
fho62mtSXi0FgLYMQJMUMF66iaamjCxuUj0+ddH98Imzi2LWN+zhBUAaMDfLI0X9HH69NT4hTbAT
O3rI4OjlRHJGmlFF/edvtIGPVZY8ry6Z8+CqEsFSsu4KEWzSdxIyRIy3XaN1xoJLgnKKzfGKniHp
MGlNqyqRa46/A55I1Zn+Bjm1rURduiT6Q67kbJ4DU075OnQAFuDgrbJfMncaYjM6ynELxdgGVZ35
OvzXUxwS4S8VW3tPZm+MkRGDF5GG07CY6t4QjUIU/2vlVWPeONKuD5RQQC0DpVnSpu7md46uTgS3
ZhMf2JCVffK4csjV38buPuTO4GsIY8lS2RXmsDxDJVk19LhLKbP0XnA2Em6fG8l9KOx1R7Kiz111
8i2EE0SiMdDstDHSsm7HB7WtOp9FIRPKgFsVxBTqUjkpBZPUTJO47hTHTRLgcsjZgwMheVBs6SNv
Wm5XnsANcABl+WmMbhTkEqdkEkEZXVw8KsA3V19EWpHM2/Mt1BVPOjSoYl2CHxLHl86CEOsl3RMf
fP4fr0q663DPBbkQjuS7c36as8sMx3n37g0bZX2k3EOoBq2y5JE/uNAFE5u7Awg1qd49nO4gCdCO
L5VDzsB5D+bkZWls3qW8znzikBFuRxI/UBDbb9ILROJrfsSPfVp8lEz2G35H1UyerbOih6wd5wfC
EqWYhXoGmmeY1riNc21QX1m0FO1WIAtpHoElVCx+qOdQ9UiJ5n2FBpI/KWGI9xJsGPGf/ArVSCz9
SUFNmaiWtELFHKkNJBB/rB0/49t0NYusyaFF8nbiGIzqIA9o+d01vjRwfVzmHLuWbzNk1IkQivEq
4fVlDO5LBY3MVHbV1pqlMT6wety9kMWw/nmJpXH1Tzib0svanDGTuS53QjlSu+WsWUeCW2yIOvRj
/ezynpMUQUZTSvl4YWF5bdLheipdoo7Y7q5bEFPSMEqv/gHTL/U4NHHM8lf3zh3qRFClUvNtU3e3
Ygp/XRKGZ+zsE/nqHQChJvIMwtGiDTnjWa/rMyi9TfJFBGWEgAtX03CEerBGpkI4cxz20TGNqyGu
LrLKdiQFOdjyH2E7C877CDg6hrtwHNxrmdKUwWiZfG8Vo9NavVhOJbsVbpA1uHkJsePtGFR/ejqJ
XbCSdHLrBwtk5wGQw9RpnEm8rQW4zX2WKiRDAn9Rhxfk7L23oX+BkXfOEcbUdVdvadk6gNEl2oIi
h2ZdurVOzb60YTrXYbHhdtBosb1i168dcmHIOLnxX5L0W+xRAKwbzjpXhhnF56797y8B2wh4g6HM
LKBu9K/zpXmRnnRjmOaTl/79AT6uN0QGZoM/mlkMhhqGoUP0rMdUKiLQczIkdfZi86/9QvcSiac1
wccWqhaB8zory62cStR8Y1Qs38F6pqwRbSuRDdF2wWOZiZd+sWqslwCQOh8MGyZzwTUd+QIQdzHa
H7CY4aYUMDhgshku4K6tz/+m5xIkc6z1UfJSYNzYbRzQ6vLMpHxDPUseanaJsqfOcvUjtbSOxyDC
EKG2bbF0mj4egL1zc/m+KGMoF6a6UEOkKfnA+CJVhC/z9KtOnTE5tpkIotMgYj/z/ehIGHJJiTeY
nDkfXmGm2uBz6vCm1fYZHuzXAAOYKqsW49uJVjdvnUMwt+SM2XntZ+0t0S4XIjBh3fezAynMDCDy
bLCS0jdk6pZhqsKmmBzmtWAB0vdr7pJhGp9eVq2JvfnH/MwTvoG7prjKcLL5d/Or+Ve8Idhlu72s
XRYRoWb7TClBI1ajhqRNWjrbK5DKhD2wrAHdOQMCQ8lYw1OQ7giyhdfQIJ76enujiRJkASxQd4fq
QeHHdmWE1Rksdht/jhFnC5WljOTM2wpnHnVHYnHQ7wc2uiVEbV1higckgxAS7YGOwbb2gNoGotyd
VKhFAwXgwE8KqjyW8qe9MHi1bDHtHjaVDuPJnr/NTwy/uYCjeQaQ9oZ2mETmZUOeegRBy/dKQMzm
AxqdtUkWchDybSEqh4f3wYfwssvs3hrUTefzRIOM8jw/uvsGytgnRN3Wjp3VeWZoB4k8dfUX/8Uy
VXAFHkHyl9qWf5M0kK4CgS8lSxTvaChA/TAocOrpYPaZ3k64hdnBLXDu1l98uox+S2D3D3I6tOnv
Kft+ysj+uLqMHci0Ee6NG/JpQhXp9RAkseYXDRNbEh5q6BlCT0J8JlRBceZPXSZDwYbIW5AzaHDt
rd0vCdHaF+7hD5iuDgMT2EVxhJBC/LsaZPA1r6GRnqrklzI9I5BqInzHho0T1pFlQ64atEXj7j9D
7M1QtlAgsH79gUlDMIonz2HCz0sh07U2euITFvOo4biCc0vE+YjvX0Cr5zq+AQUQJfGDmRtYRiV9
4SU80eqh5Pn/pJV5+HXvSW4RJH36fqDqiBdq+Byzit/pxhSo8BY8TUot5k9bLFF2XFN56SKMPYmU
fKj1yMD1Tb8+ImIeXLLL9rVJ3m3cs73x0+5fI/o3rVXlpu17ER5Ub9psbtUE35XCof8wB7Xl23QJ
uYDa+N5+X/JAxQ7Z6zDpSw4F7otlOQxlQ6FKpI2Kg0P1Oa9n8c0IxmDSrU9ZRWseqye/LjEBwpuu
VRai9h3MkmOmMWJ3qg6j3+7hzoUctUZBHMh0kEI0cd1xkXr0kTYHj5uJv0l9MqQfIY7zUCZmsJQn
RI0vqeJQNlG00l2iUO8E9ezqWmGrPV5ysERkrTAshGWRkz0fpNnVo9wKXcDGvpH/iK+TOURngD12
Wfu4ttEr64A2vz7EuyR8vfvAGDE3INpN3aNQwyjY49EaXA0yfmerZ9bZ9ABUvHnKOX72G3zfyIse
LctKooYh4AdwTun4WxB/BEOmI1pn1Qa9LUZSjOyptgNpfRFzIRGjjoCAZhQOx3vGcaThqUSXwPgz
D34qLqezZv4m4UfD23gXxwl/lAan5JqVI2ejloV19YOJBdpMY2R52dCBN0lxukDRj84/y/6AkCls
hjx5JIdGsy892P+qH3SMp3WDB72dqe12MWg5TepkQQjz8iAHzqrQxa1vsiPgHDEDQtRdX051EXM6
8n9NaaCIxjeg9hWtbuIutyiyI+wCRjoXH5lC1KUPXnyf8qJr4lxvOwNa+O1jufA45e9sq2Xdr32r
HgoVa5ygULRafRMyn7+e5ziDEZQwdWUGPYOFFcPRN/msJjXE9zMyI89mFcsPFeYCvb2NuDOuKIy6
thSk4BxhXCF3YUU7UY6BEHHJLt14ANScSKdyLpL3p/b/Mg+XmWrh3yuYEG2eUzyGff/MS/DVxdDC
YtL4rbjCCZkYK0Z4GvNLUYT+M9sef63CIn7I0yDwBD1xGcH9ibud8xaQf7P9fyCC/YB/URNpMA2W
vksvTzIVtDBxRTDJ8VSxALiqzqWWfXl1CtYeGOdxfpZJWEnaqokBXNxq5807+Aajn3T5vC/gO3kI
CmVX36rMVQswN472h29jEeRxndBds8Tse4Gl6Zw+cBB9oIeMA0f3Xm34uY5IJIMFmGdRsb7BVTZ0
r9ysln8FKx7mR3Q4Pc+h6tU/xEV0ioNj4CPHeUgT4Vgqo7/i8L7iE1MEfQ/VU6Kqjj0tBErYxwUA
mh+uBU2MUeh4fifvA+R+SjPV+AJFEaVDa5jRXrcZMC56Ho4E+40MFDee6v+ulTaDAz80X0ynG8ET
My7cpjWgRYNsPifNLl54GYNm+t2AWmGp4FrK/KnFqdxc746uN2P+ptVN/FE+BrJOzh3GJNUHp9Ec
NlOyBXOrBvPE1Gjujkth9eF1v6cpXTz36fWYZ0rVBHlmxlRb8RW5gjD13fxGrXdMgIhtD20ossjt
IxDm0GEmnhvLerRJFWadc3IpC+SVA8y4atFuajYNpigimizEfRNbcWRZYQznJOyj83qWlUNzKf42
KO/YQ8sa8UIHXyQOv6zz9w/esEvG6DPMsJ7Yxe8T5LJNeBueHl9T27zVLWmk/De6dp+OzxunKvfw
3HPlmY1wpRujI4fmzxZTke8Lt3tBE5lNtG1zvMysCEFo7dmPgSJlYqo4u6wFK3t+kGRC5n1hss7a
ZCOQsJGkY9EXFn4mQAMfCnJt8Op0NN1i5f2eZbtyLeLboYUGkfFz2DpMVv6fyqRi9+KYTDShF39n
zAqASulR+00PqDe6jwsK/Ve1Xja7scWHJulgOk5/uq/pNQs3fIQJCpQvfC4E5YVCGk+N+yU9v2Vb
ZzYPzaNFO5R1qXgy+6adgbd/lEIsC6vnHo2m8uHnUZmSQB2BeID+GoJUGEY6JC7NSdUvH7OBIjKB
B0+G3DmOPeqlKdH9XOXT9VSyENuFzVYfXMLrGAxe/rGkhwsUwqEffEiFaVO2S37kDYtYHwDjQiDX
qSDPAbO6vq+3p1W4pYGX9fkswVrNLrKmJQSAxXiG3Gap1pzfP5Mpzj5Hr+ULXCZxtujhTpmMfZi9
JO+JxeTCjxOfkV675rL1NHuT4ujmncxVBGkb5mmFboo2lzCw0UvHD/+JzZWVtn5HbbPFF5s0GIea
0Ki0ZTInB1I0oy6SENksV24pJLSAzKZ6hs1OQKd0ek5E9Wu/AszYMeFA4OW7otLSqENJxfc2967n
wstb065JIckDSVs45/pLUChtR1LI0VIOnuMdOl7vMB7ELDkexBLf+uWabiiuA031HXnEqtq+snYK
ODUjfesWGbnd5F9dg2d8nN6aHtEUzy1Q8UzJlp9F5MBUjy4mUCiW+p+uzVw1gkkDliCi2GNGqtUn
Vv/FBz9H4jQHEt5Flb+IHDTMIO/jDgJVxqIbP/gZsG4Rl4ARL1vbBL+F44KBG6zoY3thExMUDZnH
t47zwYVgDnEbfz/CINV6pS1bHqam9rgdZ32M+gTENRyneEtrN9aIRMg4NhjoViBt2cG9q1feo7TX
HWSNVBPWLBsT/jR2z7zQnS/Hhuxp56FNk5wIdlRzpkZxGO36g75QxBA3KhkGf3XHsebcUOtwWipd
v/zCXn38rGwVSI/v/2ws9CD7bbKaQR9yen+b7rPvAG+IIOHSjziNQu5TpKi7c6fWuHPfB/LB10Yq
2jtseN8Czuzqn/hQG2fV6vga2scJeSWgkZXunCxZQTeL9jUa/uw/nSKo6LsGonbDpw+VNs56CbR7
a1WiE7+pd/9izvs5Tyvwq6v+wRlBuM7C24XvJUKNyvjkxXxhnjXaIdiFMy5Da1h8Ey6b2GvwG4/Z
epJFmkk/zblZX2ZUUF5WyY5JFST3STatfUfqAg+cUegVncQlr5f+2EcgkWvZq8YWGPZgrkQg7MfZ
jMkzaMpNaeWwPit3fjSUpbIRqz9e41kanQ0Iz/YlkHOPU+/t5Hd25MCl2+s4mM0NuoaUbQwy4mHZ
r5LeF++p2QRkgUVQ7OC7O48Wbq6MPzMI7gngyjlEGSrk8ZrsyEXJLuIB1ALOQ+wvXVKTBZQSFtXo
vsQXbp0dcnfYWiqyeaer3vyHXV+Njs0FOgRfmcwlVtknWxJh27MkRl36ynHPHCD7XnSL1a8gOJS8
c0SgoCSSXIzJdGATCR+CW/BaBUI8NoYfKA6tMTqNDpHgW57tazLzwijLNG1jGCmrOfd9AVM4CXG/
r8YoDB7GvkOJhCfRSI2t5K12vfCROF+NSvvxIWq1N0yMTEql3OOBslDyOFkxSb31kF6zBqWxjrus
M/q7JR/nw1WknAu9cY0YTbCCzFz0DBwWNb8cED5t2Wh8dW273oan/zagkmzpAwsI9aQ9xHF4sHsy
2Qiyu+YcXKl+YnSyHCwE/ZBzeHvd/OYPBQoFTV8dqDfwTpBQZZnqxqY8G4MQlf/02NGZ6aGV8A8t
w7FZngVn3DqmR+w+Q0YFgNY3FSFbl5byYWDuG9F6G5vHIsQdrZCALCwIpKSRoEU5i/nCzNjc3WNE
FkToJ0VlGolGxbdNzPAEwZ4S3A9n/iqR78axcPA4/6cMEHFnLWyDfHPQXiGG0hjENa5Z6yAtr0V6
Tu38lUDToTym12MnA2CuqbFNd2Cn+ApSh1WrQTnwv5bSIqu0w8jjT17gcyvHE4G8g4SEGJffbDnF
dBB3y622vQJcoSssTATYXY+losnkhYE6MVdv+eu68r3geePlliyzr2NXNBLc7X9bV8Tvikc2p18J
Q5iYvqBJhy0G/WGMFoDwKRi74FJilG07ajhuOdQkAOf4nHMLDgUapq2XwHph+HIp9ZsaciZFRia+
kmziSBbq52glG604vIqmwESU8Y20KoN3TZtyGLeh02AnAZFerv5H5nGJ0RkjNer3rnLCSvxzVQ2J
BJN89uvxwn0cIhrY8il/Nory4KzYqkk9kIqkzShX+yO2tmMousWJNR8XLIKBvT6RFAOigqMOKd3J
SPvl1/x2uB7BUKf8BFPud/R3hJIYDPxqWXSu/7PKVvmOT7eOGfdgT36Sj10CuRybwk4/CSahsANz
XusmBzzoBzTif6zetvFeDkps9FfjDZ1/crmwOpjBD8OiEZq/441d/riuaESFVn9nLR/qkoAA8Rl6
JlVy3F2rhiUhgnrDsIPv0ZFc6T3k72uQYKmaQh5vf9uczP1RSMPEgbIDww+W+zsPlTkq/txbKNiR
unmE4Tn2iBVCYnSQwxta6UGj6t3GFFhMroO5GZS6JRzRpkePvnu/w22G3gQdwiz2jdlckgKG0WHK
EkKSOLzy+BwIAPnP+yDVddDzFPV4ira2MUrKyl94w4AO3MbRLIFMZWQQK9GnhBxeA0EQo9OUoIwo
XawEvRgrii2iQwzIH7FfUg357P3OKHjVg+Ce0HfB8Gao6aQu2OguI5R4nc6VJQqzRM7Y0EVKtHgC
zeZCiK3HPcc5IZWLS4+Cgn/+8iPl1ZTYJnsFQjB/ltsA2wbtTBxUDe+bT5NH4b6PbQ/YQBbBUBMI
zKwH3c8dCQr9k2p4t42SjtkYzkhRLN1ZTKczLyh6ngENRlqxaGqQr/XnI6n+QqxC9vIgpp5/1BQT
9ZH79vD+G/bjxw7+u+oAHUV5fLMJ8siUCTOb8UJt4FDViKazA6A8iM0HEcw8LVC+aj/EAoHBdV0F
dZwhV+/f3/vdsmiSyV0D8Si/rZfGBiTZ5usduJo8iDg59txCm9esinnjtaKeGU7ZWAWAUITkV0WM
NLB2TPv5RPYTxT6CDfNAffmd3MbVohHnYU2iDx6UvenxWZMOCeByai+6I89gBt/SkKBg6xqdTZy8
hNffifW+Cte4/nqQqeWNNMIQIsqjunxwds+6HhgFQ2PoX+UkYDTeKwYnOm9CQ+c1Xw93fsUCyRCk
0xK3AFbSuCxnTqTvsiFpNG5cuLOeqy9na5S4jFwyH0RA5gDLlaiIzzfAJRkL8s/bGtNIV5klSb4C
c8y/JflFfICRBvQj4n7+mpOmuKjBxhttREUswCY2j7mhU4/GIi3m3wIi6yOVqZ4OIdZm+rtZabtU
uVKF3gnY0VaKkGJR3Lsj/HYiimUnfXtll1pDsSycMP/EslMrjV6bbNyDhr+zZ8ow48eEej43Bb1v
6vu34tikuiPf5RR3Ly8iHSgyoD0Eo6DRM5nbA4d4WuaqOJ97Ln/5jMs1lT6y1tqEHTxbWrz+NK+J
IOw1jyKQxX1J5jOdYQsU5uYGWJMB7EUqtFM8KuaxAV1WwDEt3NxYCAqrLxxdbyqKMeXfsZJKugBX
ZAkp4UnLGG2Eppe3O7PuC1CmrlOnLy8XZM2N0TDCQhCIY8AzOj+AyEoFsbhTdVTFU+OB+oGiQ4PZ
Pv1eWdbQjLA4/DDdrSDYD6LB4JplGv0W400YMnvGxkoiZI4iLUheTQZI3SD35nBLQkApoxfJjpen
D9mc1LLwXEcMKQSQkWwy0M2kYCXMTAqEs73Y1PxZe8j+FVVS6m2NZR39YfLuIWCSy9yrW4C2K62m
y89FptjobixsHh2r7XU9Rse4A2Y28WkUSgb6RKZXiXx79q3Kp5Qyf9IbHtJ7+txTmqCcwP8wAK58
vn6/F8ZuWO3FxE3FapiSlJrIqglqA23qKuWKlKyg7HRNZRyGx0iuPlBZQ1b21O2kU0VjKFKPCdwi
wLfWDDGAUFyvaKigCNZ1EUQQd9Wy441uCP9qbugACNX+lCyEQnGXrLnE/2gtQH3DCj0eVvkxmXcn
DIt9ElcicvaBMTRCxoSdbQfCLpVvWOzhutQnxFT5Bp9Cz+OJ5XzlrKWSZAKnG+JLWAuTjY3xDz9v
2KOULVuU1gIScG8KxL2PUBkRxFK0G3zIDWc0guU6GC5WBLOJWNTNDfZveT9Kbz03N2hOjZb4O2pF
GC0y639Wi51XtMZaIkROJMWpXYUpCwH9rXZHHJk6SimwZUNbghYONWNIaCPRh8Nfark2XP8ag1gq
em8+YNkhE4XHmuLaHuA7xxeYRvzZnTxuKY/BeEIMs8xJPcc/WpJ9qjnYH4INf/usqfYgsiKsIpsm
1S+5MJFJHmf8h4eWwGjwdbh/jtD265HAeEZVp1WU4qJzg4tzh2alr8tPfgj045Lo2lQ9yG/otVC/
dEsudGjFmEroXOubz4JstoWuHdJ6oBjsrILggCb3+S9Oxz0xIewzSiFo44JZao4GY8U/KyPnsDsJ
CV0D20zqRyiIlAdibomqwYKAO6okd+lykujUwJjIsDn0d1JmI1SnMIDK4mn9lGxJVB1jaj8nl4zK
7qv1BknAM9UV00bz/ALI+ma+x4UbnKYNGezL9FvPnosR3XELHTUGh/cUhgT45zQpKsFalIREHZXX
6bhLHvJrykKT30N1ZFgsLmCzI7HpPBnEW/PwOtL2xHo85uehDi+g/LFUqEwrbLA/h0DWp7wq88OF
ocpLhrlBe0y/jMw5Ugg+77fWf9N9pXeIKmJjB9153++ddtauPuOgIeNLGfdCx1Ff3WJapl1QqmJv
+YczZ2iQIsB+A7qT8RA7pUf5Ha27peq+c78ZbKsEt/iHospT+a/kToP7D0mGSrUarcKVUmpANpOS
AlyZrBYJhdAo4yY1eBhqs2XupI5sqo7hTzbEY+X5eA7grWCTze8o7ZfhKctcZ76Pxtzqv1JYsdrF
kWCAeeqraZ9ujrqYbJTUQMkRK8X59GfhZuJaKH8fELYF24CN0jAtD+Deh8rmPp3JGDCfytJDXMde
G6r1GAvRudGjFOTWgKBZAo7s2/9bpWgJcf7FL3tgbReEkC4j0hGrite/2TFEqjCkMd06TcY9oGIK
+Xp4ixgyXsRejKNNL7qP507qyHqUz5xqvKPEorHwtDe92bHFN6LjxuXihAyOYpIJ62ggjh2qLVIv
qMu3IRyZrkRaODNj5rDqp10u+amEP1CQuFbj/1c4qQE4PQ1F3RMjsM4XgyJV7BI60IzA6MDj8tNA
hR7hpTHKFTiddeSuUuyzTh2larJcXojSXI4wanRWVyBKOt2/B4Z8UoSZntxGhMj4qYVpvoZiNwdT
mFT5v0bAJMT8o7+FvdzjfnovrOqPSa4Amt6m551wtM3kQ3h+r+uj+1I57+bfoqPKgWPVPAbmn5f4
z5akcuRAQhc229iyMjMHPNsZ+RvLQlb5piTv+KR7cOYKHcWXV8ozkuyTzpsDXuve9s8zxyN9uN3K
hCdVQ5FEbWpwUNah19Lpu8Vvcw7suiR1FkXUR3NLZB9lND78TR1QPx2Nl6T+fDxB6lXuCgA+bHaW
tvF4zny1l1E0TRNz9v9ZriBVxIvCaUXh1z2Z9yb75Dq8KSvwAfcLQgzzdxK4FasytR9ehKg3X2/W
IVt0xq+tnjK7iYxW8ZrBHE728JMDf8BulSCK8RW2RR4okAXnA+VDw3lqPcltEjFxiYCbUL0+HsUT
SnCwCvxzwwdiNuJtTx/gra8ZH/ijyRtraxIdlN6A3PsIDQhXs/mvsY6oOqseJSvSKFbVSeLpGtRY
j81Q24cBM2LIHyf8GvWrEJgevVvn20pIYe6KjaDjHkf86p227CEnav31UYngbag9wnFFaQDIbuYH
eYNIddoecP0TSIiJyla3KXttUzvn7cj5dN2D64MndjEIwOg+PVp6zKW6vhddyfPH1G2HNYL/T86T
TXfeC9oySZlnnTojiByKNsrin0GiPsbDkKIqgocR52rSgddon7UV5QNuv/speDnvnQ0wS2M2JGfL
uTooXoSWnjRb80EJtF/2NPBUHCyCrbsRpANSQXWtLtzlE6+99PUdVq6V3EjW47jsiCGtTVrk2mBp
jwQ8DQdHLytSXoyJcgrep3/yb817ePblwU/y43N0PMLxEJRvHixfTcXKdbUx02XfpttG1Zit5xKq
Ro5MhSkytNyx+PThSA6gf29t9VvxfJE1N3BxHGE4QNaLvYQcdN7XvCGTzrS+PrL/umzrj4zafvfd
7dvhShK0i1zl3Ey96cQTB5PzFrHBxZRt3ar/TR2nquLl9kxWNT2a7JJZjHBreAi5fFVa4RCM7Mya
g11AvpGKCgOr6glyNnKIZ1TCuZSNS8Td5j7uB1jNBL/KZj2QhhuY9S2AI3fb8TVsqpWQNw+pXSKZ
euuDoaUAbUF03HOcoYvqBSQTwyk49zxbZSPLB0CzNAnHuj6EPgtKyWHrydI7fqOmIRSaY5MdXiDF
p804aJFri3WImdxWU4yq8JTvPw0ulfZfK3z05TMd60V7sSBPBjcz0b/Y9Ay/5F9bAqR0zjHPeQjA
nKXP6C30p68cTTYFlyxKOvqT8KNkKZo3hDXKOYC4A/tb3bjqzilhdjEzZ/OI1iHvlQCeRasGZQ+2
Rfbx2Obf/aWfwTp4edhnxrCQNObFJp9LCeuN2nRkRUUv7cgATExvs1lT4e0ofXIHeUnGG/qWMHCw
kI2GZ6I4gCUrAxZ/nCJrKnX7CYwinvNA+WQQN5h+4SYcCUGpC5gDSlLKD7gnQtX1N0CP3F28YKhk
3kHE8kMkh5UjoHTqg6DLYpEGF1Ap/o0XBEyKhsqnfxF93HUBacT/fjk/GdJkVFsdbFpibYfE/Le6
01Q/j3Z7MAuyolQoN6kuTe1kudLsqfkYPdavznCqEO2g/mr9ux4Fh5YNBPOQop6UrjnnrORc57Uy
G/wG/cI4GBVqWeu+ulVLefUQxY3Nom+3OZM088gfdNy3hit7uw1r2SXfDVOqc6BrDHz9vBQLdSZI
jGl0L12UF8MMNO6W12HC7vYcLy4Oe3AeGv/K1/uxDPR6kUmiWeATSjhF/95ndbkETlBw4AOTXpL2
H1K3YXKcBFfaEyI0wu80TjdEh0kPmzP5OkOblBWzJO0VBcp/ijePRykNjOY3L1AYJzfSqG88B03A
SeQScXfGdekmFS29o4V7iAgYeBZmv1r4UAcNB2a2xLfbK8P7ueB3Ayvub21o6QTairmhgVobFtGU
/y1WTNY587gO1sS7Ah6R4hC7J7GO6MGnhPU8gDAawxdGCQBZz5xROKAfxLjzcVw+zhtUJQPwa7Bs
Sh/3bDGhvwaZXVhXlmY3quUeJXCktgUGos7o7sO8PMMO49x18JeS9xRnahnp3h2zbVki5gHOJcZ1
nxZ9KfmFDQq8v96UiXax3UzCXqgSCR0b3wyfYjtJUasAnwgLlhAPkq+viniqb5NJL/mFHlvS/9sF
lH56qazKZG1ADLRrMhp6dBCd64NWRqeRFKr2Z6QKzydBJOBQaBSuAuEH3c4iftW/UKOqYfNTK/7F
No8iNt9Q8CtDTGImI2Yup10kI4UIcNb04ptoG7dOhOtAR70fdHfSavev3ZT54XExwFvmnCYrfZYf
4gKG04UmZlPYiUXDSDLjO09Y7uLhFfVuglzc4zT/M0rHUOxO3OLh33hn1VnD0cxwmtSkqiEhlAtO
MarSur5mKN4hfj7SsiLUtYEWJHRfQI6cWvr3YsWsm4cO8DUct32Jke5czbV7NKGgK4oJ61e+zIuA
cAw51RQMk5DB1CG+MW3NpY1elNfVs7Ih8sUZ7Hp2yMGVYQGOogpY1XL94rYEJTSCJoT317MgiHuf
66lhcexlp/KmrjdreOob10ihbcjealrow6vMN14VU34eAxE0aTri+YdgcDna0s37WaZH6hPXWHGZ
JdK7Mlp827Pzzq5l57vWBFPC3L6XEHCqNxdrzsjJUpBmaBAWA/L4+1u8uWp85Nmrei9n7qiCdZBs
1X2OQypo+/AvirS8Pt9bK5dFIm8xIT7v5olIM8HB4c3XW8zOh1KVfwsokSoWA3acSdvmucYU2ojp
DlRri2Me3W+EyG5bp4vs9aSkFC45/NgVNjqX2Ep+Jk1KheeQX2vXjRQtYsCkyvspA9xtRGHbh6oD
WwFfn4KKkMBQpOo9k9Zgx6G5OMfud6oIyTZRke1LKRLsgZntxOe1Lj2V9R86ZHPrYvLOIi2k4TlU
x2hs3c/dwJaejifc5NyrZLt1S/fz0ItX4woWMx0ID8a7g1pOiV1zBIRsEX4AAyCvEUnZ6bc/m+SZ
CT2NaexIbgDkNJlsRLnCTeKa25s4l77PocsszXy4kOXqlUwHFeA5jDA4nCQYuVnCtGClwIhd386l
uek5X9Kv3sKbjAakYPmgpSvGwCM8QFa4Fu+aHPLL7mgI4qpuask3RTHUBc0xdnN55oxDlPff6mzU
GcqSx8ns7p/rftqXjj7Br36e3ZglmZtiUvCAJ+UVta/jmyR1OM5faHQzs1fuZcDguyt/9Oi6waFm
p3Ruzttze7XFUopqYpcIFGRduK5mNMEVDURz7nlyGGWsjK4Vq6Gvhy+P+KmlMXmInBwhJLCOQb/2
AufjYZVfyqm7OGsi8mcDMQ9SAODk3yW8jsV/8j13McrYdJDoafYqamTwOn+Hd4fOqELbIWUxSB7P
o5zt4ZQ8uRcu0uOsUDE9P+ssW3R7Mm8+f83migoHNwzGfu5tPALXG0/NWPlzf+HDRnFqeHxY+NSk
/AMPMY6bipd5EcLm7Cn/eX/owQXay60JAa0PjbTtePkbnJ2Owy9/r8u0jnUJu3vBs7ZClCRic/zv
aCFqkEvLeB8RtVRA+M/SyGi4vprdEITg4OabilxLL9UtqpUh4ktJfCuJIt0+o2yF8iKec6ZKvMuZ
QtbGH+ceFpODPqDyHqlNtOeQWouG2GMw+IrxDHtVEswVvUaPWXkLNxVau8CixrFHgREDmEU86b99
3b0D4tuZCuAGRDd/atHipPCCoTS69jllINdiup4JDmTESe72dAKgTPdHFaQ3jcTDNAQHwzJ8Rf0e
/Xync3rQwoKufMJL1VvE4X1xe7AlCNOtJaHkw5E73nSvhQiQoWXNJhBIASApKWGSMoD+nzAyLTXT
Te2xZ/wSLlTOD3Q0P+Nk1jPhcZXnAY16wS5oIP3z5oq2R+JeGIuono+AfxXb8HYtR60WVUtjol/g
KYWzWrfLiQ+offoz/r04suJD66ap1J6orpNtBj/DAxjh2O/7u5dxgG9fveYlz91GWC9ijh3tH6PB
BOPtaacbAlUd3eegAD69Rer5R3puJvXdSxmDW+iMpEqAXBMqkKJipVwm6T0GZGd7O4S9eJmIY82m
JJ0wbo5YO/9JBa+AXQNus/EvyW16StFF0SRanMf6BJCIIHTi8iwGTJHni5T3sUNoOr6BSBEsxJPY
amC3cdpRouwev4u0HcggaT4BbvXi/7arRBmH86bXXTzxl7UFJ1av3EqV6KqM0640sBOlCRAPs1xG
Xr4PtjvvaZYOgyXjohXG1XvfcZ/nzI8rjiRU6/ozf648DnMYdsfu+SG5uPqBdYKRtr5x5fDpT8v7
UHCfKvv45eZVJHOVXG2+6sstu1Kf+K6Mu+lPVM8qrZUGSYdxhFpY4zeak8eibmxkQPqSTJJ9t7lW
ud+lMA+oPi6LCt055ePAo3cvu0dFBWXd0/wabO8D7QXZVRGOssCIKojUSMQFChkkntA9FpTBa9fD
5QmVf8azTglZrseUvxMpepURVEPwWjWnZ5j1OPtNOF4jx+9Q7VOobnP+veq64VBElFbn8CMMZGE3
GH4TAshV4+8N8oCOutn62pNTCZnAaZvhClUEUCAyH8NlrwXxFRd6nIddiKWvbScA9EiJvmEFOIKw
PRgWJngcEFAfM2Jp2qbSWbYOytAff94u44ZPOzJ23qMbX4Avd4fl88QK+6j+iRXXEnqYROd+3KKL
1CpcYQSNxZY1dAA0dWhmOUyNmqUu5lfhXAl/MkHNBdq+nWaWWbsqp3Z1bYoQgHlUyiWrfzIW/uV8
t9VGMZ6Mi+HszzUYh3Qww51MsXaXUhSAKDdEI2kVb+ZAjAEjra4epSkjMFv2TRjZfR2D1mF8xD0X
NKXCa3FWF6HNxWMyhlMLENEicA4kPD90BQioVl+GWSrQoHLn5ySuIn9l/fXDy/GaTz/F9VD9tF0e
7+22QXAbtCHVoHq1njisVRqM2M+4h+PQbEHUssTQVKm021aJ6rGU/dTEtmjpEfNxLs84GEygpaaW
F6tIENk9+KtJPUIGLUD/MDNpLfhoLx02oVQ3AnEnKZyXDsaEkzpBqroel+fbB4WoU1tE6p/V/w/O
BudU/rTLcdsxzJc3TfYszYw5ieqXCzZIx+GZ+lD7puVyZ/La9P7owxRqGjWD0spyxcNLPrh4Zxas
WQNIWIKI7SPmFjHc7VJWyhUykVu5azGvEB0T4aeS9D5+7oEPfOZIoKHS0PMAGELepxkwyqI026Ps
euLZfk80aodRNA5eSGmp0oehX1cCBIXmCThW1pFQ3RJxF/6yUIaqUTonkNe94+e/79j374fBG0KM
DuQya/ScY9FoKzNM+78qLFbHgn2n6C4OJ6yx1ApVE84teSuku09nm8wDhf9e/D0aeZX1bEqbmqGs
Mqo/EBt+eCYP2TlO4KRDIe8pek3UdekleO5IW5an9bxD3GamT/bIIf2zRmqMhzjbrjHahhCeOFzb
zRsN8pBw5qy8G3YzziYKjD03tejnvmQY5nHKQZk/3W9X9RgbR2kbWIJyYrJTVhwUd/GDryD2xuAX
KKyIUIFHoe0bxjONkPaY1wI3MTKNQQsZxnV4z1wgJvtIdZRuVttFjtwZg68KZEK5RC74w9OzYgCX
rXBCgWJD2P7qk+c4NyxrnjG/WFvVeIp0mvzWKNAIJjKJKhHcXrJe47O/YjdCqp18jqGc2Q8oWclu
Hj9/LH8s4RjhyARxym7CTlz+uTc3xukweRYFEiF/6lYsyjo/4q6PfY5ZdMcA5iRT1x+YJBDWyv4U
5i1vWSauARipNroTX2Tu+EGgMS11Mvi1afLBj/VZDD0ao86kT1l+VXC2c/TSB5EgFx2uaf32UUum
02//WxQqZP5fHQmAIRosfFAjoUIskJ+sZyS2030LUpivn204Bw1B/JgbJtlCfpqMO/uHVUCDgOzC
CYEjzIMWxTMmYAYmaZ0+jARIU0byF0SeFOLQJ1e9EJzwyutrzFmPy4OZpddY4eHdECUcn/p9rTVM
SbYO3smi359K6f1IEa9NSqMmBaURZO7rTAKmdcC2rjP1hz+3wMH0DGXk5/VzdfkVtJ4MfxWGgY9S
QlqjpCtX12D/gFprwYLTkiK4zlQUD48wHMnIB+49sTTyPMOZMf8rEkxKb3oxupD5Tn9Fakj0s5re
TyfAp3LYkGe9PyFQXgQFDnO3s0EtZ3nZhi2OFc8Yi0MdAUL9gbfMIFn9NH8+GEl09e809FjXeBHx
in91h4QWsaPmzbN6phKmA0yxcuv9lKKrzGarm7twkIx5bkqJFZd+MfX+F6WEGUXADpUXykEDhwRK
z2bEIx80enGZtfFMKuZyWmbygtz63NyToE1heIHKWVJ0k8YRhFmKjthPv83S+DxdZeQSjsEtI7An
5oBGm1p/Zf4isJeFpa9Ahxy3RpAdAbMj2OTIE6Iv1bWT/J8/EriZDzg1AZv+iOmFfE8yCOoUQR+F
mvC2MxkdWxZ6v6CiARJF3c0CKwO/uX4L5IK7fLMHLg8uu2AbYWUdZGUazsZep4mz51kKBuRqDm50
WRBo+NB3097HU2Zx5dc/cEiF6NHcV1t058fRGbIHyO+3s38vFQGL62RwewRwCiZGDBEubdML8m+E
wwIL6zrsB2xZ5eEGaOdZRpqjmKUakS195rDAgtwcHpjf9RGjc/BpJ43yL5iyu4eEcrwzkFPUT2mJ
rWALz1Y7fXq4PN+EqhzJeWiXmKwjZ+dlRFLysse0IJz+EuKsP276XbFgyMAtUni5YO1G3kcF5BkT
uB4Rcw3n6L6vYzAw3fHLeBOu4+VjSVF0Z/hL4hTCEBtqlyukGE18KBAYu4eLrAue/KTCFuGcN9gK
rcaAAmxtEl3peaI+UqUqEgSSXEvzBh9D8wHK5iFgqAq3FR/BdogHpGkfItR+EpNF8kquT/gfHPLd
FE8100xrpJKtLbP9N68Nh87X9uWBOBMQAwwdz4gEZsaNQ8J7U5mRoqrXp4J0pwKB1By/Qb0Ehs+l
HWPsRVJr/MM/b+T69qQLT/8Up4z64PTXMZ1Oon7hJghBYWbynthkge+RusYokQMRTocyhTlfgrNk
eirGf9sk813/H+b1mGq/Clnw7dpVGAEERdpbQbfW5LXWHLitPfq4IlUWaCDWMw3XGxiR4ufCaRpo
LaeAGn68Tnd1FlWHfkEbS31h97Gwe9r1nunaUxN2YrM3e0RS1kkdd9laYQ2FOrb6CW2rInP7CVkn
l7V6NdcSxqDXODozZigGGdOlcCT+4Dqhl/ywm9R8/wMmPHLliYKxR6aWSmCvqdhf++V3e04RdMN2
0p0P5GLzaM3QutWVmQLPO+UEX2oK9j9G2Y2ll4Z4pVl0WU40xVsDEbv9R3qLlDZNCC4m1Vk2S6x9
XeEAxlsFbMwdsa8kxgxLJTxzEFUTBKdME+VUOk8HPbc2Nt0O9xrYDj/gDHcLx8aEtM0b7AcjVlJA
HmVIl5MUwW3MV0205mzI4DQHEh4Z7MJLu4uoIz+U6WUxbURpywdS8XC65Vt/cvuov4OGONYRiQNa
VEJVZFG0S7cFnEsanEWGzU7W8/rjV/dREyo6kiuR/ib4Ziulx3xM6Nw1XiSFc10hnSDCQ1aEYYiB
d/IrztODFBkgo8Q7VIL4VSV7wzHIpiSZxAmeBAFtI9UE75UWPvPFQlNSOiY8MteW6Ur99NTc284C
DvNepx+0Z/M0ZsaFn4uVRedFV+sl1I71ygaZZIcdu3ATVoTTd4nv3d1H/EoeXfczllj6NQ7uBEXC
VjGEAOgeNd0cdMwPoJcvY250cDYKh2F/QbhH4CHKcC6gMmvJF6R44eMoZgTSBotak1Dp7czJwntd
tYoDPzzdSnQ+YH0CJsQPd60+J7Kn/CQrE+D9DBXkyo7joGiLNNQNXP9NxMa/+Dtbs5OslfRyfNxz
ahrROVqSioCbgSBqnSOzBNje3rtn+alK5JrQ9YMMIovwy0j6jaoGdafyYzaDv2pY9dmdPVILb6Uo
8JX9DUwBD0pfUXcRISgR0X+I+MTWL+9zGb/OQ5NfNQaCjM7wtThzoljJ56zl0EFaAf0ifj+ucPff
NrsvlmezUq9roON1CMSPk9mB2J33DxIhpLFqTu1gUVf9f5xgwkw6JY2CrAQvi0WvHrSyNnWZIN3Y
3j4nx5Sp9NseV3kUAcZahmZGkmgipPS9kuWMmIovSGUiPBA63bngfoFX1FSPF1nFRmt88KN6e0BU
CnCFYay7qyXgyugWMaV/UG4xqudHxRW35kjMlk9Xqk28nc+3wB7d/MbcdPTh/nN42FNYWpE3bMw3
iFflTwiQu0cHQQ2h/7N+Eyrst8VibumWrDTaOPxSNlpxCDRwfoo4gZ3Q70WEuU2gAyF1phm1dAqO
kLNmng0dRu/Sz+I3hBo8gWaeFwo+k9G6B3yjrNKoZWx3Mjgm1+VyDcSm2YFxF1ZHNfAYMUtQOl+P
kX5YTfCn/X/n1f4YpTdp9Sq055hi9JvjBs/Ws6scdWJxrCpX5xNBaKiYJuATNlLcZnzloP1uAe6/
b7Cc6CozGbNp8vstgL3Jm6T2ggdSfeLKvOy6GpW3VDuwUPUFCBaM6NIVLFbCLdBShk0Uu8mA/Ux/
arTKWqecBiSmM8K7k5CCG1eS15fJj2r+o8/MvTLUsF058Xzj0+HwEqS82e4aBJ59PnDK3FRsZj+Y
Ik92ek8MrX4T9P0i6VmJJ+SxoCn0e/zBySK0kepej/jxD4Kgq8opKAt0IilFPAWaIElyt/gyWkTk
gWfCmtQ9D4DM5SIx1BRMC/qgcI4I+k96CbN5bgETlEeYA3rCA1dLNjPeV5NK6Om0yDRAd/BxbkhU
HxPojX+z9Mu18uzBE0MfNM4qFGgyVEJ62ego7i0vsSh47En9wHR2r7NlPh1UoaUwlleps1hHNxEK
E5nZNgzqbapXAZ2u1Zq8L0Yn70MtjZGVFr2ccXE9Uc78Z86jAe/UNWh4TPVxAkKoxbxMF1ayFQ4J
A++/dxBSZtf0SuNNusbRSYbuzQWsT5znFR/JQS7GLSfpxqRffe22ptwGm09MHsc7wFJfvHd6tD1b
SqB3m854OdXy9M4UdQ2vYdxVeATS4Eg/SKDSS9OiuYKHMp0QDDou+1j+nl2vf2Ej5Jbe/no5Ku3F
So60IkRy+WWATwuY0zdCI1kz9kSgSjPtg/qXhFtTzAic50XRpB9GjruIZihvWV1R/Mki+rrUaHVY
MR7SyPLmnhO3yERfWLGnUqrWGf6rDiGNlKJViUsTpCPiVQIaTXiIRzNodxb7CKikbyoclQUNSd76
C1lepodEKcI49MA7sVX9FqbIFO9cJyZRCI8GyGjWHyFGvJkL5A2X/GlbKyB7ZDU306QsZaZEt+gt
wYYYvOmQbjBL4ajeWCy+XOW/eF7cNpjgQnwNgR0SdfxO6GA8yQSkZfJUBT+DqSomTQGHTn0WD2OX
G+P1JL2htXc7fpWreT01IbDpMd/Q4XYyy32zmBCWzkJxs608pkcN3rarTouf2xQ6kh3LdfSg+Ll1
MFFCZyrP3N/vMfT/oJwLLUHz5SrUKH2EPh5/k3r/ItSHz6ms3tTxxL1koJPEFR4jYZk46WNg3Nvz
Da/9q40tmFISAozOWSy6Aoaq6/QGZoeABxpdPNozTw8CisPnnmWBrdl1T1OBfoJtZx5b2ae38O4p
QWkB0fUuqO7e+Zy0alkzmqAPb9x1ezMFCHBo39WQwe8Ac6Ko2dT0tTQ+bEXTgJbad5a7Vj+cRpGE
3tR3BDyNUjrvtoFPU7dIV8bnezSx94GyABJ46i++9emcIgcUDI/TYzoOsNnIVbiq83XpclPp80Ng
zX9rEy6kenLfaldSJTAv5lxZ5FIKbMbAl8+qdA0yzjd2leKgKNkIo5qi1mMLGnhujG9UJs00y5D4
OBd31HtgO738YX9JVaGMduxrWUMYTLZRJ0Cilie+d/3BDl//Zj6TY1r2TyOuha15ZlyVS8C8ai/8
DL4F8ugXCKkpfYIRb1rd6JfNoWU5DSKeMvvvd7xU9YMAGtY/xvJwjMLGXZAs74A6zh+4swdfCABK
35fJZ6jhFy1n+xFIWr1o/KjfFjOP/NM0xLD9Q+xuKCDcnTWfSPjj7CbxlhH9xuvKQDZ37Dj+uBca
hkHqHtRf1eigQTAoO5zMZylOureYsIdtbsHXgo/E1AudtU3EZ+T2uG5acy8FlLTaexi4qk5Ex83V
06XOdiXeqHmPF3et4zRefN/MSwvU1f799eNDK9rbF996Mq4DirrCxQgllU+uCPUrz8UXE0LxcamT
fbEjmAXcTq9fL0M8WywJZ3/htovZBe4eMF+RnkfaAesXAddWSN/jPx5qVP6hXByyzhmPszAlqWsZ
Sk+OVUZF1eS4Za9IrWSygh69tVnHlnSX+vEQzccQ+bjIHjt63j0xP9Guh76NYnfubcon1qkdQ979
iMcbHqX5dsrb6wemBx5nNvTSSAm2TN2kUY1HCRnovve5q0jgJIBWFQF6xjFxPIOtmMSMUOOtejeA
k8e7dO4aV1fWnA6o/Jicy7fToz19MvjaYWh4XPahTd8iBHg6EOUuwNtrJ0aDyF89qiQdlVPW4+ps
XJ5Ok5lfKhUjW2NB6LNvqUxqzMMH/Q0nVs13iiY8Er5rPgo3xWunCNYS3sGOWQf8dKXj4zkoDMyk
3Lz9OguC2NzDQ1AL76UkWNSiWcHxuJfWeP2bg9Fa/9XB3wyvVJ/S0mzAdPXIC2sanitRXToKaDQE
BvYluh4UcQUDmCj44lfIz/zt3etNTx7ohh+Xph1A8VMSGXDcFOcgUTgQsk/X/2HoJe6vYnCWWfjz
hrHyqGBwPfrxupItDyIdEGJ0LIv3ElNjmlUW9mKvuRdi9XSM4o5H+Wrb/9h8NwafGYK2QgEMYenm
MBv98w4bru15u3jmJIte13lYXnYWBQI6vZDzgKeHWvmG0CwIc9RxCEJae6mjSvK+2mFgVCNB4Zyk
mEYrH91Kc+3opNrRG8OOJ/Ks3ic5V4DN2xGycBB/zZ9CsOobGfB1Yt1Szmwv3nKDFZd1EmbpNxuh
nSyuoPSS5sZLNKYwO2c90ljX9Y0Nz2LHSqmlV+fJz1hGWkH6t7h9ciVc/326vvb3FFQOGEKVlhlC
CtRXPCW20ud9uU+1z8EI+O6KotMeboXMLfX+S4xuYxYHAurBvB52LCLPc/fo+3HJNPaFdAoBvRC5
LIMobSrjohyNxzeaBJGEfcpTXQA/elGTa591HcPaWWCFhwkxxQxr2ZP/i9nTHaqDYxTSpUncT5bZ
Mj647eM7bGuh8OZAhYQGZBgPV8EF6r8umCBA5R8N+OTJUw9VasrKrdU/idTAEHEK09L2reF7fmbd
z8uKB4/wM5P2ZBnQeJAl1XCJJlVpfVMJOcf0DygjauKNjfKN5akOr4qBjW+PeAeA7QnNh3TOFeSY
GGnap6FL0TwFCXIzCSVmoUQz4CGOss04gUNKvb36YO5wK3GMay8lCWvQ3pxC2kS5pzN3oWjDNYwL
Tf8FaLSY79T8sOEGMsy3UEW6OKYkxzl0N5u8j3YuExQZgTI4plK3hDopfH3fR8jBRPLM1LBJ4WYs
kP71xFeAWEkIlMAET856w7NS52wt8WNCNUoYZ5rE0DRSgEdU9eFk1Uk0CUaBDvg0UUHE3OMbvlPx
Q3Hzg4N6JDujEx87gfPhfWHaFtXVTAzw/v4T8bdzQr34znKA6oZHRem3tO9SiqBoX4ocq5msrlE7
bRW1HlayF0tW894KzhYzgzLCftcYDXw1YZjIYFnaXKIGFlDlgoG51L+q5OAa9WWVYd00/Ik4NCs/
tT1GFJKWIGblWSWVoTFWkhPTywR/2JocSMqhWphfiRkT9xFBtBbka9efBGc/UD19kxgb3Dr+A5HV
82i3jBf/zOhD7BQbYIA/btCukPPahoI40GNFdE69X50R96i/p1BtblF6zbm9CbiEg3rPrczrvHz3
53CtZxJ3naanOwmcdkfYNpW7lYTn2dd247IIkexi/yzwYKiA0USPbtQ1nD99AtbEmNat1cL4jPo3
QYRTSrD3WufF5+KnQrpvKR5tKL/QDL7tFR2ItxRtpvMdj+tffK+OxED1IrOAPyTyLG+/pzdWkWDE
eLQg2rMNrN/251Lriz2etVcBfl0c14jFzBD627lNpCGzjgIrewrDHupDzl2uPgZ8RL+ZrtH5v+P0
vDRo7qYMHxqBeTRnJhXmwdD5naZK05qSMwT5sAuL7lBrq8zcJRuqg0ZJvFKd8SrCgPkCEtnzPF6H
wbLow3RaiahGfHi3xE15MMbUmV5LoXQJqC4rH6NCFK59ZWWl9j999jEFU7OBI2GXPRZrsg/glk3D
cm90P9sRxBtYfGhk5GOqtKOEodZAPbrWT+5OenUeJgrE5yUiG9ToW117VTnxYvfy79pHMBe7m4gq
xsaQ/7KPO8VswJxbON3zg1KAWmkBqlvBq7A9s07ESxUDfqdsNXLuu0IjyK/uM7v0NVqa4MDAc21X
Inu4JPj15eang+/fJfrWprPtggcughHDSlrZ4guv7X2ZZx8yjcegzZyrCqkCD95yKPo1vsb/TWdo
3W2brDskBdh6LhflzAi21vElcCwJriGw8g5JLmLkzh6mgBHeapY/0q3ur2dmLX3evMjX5keYEdZO
/Ag0M1afHu+ZzWTLTo06uS27geLc5lGzVlW3ydxQwRN+AnTy9Zvtw3Ff1+Js89Zyw6W+xeZVZlGp
6t1hvv4nwB4PSwN42+taXr83rGfsqjzHN3UOjhsZu6a3f4JgHtXHmTwnmcysM7jJrc4BzsBGNhyg
in2Mut6Cyq/ZHlBLTm642RWVoaO7FIegS6UVXNJrflXIVrxqiyootxqqwvYfiRWOysHgtkdEfRJH
UronN1Z68pENmuh0kR1z07AyJpRya62gErb7B1dOPCKYzHtOWD3WnghA2/PTwHbkcRTlrLiVyGXE
usivoeM9KYAjxYo7h7nCrBswTLik9DKpShAiaEM+/eilnVr9vQr4sGZSr0nKUCfBS9WrC1S6e8YM
jw2coM6sdIvOJaMr5ILPNJVIaZlXFiRoIQlR81Palxc550f7KMiFhZ3bwp8cINduYm39OczRG5GD
a6ATUJ+vrGChZI4nABbyUrTIZq8q9JRuaL/nBVKsxs9QllqmmujgqE8hXdZZo7jIFN0MVsDiH1Li
8cgLw89Yq4o9oCzsgTxTE9YO2No0x4jy6C8OxmbrIBfKZvO+gB9MpAP+6hrG3VLQn6AxKWvD7CLI
IQmGuhtQ2/wo4m3ipPa59iyO64H0cNslS+Nc+pMML7/pzPyLPQRPrHwQKr1u/c9twAumhSBN3mQJ
mbpT65UQwctdvCVPRu58U64vOpk/xTYyP6V6bFX+VALwaOjamLFVFJO1kkR6ux/8Fs+1W3ys8xfv
rKk0lolj7lwSy7yMcDXXwOJtRZJIyeGs8GC90Xoj+wPOlSuhvkIpP0EdVGSCOuGohPtKUbzh9puR
t+r/DPquUL0G13OdmzY0Bq20+oOJRuAc2JTf35fXoVcm/7Lxpp+GN2szy3oLMFmB5bwbaaAC5MjW
w7DBItglousR+le6cBPcx3+jbwrgHytfTmlR4vxQKpDqXxUTTUvOI8Y3RHa5rMEDI3R2+dIYg6bm
tTD4FCNoIZuyKSwN6W1fbeIjFylY82CJKjNni9ZWjSRDyFwUlZw+ID2yTXu3/M2g0AJ3olHz6YDo
T1ilIPkaoTaoZDNNoYXiO4ImY369LqPFAclldlkxNbucwtKkVyh4KyTbhar7P/L4pXTbjMHxKOIa
eUk2CRXZEJ3NM2Ruk4GOlEkFyOeAh44SDSb3QhV7yDspgYFlSJ9IfU1ZRfhBzlMEua+kFys+toeE
BNgA3suYo+KwAVBLM6dsyI56/xeC2hRS9ddzzx6jzrcx/LSHMa8r66/YRYJXpan2ZSvQCgYmgejG
yHvT6ehArIQ3IUtqQyE8/fk+odZqbdvQhgHJVOaZGb7/MHzEctOChAT1p4o/6z7hVNR6XbWjk5bt
IL3U0/WFo6IoG2v/picau9z6EO3MRMGHGxHtlsc3JzZSjODJs3h2GElFFgJxrrAGfjZBzWNOjji7
vf0g1HwGy9ZHMD7XabA8OwPlvFd344c9Yq1DRS31vo7dobTVjQSajVqB1OPbat3aTDZTBlczFJ1v
ki68TQ0DCROoGzBbRMdDHYV8ZB/4+0/tw+FJBqDXGjC93Kpjecqt+p2nmv3WLk1iRUwpTVskP3FU
ZQP5rX1I8Kvx/9YrUhJ/1Vyf36SpCYc4HkdR4HlO5mw9y9J2rNOC6hIomeRIEfVlJzeNL7uKBfDX
7U3NkDC/o15Cx4CpRgphfRFfMwTI0m8B6BWyIHWoVSRIaOtGG7CCq5HtkucUgp7UEg9I7hIvS6ko
vAVSbGuP3ipiqIwx2MVBsF2LhEEmAekIsVOV0ezk6Fz/eq7xTFbT9Jfed3VfNqrf7QaploeEEx2l
uuDJTTkE6W9/2X3/s3J46IMr/mrIRYrJiTOj9d+X3Mtf0LHiCXsSzIevLuWDvY12v0RKYV+RpPQb
X0Xgs3keO38laCqjHqcBSQwIpHQsvALCZmfgUPU+K5V40pi5ByHeXgOgpCCg3QNLN1mybmb4KHPf
6ABcsWkXA2+kRTfNaOQWNpsrgeL0geI3wy9w89bjXTQP2ss8X+DqFbV+QoB0y+iS45e8w5TkcbFR
Uo2B//g7rzp7iXcjIQWCVJNqrC6ScC48qDRweWw6FzZbl9bjcC9TwVuu5KYtw0WWZQ48Fv2MXr8C
4jonSNso6iFtTQVEhgpHryTmmuyHAFQHyMQgI/MBJpalhC4b0oQ+WzsM0WwCuEqh7N3BAgaFJ8+Z
37GhFEEA/bFkwF/xum4rBWjhoz2kYPQFKTnfFkcHzy3fwZPmBWc5BtxEyLmFQ14he1VDbYM+qnZ6
ye+9FulgFybkZKA36KgcCPw+f59zSt74yBgZeD3z2Sj5OAocHOacYqN9QN2ltpX+WEhWyGvJSXw5
xjYDqDkIACEcmTIxyxcNtqYJ6Vt+auSU+clB8Svd+GCJSjcG1bZZ6hgrFc56lJMxVGvy8NY58wiM
bp1iGyh+cXiR+YhbjaEKKk6Qx5pCyfgb7tNBktofs5x8GO9kgnsKJBCA0j55uuGItCdgYYmlrwbt
EWzqOHWg1PzmPkkkNoGHL0Io/bMRxsQGg/gSvmegVRbf2HtlCGGqI9DMKwGg0GXYNyiQ+34reR+r
LUf9G1rLyDAtKqQVwepuiME5iAqu/nUaMPjAcQe6UgrqiUW2Ieci4GMtltCg5+z2GxvwnteSK5DJ
AbZpCXoMKLU1rGUeYZ4O6RiYj2xQ5f6A/i0f9zWDB+JArBFJcmdFQ3mFY38aNm48o67lYxVBtsuA
7MaoudL0hBiGV8DvGko57f/1qIHjbaPUHXW4DBRTU2ZLHoj2l2mlMPSd08ZAaMr+P0q1JUl8io6j
lo8JXbHbewbwOuh0AxynVXnh9LFa2cPNlw8vFwYdGkGn2+8YqfrU0NjCQn00DCUvqsKzeDLGdM7j
SJD08/nm6xa/Awob2Uyt/35kpnMtdsLsh/lomJr+VKIwaAbhWS2UlrTQPq/aiSfOlLxNixNGOZLM
mPnVGtX0/EhsNbkdHoo9E+kT780RHJB70z7CPevy8vm3NbTO7WJCjsA3MLnQCDTgmHpBE1c30bsw
Vt8qQdFU4EeAJtlFtJLcHKL2zIMKjJ4jDafQ3lgoqdltTqxkkVgMJEwxqljSZUdwYtfnafWDR3We
7qLe5eFe0o+dCg2eWbPKK9m3yhV+Uhj6v0iPbxQlU4iiEJk4YRAJ+CZnI9tWFpLysI06H+ZPMgkv
ck0k+/styrjMw2sbwLB/5EcLU+qP2qO7zTcamNto/Tyz3+nycETtabTGVsR/bS24otbBThu8afaV
QxPFGdiqywz28AnMFyu8z2sz/+W3vPW5a1obQOxWhuWu2A1tTjZR9E0SZNAveAI9hBaBwTj+TGRf
2hZy9kZishZA10Co7bl83TnvH99Do/bT92zGHTgh2zl9546LVrMxEOcLXMA1c4lJ6TLsF+nfpT5q
g2LqhH8/90jQ4jZYnICQzNHPwuNSJmMMXSMT+p8OCfLj6istk+fmrjgNNVE4Qwt/5qk5TP9ih4Xx
vQZjyoc02xHauFOVRDURhzBMbDd0apyoZeiJHDNvy/jcz/Mu/DM1xNKyeSnLCcaa1LKYnxeuSeaY
OpBmDMTnpvKnNJc2u+Xzp1PJ+EoYTapcki+8gGmbo4EiYlt705x1DMgqwq69T/QTfOX8q6hn1mLK
kJSY1N02z56a9zKX+T3GSNQOTs6sHqZMuwos32eUhKR2Erm+Ir+1sTpsQ0ZEcQ3x4AlPu03bSXXP
reO2HdE+QGZEWdKcPwgUfx7ZqYUicib4iNfD9R/+Q/vY1Pd7lFM6WJZ7rVBAq+IysKgeM7pNzu+y
HAMrIaK0qUQdUspOSIS1HCsiLaJQeiVWSOy5Qk2wZk8jf+1gef65OOPIDsY86fXjBnE2cubEs/rB
fk7XSbEPX0UrK6AKVU2VbFUKMutuPR5+3r6tf0jb4Mo0M/PdLDr6nLOts1e2jmrvZ+9zcCizdNTb
RF5V9hh1Bz+Rpd7yNT9DXs4MGcRjHzuSLl5MsyB09rRYg9Aeirc1Yr48kU1BgbfWHbhNOr01rJmN
Sk1PPbKYfDH77w1Bjv7YAFDmBuNry1mtygWdnP/OKQNjIJ0ZBS5g2oLzdf+BowgHX2yOAOf4+8jQ
8CpvaxG3LxTONAmMHR9YKKxGIegmxZ2l9I4tvLJQ3Inkf7haKHVFwt+jlKesyEDvFyAevWUiLoDM
H9Bss95NTVMER2cULJVYMQjH2+byoMaAfg1KIEQLPpOFyJW13HyPlQkYB+2CnIzCm/kaTrXIRz3B
MPnVjMBrYG4f/r1SldQs4L6ifxrFeT7vf9sdOZ5ASZ650kzD7aRyyniNWIYsNePLJMoJGJ/Ru4Vr
KtHZziFJ4hs9AzE7O1hG8v94h4R7BoZG6wPtlRlT26GHhwV02A1InG3O79dyZjqY1SChUQoTZHqH
wiqCoS9jkAVG5xbGB2soHBDLq5ZAKVjxmS3FmVrYAGVlXYCbFruqR/DhBWEcoPP9nPM/6b/bZrtV
DEBQFZ01sYNBmjyK3WpGqDOJVgCahocvTUs+Fw7ia3svsDCKYRGy62Gk+yE1CFT/3AwAzSSj+8on
uattGqu0i6Ii3UBZBAuPGLvhyAxf9ZPdvvwhsNRs2lDXQZDZwTHHwXYKhIcfcNa8V+QV1Te5/zD0
2Pxnbw6DBZ4MD7pws/q6oj7Kfdd+jdOt4ILf/+AqRSHGRTTYA/V3S4a79523INcVBU1fb0THWNvb
0XC4ciucugE3tMrSFJhv4MztTOBpW3PLgaZWeDDNjEiE15GVA81NUHydpsnEUiN7O4huUv9vJh7n
Xroa4/et1lzGnvmsIJ+CoH3QvoqPGAKnY359+2jdPV9X2G/UWpHZIc3ntrxFomFreNcPUG8E98YU
mJEFTMSkDvi5rRz6b7Eph0qo84cspC4mutcV7h5Ram+JSMHtJ7QZs/xPcXKdzQTOKaWPRz3j1d70
k6yaSrOsnnctF0w2kZQGzHFoqCV0QwtlXSjCTTCgMRuRLAcIqp/deEqAp3m+kDBUYo7slx7bYeH+
1utEarHMBs54qqvUuVSv3vTmdXgRD01eApSeq2U1N9YjFHASTllLYpAh2qqWKTbRRTwzRWb1AibJ
bhVlCqnECbRrxGv6GLjSaEr+y2wqfC4HGoznOXkcyIfcOdewUeTyYBFffU4FDGAkzuL32jWGphA+
9tVAuouszldv7k3p0YQZU1Qva9O/g8zeCL2sRVOXNUWgQvxU7MIs22bF6jwgXr80nZc95ol2JKwU
eQoOWzSmRVcTOFGt5K8JTPNbq7P4+kSRu2UtnWnqewNhS6dDIupE1zCya1ofA6Ifilo3115huroR
8eppkcWvr7spZYSFF7BSdZ9Z2w+irDW5PN8jSCZRzykbdRKJCgysz5j4Pznf3qhT0xnVs93bueND
f0UWDEuuZmz3zEq1GfUtWLWmXxrGhzMUJJQwCPiEEABMffEb7bZ0qG0XIVezXrMGG0XL3T1Nu3id
ENmUYkW+9elQERf7Eqec7Y/1HqKIpuSPTbNyZe8NuyxKUmeSYOhr8Bef+GwhB1w/Hxsghwn4/4In
afVqpcTN4a797D1U6ezi/X2VN5SpK4JrRL2aRmWVoDosWHoPEw18kwAyYyXxwC/QogSYQF8r87c4
zraIlXcbzZHkBNEkgPZgvYqMf2A+bGrSVT+9PFeoxW/kMYwmNKvR4SSdGGPCOcurF3Lyk4aaPnKu
bR/JgGeXlkPE+hFKGZIMhMbLoKrJe1wSmY9QU3AVvucT78TKvPg5Z5hxy2ZQMVTiL9x8Lx3ekZDt
bFMAcQoJ9QyR8tKCiWjXyzGqWlGdILW6SuebKzGfPn2Tu1U83PmDF33/ezveNysrO2kRpgHxsAQE
TO9mJYy33GCCivML8YFwb1omdE0HHMfIzNhcKpBV7+DxGFaBmLxkusCOVdIIfolb8Qn5zW4cIh0B
tRbdvZfnzJRmpceQ0M0YK9FcA06cGx+6+SeSy0wVc66qEJbfWJ5q6cVqN7W78Goa6d05jxLltuJF
5qgCXPa7fZMdI1FykWOM9nLVg6Pw6BtzzxlHSnJRQXeYhMckaqmLi1MGLn70NSBQSkvfRS6Bx41B
hktpdMbMpU8LBgm5N2opVevDLw+zjY+JtjuPoo5jAhLmg/brK4gb0IAnvj4xdGGIrJ9qYwDOwW16
25srQf+f55fMv9gFAZyRTM1M9zwlhmMgX2dlU224Pkj01dI/47hNIKde+DIUmq3a4f/ktkej166t
NLmx6CM2kbtp+unWKEmB3fcTYP0pcu2Lr18f7mv4Pp6i37S6pE+IgoAM5Uww02oMGW89FQcfu7VT
GWgbtZOTLvnHVG2jo/ZmNVp+U5dnnRH/8qUzMHazLEn414Et9ncYMJ3345Ab9WsQ3kYZ2X2zGrkT
1UJxY4zY+CULstJziYrrbjd4nKevU24qz1XFgHf/9vzMllENFAydpgyv21cPa/M6AXxBHd/Ri85U
GvHigE2uOH66R46zDVnt53TDpc3GYd1TykrjaKCFG4uq6wbp4tCFAjy6F/5HkTuYHyYw/rYG97KZ
dZuNaLVxQhuM4qh2CwGASaHPEqLYR2I//1AsWnynkZaXx/qembm1borcG7kXpj9umjugxlnSjsFj
KkJqctyt91e6qb71t7wo4F9HfcmXxl+A5IhDrXVIBkh/9nc2RQ4cfiiKKOD5S6zLIOPdMfuMBN5a
jr48CkVl8e4Q1jDxtVbGgU21hOkD3peEuc03QQ9qPniCcxravKDwUp3QaJxuus+qGqa/Y98bFKaa
N5wsGUgsy30S3EurnzRZRf4Hd1wgMbqDh/bCPBWAXJOgXoV6YB3bwHnlPJf7Be03tvq2WfoMW7+P
gGzyEwF+CvXs9KVPP1sWTz8lVpj3nmMIY5yerpbRdYpyC9lNGSDtHiAn3x8LaYMXD3EbangRPmvg
MR+YBAJj1eE+nN6F9eW9sRjMSRCtOAbifLznYpT3YkgADqL2+hvk+E23OCJBd9J6tAgQnYUXkxw2
PcbacMbtn/MC32vpMwvAmqMlbtQvURwXAA4+Vucr5yRPsLH3NMpg2VPxWniZSW036MVloNsQyqvB
d+RcAI2JuN2tl++vAy7dUvDEjjg2KX9hAP5cD90R1gmahaMA8LLsPUA4pmxci1/izczgEtqae+Ro
Ue9F9JjYD4xM2YZo4c+rU9TW8WhM1+DHphRvJLk1h690veEaekZD3rPbqVW2bXxlhetY87Wy81gM
OPnU4AyHC7y5JiS629+EHWM4l8LRi6qtyuBskwXJfSg5/U3ktsiPmEEVemrxeCYwh7yS1L4vPDMa
PvM22dwnK8rY4QBdFfdKV5qBt2gEqnCykgAD1cKWu2iMaWYH7BqM586/8QKcSj9kl9kp8tB+1dqM
j/Z9HVe/HNV9r2dlTJm5QLx1fUZIc9jZQBUKJWcXpqYBXZdXSSsp8CjwnHHbIy8HaSKMNaPtOOYQ
2fZ1kWBpErMvWlk5+1aoszE2FivRRQP1vfAudpO47pbZEUnPoSIrXZgPTaq9n13E1dFZL43jxBh6
N9nLxDPHMZE7Dmu5WDrOx4/09eZFdlOI0C8nC+n0LcsdAZj3KqsvqPzwl6g1Zw+N2BBP0orRduoD
iGoZ9mnJ4puA9ISgXIWBVpYuIC5wUX0aLwsYMN47eDrdP2wdMRiEJie0vzYktRulcUvl3yDzYi8E
Qbm0EQT3zwrHd7leCyy8hlhZabKsPzDzEVe9BQGBsi0mZSQI+UwC6VZbQLfkrZiCPTtillzME3FD
4EVRqxQv1E1Hx+4e4Zqm6dGNO1SoLaH5sBaJ3Tf+QOGE5PzZ3VRxvRrdiIsZ0JtEmPUNFezrPMZ/
j5HdaqCoGTpOub3gihId0/HKcZWHXcLVMpcVEdZ0y648Y8ukWtF4Qw6Rw3YlTeb5x1QGV1EXgubo
Gzk2NnAjmOcM99sruwfsekwJfp5pGK2kXK4d/sGQy2DhuPjmyJhPurgeUuz51/SSzFSlNoaeBG28
QiX1rhqiZRrcJJH5RLh3mcNrV0jmWlKldnRcfs1Xkp/+Mdn+ZORNs1rHCWlURJSLGzM9PxYzb74H
RivLmn54R0ex/X+wpZRziBv7vgOmXFlOQwNpos/vBlfFJWCaPDWGNnqm4jZY/Gri92Uglk/LrGRK
oVo8WujbUamGHJgwGY2q5IBAuGHj7SpIt9t7XHWzaUtxpqdN9WaVBHUT2f5ysOfmi5fiCWa5BKHQ
Q96Bygr7Z+dDYj+3k0TT2RLlUZ5giRE/EinBIjl9cg8zicFBu/5R9EXqe1fnJeBNb74RwdSxT9Pp
YCn91gf9YGZlYidiRLpfYXm2ydLGdDp/f2tDC72JD+xbt2jeQ25OdPiUp1UJCV+MWE9Ppw8WbzvX
PV3I4xHXZOxQPnR2bs9nYt1LR6iAw/H5wgxj6fWnGiEXp7/gKrwnw1zvC03QbtdJW1FAUexTYGdA
KvhO9Lt34bmX2Vf7T9DR0EYuXxjnyDuYo5QZ8LJY+tQMsm4048ACbHKutLFKruv0V3ZTX8oEHbJ1
ibSbOYUa6XVxc+uluWjo0JcZFWfGUw/AFKHjcSviJMki2P271eynpLHGv/pb8Js1Xt96MfQPR4w8
0leKyWbvBPvrhXVPW/UR6xX3/m1roBffA5It/nSz5HiEPwcfLzR1IxxzNElNZQkPVFvtjgMcC5jN
BmbL1tmo1w3I0SWet2TxidxvqxORuCXY9v8PTeCLWHGatnQhMbgsBZw383deL6O1ETGFhhUWOgab
i0QTj8MAFic2b2P09eLn68lH9RrOIWbT0rMVehsufCLxKsA1MSzIrJ/0CPM1wolpTAP+Ky+9zNcc
a4csZbvE4WU1AjrqTPOPcDRUSazbIEBDSRyIxWfJdYNlLHytEWbF0WVFPc/IKMIPTVfbgc2wsDkG
2dHUv7vkeEF2HXgAukU4WTL80ZkdlRbeSm0mYgfCHKUopcLQc8iS3JVnPv1hmqZGFe7z11jU+7iJ
bwSunOQlHsDO6IT+IA7RqxcjUDKzfZabGUmEuzGu/UY4+J1nyT2zn6+nZZm/wX9yJAio42xZE40I
PQ7DpQI2S2Ri5h8oEcIwTbclVVAgojxUXPAgjTVraEaZHLSDa73psTVQbm6UNhJPEmWbqi4xNbUz
sSWtjZrasi5UZZhxjjZsBajP3EygH1bgv7sHwqFrhBICinU7mFlZ/Pf0XaUKCczHXtLeGmtIDyNz
i3kComA4TR906lRR/82mNzycE+zdQ1eoOPtn4Zf4jOSy3noLLSLrfmcjdyvTRIs1E7m2ltw3l16t
QExQRk+r4jEvN7unJVIOu6pQtB8efhyZvMeS+ivIWJGlFhfgJGJ+bDnzMCHzPi8cL1IsgxeR15zB
/eSuzMzQKmPEGgs8tGhS2kVvYP1Zgpv8e6xO4aePUWX4/BvMh15ppxTGk0mKqIY6pR3V4p710Mov
3mToKqXei5AmrWIVDZRjPQTNRCdMDporfnIVLn5ll2xDJ6j2FiCMBNnr0N7Rx3fPPgbwtOhY1mWE
EGZ54kW36anURHK24QTaenpnv6J/c21PbPDY/91CabkFrYZ41rBPYTCN2mozg9Ul47TjacVmbCi4
dYdtSDi3nBUB5uhfZbcYY/JCnMptNKr5c2obu3vSBTrMz3xk7nGOIaerw8HQL2KoZjs9XoaMn82b
HWQlMEgvIEHCTFjZknGYlA51RYE0zuKlVuLJzYbzCB9WH3rrW/CJ3Atatn5lWlPF86sZAFez6mve
H7/hBWbDWYKOSuw/mcuIiS4Ul05Hhl1RyuT9B4aoBRB9O5CdT1iSvNqlrDWWhfqeNTNgCkoB9xx+
ZOAxzB0IjBpjAluBH0GUuAqwJNSIrYQdKDecfa1KhDGxyRc+XHwjFeKWqF7DjnIkdlow31p3/XMr
B9LwBVZjM83KLd42b274N+t2PsUXTnrXUeAGEk+ix2XT3AN+V5ge+BKerzjrrN/aiPa+M95k8ZDg
DRHZI+ZNxibFX55BQ0a87v0gG+ZxL6ucYEiqxIjhSqXwguTTDruxlilxzI1AHyNyIajpl6mtWCcH
dA09ZfogibMdwXZnCThzGoGjW85WoHR1GayscwqcTKBLZq1BeDc9LojODXSsaJAeNapg1VcCZ5T5
CX1fF96s16SoWYuSGUoCohBtX1DSpmzoaEzdb02crkE9ATKcKo36njC1iCEVjVJZKtYeLB6Kv66e
ibyJfrts2l0+ytE6B9iEBXeS1U1gXUGZp/kZLZTjwJEGBsjGGpxxlQZcS0ezS0i17mjCK0P66WBd
1b/fRCyWvwwZMiWHttVwG1MZxid7HSU0IdhJvjdWQmqYQbE4QosKx8Mz16KC6cVXXUR0E5kvpKwb
G8GksBhjh6PZBYxZtnewc67yOPxQkaFIwe/1O1u91dFxbNYm0MVSPmY/y3YoQxqY/zPFKxQ6mdfY
t2mrCpBB4SpLNFgOwVxiexXKm8g0Xrrf7fLNuPV0QjhS8XhACcpagRRhk5Ue5N4xf/vbh33kx1OM
+02VYcjxBZy/QvEUheBFB268GuKGcE3ePQQGxQYBH9VXjA1tZXnbKFEF/UfhwM5vUvKvm+rGkYFn
lzVyeb+Kvf3TFC5W3JJ1kYRQ1R4PtNCFnQz/9IYo7l6E5BOXz1TUtaJ92sZ7L2V3TduWwromwBZf
S/3bqDrdXaw3nFWtBTf1r0gWyRxBkFEHcluqtyKRXGxrHlv1o08MPEVwA4jtACPa20l2h2gCzZWj
qseWEMTv3dd7gjZz+I3i8oYjZH/srghoAxN+TQx14b1A0aX7TK5xTwWECUVRkyLFqX9OwTYyALsy
ik0EHFrhUl0gqwluPrwHsfJiffWXzSxJoLagUa5EJZZCTcU4s0/64hk3uAWvU7J28fbMe78wMnWj
zfWkZRvO8fVhQBhiJP5hN2FpgOnPKhRQtS6q3X6WTvgtJBYHMmaD2HC9GsEEgpY4vRSaAaChKTBJ
bllN6JkYa/lRY6n62Mu4Kzkf0rjQTPQHLHJEfGjOMOW8IC0tehMVzRXt/wSt1ESCaSbyCCUfQrui
HMu8Wzt81SWSgWksyynCm1UTKo7C2GO5zGtmXBLyMatUrHAG4Ak2ii2V9IdR+XO2OUeDTyYDQ6Od
EqLU8G7ZpxSQGEVDVTEeCh0mUDCUVwNaet6JBYDSVyqqJVjPyTQxXjU72LTur1Rs4dTxo2FpFj39
jC8RAybpeNxpsVEbLLpM4BbbqDImyjibEZUGqFJWwO8yxba8l1Ttks2CUFHpqxRqn10nvQScGjiw
RLhNyM8MYJOjrud5HCNXYm/ivJn8o+/iLhsK2zLlaPenDijM+eAP1/kAMdjkw/tzYyCu0jg74oSl
T0ZuOTySOgtghwMCbL3SIXzPpmaVlmeKZa+Xz6/KV8vxc2+sO7qwhfO6/KuFjRSEJbRl6o1wkPzd
KlwpgbIr8Y/ANd8M9E6OI5Z4lOysCIMkf8klB4Jgw+QP0rewHJ80iGpufK/GQwcfhyIkXbC7xqqm
nhnQXnjuUhJM3mtySVp7JJ4luVFqqwDpJ5m8b0C5ki/NsGi+wWBl5lljUMwioVCaVbcEqaCze8oE
RjRcbsTvS2glTC5JnOVp3BLI6fjKZV/iWYeYaz18rwg8uCZYIUFJ3t1N7bI8Lrd+8LMU/0HhI9Tl
CcnFjJNLCjFBAl7plt8KDzXml8n8qJc8GkMZ2z8EjrN0PM4CQuyxQEaMoKz4ngV6wkEYkkARlqNc
gZg7lkprnBqU4hqntgl6F66fpnu+xQx/sisrJS+SWOTyQVdOSVsZc7b8za5jx8k2Vtl04PqXQZ58
FN9TqxyqOvk9QIT1uqEDEsaozclzNX2eyR16EPLhMJEMMVBS3h4HotrJY3ehfuKttxjf8rU3BRe4
44Zcc4h4D9uAYcTfiwW24bezAwus8xTWMB/x+acXKFV0Rc5kgf/vszNVgcoqGG1rE+JJPnQ56Z2R
q2v572n2bnUg43ybo9IA1WhiU7hS1keXvZrsG+ioYE6ElREb99bZnILsFl6W+33zZxYzkwHjSVnt
MY3T5tsyIUYeq5vcOIrKHTxjDj/FuFD0CYLaN6kUN8fmF/V9lLLBo1piqXV2saiFGKW6f9gZFFPI
i2o0Bh0AXVO1WBaElmgbRTHb4aD78zE+VbOUA8il6HhdFz9mcmbXwldGN1z2a1Ud6ufmkODJ0UXn
W6f7ng/w0EqO9papZ0UvflodGaonZFl5xQyAzuyQMC+1gp7FNJuolnlPTr+hXFrmjKh0J2ssk//3
9FVs2FXoV1U9mbN1ZRMJdLE+ftow64NgArYAUp6Be2E88fs8F+TGuRG1971wdzujlILBJsR4kK34
vmnZq7qp3HjKzzbnSGk5lb1mfPZvPOdYiiRUQ6iBDD776/ScAnVDDTmwf4LjpjbeWxpgDfUUe89B
+N56+9uyoH4nwD1/ry2Egu9PiLklHxuqIFn51IM7CTuB27Ii82ZtcImFSF7WqVSC5iJpH1KGpUE5
XcCCi62QIi/blmPaauWHxVW+1/XxfPWW2YXMvzDzCzEHdWIfz7SjCB1XjDCMIrRibFAAg5EeNnoU
+pLQljNLaXBhdyPm8YgP9SgI5NtyZJHETIbI3GnH2CLxoAY6QNEDQkH8fbxOVXObaPxCWLSPKDLP
M8n2GO114cxwA4Okx4hNQIj1h1h0eJ/77cYRj8OlV7VRrZvav2uomhSsH7x9yCuXA9TYx7mskmaJ
n6cfGQ+rufk+TJK/QmPWDnq9rWkIJFkMBOVbZ/1+I4J9JS+LWdbhXTusiceqUdOnF9LclU+ebNkr
3d0U7/8zVhLFsquRzJ+lmEzfqkg/7nMLYzab4hn2kj0RFM/+MxHiVwgo5QXXQ9LZctdaBpU9X+6r
JOj/qdiuKKopGAoqiXbYKV0kZfzVUCaqz+yTUUrdue+7wyNGJzTbkfq6fJtDQPkrxE4XZOXdqxwn
KzmRF6DvNbqTs+Xhc2WQKraMFvgy27zDbRX1dgZ7jN5fRrdoOrVRAMsvN8tH74p3XF7GBoQX/Wh9
1j7Lcq7bsXmRicabAbeygOBIbCks2WNTezYBQaqY3sNL38yi9BK7fqw0BGZMF5suI8931dQaR+Ud
GYN/DRGy1U+zJ0+xNRGhYaQu0gV5H3S1gsar3lFWnCH1c6we1w2EXUlJQgd1gc+aiyP8PVKPqUnX
o9HfPFQNdR/yl1zW7Kdxsg86QwobsH/t8ogve4pkgfMuZoY7xFeijZfwAekh8UCs262T8BdJASq4
kJEae+w8WpY28auFuGY64fl5gRAnIRjVU38eudODEuvwHyzuZJJseJFYWb9jFwyICw224N0OfSWP
hIF9HVjZKGG/70QYXiRT73mzuxz7M0L4E7RxvVJbJ8J8dJK4jkXN/AtuEB2RKzl7U1h3xbd8IbGs
JwnoqkfCH0Oqqx7Z6DJ8hTlnrn3C8EZu+7U16ItZhWRdSkVrwcpm91OSDWhy4VLQNZbfCa+6szWI
HS8BnHDd+dJ2ap8b4/UKg9kORLCTOhlzaWshGZV/a3wNRLPzNBAVYWH1LzW8s11Z6560Vms857Wl
HVutE8BUP+DNqcZCZpGE37L2rPT6AOMkm8hr34pDy7A9n9eyTwq5U6ARJpVHoIz5VeiWACzARKbW
b9jBaawjUFAAOI9SRMvwPLC+knZKynVj7kiXlt8UnDvNrPukO6Nzwq4kT89Xukds2ued4dEQdUVz
4ARvvuqa2PUwXQicZoefKPTaL0JuwEEy4DbjBOXv3hlR2SekjPsdVrWXEQ5mCK0MXQJ8QisRnX6d
2/qCVaVn0ISZA98fJJW2XmfuOByO6nreMPqlFByUeubxxE9otd5OCt0NOWhzU3mnOV+wXkXRbMS9
ZuTjsgSHRQ2cU9h1gCHAjWgH3uQrU51Ly1Z+To0nceamjCN6k6kkr2TCkbf6KI4hd0xdeQ754Lh4
nh6Fvbqr8fLKVmaZ3+rvYl3CDWMHWrRSrN0GDzxgvJmrFIzndfftnMtqIex5JPLUZWXW9Z0lBLuJ
/Pq9E76DnNZHlcnWmihmD7bBTN0XWBKu+mFx1nkdmkltxzNIpY+s78lnNEdi3hvAVsz96ZSJboqv
PxcdDW+j2sZrZZGqyV2g74IYScRLZGdZgqYfEXW0pWewY6OIjYv1gmZGu3bOpM6WxzDr6sx8Id2v
Chbw/kjv3ucYlSGrzXItNbqpKjLyVgtc7B2Gkto91xTsBKKuYxU1Qap72JzmOYJTYAeD12t9G8+B
hRraESzzR/quZ0FepqjvSmsFEezDqaFbiPTuMvN3TyJtqDxQ9sKvweQPtot0bsokm5ELjmuDohRQ
DxpGUapHGfZiGC4sGlXWX42nDlgMRzWnlUwQ7l8tkGyBEqh1fkNgo5tFnRz9pUtnM32BB8NOJSqV
yUK6MSmucFFIPn7nPbfBAvHSbdrzglUG38/6DVnkXPal9w3hIH/D2wNY2bvZsZP8C6wAyiVqWgmM
r8qw59MJJ6oIxzGF8sAF5XeMNeauVMYVWka+i7zCwFCZztHRen97xW90kG/u0FSCq2GaHR4dRS17
gwqKj4Kpxmht0ezHMLAeQF/BM+7H1K+3h8TBzYJamRTyenasY71Nhe/gXZk+bjMhLX5ZR1btHpZw
2A9yu/Mncw8swK34XwcR8236KZEBdn19QCDDrmDtiJwB3XX196CxthuuoGGQqX8VAWqeRFq4M81p
gxeuf6oVH9+MMxke2WdUi1F+tfqeS9YqrZL2+HIgnUnyd6sCCwdMOiOBzVf598mYh+Zkk1Ka+1yn
slqmKNmzctleq1TD/PTjdlK2sP4BhvngzqgcG1xkYVYx6JfguS4wXGRewkhV86hGJ9roTkc9e9Fy
AkoFggmMnjRUd/Hyq+RF6bGtii2HR321hvsvoDLsEvD0sb6GZ+PhUER6Q5OsNNQDH4dXlYp/8la9
kijJez8EPbW539Uc2i4Fy12kQAVkTS+Em8unT8mBSfyC2gO6MuvSkTt1cHGk+KWz9TbtQACSQFFs
51Y5BAFbZ1E15RmH0p2o7txYnCCLQfJnRokjiWRLM61kFSRlWNLRoYw1f2wroNTyVR6dfbHABQK6
7ITi+q9/R0TZatXnu5lMImDSP3So5jS2NvicusGCZIpMroAp70fmeEaLClfsBGLTfZ9zUeYYRYDD
9la2e/BpkaD6qyvMnLF1CUsruFUOp3R992ygzv9hAcLOc40XEa55RljbI/NAhaDVrGWyTPCdLLvl
LpM3xR3T2b7ztY/NW1w4/4xPiTu1scdCICPPTfVDsDj8JRYyylkz7HKpDt0chl53yswWn1xuhf7Y
18q+r0kq4jI5eejA23YXsw73Lv8H19IMQm8JN2puRryXLvcs087e7Wx7YxUIKqPcMUQC5TGddpw2
uf9Rv2qg3sHb8goD8x5MvJtB7Rlg59U9tu2ccUwVAG6TPFz6BpKJGhYTS8hNt/GdBo2OdF+oXSoK
FMlz5EwRoos8aQYMtWLFq90m/Kd+Sbud/LlOi3MW1wnmjgDDEHVfHcMSbMfUB90jBCLIq0smrBE/
FEvbnaT6xHbPVfOMJfHeVPjcaMD/+W4ZcbWEaa4ZZkDU0ZpPi1PZqXXPHsj+58B8Yk37RiPVYut/
EawFrGE0NrKOv4bnnn1vK/GwjfwH3jvJ3CwMoEXW/ZMiLIhFU2gQBCm2zgAuH9E3arXmA5OwIsqk
6OHcYgbqz2w7Kzj04LPTmx+eUy7WCoLY6wuir4TekYnK2AZZRSUwTrgsrDovdthWVHPhq/fXly49
gpl9lIA8rj3o4RCWkaKj2PolsCU0jOOm+VwpWvWWLzkJpF6aZUwrZM9W4nzkV8uA1qOMdZPTHYdi
/pPWNpTwuLNEuRIfj+SZHJmJXc1T6eaDn+zfoPzh/5MkrXGpO5DEydkHYJqdbQmEBL3+399oHsJ9
iYxQfOXbK3wlzQiwflftHJ445wTTtY3Tue5lNc7DG/95vZJntznT007gKsDGrx8MnOROS4FSt88l
mPtfyovRRyZmRsnbnC+NYBgSNpDw9K65JH0THBHI5Dcz+Nu1+v/Ehx9qlnanvmCmfVeinVeZD3Bh
S/Yn+8n5RZiSg0lLGnN3UBAuqvzpnhcYT9uxKgd7WtRvRhbcHssv+jKng3Qm/FxSWQenanS3Kdlp
yTsGvbtspjDDyNo2ovCkzJygoEYV+RXmxLWHeR3nx2WI4WdPhvSw4O5HpGCIdIUTCrlgsmtJeQWH
uh49+f20fpelnS/p+ns2gmf88vEIN0TbOETU+LRLUPjuC/panxLtB/hYfWXZUF0Ly2cI30VTuOa7
dToiovF/3/Z/PWNIjET/l6PmyarxC2n5yETB7vN5foO48Q9d/Vu6AWg2eo7C0yeRdkei8ikQAI0E
/9IBVzkmBy1fE6SEuBykkPIzOfosXU5zkDf+Ks2cMJ88dVvekcQXEc7KLwuol3rvpXeZ0u2IsMAB
FyJ0x1D6NLXXgl7tJBz9y8qpcto1I1/G7LBXamy437sP4DgTT6a9Ajyjs1z68md/G7NFtPgFPGI9
VoPl1a7MsDp+zvaSXmaoFF2WtxhEZWDUGbcRvDbWeSjhcgDSsGcBxPbv4g2Z/+uKYFQ52+1FJjuE
BsbR1kU8yOvOZad0Lnj3YcaMaOPNbCD09hPXu0IaOXcAZgQniA8mFeBXMiHzqp8+toDt+UCauVsa
UoGBizEqE6gKQa3yd51x5K5BZAAW/KcEilIWIAQ1RBJSbKg1M3TRoC+aSD6wwaWGfW8jrckxO5wm
GQ/ueH4IUTJm6FxxjAqhrv/5aRKwJi3luGwvCISu0u59dLv+WLuFYT82gDcxMLajtzhVZcElYYez
4zLJUvDm6uwkOZdeZa9OSNNWtNc+gZyWuuS9TzG3PB0hXje7C3ZXOHMmMzVZsr1mBDF6+S0JRxkd
kIUjj9mCLNCLAXmrhyX1iSAVtJstyPRmgOdiQ85XdJMQljn3Dwpgtuc3DsFRR/ssxYrXIjCYPuKu
a3VFmi+kKJC7xrcnl8La9yxvilvccKc8PCG/yj4N/hHWhnWqmiJLN8c+gC93u6HSqyyrXPfsn17j
79/PwyAWHGOq9gxH+iRWe1f4yTcnIuDNkZs4Ku+DCMqy7w6F8TgB0vI7u3eD2E0Qc5KmhW+Sz4Mv
ehmIMgs7HGxvK4e5y6mfIYR5oSX7DOucrqIH8iWDoIalk5J2JSI91i4PNvFteNTeUKeoK5wn21r6
TWqSQTODpGU5yR+k7+trA/8WqTsmiFYLisYksodO/4vHISdFreBh3LYgd+2a9h88rflnOQeEsJz2
Vmk0HlTOoM8HPBYz90wjTBpSXatnDFquB8yGHeQGDJou9FuErcmRsu1xp5eSjZIqhYntLfJJf1V7
7pvMxXOUbI/n4r0wAAhX2vZ1a5LS1/68pbd5jtaD024+gx/64yM9adBTYuhGV1JIrDBctjGawRWV
5BaK5B6sTE8FlKQg4bpWYtMYI1g0669JSgLqoWMC+QGAMKyVeFGGhlczhLZnc+b4MiRKWSsz2CA1
WhP1T757lH08xYtoTvk4uRr4EZ4UKJg5BVDZnDwjKwqW++o6eq60hrwO6JB4478/offBScs7pJp9
YwSlbi2V8jrmZkrUnwCwrbBnrwQH5Pzc331r88AvnTAaIllPSaAR01vzaweH/fnNl7kAhLNA+zQe
TqWexyL7MTnxAnzs7Xs5++qzoHjNBt3X0kN5io3DoLHSe3Es2YzgxJWYcHEnlbbbMfsisZtDf5tY
C+q5cOXJALYoZGyOLiEHyQ8C0ElLf+uIHTQi2ewbNrQg+grinL2SmLySdpqURWeKZcFu3EG+rAk2
96iIybiB8g6LVDs4JLOexw3MJZJhAm4g6UeMcq3eC/CjppQHvYYFAzV1Ex93NHSw4NT9kTIz3D0G
66aXV1svbkZP1RyvOilHzVO7Zr71wLjlB5tFewo9HuRBddPD/XEp/vVwNuENEBZ9MoxkpJmwPiNn
JSPshGz60pcsXbnWmA7PsgqPVU+QcrDzc/4L4xRsaMz2Rv9coo93NJ+rXIaurgICgE2mIfrJC2M9
z3xTizcIgHYz/OAF39WN/tlw3JYr8/CzVncQdvYtpizRKyWAceikMieEkB+3OzDOxGnK87ts2ocg
luEZjoZTm4ro5wJxQRC3M71KU9Yw9yxwt9+autPmPWC1jn5PdSD5hU4nPovKBqlSRkMcj1jchx/4
/rzV28bdCqebXLZjfZuoOMqOWnZ4UzhuqTFA2hQVrbSBy8QSSg833fzvolBmo02ZkBg81Mr6r2+0
4vV/YxMZWMjFsbZbDboKC0/aVuBf/uYsHid2xw8fuNtojHDVU7WFuhhhmBSO8y8lTPZB/4UEtrwN
SVGfYf0BClGhI9qMdHdoPbVeTKhrWT0RYZ9gWvaU5vBdRAckYRg3PjTVi6+SjRpH9yqq/7KS35jI
qsIlYyJtgT27PVz8XIghhO3CnaYaXk5x+7CHnIjsk/k5WsNTnWscAObhy4asRZoGJdHSwny09K9X
S13woXoOWoXdxv/KVV+lAnn4fAiT144TTj+6kD9fVTwLyGnt/p3w1Iwj/Jv/3RmmEsyyggzVo7NU
SxA8rxmQuZ1bwDHLDtAjdhHcN/EJ7dUj00mbKCF4HhtMjmdekvCBikSF2yadtd8XKJAfJhKhPopU
ZcGdsRFcCxA40Qlmy3V9U+we+7QIjweqDaB2LiUswVCyEt3CeKPU6nc3O4SoCuUAUwzTV7htwBg9
lTGifCITiNUTaA+X1/Saw6HXSvXBd3HJh9GFdecswGg/RtER5hctnCVVYdkkLPphwLHr+HFn/RWo
CVVhgUmBH+Qq/YN8XIc4ATLkNHkE1J2hBP/f+ypqwkG7jKcszWRNeGnG9hmcj2mf1S07BCFO4BA8
13wQRfSWN88osa2ztV4lx1ZQJg8gz8bdscjRPdRrJhCS0wVFGT+tOJXao7iC/i9nwWJ6pmY6iDE4
KSJncKuj0cEW3sqIHZrXJsOe3gyOUmaWx2URE8G8TXS7udNDZDVsbAvB4SZhiIfrj3KeQvQfQUN/
zKBy4/G2/wLOARIF/idb3Y17f6evaOtXPSR9m8MFchBnDdgVS9v/ACIGsARCYamaxRSYkz156FYC
55wECQQZtDTep++17pJxsWZh0ivw79kmOnR2tePIzK7wjvRt3dtMqj8q/LT9L/Td/znLpFYXyyI2
LYIdluOvRVcSuLBWoTkd5jxHM6WzJGbMV8tCrt+cIQ1ne3UYtTHgiGSNyFUEV958KU1mbQM+N1jg
IKs3L0TfYMRFm7wJQjwf3HoVpBf3LD3GqLgi3g+Aje0Tzv7PDHwk/wSH/3QKoNt1tO5m97LDRX2R
oA7CdqG+2yNEBfFfba/eACVGXiVbseX+qPyhACetBwbg/KB/mxtT5JW9PEkVE1zGkxDT/QOkibRs
vKtpdyHWeM1O/z+xpYyKEc2J0Wvf1Ur7W08yBANHQU5nu24AJcKgJZTOaJ3h/GAixRHNhSoiwSH4
h4QtlT9lUymMQX+nok8lXQ6s9UpHvXJO/GnzrLN9XqPxPs9GLadZGINj0hNJdcTpsKnZsAhhP6kw
oKmuaQDvGON2iyXs7bq4OaFv+Vgm4T5KR7WpWAIC2X3wG2CscBBLakXjdxfQVwF2c1dGw+jbe+7e
guec0KBOl0HJ0HuIoAiUIZhB0HRHwGQVfOun6+rXalMm7NCPEr8MV9BdSKFEhEMf4okeogL0Ghmm
wP5HfCox+Uji5T+hlWOizGl/znfzBVX5k8kcSQK0jtFTdKLBaZptvZuradvbYetMqmM9iwg0kIyq
UT/E4u61eXicpMrzPeYt5LuIgeQcU6uddtXuT7+dGb9gI+vF3gsF8H4jWUA6vtIyu33ONxfT5Sue
UGEfbb7W+zVuukLBRjFZpdsNW+V1xp1wJwc0u5R/9UIRYg09uhsuFysLIFjV63935BwcOotFnmkm
hrAh5CwCVom4NtsBEZbkiCnB5hssJjXyc4Et0Swz8/K6i1keJwGJoQduWWemFOVKiQlhkEgev4ll
b0bEApndeetdwhJRNRNUFRSaC4eGx0Q/+RKv4i2nzgw05p00pmEKBe3wNVzTkNABQHokWAUHylXc
3GoSrPBhJ22y9h+WwiWuuMovJLBqaV+w3RdMTACQO+C/Bk8z9UaSFZbDOuJ7NFqPOr/PNKMeLtEy
DT9dQlPamHEKmdBUefPsiNA56TZ+2hm8AHVRYh7GSLF+mc8YSCnJcur7gF+xjcrY57x/thGqIdWp
IZpoX8o+bmvvz8moedjiON+o6DhBNH1fI2WRlSLRapaY4Xl8XuZ0KLEg/v2i3/Ai2sgqGbJOv3G/
XdHR4lFsVFKP+xjSrw2DM6aWqMZMrXCX57a1R+Xisl9iG8ZaL/98wZPbx54cGqiFMoADl2RyrjFM
MQlL/Rd0y4aX+iuaftaV/4GLWmVN0DTyr5bO+ajTr/fg+wwPg0NMRycfbdt9K4181hM1wmQdzKRc
ERHKuge7DGvW7/wHGJNll8ubn7D5hYIpRAzAauSX2vmjIQLmQ+0AQbPKepugXQuJA2gVonkVxLz4
i94++VpzN3qPNLmZC3i8oa9VRulMH/971J8tu29gavbE/qfA/14FSiEgvM7o/vypVOP1RGlBK2QF
8ojoToROlXNPSkKcs6YaMTx1OF4OPF8Pr7Vx9BevXeQAZg6/KTUeijV4yxG4SHpgH5/eN7qEq8k9
V7yAeyZ9TcgfqyGeWOwxh+ns6bSFgko177v6iVTSPuGk34NCL/F30W/7lJbiPt5VMaWa2Vdb05iS
30Rs6tS29meE7MQrB90XDkoPczjerMFGwQIDJzVVmSTK4jrR71lNs0BZGYoUCPe+TenY3bdqrZoQ
wYPY2pxwi1TfnjV63vXTqfxlMNxDKeYQ8kGzRQ5qjf3xpJ5j26U1s/mP/+Jf4vxGRSrExymxO/E+
TP3CcTVI7a7As3mKBBoXY4ymiFUvf9YYVHKIHm2T1gHFcVlg9SYjvFEDb8e4EvswfVPd9TDXsMtL
cGKKzcgSYtyPBAmct59JZr3JZ5InZqn/nLulJcLqCkM4Dcnap9Da+kjnugxPnyjwI6gf3QotONyd
KcuuxkbZD+WlsVZLGLVECeFo0ezhnsiqJvtf3gJN7CUyPrIjTj9o+EjGsEal/I7RF5yrCdOMBGDB
eUdpZ/Q9TpFxoxcdZFS9v+qyDM3dCpIzCDxc5UCpjyKMGil1kgx4kv6WBtsGm6X/RQLgwX8V4+0e
AqAhn4r2zmAltCxDH+AF7l5C3mb3GKg4XBGOyIDu5uu15NohYUj9GPdb4NjDuXbb70FzOyO9bEID
aV/B8vIOtTr2FMw+W9bWtkGF7VLfVnhD0v6uLH07FLF7dFJK1FX/qIv6SvpFqojOWLeG9vMNestt
h6ZSb028kZr6j4xoRaTnraYlisoj4AyArxHfWiZBqpfWpuraJ/KqCxbNtHI2Ie0T6JZmNWVzNhuy
OV+G6+yRd2c1x2xEq6HfCeBL3tA6OOPiOZoTRbBdV+RE69nQfAHYooYbw2tHD1Mbh9egabLL85Ys
WHXYMMBKrPalXMeMt9o/c8rmHfA8J+HSUUi3AylMeUHDW/YP/Z5Szfviub0Hzlco1exfofRU0IkG
Bz/bWlXZtYEtC0Dl0E+OWocSsB+aUCFZ1oIcJtSvvkRq1td6IHT/9vpysVppDJMI6i7R1xYqKPFK
4fNDXi/Y7iZqjm7U6sxQKtGWRB5Cu5Bb78vThT4Bt3CI7+AS2IEK1gsaeFaOitLEOa7l+D5brm9t
4YalDDdE9IyRFxctJgeU1enUv+F+MOkvG5FfDg4aRJnJBE7zfqiUSedz9B7c+rYjBL81pR8oMjAB
jOcuceC1/zNqmz5dewrqYC8tP7lgxK+S7W2sAsOCYCoKYDCaw12/krJd3d78P7teqNJqSXG/gNP3
ZrrSErd+bm87ccPico+BlG5GORB3RlYV6ED97keSd3CUcIRQmVPV4V/674DDLQ4MrAOeEbmDFmfZ
ImqAfAybQWVL04igx5P1EZb840VfuCEiFkobXPZpx7BKfCMVOQU6AY2wnDlizmofng4e6FZVMB+O
+3bx1p+CHukHUbzHgW2Sc4ZjjesXZuscOlFoxhGIQI6qg5keeFqKUyX5daVQyCd1gXy57RF0fLMg
6tN922RSQQE2qB8tvuncLeWImexZHGLdQfJRb3ukaXM5MCDr3bcFh5QHGvBvY7ye7gt5QRE7ud66
Yt1NhaqxViUJDYoLDJq/OJqusoYCU9q4rNIqsn3GyTuDdKsWDS9je+I6cx46xkQIIZYwmXtBeJg8
jxAbZN5INSHtk+18USFqN9bem0lbcniDa7FqHCZPBLasQ4VcxkyATVNTZnkc3Og/LL2oIZ7oneQE
LZYkx4vQoeCd9GTtXirY2mmx0aUQRD8W1xOO8M0vKmP7jPiV23qEUDMCR5MEolbTNcT/y85rQkyJ
6dX4PCqi0oj7/ACU+fJvPrc5Lfu/Mj26fgkFeuZVYJGgqkJ9jLTvPOd2uuiIkwT8YbPceNoKDotv
HTRy+h6glGVBh96Ok95u0VqqcAZILWmH9DP9aD+S6i/qPwO6l0Rh8eRaCm78xGo53Z6pdiHdgLGw
Iv/JYkYPyWle/LEH9txFDovLaIeTznOy5wWkIEfVAwpv9N1xGlovjWzF/0F4vO84F2bqkJFqj1kL
ZPRNeF61mp8FFo6l/0weD1XB0NzFGWgY/hjyHZ3jrHoUqkqQFbPMq0Qd7k/UydH1NszJYNbDQKDX
PMQ1TjLdTWrM3n57la2NYoSle6QYB4Nzf84SczzVgIM5mn4tftAh7VEL97V3AkCpavXphPltvakd
p6UJ+nOAWLwUJ33ZwuAZw16e6In4I7MqvhQXpbBKnfBEkAqH5f/swhSeIzCsqMi8N12snhJIL1dQ
VMx2CAHEbQsXC/h4dMlk+9zxNmj51WsfmlSWatsyidszu8rwGaElHgHuSyFldLi7hAPWqvrZZ1xI
6VfYEnT5+ipB7yIp8u6se3kRLrC1AYjNxD0Wan2dDIgbBpCEmYOD6ld+/nD6JBuVWFQsH0/inMLJ
BPuw6obtVgKXDF1vZ7s5nB+Y3WgCP/dn4Q1PhoBwX78i0cAUSPFF9SjGeUiMk5medc+7dJER/DSC
AgNVp0Uq+1ZuaF9c2WnVHaA2azXyzHvN2NgaE7yeAV7GK5A0wJh4VZ3QTIWtV+3ekXtZ0yTvlU6V
WaCJ4fqeBGeaFgCA44+VZ81J59Qb8qKSJFRbpqRiLaqpY4+Dq7QCSP8ak5r1l7KSNbKlZx42xttq
cZ1s9ztem3mAWm+KkJH5fuV5tagyHYXQO5pr/xqRZn8GI+4iic+W2p5PHvm98urqJaZvhoyXcfFt
e3xHnkbH/96AC1EtfFvWwaoJDrAEQnek12I++5UyM72S/+P3N5vJiQCzx2JZPCIpQBL/dycfKBOX
1AOrhrJWOxrWM2HmVXhAMyy/OiVqWiz4wa1MLSLrZEKPhM8Olji1Vm7GJW786U1FATquIjqVtovG
S1OzfNGKzm2x8eKa9PaWaR+seWLpRay8w6cwTWNjQf7N+stxLXMIKgIuI8WTxWLC8LTAITR0QTBI
75hexHPIPxPqKYsWthwnpnhaBH4jHGQF8O63mq+wHnipvBXrEE9s1eLSLjtuONA1jF7NsXQWndEb
PKlAB58fUkfCjW/CEzmT7bTSru32kF6kuWaSQTiYc1tINtriCdE8ROKshfEotpo9IQe14JZsBlKo
n3rcGpk/ITSZCGGTYODQ7LRMo0l3Ef56qXGiCGu6IXsoFP+bz4BWGzKSq8eUdb6yEk4Fz6U5TLm6
9wBZ0/xaKv13z/Muu8ktq3RD2AIR0Sk182zLWhsav39p4ltfV/YIup2FrlcCCR5di4mFF2njJbH8
RT+cCssYq34xpsUF1AetTWJBPHUVx3EAi+ciRFIsfJuD69EIrdQHsVpWNnlhDhG+38kLvd6Q7IzL
O8RECCOkGGYDY5NGFv0sFpA77YOke02YC4z7jMHBUiGSA5LqGyWO6PypcMnrl5hDnBfddwDs8h6o
O9+JUYPd6nTGq8rSF3QQgTcG7a1xu0tUJo50yVU6FtXiN13AOxlshtJqw+/h6/bdBLtujMIWiDzE
OREVRH6jPxMTvE5j5PZFY/YDssSwrzalgwp8S9IQSsFqVph2hUN1HYu4MR1T6gWOdCGndDqfGQNK
tv+3aRqFx3eHNGzJBBryf6d84Lap3+EZ4PpIl2TDm6J6AYMDe/cz2AzSbaBOosFQ1LjmcPVuvES4
fZ0vBkZbiR+rBGA96xeTrEcSWWZdcxhU+jalPq3ZyYvxrdoKSVdUGqfmq3PhklwSoMxSA0Gv6rgu
tZP1HqBCeePzsKzURG+6seYnO5SMRPmYYft1OPlKO7mrqJgu7AY54Lr8HIkKa/ScK4QJyuHgXVkr
ZGvSrEkgOM9dBNbAw6pnNzRMVPgIv46d0IJkszuR5dofEcDpJmwkwM27UP/7z54ggG9Y4OxQxgWq
9uhjyb2GlZoCQY9uil1VNhw0Yu+ME34gFUWl/gydo4faW3E1LyA7pUlWhyldDT6NSenbndt7Rey+
GrOpEKxLEJCzPwELmeeidzTjdXV/suc1qwQTTUs0s4k8vKBH/aoCZt7Fyzhn5ykdYfaYN0ZtFiHL
OX6QYu2+HnG8yRfQbgRFjfPhaMxCkTa+T252qqjzm4nvluQno4WOZbJcrNB482WHFabGTs5zRgL/
IZNVLUcrRDU/jUPNFdm44veigaiOJHSMjDhtHxzCZPYXeWgv1RVr/gaRlTvBoCXB5Uu/gZtZjwYH
fZcrE3rBAs6eFGmE/OdWAX8nsQRMpN9LGahefWo3ecKXV9qTwGPfWAC0Hbjh71WecuUsDQS7573r
x+MEEavY/71GO6BWFlAPBY9ylN5c0B3u66IJZHfEPM6qg+4q64itOiEtyosHxpqk+NxYZKnbDLOZ
LEDReGTxbUb7PhS5bicYHjTmYrIlrNoTENWGP4lalUMYJQOQxZ7/dKzNOM+Xf4rPRyI2sCwOd9Sh
eSwJ9SnEf4oUj/+O0iX755Gf8QuaxnHJvpnusqmVHm+fm9E58TicYQaWVElS/hll6TjNja3o1A+3
mEa2TxgHlOUMDmGV+36jy/tp5A1SUCTCbJTeyVEj46s07cTr9HV2j6YqbknzW1GvQfRyHmlKl4fO
VTsFz9lJm3sdFQmdNl6V7VUTsCJS8SmYWAxRpB+bwf6uWOTIrBklXSK2yskLmeloJDMbKRyIAwUv
d1Y6wD/sMlhpOJjaFFiVBQkiOlbmBFc9Fzj7FsyGobl8JeyWG6MGVM/H8Zgsk8yAwmeGuqvqpP3G
8MzvWgEU1GjWx9LxLM7Nz99uleMlEyTnRwy3QnjMq6xK1MjX/FEguNYYkGHHs9jsX45eyUPGv6V7
v1zBsxpC5NPnc+z9ckPFxS9UATZ4j8G81YL0w/io2XW/UtvHYSi34Yd9oCSHRmpNXUYNDOk3fpgV
lij3QEsQDkgiH58WRm79KJ5XFohcZhe2jr5HC9NtcUGHUVbqZbVn7NGe7Ard5J0uLHPNI/l67qjL
PUQE6PKhK5GYAZubi1cTWPWnkM+6imoZRyAfJ2Y3U3lgbLyzaq8Fj+9CY3gO27X0w8GGxVIxQYQX
+bka9ctO2B1pKd5VSanibdRJ2/F2n3yDD4/VAL9AVN5DIo4+2JBIiAc91o1mus57rIbOKGNwZUp6
Lp7Z4ybCngWzmUQWvgGfFyYL9HmTwcSRk0P61XJofsE6VCEx5JdHZZo71ZEA78Qs94yKYvCHsxdr
+ZOopZZzp0AjHsLu9IKZ3+/O8QfMokp9v658Hk+ZSeV7iCqtCWhG+T3psmfW4ZLJXG0Z08zgmO6K
Q+xvndf628fyt1u4BkkABA/fzyNsmbBo6I2SdcfuE3FeDaUtakXa6Zwq5WiOGhVNL3CL6UYPzGi5
44d+rxd///dUzDqN6WkBxhcy/usm+3jD76i+WHacJrqCQWr+m55OwX3h9O7TIJ9sfDfyiFr1QZrW
Zw5K2+F6LUlMy85nIYdRGld0Ne4DwxYkerUZrGygrYTq/I4Dot8lpQl1KBzvnvgbMKtVAgOFYLQa
T6NxjIioB13l3K8sCkVqoNNdNiF8Zo41rbN2cz1UYDwcNUBa0asqWlCV5o6O00bVdB8R0KdE2Qy8
oeZ+2+iNtecvcCwHDX0zjiEQCZRwbriKL2X789SumJf0p07B0ijCAWArKsN7FbH+CB31aG2ey7/S
o+ll3P2nGVv0jmLSTplSDz3y9GLZAuME/X/XMR9+MQXvtC7e83+0vgFjZw79g020tCKQ1z1ov8OY
lwCeu3TD/TOK5mUHMqh3jswHYdYxDi1gDbf+dLw2y1QExi3sU8z1nEzxS7dqla8lZlKjR+fDJA13
cQK0Y2JCXpNcymWqrY64z1AGfsrafVX0J1eBhe0tPJn/KqvJgonfukNhZPVRV6vcSvkdxbtdCOP2
xwALQaVBuvwuY9WUUcX4mjqtTlrHw16ZaGKGRTvWHGXb+aDIBWPecvHUbccgwN5c+uUToovBvfGv
t8jbjZh66BITRxoNdDeMG2NzEJFRyCndM0TFehlHTgKheF4CxZbkZ6OoM7/UqzGjWsGZAm5qyr9S
9+iD22io83zIZAvZBP5AGfTBLHvZnY3AKZGKqAVfweg5Atgf5Zd1tsS9P4PK+kS2Mv8L/133G5Dy
GYniCcplUUZkqplwXOdFMQGat756XoKGqF83B88Dtbbzf25mPG5LynO5YL/DRI84dOW+OEp9mlbs
98+ouPhvp04rz3C8vV47sgK7u+3/L5TSfbcJmJu8MY/nKFSqaUT6Q2OxNlPwCJSlOKtaP0I39g6Z
+cXiUxt3bqhB1nw4WMfa2FRMGV3We8H3YoSfs1B+t2O9jlzGnkxRLig1W98ghzkepFBLIj658vMX
e87RQql26S6SgKOtl3BKw9/oONMlM5mtRXKCqavGbmJid/gh9FTPuqFDFsK+JJ2kUjRzLdbaFmqT
uIt/G07JGX/OzZiF9u85XhMoWYeJGD1AU6++hBM1Zgys5ICCgYWMurUKrSFSwVZOPSFa/sFhXw7f
11nJKi88OeMEfZubPEhQ5pKfc865Yh5ywmpiCMoEY8nks/wVaBtFDOt/uBMDrpCzE6m6kFyZFjnn
qSt9Gugp35zwSKsCNYFpf182KBXoaeYDMkQxF6KSZPEo67HS1F4WtrPg0BXU0YbgjoFdoAmk0L3d
6YQ3+1QUADmNSyp+WFDUCY941k9aTbai4fTEk61y3o1xzbm2WJRdyE2unLs5k5SEuJSO98Qbpv2k
3Gdiu6i6tLRIbcZROE/ag8Gz8w5M4s2GDAHL0CwOo1EME10ezqeb0YXUtjCR4O6tHfWbi5KGYtjq
IBaY3Xy2xxyfdATvBeGIKNQiaazdmajKla9QJ4iE5FuraJ8WrzBzcI4fPSMQlb9YUPkCKagbwOcE
FhzKaWLiXkL5sm4OpYDOJsTLFL/FgAAJdj1s1PD9eE9sitJdUfyGYR/DTaSTQgOgM2lQcHf0ByLK
n2VaIJuxvL73rxH0XWqnI0L2ePNvWDff3w9BhKEeM7d8r8sfY8xVScYPfIdqowHhXqail7CYuMsS
vRKwxLPAqJsCTrDb8LyOKQyWnr+z0qDvJ70AMXKcH6jqmROSCAwMH8+ut2fNlZh0C69/DQDwEub9
IlFI07AUTt3fBVFXTZJyF4kD2lp92gi0n1mtmkRSlbeVNehU+OMT6M7D4GepDJYEeVNEvpxRK6zr
X+cgZlkffvfHID2cLYgkQ52zx/CjT0AcylkKLLayteRFsA5cD17ymSu7TwJrUKp1SpcgvQusaa/l
jUyM6IbmYFSthx9NhBZT8+mRfy37Po2FbIWeSjAI5v8V+M2Jrakh3ocTs0L77Cryf6nCxqvRwbWD
M+Ra+rHpwr3ZnT5r8BpWl8o7FF1HtiDUa6jGPCsUxL6vW5q44bsUlTQGRVp3AVs/C/yW/pjmATDs
ICr3lDGhEIzC61MFXrFUn0Y5ERFeWfAEPq6QP/PYRr+zIM8hLV6GBJ8vwZoTnW0YP15TO71GE/g7
OPVNLAbYXfFoIC/cDxFixP4w3YRlycBVQicf7zfpHd0zZiFpwi1I01ah+zo9br+Y39kL7DE7Gtzx
vOCq9jndYaf0ALVKihpP2OMtCzs8RAdOjEpaTpDNtj8aUInC7FhioIRoVTD9IMZh6QREdRU8v48k
5tCKtBCvJrr0tTuQa5crx9P+h5NxBjwNneyEWotrMIunVs/oUhpVr4EiQyWu/ZBMNq4YUiRQvs5U
XUFbUpHs6foVJjnhvigrTH4nDa4Jw/MSKitowrUnsg4VUFAwdWMXxqBI9CPNengOTPKpUHovrkQo
eQt3L4g9d+9xTLSYkdhP6Gq1QhVusoImYYElE9Fb/UMer8d+9txeX3Uw6HJqj/okgojv46JDPs58
bPqLeQb/oiweBsfiZOlhCZOUAcOnI84jZRXs+vV+TOUGM33v62vsXq39+gqAp4+PeVsXUuj7FMWP
gytIx2Na9uKZw7C3wsRBXHZVu6XWgRiO1Zyvpn2B6OTgaIdpjpuB3tbgOu+Y/olFRqZFJaIvzSOo
n/m2P8JwBSuP8CKPWG6IHOiXeaq6nu8b5ERzOC5DHEvyGeiSHZzZncDfDx1u852Gmtsnlic8GqvK
Vepcum54SO82vCWIIRB4h2vLVgT3Gkotaib4n2jUJQbJ/pi9Gs4sN3Z5dtMtApmk/9K3XJ+DWRO2
ikKpsH/veU7jprGaUkzxIbNbiriS90d17ihLQ6Tgyg9YtyStcfVWok9EhA0TmmTW1XvwXnqsw6YT
cC7PRScymAbhg5UcqwdBn8tKczk2XiYG9pMJ02/cjHZZlVqABscQFqrKlc32xUxHHwbkaR76Mhf0
11pPTy0YT6pjmVxX1+c5GTeOtnbeiydFsFdnOMANBXSdP/Xv3k6fJPYPvmQRZ+J9WyhFrbHRDzSc
2RkvnL6vtp6tpEfsC5oQy0NSBeHPCLMwlnWEyneXMmWVdbXvinNsg+QDDYfc/SvUCEdI4Wm9YtkO
Wh7rxvhS1cgeCfWIxHdtMaSVdpaXSPnFr25lvsO6+DNT+PH+vDeCuxeb1b95Cr8LjTlblj3qjtgf
dq2/MxGc7zbUrW10GIG5fmKTP0KC4EMk0YQOFMdtonrJe5iIP9mnU7Ckwz45M7SAOGfchAySYdIG
MMyLCexeh1+VUNLqUNMJt8UWw6UUgb9pzJvoe1MOyFDUTfGjbqdGIczlU26WUVFdEItKYfDKjezg
MumpTxObvUurck5pGAAPO1zW/geE96eiY//suMsbkTS6FJNX/am//hxQ0lAp+NylAysKaWkOispB
oEPkl4X/XoDdmDYk0FDn9kVvnzjzDZ70EXyhTlN2DfgPgSJdDF8AXhGyq0alkw+FPRdl4LWnJk+0
aEQ8MRFJ9z8vOPucfPpKknX8RdmwuxKo1/4L4dHNCSVi7oUnMP1WKkeF2y7RXJfNNqxERojW6AE1
Zt3YYWNtSn39qKVQI/YP5dzRCb0T1pNzIvdHt/nZnuwu0GGOxYNz4yEKUSEGcnCcC+rEw/TCmrnV
MHsvwJoVtS++M7jeKO4tyrlyVtpK4NwtJd/sYWPeaCzcKZNLW1CR6Lx6EvemH+za9AOR6023aTJ/
quZuE+rp4iJs1hMrED/NCJ4/b4lK4pmMAzhmcGDEW5Jk/y6DD2er+d5HudbIVu+rsdsGussGhpaU
pSKuqiMaJ6/c5mrIDtBx93OoiGYZwVw4POsb+H7UkABoLmwxSqXAY/1tbQoqdAHd9fr5+2RF9E2O
p7RKup+/henqRL+8vdZsY9E8Yw6JEHJ3eOUFBnwOv2eIP6uz35iLsCuj3yx9Qq4TK9KEbvGbfS1w
FdGc9yJhM8J1UrwNYCH4vTxzhjYhWVsEZuTyDtJ7ssdaVVgW0UtcQ09C3nmXjRmLawvtsoi5HZEP
2M+9U0D/1SpW1IAcHd04iCUIav+UhKATAV4yjDbUjfuynzJafKn4x9GQV8OttcbEXsWvyNUS9cI0
A6xUqGZdJmZPVjrLK6SvFbJbgOg+fEuUt7VUnA4RlAHpSKQywlq3gd4SvQR53fYWhSoJGuloLUBF
tMaFxxAImlTlpJ+NizvhtnUKqqaiil9mBA23/BVlbfWdhzggVTHm2tT/AkrVSRjZ4Lbi31Om2ALg
HYp8Z/YBNj8WCs5w5YixlO4XZGsJRFCqZiBC0a9r/uN7wwTNEVAdgPUKkJ929hB1pHusDhIsqwfc
1TVBApMWU3lBORv1aUmxu7URbmjdgh58gQQDuOT+fRnAZYnx+BNNb5K6ktKDKN66N9BpNGYVJowe
SJrQ9A1ORnZ1pjaeBhgpcAhN7svYHvy0wweoTnmo8GsOA/reqyMkDn8krSWgJMHfy2orqs09wglQ
em2KfIANLk7xN5hI0m39tEnYk3HV96fUHI480lotTG2y6l5YfCvKhXGzSxUq2k3py+OKe6+llYz4
y4iCOujvgS1jrbZR6I79o7jYWVUaV3+XIaU8ZEV96AtVtB4g2mY3wsa2BHtGo1rG0p0zgPjeVw5B
/SmSVHX5Tl2C7/evcr/DU4VxLjz3HvPQpzDS9oL6e9JY+yWEtHsjDuBEWfO/GkNvS7xnbLsFHZUT
K5BobtDdFmhJPfRLnfK6QIfLSVyYwxXem0XQobQgcZ6tMUO1e1xdJn6pagcb+ca5qs95rCoUP7AC
Tr61gGz8fuNSmydW/JxpbpEb0jj2GXMMUFdEGDpuNB7CBMLGYuLPpTcrBtA7h6oXfuu7t+3tbzxG
sHKT5xBpslB43L667ldpq7yDCAyL5g9HHLBqEEcTDsvXznPNLQfUFXM82FaXscQ/n5LS41XxNBVu
W/9GTaU2fyuYtZ1JCwpwWXDjAXCViY2InPfEMzjiOilUWcYcKA84GzvPFrIhO0CDGCMkOw4u/SFO
/AWmwyqc77FyAOBj94sOFFPvkimXxKIEEI2mOCu42uXu8ta7kZcUEt9vTsAyV2qfDQP+QQMFA/Ip
SbLV+RFk5nfvTzD7afeV8kIu5rLdbD4E6ARgi0QojYJw+9cJh3RyvM51W+aCMpjS6e6UlBozldjs
TlkTuN9AG1aYMMxIJlkmTzgzo9P2PXyiv0Xngrvufc0PogbKGfItRnGu2XLK3nq3jmFwYVpKeEPD
pfUPx0OvZpxuKKgW1rAC3/aCayL4veRJ3UuWN2105v1yesjcrE3yQdnm0qU2OEqmZTAq9G/kdNV8
bog5Qgd8d0HZp2jlZ8UwZE9gWyVOwKfg1tk0wyLC8hWUZh0QM+b5KxX9KALXeEXz33BWM+qYhEe9
GdXUcJI2ychLeojdzhaNLi7KUKZZunaZs/WPKlSOhvZUqFMYgwLGSAg81oflUExSlIE9ZGyENSZ6
l1Vw/WHOqU2eLqrCVKDdcIIO6pm7Gvz5krtTXAFU0FaKRQwBU3W9Zg+Vcr90xPqWdHyo1utZ6VpZ
2Y9RIY9Sr5lIh0yaImlOM5xRNaXM13gMXS4RFaNazEmz538bQUOu+u6Q8U0TI3gI/c/517pvLGT9
veLsnDmSwQO1lsxd+wvd5rBGAvaeB17yrdGqjczwj2DpuQvA8ZDVkPpE50kWE1rRPYywTbmT53Va
5CGtMIdX9i8OfQ7O3i+NTKj6X2SdD+csq2a5AqBk+qHtWhUdAb6lJzMSpRUruA67gdYaN4i3J9L3
zxJhTSF76ueBwwQ7n346Yy0cRSd9I+AdtHLv4vl1/2lC2DtplHsTxfX9UWmizfdqjjJwON3Ov/cc
gzBjM4rwDssk/TTgU+ZmX7IWHHWKYQz3CrW+yk0BYgTjrx0JYeg79QSLs4uhWTKf5W+aCYujF9v6
SziFDdaMfJbpuuS3aohClSv72nB9rKK9opTzcU6vezP0eRvuPzqp36kau5q6G82TdyjKon2fUX8x
kGTTXyvfC2De14X3RypJ728QopnDPqBu6E8R0nj4i6+qFAATEn0f5lo5ruZ9InaU7/sFaX/PqOd0
PJ8socNSExwJvjXpq//33SYFzRmfKk+Mvyw9a5xxiitxxqkUBEFz3MA/qgH7QyaSRpLvUu+hzVXT
wqj+q9VfXnPpRr/N7yyT56dTK7KvxcagqPoqiqHpsnYelunhZZLpxEi1K6D2PN7V6QL+XAdP8oT6
wil/m+KDtDMr8Wza38XyYq3/KPMmRMFRk2ciAtfQ0B1G1bnRqr6D0iRJKySQBE/KNyledMfsyyWi
RY1jyl/kQYw3q2psd15A0D6ncQ4/3d5ndfILtpEbmfjsjgAMorPqpQURDQT3IUutMtdPJVW5zkbr
NPzRGbV3gd6L4pPa25cArIV5seyQbvte76X+1mCPGG3n8X9UzClex/k1dmKGkhV5IB6jyDO9FiF9
eP6zC4lDKCuMZxq/KTQoxllwmvSsPLIuOmXm8yQz70eY63CHA7cXoqildaNVP7Ihs7hoHLc/M98y
cv5a5B7P+J+pqjLp+uqkG8CClymrWlzALRDv8pHrqg5Knk+UbwJgQjNKOHP1Bg9WScalOKKO32Ne
oeuM2TIzrArDowOegUC24szXsrMwlvLV/FFrbm4yyvp9TQi3917GSYj+uJvrmDqxko3srJTx4qp0
ZxJzUssYYAxjhQJGNorY2JtTihuNxWjBpSWfvrYQJZz1dGAEw6J95k+b26zkEfdkHJCOQhgKRcNt
6WG2973LrhxY5JFrbsDse0MfMxQCReqcgkATQPTkf4sSteYZzhU1sg455bt8Rzqn2YVpLLDZfYFw
OHQxSuZ6m44p0Z1z0cFQjaQszFWQyCJPWrPvvxFk9qjdIOGAJK94/5VBw0B1Tg9NYuYo2BM2xmD8
NwXSGJ98IMkxt+IKR50oVlwkHQi46EY9k2iJ2VVS6C9HA/po71ervRSbIsf60bDKUyht6xLUj017
nOikS4zMRTvt7yId5Vmqau6nntpT/ulE+QPiJClB3KKJVT5L1TP0vewny1sP/BNp/yR5dpCydSYz
kJt7w0MHsv+9TY8bT6h8qVKnqQHwYYMP0vmYemW28SpxCE9IKwtUQXdj6MX2LiQimCupNXZ/ymQI
WmXQ5e3mgEMGSfMbJySTt/EiMlSifi8UwsvDM0B1fSJS2WD256tXKsyAC88wEEnS2hpf514fD0mD
8f5vCAQrPQdUsP08VLbfgYgDUQPbHwFT0SGJ2/MZQ8qSsZ9Dx9KyCaRMLNwCYAe0SH6tg1mTMtNb
XBv+lwLlLjZ+YSkun9uPLir1mDGIe2xwnrv6Ff0BVmvPK9Ca6/KN4EFS5SX1l72SsqFYoZxhTBiu
+JI1aKqfV5QJn8dvb1IevSc4/TxjAslmu30XrQjQVir72C+JthrbD8vWG7t5YEUszn13ht1UseiD
4rFzcBOao3rxsc0cZGIxrWLixnP3+Kh0MerNBq3xEsXZMBgcTFeH0m9AWEngI+y52iMOyJthm6C+
WNXmzQXSzLg5KhPt5E2SybIeI71uoUUIuqdJPMFoHerBUW95//K3HBPPqH8X5MkcS8kWpHB3DVRG
7PWyOBRlxShy0EHfEM4iGc2X9LRGervkNzdjTnDh3ayqXz7fjMX5S68EZ0+xQVNYo5u2AZ6qJZ5i
meko2FeJDjjwczxJtznhShb+7KfZ1T+5KKii7NtU8j1nATwyX8sfOfHoxOPFsfRN0Em/s1mCwOpF
MQSbC1XmuPBcVSVlFLziEJbkczA7BMN6qNy8Zd1Hd2QeP4ykmfOkWpxOK+7fJwgCsoBjqCUVIxd1
GFI9+ZKOjVRFtB2PfwmFvcF0FmHqKQ5KoN6C2xSqUkHXSICCPCil3a7lh1FbyBgNmCqaHt3zBgiu
LKNxMtjWf7mjQj0mj8Ly8u1gBuAC51zLgqikCneqOi/XWD7YtZZzMLutYwEOFceIAcEWCn0ojxXv
7KP+ku00ZpBfLxcKM9IIoyJRRJTyuprGsgH28deP6Exekq0l1jYh55stN7/U3KJf7fMlvgi95TKW
yWkFdNzMzG0emk1wKVRdKXUN2ITP3tEKJhBA5KHspMAlEu8E/3OtxXIi2TE6ulNPLasC7MiWV9Vh
CfjQUKK487CymDvS5dR14XgPRfLs2UdkoXujocnxULTBLGft9z4WodBrme5/uFYCBCRr//wjeosL
1r+86A1ej+WMOc2R70ztUWrDkcuqxDDaVvxegBuTSPdslUQL91FBpQTVIKWegAJh2m01DHEDqYyM
UJ4bqt/MKpQ25WZBy+3CVcKVrELMz2kLW7LRvihaE71II9s7Ys357T5WBu8VD5Br1J29B/CgHTzC
3tpgxgwR8s6v8C6JINYPGBMP/7q+je+2w5F7cpvYrNkdGqE7f41sEwyWqyreKNW+u5CoLI5SeX//
mkx+h4A9+3XPp90/XtrrF1FfCtabd6fI9tjjlytM4hPzkClSlanqyy2nlJ6UfV7RLTMSErE4knbF
QMOxHN7cr+6TOTOr5fSQxyeZ8IdLB+eEOTAvGVoSz/rQs7DmroFR5GWGaRwdWtE1lz3ryAGMAePi
krFHxkqxFf2HrhxQkvENS63OtNGp2RRfkatABcsoexykWQhDIO3MB9J2HqqBXlzdQ6PazCcMLkjB
NM19D9Z0ZwzCczQGzppnlbyhf9JD50N9h988ZOrkb3r4ipq84BzwuV4H7dDA1+r4VA1XtlEL+QnF
y7+eUHklXTZJDoRo5WNg5s7UF4/VCCDy6P+wNSj7QanBSn2U16FaSvXvPbFgpOoyGmhjJAaEnmpA
yQEVhU/+6eYoUP1CbGqPrEcxOaA/EvAPpv/PmycavmYoF22VmJeltdlDW8YTh8Yd4nflpTV8/dTq
MwE952hYSiv0VrYR0872STf9X0/Cl717UxVtpI2NtwNlVImwNoCX4t7GqJd8xsrn2QCo4KRYi/3Z
Z1vFGz35EMo6j6tqkmFIXSEcd8xiqJFr4CDROMy4mwwmOY3PQL8/qoXjJXokAjt/rXXVr5ykw3lW
R+k0RyyK0PynWL8yxkfYdNY19aQWZSiG4PmhrLeEbNQ64e+NNVRzDyc2TfYLd6RngRtLBXbRAF4/
O6IekrdTVmEHbU2W7ykMR6QbArQv5+VfhfgP9wHWYfzT4PvbmEEi4lC5yNbOGsjjJNoGzr7Srtfk
wW7dKCeu+oNQsJMDxp/TlCi6cJNPnrtKY8CioNV5gDLufYf6LRAux4c34WnnNiv9FvH1uFhoKQ/u
fDBVBocbyyWFOli2j7+qCfoEcsnz94IfJJE+9GDzi9+rN/00OTXKoZUSsChNdAFYM5aYvwm0U0Nz
lImQtA5qGK1H3fbBYL0PtVdQqemYREM7jYBV9qMBdBJqgsP8bTdBhX4UjHRipAOEcXs4k8ycyPfU
DnzE3Cx5MlIFA93TN/PnniK0FJh/jNcxyLmGkmGWhnqpOkPaDGMMdMnzyCfirEXzN1bMlvBmtQyo
B/Z0l3JW9hvT42mZF0u779FztV8Go+ajgOLBOG+YFKiiYjqrEZTZkqsV6y+bVELz4rHVCVCZXx93
BrhsHcWdJKTYKWGVSbywpEz0YuqGRd8g7bHCCrC4cN0GgM+NbEM1IQjnJ88SCgfupLqR+faXWbgB
kaX3TdMrS6dyOoEZrHmaaEeESUeVb1exObkMSpoJwetnBi2d/4W9HeMBMRwtYOfN6iqxJbqtCwIW
EnWxOF/d+u1ZNqqgq5eN05/IIS1teQMmmRAin5qjH+wbo/i3Hno4ogzcczodi+4fgnXG/uY/X9Nv
1zFIf2pxqV8n6OQoFJ9DS4gBl+OhQIZRYD4nBU+1i+U4TvpZ8GEqJH6Yk+aqOlJtnLEaK7RSp4nI
cjkfUQGjc7a+eJD1bois6YdrEzMWLOPXyTtvbOaZIoC9ry+C7Kbz2ujgG14Ch3dgHKj55/JziRg8
Y/aeuoIltnAysZ7lJwQ3lQGsn4OEVWmhLD9a+VD3hhVNAHNv3IMu2RtmIVf5iNHxzwS+Moqpdtfc
NnohCBfvnMQlJkua1f689Tdj8z6Hq5nQfXzZi7ab2zJJSrE5g/VEjIr7hCVr1f08ZptJyteT7jrT
y/iWDdB6OBXZug+sdWmRfINcqZcpPXWHVx5ZC5uJedOxYmzu5TXMfK1/y85X0PPTUgbegZjGlvXm
rRYHSYECW7zugR55LHDvDjygQIuR/b1pPq6DdH5j43LyjhidqFMCau+mIrZyZ5GH3i2KxLshaA0E
ThHikEMtUBWFzrjNtOWF58MnTEkRbXTZRjDuRQuzsjpE7fKxc77gOVeUC6LSs/PQDQf+BCh8pxW0
DsISmfIZxR77Iag5+Tm/ZmsKYHm4mo2du5Y6S8jcesODivIHcA4iP0jF5gtSAkqQebbOqAk9hV1j
+XndXLsa3a4qeS3GDE17ACbOJF9ubP/dL9L7tiXwu4/GYJEjEzzyRDUDFS/MzGa+WEHGFSnV0BkV
X4+II43bTSonzvZKDKVThyf4xLCimCj9brbYNubnL5idRIps7dExct3dL2092L/HoRE9oAt+erfA
wGiGseAyP8JeRa1oqKnSI83Y7H64KRdqk1IIdxCR0sWk5JvsDlT0BCOaHWKUy5Y+aDo3dLEMv3Kt
npXXgi5KfJkvhP+YhyLe5gi3mZyDUhS+U50LPYzW5c8lXM4VBCmzWMcwQqiXQCg2R0OH2tRHMLZ1
R3qDiz6avnA/sQIEb/IEcWbyLmzypbywOOOuEPZzrhj5opibopjwQibwUEnpBQopkG9EO/XU7Q8Z
glYCrIHyIup8+D9O/3EXGfKTYfK+MaxAqKUZryv53SGHnQ3I8oidRmgI2z/S4mzhJBfz0ztT1FFh
iBp2t6r+Wd/6I7SYK+0Rsz3KJY+kDkU60HdokaA5sGbgmeCm7dmc+ke7Ql5Jykfqbs1XgUI4A064
fb6SArvgr+BXBJeo+uEZv0Tu938Yr8rmztVDzsn49ZKrlfrSS9Au6pO6CU5fDeK1cciIVP5xRJMR
4FG/Jr0A1VY7ZIGOFclXVpuVYiSvuWFvFPcioefTkzNSS0+jgHsrcTHfSOyA5lYB5ebMm4u5d2/B
trVfWfUF+yLAtFIZt4Knp8mm5pASB9GfCAtAn/4lagmai5I1OCM8d+AyI0wyYYsVhBPxarj/oEn8
4zMjaNgdh50UoIME3I4DkzcvyjMu/sFKXmK4KpVdOcrweRaeifcxNk0gB/9rTshNhf0KZOT1T2Td
pQHwDyn3xM+qhH/znGX5SQVBp6uS6ZtSwWC4ZW9cfNkJZXpqde+5AOFo17Yzx/rI+t6MG0qHhYCF
VBZfwxu06Hz+jMxQzvgvtqHIbWyMHMFWRWY/gngkRJvxyzZMKfQkQ/IxexAsVepc24VdShAtCJDU
RyHTFpjCUAR/GEFYyvdQ9oB5QWhQg0RA05kpDDEJR52qaMu1u3U+9xF4UNBDF1ZdccUS+0vrlzUC
HczEiC7oevzmQxoEuUP04dJM0wP6vsdmdqSIz4oo0CbFXTZb70UaDppTkE1R1MNz7d6bSPGOxMR+
9R+FuYTsNF7jr2vX4uSFuXEpuIfFmrzBJqWQ8RoNbbUlmiJfbmFput1UAXKycoVxw1jzi07tW/6N
VXl2jl9PsEkWaUzug1qaI5y3Lll07au15nWTDtSMrpk8NPBtsNYEbvtFOHZT3UIhxrv5zHFMbYs1
T9jxnw+DKmxv7Th05iyUHsFYAVq3DKyda8ktwz+RJykK0wZkGV7hlUyS9jSIpuV9n/NsrTnJoYHo
RIXMyL3Y8lPMh6sdtyK0HM11ZqOs9FKoRGacDfxHH6MFRHazUfMvFzncyOGFsU82Eay5BEfn9eDQ
C2y5ivYt/daBUzAWPAnix8S7rZKAnFAimnJiKOafMK9BHJ9OCCwOYW5hnc2dWU2rPVnKwWhb/nPz
ADN/qwEj1CITu0uRtQqvPxvrlDdKP0dd8bZIWtfT7Kw8veF5Mz6k9L0LTbZNP3RUeT+uAvjAkLBp
EHUtwT1DYsxmpr7So3kUwQEu6yP5XYG8tcMkIZBS2aFTLy5xdnWrbuLALSZ2WqB1RcWMiZeC45D1
7YkkdHWh2ZAf2XupgQzyvDYM1f5PzIiTVz0/Q5i498eiWwFu101lfT18lipnUMPmPROR2c9OmPf+
pGwBYIIc+ufp9EAnE5dorumpo8bdbHGLRQICrHUUlbZCNmGCnbqCV3xW7lqdkznln+GmIt7hnbu5
97I/rEyBU95CW9ha8keU8Gw/mQdkXci1AWlR1JZXjUqFiP1dj/gck8xWRQ6wB78xWqf8MwadrKrY
e5RCkV3ruzMLGrd6Ahmh2xtXkw85Rsl3eT7FawI64oylK1//S0XbBnV+Xg+BV1Owkgdm7UG870Wj
JwHbnnuJttk1pRVo9IS83wIvOosXChxWg1FhurQDPl9RT6cNpo+OXqsWl/uLYs3YXdEVLYb/VfMN
XbULBwm8O5Tw2615lNpckKtwSpSAgYLgIoXgeEVRNkKHmA3+lALRnUNfkfXO67UQJRjCnkDPtumw
BhTTxet0JBFpR9yiWyK+BTVWDwx51t5j2/C2aD7nnSdGWErjyLUtF7PCptQ3OjcdczwRKbzsGt0E
PLtp9yElPgQ4iye1+zDCzJ8RqHdYFVvH9Ll8BQs20wz/V5bh3aCdIVO62GUVxZdCYvh1Xsl6J/F+
MmToezEGxVAYWFaCGgykcc4ekuszKte3kCex9qi/aq9dT/fd8hEpY2N1UKrrPPIq3wD6b0D62CQN
z5I42gnML76Jn913NUn4bVaWYKvB0+2pjho9yp1zmFJLmBSx2E5/pTXwAaBmBvLT0tG7EJq4/dm4
cfXtGCevPrIrb0NkJb0/TKqJlCEkRJJOBGKyT/+SAWQMQspwd17YNNuIhX8W3syt6ml3LMeOV81p
OYyVmPUPEujSu9Jx+GjBUOQH7JF8HfaCaPfoRUi1iSzz2goMz3GUpNhljw/AVQYg39MomigxbH23
aDE94/aHr5AkyOaMf7Tq5/XbfhbF/7azTpGLzZptMgVWO5DzwDfZLWZ9n1lA/CFlaH4m1FqUaIkE
GeliesIBI5W9uS+3I+BjjKO3zZ/Qoaco+eEwc1ayvJXk4MG8PJcc8bRSEifQzV78wgios6/+MGcw
fr9T0pcMRv1MgyLd4oTxFvaaeVT/NcmNom5ZjOxg92Qmg2+5aIB4e5u+K6eMwwc9VmTLsrqi9QHZ
VpMpngEBFebh63bQBfQY6+WxXrk/6CrUpNaMGuS6uiPRNMqaR0+zpxKPyIolGKujA5Cqb/fDs4/O
XRfwJo9U3yp74KWf72vjtQW68YvHspnyUu+kz+HOq53g6q1K5AHypmxUm7qN8AN8pA87+M7nkpOl
gO3xD7xWgXrMrgzppyWa1uDKoJn6FnqLG8efOtHjSn+VVj4EOfqO7TnGWju/ZL9PtCBPZC5iev5k
kdmIWNxCrlbwZvkkbYq6HinTx2+Leo7Auh0JlbnezD60SSWmrpcpenez/Z2TbAICSdddOW11ffmj
VYsFTJvb1bid2EbZxMiNCjG957E0Ld+5MD3B6MOxjvcDjcCW/NGZT0K2eZ2m72gDFynkfc2mi9c5
9JgWhe2OBvdOsDVW+abWtKDcr6PXz8v4IMJftoZIj3Ee39g2gVMhrRL6EXjzshPID9h3VMLQ86dJ
0i6ljChaU1c0sQ5vRw8bjrG5Js6fM9aTnJNwvGhxYFsL/0LQ40rppS2GPCHvswXqf48rfuKuAFeU
i3HKssu8IFninLGEvjjXpPjV1gSM43YjiwlO0vjiEHHNHQo/vtTp5i4Ez08KdJLwgGP16mSiAEVM
kVeb6Zyj4c+lIXfNcb/lIesBadPf+YX/HhNJmPzxvO1zNxf/hUYRDWzRyeCyHJlewdOVrDXkmunJ
q6+yPj0Sq3PpN9WCTPsPOclEZOp6qSE+ScG4R4U4WWuCvHBBbPE78Qcoji3j+xt86ftmRgFCt4zV
QgpCNXxAz1sr/funI7iDyVAqP7z58BLaDKd5MKvfUS0rlnJXRLJOHzZpTVEmbnqgQcBOEYX0Fjjz
32AUcrnz1V12I4sspHwCuAcuMW/3eteGpRi6579gqqtmNgcBAM6YppLPUP/tSZPLDv1a2pFOomj7
XEeHLdLgQSHU3l/0MifGrYllqZJ7rRfybbiS/DPBjB1m59KZ3Z7D5wykST6kaMDmYpThlHa0hRmK
v2ONBXiJG/lSqnw/4tQ96vNCbtFOW/P9csn2TSnde9zK5f7jkLEw3+LXU2u302MVMtwmpP7YuA53
7ID0YYt7JtjIqWnAL0gRP7CYtrgj3dCONZGv7WN8E4LkD8o6tYKuK3OYVfz3AKMuxISS7SylPHlY
gHu6HWftJt24/CI/hziLZnlm0C7pIvNpkB6vO08YfqpdzAMDHPGriyv7LXwWjYN3P+HrPJScTGBf
CFejits4WNj/IWZGT+8pLnCMY+vdAD9Uat6peLw4PNKux3FcOgHhfB+bBJzGf1nZL6oR6vJrDtDI
+s6rNjvgj1oRKUpobG3NgkqpWurGxW8BTVFW7OO/xTibG1A3kjckCWvNEjuOAE6Acb8lMB21yOPF
txpTzU/wkJMPw5prA5gdkXY6CsWETUPgLrTwN2ysDEEDLOg9s4WGGzf0159KI6wuXlCzyldYPc98
fWe8imVmMCvXbCmJgpqp6kczqq0Jvj1oXu4E43mu17bgDhraKFdgqyt3fUP0xfbhWOAy2ZPcM7lE
fmvjqHcBrcH9e9XByBCN/mSzbPmS5/acRUfE8UuMIs2FB60ZPxQwUkD9Cd597MzV21/aoagI5c0S
2JBQG3xiaZ9IMxcFfUW4eacvAOgfnUBZX56JDCCrOzkNfoHbZEC2uMfK8oW8B4f2VWSgUOA97nEK
8qmG8hQFuYeOBrCFsXSGBSL5Gjz9bYwp5I9fCl8crDe/d4tDUNlo1lckJe25pbTRx/rJsPgmi0Eo
LSaC4JOqqMisg5vstSLfXi0OgiNzq0CdVfayI7LB0sNkUZeWnUjrTJdL2ATJskWcdIBHHDG97u+s
5iFNZgyJ61q46fQZJTuQunZsQ1PaydEJaOpHuuZ5NMACubLsbMbWwyiqqfIJAPYC3mOLKqVtYad2
3e94+ZyEdqH11ZHRUoBerJm/FSdqJk2wYIvklSox0QTVouhLwF9R+Xx/qC58bOxwBOv8rPRLpky0
R3leJTNVkx6oMijnNQEF4XJpWfe4YuKgu7K5ACOxKkmzRh0t4pHSTc+PlZtuhfTIjPYy7Nc9v1gk
4t0tDc33hZv5G1R8f0VL6tqhgJLxMVCYBsalhjfs0/BWt0B54WfsusY7brYcqRewN3cwpqfWzYNQ
oE5s9wgutybqin5DFLs9vb4qvQjNMxYnm8CRd/aXinF+qqvq1PdRVOq0+6nJqcpIuawvAti8RYbP
q6qc8QEdInyPg1aHHdcB7p0mxbU7s4ObBjz51yyAyfLx8oKfYHsMlNBkHb74ZqBLmiLSoDl/g6gJ
XyVVXe74CWu4gZJ1tfQKAe0bQGKSjEJwANDdxqNGSZtwhlBDdjuJ3/7WqaV0bVg/8WYQlNyd+jn9
FHNLySltQk/fYISFJcTfikqu8eIj5JDLq+IRdgjJJgqf1vaNco4pSIPSOmMDG4QPL7bTuWGloDub
9xcsWHdPjp/EhYrGY0Kh3r+2z2/iGI/N20dQMyWEatlqZ2I0lsyrUJqq5HghrwUqHECEk8AMAdrm
VZvGFuCU9Ruohyiv6YR1/nCJoywQbmZMeyPrLrfKOVu6YfUVjsHFTSH4JQCiZQsxTGzozRC6UHqg
86UMKyoIN843Ncui2RHz0w5in7OP4efFD0Flr1i2gpvan3hWs6j6t/uzc46e7Fg5SZIwizi44w0G
riRkugo+DRSX8Nyrx4NMoWW/VIZRrdmwRc9/GJQBLkazJpfBuG/7mJ4idnKshcA7OiX/LAszIIQs
exLGdxdQPzPDanlWsNjaA9p6AvF5A8Bu6b0CdT1B3Sn9fkReDjHDe8unYa1k2l1fmTTMdsgAr9Vq
VFkNtQoS0EcSF84e3v39SvL75BLC2mSzbA4t5r+H4yF+7wWPdGniCIR3n4DxktVbLO01FLRG90qF
j4SfRixeCmb0oxfxNv1lEQ3KTDg2dVO0tDmImdm01TfSo/qr9Cx4PgelSO/82adiJD2wg/ZskEXR
pJp1o+TfATaZ1TOi5RbgQShUt8sR5wOxc1g5DdeFOXe20vkufApbJ1vIQVzaS7OzV50vCibFQbZf
H4LWDm5n8IlkaLreJmyCvdnHP6vvUsjpJvMzM1fN06bhkQaRd7ug23TuJF82NAoW3kmKKUI2Qy6l
4UNfpwDCKDQIji005ZkYs+jVzKiteCFcgk3NVdWk2nYE1Clj8REW2N8EAmMF6kOJDjGrL2yY4LdD
qJsPh27w46vqLXX56N7RGaFIYMtHqJ0/CLUw34BjLX225ssryp1pFPy5gIAB/taEXenfTv5r0qmK
7O7tsAVnL6VSB+QJhtKNGhFIBLVDW9/o6/JwlIbIW9xigu0RLXpYtA5jHZAGf0QtEpBJQ+7Co2YF
e1McRri4L2d4E5feHqFDKywQUVDEtM6fgn+LSNaRCHs8+szpZ6MVGkWINBVLImMJUzcwRoUXYJ4Q
E6BzrBSrwuE12jaeCGKvQI6O+R8ovrVPsiiHh2pvSUxiQ8moetlBiHJY5ob3w5rFtxu9C+XPbhto
vw36/GqQZQ32Clr791qh8065xK/Zj9q5rg9027r1c71l3Il2XWyz1WZjphaPu384pDUH2HGkUb/N
lCLtACb/+eLKoGVG2xlHArMSHn4vi/urHpmdwywfp+N/6aPldsQ4i8RWoUHZ/3cYVfCGkv96s5ez
KFKxWFeM+LfjOR/5gzbUsmXDtJIo8w8pC9+FZyiuZ1gPH2VLZc3eFwPsbpIClF3XDk3f4b2yxfUZ
n+W69c8H96PIfJJPv0r3wB93hnCH+fnipJFKJhC+M+DToXmmt4dXl7iyqUDtg/fneAeKflQoxuiS
lz+qe09A3flCNy1u929wtx1sTjpdzRutA9+cK+ZgQkDPMQt2CikMHOWa0ONyfbm4oyxI9j2eA2j4
az7fmnpCWDawm9nM2h2bKmlAZ01ngUX7Non8DtZkhNMevg66HKv48GACcMAAIEyTAwKxjhgNBlj5
SAhZLsUa/ugo+NDw+XlDz63ruhwGyMUera7/DWA0RWEaPsdefdoWNcQsc7RGXNOz+gtxIwNUOkg/
85vek78RkZIJpBBMG/0/3sXNNqaZqAL7OSaE/mH2szXxOayjE768+lbF9xTwi5omyqzx2aR4m1+R
qdag5IORKRiGqhR3qBawJIpn8cR8rjMoUGhDamNX5W55w+fFnQsf5kFYdjkuVtZfOMzquTIcSTb4
u9qX7XQ8u61I9IT/xUPJS94U+NfUX8eJeL/gTFJzeucq+83VKWlj6i5rfM/Vu9Hmye3VviyjaddP
+uIfh3NJjadP9qQwPok+jXu+DXvWrOfV28Y/OhszG5KQkHJ7GejPze5/2sDEKRdMVhiEeYe+2SDX
1c9+nmXa7HglIFu6t2BTmnYTEP6NlSgcATDs/TlQ3aAKlCUwUrlCP/As/qWq5yD9AvkF1s03j9BU
KI1fR2FFncT8bAdg6uCDhqfKYNsQ89uPd3zp6ZxVvl3/q+ylbGcna29lzCx8oOOhvsXzjGXajJ5W
7Bmw0PkGUl8bYvMwsm1rDdHTN9OgiSJxbyUwczwqs0YTB4MAAOFqsfEXM1JMJr+XeIWPZ3oXcJ7E
myQSQqnmqkWiSakVIJlmFmVartTMSpswpWiFV9sl2jThORwi1+HsD0K+eYlkkfcjK7Ac/FBSaWba
IodSAcDhZc/N+PKDtrpLEjqta8z6OC2MYrfZcsHyJ4kaXvVVOq0zao7C7jHU9ylHGxiOTaSEJGvq
GhALJ4+L6ueaFIFGk8ZqLyJZYg3p1FENDgVZgDFjPP6pHXcAC3agiqAzxbWndgaaEgZILkKHK4/L
q2c1v7Xsxb7Zmsg+HVbtOnhvXFUAoQi8gz8ppQL/fp3sfcvUNTdoVBwoot9idhz6pWXY8dWNh9Jv
hhwXP9XZlqW6GzkB6xzPelqs3ADoFkPcVZZZlndyqjmxECQlGvgOzVvY9TOUVPYXVI21to5glhtI
3pNwpu7yztF5slXdY+wemw1peF/s7yvhWwWT7kxHjnzTmhSCjN/WIjsGFOvQLe60rMz0D9YZQkwc
lUkoynBjbzhP3dt2TGZfWrmNTVLDgDnk9+EC6WF07ABTZVnPvCxIwijuxrDYAtGXjZuk/JBzUNGD
lGoQQyon3rzpkNEdsIBtSrbG9psvK4fiH+uA3sZ5Do9onMebfWakqyfQ93tZWofgwe3zCB0hiy7W
K1/uMqFUuB5BJjt3uXYZdD+83kJcQ+e4UCc5pfKBh8Ga0vaMA5ZcgdQPRoT/8rsa7VtfF9dUhsLO
Kq0Ovy+Z9gdqY84UBo3Y3+Jt16eyjmmLEfSLcKQxsIgtgR700KvHHsjFsG5+8Cjj464asNH+SGYk
Tp7Z8ir2XR2PvddMpLZHc+hp86lt9XQT3j1OIZMHfIkN6RJmIBcHDhl2HsQ5ss7ztuI9JsZsKgAF
8Ec2K3/4tvsDI/xWj/wDxgAudVnJMbi9hVQm8PiLfCdg2Z0XRtBi9qifpXINiM3UdyNMYxWydWee
nKACDcq0J3IvM9weD4IGNrQObLKBfke0nzQS/JSkCSV7H2r6Jmuf6Xa39qJDK5EivDMyQ2fQfl1M
FiMCyhe88BP0yWSBL7tLa/NDDmikB7ywkaV2uqVSDEvh7U3Yw66Llo3E+fqK7kkKhLIiwP1WgRWQ
/rRziG0s7aCGBAkWIrPV04ONMCxwlkG43UbbRYJOyTIA4ywhBu/GVNZzyX1Y1qURZZ/PFOoCh5LZ
qc5FdnEvuO7aRAE48JK6SKkgQgNWg1lExB7+kf+3CROtpV+ci3DHD028h+ZJ0tHEHGMIRyTf4Bx5
Nia2IbRi1X4VHIupuMbYMv2oMs6i14iY1+z+qrjHR8Z5uWWTnfS4rNngPJHE811E/mMDFthG9UH9
KWUw/S1CmLljC7IkA+342Gr/t+OmwZ3bQ/NRrNvHV58VbW4LaLqgX1ZOFhWxjZOEad+cZpCjAE1Z
tm2CCFsp4p4GKo2sp95jC9uD/d8ZXX3PqcRlvPjxZmFtLRT57eDzsKK4g1z3g3Hu/sw8Tx2/ywpY
QhGFyb0Cb6tsj2e8I4uBSAndXo6kRvOxB2qWziofX4t1Bb0uufAe+0/y4R1mPYTHoJs3qBGuTugp
XgY4MWHSZhyZ/bmpg5ZGv7sOYHNpRSz80cY6KLC0+JoLEX9MGUA/vZNs0o3kV53EJX3H4O2tW3O8
/3nWo/nT7n2fhJVmsG8q6hDvl2B7t8Pkkc0wN1fOe06sqVWDT2I7uAdiwQhSw6g3onqPNuelmZ8E
LNuKLnJG0iwozbz3uYvpHeCdEiH6PZh8qUBb4r6d2f2mtBT0jboF11kDeeOyIgA8oNPAlVhj+bgp
C/uQXamXv9AWsn7pPMxj5EUDToQ22cYdHSIcCgpa6KnrQuOeQ1Mrz05Ce6aDRB187As33stsNfNS
ZLGDJ9uLiXjHdvu1bzNzwwrO/tlmDotB+TWd2ZTz06Q37EkBBQ4cVnn5Uq3SJDsWl5gXTW2uZnYT
7US+OUKbyMp+0ZBCGot+xjy5DMUR1+ngaTaYc2SLJF7OIkBZ46u7uSwu9xt6VWsCedbSnGLZA4Y7
zl2knHMdwq93LDpkKD+f3FVzguyxjbr0WDImZtarZCqQAaiftwBKXRcR6M17tNQMTj62A/w4G6Nt
Kdik2zfG1bTUUeZSOowhQuj0PIIU+xxyFEKq8qVmomSbb4YHCl1uV/7oPe5Saoe90TOZk+fR94U6
tyear8G4Sk6FZAFIHVw6mA75fwHyaqE49GPVfn5zbi6krxJe04ghXXyQ8lJAHEEhpa6tYittVHkt
UANkes8FwddJ9jS7Q4i+zmUOK5Oui8ZVm46d+qO71Ds1i+E4JutOjakkY93nMCj39rvUpWPbc+i1
410t82TSq9wJM+9/XFyEwyA4aDiN6H7JZlV6uVQJQVL9gEVcyMU3O3QJXaMvmMBsJxqH26lqCx2S
+QOrfL5blV9QNxM/M0Ne5N2fscg12n2m43iJhVvfHcK22aXtQ/Nt0jeQd3QfxId4ON2/N3z/Q2/Z
j9jAyROuOma0YF+qiL/Te9WY/5FQPmG1YBjVqKhANYLXrpeuowt6MZ6NtshVTO2mVn3FQF1jhusi
ubBeBGLMccTdFO1/qNnUBm5oY9/2Gi9Z9LRDfrMVppnfQzALAmtptUtJUHKLLSj2H4QG2/37bwHC
gx5uEwS8S8ylSrKBXoE7Kv+ZLdcFKeaDPv03KljWVlhzqKjGPMyq80xVEXAUIbykplQyPcUIYqcr
TIW9yJJEKNgUs6f2rQ8QnZFILGBwf1HfZrVYthjtcdmUbQMKx/NJ0UpJN+9T5A5METvybEXGYiEj
O5IH0+NuEFgCtIGDEOlk0rgipM2XpuiKGn8c1bC7jY/5Anl/RzJFkVRbYrC9qV2+j4l2dSc3Xm3H
FiFwe6ijJ676eJP0LgRCALe2JE6yZ4si3I0Q2xkxlVdbW6nPDYSJitaKPCkXsqcErO/WmDicga5A
kcDwuuz9bhqORkV5Opgdt7XS7/8WE2O1NRvyyf52CkwuGLH5CAAq6+d23zSav+ZHYj9zCGxonXul
PFKDZ29qcnav3G/yqRIf/rI7mjuht/m4Z8DLudtt49Qhvu85UZJertiT3VHnJOh6D00TUU7t+Sy8
/PncLBqTWzGvxC4axDlwVJiggIjKJgnBQcaX1/SQoG0w5BDjmnLnnPHgNRhV/ZogafvwHpbwy7TG
HGOFTqS4OA7vJgteIisBrvFpuAUeZR0e6QV5173btn7u+NTlaq46Hw4QinFhGb3KvmHRNDMYanVm
SalWChC0JJpCTOtpo/9DE8eG8cDk3NDOjkHTOIJKq+Olyh/ANM6ihSHfSDPBFTnaaVfQ+W13Wnzo
mZjfBIwodjT7oUM9InsLzWDhRN2kR/I3h5/rfHvpT1+fEORd3+xHtPwWzGDfklZi4umP6afCjlKN
Gnml6TtHR5hu20Fk8nV7KORuWEypKixiAJXuJoyjfdNEzzLJBPEF9UpDjZXRTVmbsXBC3Ku0Sv7B
pr6MxvvZNqEWv6nqU0o8X3I4Yhf03zpVuzoRFqncKB8Dj8o4Uy/22Lr2fbv9D4uC+/QTuF3pNQai
JpIJcarz7BtD1QKwSDIy/de9FD0yT45NVgFuaNMoV8TKhl8onvEzAwl1nZ7Pa3Yj9k+/d9WMmAvZ
0Mr195SAadUfTO1Q+M8Ong+cDR0JHgFiby3BnI/WT5rd62Q0BMTd6k6OGIyrnHRUltBr65OgYCtS
Xd645XlxwMMTSjCeSUAmg3TZG1usFnLg/35Fvaww1p7iXi+GXt/5Wyr2gCdbZyy67CvC1gb3K+FX
Oy36IBZwGfBSIPrzmNc1dInXzArAWkutYnSBxr/Sal1EhJbfGtbbNufNfF+dimQ9mFVayQbV/UPc
oo7VoTTMyicrDRwbk+8okjnv/slEfjy4c8ZJ4V7QhR3o6BuLD41OsJu8d8pOhsuhwuziPFRNRVE4
tHVHIBEYXQmJtiIR9Uz8CqkHSYfjgUinYk5bmkLNbGM3CV0WSUKRBlA+Q2kemOp6jldcGBH1blVw
ayy5P+G5OaKjLYvW1qLLNceWppBJ8r4v6p6htaqfBT8KDmA4sD9gPJ9+PpRC1v8KjatrV/akLdvq
bCR8y+bW9tutxcGlUe0cFpHvRme714aIQ2aokQvoO9LWFZHVaTmkhZeUukVHAH72GwV9oZJnsYbi
vGCE0UiX/N8Kgt7SAeDuQGnw6YNOZ2Y1DUDB+Yag2Guzifpds8qa5PVK1TyXe5mUGbZnT9oBBZCd
/VRS+14G8/ihg1IjdMcU8EuV/DWyQMdqIRBXG7ToPF353sY1i4+ls73IU0ImpLvFvW94lAe/5V5R
heEsvN29xozBAc4JyGA80fTN7szcnI7X7psKoNw4fsVz9kwUGl9wXOakIDUpU0guqTyU1FF6+Ox1
ULUxM0FgBJjQG7SIvqz+fpfn2godHHMOwIvYERBhTnMo/d+3WUGigzT/VeGsPvTPLnTj4HsolFGu
UV5+cxC/SdnbVx2rNNghd4oegXvj7rKSnXStPcSFFxirIk3Jx6fqrQrV2LUBmGqPg/WIzdqtatw2
9eWRs+GUxnc69ofA1SRAtVgFBCgEQA8W7yQw6NFQYKHMNQsxqHFWiY+2DmQ3nd4LjHkx5bXGo0kZ
uBze5rxeSo7naOKsM/nORhnW5WSCZv9MpaFKGccLv3hIEYifyg25ETJm/RZLdcIU5wOqm4aEYx1R
rA9We1Thet/NNih6tXCcXoRthddgWZlSwpp9HILMxOmBTafZdLxL8bXJxw5iYP6IE9G6DvmkgnE/
sB2wtoIm2z/NsHijZOwa6XsTDDjyGNorLT0GbbMbmPFhtPUFRMnyVT84VnDltQXZvF52pg0XSOHg
07En2nm2LtxapOXP4/NA4nKbudpfn+NdOAH/Efq81cXregocLLpfQKQfOWnTolOs3++IculDcMHI
aUUgyX1jIq27h5XmT/aqOAr4fLkvAGpoKS8+zw9wPIHcQiSpuuXcQ2CZOJhApeQ4ljU8vz0iqyR4
Mr+An1uDTV0sBQAV9CTgUSq3Wky/BKt37h8ipnc3xR82tNl+0aJHwM4Ro5nNh/TzczSaHxAbndda
V5U5fTNDhs6xGrx3JZ9tFiHZyS0K418imkSdkpZC2M+YCx3rIl3iS8PjyEDdNqJK9nocBPYevmmW
sSyIxb63tgwIFdpTh4Y1Jz1Nt+aTLZwxzotMunyjkZapmealmpKgf7ejOuX3I8DAZ2L7ckRTrxOL
7xGkINmljj33Bwco2jfEdKya4oEc1BpbRJmI13AlY9jSgRcOKH2jTwWCrsrdUqDdHjJSruevohA0
Z3haNwhe1ZgC1IRPU+qp0riW4lhsI9D6B+Po33LmxJI/8/s3LwuuoCrO0WZgHossC5YGZDTxgxz6
yrOyCuC6NYykO0ji7ihd/qvPKKaa2x+U24V6A2QuvZKmysbH3tWAeqj2o4vbXZVgn/zVeIOyiRDQ
TUwthQvLSvf5Lw5R18osYKXjO2nAl7YOOEMXmBZLzK9XChnARDZPqMrb8OGYB9OLS0rSgqXTYYUW
1Fdp461AvadrQQZM/JRh51Xq8SuNie5kdmx2nYWmCfEiBF8BuBZxyicWf0K3hNW/tfFv1SzbltoJ
aWXIJCGNBpOlbQ8xkMV5iyenISvrGcyHXWXBScQ/YTRLxEk96HOPrQP39+l1q1zRT8/UF8uYh/B6
d4vlFCUVCFZyGI8z+QRKBb2WI2fI6WdRmDZYCnVUK1MxlgoTSS1EtY2bODZrOZP/xazLzEHIhNVZ
vbNNwP0ZvvBuerR7pLFgZy3p40ccciOO4t9UsjegRqdPdIVeF9tIvv+ayrKF579Dr9sNHHVeRyTz
W7oLANV1bsGUiR0D4sfxmya5d9SqwaiZn+f98evFYW4fNdBmhYtdttjspgRB8fHSIY3QfQ0FGqHu
QiNylmGErQEra/7sVkrNTrmmYdIenqb4pm0cxcbcp3eR1P9IrvL2keqHZaAjwfq8UBY6rxpIgg0g
eXFoE49r+AbxYOuC/m7KzaulMpbX7DYjtsFpzDatODv9cJ9QWfDRoI13PU/XXLAbc8jRDD3WV0RR
z1vyyRyyU+oAlr2F+qlJvnuotZ2x5os4bzU+FjALzm3abLVr/vUB0B/1gmI/0WBuBotHCNZit7lu
ddXZqgK3l0vdlsTNMc11jysk7ddFslnYHI2D4wi/uq/HPcjR/IaBNa9F9uOLhS3e6b0M2ZBb5NGt
CitSVxXzNBgidbNwF/vmp1imLGT6WKuKDZh2KUYvEzS55EcLJd39bqb5mv92MCHHj80i/Qk53cly
e/lxSJvc4nWt606FdnEwyJSTM6Sk3IXFXi8PhUhKt7TGkTvWOQ+HVOyUWAr9RP3Qq9W9wW8zmxkn
ojbUOkOjpw/Qz9BZH0a3PfpZL1PU8JfhXMI0sb7mlwQ5YlRg48G6QInnyeQJGZWlUahRisjfdi9Z
fYc9iDU+zI7jWUAiMNY3oYZGX5Z8Y15cT8J6jU7MSyehAAwH2M0qM2ilkHam7FAxLbupDTpjY2Rh
myK3ZNvxsbTte2EUL97Limi7qVFdKkwrA+yXgfVi0dGcgj+vbyS1ih4DmG0U3KrfSghJ4hxOBhq2
9bcU7LoP00xzuvFllzBFHdozASRyhzRkex3oswD6YCJ+VyFuOS2QPMpAJLwpindiJmdu0vlYTt6q
XTURuG93Rs6ny62j8mI8YqGEDiYMY4ZFmB7Yu+rglmun2siX9kZzHH8AIiOWLsIGZFuIusx+2PCC
uzoZ0e3iNCDgHHyjakwen5ig0Lzvl+p145c6Vfo/y5c+1LMBzxWcwmcPxSLxldlezSgdyBgJRIGp
rOi1Yba4x4bew3u4Hc5h3L7u70vNNYVKTsNv4Ta7iTZyoLod18SF8kt2gdS0Wmri4lqt16h6c+JG
j5cWgC6KHq12BYttjYtK8/NSRI8Ngxfc0NAi5wy5JukIwOBEUh//M6hISUldltytWHPUh8uvKaz1
s78GbdVN70hN/N3czOIO5/WIbl40yqaWyn2pyWYkVZgiVBMvchNIklkDCtZB41SLMdY0p2BZZ7Xk
HtqJReF4lQ8JilgWdr5uYDmsGgTlDTJ6M2VOt5jPSwqyyGiWrjgYFxYnS5obQM5j52EnYcuNj7lr
hbHthQBVLGvpNwkHcH6rj00t1mO+1TMfkjNQeyPFRmU3VjZzimLHAAa33bNhNM5MnzEXbZNXXWjd
DCgWPN2W5Ze4iQQ9oKjWpuPN8JDAb0+jgMb0pX7pfkz5rAtmYDhcoH9L20lTkujyOWvdodZqSpaL
wGSrVlgba+xmn1sm570PjAkh0VfMz4ZExOi7YS3lXQWsB6QN12+oS3VZgF8ocn5If7oXZddB9UAf
Dcf2IflNWUy3pZ/xGaLmjyUA63MhkCD+42jvVUrw3gg/odOQ7xBc3Wfv8FJdMHFRSdIEOf6oDBTP
jZquC3ayU5B7CmWLTiT69dxdhf3HAns9TS8fmmq/5p323oUuO/x7wSF8kzos+f2ceHut6zJCdA5B
J6kII7/VIQru+9Lip7tFLIa/skVVywdXEDiLrxt86xY76nmESKprL8PMzsS+WB6gEMNC2QUfAjr8
/Ef4LrFOBBi6FmxWN2jhL8dfaYrRIZizilbeMiXmouBiA0wtXqSX1etzvp5pxyfHRByGQcUxNK1e
5klR4lH7I/sqMbRmr8Uvvb9ggMHCPuIVY03QVfc0MG+IbQConf2uze0+orWgz1K9B59n+d1AD+2E
t+Q8XpwP/rYyR09gju4q06zK5oXtmLsJuXIIx+943uUGEKWPxBB1NdUf6QhFLSoli9S97uAOnmy/
7yqTOR9OSzRNX5ObqzlrGlmxW3u0I2nFueT9Z6gtAeJn+RYroEKjAsfzU5XQG7WeLhieu5UWfiln
R9mgz96OsTF5jvZUUm0jfjYS0Ro1jrCWAJmv+m32/0/9yME5mqutXK6g0a2ZHCoP+Ikimy+PPUg0
Prxh9eizp7WXzvG2ikNF1VmJzdrYl5svVjLZZ1MQRl2tPqj6vb6fd8RRXMboIxDb/qva5R44uxbs
+YTd5/LJu6F4lgPB44j4yrcGMZMXJLCZVktnvMmiRqe8FHyfRT10jGJdEFWWtlA5o4pPoNfqJKMT
+ErzGsfJk4M8NRzIibXBOGq1i5qORlDHDAZmCxYKhBVBY5ww0cuL8aAD8YLf3qiEfgNeT6SeUGuM
nMsiC/15Fr7Qssv5f7LU0fUmbNS42DjgpaNAb7WRmZMz/hK+wNY5MKMhlMV5FALUbysPMKbNKEXi
WCKtw3o1zojyYP6SiY9/t9TFX7Ovhp6R4bVZDiyHHUNRbbHj7mbj2YjihxXIeTb8i980pB0Gr2Iy
oS11wBnltebxinXAz4hiKEo3ajYEeE/LpdOfccYp4QXDH628pCwMYHB6PiEc/DsSesGwJnzB6Hvw
+5j5qzCSgLLhSQmTsT92/he6OPySySkA7eStMxFB071knsCO3maILdrJuqoBnS5/iFliVaJNPpqy
a+n3EaIny+7kzr6kRaMC0YGbtW0hnNy462DDHAcI+eDCRR7ouNCH0QoMDnr+uEAgrcQe7OMAI9eP
3bxxkXjBp4qDyJZlNva7RvjpDi2mSI+sq2ZDtO7ChouxE8iMjMoOOQich8kydqXqX/P1BHNfrlvC
hzNi2TyFsVH7gF+XGroC4FP84edsrL6U6STp/vJ2P8pBNY6H0lq5Tl2CcOvv8AUYrEN6CkZQoMJF
wwKn2QenmxfJHLlor4bM2Vm2Odf8i/VWCQDdRI0tGvV2cXc0ShxKTH6WkYHlNsUH3Qf4d1KejRrt
x07l5DqC4zpPqBsadozdJ+spgnd+ZyFzsq/p8G2KEDHXk7YBU6Lzgv46UstXbTgbo2FBTqiiZBqf
d3cD4g5z+kCAgNcn6BHhHyp57jBh2Dv38IerHoqzr7WxNleoqp3fJ7UT28bSk3WeNNpBldbPZgNy
WTXtg7OrD9/AizUu5WA8UsfgUeOzfCYNjQ+lkZyB8yTtfam1mxViWWEM/0TNpJIvo890adx2XYkw
31TmNDBwuy8XIZ9+EJOpKvfxvpfwn17hTE80wtcpDRGxoTzgol3+MLhSbiHxwzThcQS/UmOKrUyb
Xc2kQTG/+nM8YY9pAgEKaqR87akizG1aYGUHrPgL95r0/KtvBbSgzrCcGmLeOjtSShWUtKla1a4H
stz6HTBzfLzMZ9gFb1nat/TPRr4jflI+H6z5fmewAgJ/Qfb2FG+cisVAwuCWumr9QKPNoRDXCg8L
FVeOpaP0B9lVqblSMIicucYK//7IKGqGOkRFs42ETuAPJQERvaUmPr/IEsdbL3O8SBep/AQhMoG6
0ZSaSBnLoB6nKLXiUXOoE8YAwYMzAhhZcdg+Qg0SgRHSQzTFe8bsFeWgNiIMb4xJCEBrkYUBDj8Z
Q1am41Uou6cgeLAMv9SEB0AM1J8ICFEWukU+PaK0wqhWO6vjswd0nrBobF2a+LU6cfYbDHGFNG/F
7J+J7xD3PAdLkAghzolEpjU9GvXyL0buI/vRuhFCpaqlaTL4YiroKPGGMmaKUL8wBzbhzYtJS4iP
ocLIC+x6t5YCOnVxb1VbhWUBbWFoa2pwqcwDUzkzS8+9HcfzD20Kz9ciBQYn1taIBH8reU4PGiVP
lOpBshdwH2DgW4OlnSRquSrWqXqlaS9pNG81KQYQthWTysTu6KhRoSclEPxJXw94HDlz4jLW00zy
/Ox0urxEGkgfn63cONBhJgGVHn4JryiBtDFFNtQNEJ4BhI9XEy8dvC1SzEtk7ap+Jn2MGyvvtJai
3pnrPGmiHvRzHp0yE7XKiPe/atBI0fpVMzhvo2DtSDCJi171b6LiFjV/9zb5tFb9fCHBlRReZ6zu
khBkZ76xaE7oEkvRzAjatcNqJhAc32houT58TG++wzQENbmu6qELh5XfAwHjBENJvFw4c0RSslZ8
EZl478vDEPMG2SNoGaZvNlyrAvjPUmgcYGO9+iPV6BHGXkHH28zvVevn4zpAFerfeWIgu+aqeySX
bJqK137dOmYKqUzNf+hY21RwpVNGXZ6VHSlELHtxrSin+3YhzrakBW4Dxh2V+urGpKPXxZeJHv9a
sXMvDes7J3GZK/XWMIct0z+y/hTTH3QZiI8iWfSjQcJZybA/SQzjKTxoRYyoedvFYljYj5tdcCs/
JE5jC7bLLmjo00kA50FL3UiElRTWr7INSH41Nrjm6D8mtzVheSB8K4uE/iNVx7hiFWkCtmZeuU7G
QKCftjLohAgBbQVpWACnTjq/EJXfSHPsoevTzewfKW1PXFhrt9tciFFuMaV5nwyjF+QEbYV7MaKQ
7TwJO4R35QhdvlEzQX8d5e98j2vZoPzmu2XCjxbJrBu98MGz95L4B54nYIasvUONhEy8+hTONv2a
2Z9QYC8Qc0u0QuTOsC5K6jJiQzr+OnBdmwTim6HijjxhgkiuQWqVElmnVpz+xngBjCfJokLY3QRa
RkbSWGuCSEmSfc9Y6aEYXT3kohPr9oaV0qrQ4ixc4pTV6blHNOHbiRB//+bFBpq0baWHeq1LYBB9
pfsV/+gtFPxV7hB2fdhPnrDrOBF2poW1K0rt3kyjIJNX+gSTG2lHdIgm83Q2M8HzvUorxm43jw6P
PLq6Ul1OYvJPRyyGZbpZVW4kdc7VjABur3YaeKqjxr1bUzUldSaybZBUgDxeXwaJB1f0s3s+Ymnw
tCPmYUqdgCRr+lVMh7X9bR68lAVDH1SGauY9Ao1iN/Q/acAVMomPhzSVlmqi9NOcl0XStelZZtzJ
7l3pDAYfYkF+t/iLT5l0GmvVTvJMO0eguee+HSEf0496jWX9XUVzQIBUT9G4kkONpRpskmE8s3Hl
ZWLf/JCd4IsbveJnAEsWNTKFDOkzFKI3yUMOoy2VciqqCy0q0cnE2qc9K0Hr8Ts4TisjtQNwXQaq
K7C9myiRBvORsH+EvR9FBqfqsDEmDlJFOqjW2dqf39BJHZPba2P31kj2VM3YNF8smdQq1uKiFEm7
BzMXOtcqP/e/bl57Hn4YZTeAYY2DYN8TvuDgUN/TVKmi82qnczWJubC7p55XNg0KWJoM/TwF8p/C
0XyyvSolYQftiRyaeu3/SdHyEf7TXoPoY5dZlpDIpdMnEFIuSmMx0qpt/+QMJN6QeSOLht+vBdlI
LtknYFqK9XYiL7LG2SYNbvGWbZVzex1X86OgNAJG5TlMHq1PkcHN8vII5URQDEov2bNWUPM4sVMQ
Mv5qimTXC1kpRPB3WVkztHHUGVGFXb79LKIFKlMLKbCZibbcG0mMKeBqZoU+5gkNjxsH5VDfCqLA
TXkIJiQBoKMacxTXT4jFCnLVf59zoLyYOZjzMy/r3q004l2lzA4/+lX1YCPD5Un/TDThsxvdVv2w
DYxo4ZNgsRnl12HSOnpGjAb9TcPRDZBH+Us4R9VEoglXOxUtPDc7CAFZqybDA+z+tkP+xRXDUuEt
apMNQJworso0Ym3tiS8QVxzguaCmoth0vuo5VWaI9rUQx9DJKjgItt1YHO/+iMy2AgKivyaOUK89
x247Vv2Fb1McJ+prCl66OJbsmODsZcdfHoFX+pN0Qs5RrZ3tOm+l+Kij7P8Z5XOA4QQ2oesf1MbU
CbzLGT02i7cD6/gZDd2DUdxwueK6QT4Q/q55h+4z4s87zuth29tkrVea9n+JxPsi5sTVZlBjYX4T
CD6O04rdBKBLIeZn6M3MlfCjRZ1VevlywiY+cs6GNQMnoPYZTEZ2beJ1aaW1H5o1qdPPo1Bb4Jja
zm9/SDlHih0LnTzA7swvTGrC8hLuw8g3xth7XN/i9jmCIYAfP4jcB2zZBuhLV7oxawB8SlOJ6Yq/
8WQ5lV3u3bFpewU4fETrl7I097aXhAjSKfzl4YVHrhwFKVqgJ582IK9kiqFd1PKR+434rzavw1bN
sJYyU9QxuHTNQy3e9WTr94EMoGAzNRh9ce7kjwA5CQtzpSBNcI39N3s2CBc//Ez/g9pu9FbDYt6R
2wbj7d80jHs6jJx/IZsHSE8DJMRQvMOaehUt5z+uDHkrfC6K7w8ouBalMPBQffhHpG29ynTRyN6z
2C23BzCDWAG3zJGaeN6j9UHp8ey4Xoi6s+vJMpmPlEB8q5miikLRLiU4Ere46g14Gz/+lfCdmJww
4qBT/oUdtItJoQGWzVVBLmXXz1iXRvVFs5yf/v9P7YnbstuhtSL24FqQM+OM5OIHpbz5277um8JP
KgSMUSssVH85rxoh4ywsUyEFBHc+/NZgSNRcUADklx8wgSVjjGHBMe2w0cBUFEjzXtf7HnH4LKGD
JOuq59Oj7cFZVauKzXS5ca+/zsLUnwQMHnQiYe5aXv7I3vYsXJjiJ7YpzW9QxRmfZs3uR3O3ighR
36uDkmgyvj+3L4O/XLB6vvWETcWwR1VR2qMrHvsvwZ/NXLJ+G+GRgzcfvbK9g/6J8YTRb8vD83lI
mhYYF9lI/XUm5SnLIxp8atLRWuHtICUy81WUinIwYHwtpHPA0oghD0zxAynnQORLd5hOhhMRbiw0
V2HgI474TZecLIrRnSXXx6rsPOVnwryWw52cOvibOSJPNk/MEfg+9pSpA4Qqro9QeofN9OCj/oUh
3Z8lYgIe8SD9GuBMdJgDlsWa+4OdOBjnKuZpIzkE8+OWjPyr8QJpfgw/NW187NCFYzjgDaN6fjTe
zWcjuCTpc9wTiRC8SZgEZQqIw8DgOFFeBkPxuwtzOC17qJGoFt69Iahw73oefSpBsTKsn3fLkzzU
nciL/LcHbuDmihCsLPbXUT7NSUeAqylgQJVitKZLF5t+SHC6Bpur/JY9FFE4fDduTGuB3akv7b7h
1VzjQ0o/gxR1MSBZxpVp+8tSxWwJ3V4P0gBIZx55juKduW/J+PeoER9Brk8B11NPd4GFOqljwLIx
fa8zjI89Io1jRKF+bAW8FJQTxHC+J0GXtTRl/px9pwvojXCyeHbf2IXeNA1DMcZgzgH+pOg4hfhb
lXOcSSRRipSaWDdmacNW9S8FZdBMvKCEZFHZamSwmj1ARzGsEaLmofIN8Bu3qluCCXvx0CZPFlsS
UbzasAAyga831NZnPmRYHu1MAaQ1oXFe3ANpIWf99AHImBflLMw2Fqa1q6khGYRoxjV+86lP1S4p
EE2N/xzv9AKTKpLmWVb1vvV6oF7l4lAtiqdX7yL1W+i14GY3cXxfTS6G+CULEPz4/SzeR+JeQmAg
isJKmMnPmkPxMlgVh3NwQzbVCoD4sQMzZgf892RTQuyCLaOpdhWMkGkAWiWMgMpZs61w3fD7IE6b
Ne8EgS1wUxh/prnJgKUQ8HPCpsxpHIfmuy/lrG4QdWh8YWVDR5boapwtwA9+ORjjp9DgswEe5TV6
frGIht55hHKVw3FHJryYOvt/ubFdUe/zxoJjs+sFXD5959sU0AtFc3T3jt07gzEQhXRYsl3ziU/m
wTlyhBluaCw6ngFIkWYDWCsAc7QX+cwRpT4uW/1rAIMFb0K3iI9lSoRWwJC4FVjHIEc75ojvoZWh
PboauGmDCxW0svZdo3rNZ7kIN5GmSX1t7Hw4T2fl8nzZe9MQNc/slnKv/OStX6LBFU80phO8M0Jj
BJXlLUvRARppLCWiG9H0GTR95qnGB2Fr5tZp0uxZxddIgI3BnS9ELEWXBwAQHjXGktkdUX65UkFN
chufIQwBoVgFemUANDpOxMTE/Tb1dUPohfJHmYeCrECFhNCUnm3dDTq3PxOhE4tOTXVOZiQLE6+y
r9eEMc/xTEMNCw6m3cLzH9k1YN0AxbNDlKhi158VRveLkFzHMAUyMvaO4hWpxl6ZWyumHaps1gbG
1vpjwl9/K9wxmkEpgC9QBA3t8rH+2cP9jZRdw20yzwVrrtdUXY1nlG5net0mGKDDfk+B87z2ohBf
igHGRYZbsfpsLVh5IzmpO4whmwRN+3g+6JJ9lZC3AJEtzSobqzsZb3UfAZ7np5EWKKOj9zkSYD6J
mtCLIueYTna/e5U6pSTPxgA974+bjN6hp1wPcpj1E6PHhWK57kRmTiYnRWtzhkxpbsqr3e0VRtNy
JVof5aIFZpxTOuaht/+2DL9uYM5g73zlRZiJ6Av1qHszCj2l0z3BohD3E7aE6GZVL0UVu4bOZ+tl
pV0P8AEwbQDYWMhaPa9vrA8zS1AzGHyk47oDekJDB6/CGfaFlibgsrOeiFdxwj7wtTEoxKQeJWPx
d6Oy0+5kFWL43vIRkePUhT5uRubli2xwK1uk4CwukGs1+wZip603qp8qsSYN9qoNORVKArkkvROK
86UVD/boJbsi3eUOZd3dgkBIHMtMXqU0lhacEdK7mS2xl8A4/1MyBiu6FncPt6ohBaj9muoYSuC6
v9S9kiHZjaFVqTA8XF5Qi8mOljyxxBZXDHgxMgXyj9gxrAQxXAPGjltrrTxh/y6wPTbGYtqyGb8N
j30q+iSVdxgi6n81cs2/XlAhwxQJ4rFl3PJkpJOELofD9Sy1MIWfAzoL3s3Uf99+6g63T5ZhdECV
F1ZNR4P2n7crVFMRZesycGlqVpaTxzvnPaR1ujiQiUcoAJ3A9S03V19a57gky08Kkukt0CqHzkyt
p+NRYUf3jK9aUjqCkTNjjS1ep2A/vggzTTdYcNMIioBAzNPOwI8cFiNZ2oRV5mTkVxGEWUjDN6Ep
02oVfgmhtE2gkbLu5MGTDxinqEtKwsRmDWah4bC9MFO+WauuONQfZJg+zvqmrVlJu1plQFBaAwDN
M1uNdMqBnEw0bJNmiPKSW/u3zDQtsVIScu46fYICbo24WtMKSFF+Dpo6HkB27t3ci+Yy/p4ZxnNY
L0+rE1LonHVBP749WyiC1b6hxymbF1a9kGtNaYWjsuJpQ5NEsrcR3jAYBh4xGve8FSFauU0Xcgbd
VduY9kZ3j2Sra8Z80x7NqoNaUc8IaYxEpCZQ3Ilow3mCJSQsc9vgkAEANvthqQMtxHsJDPcXYjd3
MhYaYUvKMeO2s246BYjknGW6mAbyFFJxn7/HdqohS7eHwIBAl8GPO81jLpNPFp1CZO+ugRKGnam5
JHZHAcu1ItoEHse6v49FcpQgObYzg+XVvMauLc8g7vtbx4Ibc0/xffk+GDAW822rdgAfvoK848r/
fp3Red/Y13rTWGqLMuEVAo/+scZkpqWrTtHX1XcwhefvbDfKDJHSmwGzTShWrvlGxn9HkR636O3q
uhz4ppjnfeJV2Xj4Fx5/hOnWPwuwZ5jctMU3WMrVxyty9K93TJIvQjfTZkys6sDAdvJ2qUQ6GMAF
lx7286bCqFCzsNb+kCMb+N9/gf5B8rfPxadoL683jjoTmnceOfXtiUqHQ3MEjSspuBLzYpz4Hyy4
NLQib9Bbl6pahghGqXQu/vwnrlR8svOrcUSQQXyajuO4wb3dF3vQBkZmR5tQ8/xPnN6s6jmb8Y/H
K+RE38y1WW117S1JyxwNu4lHSUCDaQQ3GhL2rEqBYtKjrRIIh6L3XLxRGc5J0Ae8BjxVMgc8e0Oa
mMf6OyUE4AlcBw1DAGLDCZTCjURb5+RL4RF49qhlzWunzCm3xrSa4JpjL07uAf8Ot+syIg+g06dr
rXixD7tklFHcTPkcMDkZFhzCpvnx9/bXakd0pI4euxiKlFyAS681Z6YgseW1+QRfn881kh75xxQB
Tnt3YF7v5/r9FBNXr4xGHNklH4p1yeTSzzqt9ruFEug7tg8DIagz/7g/XbXSpRb644fM1Whli+DX
PHzrc1qwjdiGDG0wHwfIhYmm1Wb/+hIxJPdcdfuOwLTgEJB+u2QSk1gsGJC0BRJQl75GCGfoCuHM
3dAJJvAFiUTLbzQZ2vtVssY2p3aB8s0nhw8KcGkDey5VHxwp6UUYOmWMrouTnU/xSNir5T8e68EX
K1mrm2iHgUaMjlnVvdsb+ErtkHdFC5AfD1Q2lA38bvkkLCaJUrZNZpI0QkCf1p9o6TAaLxAwwMTv
RYBnEJeJfzUi0l5EJ1egrBS6cpPcVchfSYBDc/Z1Q6JQhEomtG0vuoqIKo9Z5npKMriIZCwqlWVq
odxknlb+hBcnj9s7n3L2X3V9NxgOQmZF0+vjid5uMlaf+1ClvTsCjv4vhk+tqjVpGwcRMVt0P1xI
j87v+B3EPegeejutsC1cXzMmgn/rDNxVfmL3B4XWvf+CK6EPN3aHYrvSIN9KZ0nZ0gg5EoKSc0RE
uKkCfJE71vKvBZjcG/ASOn6Qr+b4DuryzjiJ9W1fC8jA5bh3PaM5KgQvMCpIxv+P7GcgRrOoxpMg
PQHlEvtE68Wjl0Vg3PXMXEU9wFH50PgKvSRPHgJRxG+3mSJe0A2eDiBiqBd+BS7Ub9Zw8eaTwc41
P0eZ3oKiNUwWzzGUsXnbJIgE/5BMWX440HAOH85tS6C4gzg2/+SwElWChizySSV+ur09z0b73RXq
YffkTVwZzJDwElpXGCFygbU83khWoDifIjXmFqrn8Lvu1fDtHXOPujFQZZNG5hghMIUa3G4oSrRv
/BBiU24bXOuiwfDLFB8MJ3bupf52hhn8gZNmzsXBvQckXJej17hMffKR1G2TGioXHd8MNLGIWApX
rvDD5WyhJuh9JqrLFZXnZvZR4wGcHCm4OwmXtwLkCtZ2dwX8dawJ4b8HSZg2dF6JnNWPnJVX1uX+
kEXplgHOY3RtBdpKyZ9RXpHgoSuaGIKY8++b/stCdTF+ANLWtY69jg/0vC/T6MqVVhjyYjcEvJKq
rJtqKlgAbyPWaM8VCP3ustgv44Jjbmr3MYDuheinWIybHWyufIHuDBwsPb+W4P1hPcxwf/yowKgm
xO87ul22tOSNBSTbrTVbsPgNvjtHjfB5tDzfkzt/m2ARON/WNVLuUIMOc3Eeh248SsD01Z2YVNO/
YBziD5tSvcMrQJgH8rPTzSGSDg1nsLFT3X/9GFPaT9vOuDZrKYP81ezHjWF9wxBHlrNFRSdeaf4D
fSTJvEyyeyLYxcbxteArJV3wrFOGJaJIyMKALeGP9uUg6ZEjM0GRJeb2RYlP9ZrqVvcR8JTg5Htn
Zt/ssQIXTir2v/uh/a44cDh6pmMgTIFqxEdA6bbQrGjJuHqrI9jIKtdAuLNzBgJMv4zyZQ7U0yoG
2nxg4b9xekoJC1dER0aPVB4CVjWHi0/xr/wDHjZdv3TFkmaiTHE2nSRZqzv+AJ4ke+O4V+pW6tj7
gz8529+d4LWCiNxAoMVQFriM6mnXZQUc4SxmtB2exri+qVVZX8C49v1Ck07GQdE0WJlevg10MiJ2
rSDyePky+nzWAFkwC5HA1Zub1rGezPScKEPVyhzSDPHIGyUw6i1wv0Yjb8McTBAG9X/mN+eXElQ6
9PxoG2h3yk9nuMCzwC2jP9pErNfnvHo8Jdj0HJyECaiEbd2VHQI3Sl6CwYSbZosB31S9Jc1+8Za+
Aj/plA8Aah62YXGVgTilDjqmb8mOD0GMQgN2XZS/g9yDrliWTLJXEI4wC/reHFbrvxvOVEvx9Ln+
7phCuTAd7G1KUCBlXH0jAGe5Vve4EAWZYOpe1f+QwKyVqHCchQMybDB0aeBz0+f1EhNzw2dCodlQ
vbmhl+RQ5MtFEBrTw2whJ9pCaU+d040fLyW0H8xBPQ/iSZBxFkOHpTXYhQyy45tSxuBjETFUQCcp
zGSJKQA/cGEfDghesq0vWYsn5ZWYA4Tp57B3gZr0ZCQhW80kpBw4gWKPzNWIqkJbfI1XuXgG2Tug
zmmqRD8+BBQywoYu3iminLJ9OB+J5F88nkffl5jrBKr+kB12Tr5mOU8V0KFCoB2f2FpKeb92KAAr
2qTlQfejllOC9YWAa5sctd0vw8CwnifjN3tjCEHvSGwnGHZaLsHl18SAuEzdVVcmjEnZAt8Dud8t
B3+DHv2CrYhlnqLEijWi6D+9qBNuDbklQUx5Z9oEoKlN6930r2kpFM/GHUOmF23gTerV/v+30Dlj
vt8qFOxm4AJdZHEubEKqD4P7OIDjZ1E6UaMgol32KnxfUe/orM2HHHFDTQ6mMfoyAhBhPQqokxOy
t0B21UwuSUGVHolSAn4RlLCmA7ZixcytLna05tN5G/3HUNONrFFnFfISCdEpMKOoIsTAmU17Aogz
luTXhm57+WaO/5oJp3L4LITathhPh6N2OvP31kWnvhFGe19s+3PSI62TNR0RNWu0ovNLwYY3wJ32
tY5e9+qkCv8X3Q+1AirhMH6jyqJXZdfv+rgTxJh9TSiycPYiKYtimSJMAxrvk0qfplOCMUhbnayz
MTpcPPYGCdgi2OIUee9f/niXk+J9YORhJ61Xj9HBgi5KsQ8D/OAqGErkbvjnwiQ4bJATu78Sd89O
ao/UKnuJ/2QymoU+j87fnwS1XE7uLo6zzPnXciF4EgaJwS/VFyA4nj3OYpzHGGSuVFf5mnUi22tN
ZuGyflaaOCoqKofehqEZReP/M6wIfyenFJ+gYyrb7EKIocKzquWSo/dzJJqnb/sqhaG9PcVC7jd4
WkMASRIqrb5Ye6sJkcDWMoitrIh7J/YNhCIrpJ9TG+sH7xjgZYZlyTWo7U9IeXa2i62ZwBIFLpps
v/OhXg2Jr6RF+71b5A8xhKjv69FXinQH8ADEagcyNxi8PKcDkjz+7E2sR+F+KNusbDL/1CFIQn3y
qxAQNyVugH/CLq3Kqdc5Y/vysYSOn3INeYAdM/bvHzCdxRnaz/ZsjUTrhezYMJaKO6nIzVYUeDB8
RtPnwr8YEkDqUzoQSQ0nsOeNyzHIUuXdU16o594hm8gfyfhsYkicWN2rSsUb8+etLFkQuv7d2yOy
2EM5Rr6nE1rGFR8oPs1gTHGwCt9nyvbfakDSdowK6Hu+PZLXFq3ayR9CfglWToJ/heD+h4CaJB3n
QmqH6wOXvy/gFZoaaubLFUaDUCw5jRK/vycZ7DRZm7fyjmwZCPZyuH0ofjC/u5OPuQIfucyaM7Ic
jF+Qei/LTJxmF/nD8WAtmtpS1cy6R1RIKg/hgqxXKTXD6PQsGLfrzNifvqEzYOg1iyLrjRJp4I1r
/HlrmYHkqWHseD62UXrf2Kll7DNXhpZb0hJsMp5pXHJ+OrBry7h1ecOFABHQktCe8kjG6s4tp6XB
wYm8ybsYWE2lhaRpPhr7RuXlJNoFKCoMUIZ4sgo4ZRZ00nYb5OXr7Iud1A8FLNNEgnsCXr8q3Jx4
Mmkjt4dbX3Sx2ONMX/X4LJXWpjiN6Hc61zdyBEeu2qWJuAR0wKY4jL+CzwQpHMY9UALdiQ2NjbQT
B0Z1g/SF7Pmd5YNECeqrMiDGDwePbH6YGEw69sFreaNOEbd4xtpm1LT6dTmlZvy6ev3CP6zfT3SN
2G1MAFMKfQoWKK6FDPbdaIy1LDjW0bxkY/T+KtP7th4YntVVgXT7VGhP4nBEPBQx1xah3v9HiQ+V
7ON1mSC+SaJuAqFVE5Oc+xFjNWL2Ex6z41ZlI81mu1K4I7s+2REk7BosgsaCLagl5HivUpEiFbNg
yAcf0IIiRiRuFyI2Y2MtQIlny2cQHDVJC8i6R27/tttfQUL4/9L1bIpdFaA+8cBYp5Zp3Hu4E8+p
gUIgOvJnggeotePoT6gImucGNXdw/RGX6TCTeACVW2r1+HYmmQtZ3p/W+500I2qJ95TDmmiqf89x
AHWBZApPspMPHdlS+qyJxIVRpZA8h9RfGqdsUHGVlsvOl56gOv4dIbTKPqT3vgczyytuuqwka00m
Gz80Wvp2Fvb333kD1NEg3JL/olk/Vz4uWdj66mL6BC2dW+A9yboaSv0WHoUxPia1CAAvDWIz5WwI
6x6RY+9kN2uzS4q7yaAV4ERrlq1COOa7uFBngT505PxlNi/ZRLcZ4rLA1oQIiRFJwywTNgvsqwTL
Vjqi1U4qPyPxWQM2RWNs8OgJ/LXAo5edDGi6W1vRc61gf9MCmoB81Hl9rILeWxnT0xhRlrQM540A
xypcfQDxSZ2g6bpqX6lOzjWjeUgjlhFXOWcmrNXlGG6oqytOoqnt2M+rcsg2062fRdtwZAu2THFA
Ag8aF7MhYiKSb/UbdG+K4zz0eQjuSMQl9IGiudQPoTl69et/vhy/dWBAfHkwL9rRyiUjlxPciLT3
lnLUE2FNNQO6cCr75F2mjPRV6CpJwdTnINwD8rNFa9XrCE/qAsrpXz7eFM5ukj83NjuMz3alxSM8
iLDOyJm5+ebRJyCWv+DdRPudDudfy+0jfWFsF3sdcu+UiDlZ8t3OgG+2CfcJF5ydLiGWFe9hMv8A
4OeNejd9XxiqrGUdj1tuqyykfgzqahkWw6tzc5VUMVprn9DBY5vMV5NmP30r0KLO11PqeAChuMN1
jBSf7P354ZKsq/Q7ZKQBjsiHfAq/ebzJ6T9Sjd18QsLZcPAU5dzgoSXUZNQdfbyId9yuMwWOIhDG
1kw3qSljaRe/cZOru44oZ0VhsmA8Z0GSW13CMZBBZ58x+2oN8DA9ibL/ZbrO6z47FGnAr+rur4to
lMx2xAon4EjuYPR1KXdKl+Hjpbf9dtM8x4rI2hOJELqqR0fXCMmuaP90msbDOIzeMOAqBS0nZN3K
DVhcTz5e0SvFeJhRY49x14vv1bGs5qw9vPjVaHOyqOnz9dbeZxolD2gOOSbO+L2+jiyEUd5f5xRx
Gi6nIjENmB7SArM591E9a3GwPdagmxd5Q+vVMrfeiE2okGkIq06wAeAB44Z5HbCkxGnvgPZOh/1Z
W+JdbwdIsb/YCvY06onIPaM3O9mqA+Nmh3MTMfKgoCZDBg/+ZV7C45kw5uett7NYP+CcgV8c6muc
FIPSbfLlO7p3vGQRe1T2wtgugbcxffr6K+umLwLIVVcUZmndTE9LuSwCeOZ9NiGbBiKxllb2xoZL
X7NDJUsPOvGl+RKVT3zL60CWszEmH7aja6BgyshXMDTAWpqyxEEWunNCRox74J3Dj3ws+Nd6QCz0
Mq8scFxBdMCED9HRJCEfxykUAdhhuuh++WnREc+Vj73e9x7rZeUZH3eOY24iQusD4MtxZdFV3Vb0
3AlgND9UpAmRnLnMqSWLdw1/CF6qUNs7rIlv0DeQ/jhqvGY1ixx5hxCW2EIHkDAVifdx00hGxZF3
2S60Fx6PSDekTxPlm5sIFTIPyPM3WTmoHK346FIoiXRIFmlIPJcNzDiLrF5Ag7nIhhZFpJFibH6p
F4oxS36bm60L8+Zi9O55F7Iz7miR7mhWs71nM5BZw6C99lK6OdtBhsi5BaMk2cMNMWoJer0OQJDC
8913jg74RkaeuZuwm+8B5ZUcgl8BW3j+phHO1WWIKVeoN7Obb/0VypwbN9gNp3aClWauDX+/Hv25
dGjgjaqeDdc460qpAYSqImqXeTB5kACwjQOUpRNstmM28vk87fneUqJs47s/dyAuGmcmv4IoXQCD
31zJ1jR2qfH719lwnyaycGiq0/bnPIsQxM3d3YGWR/jriJXbA0FNa+TFj2m5oYHJ40UN39xk5WTO
E2234hujkXw2Ys5goUj/YNcYwfWbmy3fkutFTKnfk5Tne+SHpNQqgg65CvRH/cAgg0+NbhcJvzpl
UZUHOIipKLBxBdHZRQvMGQ8nLMaTUaS+u90nOpJhDFXjwqFF9CgVSOEXz8U+9FQk6qdpUFbUVHLu
cQBmrM1WqPoZHdodwB1IqalqFXjCa13S3W5TZN7TlzZMjLWbqu1FTp3OXP13Mim+EDInIR6RzoZG
F9RwpRLiKXfVG3YhNx50Tf26FeCP1ga9bkC5DMuSkvCJOwgIxo+4lbXc0W2ChfgI+ZXc1n+9rqL2
ItHjw5aUfWcZB0RXxmw7G4OCCrcxKPE/mXkTWJ4t/IcQAecWk5M0quGpFNXuC5tNtNOHxA/ahgJc
1YmEa53VQ97vO3WQooCoPJdC0XhilYJrUOrW6eO8+zEpthyjHVZAoLXSDXtz2U1lJ3fTsXs35TDz
3GXJd07/NEg6cGVWrIN3UWjnHf8iJahehM46wUc+MCbaXGjfJoQNOY2F5yk9VW9j/NgwIiGZegRx
j2FHdX1FouurKfXKgrnd6FWOESE5E/la3z4FuwgC/IuhJk1cD5M4VjJls4u4JJFcWoa3EhhSOcPn
Tne0KzDjDZFeb/DWfK6MhilwSoSN1PR3LolWZoMmSSd6UtLBl1awIIAcXQrdhnBkVI8snZu//fs4
HQkud0lhue7zpn7hKTIojjIhieKN8f+SJe+IxDAx11UjOfyUx7AiXDfx69m+ji1ZrRHYESQPRrsk
/QdIEIE0DJTVt77qLqO0D+CUB3MpSDB0J9fpIuDN/61Uy4yXrJwqDri0uiphQ3fWnK1WpS2xQwCV
oBIBwaBJlPkhZ3IhyTz0SZKwvxJXL7ZLXmiBLLCw6psrJ4z9LOjkJWyYqQ9LKHaHOUOKadg8iciB
gW+KeHh+OLgltpHatWgYjjbkPXS/lTCUSCMV641sv64yB3EXCW2xqoDaO3vI2FD8Zi5IwmvuZMDI
Q+ZEyqUWiZifWhQeo7Frmb/CsLDT+OREzJdY9pbeT4k3oEt4XFFpu6rKzzuOFR/Fme7ZHYewqhHk
v8G2ZkGoOhRXIreBj50TIW6XeVZBlajof8aHCvQwrRYtlpKRN0+O/7a9YyOwKoTJEjImqaIdWn7a
5tUfrcl3Mu/HIReJtAspsGBJ5t9Z9OUQjxG4TGzldBrWf5WDmoqzWjro64uoQG5hYh1JYMIRDQ2m
WjeHhP9HwzMSjB8uVXTAQpTrhzUe9owiV1ClQQn3wrQ5h2d1vJXWbvTbXTBlh4IT5Pi5YIviie1Y
2DjmSZ2MFxcBm57kAcQOuR2hY+CLcxAGSwlurIncNLEUJF7vMG2O0C98kyNJRG8IY6CdbhUoiOSU
hlhyQFoEYI81JQZxEYNaQ4mmSxNLPPe3nM55DGIUsE54eYomhzBlOBp9bjV9biGp+2d9NiaHBemd
tcQBBzEBi29MCZIvpaykSpcA/oY69EhBNNSeiNrNW1Q7aVaXzttbzoas5jEA0VleFtKyLRWu+OI2
mVAtb3UhKUZDs+2s91y2pi9umVdeD/Lj/qDhupEBX66vmBAA9IbnNSq/8TZfPShYKSD+c0sOvhvI
YX7fJCWBPXfy/SlufacH1BSeQ4MqrlrL/d/rYQytQX9Umupwc7BYcUJIJFfa7s/u2PMAtj1Pf+1X
Qr19OQM/C+iVIDCp6TSAMObENqbeLXgcuTuzY4dlo0uUvXPyXgsK4b1vLKxQbhhqTd17tKZBWQs1
n3qBMVWiMfrGiFOm8IifalZx4QlZeCnXfQRtz+22z/1C7ofS1bsplYrZjWtX0KDAeKN2GVjP703f
EUNzhKXElsh7MxTtKlIYcdla5inx/Anh0awNR/ZMfoQ9Rj9t0tl99h4HrkQEwri1o+wsQtNyemIe
0UNm1zGoJOBOViTWvdre+lDi669uVwQRJp/p0qDIgiOhXC41zoUpiJ1mxq6vaFrEDPn2T8/1ycBU
kWfb7gB1SUPap10b8b96+P7Sbyo5/5L41AHyK2MR6vcEMyN9waX6zo19pOtyeXC+WMBv5YW5uEsw
nThVjjVYNVIS7IfieCbqIJM26JFq5YmPQh6e7tmmAMHTHlaJ6KCec+rR7FIlkIRTGoor+5CbvzHn
OhtZhxgHQ9FWMUYPlIws6qHyZjZ2ea8BHFqrCeI9OsGAFzLSBFugcvv3G09dhGo5c0lY64+B1d80
+T+CcP3swppS2C7tTNwHwy/W0ePCLr0OcAPTcXd7HFFA6NjELJGAY46SQuGOnQ6Dx6iJzVTqDQl7
sHpald5Wmajk1OriGuPXoggfxrSPvyRiHEnIG7eXjj+omLgRDmyiXzIEa5oWkA2+Mn6dB5g9Lfxi
5v3UgyA2HucQsWkMI3VkhcyYmB8eN3akcWzONjizWnqWH2ABXTKNAqawFpqq/4bciInZSc+yi5PR
7BxP6J2chgFt4pWmvx7Ss7KfvEaKNc7XHq73YNn7DtczBqMhJRVS7y4GgPydsNa4km4crleWQlHV
Q+D2NJa6u4aZdetL9/pHNgNu4zW2jZ+yFtGIMqKqF8aVNpwmE3fkYVQc+h3V58j9+i4TCFaHXtHr
ae2/JWF/dXqLYNXK2B5bC+2qdBSlpxhL85t6YuH9WM0xMgwS/nzFJZat9lJ2m6DmDjAySITbWjeZ
eLIUZAvMVfhLHCFktZB6GLW7Ur0Hq/a3rpZqnWCxZVrVbihQtRb/MFXgineHCtpz5BAdFQkZDgdH
09UxiDukGsv1lx5xc0rgoAo9Wctb+7Ct/tgJkvKwQjzkHNplHHBEW5NW92Atfx3/RPxwQCh+O0SB
c3NExFV0HReQrZRx8IcLaZBSFLQ9yvtBQMGkUYVSHCwh7JDmn50ppb37V1aDu1rgJaoYyDWwkyYZ
sx6PHZELyUU7pVUT9I7QO9AGze5rQ9iL+TzjDGH8keX60O7M8ffIXhnNBiBHOxRNjaVY9hTdNP3Q
l5fNtAs2+TjENqx50NVV6Rs34kUNoRbAurzjoDO3ZNQBVmQsx8iRkRHFQtcM3IlcAjS9z8e7tE7N
A5GaWz4qb4AU2mc4AXWNx+T+JxYkRIFEeDTQkh9lN2BOx08icIp3ev8c7Mu5Klu/hdS8RO0BTctQ
SyXflWIbRPRSF+VA4zodXQpS8fSJ5tVopI/rE91J7KFmYHPbU05a2IIWYiXIqsaghyjLxZlQck2J
ro3v3/34m+7ISZ3scpP96Kd0PsvzfNB5q6mqpBP1ctNuhcqqjG1ODEIx8J6PGN/qHZsD/ApPQQMJ
USM1UW0dZgDTMAWLq915lOZdtc5UP5BHGRfKbCVHEGA60OSqdyXsgnbXX2wbbrp7N10cnsK6INdL
54Xsz+Bj3jSiIBIjg3cOvV7tcug7lXKUotv+pOcbZYfWylSdscpe1l5cuMAQcrlxBIaLekko6tuo
bZ4NlmRwyF7XE7xgMmBGhKTKkXT3BdbfcMUJPXyBry49t85eZqeQK+iWlRVSt70jTLMVDtMNwIjJ
sSyDIptZs6gT5QSDw/EBPCf5jFSBNaNIhNsG+ggzCB48739br5o6k+U85VuZcd/2jbHzvuIGNgfM
7Ve6/N8+Yfn9ovKiO7ewBLk02COsbKfH0ILuneQgmgIMFL8NRDfoDNoum7J7WURSZkGvHzhRh33x
9/jTDbAWoxzbZlSoXisqyXlauTNisI2bNo/5o/G76N94fnhQqtneb97ld5laIVbFtw37jBGcuSWR
djZLGgDtUp2DyiIku20r45i5IjJ350AylYLpUe+rAR7HttNn6inYt1xB+/G7ITA04ctHIhAMQFkx
Kcj8TQG2x5mGaoCvG5D9e69ZeyVoQKMMfqXK71O0u/RGl9/dnwqr95rg1j1qDz776V3w6RVq2Sj2
vrfgpgUhmCLKfGaHXaTvYYJa+mJb
`protect end_protected

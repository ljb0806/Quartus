��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB��1��F1Z\�IK�8ib��!���+o9�%zM�%���U��(���0�|���!#���y�.z��c�%�>��������Y*Yz�?�����+講�R/� ����ݑ�W!;ݰc����К��i��K�9\�� aO!23���
�1f��)���R�:�!���P��%��r$W6rm�M^h����*&���ZSì6����v�2���P_a�j�)�r�^:D���g�A�Jܸf![�����E�',���혎}7*<�eJgS�8O$g��J���L*
�k�f����_��!�ɰ�������j��� 1��Z=����a
9l�p\n}q��u[m*��Vy]��L8�9*"4�k�[U�ߒQ �.9������B>g`_��-=���&4O�8F�!Q3�m"}�H"n���G{�wu��Dܼ��!��	/��ϩ
�\֨���q��8��ͩ�|A{	?{�v*�VUa��\�/������T3|&gI�< -:�A�Vj�Z�Q��f@X84w'�I�$Q<$-�S{�6�kV���p��m؍�<��~d}@�i=RXA�x�d�Nr!,����HG4>-���=т��(pW��3�Kq�}�"��N�s!��틿bu��M�Q_��:Y�3��i���0RZR�x�;����99��|/k�l$��D���^8�ڏS�/�"��p�~C����k.�m�i��Y��#Y$m��O�y���҇��਎GM�\�hr|��]�3�>+f�=�O>D����[���k�V�oM������;m�%���ӉjS6�n�E����E&M�3j-�_O��BL�`/٨�i�Ξ��(]�hȕ{=�')�I��l�4��I�\�t��P�,l���ki�S���&�ش-v��>BD��f* ��x�&��z�<�L����-4�,�ߧr��H��Ws��B!�S5k�"�Qm���Q>�g�KA�4�E9d~��jZ��w蠣A�EZ���H}�3�h���N4[B���0���U9*��8��7a�	��[�{<��7�DL���%��}ۍ��Iy��Im0(�U���s����banH�-4�������~+��H�G�	�~�I!���B2����T�TUW����7�2Fs˼�SZ�=����b���>�lD�d%Ct�����ĵ�Т�*I�ڲ��le� �s��t8����x�<�{�q�x��)
Ro=8���v���8fI��_�g�x!�����C��pO�kAS��T��	�^(���7_M���`��V&y4�q�k�2�j`O�*�"Y�a���鎒[H>F�iW
���A�W��^c��a�9���"�f�㿡xx�\Q8S����}���܂�t[�u�����N���qԸ�meW�Q�-g.�#�E]�>�.��n�1���#+��(\-�` \Cr��,l&O@���.��TA�ڮ9e����|�o,T���&M�y-���9ȕ�}g�n�-�����J ����.5�0�N��1K��EY��$��l<�X�tִ~bW�-G�} �e�g�[A��O�T���h���l�v�_�6���~�)掴�������CJ%�.K̓�J�Z�0i8��k���|4�F��zj"7��ۣ�/��f׮�w�?��^$�n�_o���_��H�ܘ�dh�i��F7W���3�+�:�Te�J�T�qc�q��޶��5^��[�3pO�𪥫	����hl*B>�����O�(&ßw��w'��dq~8f�����b{C�����@��v� %�$��с��B_>$�~b����N�M��O���xi�K),��1�H�DtXL��B����O����w�b���"`����J�O�q��C+�?�O����4P���Th��� �W���Wn�����J#j�?9or��I���5��A����b�S=D��BdOO�A�+���8˂�]���J(��x�;h�8+�J���0.M����R�M#�Vyp�E*�)e1�kLw���fj����.�$O�����̛q6��Ѕ?�v��GyA�����NE�i$%/��R"Q��Ab_@���)X�͵���?Eg�#^rI�q��������G��m}}$5�A� ,��l���_�a~���ڹ�&�JE��j3�*x�\�;�d�>n����'/�\��ΰ6YQ<��a���m�ATָ���&�HQ��^��=߀�~R�G����,�2�u��P���V�u�� �@�0�Eq��Yx������h�C����ιi��g�D��S!=��.v  D���ػ¡Lx܌*jt��A��5�Nm��g���k,�R�zN�D�����P����yE��i�b^��	��	�N.�l �t�*�SJ�xC�6�*�s�d�O�NC<rX��xh��	i&B�cCPy(�[�
�͕�������{v�O}��<�p���
��0��=��s7�Ư}.0p���Ρ�-����D& 5;���M�J���7�и�9<����r�O���޻�,< ��2�֒
��cW&��,���giE�Z�s�.�n��6\)k*�.c�+G����Z� |���h�+�R��r�^'�ڿ�Y��A�DW�| \��ʒP��X����`���i��t~�Ylj�	��E^g�͏ �ǑT�␳4K1���V�k�?��]e)�g�פ:�(��6(hL>���ش��
�'�t�\�탍I�}�xU��PZ�󣜀U¤�ёu�a��fx_D�H��a�B Tb�^��\L̓#g�{ƌ�rt��I��BO��I��$���	|�G��ٹvށb�ɤ,d�@�`}����"�.�1\�fԡ��,�躸���6P�d,�������ڄRI&�����^���9��TZYkk /H�[+
�(�i.&��.�pUm�z�^\ ޓA���=P,��s���4�j_WR���s|j=��A2\C#��``wJ��t�`�;?;vk��Љ�A�"%m�:�Cǋ!㤻g�j��1�h20�fk�huv�����g��Y/I�?������t���
�C�A\�JR*6O͸,R�O2c#�9���E_�e~~�IK^�B#�D~��D� �~�8�jh�P:#����6�\\w{��b1��C\��L�Y�����H�߲�IP�<KdU�Y޾߶�=8�e��Go~`ѳ��I��?���*Hi���-��Z�A ��#6���m�,{�ڜ��Fdq���5(��&�(lX��ȩ�Ew5&�����҈v��Q�.t�ͻ��b m���.�&�4�Ǝ��z���+L�҇%���%��%����!�8� ��Iy�J�t,��k�c��%��:���+"�TFme�'*7a�hd��"'�%��]s�ӣ�>#iJ�-�!���nPb�vgD�>�R���7�e��$�: >���i>S�) �YU8T���o'C������{_-C�5;7Ȯ�����롵�pUʏ�W)����y�W��c��G��쩥|��C��-@�Y�k�D�ж�-:6��=���9Xm�c�n"��cz_ݮ9���c3��:���a��fV������!Ok��9����l�p�V�5즸�2�����!lJ��*�J�D�U�Н A�Ö��F�{W2�m��*!���tu5<�.��>�D�2�Z鎰�L���2G� K��{Ԛ�� z��x(<���q�x~E�90y�g��#��G���v\޽ܻ���Z����0��1��`� ��ř��7�)b� �q�[N�
�f��������Pa�|��@8��ND[Pe���=���t�(���ƪZ�b蒕Gm^�M3x�S�^dW�|�As��la�eF��"l���v�Q���XŎFB��Bժ����9���n�Bb4�I�ք���$Lp��4�����h{�;�}u��/�ǩL���-�M�N$��E��4��?���9���9�����N@I ���o���(�K>/T��5�6�0,>/_�	Q��"�=5ڔ�S��|�`��S|u�5$f��DW�cղ��tO�A��Z�7:a����
6� �����k���Y�7��o{ݷL��L�J(ɯ�B���i�n�I����|rlz���� ԻM�FekU�xv��h�y��i��$&�c��ך�G�����pu��P����^��]������b%SE� -���!�]y�&l�8�X�FG��ABR�#/���/m��~V/p��2�8H�剳�"b���c�@Ь!#���ږR~n��A߳�e.�'�a북��&/�r���h �2T��H�7K�ϼ�M�m+څ��Y��v��hם�5[S������)�cNS䏱[�_���z�H#&�I�k�wLa���'��25�-w$Ie�C΃�hIk�x�V񺁷����E?5o�3.a���O��3':%6tv.��(.T�$k� �kVq��&���T�в� e�hҿ�u�H��dN�4c��r���k嗟����c���;�`�V���8A8�u<�����Q�g\�`A�h���\�E�2�͖{�=�=�NRV�B����3Lr ��x��X�J�cJf�4��F�h���3�����@�'R�Q���᎟!8zz��@Ԉ��ٿxZ�o�&�1�2�%��G9F~c����).i���D����F�	�С�}p�x�)}������Dy��w���{?����~;j�qv(	V�^����"�n.�qP�īi�G��1��+ɪ��b\t�B�#�´������a�WBȦ�|6|��
x��l{wPr{�i>���c��(6l����AIrc������K+���=����:fi��J������!�:�\��>�E�=�O������*�O��ά�]/���g�"�O��ݽ���+G��dL~dË�؊�*W���-K��%���+퇌��,��ô�N,s~q��7��Ì��+��J2g[�8�]B�D	X���#e�/��]jVR�#��|�����&�X�`6����`�Ye���-�[��A�#Ƣti��g���v7o�2�C��!��o���T%����bS�ڋy�s����I���B����
}��0�jI���?����1ט%8/�_AW����֖�9��K8ۼ�Uk������\ �yl>|��%��q������X������O��4\c�-\8� K���F��vΈy�#�[?(ac��j1q@蠮 jn�d}�6)'��S\F���>h�����N�X�.b^���_C��;CcM0RF#�u6�d��D!���	��y�����p���;����%s㽴�6SĎ�� (hi�=O�!ZiH�w���4� `��<z�E3�}k�ya�؄��������2�&�
�a���)NGo��QxL��6�+�~���~��g-�I�1~}z>+>V���>��l����!�*�RF%���|A�l��5Y	��^��y�W�A������[� "o����-Rƌ�'�3�Z��:/��q���G�sG8>+�����d�GVdQCt9*ݰ�2|<�����B�����y���F�f�O�mW�.���F��,�t���x�@�Pv��>��#ɂ�D?<��ݓg6��w�	��؎k���YƱ��"jN�����h5�Qq�"@)v9=���ۅF���ag+r��B�������N�-v#�ͦ���LVr���XaASK�@�3M)��n�&3l�S�e)�|Xۆ �q�����r̕S����J��Ug��`���l�Ϩ�FvQ��؛�T�l���t@�R�>��xg��Ȩ��A�2�a��	�OP���kz ��'�ڤ�&�x'�-�DUR� �+�cAo��U`o^3b�8�\oY�X��(����s~a┇)�	2�FM7Zp�q����~j���� p�c���S���6�e��z������p#�+v^�����@���3l%b*B+��%ш��� .��E��zwO�����A7W�.�GO�dKJ�Z������;Nב�)#�[$��wB���P�F%"SF��)�?��U�����鸥p�ijd����ap�|`�X��8�LN�|.:�)n��۲�sN�.���j���*\l;�.l`U�V��ts��|�5�2��,�eS�1D�p���6�M�tg�,�,dnD�y���Ch��9��jg��I/{+�͒�؟|�y!/=�T�:b�&{��	G�e>-wL@��O�;�%B�U�����K�ݣ�[������0������__���l�%��:��!���"A6��jW�I�yǂcA��Jw���Mhf'��1��JQ���3�F�2!To���J�Z�ә�R���z3f��bjS�\��J���������(�2%�J��M��bi���fn�o^�]�n\����ȯR��������E�W�a��"��/B�nm6�^8��7n�۷�璵M�)�"k��g;(	|�Ų��6���.�5�Z`�ׅ�\`V�UtL�8Z��fU��m���Q �VN��D"�>-,xU�:�:��P���e�mt~Q���.;)�gv��9��;G~ܓu���*PNq��K1\��)�~Y���n��Mċ֌ڸ&a�_І�ܰ���iC�Y)���	��ȽivRkF�5��Z�J?_�D8]�+v��^�(Qg�Ω�3�^��7���z�@�y3P�:�cHH/#N�?]Ňd�*�F��{i*�ld��!c�����t�D���@�{%��z`nU�������6a,�`�Af<�}����
>�9���!QhsYJ��O;��oV32Z���b�~��\#jJusH�����&�`WE�ce��N�Mu����o�_7�]��TVq��yڔ��5('m�$Iݯ�a���r�!B����K��]4i)w2gc�q�c�Vy2��!ru�skWli�����Ɂ@p?<���g��t�]E���RI�πے�&�f͑�謽:����E'yL?v�?��k�L!|�Y�=%1�f ����j�z����7���IK��V-��Z�i6W�[E��=��?�&�#��
�w|��d8�5j.��H�][�cȟ���l�ya��5 �����gՙW���~~Z'�HU�^ç8�k��4˘�c1�0�x^� �����?T���d�o�"6�ár:���ޔ\���e(��[sw����
䦈��y�vX|1�v_d�R�`�P�j�����1�m��Q�~�_�S�����J41_rnU7��m*��ApN�ѡ���5՜����5,�tr�͍Ē���L����8
��a���`���v��
`��j����O�c1��D��+�{���%z���#&���A�3���e��|i*[�L����2�B���y��RI��F�(�_{Xr��ɤ��1�	��e3$6�	t�wf���k�	d���r��ۨ&�=²҄��\�3���_��=#yi��i_ƥ��x���ա�nx�Dd$?�՚o�6zT�_a ��5p����a�����t�[E� mZ3��f�uZ=w%�0W��7�مt�jb��}�m j��Ѻ�Y�1�"ٍ_���j���aPlPy�93g�A\kD����/G��,��E���<Y�����X"*^�|[���F��G���u'��/ �-���ǘ�����'��*:�m��0i»�2�0����8VIo]�cC�����?���U�Q��
�jYX1�x�DlOL���c���)�,�⤖������C36	����Uz%[��a��<�_F�4���ISl�Q���?�kԔZM��X5[��(���ź �K�aQӕحSU7E��!:r�����f�V..ԍ��K�:�4j�f�E�A�Gxw}q�r?'@F�h�ѳ��q�3C	����}"7��.����Yk��*!�G�w9��+8�Ə���\�E��{��O��8rђ�b��a "�=zf��Ÿ���t-v�F-Gq�6�����[�}�d�̜�Bu%�($UZiG˟���� w%.2�Gz�K1�=��j�eH�a��B���Te����4a���\�T����,X��;=�� UY�q�A]��XoP6�_�C� �#�>�N����4�l?.B�W�S5(��F*p���L���9��*{6z#t��x,r���\����@���O#�*$5�|�&I{�d�����B"�4AEO:��S�_p��_2����������BgƟC��;���T�MO�����W�_ �)��ź�����<
C��Y��!�2���<�J�?n=3,\��3dISk�5:v�+2�ɮa#22V���d:��Wj�Y�mo���Qi	�#��~�R��/�K ����5����|��� 0�Œ܄��N�	�����9j�F.�&��p��$'2���h�(h!��7���	�?�e��Gt�79m mxy��'W8�`xE��{�M�}c8�j� Y��+��v���/��U+�o�T�9�I�$�P�`�ۏ��8����۶�G(����d{�|5җ�a����N)��aJ�1�u�gvF��Q_z��!`���/ئ��z_�mn�(,�{g"���!�[gW�\X$��Y} ��w(���6��B��=���%?Q���O6��P�4��)6/����9������"�&ol�Ν������
jS����xO��ͧ��cT|{N#L��d���?2��G��5���c���A=ÊLf(2���d�Y����Ţ+<5?Zj�(T��Y��B�'F$��aE
յs4\���,�\ݧ�
����!P-�< �Yؑ���1��"9Vb��'OT(����HH�'-ǽ)h{[:7�a\��E&�/\b#p4�ǂ{��~~!r-�.�W�|:�=b5�����B��ȷV7��#c*eZ�*K'-j�����O՞^U�M\�*	�D��TP�W~�f�ߍY7����R�ĥGS�r��t�z�0@`,�]��@������`w%Q�-X<:^$���ȅfT�΁��*������&��������!��p�U��\k�_�*��RƠM���/�i��@c������ò��ͲS�咡(�������t�kp��%���I4�5H���,]?�����/8up�8�ך��`j��������|Ԩ^?/%�"y� �[>zr0���vE��@��n]����ĈǠ�|3�����lwd���S�H7-���I��+������KeR�0����v?����0Fb5��Ǖ���?�O�C������<���!oAKl���B�` �R~S�@1�����E� [R�J>?k�Q��TΠ'$#�L�,�p֝�CI�8����i`�b��r@�1�z.s̺�yt����5<�F�����#x�;��[�Ô�U�Y�U��F(�YBJ*��g�XΥ �
�w��9=34�D��y��4By��9� �����cjcY����x��ݜ���P��&������N�t�3zV���!���=�J�I��V��	�k��XH���!3��Z���� Ċ�3u��F�
Q7�0�1~���᡼��U�>&/��Lo�p0�Bح\F����(Y�ٰ��!�|3�@�S����B'�Im?�=��+p�뿫wi��P�S�^�s�����)!��<�8��k���2b�B-�_�a�<��u�>��9Rރ��ϒ�����@�݃��\k�+�h����l��9�\_���<7��m��WU���L�t�����y�Ow��@QHw��]��HKt��2	7{Z�Y~��SI-�Ђ�G��	�rEX\�V�8_���__�Ү߫�||�qF�����Ը��M"������v�P��m5E��z[�;8���!�>o��\��ӓp�k�Au:��Q���q)�v��o�ϔC6P���E�|<!�tl��Ad�h�{���'�jY�3�T�Թ���v��:Y���������f!�E����b�����b��Z�f��6�8�wP����(���qP/�=k�����@С���p��E�<�ᔾ ��t�飁���ˬ�|�vvi�¨ځdz��3j��\β�w��*.Un����-4�I}��Ӷ�I�%�u�ϤkC��a<Úv"R�0^ot��V{��]�^K�%h�t�:/u����u�A-�J�(T���P���D�C���˦rV��b����T9��H/
uCA��"s��2�YYhE����y\��
�>@*b)��*� Ȓr�$U�9�����sg����P�:��!�'���$`�z�r��'.		�=Yx��ݨa^{�v_�eeh��d1��R:����E���V��3�ȵ�Uf��6��疤�~��N觑�P*AX>!�Ӽ�Ti�8�a�,b�	;2��>0`�ս�CXǍ'���lf���mx�a�^&���I��%f��Htn#0��_lVXX��AH:'Q5�Wl��~>��-׆2�'��j"tBh�����VY�����u����;���v�����L
@:�ɾo��^#Uם"���WHGPCO�2���>�yU������X�6��U;(����9�}����j?��'�v*�ORU���'QL��dW�pBP���(��ҵX�OFǊ�نb�4 �	�	6*�p�:;1<�u�4�'���y,�p��y�4f?�:�:\$B�EHEq���ʕ���?�ܡ'�D?��cv��k�V�~LZ
�&{� ������J���Fy���;\�EO�2R\�5 �;���_�w�u���V�MC+�u^��P�R�>8]j�K����9�������St�v�tEc�$�XB�\�k�.�_}4� V#}<l�cWgD3��J�WZ�fC�T� ��[��ŁS��G8��|Ƞl�ʺ��,��~��
)s@5��)��ۉ�rkV��ԔM=�׮��tE^v�*�b�Tg��*̓P|��e�������'ytBV���7�aqa`�{)ڌ�S��kh��X A�r�E�+4�������?���#ȣ �2+^���+otgUS3��@��ԧ�b���{�xX�W����`��'����۔+���d��{�0Tc	OJ���VG�R��tˀ W�Lr���F <����F���$,�b��]ND ��y���|y������-�n=Y����}��!�˘�2��Z<#�
˦CG��8����߹dI�d����[���Rjc����Ew-A:��E��e	v�l_��Ŋs�FѪ{�/��B��m�$��H�N�5=GVJ�`���lp�עx��6����&U(��>J����:$�@����~[�G�L��I+��K�*��+�cCPf��7�j��05����w<&s��!�(�"�2]U�gB��}a�S��7�j��ll9땧e�(��S2��y/��x�����C�����Yz�#�Qx�ȊS���9F�ɝWx �q2
�)��O��X�:��;����xf��ςYE������2��V�RN�˰��3Zb
�s�'1>���ǟB�c��"���;MgK�E9�e��[�,tm��\�p	X�c�p�E� ̳=�(F�a�)��.bhX9�q2г�5$2WKz]��z��%8�V�]���1���,@`g����Nf�V��ج�����\e ��{���e��p;�r{��BF*�KG�z[Ң	��Kh4�����J�D��if��ܶy���+��V̧�\J��h����y��>���D�K�	<,�m=�iV
�p��x���x/jQ���%w.�MG���0A�F�Y�|���C�6G�j$u��[�5�(���?�7� �3��5/Y�ތ1�?�׳��炭��1��>�ܛB����_���G��F��u���hr���d��&̗kH/ʎN�`N�'���_H�p%�L�^dG-��È���.�,ag�گL�vr�q��ETv68���������R.1o!d��3�+_���bW�U�]r��S�(rA 
h3⻶Xv����բ�8��ۂ�sπC��a�y� �;�9�ߔ23�@����I8A	#i���WY�]��bj�z��ջ�ц;���|n�!5�
�|gB+~��R�Q̯��P�}C(pN[��t�(~��.��r?���l\�v�;�Ū��_�W�7A�JB?7�rWh�$H:����W�r�)� �~O9>�^���I�� ���+M���G�Y������Z�P��;&�p �H�:�����X���1��-��'C�������!�����b�B(L��	���V�,T'i2�≂
�N��� ���LS��;?��eY�G5���\�#C9������1�k�g���Y��	���&�QƇ��]/�	|�*��s��p����&<��;˙�z<T���cÈ�C�2�%�hn�@�����P���Z"�|��9�X"���Z�ɇZW�.�uA�8��~�Z�r�[��,�_��O����v�%�8�XQU?���!�䫺�rONE�|�U��#}�����)�&��Վ���#�p�8)>��8*��\E�9	�4Jr3����(&�~���BA}W���8��-Ql�*r� C¶�
s��b'F��K�|/�S�j�{l6��WCrl4ƙ��C̽�m�&�)ax�R��Q�&Q~���R���dZU7憶~%���O|g��^`�@���a�0��8 ���eT Mj'����VƆ`�eǖ�G;��x��0��k����ma43����ȗ������%jV��Y'�<���jԪ5���jc-.�z��{Q8k5������� Q����P{�[�.�����N1��*�����7�-��:�+�Ł�w�Y�?y;�Uƥ�ů,�$��������W:��
F0�TU:;!˭A�,�~Zfv���"'fj����bôA~d�8���¤g.G�į��rՅ��:V8�2��貜�}Y�l���+-�ezta?l�H7�}����ZZ�7�:�n����b�Z;�!۠E"���x&���ęXkk�7�3����_.S2h,Z@�UK{�
�j�L���)j�5 $z�!�W���:��O�V��dP�p���b;Gʥ��Aʯ/��I��)"����k��s��		u�Kڊ�(��փ�%�q��HHQh�}(���Y��=�i5F�����`�M��s�=f�9�\�?A�dv�і��h�0�f�<{�RC��/-�8a�;t�h�9��Il]�'fJ�쉭=�̻:�;._���?Տ����‰���d�Ȉ���]�g/C�xn�DZs
H. �^�]&�6}�bY.�,�LGy���U˸��Lv(���FY��P�
�P��	|u��c[����?���o�?#{}�]�b�1�a��´��諕FV�!��'�H��o�i��7�	��In&�Ԣ
�:;{^T�e�
��m
Y�,�*�\�s�Yٴ�'"�;���w^�~c�M@J	$�x˸�Z8�>���%�OE���q����'&n*�0���J�[4~�^_	�ɛ���/ީ���,�+�5�R����,u0hG����h�����o�9�yx��"�a)��HQ皪�N����x$��̍&��3:͈��]�~� >˒�j������l��lڞ��Y �ϔS>����w@ۢ���hMh��d�</�L��Y�������}
�7����H G%��;�Z�UU������������zN��C[ ���x�����'W�s���!����u���`�+/B��][�X�s��k�~B �.�@�\�SB��;,�˴r>P����_��r����
ތ�&^6a����4�N�\*K\�nP����nl^��T�~>9�<����`52d��2�U0�̡I9:}�����ƭ�ےv[����8�<�k��À���4�Q�����}��(vhj�mvBdk/�� �c�$$v���#����F��ȫw����p
Օ�u�\��/�|��Q��a���1�D;�к��J��>�G�*�ic4T����9F5��[�.6+��a���9j�/!�b'�|�+=z�[Gt�a�	�=8qs��E`A�GB�XG�螟�W�P�[~� Z�K�x�)�HݲX�}q���K�{�{�z���J�BWC����-� (@��a�V���v�d��1��U�t:AD�"��+8־r��⏮N[Ed ��Z��}D�D/� Vu%���͎_�ԍ��(������^t��w�Wm�)���U%��4��T��Q{��:%Z;uU�Aj��,�7�PT#h��ʈ�7�Ff#�3 ;�s���Y�kw��<tȯ��O�rnr�p.xX�M��V�|i9v��P�Q)puy��d��V��/��]���C�C�+�]X�3*��?�)����OG��SOCRa��+�b;��9t�����6B<�B����v��}�F�HSZ{��/���w�ܧφn#0��L'&�� .����Ц��ʤ|�+=�TlZW{�3��/���_�z�����_�o��c����`�G���ˋ�V����s� ���:�0k��ԏ7��*j�96�N$̆���].��`:A>|\__nqPX¿Us$f��2�,�* �Znp"f�m��!6p�pϒťxS����D���:{7E()���R�����2B� x�MiY���^k	�jR�V!��U[-^�3Og!D�+�?әdۿ\����h0W�W��o�	u��c�$Gx�k�p���LBc�O&��!�>$����dH�T��v�5p�����a����1�:��V\;mT��f���5w�O�kWR��jp��4�O���ya�= 'W�	ln�.�i� �TQ�O[�~��x)h���Z<~4����ꅤ0�6|��uR��6�3U��}XS�)d�1.3v%F��`}A-ǚx��2�(���6�KːR!���*�#�1Q��m�[|�|��wq�3W��"�����V� rg<�z���+�~FA�R��,��M�Q�Nn��	�N쪭$�;��fZG�!��E���goc)!�Z�K��$Z�� ��@C�͟����įN������/e������4j,�ط��?t����q
ܡ}�87��'�N�m4F�罃�h�������,��sWu�9B��8A瞭���׮�8���ȝ���;'�hrId�ݭb��ss�s_��$�qsԥ��зw�~��`�ɒ�L.���ԋ����fvl���0�.��q7��E�����N܂�2x�vK@B�l�^�n�`2����[�m��r"N~��:>tW��,*g�f^�q��	uPr��d@��c)���2g
&�H�Zw+XҾ���*c7�Q23��:`�頫����r�)+d�A�j��Q���3��L�N�D�ƻZ8RgU62�+ލd2GNd��$������EM�h�jQ��=��J���-�-��N�&w�@��1St��"(��ɋ��:�q�r{���0s�۝\sq��mg�C��N�e�E�����>�F���l�<'Ro2B)���qG�����/q2s�5l^�I�����,K�t��T2�9R����������{փed�u7��"VF���XJ������;!��.�h$+�8	a<�cH��	[݀�S����l��'��ğ�*��!�Im�#��6��E��O����1ؑ�@pt��O����4�J.�G���j��[� ԑLS}�-���@+�o�Ѡ�ҌBl�6g�IҴ���C���ʺ�	�v�Ǚ<Z^D��UM�5��:~$����>�#H�`���Տ��ۢ	뱚�A�G4�p�l�dS�7D桪�?�Տ���x�5��1}�9���1g*�4&�߅��1�	cr��2:��lrEW�����5u��c+rӞ�B����BE0�M�9��ɤ�����F[�i]2)0/jx;�~꭯)���q��H=�"F����";d��EE��'��������p����K}���'��+N+�и�%���x�+��K"��C'��y��*O.7�w'+\l4�&k!���K�R��n2���b?eZ��!4�!C���'�V (�l�M�(��Uf��R���u�y�g��h\Zk˂��X��1��־@�k |���~����ķt:?��
�j(S1p���.�yќ��xZ�0Q1���շK�r^�ܡL$ổ�<����UE��C�*x�÷�	�����Y�����-�QEu�%�O�1jm]����� ��}<�˧�ދakʷ.��,�;�� �m��#�e�k��mD/m.d�upd@z�罨`��խ�m����5�ܴ���_E�ڥ�����.���k�k 5J"�%���	݃��Pt6ǧWM��$���ۑ>�j���ɇ�4��ȱ����X/B ��k>4�(Q��M�D��pi 

D�F��������{�� �wQj��fN{װ��u��Ĥ��Iu��4�=Ω�&/f����E�_7��x4��5�.c\����T#߸McU��y� ��4�l=���?��tmr�Cj[m䧍.�ULQ�7�S�b�X/��#�af켂�+��Y�N1�,^]X#2�5�Ӕu�f�����<�%e{�Uu��Op%�f�E��ݻ�XU���LL�AtQ/�!���Cq�~t�p�ŕ�^�2u0Q�����SlN�E���P��d�5ƸE��?>����ZXv/����*|��{�1͚|�Ӳ|��k6��քx�%���y����Lk�(PN�l&���΋���+o))�4@�as�i��Ja�fx ��cq��A�'D���ET��o +.O�sok�Q����A�\�&{5��������c�ũ��5V���W��d�������x���y=�$1�3�7pC?_j	)	ώ�C�����YU��f�U �W����J�z
�����i�ܹ3m��nM�F:�A+��*Fu$HE���ډ͡'%��i1�-�x�pPµ�&�l*jOӊV�������]��H$��Q�ł^&T��9i���<I�$�m@��q`��� �+���D���(����B�[4��U�b^�^uJ�&�ؿz��}gί@��sr��v��5X�/4�"��R��x~��=�/|<��m]#.8����Eq!~�D�'�Ri0e��L)pi�owY646�yk�� ɛ���U0&�@���jW`	v�~ �N���Ί�-)�F``9�����?g��1��Ex��0Zr���*��1a��4�ܖ<v1	|O�0�O�QB�,�2p��/���v��u��@�Q�ن���T���3�ە����AeY)����e;�`q�5�wr�-ۈ�.DX⊗�F�ep{)?���5{'�[�Yv��7�.�����b}���#�GC��ǩ�[v9d�7~j��L��eb�ȦGβ�s]�(,bh]�Qu�	O�+׺o���(�Vu����G�Tc��/`�z=�6m��xP���Էw_
Z�v+؆�n%4�q�X�]et��ap&��<�u-�[��������ҧ:���,��"�&�}9�$�r�h)mϲT��D��ƺ� ��r����m��a�[�zofN����܃i}7�j�l�ד�@*s.趁5�b`�7̖����OZZ�����9��R�O�Q��2�u��}��ۛ�c����,�ݒ�A�7�}[�"�����| ���,�٧1��<�_{���%q�3Ι��7���o���LJ_x��y#�'��E�Vv�`)���YaC����]8Y�Mvq�G0&�y�!�?��dMf3����Q4�/�N��˫h_���0�Tُ��
v!���V��B��c�trJ3r��і�\�T"��8�]�:���������sR1����~I�6���oK�i.��$�����E@�Sr���"
���h��s��+��;K��Oe�ܚ�zI�{���v��<��"���\琱{އE��iı�O��<)�r�.��]	�-��M`��/���DL@ݝ�-�/�����Q�D_���{���F���X@��_���#�]Q�5/<�d��KHi��^$Cu���v/捪���?���	9�~ؘ*��i�(������0��������1]+p˙�����d�E֬wҘ��[�~�Rfx4}���g�۶?
Y��T^Ǩ�t�9��Q�Z���i�� �Sv��M�������er��
�0��	LU��%��E�Dr��&��2'��Q�ߨR���#�Tc��;Ч��]·Z���ɗ��n��s|T��Cj���r
�i�%��������(��c�_�u�v���rF9�f"�%�%�Q�أX� /��n�UVu�%a*��n9�~^ 7U�I*�5�Г<�p����fª� W�	X��F�qЦ�߻�#�/y�Ų�J6=B���>|���?�M��!��1�h�3�Sh?�>þ� ����
R-���q��������O�U&cT�>-x|CC���It�U�?]�Ã�#�=ѱ���v�_j-��2�ּ���YG��~dʬI����.�l�o���}�Y.�w⺥��Υ���e�j#��)P~z�h��K>6q�  ��<�n�N5�yhx�O�rZ�u����g���.h-T"vd����],�CX�E@��F���	�]�U8���]�f�|���!d*v[eBoH(.AH� ��iv+�4<^O~rj�0x_��$��ܨ ����`��C\�?7~���."�1��ɉ��Z,�Ì8��|�KJM;~�&��^"�$���W҃��;��a��s����<3���(J�"�}�)y���o��o�����.58`�ֽLQr'otI�G{~+���*�$�ۣ�5��<��6�0#��']�	�D)YQ·`E�����x
�g�[V^���F�4 ��A	�`�_���hj��AQP��*�[���c��a��,6;��1����� �w� �
�d�������0-��V�W���\y�����H7 ׭��_�0Vo W˫� �F�7����*�T�G��ޮ�	��=cB��@0v�c�~E[0��V�����12*[B%A�Zh�v.����%9Zk3Q���.
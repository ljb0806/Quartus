��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y���U� �ܮ(a�����=t��n�P��L��q�\�����
nZ?v�^N��bYJ�3�e�9�<[ey)�Qy� �Ƶg��> nuܮgש���F;���F�Ή[����wQB�ȯ'T�u�U��M�pI3,7��E�k���m��~��n	�D䳻�	V=v���e�X��k���#��6��%z
���U�L��%�����	��K�	�{gg��yE�*]�ݽ1C�7�>�T��H�I��1�.+g�4jTl�D�6pX��9.�
��%�Q�m���$?�Dc8�v(05�?M
QV��Ce@���/;��1oMwhgU��+X�{C���{��厊��(��$Ds��d�떦@��|K��G�5 ǪH3�cWL��ռ��I����ʸe<7�x�]������3�����w���L�@qi��wJ�vo�=T߬��5��0˜$۳;t�|��p�� ��m������F Ҫ�}��9M��4Q��L�H]9Ѡ��8m$�S$�w�5U7#��	����0p���zj��Y��5�С�c@`���8�͈��N='��M\��U��BE:u����qf�`�ڎ��&z5^�t.�w3�O ������{�e�W����Et��4c�z)�/\������#lv��B
hFքE� z߹-���ݔ>��	FSvY�m�E���9D�c�S�<�}�覑o�/@vC��`FF'=N&]xr����a��w�7�4���a��3���a|�p���3�G�z�:�E�s��D:3�ٰ�<rŁp��m��5����w�b�%�}�:y��Cc�u���mbt�=��#+�F��]�L�^ t3I�a�Ņ�[A�aB��3
�����#$��O�o��p=G}z'�l1>�����3ؚċ�iUO��|��_�M�%ǩ�Ǐ��-�ý���*��(��iVT�2{�x.^N!��3I���!,�O)4�JJΜ�ݐ��K�$��*
��
U|�
�D��vhi{��(xT;swV�)�6SA+�ݾ������}@�h�)����e���Y�\Z��٘��l,Ǌ�͢�N��5�#ͧ�0w���#�{��VlA �q��Z���_I6�z���}5���ZY�u�9� �H �$�l�Z��L���������`bܪ?þ�`L-� �3����٣%�Qb���O[=PcU؝ZU�������t|BU���㼘GH�u���jh[p3��|N�C� ���$�W�$0�!�,1_�`�
4e�������|��󣼂pWb��j~�/�:t���6 U�K�:"� BY�1POm�@J��"���}ִH�%��e㔇�͹�a$O���J!0��I�a���)*���3��Ƃ����2	y��*��Ob6����w���b�x��?�Ý����ZV�@Po,�/@,f�/E�x��O�V��2��+;h��hf��	Q�h�a��Fc�uk̄Q1N�ur]��O0���k� +�����#%��j�ә�E|���6��������]�$4��H�8�c�`C��g�U���TY^9���LO�T)c�����p׺���{�}�jԅ��_� ����s��3k�/6r���E`l�&��
��V��Ơ^Ժ��tEP�\�|]��Z���ѧ��_;r�z�c�X�y+��Aw{��d��� ���4���O!���+��xl�\J㪂�bn���C(��ι��{"�)�5n﵄&��x
��3d���t�+��`Ǻ`���j���<NM��c[e0xX�ݟ� �Z�ei�'���8`:�3���ĕ=9�?JJ��Ƶ5A ޅ7A5��T؋��g�Eo�]�X��ݸL�0؊�&Ej콉�.
���[�)؄��7;�!�)8�~�{�D�#c��_G�É���Nc��"吘0��u@�%�$_��E������0��a�͉�?�%=w��*�l��ntw"�OZ	i��4�!�`���`'3
�������1?��Z��;�_��S΀x^�o�nUf�K��"L<,���G��GJ���wô�K@�T,i)B]���G���5��s�]��*�d����~�Y�]���os��sq ��(��>uf�%�(�����q�߉����2Et��e!/�I�lW�$�˹@<���Lh�C0ZZ�(83!�1�1�A��*�֣6��Qp_�d�!���~��<�f�{�hŉ\��.��<�C��I	����?K�)Ý&�0��t�B���aEf�j��/�5/�Q�=
�
'Q��J��i�;��=g���n��'���LSj�ؽ>&FR�j#��_B��$��8�D4�lYZ"F����Q�"�tt<M�b�D�υ,�(�(��T�D�G>�`�u��A�Ql{8+1�iK?��²�t�z�q����av�6��Z���q��t�I�~�:�.�p�����[�3�t�̥�Ώ)�!0H�iγ`ߪn�#�,P�,�+]�EgY,:)V,�r��޻H� y����&e^bR=� u��-Fқ9E�.a��G��\���UyZi�����r�D �ѣ-0�GG5��G�}�1>8�ʔ˔��G ��O�z��Ǯ�y�t�ɱ��� `������ST�7ϖƽQ��>v"�"M(N�^سN\�*\���k馤�dh�O�L$�S���R��8�	�X�7пǂ<�Ws-�Y��H���Y��T��y���>��wM��	%�ٟ.$-� �x��b$�z��3��`F@xSRTZė�9_X>Y�->�K�D�E�=�N��SeUזM��?}��-��=On�{�6f��[m����G2�B&�v���9���rL��.�FB�����),��� �Zs�Z-~�͠����"ؿ��,X+��t�o.*�=m��@cf�8`��J2��za�w�E{3�\�p��a����&56ΐb�lօ�I�m��wJ׌�&��/~�ce	_�����g2�R���+��۵�ެb2\�{�p��8�5�ך�z]�q��b�L�����8=ٔ����^���]��,t�913�#֦S��XEq� Ǒ;v�ǉ�a�&�o�/����=���������Q|_U������K!�DƧ&�q����F9�W�[%3��k3ﰮ��w������}Q�d�(8%xJ�X~�(6������'���J���<�fV�]E��x�g��I�R�T��`�#'	!���:R�o��h鍬vzs�-��5�-j�FSږY�)/���Y�EV)e6X��y/�E�1@#H-����6�Ǒ�q������w�����w�Z@L��	���G�6��'EU�c:A���4���� ����	;�=C�Hb����L[hg��ln���� l,&���fZ؇�;Kt���D�6/PE�Z��k[n��_��/hV���� �U���h��Uv��m�����Dê<,���x���?:�o�K�	H�]t���jk��l��S$
�~�w�%�9In���[?ă����r�o���K��b���d/+�����%�U��CǤ����0�9'��KI�ȍ?l�ץr�N!�[$J�Q*2����q7D �ڽ/�p�\��0[V�d�0����*RAbM��}��V��׮���޵�p�����r��$�ϼw�Ny\Y����=���c�0o�u��^�0��Rs_�k�)#�&��[�ȫ����(�6�Y=�,B}��D�[?}���a!�<�,�L䔷�Z�F�! �2A�i�Y�xC��Y$���瓔���ʣ�ĸ�b9�}�G�A���l��8�!��.W�t P;9,;hx�N
��v�֋Pxet���ؤT�>b��ۑ�:�W-�Z��r�5Q$�1G&ݟ����rI|�Н���o�z��#��8<�FP��1@hOPk�W�匃9��<n7���%��B�)�ߎLD`)yA2�S�~9�d�����Q�KUX6���Nh,3��څptrY�N���
?T1����+��,h�1ԍ�]�uN���#{gL�Z�o���e`�5=�6���ɾ�_S^\��|�����v+�hI'@�n�|��_����g��P�ے����7�k
���W�H�(t6r���4[��Y>��v�х�r�� ���J�_�L�K���y��vK�[�MK�~I"�ZU6�j?����B�<!S(�$��;�,lm�7�i�s��mb�_sQ��М��L�]57��s�aZ�Sl&����6��n�;u�G�O�ё���{���8���槸Ao���2,�IT��A��Y&��� �ƮU��6ow��F��N��+L��&2�)aƤ�����|�:��P����gLM%0<��x�����A�S+7��LJ���v��H!Z�G&#�Wt�t��Yq�n�4��b��S�A�qT�fj�$[�`��q`�XD��������9Kd��1��+� ���P�������cä����Q�5WL������c�x��)g>F�"64N|}�S<@���f�r�5XT�).��{r y��&�����n��kg��'㥁҆�G�����\��NT-n��C���~��B�xj"k��a�L��"���B�)�r~���E�kϜo�|�6�ˑ޾ɞS������2|3A-�ߨD���l^¥y@�CG����t����蹳���z<:����ck~��L�]S	\��J�je�X�R	_���,R��W�s�'/p��	`sl�t]� 08(�N
q����oC�"+��%�M}��)���>��/�z���k�l�z��C�� Y���Ȓ<�c��F�]�I�;䪀G��$jc��Ǎ���niݕP��HK����4�`��b��e�\rL��&�lO�Ov4S!��`$%��#]v�ki��0�]��χy��L3�!���X/.�	��IEi��.�6&0��c5!�i���z$�=�~Y1�[7q�"�l��c�H�`$��QD/7�~���2�13�x�W.Z<I�a����YDwF�cD�୶h-��u��Ľ^�:���Ӈv�a�<il��⽑o��P}��x�(�ɓB�9�UxAS��Xn>���j�?�U�=8�>&?�|���7�bk�һ�H�1S��Pg�d|r��9q��5��"�5�(6�%U
���'F�vMl<��D&���J��i(�&�C�C���|V�n��}��ܣ�]�U���ZqWw�s����D�5)���,���	;���H��Xe����]4b�������ʄB�*AX��K9?�?VНh�U@_dͳ�Q@�c�I��0���n����cBf-n��2��wҌ*�,�'�6��=��X8 ��`�݁��?Ž~$�Fr1�[��.��\7-^�P�Y*��-+*E> �
�*.`ɨ�M�t��~HEEא�7Fho�����L��P�Ó�5ٶ�i�bx��VP�Uyݔ&9�����n+z/^�F\s��m��GcJ���^G}b���XE���� �>��B�O&DW���u���������w˘i�������W!xKA�-����m�p�W����Л��_E�캏�� ��pi��agm��8.���x�h�e��,�Iq"nj�Θn����Y �IY�g�.���8}SHy��H��瞳�g�_su�=Ŗ�iT�q�&�q��m8����-�����WA,������: Y�E���]-�k=�m��J~��j4$W lqP�C]�+��@v�(p��`3�:�h�C1Nfw�,Pa��e�#��Ì�R�P���Ada�&L*�K/N<�Ek�v��NZ��}��)"�4u.F��U���'3���[��j@.�cg�%E�<8a=2��iڨm���N��,.x9�B�Y(<<k�Wd��:0�{�2V~���y�TϽ���R�!x:E�{��ѓ,�h5&�I}�ʡ@ȯ��. ]�g����J��[xt,��!�4^u���
�^<(p�/&7���}Y�_U��1����������a��x��S{-7�%�D��XLD�7��e���e���(�r+�_��u�vǼ��Q�������ɀ"Jy����{"�p��� -ğ��}�FX�� "��"���d�����q�s�{��rЇn��-�.��!���H�/Q���PjM��!��H��D�B���� �i�[�f��g�m%Ӯ97� �o�ƭǚ�`�}��$o77�g Q�v���\��ˇ�'��ڔF�g�Yc�]��P�� w�baf��]��\���`*���܏�/��Vd�����_�}���]w4�+��'|�]�GbR�z��K.]���@��PHҿ�p���݋;]��c�"�_��w�&H����Ԥ�?�v<��hR�N��QB�M�mc�vd������yEW��zk�	F,6&�ք2&z��X����z��eK��-E��|�c��1��3/&�܈t\X�a�؀[�o�d�� P2��A5j����B��m�QSV5�::B��'q�K�Τ����731��A5rJo;��`{�l	�4��=7�N�����6�K4��ɬ��m�@ jǂ�ݥ^�L�]��V��\�������({�~h��JtOXH��Ig���X�̍����b�9�a�� �֛8)y��LQ�F`�6�su��í��d�\�C���fu� ��uhP1�S"t	!R����Ҷa��ީ�,�`2�]�����ShN�Ꮾ�s��J�ȭ�@��>����$�M��f�h}��(2��Վps[���{�������#+�@�L��īu'Ϧ�u�)=�!�����������b=h��u�H�Y:=T�NI!�bC��<�ꕃ!�K������]�YRXBФ!���YKY���=�.z��T�� ��Hd��
�A��l�<�u�Q_c+����`��:��z��W�|T�Vy60`�d�=���e��Θ��.wIscA�|�"[�Zt�ӷ����_Yӄ�CxNc�:F �S��e6hU�Z?ʧ������V&z���jH:Hq+��\���gf{u�g(.�f�S�U]@&���A{��db��Y7;�@ �	٭�rC�,��IE~�)�s�W7ش.���*��:�o�=�vz�![�[s��׊>�9@��E	i��0ڎ��U/�����l)Fy�B��EC���)�:{J��o(��w
�Q��^�Q����t�>�C���������e�V��(3ж֠ght�~�H`PP���Q�Ab�wj����]�Ӹ)i�МYb���C����/s�X/�Td�Oo�VN-˸�7�����Nʐ�"=i���,4�Z�r+�Y@���'3���.Ɯ7�خ��M��o,Ǉmj3ï���X]|�c���#$D!��P�*剽;Ӛk���9(�3TL$�L��׫@?��Y��
��
���O�z��շu�i@Bj}Em�y���/��[<f@}�՘*����pQw~���#*��r���}�ǫ�'�,z�SmT���&%�e��\�o37�3�|H�����J��a�o��C�NfL��顗?;���3����Ua�R@/�,]�HX>xL>��S�p����ŀ��<X�$��x�u��n���Fę���Y�[)9�J�|�l���W���-��&�X��%�2��9�|���G�_5�R[�Û:�}�{�]��B?&�۾k>���sf$�gq�y`��Uܫf[S	������T9u9Ʃ0���ƻ���B�S����`���ĳ�XZMŀ�7�]�WP�b�!��u�C��\hε�H���no�b- ��tKI��t��]Ks�w\X�D��q�ư)���GK`����A�e�	��x^+���9�>kJB.s��ub���v��]ʼ@P<�]��&�U7��ߜ���Ecl*�I~>z.5,���e�Z���D0�x�?�ǺZ���~�F?�fk�o�O.�/�zcK$����bQZ7jK�/���s�0K[�E#6�ACn6(��e�Ԫa���6몣�fR���m|�*[�F�̸>�e~�чz�,4�2Ղ �L/���$3-���=�:�\��7�[V@!��+y�ԁ�����9�X�7���:��#��	�|�=L֩ W�j��U5�l����c���6dj�g=NK�wD���^kVX|T3X�&�[�w��t冀�U�h�:����lA��5�IIQ ՆSɦU��95��s��ѩ:m�ˇ�4�j<8���'y!�Ho��[X�n{��B�[�M$\X4��6:�>_��;�S[�Yg ���嘵�U]գ�im����_���D��9b**"yX��3���Ȇ�PS�Db[��%��$�t��H���f����$. �' ��)�v������
O��%*̥}���qyP����,�`���5��2N����?��� �'��@`��Ar<��+�i�oI����!C2u�/6K��cjT�xl!%� $�,�[$Y���n���� �����8uo8�*?�'��YzGJux	8�?.ǎ�|8��3u�ߚS�f�U�G[�	C��M h'��� "5C��q�Y¨��}�$ҭ�@�0bw�nh��/�Z��Y���Ru��v�eQ�R����8�?vzT���?�S-�W�ʚʵ��.?��jB%�~��^��1,R��L�C�H#?�3�ЬZ

gY�Gx�P�]WG�%����J�P�u�(5��g�8�9���u�����!�K��廉.7���[FA��@6�'$C��@~[ܝ�� f���� X�V��*�/;�g�s�2JQFe��CP�.��n Z9��]�P�j��'eS��Q4&��"9j�I�Ģƍ�6��;y�m��<��)�Ӕ����>�C��#��t�p�#�f�#:;�f܀�:m�Y��z���ܠd[�M�<�-io�ՠy p&�$C�h����R�˛��ϟc�%%jq�ezPL3��X�8�p_�&"W5��o"�҈�*@�vRs�lA�򹆻�!LkӕǬP�J��%����"�����DT�gRm��$��$k�q����15����_��|酺͎3���"������J�lE-���
����ޟ�e�}��W��T�GC�|<8@��lӢ�vT�[`98�B�|,S�����;�,�l����S�q媂�����;���9�H�<�ག� ��e	�a-�*-˔���w:{�;�#"bU����@rY��s�2�.TqC �lz0�h�H�>!pc�����x�SkLg2/��]�2�L��Y
;q�t4��G�B�!��*vc��St5j~�H`�]Z��I$��$��t37��u���@�m��k�k�so��v��+���C��@ݒJ2�o����ՠ�j(oC�Ne�Y�^���(��U1�a1��]J(��q����Ԍ�� �����J����tp2 T�$#�rM��|�r��JuV�������a�)��ؓ}MÅF�X�4	�8���j�dS��r�.=Mc��8�����ĸ�Q���,� (;�Ng�ʻ���0��H�*�9�^�$�R������C�r�G�9�~%�E����FBM�E�]9n�T��&���X�j$t��4�-����S@�����TNm׶(�����G�-�<����e��S�`��	�E���mg7\���F�	I/�y]��^WO�쫆:�끗��������5�\�3o ��W��8s"50���K�Ǹ��&�wK�6u��+�ͳ@��h6�}����� '6����#`���%��hC�&��s�s�mb-Djє�ϔ�8�ݲ��f>Y�Љ>�4W�-�x�H���M���8]_;��C��aK"HZA��8��+�(.-��e����X6�¼1t���!���Q؍N����׳��2|��W�"  e���3Y%˗Y
�#�r2���p����'y�.f IA@r�%#�^c�����.������&�|v5�
rM0`�jSPoڝ1�ђ=��ؿ�}ϊ�Q���p�puO����Nї���+����q���{m:��$!C*��Xk �G"��D2)�ɰO	������V��.�� 	m���T�/��_���J[�PǊ���a��X�."&��A!��q�U�锶�
�-/���1����~ �3���V&ѢD���o�����T��m��?Hܹ��t.�(V>d�E�n8�F�v�a����r�Q�C���^�0�jQ�u8�a�����~�9�/�N>~�F�n!���珗 ���QZu�����^C1��#�6�ؙT��✶�C_#Q��s|���_�o��Sv'<��/��֬E#�q�ǟ�[;Wr��ӿ�Hvb�L�5�743;Bq����Eﬨ�����X�˔�)��o���q�b��/F�E#�����ky�p��/�\v!�x�Q��N>r|V�I5�<��n��HF���Dr\Pw�@qY��$���U������� �$��G_�76h�۰a
o� ү[�-b���^xл\�Áu�*$�f��E��lA�,�mx�ı�{�D���Q�7.�~���m�jڋ�y�{�\�U���v�m�1{y��u���L����B ^̔q�dXܡ�V�]���w����h��,�^�T[�7H�&f�w��,�库И"LA��;+��R�� Wn0�I�:�l���K^.)���?��$�<��",Ku!�E#ތ�H�e2tL���������f�)<�u�d��jw�5�m2�i���R�_g8��*
����+b��?�s���$�Uf#J���=r�u�6�٧0=���`{w�㬑��P�F�2V�j��P>�';���lu��"%��~�1V1Գ�
	,i�%��p�\�>�D�8 ��`�>��t'�l{�����^��	�a��	Q�G�K�4��fw�]��<*�� !_ʍ�YP6���ٟ��t�~G�D:�SQo$�A�y���
���/&�3����'Y�2�)b6��T$cFf��i�d�bqv��1���K��7ㇾ�Xx�������Zs��mgq���ۖj���oY,�*x1$�Ǩ4�  �p����u�#����kwF�G@�F� �}vO6rbM�-\q���p(�����]:h�����h>��v&���»�����wY����[�� �}�fAʦ��܃������������{���>�f�ߊ�S�1Y�sH����>�-���.��(��ܽ��$�)�m2��D��笜n���;P;̓��	�Y/��4�\`x��5Ա��/\�aU*�1���#L+����I!�~q@�-3&Vs��q)B^a��U�G�%�G�� �w�@��Э�w�B�$��q� 鯭X��$��	�O� ��K��X�oR1����.+��BE�f��N#O	'�b[�T�8��|td��KLR��N�5���{|2i�9Qs?]FO���t�,�U����D|�a���v#��u,ut��3A)0}�PjJ��6͖G������"��[��m���]�XZXN�Y���jR�v}/��'��7'��O�ȟ�O]���qݓ�u�.0c�< ��֮z�qb��'���c�j�%�=ԅөUEp.�\�H�-�9sL❌�r3���Eg�8	.[At	C�m�n�����dGA�Q(r���v��̓�dA{K��>�U����8)��|��p�TA�"\��ԇ�ƍ�$��밈�Ab���d�h�!���E[�8vK&4Ԛ�!�hҘ�<4`��c�򀐽�r����`'l�>}g伪Ld�C�*)�ƹS!��z��2�ӈZȼ��βmĊsw��O�|��F�[��ft��	0-�a��03���3�����{ʬ������!�"fL�l�;�Pkd	c��K�,d���n�!���OG]�^!c���a���\� r9@N������k�p���><�,u����@	Ɂ�3�R�(�Vo�O�w�C�=t�/��d	v���{��M�`w�>��?>��\z�p��o��-�_T���K�n��\��lg��MjRs��p�6�s�xՊO��y�O�s�	&>SAC����{��#�w��l�c%:,��P��z�Y4�1��:�Dx����u�J-�=N�q�N�U����N���Y8��j%�B�gU��7����5�z<Dl���I?��pT�]Rk�f�а�J��ܥ�	�����*�`;���ޅ��X[T�@�IoK.���s}{���OD�h�]z�'���#��p��a=,5���zT���I0�e�h��
Mʀ3n��6�Xf~�<�Un���5@�.�-���t��%@�J�ـ���O�3C����Z�4_Ύ�R�W�5*�4�S��9D��йb
��^��r���W�L�vQ�1r�#�*��C ��N�������"�}^�z��d�60��30Iu�'�c2�Q�<�]&��f3���C�O����0Y��UϺ�F�eZ�b8�c�Dww�S�#f�>#[�ہ"��HB�B�Ǎt���(S90Ba~#������E'�9�$�Bom9ڻ�[	�PAC��HRZ%)gGx��ݬ���A͋�u����8m�5����6n#	�NEu�.R����/9��AG��E�Y-���\�G4�	�ޛm
V>�㍧���7lWx1�ap�7#G��#�������e+!���tt�>�[
����+�o����R� ��	M���k��tJ67
��V�wf_�ڭ�e�%���3Xǘ�98��� K3o�f���]+"�J�&��l�_�EM�mX�VO���a�~јNdWg2֓���]�q�ܥi�,O���/Xd�1~*)��WD�>���y���[��W�����}�N�u;����L�Y�wn'���g��	7\�
��
R��J����(����sQeF��O����۪2�Z��!m@�(�ު�I5��VM`�a��;�X蘃WN�O�r@�Gm
� �N�w���T�����ݜ�'1> |#>$<��;�
9ɀ2�Dl?2�S�ǩ��������p
�4�ĸ)�7#���Q��跢��:Ӹ�ۅo�&��й�(a����.��]��*�.�I��,���p��%3еaYrw��"���&s�,Ζ�<qZ�|��aX��b����AHd�>�H�UO�j�}H/�Ñ������G[91Fh���E@�K��wQ��-Q�a��[�9�9���x�w$�^�:��Q��sf�E�_����NO����qRaW"�M�:֍������i����QV3�
#B��t,r,�Ы�ePX��^`t�ð29Ӵ�E����׀��K,�Q�^K6n6&G�ַ6l"M��o]�j�̌uuHcWz���h�0�/ EiO$NS�c�>,�RLW嚞�v�h�������e�lė�LZ6֛��f*2;��00l~��*PXN)I�-�@Z�h�G�o�a$�g,^ �8�lq����;'�ީ"ܾ��������Q�+�9��>�^V��d�6*Dۉ6���m9A������j@�Y�3Q�=�*7��+�H��K��H��^݅��a��+K��Af���l�w0u�4u5���6��:u�&㎀v_?�٫9|��F�ћM�<	�Ȅ��,�i~��HĚ�"�s�&Ey���;�03�G-\�{dl�N��8��C��Q���4�������0�F5���Bz�;EWp50�ƭ�戢����y�v�Oh�+�p�����<� z�&iG dV��]/��:��x~�A�E��O�8`�?��bC��3��fK�����˱�yx,ũ�YL
��Tq7��]l{��!�&�,!�g�/C荟�2$+'}�r��O�#�^�F�����O8���2��{c�8o�̳G������a	�.8�S5��D̳��D@uu���cb�=Ĕ�����~`߶����{Y�h6l�x�C\WV�/����	�7���Aԓ����f!<&~Q\{���:v�i�.&����2�6��Üt�o�t�� � �k�ꊧ�oV#K�V���A��>�w?��"CΨ�s������� �e�TK\0�s,΃��ށBm��`x�iZ�ן!�fO�ldi5oNW�`�a��`����?���]
�8���A�I��G��6�p�(�XvU��wZ�@��.4�V��vb��?P���:�f�r��'�rFi�|'��qC&�Fd��/!��:m����-o�3r�c��YuZ�ߟS��^gV�>�-_]����0��@#���-~y�������t���OHr2&�X�>t[�����j�)ED) {_D�k�s*��Z�Jl.�.�7K򏯎X�$D�	U��	��i�4�4s�Ͷq����������|�V_m��aIy`i��C�к���"(6,��U������ԟ��v�ɹ� ���x��ᛀ%���v#1�-�[�a�r�S^$E��Ԗ��.� �A�W��Y�&�#όTҕT�T�HY}]�ҨR�9)��N��f�x�MQ�[�6�|Y�svŘ�Z�1��)F�N�@�:�w)���������b��FM�<����v*�bK�a*�َ"�����ꛚ%�<8��h1MC:�7eF���H�t�0hJ������ka�S|/��x�4����m�h(-��1�x$�D�.a�Z�-r�ǳ�z&�'K&��s�P�8�z��F��YуA�"��\{���JH�"��plsy�֞�>sSA���'�P����5=��e.����9�	`ē3;�������^���Y�&l˖�u��Ȥ�, �P�$92Q�
)���ޣ㔌�Ц�T̿P?f,�����7�Hp���Nh�af^�u�,�t3�?��7h�������������zڗ���=y����(}�����}t�E�����3Y>�|,04�����`�\%���^>\�/���78*Y"L_>O�ӷ�kĿ�w�"T���x�AGom�k�E}	�T������MS���nbpiO�s��b쵠���t���<ښ��Gº���R�c+��!�@+���4D��u�S���mӌ�1]GʠL�)���B�}�:��imo�Ė����>����C���XK8�������#�>p�5WD�(/)FrQ�����-?܄K~��y^k��'�q>eLo��%�ɂ,� �Vb�=z ��.��;D�$K� �!�V2�Eը�}����9��a�N0���v9V��L�-��,ݜ N�ǌ�q������{dF�7���gI��p��\(���W�hԝ��w�[guPm�_j������py*�2q���B�"�(E�xx�qZ\��`�����ZU�ō�N��u�F}�Ej����u��0O	f�OhbT-Ƣm��E|延9^�ZB��՞,��]����,7r%K h��KlW{vͱ��eP�	�п�Κ�V0v*&��?���a�U��,�_⇶?.&�Po��N_^t&8(�nK��NJ�_M��Y���MY�Pk��mT��L�>�����b)g�PD�0F��91+���m>�𵪎IbE�sI<_8��Ў ��p*�Is' O�5��S�\Z��Ƥ����3/q���`�>����f�$8y����ׅ�N�`��98T\�����rcIT�F%72�ޡ��<�Ѧ�ТA{Y;�n������Vߴ�������jw�h��[{[u�U��0���7�K�������*rZ!�{
��,�Pnݣ+�
cX�-�u����.Qb9,X�r�N��iQ�~b7�.�ֵ	݀�^�����?���M)��}zEm\���5
�z��p@ӄE�m �^|�h�?���&�Q�o���x�aGl~��]9i��-���qOڞ?o�K�+rO����9�Xk�\%�V���V�ɜ�S�)�D������3�-S��4՚3(�-�D�w4��♑�r�t��~0"�0�����}����M��f�]
lp�F�o��T�Џ� 5�S�]zυĽ����A5C�O��=�
e�Y81E�Gy������R=�O�:`���J&(LQ��
\ �V�k�/��uT��x'����e�:�[a&A��j�r��<B��	ou��CȊ'Z�!--�'�x�"&{빌�yVox�z��kV�>If���\H���`"�"ucU�9C����U�7���o��UdD��v0/?�L4}��A|K1�|�b�f<A3:�;��[��ƌN�7�--21�{G��#	6���-!��Rަ�Rv��Y��g�b��Bƹ���j��p����sd�;~����״MaT^����'ó�R'E�O�Sk#�K�\ˁM����"���%ٟߊK��k]
���0��W8�0����H��s� n��ؒ�)9�R���J5<_@Šn�ɠ7|�&Np�M�u@Ԯ �w�	&�Ƿ)~0d�z aA���O��/5�SH����X���,}�a��CD�hJ�ҷ�
C����^�]�|�,���'2B�q�]�Tq���6�����ԔV��������y������%�)�p��s��Ɖ�RNgܬA3��ʟ�i�r�&ֆ�ag(Hĺ���U�3�N�k�� ߎ�q���%�ܯJ|�M�*�Zԏ�Iv̼�Y����h3�Ss�C��������#Q;�G}%�m*lt$,���������i���^�W����A�����t��&��K��9���E�iT�T��i�Vnll�^���Yq�i{҃�RB��փ�H}(;ۡ)�RO{����D8dhX~-	�rb�&YP'�~�ڒM��]��:\E�������p������w&��m�ky���.�I�������IV���ra�+�%}s���M�-׌S�p- J�S6K=�;����%�Y���7� ��,\���Zn�33�,/Qފ)
ۡK���x��5)����Go�j�/��9{"��T�q����(�'t�ٙ����-x`�H1q\e�k�h��dK�e|@�Է��FoL��R�x2S/�v-F��T��UQ%45&>@����o�(��KO)0�;���j�e.�z�Gk-���tt��6W�^����FL����&{\yo��)/��1���}\D��=I�P����^WqO�$彐g���M�AR��.v��VK��bl���9��������t 5b��Jqv��z�H��[��e���v�$ҊbZzŦw	i�b��)0��4P�����F�)|ܽ;Xy�(`h��}a���J��o:��r?yO~��@U�:q�.?̺�a��,�O}Ϟ�+U�O:7"�#�m��"�qu��5���	9�O��׽%y0N�}�Y!S�m@�k&:$[�ǡc"6�:���&{T���	i΀�F�[�uU@��@�?�_VoZ?���=ρ��$���	,k7wm���O�}�_t��+(�oDaк�s6�Ģ�w�p��TF�|��K�G���~3��-9�i�����QU��B�n��7�P�rq%�`E1�n�:Y�B⧡ː1����h�u���hT�'�ZE+�̊��2N�����|b#�<�;��c);�k6�Q��h_J����b��1�|�n5FbHBp=+T����]v����v��cyd1O�U��<tՂ$���T.zĨ=�K�V���=����#~��s#��u�$ki4�.ǜ��E*���y����굓��;��OpL�4��9#���==ɍH���x��g{�!���|}$iل ~ᕾ�>b� n�ջ�I��������p��4����.�R�o���KB�e��8�c�6�n^�
q�8�t��ja;&��U�q8�}��j�,����I�4�:��N���"N#�R�$`d}	�X4{����,5�'W]M��� -�a�[-����)���IR��
x�ڶ��(N��i�(�c���
m8��M�&�_&z|F*i����gGpdeh�;�La&��K%�*+�W�n莓�)A֡�̘�c�5WÁŬ�II�m����G�{:�Ğ��ɢ�U��&��4d�Kweݤ{��IB��`Ea�
��"6v����~�A&;�_����dQ��1F�S�
�$��=`\����!��ު�]kN]���cէ�c�tweL���˺W4���)��i*����~�?H	ѡK�A��5�=1�J-*��|䚇�t"q�.i�����#;�1#/0��P/����J4�ʠ�kr%��(b�/ޏ�~��%2��c��I>��@�5)b�� �ԋ�����.�%XzՉ���"M �}DÐ��zG���uHtS�f;�k���:b_��l�^$�C.q�P���փR�����نS*9gW!�@���i��kn��F�X^	�/�)�^��GWt7*�&�RW��"��q��nr8��S��#Q���� �<�io�K%�����ŉQ[\��M�n��t�>������ki�s
��A��D4�/���>��ѵ���ڠu�	C�a�FX$��˳���!.��M,�ُ�}�8�\o��pQ�;����<{��$N���=sϢ��zX��z��,~�;[P|�ɏGY���MwR�V��rp���G�%>��R�f���s���� [_XĨg�1�;Ly�;�<{�;�@��,���T*&I���~r����e��$É�41]�@�O��,�f�{��x�cm���0ӯ���Rc���u2�v
����.@=]��jt���pC8gf��b�}<|��&
@_C\�*g+��3Ȩ�B��>
>�+�8~�9��ܨβK��V����>8���~�!q TE����T#��D+>�vA�����Z�so�\
nU�)��I�o̠��@����ȹ���Y�?�΂�:�2��{��.\�ii$���g/�m�	&�iR-:�avR�I���	F��͞jGj ��e�wsug�^/��m5�5����=G����f"�h�zWE�F�;�HB����Vd��τ�q�lI	zL	��!��j���IU� �t�e>[�^D(齮�;�G��Hf���?9�	q��]���"��T;��dWi	^�&q�c98��cdj	�Y4�A{���Q}�I.bE� �;w�/���

ֿ�^������fA���n���5j�	A���+�׽��3�����nS�2ê�*C]
��h���̨&	~}k�}�M��7�J�x��0a�j9��?Pe��O#-����$[1���>˝���+�ԃ��J��i�T��E6���E�G�M~q��W��o��\2�\����0����2��#m�K�BF3��O���_X��*��RF3�nXb��(h�����o��-��ps�� b��R�Dk, &u^J�'tNI�E���w���ȼc߹���*�<��=�@�5���W�1�/�C�7��w:IA9%�6��O��7��鴧�nq�?wD!�{7`&��FF�֣|�q�����1[O���
�5������k�L6�i��P?$J�W�Z�&O����Ev�����uv���N]	t��煎����בT�D�&�c���?Xw�d���>;,֦wS��9@�/__XS�]������{�*��m<H�o9hk���uSC-�m �ǅ�N_ߜe��������Ӷ�1k�ȧT�S{i�W=��/QI[�Y�t^���A92?�b��ƙ�>�ђF9�Ϋ����?����)�̜��r4p� y��z �Lh2\l��(�v+7'#��EZ?�8gDK� �^-^�P$��C�@`��Q|���S���6i���ި���϶uh��k�\]���S�-�g����\�[�B��|{-�Y��_��͘g���g�N<�N�>���A�&���x�$tbVi����Y��P�Q��4��C���JG�}_�d����Ρ�@�}6|�T��,�Z�#zO$�S	�t�[(�U?`҃Mg�_l��,~w Ek׉���[�`�'�����	i�k#w���c9sl$��!`�xC�H"E�˵��R�������7,�C>���b
�ǯ�k
�mF�����ƌe��� ��h�|}���!4\ʖ�Ȏ�$p��~H� =1b��2z��A�����������%y�^�T
C7���N��ht����V��ĵ�r�/f�V�X��2b�E9����g��-��-F�QtR��|�9,,�Z�1;����NP�˧ �G�r�E�Xz��,�&�by[1�0/{>�vW\7|?p��;���ʹF@��!���(�>,6r��!���V�[�#���s�$|���{�4զ���b�ߙ��X���;u��}��i�vO�kG#k�]@GxCϗ�C <Eݜ�Db\^cL�-�I�j�I��qA�l��R����E�uWC�C��=z��4�&/��QZ^Y���w�� kE��/���=����UЗ��g�U$�l�L�h2ZN�{8��3�J����H+C=6����%\��!'U��ӏ�x�tWsHyn�LZ��Z)��A�%oE��Q�}�����#�яrAn���&#Cz���~(�'a����2��h@p�^c'Rh/"��aE\�!�u S�YA*yT�a��������X���S�_VR����NH�p,�!)�!	�� W9��R�R���m	7��	Up�﵆?�̻6�A��9�h&^>�^�׆�.��Y��u��=4�ikh�w�L/Q{���Z���<����F�dR�Wj;Ț����دM;M�7���!B7���pJ:ډ<��Pl;ƾ���%'��>�T���bD���<� �T�_���=�;Q�������\ u��Oz��w;)<K8M��ef�� J6%�&�^��X+.S���΀O@8�F.17������<�d�aa;-�BPy��t��u^/�l����ny�W1J����|��%�>�#Ku7��3��K�CEݓ���=]-��Ƴ�ڈ�o�+������ye��=�9 �9���G��~�dHy�l���Á�e7e�^��{NG����dF��n�
^.q�|��j����ޓ\�{'_F���:�P��HT,��+��*��5��>�m$��w���h���7Rkޅ-���;�V�Ծ�k��j�₠ ��Kc�vO����%|�..���#k������a$�xh��J��Urq��\G�P(zV�.�.	A?J>����{�!kĲECut������j�1Rv�
W(<O�/e�o��
�(�YO�9�6��y��(	��}�ikn�4R��,���r���;)_��ғB��e���L"��@u<@���:�IZZ�D9�1��ńl��0�D3�<�����y8����"?�47����{d���:�HvX;F[���:z��D�~�CIW^��U ��qӜƜ��N?H��RXW%�@�%+��;,��O6Q"��w�!� ��
o�	��s���+�	�P���M�Wf2|�����S�Ouو���@��
GN�֚ەx��0�=��b�Aٮ;��V�����"ȋ��=� )�E��� �z�O�9�����|�?�����}��=�{�5	�}?�Q�,��6����GH�+]�ᘬ8��i�&��<�H��b�Hm
.?�Q;��,���G�DB�Z�B-�������MT���mL���<#��Sjd���~����v���$s�$J��>F��[�,^W���2Ѽfς�0)�?�B*c�����>�tCq��)Z�D�7���ڃ�_X��H
pAFU��f
=��+����5�[���4�*���O�F�Љ6���B, ���I��DA���<���y���k�����*}�~xQ��H1����P�ǀ����:'��<��[Kh��G}�%�1�å�|��fu��5\�|vj6���uyC��~�LQ{躘�!���8�F8�-��,4!�6��fߚϪ��\����]Q��/��x������6�Aux��e�D��wc$O���j;����Q��&�7hj`G�e=��SQ�e����n��h
�-��x��0n�P�N(}ƈ��Ѷ��jd�����z�N/R��#�N{Hpݹ�"J)�/>��?��+�{
j�����,����y4W3`l���$J��
������R��?�)*
���1A<}M���K�C���!�M��i	Ȱs$)�=43�Z��R
�5QZY�[`�+���Y~�d�B�}ѥWǉ&� Oq��q�g�^i+�3�����j�C/��O�)ۚ%!%�݃>=H�~I*F�[��Ѣ���_G0t�ș������x�?�"��B_	h�PHo��{پS�gg��-}Q�q��� wNR~>�smJ>
�uh���M����1Y�ĎsB���:�l��bQ����F�hzz��#�r�^r��$�Pװ"������l�jS�Hn,�نL\9	V��b��hé�_�U�E�1������;�4��~��\gW��}5�MS^�,Y�X�Y�m<��Ԇ���`�z����:6V��0���f_ED��X;��qV��lo0�1t�,4�>�����y�'6:�ܽU��-�v1�9���%�q2~�$C���B��(���U��	��ʅE3��T��*e�HP�]�#���F�m���y�� U��쁓��. \�2�D�>����l!y{�����&�d\ג�׳Nª����)e�S��bD-�c(��w�@Ju�8w+&2^�8��ڈN�؋�w��<���%���b�ӷB*�X�d��]���R�5y#oE\`Ƿ	7Y��!���̠fm�o�g����=P�$��U�7�0^���7$#A������XG0g�n{R������sn��$����cr�k�$�ս���AJ.��$������s��Bf%(+��X�����k�Z���?�M�P�[|�s��f�σ��`Q��.���j$Q��j�&Yߢ4�;c;/�h�A��8�����箚v��SX�����~�[;��(���z��f����t��ܸk3\o*ٗчa/��>�Չ�f�!�»��7o��i��s+ʹ��Fh��Wo�7v��D�|�]�Z+�@j�肂۫��'�\��d�t�y�o���o
	[	>fL��s#E���#�R�So�gmw�	�t����KU!b;��k'�c�x��wy�c�<�2~K
�]���NQ�c�?����}y?��|�ٯ�g���Y����@�KK�����0S�Ŭ�a~�����:��w�	r�(���r�%J�`'�P�U8��ls�1�}*RPl %u��*�D:W�CyS�!�҄�m���/�~�2*�pb�=�!�<Q��v�����}#�,�W0}G������{*��`�8u�Aas�� �	6LfJ�v�nÐ�hU��K��㒝��r` F�8�rw��q������
K��f;y�o�;�?���%Dv�Aֵ�`j���'KE��9���`���8���6������%�45$S��J:m���J
/h.�X^��W�����@��"3��-�P��@+����K�
M�ʢ�=@}�l{~=B�k��JW�E������V��Z@�j��(o�ٶ����|�9?�� ��>����1L�M���s�oC�Jz�q�@1�>�s�J���kӛS�ygL�ǫ�*
�ji�3z � H�I∱i�:�FF����Ă�{��aG�U�w����������a�d\�K������W�`vaΟ�!�!�;���4��>����F²
J
xߺ �Gs���;��A���ݢ`s�'��"(nb�c��V�V.�wM48�Ed�w�#B���(��Y��≽啚��qGa�8��\�M�[`T�����䓊�4��_Wݳ'�����f�,�%���b_�6�,�g�C��w���s�P'7���m�v3i�eT8�Q���r8$`�ܟ�Z�*0�ȵ{_�؞,x��M�@y��P?El�����F�c�^P��[J�c?YRڄQ�4�4��o�<1%i�I<����t]�q������&��b+Y�(
Y�!)�,�H~<^��z�=�'�B�%�����_�8/��v���wJ�`��͏��I,Zt��X6l��RiIh5F��0�Ǔ�ӆ%�4n3� ~�4eA솈�W� �s����_<��#��n/�.��5Љ�]�>R�Q����K\����5ؑ>��Tk��/�(�؇���������EИ��[sU����
HM�{�
uǮE�&�?�x�I�|gRA��:�`g�刣�s[�"�@���I:���Zkf
�r��%jCҞ����=��f�%9�!��3_c\�K�;UÕ�5�u�Q^߁��x��ax�+$dk��W�'�$�T&�����`��[\�<d0&kJyd�����yE�¢D���&YK�y7�a��E����a,���r�|C��6��:oOơ*��j4/-il����h�߁'a�y���܎7[;}K��O�����F(w!�h����������l�Pc���o�T"���z����d~��l���
�.����E�X�Cz(60\���L��;J4�X��;�!g�9i�ïx��dc	�_���f=�u���*'}bW�#b3)��,�f�މ����Kp-��}� �2�O4�c4_gXB�9�5M�a黇�r7|�I��
T��؄N'sT�\�u��k�%}s���j$.�x*꘱���{=��H�+�iU4bXsϚ��S��+K 7�±��R2Nn�(�C����)$�hp�$0�ۜ��g(�Km��*������I}�i��N���8�2o�/I�' LK�f���N�ݺ
iu��W��(}�	�D�ǳ��<�8�2�`,���cS҃ ��M"�?ʏJy������������]���Cv���?-P�̇������[ց⽤�U�拴͙c3>O�������8\!a�9p�\:�n���k�ܐ����+dxy3�dr>�$93	�ʪ�۲⥪��Hv���1c�;�w�٦Ou�Aw�ʶv\��J��=&!�.w~PyM兀	n����h{��6M!c.��b�lDe9�(�=\����ϡ�¸�܀/]�s���Ꙗ�?�TlC��r[���%�{l�BV�z�9:L��#?�A�:	,�г#���W��� j�l�dX��/\��ܠ5_����iBSz����
2AIr.����3W ���0^f����/6Z��z���L�ʡ~��=�ni�,�{���,�m��|Y�C7NpQ��	<[Н��8[�B��`@	d��Ɛ� 1��G�������[�@F�}�!����L¤��63���e��� D��Ǌj1�a�ί���?9��ԯ�1��]r_��(�Βߨ���(�HM=L3��ɯ�!$�Ò��J,ؽO!ֻ�J�gX
��@y;�5�P�_�[j;mK����sO��,4����q�.�0O_:Qľ
}sC<8|�
�2<?���6��0"y�ht��|����q��[I�*$�qث�\��]� ����Gހ#*�[����-v,w��_|Cui�P�L:�~�P%Z�˙�Q0��GK�L��]�`r�U.Ҹ喅+���C��Ty���%CD��
}hxR�����ɦm�B�*ר����/x�l��v��U�Ԥ���/�F�X��S.�3!GHD�N u�H�f�C�)�Y<��x���}���7uĿ�mU=���JS���Ȧ� �A5kʯ�AQ��k�8���,�L����E�"�;�����}m��i���L�^٠�Rr7��W�����-5�EZ����9R���60#@F�2Hw9F����`�%A�\�0���ZbG�3���f����U�=�- ��q��Kz2��8̵Y^rVQ�J����ؒ��ǻ�����+��G����qb���|�^�*D�D�B���?�w$�þ4�������:u�{�8wV�$C}5�W������L��H�
Dl��->ou"��6�sk��}���n5�dlo�Qn
7���M@��.{D�
I�0\�eJI8C�®��t�Smك�#��Ū���Is���{�Q.f��tA(�t��I��%v',�Rq��u�~�&��в�/���a���T&TE:O�^�+3�������I��U���4�&oxg�������k,?##�ozi�Y���?���B� ˙���`�LG��;�,W45P�`�#�~.d��M�?�G�3����_�L{�t��ނ�� ��i�J�e�$�r��&����s'��
���(�����ְ�n=I����	���qx�r�%�/�V��y���A�\�;��2�Z���|Q.�E��h���V���چ�]�a�T�C��xb���P�o�Bf=U�V�!i�SB0އF)J��;x�Mfj���c���R|0�y�����ٔ��� �
��<�G��?�p�;o��F�S�lث �FC5��L��O������YEA�ڏя1Y�e�n0��J
?=(�Uy��}���45e5z][�2�s��~�^7���n��m�<H^S�row%]2���{�A��`��{\<y?��uV�S�p��/��?@��ze���HY`�Z�oxMYv�c~����Zuq�9Y�Xhc��Ta��h���v�N幅f��qė��=�x���3�I��۾�s7�@ؼ���[��-�&Q�_9^Taʺ�X�GWOL�h���@bZn����H9*ĩ0�N�]������qǽ�ohϤ�Kx���=�������@�q�<��`�/�ٕ%�%�����'���I��x��8>� ~�~�r����%@"�2� _��D#%��d�I��j�<_t�--h|4	i��޵�j|9X���(�����)
.�%��͂0 �8�;?��p�O���*^��#4�×��{�c�O�>���h��3��w
�`x�!bc���-[�T��R��o����շ6�G{07��D
ܦ
f8��9�!�w���9�qs#F��*�7�7|�����)�@�_�7�
$��Ai�|v��w*�a�)jL���+�?����J�%c���U�������M��}u�yb3�i5�FR;� Xr��"'�����[�=�0��?�W�w\��Ń{9R��h��s�|��$��Sϲ� Aԍ����"�멧�4K� ���\⫂���,���<��h��]�6�_�!��4n�~������C���<�X\���s����Ki��<Da�Q@6�w�*�TaD��J�3��B��z��;�t>%^�ܝMίF�T�������B�Q��L��������N��2wC�WzF���W��@�hUh}��Q��*ݭ��w�=4
�:�T�d}fa��6jU�R�U��Ewʘ��n/�{����h���Fϖ
߫ܘ�XZS*�X������=sD�|$��:����SÆ�{����o�5Ļ�kP�t)��Ba'�Y �$��!�&H'O�lwaA8 �M���H-�|-����mh�$��y��Ξ�4t��"ghY��8vue�%a���m+J�������gc�c� O��y���$�x��a2e:%�T'�_��0�|+Thp�/v��v�g-�{�~��P���e��>Y��m�$q#ƫ�r���>��F�'[;���{?�^4ָ��̿�)j���	�h�9.1�OY^[-{B��Q���@�W���z��ַo�^�`�E~ˊJ���P���T�j�����O�}��y�pg�el˜%2�"B�4�5�>���+L1*n���9�]t��V����$�b4�����RY
}޿�~����Y�1(�,ײ�GOE�2bf����8L�~��T��[�$!b3�[sl5�ĄKq�?��~���h�_r��:6T��P�=�I���ו�)��a�{Aa�u��ȅ�k�y-�$�j�;��5۩���2����������w��x��h|г^U
0�d8�?�^p�M` �An����-\6&źh�s�H�@a_8,�o�d/�<���}O�E�xpu=28�R(2�y_��o����O=�Y</�o�9�J���7C\㥎�pg��>=:������5���:!и��"��l!�x$S'���g�92Rڟ� )|�.}tf���h
m�Є�nt<���LK�&��]`m���� ���7Z��@�B|G��n6I�5�9�	����N����k��i1v�1R�v��qM�Di���0��b��}߼�%Ki�8"�����z���ȴ�%o�d*Fo�6�b��j�C��#g�q:H�-S+�T R��. fa�Z��RHx]<�#N��u�������e����5t՝��4�<��8��y6{��bl���Oλ�w��c�YmS��g��%���ߢy���[5h��({E�A��g0r�h�K�AMp(����oL��d�@���KO�Y�np!��'G��%ɼ��EN��4RO�;4��wad��2��!0<��4\$��U�c���k�\R������+��UDy�@��|��H5��{����X��ȹ�)N3�_���Y���Fn�� r�q@W��C�)�?,�� ���qD�v[(��
0���O�Muc�.���zU�$fK��UR1�E�/f�"𖸧��C��߆M�hmՃ-c�<����6�?�&�q��;���=}
֋lƪ�v��S�R�S�_!�r$.?N�X�i�3�Ѳ�VQ���>ée9�4G��P�nLkÈҩ'LZ$�|�D�ͷ�֭c(������-�QK�W'KbZ�ó]ύ$��[u�����yD�����pa4E����3��KVQ�F4�񆜓�p����"�@-�_��q8=��ⶢ;��a���jG;=139�G��G�F.����"��(�5�/,Y�+wc&Mǒ�>�g���c?9��|H�[�ϻ�Cvlg��ĹS|�#;����8�z��(2	!A���k��ѥX��:0Hx+�N��i��YQ�p���d�L�ڙ@���x�mKw�H��URNp�:�
r&^��,�C���~�tQL�b͘�����l�o9��̣m9�g?��ZY6��ژ�z[��˔jڽz�������c\ߋ���h>��'n�bm��Al�f�y$-z��RV&E����J��M��Ui$.v8���RX�="�6��E�L���4�=e ���@��Ĕ9?���r��At�%0Nwb�(<*:�+NR,:箂�:朽fj��r�A�}�Q���&��dWg��`
�N�r��k��;�!nCU�%t���9U��{�IӺѼȺs\
�9��*W7�'4E/ƝI`����U�V��Mq�pT.�!�� 9D�\
O_l��hn8�T��1j��!��mMT}7��w��cሸ���]� �pۏ��E[�_�8C�c��vS�iH$X~^���>�� �:~>�f'�[��P��z�ڱ�����0:>Z�*֮�I���w��5^�A�g�?��`�\���"�.�wH�;�3�^ ?e�N���	F�謐�$���?�g� ��>��q��^�5��dgv&��X�����(���������A)��z�Nҋ��~>r��?W���pǛ΃@dָ����c��r�'e6uf��?��ޭ�PF�&���KLAW1�M c/��8X�>����uov4Z�|�d�HM�sA4x�Hlzy\n�X`ݮ�1�R�e�ˎ��~�{���¥�,�B-O�v��O��N��,��&�XI)�
�Q1���R�|�,Gfڑv��:�u��FU�ٸ:���������4���0��>���!���;,<�,�,�Jw�4������� RDFk�2�zf�H$���h�:̼@���!b��R�Uji�\ \_���7�
7z~��=\H���B���=Q�#Q�n����tR@Eêo\F����oӣ"�h�Mu�r�N�d,��8+Z'�xhc���%�D���˜������5�q��3���% x}d7���1Y����g i���}{«jp�x���/�����	t�T/{��C[��~�;�W���� �����٘��jBF$kw��Z�[&_�F ���V����x�D�^�	��i)nd�IT Ha��{}{k' �=�s�����g[�_9=Q`�tK@-�����_�$�����6�m��v�T�E�[��]��A���l�#�z���"����@�UPcCpX�I(c��P���4F/���˵�4��5.=����1�j&�iZЗ�(l86�H��F��h���/�,~˛ �nZ���hؔivP���{�6>��~yt4�^F��S�3J��FV��y6�o�O�PشJ43(?�(� %���
���T�Ix�CP֊
ӾNt_[��D����L�W�D���z���]m�z����Ⱥ	������t4��X�tx���x~��;��x�D�.f�'��p�R�!��@�Lh�<}� X7�u��Z�����Tw�Dz��ؚ(Lڐ�e~�/N&Ws%4-�%-����@�������{�hF�Hq��xF�Z
ͭ��΃b��C�S�D�9`;�U����Cv=�O�R_(�0��0m�U��c�/��!���)\t��.��^_J����\�E�b2��ܣ��������DO��Ԓ3b���y�J�XeҟL���E�TI����H@x�9�s�A�7���1K�\�`0%�ji9�܉t�A:��-�P^�qp��)k�|�sO�;��,�O���ho�Gl�$�^d�6�!i]��_�[��aF�h�M���,�mJk����m�3��<d��Z17|��7Z�Q���	�7�t�f,`2�B�3
�|����M�ЅP4��ҿح��T�`�Xlu;�����P����g�v{ǹ
WM�|>���ɪ�aӀŦ��0��Rw�p.BD�y��J�!�5���֩�NWu���U��Ȯ�V�̟��,<I�:ߵ%�^��p{r�fHUDQN=�н���[AZ���EP�ˏ�r�
	M%
6��+?���c�t&L=�]ߚr��rc� �v�l�p��	*�#�f��uE/nu!�v|UvS��/櫻�'J����֝�0��t�.�	�2�������ݜ���m��E�*�Q�?{*T��T�Z3��x�{4>�&Xz�v*�n�⚟����&��:�<�48$$Q��g¹���_�/Y��<�J~A�9}�̭Wb�|@��s$�CT	Y�^9�O����q�Eyv��;fw0:��p�n��P�Ț��D��z�6�W�kS����^4),�,�y3T#$�c%�g��L�.3�����X�?rI�������@y/��cz���mj���x�u꼯؁�ϥ����ƞAmJ��WE��,MW(���Ő�)��������yC�a|�q�V����݅�>�qGZT:�q�_�^Q`!�^��"
�`Ε(�(I�<���
��I=C�Q{�Q���{O�[�����78�4vh=���2�����""�1�:hnK���澇R+��7��Jn[�q.�V�N2$RR�4�X���g7���i�����+	�(,%�z8���`^0 �Ubg
T�ʟf=!�X��*

�/��q_X+!�����>HX�S�c�>�+c |(����:�A@:�驃K�9��.����I�:�O���QzD����rJޅ������v��@���x�L��UjF\^tp-8�V�����s��@S�koò��Me�H����B��[O�����l�A���� !��ZH��n�J���/갶E��`��т�H	��4�:�Lf�O��G��OlȆV5�A��GйŐ�c���j����x=�̝+H�`Yυuu�h����V*�떕G��QU#�������|%��:�z{��"TwG�d�O'�&9ԭ���{7u����7�)�f.]��X�P��_�*/��Y����!��5bN��EJ��E]�N#X�§t����GR�o�'�}�o`�Cւ��Ր�N%�rZȶL�҉��I?Fjn�w������ (���{]�,��(
.VCR�Lf	5��sVj�S�8�Erl~��N������֡�d o���vƂF���³P�4~sv��=f����w`R�g2k��j�s��P+��1�V��>ݸ!G1DC�AI����E��$U�@�fmk�=��&��kSWe��e�8��ED&�NJ�)�i4�|��$7�R�C�<�fy��.��Q��fazFD�}����	ȘȲ)CX�z6:�f�P���.��Ŋ�ٱ�)s�r߳�(�|uJ*l�S�.1���e��pi�IWY0g������!	����̱e3F���ְ��y�埍�'��q��̳/��6ë>�l a��~�M�]`F7�ڤ�ƾMS���e�����!=n�ģn��M���X0k�A�����_�KV"���gRKs�*L�(J	��<o�R��}`'���*D+�l��R���B����N�%��0�6�ע�p�V#�F�[I{��՗�cr��A����F�;�s�X�'+.h'M�3^>Y�p"�����o���\v��kC�i#)׻�������X�v�&9��2k+��Sa M�� B�(���������1�rRH�@.�]P��;~��S]�y{�$�J0����j�`�71�iJ�mz�(�0��B_T?�3�LZ-$��A-����֛ ��₂Y������}s���5vp�N�g�P(O��ϊR�]ck�(	k{�tm ���u�RK�
E�B��,���W��[�Q?v���H��H����Ɛ;Vk �<��!�V$31.�dJu���:�s2w"�qIfz����{�{��S�����du`���_kES�W �l�D�Ѿ�I��Urɯ�S�K�H��7���ɢ��;�}%Cg��$$,����	V:N�瓠�]�a�v�V@O��TJ=pl�D��A�;�ID��5�I��S����9�.H���kO��g���[R�T#T�
�ܑe��yb`���ە+�&�	�P�I�[[�%���IJNSlS���d���qL��/�k/���\�f�ŉ&����}��S\�7�_��=�1 �"��CR̓�ėy�l�a.k=�	�TМ�M���b&��E���~�<��fcU��5��+�X�a&�\�s�I����zI�����b?��Nϥ81Ҍ曀�ٚC��FZ�Fv��:����ܩ�)�_?�MF9~�'h�{resP���2)82Ik��d��[�����ڥk��m�̂�q�&΁��sw�{� �S�ʏ_�Ma���s���ϷG[rx��;r�hʑ��n�7]Zg;?>{`.�̞oY����Շ
�l�[r<��M���%�cԯ�U<h���W8�5�yfr��̝=���tn��m�ɖ�b�,�Xa�7�3���b��)j
buff��z�M��,h���#���)#R1�Y�o�x��(ə"y��s��y�\X�Rx�%H�~}ܳ(���Ֆ5R'R�Iq�c|�����+S
nI�ˋ�*�F��j8ޫ�U�%O	�^"���esF�抏��ny�9����L��e���h�|k�,��H54��p/rQ�!�~�8�T �zY8^��@�$�z��\�fF� 4�� !��h����W�c.��k�ubmn����KҾ�" �Sx>%oC�E$��&V��������Y=?(C�.w�a7�����c-r��>6�j��ì���Ք�
��M>��\�C�t�ǿ8����OlĮ6��Y�C��5˞�x;t�W�1�,E��ۘ����m�;�%:o���{y����vx:<%�^:�+���Io@����J����zW��&ۊ=��*�я�=�����-���.W'�+iǞx��0��5,�#�	w���gS���(�_�n�Ďg>Ht<���w*�?u�!E��ez�Fh�P]T�^ϊ�����ԮC�q�q�g{�Q�x6A�?۷1��g:��,دV��1Y�"�����.]i�_<��R�xU���3�S��5�Tן��h,���o�k	`9٢e�ڝ��?�m�tS�_Nu�=b�ĐV!���MD����և��a7�&�r�Ղ���Q�&J����<��x_ώ.\v`��o/�7��%56���{�7�i�Z����X�<_�'�;K�?��eCj<����Cʝ!bd�
���� s/��%�t�������x��eO:�VX@��r����3��%A�C����S���TE��#�)�\]6���H�^C,��~N�R!Z��U=��F�r�Y�|������<�f,ꛎ�(�g�nE�s~���:+^(�aM�4Ƨ��\�0֞gфDf�����f$y�X�e�EF$"�uC*���8o�}�	o����m�w.�������ڱ��ZM5!���B
C���6nӨ������@<�� ۨ���8�2;�1����}��=]N���Eڎ`�-͵�L\�`�,���Lb�%��:��e
_��jO�3 e�8�EH[7ZO�D��hl���������q��.��(z�|b�����V�RO���>�-6- ���nC�V�~��x=3Uax7�$ߎT,/#@��˙�@�K�{�����)�`�J,=IW�fW�ڬ�Y��v�.{D�;3��I���}���������ѭ儡���"]n�z�+�&��'�k�M#c�lF(�ޓ9�f���� ��������D�&�ky*�>���ǌ��⼯1�<��7������"m�,Ų�G/���B������̤�'�U��J�a�`��q�3�<��@C⢣/�QvL:�]����y�:]R�`	| �*�bW,���u�z�O�c�lݢ|C�lX��� H��_��>K�<�a�%�-�%���A���'mYS�}86��Ng�̐���;j�!>=�
͛������#�-��@먵�����O���Ɩ��I�d�c^b���@�Fv�b�G�5d�Z)Fj�OT���ʺ����������c�J؍�ì���̞�ۻ��.9�s������1=�� �����f�F�5W�p�IЂ���w<w���t�}3���
�B���t ��b�Znv��}`�ęmIv3����\�Y<����AX'2�|H5L{?'Q&����?��Հ7n����o�[�á��Dv��]_�b��J����3j�T�	����H�����q�S�X�*/چ���
�)%�@I���I�X4떉H��YN��A�]M~���͌H5-P<�z�dT�ܝ��I,�h'x�8u��	�Tm��M/U�p[��\+ g����+�J���Œ\T/����r��� 6���h��m��?(+"  ��g�tĭ���@<���#j/��7T
ydQ��}3��r"̣���.�?�5׎�2�-&�M:�7�2�DG�TZ\� @�MhmZ��N�\%Ng �R����wa�*��?X?G&DR��!�l���8�E�0��@{���N Ry̎�����L'��.���,I���ٶ���(^�B�*mwiS�p���~Y�.{8��WE�^� D�H�QJDH���5.#�E�}�d|%f=�D���EWt� �8d7~X�٧|=S��!\��a�t���Ir��p�G[P;>ҭړ�V0��"�{��B�?���]k��>���QU�����	'h#b�}_�(���dރ.��60��'��56+͛tn�$2��H;@�p!6'a��xa41���<vhu���p��� n��׍;p��p��Ev?�5�N�v�}aM�?�)_��ġd�fJ7������~�5?{gtzپ&c�e���(aitQ@�q�H)ͦ�v�W�+�6�7@]�G	�K��Z�xr�ؙ �i�ܷ8�~�ACt�xb)��VS�,��K�����?~T��a_ZL�`�j"���fLf�*r=����x��~A�{m�K,t*ǠS�ec� l����WRB�8g�jv�����+�1�[pf��R�����n�L5�2~�%���0�і�`oX(ņ=v'�>ۍ����#t/�R�	��Y��|���,yYǱ�8A����8��q��(���������Y�0^����)l�Vo+TY:p�q6��k|ƪڂ2Ύ"�UBJm�� ։�pN̳�����}���nϒWp{7p��Y,-`�(X"����g#lj��a񕢷�?�.GZu�½�V�޿W
�^%,=��<ٻ�t�4���>���m"vZ�ρB.ӽ�N���.���O���$�)�AG�YV�HB),��8�S�6{D�K'���V�b=���B۪�w�����J��<v
��}�Oy�2����L�G��h<���ߐ`�e cz%�6:�΀����[@��mɀ��0��>��x��I8��ڣYl���ʿȟcx�
���L���4�F�d��g��B�T=l�ZR�����D��*���`w�ì��Ua�3��%�G������ ��:��o�7�_������D��Ù��>�vM�SO~{|���
��9��R���&aռF��e4�W� +-c�Nƃ1^I\GQ0��[m·��G�p���Y��R�K6(1c������_U:EG�?/[����!{��Ǽ��r(-m�"�7���z�� ����MP�@��NR�?<-�����K�d���e�H)��&�KZF���T�Y/m�K#:/5K���Bk�d��J82�H�?�EC,�*i����>Ⴄg;�T��D�	��E��L#|H�F�tT�	��΅���݅$s�&�'��ֵ��i�t�N�ܟ�Z�{�{��]q��5`�/p�[��Ĭ�n��J�hk\E�z���?��	�Po?���~���O��H� ��Z7YSks�pC_@`a�-�֊Hnv������]jr��S��s����ԛn�,��$��e&���s�▤�|�Y<q�L�	�r����wwY<�"�3F���רSꬎ�!/o�
GU��;� �RI+u�b�(A�ևj��l����Ւ�!2I?��4Kd������1�]�E\�s_�.p>tI�=�T��
O��bHø��'`c�'�>Ϋ�����4�`Y��E�,�6j��d1���"���'������X��8L��O!�5P�����d������sT��=�ݫ>�p�^B�Ǩ+��Bft�� �`��rCh�l��+0ߴ֥q'o�.�u,��*(�핿��?��H�>ڍG�=Hǳ��;��D��!�)+�����jي�p:	����ár�\������m�$�i'���żA&GQץǆ�Z�X��ԔA��&J፾O:+�Y��&ݛ�����ɳq��a����1��Q�٬������΢\��8��a�����)��V��8)���p�G�T��uo�l�i�Bϲ��S��J�2��(WU�L^B̦{I6�P8��?e�� >=�������g��єD����(��88��a������^<Č�l�'�@#2��.�)!�W^�E?h��u�^BI�����X�qf�,�8�Ȗ���=q�%���%Mx��~���YRS%�_���f���]�%y7`iE!:
�ԇ�ʚ�W��k���ٙ4@��̹���^������h~��@��^��-{o���&�)Y��X�u	흕��̹�T4}��yu�?������9��8�<o�� �'�a]G��Sһb�$�!���%f��i_K���l�S�D�� )aR����0B���Γ��d��*��3i�7/�H���
T�[��t^0L����P�٭e|qMDҁ
��Z��)�7-�Z��.@͈���Sx�/2����*�H|��&9�a�MF5��_��B�6 ����m�Ҥ�s�e��,Ud�6à��\P�Nϖ�4$�1�g�J/� ��+�,��B����p�wM&$�p�YW�C4�(y��c{bhS�.�d	gL&������e��6��SNe�zV	ˊ;���Nǔ����������-pG�{������@��Y(�;�$6wͱ���Z-]2�r()5hq���f�^��9��,����4] >|jHBh|n����q�� ���S}?����GV\��%�{� ��-@�$!rj jZ��
��K�r�^�ϿT{߳ݑE)� ��fi�ڊ�,�?h��߾xY�&�w�_���̊�j(�rE��Y۔���H�5���f3��m�!-=_����5%����0v��g�Z�a/*�E���|��*���q��Ȧ<����!���M,�!t�v�uHp;�-n�=��IQ������70�MF�>�i���?ҰFfg���j�`'��5L-��[i�7b�?�����U-B��xY�0"�����������
4�����������rP�,�� D[����
���)xZ�%�TֵS�3�·%��i?��'K�V"�B�k5gi��#�� ��0W��`2��uY�k�]����U\��|�<�`Mݻ� С�ݬ��{<ȅI�o����_�w�FO�:g�7ě1��Næ#�*� 8nJKdg�X�6���M�埪I֮մ�1t�x�kɀ؀�{C�X��	+'p��QM��6�o����9]��$��~�o��A�`\ko�@~;FU�G�����GqGw�rYIa���j$�-�t�Yz�Y"+ݟ:�;��WP��C'��(�ڲ��P�p˖��1����(Q�&0������d���3�ǈ;��?KA�d�r�(AY�6(����f���#J1�F~��=Zz����B�g��'��"m1t����1����@�4�]�VX�3}?1j]/ؖ"�R,س���GU�N�h4�������B㶳�J��t4��Dȡ���4��E�e����n7�-|�?���H���kcK]����`�)p��ZR��[oi��0��S$�QV���@xaNb�e�e�;N/Iig��2g�� �w�:���3���{%�#t�?X�w��
�t��*�3��|���D�#�Jiqh! u��r/�0݃jy�~��}<�t�t��H�Ea����Ԕ�|r��T��0)�s�sɻZY��i/����+��a�]#��5z�����[���º���Վ*���w��߿�_���z "�K�BG�-Q�z�w~�~�ǭD��~i$�(�	���jP����5m�M��K2�^�ޓ��h�?�6�Uu{�L��N�����Rw
`Fe9�E�F�<[� �2�ۺ��/Zf6K�m=nk�_c��c�	N7G��I��1�[��*�B�{�ƣZJ�+6�� +s:=7Ӣ� ��13�#S	eb�nb���^_@H�=�v��j�[@jy�oC�N��o�%؜���'����dXV[U�v`����@Ə��C����R�h9��@���{�j[T�w��Z]r����q�ؼ
�2J������Z�Gݢ����ǹ��eb0�(��&��G+�?`pc�Hy,�@׫ ����Gtl��)��{FL�H����}�O����=�h��<���[��&�ă3�1�)&��ҹ~ t�8?57¦���\��� 3�e�Lp�a��72�?u�l籈�4s���KMOЫ�J���ڗ
��w�_���d.3�Q�m�[��y�Q��FV(ṰX����ꜭ�pý<]�!�����{R��.7%�[@o��� qPH�>�[����{#�s�ʓ��c�'`�ab*c:��y�Pg]2 =M����ہ�~��HԔ
}\��&�t�57g�/�/��X�rWv�8Ѐ���A-�Pӡp%꥝�&WHh	��sO���������#��Om���$�o2�i���@�� ��ɄY
B���C��ʀ��(D���g?pb{�غN�R���e�G8)���X_� D�%xq0��3?l�O~��k�=F]�æ�Y�%�6��7&}wGJ���8���i��<���t�'���GH��Ԟ.q9�4��5T#�Z	��V˰u��Y�\v�, d|c)`�N��CJ��띅6�R��a���t�8�o����q��բ���j|n:����M�9�:Ud'ǐ�h��P�d����H�>h�^UwFcf.*����<7)*R8B��x��N�8g;���/�ޱ��� #1��� ����ϴ
7�*>s�{�Q�+9�ky��ؑk�ODZ����8Ka�)Y���F�G�_
��>�8eJ*6ډ�J�r,AyN'3Iü����ןU�Y�=�m:Rc)��Pd� ��bԁĤJ�t���xRuS����{��0�vWj�SD��Xd����2�	�ж�&��r\�Y�j^K�NCT�^�8�T[4$�����~d��%�n,�D��3���L��F�H�Qnxa/���C�;���Bj����ge����++"~"oȥ(�^�)���#vru�`�_�:og߻����9�-��Ϛ1�xv��_��4�dd�V3��=g_d9[��88}�Ba��[�mJf̠���s륳���s71��n�e�˿���-..��Gq��W�J1�m������U�-�􈭥�*�l���aU9�����vJ*�&�_ϝ\��;� w 辑��*c h�ά�%v�$;��;��e&�;j[����Ô�A����޸�D31�ӱjp�Nb᧺��͆�O,��,���?r��զ�@�~oR��n0] �[��3�+t��>����1�p�׭��Cu,��Z+�Ng
�\��$_�h�Z�if[(e�)�x��b\j���ҀaE�n�<��}<x[��)z��`qCҬb�T9�ޑ�Ⱖ&���1�2�,���]�c������<.j�ahT��O#T�py;&R�ʡp|���03�W�X���� �2���w�ؘ��R �L�h{)VS܎��R�ɐϚR�����y��}�'Ö����/p`��h�ץ6ÜǏ�����)*���d?A�A$wd~ɠc���[U|6��M��+f4Mm!����rH�w�o��ѵ��(�xw���}����^�L�4^*+ssA���j$� ��Z�޴�S�4�3k�}�g��mm�n�A!�Q�vX�z����C9�X��Ძa�=�d�b�f����>�HP]1T
_w�^dYgi&�Y[��R���F��C
D��r ��	n�/<"�X��HOxCğs�9Q%z�$x�֖%!�q���d]oGs$b���\��FW���V
��R��f�P�1fA'��Yw��"FgV���ۈKo=�S�ipa΢Zr�<�(�)
(P0Tzx%�����P�=*p���ʢ��*�Rwi�g�o��D�Rxݯ7W�#�}��Oh�^~��G>B]#�P���!��6����|=�S�v_�u��)�w�ho�-�Y�BzWf�<)GrM%���\dP H{����/�*��(.~�್m��-�������-yΆ�Jis�IP���dא�g	ZR�:��i{�R7�-N�L{�%S򏠅�y�8��0����Ld�B/� CBj���-һr�����<}��s�mӾ5z��v���\)`�陆����G/�@+z�)�#;��W�ܶ"۸;��R����y�-g���7S>�@H(�qkxVPX�.4b�k�����=� �P�9s�2��r����$�꞉亵5����-I��w�y?�D���A�]�$S�F�j�c�-	�V'?}�	áۄ_<,(�E ��OsX����f��|�x�����ã�C}��^�+Z����|���\�4u���i%�)��Cr�D�5_�����l�4�QX�j(U���͹�'3bY��Ĝ��_��^I~��*�<�O�F[�4�ކX?���K�
�C����a��M9m==��͕�Q��	�5�Ԍ���<�f�H�R�^hk��0�eF���s%{Arv��5��x�5�d�Y�Ͷ��A���U9cǖ�E��I�q�Y]���m��G�F�z0i�����(�x��9�pM��M�|�_�G�3	`fz
sڽ�z¥�e���֯�%yk�j~�T�;����s��3��2[����'��>�p$.ן�܍�� �g\�3 ���o`'0*�I�؃�3Q'�b1	4�널C �fJ������mn��r�X�d �����sr�:�a�RU�wC��+�K�
w�������F ��F{�k��8|9A��&�J������v@6h+A!T���]��L�C��?gt�TZ(�r����J��)A���)�_]�F�O.<l,||M�o��Xb0sz����O|'�ˢ��F
�8����M�k�)d91˄G
+��8[�	LxV���_��w ��+K��p*U+��y{t�d��lԨ<�q^:]��.���μ�1��+�vCuIQ\���>@�[�0���7·���y-�>����<�#��=ԔBǯb� ����-Ĩ,�Ȑ���"��b����2*��Wǯ�@�r`	�8XȬ?�B9�o�b��W;�D�Қ��`�`(�4>�.����]��u�v̺hCA�6�H��`P|g����٫ٻ�h�T�q#�y7N�锱�HΠ�?�X�zizT����������h�����L6�{�q�/S܋��_�����.@.��������b�|���&�^Ao6Am�Y^_3Q�P����6���_{���)|L�.�S���ῗ�8^�8��Gc�^i/E�<_4Nt�8������j1[	
�3�О~�yOyStx�"\(J=J�T� qe� Z?�3;2pm����~�I�I4�Fة���[�]�"�w�-k�3����!6�I�)nc��$��!Lb�U~	f�;i$in���q��c~Ұ@���� /?�T�!�*�m���@�M���$Qƚ��A��6�rhX%��.�/S�%�4����r�*��ƽZ1�)]�i�i���\��Rع�D-���~.1>
��D�E�{�7���`Ě� z+�m�{�I����ը��!��w�J<_�jٶx
��%��O!BN��}y�
`��St�!���e�YȪ�Tjv��lt�|�37]Y{�4�!�a��������Ĕ%���_��ނ˿שl�b�U9Ԥ(�]6���h[3���o��C@]��j�n�d;P6�-gj��ڄnJP���zoK�F�)ݢ�! &P"P��8o8�ڳqP��[m������ů$u+ygL��Q�)U�䞆gM�r�ij�"�����͂޷1g���Q�ԄR%�r$?G���0�͑����W�C�A��p�WS�H�J��Ű��]�C��D�s8d��鹶w��~֎����OG(���Jb-/�aЉ
�g�k�(�<�]Q�D= `ĩ �|:ʵ�tb2��&
�HP}�1()상k��n�j;�������� ��{�Id[Yp5)��9��l	�^%��E�|a�� ���m��-�{�D��d��"���2G?����.Kp�_~t�gOM��H���>�S����
�Y��]�1?>���>�)~(s��3�{����T=�܈����3�Q��ڥ��W�<�_�������* �X؆�!�����`'���U��4�s�����5��ֶ�U���r�阢����������;Dm���؊~��.$�~�J�$I�5P�7~�,��9w��T{ҟ�o	7q,��ؾ:\���>��̲CVz�_-v�>L�#׏�;�<>,9\hb�^�����s�%N��'�6n���.G,P����tssZh�*[�S.'��HѴ^Gf�%^H�ݢ,�7V�Y*���ǌ�s[�`l�F�"R�3�Pc@5������#�b�Ӱb/�%:}T�]�����`A��f�HL0��)M�s:3Q�5�s�����H�	ѕsd)�U|ف��m�6:6!��wP�6_Ҿ���ʓ���A�<�����6F�m�&
������/W�Jy�#@C��ة�8��v�<������RR��-��I�W?���w"s�!�_�����c��f��OM��ƹ���g/�f;��Z�$��VB&�\*��("%9�my�*VnG>v"��[�ܘT���lg��t�</b�:���T19}��N���=�%��+O%i{�{�P9� :t�ÂP�E�����}XR/G�� bⰊc��HQWH�G��X�r�����a�2���k��N���O��{����t�J����X�p|e��U��OGY @�C�ct޼̵�B"�:��qI�e�|�QC�M缺��bJ�n�=�c�*W3�t���2���b���x��8����7�Ld)�{~�'�kE�4���м�ʭ�t���{���$��A�bh�Y�Uv��g����^tf��+� ��o��J�\{UO_�H���"�s&�s�P�D!\g��A��\��>�zj��&��.�
��U�^�;i8�2`z0���>�z����o?�V2%�4�
z�3����G�(�Q]9&{<��T�4� ��)OzXm��G�_�&�V8z!�q�,���y$����T��Zz�h���t��@�lL)">m�9�Q��.n�,�n��4�*��a^<�`�o�(�ŨgPU�vz=y��S$��O��R�R��}w:I3\9",չ�h�D��]�Ɠ���:����4ɡ@aI��,�	^�qC�!x !K��� >_���9S#�$sv�T4I���N�xĲ�@e�*�?Z�j�Q�BB޿��~xY,b%.�1$\���'GF��h�����<+\��Pl-�1�tҘ3�cG�h�_��@$���?���&C�(�Q��#O���+h�O�,���z�/^�T���MQ���PZ𸾃��&���pN�W��Օ�gJk�i�����͛�FC[���:7r
`Z�HF��:$+FD:\<*[K�C����㑴oZ�[��k��c~��B&3g�"�����ov�$/�{����3I�pyֵ땛�ZTqbc���]�~3'�OX��Ʋ�X2E�<3�9Že�&�+[*����&z�.#jw��H
�e��9&{O�Z��������3�hդ���D��g�o�-�J	��f��+�_� I�}��Վ�iR��G�×������A����������aߘI�{;�l�ʷO�3��-!�.ߚ?�1��)X휁9EhK��˒����N���idK礄 w�G聼=�e�d��O5v���~��@�2�:!w���Ww/r^ۅ2w	c����Mb���։=-z��)�ʶ�M����y�>���n��\�#x�M�W���U�_���r�:�O�oM�:'3�A�v��E��(a��R���+v��D�;�Z��4"�𜞾\��*��6��f����>q�h�]�S՛WI�oi@^� 3�Е[�	��;����9��|����g����U3yF@՝ }�N�RI�}�N��f��7�����.>�RL�m4+�o�7ᓹ}4+E�.��q�Z��$(4��m'�4%��[�1�_)߹R���P�^�6VgN����'W@�?]'�▎���t���X�Id���n���<�GH�h���ЊJۙ'UU���W����F�I�bƄc������[a\�;m��(�n_����Af�Cֹ�?Gi�b����w�V���{�N�E?T�~���/Ui~�X��Xr*~�l�}V����e���[�|�N�]n=0�[r�V�t��k F��_>q�M��(\���$F�.e�<5 �O����7դ90�j��S������Al��?�����v�y��7�9��^�G������%�h{�xqm�^�3+�� ����S���:�/���xF�*���d����'�G��^}�0���}`0�b��������eX�������8Io������td�ɖ��9�W,ç����G������H���B�8Cv���%��\;x#h��[	��{gkBGo>��:݃��!� uN���!!A��^��y'~)p|���=��']���l��
��c	�[e��:+4GWuT��*��{ׁe��sI�s;���Ok��@��Ò���~8�r��{���{偡�b ^�`�]����sX���ͧ���-������'=�>Y� 0�˴�Ƅۻ�@q���aΐ���@z��4^s����!]�֍�̀���V�nUdz����0s�U|��t�� -��/[o��{0�����	���i)6Π�@X�:�nh�$��9(��|�����J����O��c�l
�C{��~ҥ�=]U�����5]�������y���9���cΝ{�3K�l8�$�M�Wʩ����,����_��}�Zo���b�I��f#��S��B|./��7K����Po@mog��N��V��I���k�X�j��Nk��C�8�d*�Zr���B���W�;�r,�{��x���];���%@�-!V���O��ld��rt`���4�n�hw7zL�Q��uE uJ�rA���y.Ut4�A+����ٗ-�8�G����1�/�Q�8�2��ֱ[b5H�Ws�L�H��kJ����npz�,�fN�fN�k�.IE|��X���`Fn��͸���b��D�'�U���Kd�V����gW����+���w"06��I~���Yf�	��.KL�y�p�Z��[>9w+�cz8���O���B�_8+���@5L����%pPi��˿Be�X�(#��i�7 �
:E��3j��T�iG�@�u����l�8�����U�J��1�&M��ܛ���+�$fކ+<�B����+ʢ"�dS�V�b�3J�.����> �RQĊ���̍�.n�qJ]y��~9���kb�sg�)��=���%���bɾ����X�i��F0�bCbf\�*���^|��Bu���̦>���4Îw�-F��̥v��3��T�����_nE�����A��ԁl�n��ՠ1_m��,�K'�z�����������Ԏ�G�*���\��"TNS�g�G��DN�`�uJ���;+(����,O�N������7 b���ʸ3p�5.e�|c.����f�K��������(oP�9�vF�ݩc.�߃ν����S�/���It^��|Nµɧ�@B�M�� %�zP�zZ�!��p�>dekv�R!�r���, @��՝�NU�&X���֕?�i���-W�+b�HR�oc*aH;w)5��ZrqZS�.��>�?�3�6��o��Wx�O7���,�K�v$�+Kl�nŕ��x)�$�/��0�<��hB{j��u�ַ#�>""@�C���[D2�&��bv��P�6X��a��UÂ���>�5Ÿ1A�x��
]0���4�]̻;_����
x�s����\��{�)a�Yk
p3$�u�9Qo{�����-'Bt�
\�#����/�M�%��^l�Lp�����I�{/����R��؍��JTB�)�a�k��E�{�%�.��}3�7���^�zw��M����5�Ҭ������I��5-t0���l~�O�_�Y�?Ps4�`��d��WT���iE~����`��T@��2m��?��pHI�|Nǭ=�b��b^���w�}Z̊?^
��z���Y5�$ۋGJ֕(��Z<�����ܔ6)��ݶ����:�6b���L�|;�_�AwG�P���&I O|&2Ƌ�� �2B���Q�N�,5�i� [e����1��:�S9��o������ӷե@:9�ߑ="̿
V��J)�f��eknGҽp= P?� �gg�ם��̩(���J��oX�0 tp�|��ճ�v!@RN,Ӭ�@�=Wcp&����A��>Q���gzW��ro=c�n}��hA��+�����F�d�X�g�J�fh��O
ല ��Λ͢4q�G�|ۖ���Pi�&X�>/�ifn8��@`2�c�*j#����b��./c�mV���~ó�l��ʍ��3@��㸸t�1��K�҈Gf��u������i+]5�5�^�^��[�F�`����X�\z�O_��ǝ�>C�>��D	�Λ]��:�!���O5�mA��b���BN[@Km��A��-x�w����K\���	_G#Lm�{v&���>��2�_�OG��M;�m����$^((1E�t4lRW�id���[�
H=$9�m|�6D�����G ���C��>5�����I3X��ˏ�b���N�F��O,)����i�<[��h���ݫ LJ��X�Ʀ���P�n�g�w%'�֫����9z�B���A,�F�f�lA)zR;�M�m�hFAU�s��27����PB��8�tr�6�����M���C��(;&/ ~{ZH����;�E�m4J�W<�@�W�����zã�X���������k����e0Yf�]�x4v�]e�$���O��۸"3hِ�fW�AP4K�Dfj�G�n����y��sX���r�)94z�^�!�4�r������ʜ�������؃N�;,ߺ`=1�;�b5�_J9J)�٩N��#��F��ki%g��p��`��U��A2�(��IC����wT���zӟYŐ�G���;J�ȆƱV�A�>�"���ъ|��'1�9rC^�̌�%b���1USX��')�+��.�a F��R�@m5Z���Y�(/�������iH��
/�/��Ɣ-9��o��*VJ�J�O|�wQ	�~B�f�%�5��tm�� #���_o��r
���aQ����<�q>K�r��jMe�i�����T���׸��S-u[�=���ER�kCUqTo3О�N����D�����	|q��� bh�&1$h��Sio|�'�x|@>�,gx�,fD�j��+���B�/0П#�a����{���۸Z�o[�.�_���0Y�s��@��7Y�+���zCoj8FX`x��x������l�S����PɷꈹrX!*)�$߼��>���.�l��Qx���ې��(��xa��M���I���5��է����?"����;�l��u5R���N��/��@���)1�}-?�����F��C#�9�8n�>�w�6=��x��%�c��۞z">�����5>�&�������7����F��c����,�,����{.�(V9+�6�+��	?z	�y#7�G��d�~�(s��@l���>���Y��5%�����ɰݢ9w��1]^����r{W.��Ǻ��<⅘k���	\v���� �Tx��C셧�����·���i��Q�~4��*ѣ!����ȯC�>k�!A������f��I�Nz�x*A$���a:��ӈ�ʧ!�WHx9f�_�bu���P�f�/:'F8!�j!���D�A�s.�^���ܩ�*�Lܳ�b4������A�U��� ���2�}$�kM?��7�k�g�qa�9X��U��a'y��Z$�����-�W�o��^�
��+n<���3���9E���s��.%�50�O���I(A�K�#�*a�}��J�>�?;��\�K8KO���󤇝��I'�u[�� ���(��C����%j��:�Ϯ���,�rϚ���A�7�L��$�u�I
�����0����팑jML<	�6BL4Gz۰)I�E��+��am���.uS\�,����l���	�/B*���Q\:1���f��A}2C�� �Xt)�\c�C6G�e�R�v���Z|�N�Dtx�����n�a�z�{�(�͒���������@�5�A���R*(W0��p��p��p�Oo�\����~RO�д�CԿ����5�Kk���3D7��<�^ʪi��c�ة-O�������$����}�#\�1��k_6���T~�J�����1�jRⰷ�bn�!��X��$�vI��R��8%�ݸ�:��M7��d#�sLF�l�ֈ��բ{����d�/k �X� �v2Oݜ�n�r-��x<Z
w�4"kXܬ��G>�Nuy���i�h{yH'U�ȅ�=�'��9�IY0H�J�M�9;�s���jP�'��*`y�1�|;�\K�^�3r��aC�,�� �~�Ca�ii󐁧x/D�r���QS��̥c�))F�0�
|��928)�$��h\��R�����/<�,��L��Z�^��O�9�,�l%��~}�Nm�O��'�s��ebuo����Y�D�4�y����榵�
0�w/��b¿yʎ�]:N?���I�-�K�]M�����6��D'k�Hl�u�YE�:����}�R�l�e�h�V-Ez����e�y@W�p�|�}\���iV�oC�����kEW��+J��Z�jQ��QA��<@
����\�9n�Ǵ����hL��B�O��f�Y�<~��G�Ao�{��Ν^�?�#9o�=#�A�Bg�T�!�,9����XT�)�K2iy�M�#[H>N\��������cH�fZ���
g��fC��	vC�l�\Y��P"&���>J[A/)�Rن���f�=H6Eb���G����Wr�,�g��5qx�,v�'3R���T$���\+�.��S�4R��ń��B���>;Db%wI��"I���?+�Me§h�ݒ���~���+�tz>-�>.��Ij�� ���Ɓ=�]���4�u�P~���=Pz ~ꁶ���p3s��3z[3�U����V�r,�%�L�Q�ވż�O�P9���݌��cA����	O��M�s�_u_4�I�Y��>M.�Q�<�k�yE���L�ŏ�������1��u�p�H�-R�}7��a"�і�]�d���$��VU��E����PǴ&MV�[��\��sA:����7�k*����/��S�����'�"u�fȀ�2���v�=��ȴ�bA~�Q�R?�MKl����r+��&�O�s �M��x�]��Q੐RX����Y'D��zaeB�f	�#%'%7�
[��O��IU�zy�����p�p1sH\��n���ە�B�#��Gc�Vc��;���a�h��ϖ��1 W��
�{m��l��k��N�R�>�F �57� 3���{7�@:+�ӣ�tԲm��ݟ[e�j�2 �Y���f֡ũVЁ�΃=��.e�P��I���)S|����Ԥ�T�0��A�Nq�b�:�}�ձ�!����H��5##ֵ�d��M<�w5n���GwA�	��D˩
BU�MQ�,�S$^�60�E~I�ow��>qQK�7%~�+[=vO|����Rp�޳7�em>�# �}�R�s�+��-������ۙ��������������XL���3�Aac����ik��a��&S�2�!;�Ķ8���e6��.9���^�洞|3v��R�.??���f���L���wGR�[���:�10�/g�=X�Ty�����Ť���B�+�h�0��5_7\F��"��@�Fܫ=�cl���Ѭ��y E�	c��No��gK�w�̘�z���w�P΀�V
D%6.�*.t.������q?�ۡ|D�������s���u������������x�3��P3����ԕ�	��b�+l�D:dN��:m�v���ϟ��Q�HSjZ P��H뺶 �(]��A��@�5^�# �~����F/9�܏�h{y߄S�M��4�=ի*�˃���6'ӓ��]�!o���j;Ak9�셁'n��2�k��:�/��
���׮�ޤ0�jY$��s4�Vq�D���,���-�qp9����-Mڵ�w���A�0�!�29����G.���u���z9��Wv����Y��y����PLo6��SE׶�˿�#2�CL�d�=)�X����?A�^D]�D`r�^�U�Gf��"��7�SH�~�M��ʏ6Lܟ\o�4�VA�h�����Lq���݋mh���s���(^���$y��L�,������*C_b�o9"R����7�
�A��˝��|)^������C��2����(��bȰ�e���5a�]u�o�Ţ�Rn��R�_Mk1dǕ�۹�Y���Lćo�n�A�e�\��`}	�j��ż���%�J�$0C�N�*>I��OH��H�v��f�=
x�_���+��Ja$��p�S3:�J#o�8zK�.��y8%����4n7�S�hLHQ�{� !Nr��֦�86��0�ql�<�e7�q�	�L�9ҠPڽ�t���Q���%�!.�Zʶ��������+��?�!&3U�S]����չ?@��-6�C�:=b`���׾\�'�/g4c[��<љ���Ce�j�Z�8����߲�u���_;�~HY������;��^k_m���PxP���J�����D�T���@P�T�.�g;�mi���.Wu1�C�M�؎��0�Ǻ�|����"L���` �~��]�xj=�ۋOV��=?Z��Q,{�G2"H�y,
i������!������^G��HZ�ԩ��^�ț,ꈼ*�A2���8b	�7 r�Y/hP�"����3[v���1c�T�~+M~��@9����D�L'���乡��Y\���E���;�Y�����ْ���QZ�k��~��/8���"����*R��M��Da�)�H�*���d:1s�?�PKE �LBgp�2�t�nn]�^�6N���S��2�d�:�/���J�J�a�z�ï�lMT���(�w6���@���h��:�1)+	�Y�:K�=^�C��Q^F�R VM4������L���-��դQb1���se�?Y�n�.,xO&<��E��W�|�K�w?Zz��~>�\��į�ݭ�q�� &��M`�=x+���O� �f�	I��׉S� /�P��� `��!<��	|y�������T��TE>pĢ5� 
�d�u�23z�⩇���[����������r��
�;F�ڙ~&e�l�̨�?=�p�g��s�CMt��O
��M�il͕נ>�l�n�*�!�]��z(�	�L��>��������v^Ք�y�jR�/������	q�ġ@�Z�V�1�SC�)�^�9bez9�ES�k��2�~�I]�m2k�a�w��]����$g�)�Y�ڡZ$ƺ�>3��7'x���M4��7�;xSO�%�� y���i�B�;d謶�܋�	��
���!��:��"���� o\��u�Ҍ��I�X�0�<>�;]7��fNҪ"�R�+t� ����Wjظ���F�-w����{u�]ݗ@ 6	P���O�jU�1ٙ����YD�2z��?i�H�N^�Ѱ؛9�vD��@�NM�2j�1S$�X�k���`)��B������>��D�s���U����lOx�֒J�CC�PoE�G���kCo�����C~ĥ�	~�r����_��ܕ�Cq���{�<=�A�͸|ܳ^��=�A��������]�û^��GS�N�'$?�}�l�:� `�ZW{N�,^I�t<��~|��)ƴWq�
ZA�I^Ը����	���2)���&H��#s�����q*K^��G�A�D^����k�0�����70�f���z+V#m�
�e�ib�����=R W�./��ѣ�oR��_�ޗ-�)4A�f�絭�˛q����!�ܰ,��?���fI,{��w[����� 1��'���o�|�6	�%���1�EI|"��\��1�kj��5��q��9�M4����ݗ(�p��C���o��9c���h�Xʣt��c�o/��Z�i�֖߰���db*�v71Ʃ�t-���l@e��U�y�M������8u��������`���E�jض��o&�&�D��K�	����>&��3��禾Pm<���p����d��mT��Q�Z�5 P���rG�����~�Εzo�Kiݯa[U��X�~gOvq4������d�05��MHo\2�R[�ּBq1�
DH��3�.��,Ԛ�4҄�΅��[���F�!����L$��iQl2���V4��Z]�T��A~RV�Ms��q�|�p��0p���G�h�����N�/�^RY��@�zg��Y,���x%Ns$�7U����Ct�(�(E��~���<����9�Jγ�i�'�Eۉ�D����Є�iqu�*�������ڵm[�j�(U8�V\Bݩ����P���{&�ó�Բ$�pv���x��M��b=�,& ��.+�j�'c*�듉_K>cf�4����rѭI�m6���s'�����ȸGژ�s���o�mT�3��p���a�w�����MF���ԟy����1s|E��DFwe4ks�M"]��9�jWV삞�H4֨q3�"�
k"����p����l�m�����S�^g�,�g`�Bϑ⯐Se��b��jh��Zy��MHo������Z���;q?�C�4\��΄i�D��ǩ��'u�,w����ჯ�,��o_)�ɒz�d��ԥ�=�h��:�����	�:[��"S�����0ʆ[��]��IF6������-��BB����{ճ���J�Q�X�]x���I�>V��qB����K1¦���)�K�j���)A��
��y��xp�7�x����~0�A-��>j��DZZ�`�`_�{����is�����#=~�v�M���`.O�+�em�� ��B���K�a�|�ڳ�n�zD
辰��ʸ2	���}�����G%&�{��%�9R[�7X�7;��pa���7� N]@|bS����|�6�.6��v�����@�a:�F����6�FP�HZu�����Se��\��	�)'q��y�V����T&��v޴���Ր,��'83h�܎�Hn8Z�^���4 �J^����A�1��X��ʠ�d��y7m��޺yK��J�n��l�slϯ���0�}#�6P��B����z����w4O"��@�Ì�\��N��.���~;���(��+T��[c�jSt�خGFϚ#t�uЀ]�>�F�6�D�*VZƼ�LR"D,v�~ޙ��\�)�R��x"M𕗨9Z����ٶ�5G�O����δ� ���բ��2z�8�P�"e;�\@QF�ΜJk�ب�&s2G�M.�D�F�� ���n�1�۱5��O���� /$��V��v�sQ���p�[�������9�F�[)�K�h;�2�10,�"��n�����krM�[G2+�Y�����4�	v�~i�B$ǹ����\�)LY��]f�4��m�De���u�6���,����dh?JUy�0rr)��!0`e��&V)L\��06�d��if&��Є���
�3�����D: �Q������"/�y����j k�x��Vo��/�v�D��7�A=y�a��P!���ic��\(�A����Īq�/Me�+�F��WKu�J{u��t�X��og*|�X\�Ҩ��L�����}�°S�l��Z�o?d\�)��b�_��6˞�v�!����,�Q�����������H�jc{E��#�Ѐ��泗_
Sj�n�$��8�� �fy���9�Z��ðF�ϕ�"hS5�v׬����?�-�w�[9}�D͓�G{`��\DM���-u��>V�&����R�8/�XهVW�R=�|ԥ誯dI��!��R�u�i������Q����*o�����i	���͑�_ͳ��_��_e���L�.\��@ˉ��#&cf�1`�S���G@r#�"lf�	�R��r��W�e��#�^�sK!L�`kmV�z;�/zS�+C �DFx$'*6mn�7/j�9�vk�U�q�z�\�k╴1��8-U�I:/�m�YJ��N~�y�Ԛs�;�D���<�����VT�p+��ioLQ�./ �ݓ����Ip�|�S-{Mm�)�zaӿ��q9�WcV�L���J��-��KZA����Խex��Z#�蘹A<=�񶸆V�����qg�� ��h���q�6�|l:��ׯbG׬�[�W+�02FD3b��w�\3���!W(�]�ݍh�ܐ��]��:��IZ3kkz�#��OC!�[e���*R�g�=��9t��>��Q��ľ��%�Wb�k���|E��@�����Do+p���B��oҶ��(>�B�uR�>�Qi�0E�́v�����j�*��j���7{�NG�=��9ߪg�ӕ�ڳ�]����!��)4I��3�Wh�0�QM�1�R�C��G�b)d���=%V\4���q*�� �����|��li�^G���B�v3�,�a��w��Uq��)�3��A��8&+8����va7T�����\ꐩ�Kz����ȿޝ�Pt<{ЈF��1[�V$֨LrE��-�=�t?�[�ώ���o�;���u;�[	��Q�:��s�u�٫�{�U���IũBI̊�
(㾮�|i���b&1a�ʚpA�U+�k�a��v��� `k���H��y��bc�c� H15�]�˼���������3��]��˄.���ey1�7g ���IW+b�n�{��6_g�&����uHj�����5�^q�᰼aw}Uʞ��/%�qΥ����+GT���������-W�B�~����iD���,�U�7ǆH@wJU�j\9�~]�b��{kh�]��G��!�c���Wx�Y��.R��N�Hs���T��CkD��Z�(O������V�e�Q����U�Q�i�t���g��s�(�#�=�� ��%6����p��b�����M�՜2g��W䴍6�+�ke�7R��-mjN��X&��@3���%?)�)'���]F'��p+4Gy%��f�t\}wt#lIFY*��,gl����,���������ٔ�y{�D���j �9���qX�#����!OZ^I%\��w8a10���D�t�7K�6=�k��sz &7j	�c�K� !m\�'��{?�����TM}Ҵ�͓Q�Wx}ځ�i�-P��E҇Gg�{g�}}7�l_6��'��H\;�xL��N=�oh�bc=�&�C�!D��(�|�y"�S��4
�!��z��	B�-���d���{�/+�ʂ�8���ܻ:/"�|��N5�=�Sǝ'YM���x��8��(�̙n!D��=� :����$���� R2��������bRG�f���Y�gV遾��MQ"��c��ϣ���0�x�1���
��Z��ݼz�B̪"W�K�O��U��Gq��)dp��&.+l��Wg�̔åz���Y��JU�%�߀2O�����/�����ND��5��tH5-~9xw�Оt�>�s����J��I�>M���g�r�Gr���0�Fj����s��p��(���N\Ċ.J���<�}��C�	.���c�l�ޏ:���0N���Ji#7�t�0�44o)d�	,�m|��j�+X�[N������/�<o�2�zg��B�?��W$qf\����I1�-H����s]�zCKy=��	��znw�S=k�H��4�3�Q��u�l��_�w��1�ߴ$BL�g::
�ԋ�C0^��_C�?��?�G�����Uݝ"��)IB%z�_zo^��"�'�R��� 3n��;��m�k��
��T��j�A�+��n ��V����/���T��=	K�[M�]-Qa"L>��Z��eɥ��Z.!�x�����;�� ���'딨+�өR�ܺ�&J�Ț��q�p9�@��+:��<Q�L2aX��$�&��q�u�����̑^�5���A�p�kKX����Ӿ�lQf�q:s�b3ҧr�����AQ�4�ğ��D���16���;&��kG�8���3�R�N��������4z+���'���ॐ�w�f��w�Z��$GG`
�b�	G�?�a�LÀG�o�>Z��D_������'<�ރ�TL�������i�:�\f�����y�]�U�Ü�������8+>�D��Q�\���;e�J�]AA����d3J�����뷽H�,N2�9�$�K���-���m�xqSr����U�,��c^��g�8��]3j�/���J<�?��JpJ�4�V�BH���E����e��� Iw�$����Z��^�l�H�����;Xg=��R�Cp�-�������D�`p��
��M�5�����ߏ
C �	��{-�ۡ!�v�?%��*[��B<��v㺥]��'C����-�~0�aC/�4E�� ��H7ώif�z�D��ј�趮 ���U^_�T�Ɔp�7�b\ �Df���W\�Tn�L�wl!���j�����Ϋ��4W$K�&�Ux�hN��R�������w�<,$�n�D��ή{��E����2j��Y@���<?,s�v1W��SA�m�@��G	�t��|�Ś13}{5'D��:���KF�v����)�"��#�y# �i���=�F�`#w��S��\U����L���R��2$¨Z_��ҳR��G�܏��'�)j�ޭ��)�6kK�	2��l}��{�y�F�����Э��B����"fe����Q8��1�2C�C�i���X$�\�W��[B>�?��׍tqI9�}-(r�t���7�g9ĸ���X/x^���s$���\���Ǩ��\����@��SY�-�z����,�i��zy'� ���!��-S��n����C�z�[�>熎A/Z��9~��p�|���v���]]0o��}x||c�[�7�U|���{�bF�����Q"�e�$e�����J���-�wy�4_|�]��7)�m���؝�L8�%�O�p��2�k���|+V�Z�����h�y���_��nGygx$\��t�[9D�o�R�����`��`�Y>_�z���Wji^C"n���}�=�)�=���AwL����zm��=V)g�_�W t��(�� ��x5���5����5����bA�N���
ϷV�G�,d��v>	@�v.��좘'v�`��d��W�.1I�3���HO��7+��wp�5�;"dG�^`�%+�ܾ�!oڒG��*ū�w�92�/���	
�M�����K����8;�Y�M�W!ao�ǰ�f�~��|�7�J��G�hZ�<����m�vC	�2�q��#�F�<��Kߩw�����p�m���wF��s��IP#�ޢ2�P��u�����rbV_���9	mq%��yY��R��<ʣ��:P�[U,˸��ߡ�}[�p�
�Ϯ�}a��T���Uv5��I��D�)j�.�����%�m��'�cR ���ڒ�WF�&�'A.��é��=��v�Y>�l<��"{�w%����C_$2V��-#D�-��M�A(D�Y��x ���C
K��G�+�-��!�KtZ�e����d4G��A�4�S�#*u�R��liip�5����L��0�~f9��f�1�0,����Jw��n���f��0�\V���mǐ8�h������w�<���f� ��"R��S���|)�%nH�^�U��*2��1�=�_~w��;�}��`i�J�Z���A��Fj`*����	�ٓ-�!��*qj�>f0��(��rV~n0����m��5!R���#��O{�
C_Kͻ��O����,�����<D��u����Ǟy�{�ݟD�;f�8_�9����a�ab��ե8�0Ğ�:�qC�`%{����M�_�+���b}����{.��s��ݍVC[�:�,Xg5�p�V�i7�M��S}PG)0�O#��T�'A����v�g��^l:�X/?q7P{X��A�������T���h�{�����tN��^���ɝ�q�pP2���O�g�D,��<{Yڡ�pDY\���Q�T�����t7�r�5�k3>�X�S�$T5s��������I���-��6�r�do¨��C����7*��W㥄o'�c�󓽌1��D =��<4`�Sw����l�v�{�R�~��#�5>H�����$
i��G����.,kX�Ia�@Chi&S�Y�0=h��e�[��H�p�y�L�E=+�38�t>�f�D�! i�kk��q�ez'd�c��+�~l��%��"��)�V���[��4��_��	�ۙ��� �A9�/���0a
�`#�~	)�#*�>Fh�Y9B]��|�#ZNB*���P�P��r����������#��ܧ��
^�\�T�(�i���,I�Ei�ht�qᎭ�� �L���x?Y���:<�?�2
�%Ut�m[�L�b�rp9N%�����h�%�V����F�r�#���� B!�8�\�	�l͉e��:=���� ���`��g]6�n�D�>�)%�#훩HZb�_���B��{��m���ߣ�T��mz�SM]�`{��oe�_zi҉+�X��[���E+��fF1$b�&z�8�F8܊���vׁ�ֵ����h'��C���F�3{��}=�fb2��.9�E!e�@�P2$Uϡ���vO����	�����<�aibB��}�FC����mS�!���!ŦsOǓ�Kʪ]{�Ti�9�G��ry�Kl�U!©˂��\]c����w�]��8&�֨�W�9�2�Φ;���.�g�0Q�S��*�iÏ�Z_6=��azLiOv�Am�c�/�{;{E)��7�Z]h_Zu�/�eL
z�dg�n ,���K���Ԣ,���8=��O�����^����On�D��8CB�"�uD1�	�H�[v�$��i�RRk����l�y�*K;E���e����D~X�Zh�ty���`�G���Fp֚��`�E��~=��i�:�+!)�d*�=^
��jkGΓ�օ/ߖ���WBh���ޞ�Zƅn�1*A�e��͡iC��3�.M�i� �;�0�A�%�=,f������!�Z���iF�4I�ӫ�E���⎪|��(�<ơ+�C0��8��i�@��u0g[3����CJ���}���b"0���,�ѷ�O1�5�����V��Xr2����+єUa8���W����`A.ޅ?���\�#	�$���)���.T�A�G����h��t��n�6n<a�ᵮ���f�kK�+._�gV�}n� z�p�h��<��sޥJ�AA1��kHS��p$D�܆Ό-�b��J T��$<���)&�A/�P���~6��wp��T�.�m"�0�&��v͊CM��S	�ɌL�7�8�4�����h	n����%x��V�kME�Nיn��UVDx��@�Y[o��	?(Ȃϭ�����&b�� Q���,C��ձ[rUb`A�@>�M������s�I���S�gl�E�����~*m��6�n�Y�ӊ��[�$�e7G�eF��vUx)w�4�p@��)BcJ8�Kk��π7J� +ַ�"��N�3B�>|q~�4��ɪ+(��]!5��`���ķ�Д�'�k�m8�)��Dbz@݌K��%�����+�Cw����f��-��>|u�l�X2.{m|�T7����i��F�2t����*�fӵ�"��{�>�ZDmSs:x~r���
#��Z�D� x���1b�}�Ux�a {�m�:��z��4���]�9*}�b8/i�:�w`<ev��1#�aT�B��iD��}���f}�GW�ugot�����'sf����<۝�*���v;zJ�Jq�m#�+��@����#~(I�Y��N�7ro�%b ��v��}�U�R��~�ʯ~��oO�(�ȟ�m~�+0F%8tߠ��5}�v,�ߘ{�j��*z����<��kd��h�0�`�o)o�G龛�Vy���+�9g��\�����䒿��	���0m��u�Хʷ��z�� �露��+/i0E8�W����*�@�r6<O�7.η��-�i/����M�´�v�pJD�&Yؑ7���t��-�:�Vh31�3�J5Ph�lk��3�	�]�k��@	o�f����VXg�w��n�O{��l=�6�(��4H�+ �vƼ�5����#IF	���7@>�r��7mn�M���q\1�>���,R��PĲ��r�3�#�+a[�7X�&����7j�E���.�=�K�̤���\d�.t��h֏B����f�����0
�o���F\L�V٪��q�3�FIRk�����R�;�9��>�Z�	S�Q0v��'ğ33l����?�w�J)�!�.7��Z�T��us,V�N��n�2Ks�:�]:�M��TA��"��,�1�z(/��5�w"�׭�c��F���R ���pb`EΞ�[t�
E�
裂a�(\(�Ral�b��g�^��erP����<��ٵ����k&i�Bv�V��I�ЊHQ�rO�7#��|I_�a���X1�DDB�N(�հ�Q$��;}���_���9��ȷ�&�U&�J�h�9��;!(�-�w�J��-
�Oі#e!�L	�rw�<pc*�:��?t��4p[^O��'ΟSS�yp�p���1�,� ����b�-��㯥F����^G���ޕ�[?]��N����zX�ԭD�5�T��~!�v!����S��Z#�ήA��R�ŢCY���&3�eC���"OD�o��0��x�j�c|#�O7�O��!,�����-V������YR���j#�Y�z>#OR�Y�5���X~l���6jU���Q]	Gv����v`����xR$�P��zG�]��tsa�U�ˇL�����Z�H��e�F�7��C��컩n\G���Y|睢D}k�W�.S��9JF7���ە��!dGC������7���}���?��F�h!��0J7F�b ,�Gh���y�5����Ӯ��/�/?S�D9Ʊ�ff��3=�>PD�?�S��%�M�4\�Ր&�e��'���k0o�Nn�x/r��}�rJ
ê���:�1渉�K����w�Y4�&�����Y5b+ͨBJ�*�6?�f��{���+A���lX ��&��z1JO���!� /Q���5�>0'ɸc� ��VX�"�DQj�	�@�:[�� x����[��7��#�:}�d��b6K�}҆_F�F�����d�)�GP*s��#�����47R�t^��J3L�w�����ତE�Q�s�ȇ��9O�9H�@�8wʚ��G�%���c����ᅧ0�>���L��tK|ް�S��V��n��P	QE���.�  ��l��Nv7�6����@���2�͈7G��鹮#k�����g) ���*��XX�u�o+�f�?<�qPj���%�d�)Nk�g��?�3�����Y�&�Cey��F0|K[��<�⎇�4f0D��֯o��nDw+嘘�s����3I��dN�;���a#����&c�*tBZ!�: Ds%@>kG������-�e�������T_u �z�d��$�d{!D�wK?�ki��k�d6rxj?�k�!��aa��,u.��
䴠m,J:�cHg����,ǀ鶁�����f��!�f$�<JV���h�(��g�ͳs�@�6���k)���	3�XD	�W��C��V�X)=y��u�Q�ht�}$Ƞ9D@�ӟ1f�]2��V���Ӌ��;�֣ֿ`���7XK٧Bo�ư���4]p���-��]�B�+ԦZ����q���|般��NЏ��F�,����:��ޫ�[`�f1�WK�;�VTRF��z�<Ď�����t2��B%Q��]�gC��t��f
58f�)G �c]�w����Mi���r�����z��j;
��K��k�8Qj�����Y��(�<����h5^^X	�  ���u�>�߭t������g�x-X�u8uN��Ty$7�"�wٔN��Ф��/-�14�\���z;��:%��2ȺQ�k]�A쓅ZL��f���nx
�H�?bvvT4�(��P�r�B��B��ߪ�<y��~s;��j�"�����05&s�.�^$� 6m��2>�O�)܌6����d���q3�v��ET�0"
b�=HV[�ׅ�I��5L�评��9H'� ������T4�ܩ?�-o?/��q���
WsZ�=D��6=�s�z��Y;E��G�Ny��,N�(�Wp�G�F�J"`��4�(�`���'�:��P贘��h�k2�ۈ���%�{4�p�=������I�{*� ��V��v{w����t���k0V���¢SB�V��`E���q���c�Ĭ��e]�?��<�F$�62�*����	Q��LX�*��c�}sG�o��Bt�k+�Ѫ��0�d/dV�i2��K�:��ҡ�o��IS9�r��
ŸK�o��n���ܑj�����d��ǹ��Kgi��y �s������b<��K�WJ����÷�(�U1�9���q�v\�A>"���S��y��Q�x�O�k�EGˬ��7��@:*�P�#�꼪|
Oӂ�ui;撠I��d@�	�_)O[�In��(�ct.?��*�ū� LT�7m��M�
�]�E�Ĵ�|�L�آ/��?�
f�i�j��\�EA3]���3_��ـv"���WF��f�&�r�=-����;���V���-��>�s�<A���4K��-����C�?q�cg	��tX��	J"�􄃉��k-?�CO�2��h���Ǧe;��p�Hq݆g���.x���ǌM���)2���C�@,���t��k+>�y؄�������~� ���B�W�|C��<��Μ�)���ܭ͘�,�9�|
f����Ybf���T��o������j�o�*���+�8LȻqWPm�v�F���/�t�#����I�,hIf�ԯU:��^�=�5M�<��5%�e�lO�$�3���:r�ZE'Mnb�ӄ)��+z�A��.��~@Q	��9������b�ĩy�D� .��@)��m�h�0,�ّ�5(
���[��Ƨ&.{D�yX$���Eor�}���!�A�������7*nUD^������8Ϳ�wgC�׌�@��'�S�7 roD��^��pgy����]%���lJ,�OM���*�.p�� G����t?�b.G۴�f�\����>��R���oC熦x��#=v�J��"G�Ì�	� �i:2���x�	 r{jj����}��Ӏ�ܫ��!5��d%b�!
7��� �D�b�cH�.D��o��h�cj*�*<��|�A7g�fP�ZQ�l!�XB%��m>� !���V�Ԧ���~H�.!
���#��v-_@c>Ɗ��&yZK&S�㕓�#�A�G�AeM��(���B��w=Υ�;�i���S,LB��ɽ���cZ*!�-��!W���Z].�hzH�d�<;��%��\��{��@�S#�i�,)�i)�r,�H�8Y��B��ؽ?�2a$:��h�=�/��Z|��G�X��7�|����h�*�<��;PjI�/Gg�s��*�SMp �?;u��d|�����ϝeOI7R�H����͟6��3m���ߘ������0��&�G�c��� ,YD(���j4��ϔ3���m\�;���Z�
C���o}!�j�vǌJ�f%�c\�$&�r�a�U�j)W��"J���QTY��\봚Q�[���	�����+��ϠY��u�ee�g�w���.�!Dj�������	����d�C_՚�����B�JX���&�Y�׍���n $d�R�����i�/�L�����M7��N���%
H�i�8�xm�l���Bo��)a��f|��7�b����+��=�=(�6�G$h��[�	T$;b�����3~�z��QRZ��!o����p@&U2ⱄ�Xh�[�C��"4����]!~�<�w3�P��?�^^�ه� 0���?�ؕ8�>�m�p��1xaV
��D,-���Rڒ��'*s����å�{�Ĺ���z��_����0b�_�cj��z�@VAQ�\��9��ベ_�:�%��#~�7ha�( ?N���z�a��V���w�}姈�<y��U��Uf�})����/�Ƿ�G�Vt.���w�$���QP�'�ǭI���v}���Ny㜹?���e��.���$x��E}|u-�-ߣ��F{���i>�dg�K���_�Px�b�[ڸ2i3|E��|� �v������I+�kĈƋ{���r82$�X"V�n��sN52��0Ҩ�|�dB���|��G�2�36��
&�p	Q�ABi�� f��ɘ���Y�֥�S¨�=���D����D�'`ډӳ��*\��b���$��R���/gB�bP�A�t�˷���n��� ��[�X�N6ïnE}Ɂ���]����8*�|���ҽ����&q���6��O��L<��E��N�xADM���t���Ƚ�2Mܫ�V�NJ�����D���.ct�u���n�	���q���x郎7�%�$]��X�3έ�W����n\F�xy���^�V����,;�SP�gO���Fd�j�]&y�1U]��n��y�o��cY��T-=GI��Ȅ���5O0�nL{L%2����ͨ�i��#t*���V�n��Y�WH:�]�Q�����$�I��%�Z۰� �^��[�Vg�u`F{���q3��'�E�u4W~����w<�~� ��,��������,�-F@�+��>���]��aG{!tq5櫯��i���
I��?�f4�<������	88�'Â!�:=��\�-#ݎ�C܌���%M�ҏk/�c��(�|z	tJI޷��
�c<���=\�ٓ#]�G2��T*�X��ѡ�Q�r4�q#�-z��C�@�OP�Mk��%I9>��[��5�b��R��Co
,ܠ�z�_ԝ�'FJ���s��B'�����(��׮���ѳ���c�m۷rҰ¼Bt臾� _�Ҕ����� ���.r�*�����@'���MG�z!����%�y�>/��p�i���.�l�ij W]h�RK���C/n|2�]lC�V�t ��[� � ?5*�U6� ���FxmRA%a�����S�a-0�%���:���>�еd�v0��t�����y;B{����^AG?�z�J��$���TW�wG�/x.jǻ�*~mƪ�ol���G�+�����;Z�{�x��jDS�G,^��.H�5
���� �kQ�2��xe*j�Ng!�7G��Y�߅�k�s. ��o^;�BFM��<EG��* ��mo�Q��v�.���������G�� τy��2�z��</�-6��0!��\Pܳ����C�Kݕ��~1<��d�[D��#���Vu I��^� E�SX���y�R�����j��B@Sg���ϔJJ�/O䒻dR�^Xawȯ�"zg)M4�67ƒN'VÎ�����MI��tj�(,��7u�T�� PjS�����]!�"o�Z	���
R��\C�a����������d7�6tOE��u���31J�&V�kdKߏ?�-Ab��:�����f7Y��e4���������4h��^nV�����[�È�	o�D�Z	O�����U(�Hb�Ç����V{�<�Z��;����)��GI��'�ͺ��2�Pɼ��?����h�C�w��^��@���_������=�Q�OO(&1���|��v؟}ȩ>�.7�������&Y���)l���y"<&��݁��N��S�{����H�k<J!��J ftd����l�VŻ��9@�����Gd���7i/��M7��z���Dn�i�KJ���;ďy�����!	h'$��t����\�lĹݢ���ғ` W	�6���dHN���X�I�'����
 ��L�*�b�G�H��Z��{ n�ht�[E)Q�6�;w�Q��fԖ+b��B��rW"\P�s܋�]�Y,��/�Y���W4�PZ{�4�J������\V�K��uA���Z,f�t�2���cw_��{cF9� &zˉ�8��˹X| �<�Q���D�-nTʔ���!�ր��Sx9*�����AV&Gs(H���G�ǅK��U�0ک�)�4-��4����99�.�'�fj������J�����2�[-�+��cs#��m���\��z��:x��3��v�M���0�uP��3zU�H��{��t���$bȈ~�.ep���dF�B;�*�.f�8��0����b���������8<q�>��pW\C��~��K�M�3�*��b�NZ.�����EjV@]I�=�����R�hல/gl��쮙��6DR��9T��6�/6�Vɲ�$���N���B�ڷ���&^�=}��g�8L�n��8��	װ�!�?_�f_�L��=��3PKR`����b�F����L.��1�l�f��NA�r�+4���"Z���mG�lگ���Rk�0ۋ�̜�0�<�p��HԧIU,�V����oKc������L��5��V�c����Vh��T�;�Ys[�Xt�-�|˯.i�򌴬_���編,r/�9igd���RK���"b�,m�D��ǝ*U�݄}�?P���ӝ(�6ce�0%G1�?�����˱>M\�H��=�sg��iUM�.�JmPLq��N��k<Ћ��~w)�+�;��q�2QڞXkk��c��*lp���E�G��z��Bz��0���X�h�yb�Rc�v�I�8}:}V��s޿�BRF%Mjn�	Ԕ<���X�}缮a���R�����"`�+�6��1�aƆ0,;h��wc��f
V��SSb�� �E�)M w���P��B����6�^�1k_�*�.�`�NI���7�8P��i+F��\]�Q�����x��#]�UK�!͹�9f����湸��z^:P�1�M�1)���eZ�"�z�?��r���5���WPL;M���E��f��@M��E� �5�}����/�Aou�L��lO�=�[_spR2N~g7?�_�X�5cJ�S4����i_�sсō�y��+&U���ە�\�[=u-���zx�&,�����^�_]Lz�
X�j��^��yJ4�A᭰�D�.��nH3i�dY�4���lA"�D�n�L6Mb�	��N	+ThC8�P�c?�%5â_�[�x���N���{"Ϲ�3@��\��*mPH ��o�J�)j��*��z�u�.�E��0��MG�i.�ք�����gDzXj}�>Mt{?��Eͯ��Дɭ�4#�1�����|
*��Մ�Qd���q�ب���ET��|85�Q;~g����f�J�s�l���bX�X���|L��u@�BrS	�p`!Y���o�5t���i��l�!b�t
�H�%Y��$8(3�'E��2�/�_�Ypa'�C���'�x����	i*�/Ky����1 ��6������+��t��W�J}����׵���+;�t�$bk�^��z�i�0�P.Ff�*%� �������P����:�h݂s�R:��Zt{]��42<G�g@=d��	��/���t��&͚��eyǠ2_C�ᦿ*��y榡������24\����UX��Uݯ���탃g�EXhul�Zlm�W,p_�)%|y���`��^����O���=��L��}�<��Y�|��+<Zמ��<����2�pPe�>tq��P(H����u2�8��X������݂1�9o����x����75�,�*����)ۦ��TQ#yʡ]G"�l1��Ǌ�@m��1�l]�H���NgY�Sq�����h��9E=��Ey^��ka���_4�܍�S�=��H:���bP	��w*M��^wl	�3�A���!9�g٤���#���O��b�\C�y~\=�J©�:3�y���~�H�GU�s� o��x�3�Ug��b�j�bؙ��@��+��=4��x;M5��{�;.`"��n��V�6���B����²~�hf�$�?BC�a�X�|Q�p��ġG:��۶m��T!h���̮�%�eN�}rs%\{��wn2է�G�8ኗ>��]鰧+ �����B�2���0<> G0Z����mW�t+�E����!�ɾ�
�϶sc���0$C���o�?P�<� �%�+���Ԋjrp��Nz������kHMG���H���,�5�Ý>q��L��|`+�����E)�yĩ��������-�w(�0���Gg�Ƞ�[�Tlb'����h�=э�+ʻ������>��΍q����bv�._�wr�W>� ���fI����V����J����^����8"eo�z`E �����S �K�l��3�����
�DʧĖ�$�j��:�r�kИ�u����� se�F�e �V��U��qu��"�2*z��F�2zMb&X#��-Թ&��4r�S6�d����z����2�UZ��}$�<��S���5N��!/W����2��Nv�IU��}��v�s��PH�w�m�G�Ɣ��g2���R�7���W��-���F�h;����9���ډ�P�=3A:�$R�����vA��S|-��RA�Y� '|W�7�9J+T��(G�`�-�t,e��*��}-��={܁����^� ��z$lOu�|A[��<ڀg�I)�pdJ8Q�9%��2�Y	�j�����}���v9n��_.��:�:^j#�Q���!Gc>�Y�p�=D�����������ԙ��{f�}��`jzl{S�U�L�ss�'ķ��c@�b��}ǓH�t����G���6�2�q���"c�����M5��^.4$~)���_jXri:7��D��Q�WxN�,��=U���c�Q��=��ӱu�	bbs�W�YuƗq_6��ۿ�IF]�t:��9��(<f�`�W�W�)���a�]7� |�^��N�Q������&��v��R`��B�W�W��@��)}ۃ�pv9^��~I��]U�p{�|A�,��~9?:�����£��+����S$��ra����Ņ���If&���S���8= ���q�ҵ���-z�9i�2�Ϭ�%�}h�|u"�a,�`��'9�)j@����?�Ǖi�u���Uw��kH�I��ǵ�4���Sޯ�{%>�o��\�A�T�27���
#���F���������?A�.�"��m����8aZ��Zsk��A�eJY���q��+�u��`��qE���	j�;q%-�����ia�=nDr��i(�&����Mp���p��Itcd9n�Kv��-��/ ���Տ�Nί�q.<��$ǫF�^}�Q�����e^��u\D@�x�}�)#A������9'�l��c��t}K����t"R���r����i>�l5�_�|��I3�B���9��H�o��B5c�^7*
���rC�X���8q^������L
���E��V?;��r��3�?�&Nt"z��c>�{b�Ĺ��m3a�ϧ�:��,И(�f�י8�E-������>:N�C
N�V�E�����E��~x1a�e��eT� t�(�J�5�����'41�A�'�ܹ�?)��,G����zW�&�O�p	��p5����-�4�k��lx��a�4.z�*���9�*��7�ׇ_�~�w�uY���vP���n��I�w�4o�
�\ɚ��c���HWj��R�8�?=��K�����VPy�x�w'�_�����p�"
 ��bvC!�~8�}�O��k���
�Y�ax6:u|�U̕�#����黽��W�	�1�<��33�u{�q��͐�����0����&�S�Q��\���d2�8EQ��b�2_	�ŉU��=/��So3�LLm������3�um�\3R���Rs�M=_���]��ckM����+~�6J|	yL��i[���SB�K�<��i+���$���2L�=�z��{p���k9�.T��.��F�M�����]Y���n�٘�>�g�拒JoQ8����E�W���<G��%�bE	��R�?�8��P�n��0Ԕ3K�
�V�1��.Ǳ�=�2���z_�<��=_)G=�[e�:�������H��YQ��B~GZ���Ke�L�4.%�H��$M3�v����5�4���4|�mHq�u�����Ѣ�	��HY�L˹��HNF���%��we�l���A�a���g� ��2�HR��^}�Y0z{lpqqte����)3«̹��m�^%}���9ɇ��t����-M:ް�Pb���+��������B]	9��eM���}r�`��D��a�G�-�r��#3׊6Iw3�t��1��Ȫ���5�]�p��Df�tv57�<��+�r>9��";�r$�x"E��6)���=?�-�p!���,H�y��B��)��)t�ʵiQ�0�l�(u��
�G)l%I�ה�*��~���#=0	=]GL��p�ӎw�M8����8o�����9�E�pF�l`�%�Y�B�󶋟��$��~s� ��-1�FE[}/_Lj'<Z��� D�7Kuy���e�l��_zZ�ޕ���%���A�acNٶ~i6-��7*�f�6����/���/ۡ�̚���a��Ǭ�13�DY��u7> ��?��7�ǃ��=f�m����|wy������������B�:Ė?��Ё! �!�[A�{����jU*j���pC,�.�>�De�m���9"�6���I�6k�mPh�P
Qy�.�:[����"z�&�nz�Ý&ܭX��l ��1@tS�}t����e�Ԩ��>#��&����ᾣtQ�0��3�)�����t��n�{�q)�r��7�*k����C��魢�6�gF{;0Ĩ鉌d���0�J��ν�"�����`�5���ܮ�k�oH;�.[e@zr�Ǩ�%�V��I�9�FfS����8���҇t�p9�"�l����=%�4[��a~����*�����gkt်=�. :�n�!�Wg���~�X����2���7gL/V(t�x���A1��Y��N��7��WHʭh����t[4�i��3	�4�&	Z2N9ğ܁�Dt�U\7�)缈��4(�nW�P׻����7Dh�!��Wۣ�`]��u���9(���u	hdJ�㫄4i����"�Qba0��z�
`�]���� ��aw������B��~� �P��9�����~6�w�
�����P��ϔ:�HN]�<
/���S��I���_�
���[&pf��������=u${@��F��0cb=Y@#����P��X�"���ܹ�m�QzC����=���^N�Q#gR��X^��e�r"b�P����@�e]s�����E|.[��/`E�ޏ*Lvܙ�����]���OB��γw�idf�4�jj�1��L*��ŤR9Dլ<�y�h�R��mlI�ȏ��y��\`ۭw^O��)j*cM�Ag�R6�S�_r\킹
��\Gc����9�s
ɑ;Ѿr����2�|$����Kӥ��9Bra��14k�
	�'$8e.�~���Jf
�qFv+=�� Ȓ��Y]aæ'�S����hc�~��׵��T
1���؎��g�h�}���̭G���G���Q�� �`sY1]l��+3W�~��Ǫ�Q����H�xVV�۱;�c��g/1�����T�qn*����8<�!��ɍ���"ߪ�=��+�d���*����}�*᧫_W�ӺsZR���z��n��![����@>z�9'ڪ�i��ݷfD��5��/�52��H�G�M�lSWϖ�)�Y@���BX�R5Y>��d�^ủ�%�MqRdqV���2M�0�@e��D�+	��c��nF*��`�Ì�E�tƃ�o���Q�دL=�� 5�NM���nGԀ4���Ļi��E�\^�3���Nk�r��X<{��o@/{cO�9=��OP�Nkay�Cy�[���}G�Hj�ɀZ��D&]b�j���惹�BЇWu��ٚ�E>(Ѕ���i�%�j�9�"��Fh4��H>T�R��H@>8�}����4��fɾ�"�^�ȉwM'�DJ�e&m2�"���k��(�X'�i�vn7�Џ6<6[�{��̲�ɜ�?�dùzL\��o�a���|~��+E���E�%�tq��iϨk:��y|.����[)ӻOOs����q<;0X+�64~���k{IG ޓ`���\��x��;���-szݗ�L���u�x���|:~�	A�2��x���l��y~e:HSG�k����_T��Nba)���d-�US20�D��� �<ۼ)�W�<��=#Tɥok���B�l�]����qX྘5�W�c;��K(�}ܱZ�k�,F����zb�?�z��A�O�Θ> �v���p��߀[F��;N��߼�r0y�ι���&�fL�P�{hLt�� h��k����� =_u�oESM�`[�R�P�u��Z������+mbA���)	.�`(��I���
.��S�B\ã��R0sK}ͣ��BE㲝��e��Jhsg�؍R�u�=�~�,�/��]�u�^H$C��Z`y�}v�Og4c,��We�znWg���_��7�WG�Y����a@;Ԕ�ݭA��@c��稰@�"�]yg�i�4���b�%�1�Y>LZ�&<7����0q� G�����qP?	�4���-�B�:�Y9��iTS��Ȗ���k@��r�U��%^����Cw��ɌK����cP�m5o�y �|� �bN��X+�}ѥɦm�+SΜ�#z*נ��/V�B��;���o�,��n��?����0�����7�呯t}����Q�t���͎c�2v�/���ܾ����h9Y	P��<ߣ�S]��r�I>�YjG�=�M�S�#{��o��6{�c� a�\�1�R�rd�1���K�k��TԽ�Lt�W�o��U��F8�~�����[{,SК���򋴪,|��3w��!�V@jm͈J��k�Nq�g�xx��'��r�Z�����y���������RTX93ځ����=>'�+����m��Q�G�";�Nl�e=���f�����]�� i|,��l� qإ��:ә�IL��g�_��5��;�6��Gt����g]�$����<W�/³V�S�ǃ��{ֵ����B�4���]dJ�:�)C2�Ӡ9��i���Pn�$rR[����@��Pk���J~3�[����ڡ��a��~���N�R�!���7R��ʅ��r%�kk;�����R�M�3ȁ�Ǵ�K�X���E����LN�^�g���`wS��>"��NM�n��:�����bF<�KEO���K���%@� �=���M�Byu������nt�>XD"|�K�\-���7<�k�<C �b��?�qlS������fأ��V%����FO\�+4�����Żb��>�T�d����u�ȉ�J��]%��gn�K��$�.�G���z��u�AJ�ݰ����d⤍+'�%r�\'�Sю�k��q ����+����w�dR�SxͳPoɴ���ZU6�$n�k���4 [��D�K"�v5�k�����A~�e��&������{�����8��W��|v�4��}�y���Xf
K�"��}^\�g�%#��4��\ܢ�����W
�+{9,Nϼ�9%l�8����n�r6`�͏�� ��S*���D�B&�����5�_�����/�\چ�� {L����v�m�k��ތ�M|o��v>����s9Z��ؖ3���z)�1�I��6�7�,x�},��P�*pA@b��2{�VY��qe�Ao%�n�����+z���Z�EJ�NXm]3v(Y_��yC��Q���2��I�Ë�U���5ی���2d<B�u�1"�?�'�w����������g������9{3&�B`Q���l�:uh�l� 4
��p�̩it���R�
�U���pF���N%���D���ʻ.�礓����=��[9:��(��/��� -�࿰ &r�@]3~��Z�t�҂J�4����i�h��r�`�*�@Ms"éz�t�Ժ�ҭ���h[p�Mc=ڔ6sj}y�Do3l��-��Tx�u�#s���O$􉤋�\>�d�좸b]�G����~qey�N7u�\��F�g�}?4�*�Θ��7�^v����_`y���"e"V!��ë}ʼ��쐵����]��a����|w��(jd|��-a!��y�N�y��S@>�^#+f�����9<ݓ��މ�s��4��v��	CG�_�g��H H~*o�_N��u�CZv�{��3_<��_�I�q�O���*�|
�>��?���7{���,�)�iю��Ľ@U4f�\o�(�mɄ-�Qu���@huy��>]�а�)��)���)o`ga���zbG��[�@v.It���ψɯ홯���W�8�n��:�M&N�@���@Q���I���.ؕX�'�S�!�bBl���dy���ƞ�8l�ç
���Ư����xn�&�p3�;��3]�\�@5T~C:�}_���^��rG�Bc=�~������{w0���m<��%ז8}�����C�\��苢�٨]�g�/}���+1�WS Yd���y�a�����E=���P��"%��,@\	Q�\��ؘ�h�J�`��$�Z�"CZ�u���CFy��4���qwb�C�y^)�Xt���$J�!*G(��zݜ�x�k�zL̓*�/��5�q��|��^��@��S_U��ŉ,�t�-1Pt�ۣUT�GYvO0K�E\��@ϓ�)�A҅;��FY�G��q�!ӣ:��e9o� �A=�7�44�*�C9����Sr���Ņ 4 �'qN�$%gx0XrL�5�AgZ�����e\�{ZӸm�YYd�T�*��yب�WU��Ό&�Ϣ�ӊ�Z��ɰ$q��ֆ6D�w�LQQu�P�6�TG,�c�%�Z8���>���e$*RdH�7�������g.dй����#8b�\?��,�$�f3�pD��?�7���]�G�+`��[�UE���vU��4�HPLN��p�A�1G��kj�r$�t�^�P*�>�χ��_���(�pN�f2Hz$O�	L-�� L%Qcɓ��;:�=sH�yy3��TD i�]fҬ%�\F7W0���&�2�s�lN��,�K�>�31ꀭ�/����������O�}��̭m�$�����?=u�d�������h�Q��|G͋�&����[��H�@��¸��d�D}jR�Qd�"�&p�!���Q`������$	"��(�Ϯ0��B���co;C-Pq^&��v(ݣ��|���gG������>]O��9�F���Bni(i�N�ǯD�"��k�6�����*���N;�s��A,K�,/��D���R3&�bW��Jv��u�-|H����zb�v�E��y߇��(�&���19�ޘ<�Gs�ɚN���)�p�|A�\fa���?��z$Y��rs)�ËL.�����*�bX��»�`5�/U�IK��<�l����E
D�/[Cd$���pI]��èF4�錋>�D�-]�z�6�Wh�V҂�ƿp�`���&t����a�g���Z���3w-'3����Hk����v�HjlA�
��S>]]���I\����R0�����+��bh���qQ�a ,��)p�y����k78�K*h=0�����F�&�+�p;�foFYO"���YE���GE��d�Nf��o�;�*
�o�yyD����Y�{v�>]w�jg;Sa��5��J�>*@v����E��)�f��������4�m�^��!������5Q�"%�U��^�Dܼ"�����Cph�=`H�4�Wι1�z�%���[\������P��c&�:e%u�z��/]qw0~Q���O����ۥ5��Q ^P"�׬�0:ߝ@�E��c�w/�������Ȥ�k�>��kQ�����2���%=/�+��jY8��Y��ɒ�P���ea�T�5�#e��O#��y��Kkt�z�/��Ⱥ>i�*�}<��c�@k�D3��̚T�����Z�?F0���K�,��ʖR�l�beD*j'��b�����j�+V-m<�.�����(/h�~���ٺ�꺇g̜����RЗgG��-[ Z�w��6�a��c?�Wo,����;ل��)4�⥘n�F˲��*C�z�m�:QI�˺�~ҏ#>��8s^9�*� �^��9�p��W'�
9}h�M�'��H�I��y�RAUf,8�&.<�{�>�ftǉ�N�La9
�g�'��_9=+���J5g�K����Հ�p�3�lն�+ʔ���u�\��8���[��z]9�����+?^
Ɣ���]p#٫���xQ̂�,�="���`'B�\ �>z�m��K0�2��������o�����:b��k��(���ed�s�Ӳ�Xk�����6��Qb���#V�GH1����vf��S���h���_��J�^'��jh�)���V�SV���w��;4D�?	J�x�fe��"v|/.����#u�u�`��2���S$�嵅pB��k>L�7.a:gS��~���h�XΆ����]6���;�-,�Ǜk���M��b}��n�ZZ�b$0�?F�'���y���wA��L�~T��D�����?�+�[MCS�q��墶^��Uz0#+�3|�pT�Ϛ�A�7�T>�[���g}��9J��.��e��)��0��I�qZBz��\��9�ΐ�E�0U�`#��L��Wu�l;��a�7]�s�����1���j��F-���4$�3Ҙ����]�B�>i��m8h�G��Y:JV��(ڿ� �;P5��H�6B�x�e��ˆ�W]K�P�z�&���?6 �cO��L��v��)�<GD��5�ەf�t��:=p���A"��p,9��~BN%Hv�_�;���<���?���[n���D���� -��V�"��K�Vn�l�YZ�{΋�ӑ0݄t�O�e�q+�{1q �
�&�����`;x����G�U繫����̷�Qs��?A�6	�
�6	��t��9#�˺�Ŭ�]އ]v�z\��h�f킳�Y�w�}�NOȉkb�	�g��LoT��G�ڲ?�W����Cu�P�#���YڐE#�p��d��E}�����˛��]7:`���X��)�lT��S�t�#��+�<�Y�x�	2��j��Zd�ǅ�U�VE>���h��C*{�b��B��D�1۩���9w8�=�ɝSl�47IB�ưc�C����H�/��&�A��(�.H��3O�ܦd�t�A�m�̨�u��7Ҫv&�����3�9_ƌ��d��+��V��)6��E�Cyv}wy��mUOh��A9c`��CC���rf��9?��$��}�.wr�`uD�����6$�C]�;����ˏ
88�i(���q�]�����U7Ѿ
��^t�lP��r�Y��2��;�d�@H��4�~r����K�¿�$4�$ң����ח��}&:y���R'�%��Ks��"敍���6����W���~�,T��	�����7�`[5�Z2ժ�M0��46�݃@3�
1>�N��7� �1H�V7��ߪ� ��9�
l_c����|aq:;�|��`��~z�ji��|s`կݩ�l����z��p5���/vC�P�?|?.�>�y${]#�U�%M�m��*L��1����jqkF��U��m(`z=,��*W����ϧ6��Me07����/�5u��~0���ߵ*�bz�}�ٳB�@\�Xp��<��c��_"�>���1\G�f�v��,�l�:Z���-��f-f�^���	�|/Ю�ZCP	���F�'��k\�%m�]�ij�I����ғ
0���u���@~��D��m��-�Q����rnټ���������q�ߤ ��Ăuj�X:��y1���t��ʘYtQe9�
u�)� �C��.Xp�M懰��sm�zA�v���O��hm�o@���q��Z�|7�/*o1=?Z�望���J�`!�@S�
~���7��w�JLr|>�p\�Pi�KZ{q���s�"s��_�$��DYo��ÕvՑb��!E��9�0���?i�"�3A�����x{�S��b-8�y�ӽ�c��WD����Zo��9ZL�-�i��m�D� Ѽ�ƾ���a�<�Z~3�;�T)lq�?nc|�A�̰a��,鏄��E`��΅|��k-�n�i�2�;�aF7\c��=t�y��������(:_By��۠�����
@݄��Jִ�tK�@0G�Q9l�ٓ�)�����2M����'�H�U�T���Uj�
~c����L�v,�:��K��g���`z�t��k+`}�F��8���<���)��s$�� EnD?
I��t���tV��x��Z�fR��e�ZN(Pa�W��p;iߎ��M�0���l)>��ri��`�r��eNVd����t6��m�~h��H��w-�NԺh��5�x�4$����cL�kCQ�QBˌ\'��H�i�Yƣ[�h�[��+���*}��D[����;���0Asb>l���6BJg����\�ָ�4l�	O�r���{M���ߪ7�͖�rD�[Fbm���c��z���FM���s��i�P��N����;�9X����R.�G�{�@Gf��/MJ��S��y�B �����p,hq�R:U�	}aW�os�b)4�hX����-��am+3���0)�j��Zv��q쮄Kκ��-{���͗�e�R$�6�g����m}��Ӧ��t�W�d����%B%�iOF,���1�ԊT�:DF���u&��\�u�����ई��j���܅��(F��^��&�V��S#%w|-%bW��PO'ˮ�\F��ܼ��MV]��Lu�>2��_Ӱp�*�VA�"���>)�]�'��}IU$=�����y�r"3d5Y���������Z����p5�K%��c�j<c��+ƵP�d
�k����ckB��W�~�6�zWiC�5l����:Z�U�k��� ����1��8_p��*8ɚj�����]�q"���Nt���ɔ1����&N��8���9&�E+�zS>Ku�u?�G�*`�,��X���f�mЃ @g�n�Xm��r`���dKYԐ�H�2j�ۣ�xݠ����]�l��&1�Pי<:to�>��y���˲��e�V _0Z:�[`�����G���w�8vq�-I�4lg�}4��]���;�FJ�^L��F����̨"�~�����;����A8�!�P;�jip{ƆQ��:��}�#�����ŷx�SgbWzJ���;��E�_VW�zY_�Y�D�,s�j�	v����ff��*����IȄP���p��ץ=�J@��w1]4X1Y�]w���A��R�7�q�؏&^�Đ��f���!.����߉!6n��;���U��H�BM��YTo�,�$yg�?i�l$ǵ�
��I�ˈ�~w=l	M��#�465K���yt���&<�;P���&����r�Ї�̹���">q_k�F'����w	^I��u��m����UeoÕ�m������IFe�qꔉ��=>�;+ௐ���j.�l$"]e�(�����0aW����1v�꒳i��� J���B꥗�r���p�W�tJ��ƞ �v8�}�d0ϓ}@|�ƔN��YvX�f"���@��Y1
���ro5;c:w�눹+��*����g=�mI� 5���Ն͜�+A�}���e�����9���dچ�A̓�?�FK���F倕tR
R�
Ǔ��_sW�(���kLLnXz���$a�á�J�^�9�o��/0_�D3I"^R���"*d����zї���~Դn��e��ȍa<�!���qkB���^F���n���^M�&����C�������iZ��M���H��B�n�O�{�L�N8�"�[M���^u��OD�k�l�4�H��a̝��o�ZN�l4wP�Q�	Tc�'��;��%+(֣�)�EDlp����Iإ[̾ߐB�}���?! .��E��q`,B�v%E%)�3�+E��oM$��̌:tzM���[ �t��p��wnk|�6�-����܍[ql<��r�_����ī?�,[v�?p��i	��C�xw?Om�-zB����@k�i����A��ϟ#�ɽo��͖;�M�/���.�O��z)x�ګ�C��*�Y�f���]��c�1v,�T���*��<�T�'먀"q��n.s=��DF=6�H:�$��W�|�:9f'/��E
�t�,;Tq�������<�l�c�k�Q�ٰ�}�:WlN���u�� N�l��c�@_������*̱�<����W&�h��]�ݹJY��qZNV�M�aA��?��!�+vs�z�T�s@�`Jl���8���I:��7�u�X�H�����+0��d���r��i�M�^�������"��ݓ`���h�'�-]�l������P�����(��	o��׹c�,������V<��į�� ��\E�7��#	V̚�5�w�:c&��1i0JRQ��((�H A�L����`Ĳ�(a�Y�^�|�Rg�ւ]��q����"_8ȱ[�y���|��c���ފ�˳ߊ�W8��O9oO�b~m�7M�r�!D���y*xɑ�OѦM�;�R)����S�R����=�V�+]���=TX���e/�w���G�AD�Gr����i/��_���t�`hܜ��	|d�ʵ��96�\�B�㈉���ߋ.6]�0�d�|�4���m�JA_�ơ��{`�!ne��!�҃����(��JK�����>���5V�8�J}���K� Rf�P�2S9U��m�-�+�;N4��i��T=@\������E�ʙ}TRD�]�,a+���E��9�[�f扳��w(4�H���f�b0�0�
����C!� x�t%�:��=�q�K�RO�/�����ږM׻��9~��!�ٞ�!�ǷV��s�WG�P׵⡵L�i�������ucr���!�����A���F��9�H8d?�<���	Q��ɔo�m��Jux.WFy{H����H987TA iF��b�+�r[�I�_�Ȳ���S�w�{ 	8,�0eA09�b�
C]o�M�t�Bc��� �K�hi�Z7�F.��h�+��	�;�[夾���=_9���Z"Ò�����Ƌ�(c+���S;ț���I�.SC��/���1vY�������__y�J<@i��e��R�y�h{sE?z+��$^�;�S��Ŕܐ�!��@{�|"[��t�#��u���w��MͶ�v��xYo2j�<u��E�81֍WTaZ�mi����I�漘���
����"���ULɶ�%��so��u��Í�< ?+^q�'�`�IW�5���#gH,���̤��QT*Cʽ�&�W��.����/Y�Fb�:q��?�j	�>D�<��T����1آ�c�P}J�ɕfu�^K���>������^�fm6.8'�s�f�B�=�t��\��C��������㡥4x vq��xV�����^����f�v����xY�^�N#�o���ޗ�G�q3wX��Z�Ǧ�Q��;��n!�F�9X�A���qN|}cK�0���{�
J����Sg�g�Nc�ʿ����u��~�~g|����sC��Xj���]���6�`�)�5'q�$#
Я p�?�|��s�gN�ܦ�����Ӹ:�U�5JC��y�l��LTI��Q��(�~Ԙ����h�C^+~H�ҒZ����nD�+�Z�Ž�8(��z�	uRЯm��8b�:����
7���T����9s@������C�&��|*֔{�T&j�2q�<� g�Va�?��]r���r�u�eD�3�eݻ��q�O;��S}��vE,��"�f���ِ� w:����)>��"��y-S���7�%��G�=���y��s_��9�{�r�M7w�U����b91�.���s�Rn�#���g��O �y���	����	@|ݓ��O0������q4̲��Ӯ_& ��v�sMB�2��\�����C@��ϗ�k�2n5P��ږ�5��^����ω�Y�%�[0����A�#�u��D� �8�<�L�����.�E����t�P��r�S$�i_����f^#tb�h�H,�H�o"�<9Uk�Q���":��0Q��$.sz1�A���gtA����0�{7L����]�2993a��x�W�%(�;zw&~��<��U`����&���}Pћy=%��@]`]��!�YE����s	,��z��|�܋��0Rvײ\N�'P��*'/}<��xXN?8���8��gz���3��흢���7B��m�$��<�u��>��Y�ۉl��J (n�,����ub����PbO�������̷���CV\H�x�&E'��EN�0���\�����eUM��=�6�~��Xќ]����||\���ܡd�y��0���k��n��9SS����"C���D�~t9�闇��c$�ə�YZ~�/l�\��B;�����82��~j��`��eE#��;�b�[6�5����yF��A�q;��"��XQ6�?��F~zK��K�B�V����%�f)�DͯPj��~qA[�5[$���M��p	H�E�rh"�[E�Ƴ���hztg��W���@�T�0[�~��i� SQ��?�����j���?[>�o�"�Ir+��]@�*m�s�SJ;�(�j&R�~��+��eQ�����r�o>���8��m������1����� ���§+�*G����(׶ �:�װ�ʿ_"s�Rg�9iĴE� <�9�b�5� k�щ��$o	�@"����ўr[W����s$�&�J]M���K�/p���S}�N�Y��Y@��H�骨�N/P�y�?�T�$&9���Ữ�����+69��0 !� >j\�Z"8��Ҙ	CCKX��j�,�?�H�*�'׈�:�`z9�X��2T1��.� ���ʷ�r�����U�@�v\�Z	��M Q������胶 &Vb�Õq�2&��\��.qW����'R��{���K-T����(|?������w�h"5SD�M�g�'����>e��!�d����v�p�'�6r]���ƹ�\s�x���϶t�Z��J_j��!������;�-������"�<R��B{����򑦏�~�h]_+P2U���)��ۜ@��|:�gS;�9�X�z����m;��(�mr/�:�|��I#"d�7a�r��r�m�0��ɦDQ�W��Ԁ&T-M�d�<��HA6\�+9�����*�
�%9g����@����s�����]Ni,!�b0�3.w+[(�]�drt�V`��@t�<U;٢�u`�%ꞝ�jaD�u$�u`u�����Z�#Ug�.��d�E������W������V�PsRr[c�i�peՠ��.��� ,/%���c$~
�&z�1h��^�ʬ"�,�_DU�� ���)z��Q3�����v��Y$T7�i��N6���D8�~\?�AӨw��Fo��h�j��w^l�C���d��!��rǊ*��9�TȚ �FU���0��ɼ&F�ʪ���̨<sJ"��h� �O[�*v������DxJ7Y�<�L�C
�Ӷ8�a�C�)�P���[�>�Ť!%�j��C�w�k���j�_/ڐ�W��y(�4���u(#��w(�;i�(�c#����F�`d2?�i�rw^���^��oF�j�c�/~�9tsj��w�+�:L'��5���	�<^{Z��|�Ɗ�qrKM�9�ޱ9#��n��\٦Z% �yX��f{ؼL���b��*��
�P�ohp��k�~���7���C�gx�Cڕ>|x[�Ç�u�����p� �P�J�&�Ӧ�O� �z&�rjZ�6h�1�>\tߍG4;z�)�-M��\���s�3\�.��b[�X;�Y�����E�Y��Y���2`�R�ߜ����3�EN�HB����a��X-ˤ��#��S���s��f!�����n�LDe���<�Y��/�g�\��WH\���bI�=��T8/�('T̀;�[��0�)�{�:#]���Z߁����W�qs���Xm��%r.�	m��J�vC�^�1��E��~t��%i� �0"?�b�!1�q�ח&�WI��H��:�3��;��=����'�Q`Y��Z�Rx)8�1I�)-��������̤��8�>�m�A�P�=����(~���ܑQ����N���N��_ZZ �T�=zp������ޫ�0�O�x�U�~�(7	/nzj�Z�oR��uu��-���i�ظ��C��R��r�AM�<�v�aYi�.��BYl��v�����u��L�����L��^pX����Op�)N��7IR�S���q�U'���D�&y���yW/e��GM�0!�7�εY�XP�= #�=�n� �m����W�4le��f�����!��jN��#'F^D����?9F�c��Xh`Ґe��%	��]5��vrs�����ұ�F}4���<��|=��sÄ��B�5��ך$8
�������
���I���H�^�1�E�����_o��̍�����e9j{`����q�~\jg�՛@�y� W!���� Z�(�{��#�N<����״b�I	����XHH���>n�����WR�Djk9Er��_`�Y��� b�r���M����bެ�+b$G}�b&O�X�b���x%P�M��'f��R������Z_�j�������,�͸r3��0+�Jt��Mw�HW�ςց�V�g0$�$-�k h(������C�c��ľ<|Z�5���w(g�yPy�b�9ێ��4S��S�b��>Vx=B�Ǐ(K̰&�����Q`�+W��肐c��q%�-Hu���WI��^챙����S��>9�F�*�"��jD����hN����� �94��>���d���{��A��d[?���!�w���F�1�%=?:A4����ώ�������c���^�K:�QY�iO���n�&ƴT;I]�t��f���n3^g�h��*�Kz��}����
���Lނ��}��)趵s(�Υ�)��NL���
j8�$��J�
�j��@��I���c����=�&m�8���w'Uw��;�s���?�p`1�ؼ��	7�(s~ �[p$w���q������|�KQ`�}T�3�����9�t��~�c�r��f��6��n7�G�=��ȟ��mA|+�?�8�Tu�E��$��i��}̭}�$�m٘';�ZJ=�R����?ci����+bx�@�Ru�p}Ԯ������4	F7/EP�)"'��m4������$��O�R�U|�\�Kl7������l�f]g�s�I��ّ�w�5Phlp�n��}���&�L8�a7�r�k�>S5���Y�5U�E�eG�?��v[�a4\��W�j�e��,�zذ\Nf���\���KH�j:��y93�tH�Ә��{tf0L`�@� |4:�F�HӴ��s�:F���L���d1�����(�]c2s3�z��|�g��;��;�s4sU�X`?�#+�`��4&p��X%Զ@��ϢK��ˈ�g��g�`��T5���W-�:�)n��2l4����Uӭ���f�h���͖��IX�A�`9U��f�>���BP{m�8���O V��5�w��n������,q��k칥ݟ#�x�g��7� ����n�_BT�Aṿ�r����c&~��٪ξc�γHC���,�	��Jc?Z��㕫��%K�Z���cv+�<�`F�|UG<H�@�&�)��9�������	���7o�H���	��	cx��V$�	+w�pX
*��m��o��X�5��(W=yPT��e����u܂�1��ڬ$�8)ɐ���Pt�j������v�D�8>n;��HE�.j��������Q	om��Qx������<��u�Bʁ�2�O�0g��ȜCwj�T(��}�xD����f�h�ܐ�t��_����H��Ҍ���D�^��4��R�n�������\���E��nLCd���:�]�sBN�LN�*�>�=�C��Z?���;)26�nI�l31F�tm���q�`�ڜ~P�F4 n���R0V���	7��L>ǃF��W���[�aիD�|u	����2x�	�������Eh.x��	��a�Ǻ�ksz�_��l�3��Ɩ���g{3W8���Y�ޭ�̧�^�u�W���,���ĭ����7K��ЗH~����&���~|�1�򡽃�F;̯��\78�~*���e�XF��q���_v�8��n
�t�������
ɬ��ؐ�$��v^�j����a�N�1�yeN
���ɑ�|Ey�8�d�_�Y�� ;�����IF��лF�GK&a�ٛR��5Έ�ۼE�R6Q_!W��(�)�t�Ŷ���Np[\��d����)�mi'}���L$*1���h�]apQqs2�Wd��ʥ(��������-�Pd�}2I��5a����t��z��U��fў�n�U�����b�O8S6fqx����e�k����_Zre���p����ATF�*ӊ�f�lH��|��$'>t]�/�7�Gܘ_����aQ�`�ߠo��P�ub������SϦ��O����[�6��>��T�z~��ܑ�Dn-+ ����e��Q��J��WfJ��@�8��+�-)���yZl���,?� mg�o��Zoפ!&�)��0hV�Bkl���aG#�p�e�����??oO�q��[%����XWR �P�d"Wp[gm���'�?N�-&�+��r^&�*�����ܩt����s=�8K,s�ǁ,T?E��2��A'�����e�X�."mk�jkl�,��Z�YD�y�<�"'��8����g�PA3�#r($::ۣb�S��2�R�(����W�0I�����\��F��Y�Պ���Ls@*�$�.�3a]J#� ���=����a��ד��;���A�pX��l�_���k�ثz�n��a#�y_�:��o�s�P�ش�e�Q�Ժ�"Q7�6�q|����>���3g�/��v�b���L�OJ�'�=dz+ib��gV��5-쩨�=*�H�M
y�*�~�[Ж0A��2i�^D�!��Ft�ť�d,ld#�U9X�8^i�&�9����!j��eϣ����w4�q+&T�ز<�a8��Lb5ţ��HC�%�����5�cT�>�/������d/8�Wq4�"�\:��JU$)�8�"��J�H �>�ʹDz������b��`3pyߚ�g�{�Dz�M""�H�����0�Z�K��b���ej�f��A5/3μZ��'�oHT�6������T���ͻu�p�K�z�=h�NosA%�
� ���	b�R	����3�W,б�I�U���6=$�J��6Ǖ�A��-�!�+w�i�u2��v���[ͻ���OԈ�y�7��'��"�x�:�Bc�'308Ry�v���Xg%T�7�ҟ1.�'�\�[��r�Am���N9ynAud��+�Jm�n�60���L��9�ڻDt����'��L��)@5Dܿ%�Ht�c����.xUI����r��y��yw��ҝjnq��!��T_j����sp%��2�]��[xu�T�wi��,�$� 'G}I�@>4�`=�t��Z)(�p9��;ۿ�wI�^�}e���/�m}V?:41��ڡ*!&��r,M"mC�7�C]���`�?�!�y�PR9�s�Nђ��,�5)A���%�!��3�@]�&�O���B�{c9�{ A�M���A���t�?���&p6����!����=�z��M����co��y��s�mԎhk�E�̃�?���d̢�Go���K��A����(��ω�3�ERr�$�L�Ƿ���BJ	-ԭډ1�R3�id�=����ݿh9�����O��2Bd+�!�p���:Vy�s�I�t��f��{���|��3�!ֵ {��;a���fZ&a��f9��m�<�U��k���O0�N�>��2=ƨ�t1T�P���z���M�B�.\lh��Y I/|�g$7�<�H��C&�=պ�C5^TRyMRlMZk�C���⻋oͯw��������L��,�jRd��h�1W�kWr��D%���M�4��"��f��,Z���!h^�s�T�+�L4m7J�{��%D�r ���IX���܂q�[�ep���Kz�9��n�*E�I��br��˿����&���tT�P�(�T��V
��!�ʐ�|�<O�m��Kph�Cu��2��_9��|�ڊ�^.n]�DC�sk2��DL.��}�����1�6B���9��e2�K�H�`�~�߃��౹��}ǛUZw��tM�iC�X?�v)�z1�^%7z7a%ut��
Z��n�o^9a	��u�����i5���(�!�ǿ��$J���I��ҍ��$بQ�G,�[�S0��F��R��j����~��=^�L�B���y���	Dg�3	�Э<���w�� �������a&�̲)��0�Ņt4�b�,V�ɑ
�Ǥ��fə9�FƩ��h.�tL7厦��/���R8�Y~4ϻ�B�j��-����<Gw�
�O��v�& OK����R��)���腷��E�����Ͽ$,�.ڃW�2����6���*���D�SΝ���>�<�ޅ�Gp^4(F?g������%���*x��y=F9�V��{��D�����@�vԺT� ���f�� ]�8,��v�-��1[%�r�IY�s����~8��&:#���S��h��,2�a)'��7��ZG0^����|���?�&�,��.��Rƛ���D�˵n�ӡ�����u `L���h��V���J!�n��9�lݘ���jQJ���Y��/4�����No�7K�+����	������s��
��c<";����8J������je�D�w��g�Ab ڱW$$1;��)��@�|C���rp C��등b�kJN��ss�u�����T���J���4��-s�����N�K����C<�=Ҍ�~zH��"�t��|�N�iV�}4>�U"<�`�����>7QD����Zh��y�P I�7�/7pk/�i��l:~:mK��J��<�0	z������g���_��x��4�hYF���n{�C#t�|�x��h�D*-A?�l��d�V0��v�z#����m��-��I��{��]f�	��_�a�ʃ �l`�����g�`���G�q_ri3.�T�ro��y�+Ke�;ڦ>��@�D�����^�5w�˥�^q�2��V�Y���t�P 6�$���p�]�N������iW���e���7p� PeN_�$�� d��?�
����VA�1� �,�=V� �^D-�ؑl��ԗ�:��ZRɬ���Z}2;���ܷ'0m��*~u���^�<P���~4�\B'�l�bTTl&u~�K��($lV�ުLt��I��ٷ��X��E{� �w�_�b�=صm5����2��ӓ���Z[a�$�J�ԚdNvA���**I��������Nd�Й�J�G�&=q�&�ڻ�+�t[����C&���!��k֬�7��{�4�丐�yn��%�{�4P�{1���)�uH���/����q�.�����㭭R���\��ZZ��VR��.�S#))��8:"����3�}��j�I�Dk*�a]������$�\���+|�y�((�1\#�|�K8�[�a�c�C�P��)������Qg&*��}���P*p4T	Xx��}��>�#m���x���>;�:��h/.���7$���f.���?ڳ��GO�zթ��}���Cp� |�C>���P��$Ý?�AWfӝ�~ߐ��ڠS��?N���zIWn����]�K��"�X,�DP�e���i��3a�z���&/h֮l{�O
`��@�4q`l��ǒ
�8%?|�S���=(��ci6�>v)�8�p�?�c�>�l���ep�yN8�_MK��cE3�0�������ĕ�F��]����}/S �-~�`�b��i����*SJ:�j�H$G���ig\��Z�8I�h�rtJ��Z�� EK�a�h��ȼ�g�|��v}ҩ�Fy�d��ȗ]ٹ���fx	6j��4S�!����/z$x�S1>����Ch�ԋ<�5���b��x��ǯ�핝V���c�w��̱_�������ӲMvF˻Ĩ��)�ƈ���m"��)�'h�y�l�X.8-ٸ�J���G~�<:G 4��_�v�'�Ɯd�c�ל��
D��zL��*{5�g�.��z��]�u���Z����PC-t�-���*����^F�4h�o�h�D��.�@�u��r��O]Iy`��&<��mw ,R�=�p��/$/�_��򉣠7[W�H[p}�&Y�L#�#}O/͗V1��\碞*�I�"X_��;����R����G���~A�$3�FD�r��t�@'�r�'��|���	�Ũ!�f�B�.�[Y���)cjmkt_0���0�0�U�]��@�4N�!N��^����	��"-;��͙ �J� ��a�>!�M{����{7�0E�zX�����7�G��S�9-�9<�u����-޾���k��_迅~�h���nǖ�#L�W�>��@о��۪�&�$$+�����q��#������W��g�_��
�Wٙa��'�����'�
2���`Se�m<΂o������9�=S)�Ҳ�ˁ?�6���`�)�`>�����'�y���b��M��K�A^�U��|{o��ݨ�ǟL�U�Ct2��O�03]��M
;�qN'E2Q> �QdPtIJ�ITL�{��7�������shp��!��I&�uO	���*�a#能�	'm,"อd�rը���N�8>���1!��	�l��������Wb��r��f��9�<�j��+2�M��'��|�'�Vɔ/��kw�
����##��W�~�w|NZ�Ü  �XXq�[�[m�x�
��o�1^3��~�)������^��=੅�i�̒����j�.�(�ޞ.�ܔR5���xM{x>j�\��]y���=�YD���E@O7�\7GLnk�h]��+hE��0�� ��\Jo}я�i� ��G���MpR/a�qC����1p���B�#�-�*�h�����4@`�zƾ���ޮߎV�'��=��e?�
K�`���Gw��\�ۜ"�0Yf�O���`�X-��2b+2Ő���প�Z��5ʬ�b��C����jnz�v4ͭms�ː������*Y��߱�����e�Z�TeFe�a Jݡ���uI��������Ń&r�(�j�����N0�s0v)�\�|��W�l��Se�$�Xq@4��0�H�}M��q���$I��^Kg�.���Cي�s���;�����5��(|^�yA�X����%`&O�����K#�>������Q+Fb5�S�@a��)>������K!pg6
�w��Þ�����ăl����6��F@�loG��+wġ�'I�9;K#G��������.U�����)�JM���C��Y0j��������]��ɹ�sf߉&����#	�����l�y��X&�]�a����+�0���\��	�ƎX�>UH{nj� �����,�b�_>���'L�I�15f�v�hE�� Ma����OE�א�gU>U�F� H�/{M�^5vƅg1k��wm<PI+��xc�}d�G�[ٖ��XG� �{�i������对��i��wďh����E=Wˊ�A��+C����;+E�軞 �h%�;�u;G���uRK��$�vA��O��/b�q�'#�'��u���.�氒~ςͫ@P�5�B����z-YĮT*�	���>I��>���(��F~��a�2HD�xuG�����.�iI����#����(�u9��?�6�d@7jk �O#;�!�Ac`�9oV�T�M<�����I���Oq�6�LC��Ŏ���X`�8� N�sn��wY�$Ք5	_�ľ�c��Q��VS~���p��4ǻ�!�G�[�U��6��H���a:��t]f����h<'hTS.c�_^�w:���� ;*C�m$� �g\��������}�R�zO������F����\w�����웓q��O�+�!��?��@�3�����;��fz"���Xx"�{�	�cG�>�8��-b�����<"��(m�1R`�oA��z�?�.�`�@��?%̕����ݗ0R�� 	���.r ��&�%V�:���g%���N��IA���Ưa�;Q�]���ڧ�9&�0�@��a�X5�J����-�O�o���D-#���b��\9��Do%&O%ٰ* |r񄁻�����J`$���uĆ*�Wk���0�*��KTdS�7No����S%dBW��Y!L(��r.wV�e��P���|6���x���W����@c�;+���$�ft	K!������1��LUV�p���E��J���R���S�]�� ?3K�#}�z�F~>Fo3�k/��5z���h���j����ǔ��Xj@f�צ�����l$�?a$�EZuKz�}%�e�S�+�ٚ@���0H������������"�z.!gG��~���j����I�^���{R��.f���ƞ��^������M�3玜e��VI�?,9IsJ�yKA����xȵ���#��u�����\I����!�;�?���`?��9���)��)�
�۽w��eO!3bNɄ���J������0�7��ot?�&835�3�*�u��c���~�tی�s����h�0N���0�9�OY�ϼ������U�J�p~��@2+`ّ\�V'Q����\�)�k�&�]�����}���t�v�ߌg;��/*�TR'ߧ��ċ#�P�B�NCF������ĸkt#y���u� w�o|�h�DdKu~����[��j]	��}�]^i���.f1.ǖ���*���%���T!�8v�Oȝ���F4�@j��z����H�:�==	,[�Ӣǀ1_T�Sd�2cD+S�]7�u�c1� �6� ���'|�E���	F@��s&�9���Wȶ �V����!��M�D�琌)��.}�?��pՆ\K\�2I��z~����Rѕ_u�gE�,%+y��v�G*˛�Q�s�U�������cg�#�=�?������H� �]���	�8��x����˔(� �<T����m���<D���k���,w/��}��m�{XJ\2�m@Nڲ����3�TɣK�R����ޮȬΧMjvj���8a��V�!�PC��n��L�t1co��t�?��@XŶ� �f�7�-+lh_e�D�i�>-\�C��A����<'���~�{_Ƀ��XV�]��я^%n \lL����i1�?�h1f�L��ŧ!�Uj�0�y�������w䲜Rk�gR��R*�O�N�
G�Wo�/�m�e]�꒽��� �+c�upW�Y�k��E������6j��.�� ��md�Ek��8����T�\��M�9�br9��B��!�x�Ʈ��8�5���=w���u{�Y����lU�OD6�e�E�i\��Tީ ]i+ʥ��՛uu�ЉUL	,�+�n%���Lv=�U��PEϼ���D�E|��2���>(��[���+��a�b�Z&��?KE=������-G�K�K�l��RE�'��U	L������h�rH�x�]��6]������N?F��[��vٿr���gl��>�مUx�)�
���1II3�_ .ח �W��cGf��)�4d��Yx�xdp!l�9�����G��/�f�#��e��it�����v�K*jt�01Y����F��8!�&� 9+��n��5k3���b�׈
G#�Y�Ǜ��G�ZVAik	�d����ͭ�<����"Dw� �m�6�mGʹ@���r�t��Jѽ5���42��Ij�f��~��(�����c�����Ġ�Q�ӫ4���ZZHf�zw���<�����Y�j����Éwx��,F:S���^G�x��YTA�JƸ01���or�S�A��V�������`#���7�L�ȭ��{�K�A��Aq�8��pU�Mz;��v&�D��/tm�y!I�E�hz����v�B�1o�
'�����ݾ���b�8�:�Q.���R��(!�r���(�����3�ǰ�Z8�����R�p\-�*g�OW�4�!�N+GVۀ�����(4� �/f'�>����JhI0n�1�k����pV2����ll�TiW�U9�m���\�_LHw�9�g���I-^S�<UR�ٓW]�^K�cNlgv�ηYȇ��_�ެ&Y^V��s�Iʰ���̣�����>�f�B@R_�U0���UO����_Pm/���=��ZA1�r]��7�)A�⬦�Ϥ@\��.�۵S5|�
������i�H�B�2�����,�ܖY��V���=�W�uB�8)#�$�� S*<
۰�nZ-T}�:GGx�8,.�� ����fA�!�e
G�?��u�k�6�R�աl�P��9�z��'mu��Yl5���]A��i����Gr>,�,�e��V�61^{o�
�'����B�!(�M�"��{��K}K��"7� �$�o���"J��.�.a~�>�O���,�:'��:h(��&�Gi��9M?!`�f'�c���j�=@aSɵr�#���$��1:r�"���Q���&��e�2�g���F=��5S���1��UU��r)G�g��SѰH%,�i��d�dI��ȧ��X�L�-!����5z`�bO� SG�_Hs����xJ��ݫ�:[�[a-�b�+�?_����Z9�0�����o(���'�Z}F3���^���xWke�$���Y;2+�["�/;;��wq��D�e�Q��5W�(�HJ[G���r�{O�wU�N�����L��s.��;�(�/�K�h�������/ЬV �q��Aδ]7�Vp:g!P:>�F?b�_�%�c'-@��w�~Ed�c��h�	��~���h0#`�z|z\t��$w���q�j��B^y1F4���
㘆g�?�4�B����ٰ�5�z�2ĪoH
�U����hҥ"� � �|5�7��1��� ��Pm�J�?�.�������^� aP���7z��p�X��'2���
;�qi����&C���YI�O����5�=��s����m�xĀf��5�)ƣ�kp�G6$���`�vz,�5s���og�Ϭ����y�����|zx�YP�b��=�����t�("�oe��C��<E9���s�v1���a��=�F��z	����B���pf��3P�w�h��)*r��3���_��S��|��_k�*z-T.A���%i]�¨<�@�Y����b����:9KԻ��l�"������<��}�8@pl�~�1��~F���f�&W{t�w�lhl=VK��]11�&����P��N�N�#�j��A�h�?���QR'�u��Ř��n٥�5#���,>������C=�Τ�Fs�G�Y[��t���g�z��k����,6��W��O�I�؇�߼���l"9�솊K�/��hO���%NƼnrfL#N����۷*	�c���[���X���>���h�`��Z�*���?�K�H���j�Jע��
���r��
�x���Iꡃn�yWA@���J#6u"�+X�y�%�$=��b諭g&s8��ɫ�ET#�0e��.�;���5P���o�@Mß�7��1�H�9����@�K9}~�N�����J���B�_;��L+�d�Ly���_��;דG���~iV�e��oN���A�o��
�2���A�G���`�+�LcW5�� �IU03���>%t�o_)�E7��h1wj����K�`B��/ �O�^�C�	%�2�:K+V���gmub]`If�ӗ��8�����'e�߭�������ñ��95$q�}&��-���Y�$р��)�2� ������V���_Y���8��9܎�/Ӎ;��(J�z&�E�w(3��`wZ�T��(�ѓ4-�)6bŲ�}E*�� ����Tt2��j%��R�+3g�����1�e�l��X��Qx�I�(88z���3�-#��ڈ��I#O�b뽬;<-�7���3E��de�R�sPӶ�fAP��C6d},w6����
������6"��٘�>B���r�6��|2ԗ�*i�7g�g�;��9#N�fi4����1m�'���RG i�]�\%�g?!�Y�)C
����l=��^��~�!���.%�!=A�}�Q<o��xOn�=�ƶw�SX�\UB�%RW��l�7�����6N��U� '#��6B�@�����&��ZV�J���S���>�˗9�����ƪ9F�[#�`YbfXO���s'�ɭ~�,&��'�`v���w|�Ĳ=8�f�d	9����mE��(c�3e�S�N/�4�F�������}�5�I%�o�8c	 �Mґ(�T���hm�C��y����.��P���m[�#�����b���?���B��I��C	Ƨ��ͦ3��54�~���>	��'�^��~��D�����y#�u
��,E �,-0��o����iۍ(�8�C���늼�^�L���4��j@-}:CnfM�U@��O�#$|`�Uaa�ٸ<+�Hy�W�"t�,��X�Oh��`���H���Z��gjCw��VY�A߶��nv�1j���ʁ*D~-V�	��<�Y�*��&һ\�����X�7N��bݿ�0iaB4[F�s����9�ά�ጽ�2c����g�ڵeY��ڪ���j�<���¥�nCY�i���S���8�0FRQ��.j�UGQ���Ц�wb�-?Hߖ����PAH��7RS���9�9�Rz�mȝ�b&4LXpl��1��,����0��	R���B��*��1��ǅ�|Kй�T���Q�������28�.���Ԓ��^%�Cb ��/����\�5�PH2���LMܹ =-!LkbOXe]��v�*|?^�7����B0��i��\�:b�%�/!����}L#U�<nPaóe�i 7�|�&�k�Yo������r�Ņ)k�NĲc\K�s5z:-�zC�[�&,���x ���y�x��;��p�^�{�?md�t<G��㓌�	�=;�y <��l4z���s�W�R�Bt�Q��'���a� j�ڻ�N#G`�(M�����!���o;?�&�]^h����E��"vK(G8��'I�L(pռ��b�$Q�󗿆ՊS���~]9>`�f�:�k��V#��H�3�h
0}O��$��﨣ۨ�9D'ϯ��BS̵�[pԟ S�^�>t;H���'F�b
��k�O ˄����`~�?lM��G�W!�α�5����!�1�h0�m)��<�RY�T�� ����+�26�������ya6��!�	��Z�l_���ӆ �!d�����ii�A+�0�-��~p�y�.n��P�\�`5��$>��r1H�6IT&��-��Y�:/�!7�5t�͟T��["�=�	I#���Z�*֧�ş��+� ��0舤|ԑ}c~(�E�D���98T�tw�߂�f��)� ���6H�u}=_V�G֒�P��� �D${�����U�K؅��t3xӇeZ�^�x.���)��'	�Z����0H�Z!$9�����Z��X�������D]V�}�ġ�2Âè#�f�!(-�&w�踖:���u�+[%J95�����T�ud/����Ze.�F����Aڬ����������uF~��,@�x�z���
_�h�]��oxرM�g�X�g{�l��_�q�T��L�c�.k#uɣ�<�����v�#�p̤�OC9pŇ�Q��t��d[6(Կ��B4������tk��!�X�bd�A��Q��ҳċ����?���SP�3���f�o�w�>�PW.�([fci|c����$����}�>��H>�L��T0D�˔��H�{Rq]0�9Zd��{'G��S�&�	+Bxo�1C'�U�R��9��F�u�8P2U�I��-*�ǰ�����U�|��t�f	��֐%��i��+aj��y��.�m6�~%��W�)���=��=N'�%
K)fjK5]us��IYM�[ۥ-�QY���3�`\Wd�Ÿ�,��mQd]��ﺮ*b���y�B��;�d�p`�x%خ��P���:�r��l5��D����8zzN���9{[@BJ�4��"����;��L�
����� I��'�bՔ[�T�S��D �+�l,�&ڢ��Y�h�0��2�z��Y�Q{�R4
HYAj���vB�DG>�܌B��b��K��ʺ����ln_���z�9SC�s��ե�ȠCX+�2@Qi�Yt}��Q�T-a��q�I��]_K��BVO�a�*���/�U��.de@�/�1O,t�	i<���D�?#�":�D�*����Ǟ}������P�e�@s�AU3�WI�)7@3��t�����W�4�s�ͫ�yj�K�,���&�0Rö��~-�N��P��t5���R��
�"�F1��m�8d\WS�F�� |--���I ��HZo�I"j%�>"�O�<����������o��#�\S%U�� <�J�?��	k<p$@dB�V��7����`�v�0�}R\l�bJu4>����{���9|�]JezZ��qj0F�P3���Q����-9˂ĩ^U�D��QУ��E�ܒk=�p�&K��n7���L�脛�<V�s�p��A���G�Z�
��-�s{U%�OTy=K�t����"O�%A�>M� �NC���������֧ݖ�َ�5�x��0`h�d*ǈdcy�"�C�]>�¢�,��yhJ@g6	�.+�{�Lv�H�����nk�څu_�5l":�cl�_iġ؄��,��h�Ey�z :�X�Ε4� �������c5�|3��^�yh�5��I
����#֯�M����:�ӥ��$�r��? G+#���pZ���a�k��ƂI�x ��K�)���֙�RV$Nc�^
���e�F���=��-|�}�Q�+��)R�����_n��(�fI�055�-�cl*"���=q�X]�}��8�c{Ԙ��6i�k���I*e.V�%�d�x�Q��	�y�)��>Bn^7%�f�ݰ6�4��5Aʀnؾ���w�[�F�hn����������g�������6��]�>�&,��_w1�xل��<?ϓ1�J����.�n<�,��Q������4�hp�̠��Q��Տ�ZX��w��kH%ti].c/��:���K{�etWF<	�k1}�q[���� c+��8F2SU�����3�V�Sџ:��V�B¨ھn�����se8�I�1U'8.j����w�#�	�A��I�sw�LL;��1~���bSm^���g�������Я�;�M`k�&��)�O��AFДY?��r���|�E�����{�l��7~��0�-u�9�wޥu�h���Z6�O"V�s1硾��L�6d����U�J�Ct���_^��`��<�8��4���D:���2J��\8�-�u��yV��,�m�n�dN�Z�-�E�u&>��ɯ��)��c�+F�f3+!�tzj�8�d�d3s�[��PxU2��$ ��룦P�.�|#�� ���	Q*rA����� ѤVX,僷"m�d�s��o�V�'/�K�ڃ{�J2;[�)�K�����=��,a�%l!	�ͩ5��D�Sl$ۮ]Z���!��Mc���������p�sj�w��eܳ�������j2xd�1�1��y�bVpR�;��s�(�D�6ă����P��$R�$�-?L������٩2 ��I�ZP��P5yX��{������OU��!���v,���x�y�!���k}�[�&��8n�1 )&Ϡ{D��ކkp��d�eߔ8ZVr]�B�FG0ͩ:�Z�:���������.�h;i�m�3�
����0�N���M�3�#o��5H���"e���$GE���pb�N�ly�4�M��ͭ�\����k	�D6]��,�t!�G�=��nJշ�nw[�"mP�ҤY�ML\�������H��f��=����=4P������=�eD*h�,�E��m��������a�s�Ct%����γ��g�"�ӄVc:6a2�j
�<l�.��AYӜ�=��e�X�8.jH���:-�6����hJxi9������d!����,��jmgs���P�����\9h���Sk�������m3C�&���:
�r���-��V�5��0:�����vc}�������:�r��4)*ʒ��{6c�cz�Ų-̟�9����7��z�
Q>7Th��oۗW����Г_�٤*���[	86(�ڻg�"+��L~�GE~�+'��Te ���'�+�;�����d���f��pu���}:W�7���b�0>v(�����_O�@	�<D�����d�8]5���Wo,.�x�ќ<Tiϑ��]v���S3"ئ������7\���l8#�FJC���� �؎gN�Ծ�J���#"�^e���b�L�+{(v�����u�%��O@��C���/�]��Uĳ3H�U��׸�0�O�}`�1���:ӿ�y����� L�1���w�=,�Z����`��%a���v�`z�\b��6����%.ƹ��rȨؓy@�-������ͿBN��)�$�I���x5��M���v���)����օ�ɒ��τMʂ_wq��͆�I�	�r�$uk=�r�մU<�%��4}�je�?�����(���u��^�WN䭟(�D:NIv�3d�X��������ZL	йU�P�Y7�F�)��Ӿ�W���(��`����A�2�x#��W�N���RVfi5�Xw�6��b���j>��Sg+��3��u�zA����11Zcm1���K�����K�\@Bd���n��-��-���ד�����ˬL.�+}+c�j}n<�k&z��~
���8d7K.�������� �ʯ�Yǰ��(?(�~����|��X�:w��I�	H2��~�_���Npޛ�{�u�espF+���H�ֆ`���.LO W�fz.���T��i��#:�8�K�)��LQ� F�oM�Z�dЦ��9b/�+m�=Ф��;a�G�����҃y<����n�Ҙ��B���5$�}A���PF�L)iƉ"4����i>HQ�]�T�Ya����Sh�gj�V���_�K��4ћtT5	������˂�7��Z�α��?��a$S�ҵ|eQ������.6|�M��IL+�q��E�ĉf9�*�0��J/+#�c��d�� ��-�5�"�!�eR,L��k�3���3P�u3~Z��6�=��^��ւ}H5�m3b�b�#1�R�o�}p�U_��g�=�x(�1֦����v��BS����EF�}3��� ���Ǆ{N4�wu�(��W�r���.��	T:��ݳp�Tm*���F���f�� 2���o��m�&�y)'�)����_w�'�b|��STn����`n
	��[]mtD�Kp�j���50yFD̔���u�4�$^~j�o�:�m������� 5�l+�R/Ϻ�v$+o��K�W��~�-eF�����cʂYT�M�XG~X`����*��v9��a����O��/2�xR�A���ٞ�)���l%���yQN�7�Q^��r%S
�٢��������I�˴qq)+-�����!BΣO��"D��2ߜV�
d{�m���|0��n�a�]`�I3┬?�=ů=~mB3����&��7C0�R�P�ß�wknzm015�^X�_�帝�3��h���JNS��^���u�ǟ.��i�S�����CX�z��˗X�H��ej�:�A�ɛ����E��?���oy$�O�,�"��*��:�xU[_�=G1=��ɶ@���m'mh��)�/9lr��I}ł��͋�.����A�:����=h槶r1�k�L2[���<�p���¾��Y�A��pa;H�u��'��>/1�"��cG��LG�l�f,p�&�U?����dѫ23i�S_�L��뎈�5�Ц�l�c���ҷ�LO���`��xH�3qg|�C�(�+�G�ɐ�u>k{�
q���5�Fѥ��� ��������ֹ"��q�z�"�ʗR�Rܸb/�C@R,e�]��xD�U'B�^-}�l���=D�!�H���	�d�yו��],T���Z�s�o� �׉�� ���,�/��������BI6���u��d˶�yܧ����1��V��S�N�KJ2W�)ȍ��GQ"����V)�8���G��D����z�����lVHE:�c�<���7���q��ȶ�r\�{�n%\
x��8Z�I$f��K1Gb���(,�_��O��v����*s��o2M��VX���B��kx��<���#&<K:�K`2�?���glXu��cA[�%Sݯ�[k��V'�Yo	���ݼj��w?�>R�8#���&)��R�./5��(��i�"��$�!��6��P������6]TY j�N"���Eۤ�wdMwE���Ԇ�Ln:[��V����f�$�\OT�WA:���ng�S��k��UQ��v�o���kj>&�)�4�Y����`�]�I��°Ϳ�g�t)���]Y��$TC7��[cpV�u�)mv\b���%�m��h�4��3�\ӡ�lhO�N�dI^�Щ��܈bA�PG��L��J̓B��8�9�J��L��8*:��LA�/�Y~� Y�k�ĀVR���b� �7R2���m.�E�Myo=���a�]�|��u&�7K�`[���Ō�t1pzx����+wsq�h�B�Z�:�Y�^	kT��*�a����g���F��i��F;�%g�������P�l�Mh^N�K�}�LI�k��j���V/� �B4ڐ�=���!
H����Jg.�a/�=�����BB4���'#U�UJV�7��,�!ř�D����@2����X�Е�w,��f7T�/�[-��V[K���5Gq���([̖��$�Ὼd��1L0���QE�����ĴS!0B�)�!ߘ�'DI���Fa�}X�S�4T�qű�4�E%KOf�#O���Qr�b)�2��^�[.�8�$���]�'��n�S�S���T\(��2��@`�(��}~F�&�ɸ�hp����Ȭ�8@c����oe����l'GY�T���y�@��TY��%rQ���(g[dH�\��k� ��v�86���Q�3���ef"�4~�2��F
�"#�)�g���������-M:�s�+U]�|T���6��� ��I�U�
}�޴g�U^0l�.B�ue'�?xڄ�`�	��0u�����h^q���9�e[���$'�HR��'W���\����0�oߖE�r�LN
����κT�?
rş֌)�3�yo�}ʻ�A)������cf��#h�$jԛ��;l�@̭�S?o[k�9��B��1�������5'� ��2�U��߆,�i!e&Y�13ǒ�R��J��)�]�c�by�i��qV���׽�������?-�§�E�*�/7����wk\U++]L]HH�ɻ�|ۼ�pk��Y�y)w�6|����
4�z	mb��#果���ړ�u'j�@-�=?������A���1�p%�Iu�;����������o���G�G��p����\�m����
	+v�r�&�:a/��<����~4b�	�J�$���Z����R��iD^������DF�M��}��d�Jz��ˏ���࡞��Hq�Tid,���V�SRl���Jj2N<��Xwl :�!l�dT�\��9NɊ�#)]���QN�^G�b�]���vۺsG�ZYa�ܹ���LGlgu��Z�,�q^�r/���6P��5�*�YM}��"zTt���f�c�!^���f�����S4f^Y݌���o���es�	��ױ� ����v�`�z�|7�����G�`Q��\�P��c���~����h.�k��֡�r&`o����}�� %'bO���Fq+^�T,�r��I���t�ML]v7�@�F��r6@yA,�]F��w�Z������E�;���\ y�{Vt�߰�6c��n�;�-�!SXQ����É'��-�;���l������
:���z>��%�˴J{	-HI�9K���>4������w�eVm$�z�
�&NE���ZreE&��CZ�̵����R9t��Zjc�ؑ����QS�C��@j�¥3��ϯm�Ӎ!G�@���5;�o�-���ri��l��1�E��N6����A�F3d	~��T(��3i��r7W�:u���ɏpc�z���T�ݣ��xxx��N��\y-�h ~/�k���R�3'g�ݱ��nHt�0,2���E>��s��3�M��LةN~5p�qU�$��Kn=b�8��nt�̲T�>��^薆���w2��p;���Hdu�<f��z?�8��x-$���9�WUoL�}�%ҤD����y( g��P�+z�jJm�%!�ڕ8�����c����Hb4֯�,؆^�[Z{�f]�{em`8��H1�
޾��EL�8�d�^��jS�ބ]!���O�NQ��͎پ� �@�k��.{{!(��%�@�O����:ذ�ҟ[�McK�w��N\�T�(�uK�=QĬ�oU���1�Wʣ���5��kD�$��L}�C��I{�z��=P��]�Agͅi��PȮm*��y�w�s�&�
��)�髣���3l�qI؇���}Nf��B�т�N�&{WICB����S��� �^r��htK�k5��h�6n�s�%���ߒ}O<�Vch�M�7�M�%������$w���iͥ��O����J���鵮��n�����BQi<L�����2�yn�y����|��Wo"d�)�K��z�v
���	-T��^�oxtK�,�%�S����{��l0}l���ri��M#'��|k<t��wau���n���ƨ�����������㓋��5��9aq�z��_����"���Wk�#��$���n@���F ��؛�
�L�]��q�.S���B�H�{q��;}e"��b�~����xh����C���痘�֛²�a���!�f�_1#�S������;�Q����t�璗�1B�=���^�@E�CG�*B���v��w1���n
�W��lC0?��.�����Y�#łQ`e�)W��6�B�?�42��ZY��5&��v�wbO��ע�I!�2C�MR� �Y�sa�k�
�ҏ❶�;S���ǒ�TOir��*���&0pg!�\�v�P����a O�OJ�ޜz�ƃ�M����G�g�\�h2��/E(�!�{�/R�g��P�� ��MGG��
B)1O�`����έ�$Jr��b�ǇY���u*%���h���~��"�������iط6J@��q�#�'a'��[
 �~�4P��p�$�7!����Y�[��XdvvId�U"G5�q:���l@Ȅ >jt7��ꓕ�;��W�/4�W�/�d^��Qa��{J*4>��7�o_���O�����@)�+�c(O������R���=2��?|C�Ө!���֟e�ݝ��f�_=p�qc@��N��+fl~}WU���}uu��s�Yv�c^7�U���C}$%���t����׬X��X���ܳ�:,3g-,Ŭ�N5�8������v���������1�b\a��P�,��e��'��^`��Y�i4��g)��	F5�n���ލ#��X{3l��@�8t����5���K_H�^Ј�ZS���~�����|:r��Ks�dK��ȁ��A!�9���S��ث|���hXC	@�Q"I{�U����{��gN�q{�`�3��}#i�>�H���4�����b��� k|aT�����n��9��<v�`�I��X�(C9�EgY��U��tE����$�7���M��P��^s)�V_�.2&k����D�~�:�Ȥ�};Y�D�%}d2��k��~G�\$�Ġy458��{
r�rg�w� ���|�/Yr1`� Sn\�fA:w�!�o�FR�o��D���og����a\�J��՜m�Vr@��ńFGj�e�f�يp;��?*jG�(D��P�fѬ��a�u�R	<�z�3����Z�8K�a�=l���e���d���
�i���&��0� �}Ӊ�N��&�M-��9�ȎW(L�c�:��8|�(�}j��q�w�_��ݵ��`+1N�L�9��%w8���X8tCJ�b0xl1��U�a�!ⶄ J�|k>�� lī&�w~�J�?6릿$g� ��r͉�FL���%|��F�r2��N!P<ֻ�m(�N�ڐ8]ɟu<yl|�
zl������x��������;����A�b&�� x�݋v�O\$�V��@���.�����l�z5�e��p�G<�\���S�IC5���R�=X3�3��U����?\�7㌆S���Z�i+��1i�����+�"<�/��E&��߇.�k�XS��H�Q���u�])�_�>b�����i�?���}Y���(���'���bea 7�r�g֛>����#�S2S�FP���e��2�.pTHp�T���(�qm�Ũ��%迱D�n�̹%�>
�z#�Yi~�é���`I˷��� c��F�Ɔξ�׮�~X�JQ��{��;�z����_��%
�WM��m����
ٴ�[6l�rI�*�N�.7��	���-��{=��Q�ӱ{@:�QZ��8��	��X�|�9y	��٤��O�0���MY�1z�5��e787�q
�Zz-�c�����g��E����:���Z�Gg���_na���G]K��G�~$ey?iuo(�7����b�2ė�[��&��7Lч��<�i���΀�*��'v0]��=�4��G�в��@Z��Y7G�4�[x�Z ���6Y�u�f�q�?�H���f�{;dJ��~؎f1��_���t��	mn�pω�/h�a�6�^W��yX��y΍~�T�C���F�7`꺠�w[	1�.NeeY[/��f��?�{��ֈ���_��R7�^;��]�I�>*�o�~vv7Y���!|��`U���r
��[����}"apS�n��)Y�*.P�hK3e���`�.E�m�aiјD�7*����Q0�]�m��$�HkjN<.��e]P�u�`A�b��*��2_0)��޻�����f��+��:���t� �G��ʆ�����w&K�:7AAbv}����x9u���`�,�ɻ�`c�F���	�_4�'���p����#.�)�#|�����j���5�.�x����/-���r������z񍚇6���<����M�%;����	��z�nc�lXU�O�/u玛.jA�8^���T:V�g�q�q7knF&r1�dD_y����Y3���ֲ�e�<٧�wI��;x�w��0�8�e���9,�� ԧ]2��L���b���(w�U�/ު��B���8ܷgK O�D��O��<N/(�D�d��F��t�u�yh ���)����^�{���gL�pyx!JT�T���tcHv�9]�!��3���������v��� k���k2������O��a����̺�$17O%S��p�?o��+�y�<gunK�c3 3O��<��x�b�U:d}nJ�|��C���{-t��V~��53��;�h��4\2H����T�i?b.��tb�J~��P]���S��u9��kNQ:r���6� �.T#nE��-*{����h69����*M~u��5�����[����ҁ�d�n��ܬ�Ys��L���-SF����֕�Y06�Hp6mڂ��>$	He��Y�;���?g���*X��r����H�)�(���8�x,xGG��	\[LG��^5Z[�����*0!���D�;�Q�M�
�?��9-�~wNPg���ه~��}i��.J�颀@��$}"#H�!�$ŅM:�D2�T=�]�)7��e�s�t{U4�T�g��C"��c�ɚJS���y�d�s��Ң\XsC�s��	Z�
Y�� #å׍}G���� +��N���(&(U}��ޠ�v��/a/?&Zː�Q�x��s��[�|\A���v\�{��n�/��~��v5@O��Y�.��C���\�A~���IWh�B;�7ٜVq.?�vC��[X!������c116c��q?�7��%H�T~�W�=I��_���寪0�z@���v���Ju��=e������I�[D�v�\�T�O�'�B����&����p�{�ŲP���
]�4ѭ4ȅ\��~�$g3�"�6�X_�����K��ʯC$����Y167��>��_�CA��$4@��(C�p�K0��9L�`��]����?����E�L��zd��١Rt���o/$4�Hy�-�z����	����%�=��9����ZP��=����EY����竿��%dm�>��R`y�w��[k�^<���@+�W�2b�C-�F�Q]ٚ^#ʕ���&�5��=gh��$��D�Fhu��DoGI*<GX7�yp%��ķ�Фפ;sl��:x ��J����F^E�z�m|GH��t����?����$�CX�C��B�#��f!������"���e�����"��%U��;��D��L糗��ft��7�׋�7r���[��r��癦6	+x�0��c�`Æ��+_���x��QV���Y/Fާ�V�?LP/|�'`�7O�[����xayU��p���Ҭ�⮤�}F�Xƪ�p���8.���~�`��H.��J��H��Jѐڃ�\��M��P�,����~�v?��x&�,Bc��>)\6y��ʬ��-��F'*�Ʌ��W_[a2R��R�V��[ˉ�U��\D^�<*lW;�T�:}+Q<(�y6���NG���6��v�m�k���kj�P������D��-���Pv��^J�zn���r[�z+X=Ժ�"�~y^�N>��K;PQyg�X�H�#��a�I�.*�H�w����g7p�Sx�n=4�ӽ>����>�^�Gz/_�	�#�����e�ڈ��P���n�Q��̄<�������I�Bm��H|��_T�D����#�/������&�"��P����9|��^;!����y+P��e���WQ���^�s;Zc
L��}÷xx�'��Х�0�i�>�[��L��~��x�9 �#fy��P�
CF�ةk�)f �M�M"��.\҄�~�Sa[��$�����8�&�JM����hL��t�ts�}�]`ʮ���o�VQ�X����M���|�l�:��>"��3M�9�#�1g���k�����)�F��:�姮Q���6�ژ8����6���+U��:�~9dؒ�BvJ������<�T�ɝV7��3{L��K�C�©;{˲F���a��
��D$Ҿ􆍨��9�8��PG=��~~;�t̢XP�+���<�vƳE��Y�4�����?���&�2{���1Xgp�ݨO�2A��V&!b�����rt�lV���^��$����5q~��>�*D^�o�R�c�(�׾:B��O j_��)8���Pw���4����P@m;���_�d9���?���.$���m���Q��*^1�Ɨ
��Z*UM\K�������B������V��3 sᶄ��t{E�^5�`v|N��������d��7�}�G������1���C��/O�k_�{���d�4��[��v����}�G�4'��
!h�ײs7��
�ŨB���𨰎^�����C�c��a;�����X 4	��H�g)��%Y�՜`��$��|T_uL�K�β8Pn�Et0�2b
E����Cs���������j��\Ğ�qS&��پ �Ӗ���Out&{t@�/����i�����*Z�����n]C���&�c<�2<��!Sfy�����4�4���;��qp�����|��-��9��Q�4�F+!h@��ە�C������D K�
� d.D������I}H�7����iʬ;9�`[�R<'��a�z�DǧrTxHsєQ%w�fB���\�Gp���dg�ɐWm1G�̲ߟ}໑����E��=��^��A�5�ܶ_�Y�a�1�.��ծ�C� /�eUY��A��&Y9�`2�j�z�k��_��<�ُOΒ�Q���:���{C���{��W�TM�n�*��|ț��W,���M�n+3 ��ȼ�ֹ5�l�����i�����0[�޼����	�g\>��/�R��(Y=��1�H5rэ(�>ӗ	�6a�}d=�T�r���-�p�#Z�َ� �
)��]v��GE?J�VpJ�IBⱢ��7:ϔ,�*��{�u��;q��_웢2�0�DFH�A�4G�
����d=�,&s�g��΀�|�c��ޔ�Ba�z����I~���?,�|���X���UV��K�l�����
�v-��;����d�@�+>�����DMۊ,��T�+Z�>�6�צ�+ުR���>�X�6)��CiB����û�R���O��-� ��W�x���3������!����&����*���)��%�{Gu�+�����ߛ�M�+X���דe��0��(Y4s��ӴM�3OR���jD�r))��x�',Ay6V68�����m���B=s�,��6#���%E��"�YM��k���:��<�ۊ�J�űg3�~�4�l?r���[�����9+��gx2F&9!�zq���W� l�=�Q�@�`�{���csɺ���O�^�����	!���\�M�$pK	W�`���ׯ�U��)�cjJD{	�N=��:��Y���!��^(u�-�ý�]%#i?�V%w2'N�%-�fS�n��/���ߵA�����\���ƿ�Z3�?+$Y�T�'6~!�.w�#�GIڎ�{��-�'<�>]Q�+�4��,1U�^�^;@���FZ?��<�\�5�?�;c�PZ�Ȭ&��ˏ��b�Tw]W	�2@��(�%�R#	.�tUK0`.Z��\�BT��`�a5�By��q|���Ԁ�{n��d�u��e�tq�Y�����[�G4	��ǋWy.4nF��y�fF��k�<�z˦��Q#c�ul����Ē�ֹ��A��s}�ɂJ`톂�G���� S,'3O�
K��&���8�:c�	��Ľ��5L%{�Ҽ{���])��#���h���g�ٴA��ê�f��6S����K�ʉ�̩�om�7D� � غ�R���-���L��|oػ{n�����\,�5��Tm�A����v���0����)����@�M�@�>\���.��d�N$�%�]7��).ng��r�b����i| ��~?њ�}Y=Y|q�8��/�C?�RZX�a��4�xE���tc��Ȟ��Q@$|��	�	BL���B�)�|5�R)�x�3B9r~�&5	�R�lw:�Z&em�mh䀦e
o��������,�2TA�i�%��ԭn�ds��;~��h���
�G���%(T�v�z���f2�qV���VP����-$��k��%���S0�>=�2��؄mz�|pb�����b[����|Y��Jw�O����kew�d��?�������A���^�*����S`w�H1��a������DeI 3 �㛩;��(�}$$�Q(�C{G	H�sݻ�&&�R���k̴R��@AЌ�\n�R���ˌ��.t� ��iי�Y���
�I�P��G]���OB*��5�k��ߺ�O�E�>�Љ����U��%q���r	�h���p*-�o�N!��S��v�,��{߯�4ނ�~�H�w�m�zf�ӈ���~`qtݎ����R���
e��,u3������P@�$��zk.��^�GCW�z%��\���w������v�}a�DH��|:����*�=��ν�X�B��v�V��F��Y��z�;�$�>pf��:B�I����I)���/t�9��|E�/\��K�Se5�۝G�[���#價�������i4��,ޛ:���u9��
�@bW�,��|]�Y}�c������I�#�E�>t	k܍I1'�0�b�TpK��1$�&sO�P��{I�����,��/_و���"�L�����ۑ�/������-	OG���(��љ��5�I�Vͧ�����8>��+�)�%H�l�S]��{��j1�m��$Z��:��&s�/��S��1z�s�bR�o/ -M���@-�Y �� �'s��@�N�+G�x��'�*�����S}
r���3���T�|׶Թ��Y�4�^�YK��/˶%�T�u�	���uо�Ho�I��܁�܋�����y���b�R[�٧��u�	N·F%�a������x�~�C2T=L2�$�h��mr�m�2�q&:	�M�!���J&�SmҀܢ��`��O�܃ouN�dڶ��ii�}?���=J�!���8�՚����$��l��Qq���>�1�#��A�nB���K���ڷ�#��0��Sj�*6�zaoO�:;~���H���X��rZ�4�2\�e�Y:����0l������<�	(_pp*�j4T��'��R󽞐}��Mކ�_*���E�&��RH���x�H�,Tӣ�{���dm	٦#�F�.vq��h
�r�PiJ�ӏ>��y���8G=���u�щ�e�^�aK4-����P�xg�����2���KƉ��w����>��C��@���T����<�l\Y��O�c��`x�Sq=�)��Nm�S�)uٴN�TB�):`�h��yEYS4�
�����j#e�FP�躠�̿i��N�ь�{�A����S�}(t4�#[j��*#{)���zВ}��A/�r�D{�=�͑6�~�b]ϴ���%zMӪ%��V@l���޷�'R�G�@LG��ؙ
�d�,:�E�;�����������,��� ��BG
�8�j]��E[��F�&���2&�02t%NaA���^m����-�,!k�K):��B����]x�aRw�����Z\�K����pJ%j̛Z���Jr��c<��r}�S�#�Q4bI�4K���a���8�n�-��X5䰍��نX�$,��1�\ByG�^�=xgǓ~��Y|�E�I�M�.&RV)k���<�x���'���]� F�����9ڛĆO
��mS)q�&_�]~ 2���Zc%���2���7��QVE��]$�����oN�Q�$��_���w���9�OJ��L�ZR�ո��)o<���0d�̳ ���{|���υ�zh4H��U�(5+6s.�>��T�
�K����j��˝���zܪ�<���Ə�J+���@<{�/�Tnb��bGg.0�q�PD���:4��4�,h�Zǀ�9��\6��@���B�t(c��@CH�5gp����R@��I��2�����+��w�#������?�g�A=��P�(𙼢/�l��K���1kn�~GU�=�>�Ma!��Z�&(Tc�����'N%����W��Qa�s��\v3Cν�҄��� �y }�kP�����}7����������;ە��oQ_ti��zSW�{lヰ5�6TЖG#���'�f}D��|.{�Ԛɷ��u��2^J�W  m��&�SF4�Пo� �r����������E2(JlB<���t�t������hAI��]��fq\��0D2�'N\r�C@�C(�`���Xx��ϟ5������3՜&�������Pe���٢��0��Y���O�3�JFy�-��y�:�3��[��M�Jt�Qf,�(���؋��Ǜ��Q}J��$'��KBf�d�G"��Џ��/j*Ɣ�͊�;�#��>���e
odn����57I���5E���W^�(��:9��JsN�Ľ�m�?C���\�QD>���ͣ[��fخ�7��~�7®�n8B7��>�g�%a��&)��s|�-$��$�掠&��*��u���'�h����ͧN�!�  \<V#�/������ Gv��TT�h�N|'�/Qg�D%�ca)�אT�aΐ�����B��:�7��<��ّ��!ۉZ]:�噛�
���0N���fe_�!�f�������P3��}���Hؙ��>��/�Z��hU{�q��楃�8y:-gQk9��B����w�����-m��S�ŵ�+�%G��id��� �9$ié	6N�L�q`����pF��H��%����&�Psx{��}�l��a���G�$(�F�TJ�`��ZC���W0��OpQ_NI�y��7�놕oˬen���?=^n�����Py����x�"�C���:����H��pd�9����ׂP4t8�� ?|��u�N*�A�_�E���+��Z�=J����W�-�Ve&݁��I�6����@R�q�AJ�J�	��-�ʢU�
�#<��XM% ������[À�]ݮ7f>Ke!<�/E(�k��6�m `j��2L���Ԩ�,�1Hj)��oU�����g�wΉd�4�_>��G�H����w�q�J��ǣ�R����Ō�'B]�4�Ƚ�۠��A�K�3�M�7�"���kMlX)�E�E@�ѣ�h�>�Oj~�o�*�W�|��7�e�JW�w3άaL�xͦ�69^��"�n�ɹ���,	��]�99�}�h`g&<�ײ��~/*�d��a��~h��7 Y�dQ�T9�y����J���E9�����lTE>6W���,䰑��c/oh�`�[�ͻ0%>�&��{��R��׷�N��F�sL'�g�7=�\>�ϡ�,��Y��#��6��m��F�&m��~��[��TK�&#�zZ15��6x�OZ�FC�.J�*�녮$�	L���<W�`A�hd����DVyH�/4�
�jK_y7L}�1��k^��Y?�@�gm�:��������Xzr��X&ݸi+��A�ch����O�¥�T2>���0�j��&�(^u���O�Rܿt6r+����'Vy
^�=�O��0���e�(���sGb��0h;5�Unɂ��R�����'H��!�J�xi�}_�����d�C*O�-�%ðK�Y��<Hږŋ?��G��n��|����=��gP�'̗E05͏M'��_"j\��D"�g���� ��=5�g��
UQN��oR�lP&�e�,� (�aa�r�Z���G2�1^��s��G[b��fD&>s��t��ͼ}����Pu������ةV�P>FЍZ]�L�sj�j.6�v��娖O�w�=��Tv����3��i�O~�Aن�C��!q�\��j�.�7������u�b>��%��D��cNv��ʓMz,�Q����_�&�G�E6m�Z��.x��P63ˇ����+�^,[�?�E'�� E�d�z�|E��Gέ�L�O��Ŋ�o)+�8��ؤ���]�O��C�`p�gw3�9��!|�H�e(��V�/�	�u!HS���9P�i_�	0���2#dLn��D��R���u#���!�8P�li�o^�"�l�O������K��ܐ��AN1zȏH�9T��("p9+���X�s�j��HW������r�T�d��5�����|7Td�չ�`b;�:>@{φ���� �4?�u	/���%�����Oo�%g�?��~<���t����1v��p_��j��J@��|���V�W{z#'��uhD�Y���Grѵ��:Z���n��ȝ#"�U��<5��w�7�Ƕ��xo[21��=L�7$E�qŎ`|:��^��q��e��Vߜ--O�w2�jx�:@��.(Ҷl5\$eT7z�n_��&j�{��t�woŧ��}! p=Ob�
�5XK���^ğ�����HD��(�Ż�2g��2�'"��Ny)���c�r${I@��d!+�aC�u=��;�%�d�h.ܜ�wx�s��7�X^�
L�zP�|��g��	w�d�i}Ę+w �(z��5����q�Ñ8�O���~��ϐ�k�ޯb����V���+���E\��)t����D����o!tn0�Ju�HK�5���i6hZH�|��Z@��!�!·�������r;�}qZջkN�T0�9����I����gh��� ��k�h]	,���J�������8�{p�������	�YQ�h���*��Bn5��z/�v�n��q�TZ���u��m����5{;���Y,���}g�;hdP��H�6���-��Fn=Nٖ r��2T������٠9�J`�^�\��l�gD~m�)l�` b'7�I"R��0����SЍz�xS��2��$D&p����7�tl$�]���-���g�p�������z�V-聆��	�[�
X|4I`͡�l�'`���Q��F9 ����(_�z���!p� �,wb�<c�䕒�&�m��)�\\Ȍ!���A�
����o_���K��s ̹�D�QJf5�dշ��!!ދ*�h��6ߖ���h?v��K*ɝ�o�$徕���Vk&<A}M1k���ຳ)+�J��N[�ܞ��J���g�;2O/n�:Vpϰz���*���y*X��Η�4�Bד�N�s�_�m�>8�y�d�~�S��<�Q�*��$���fH"L��Hn�h�^���_��o��4�IQ� MI�]��ÚT����t�P<���Gn�Z��˞6�sj%X��5\N/i�t1�J��Z�����Ԑ�#�E���2ς~�_E*g/��L���xJ���%43v�����l�"0QA5G�����8���^}�
�E��wTo$���;��1�Brr�寣��o�1��][�o��xH��&�;T��w�8���8�w�����������m����g�3�D��%\�I�7� )�dx@�4�+u�\a���3z:�ޥ!9����NR����謝+�k�c�S�m@FvI☲A'�N��f>�z��z*wyĒ}�vo
&�?̤" �mi�
dn	U��L���ޖ��rQ���������3s�����z�ld����g�WB�	t�T�2��{xד�>����N[�?�Ù˽��W�|��o<�VmF��5��9T�:����q���Hf������b�WU�������5dT��~.�=���-��*�G�@�qg��������4ϝq^ᱪRx�o*?%���"*#�(� }����n�񍎿���� ݜb�w�{9��*����F툎%$\
��[�)�q$p��-��m��:(��9�
"��~A��6��7s�U�ߓ`�,�m�����֯qbB�
��gهf�b'���c�/3������F�(\��{<7��Ð~���΁<2�Pi,�8$�IQ~�F��Y����7�(����x�ox�Z�Z:{��-�"[]֡�#����{�G�|ߖ.zgjxڭ3$,��:G�l���LV�:�e���'S~o��\�b��	����3I{.6�*4̦�G9f%�{�����--;Wp΋y�Ӳ����������z�Ft��ێ׭�WU�1NA ������-̊ǋ���{��; ����}s��z�Ͽp%�kTK˧�_p��G�<�j����^� �,#����!0�P��M��z�n���T�����6�jۂ9�πy���i��֍�ǂL]ۥ�/w_^�,���t7�{��/5�a�1[�-���I"���"jս$��b�Bsބ�J�ʪ��
�)�lF��l��>C�Ǳ\s�>��D��-W�!�"���_tr�����d���Ty<RC��)/�~´�D��Ix��on�x�,����F�~��m��n�<EZ�nˤ�O���4�bz4��Gب=��� ��q��)������6���A�`�XW٘�+_�V1�AC�8�Yq��L���(m��z��v{��ӌE�A�o�v W:q;jT��Ln�.Ԟpn�����B�\�L`g�7?�ݕZ^%nlAgL����0vU2_�v3���^��Q��	������ ���8ȡ��ϲm�y�;a��joh�p��-���;�8�hg@�n��;/��\O	}s\��z�咔I��9�n�����>�}��
M��{�!^�2��?j�v�[<B>k��aPo��}�>�VаSԍ�2u�� �W�W �$�+꜌OSiǐͯ����ʕ��`F~m����
�(Sa�]�c$���ʞL�D�Ҵ��/��[��΂#��0J7�70*�����n8I _��q��4˲q����[�����du�*���q��_��'�O>3����O�vh���[�e��C{=���xu�S��O���4<�����
ť��H�����.$��+�m�8b>U������{�r�Y�KL	'rw?����q�H��C�PM]lq]g�pˋۢ��	��V�dlUb��G��Dw7f"gI��5T��v�g�W�ܭ!�=0ub:��-���X)/�Tݠ����\���Ӯ
�2ꯌ���0��)�Q���@ķ:B��1�i�%v�<��=
�oF��Vz���EqK��O�2����C���Y�)x��`�I������l�ǥ���2LD���ܲnRp����q/����ib=�_%Q*t�vi�(�̆{�b9����'�6W�������%7�1P�0�ԫe�$�I�1�T���e���ma��/�������-��pK��B�����4��]s��*�[4Q���V~%IUN$��2)�ݽ�8M�I%xq�5Q�G�|�ޤ�ug�݅`b�=)�t)O�zj�p�Q��v�|ʴ���L�����x�jC���UV��f �w��#�&�'�ë|U]h!�<�r�8�*�;���gݝ�ɰ������g�t���G�,���A�V�Ew�1=��f0A��T�-Ǭ�G�i�I�(8è��	�G�n����×Z�v�D�Y�s�?���'�^]�s�H=݁��.;�9���Ǧ��t+^]ݛJ^ĂV�^j�LR����=05P���5���:�q�?z`�+��%�F����-,Ry��0��ZB���]����ٝ]>7��s[�Zi?P��_\�X
�+Ŏ�?o9��f�CE�ճ9=�����#�ѡ��������}�z�§zFT��I���m�X��Ct<�E�滤V6<��/W��R�k��E��D&?�;^57I�*�۩xn~2uZ�x;����@f�MKd��Pd2�C��n������42E�=�ic�*�G�:��ؤ�k�E���T�z%y�xlsL�{O��(4H��$D|��%�xč-GP�_u����:e�/�q�ɪ쪓�;�`��*�����A���ٻ� ���%OD��ԓ̎�:����u�x�9��v�(� (_���b���5�ԓ�����d�%!5�"8l3Z�_\���lڅ3W��M��h�'�6���JI�(����i>]�~[J?���o��5y��/�n�/�Jgg�gx� q�@T�i�&���W������K��kG�b���iD�������!���с��[ו��>Q��P�����1̐�v ���i�9�����������um�,�{���9BYy�A�\�@[Mdb�ky�X@�5m��9��G��?-n{8+S���;<���鶪�O4��@^V�p>�0|�oV��M�W�,5
�s�����ŐB!�,�{�E�,JP�VԘ��B<|+����V�V�N�ri�h�(ʉ�ͮT�D���fhBh��P�Ɍ�W�.ְ����
��&J��B�?pF)�����8�����Z��9>���fT�6FNf\�	?uT�#�g���`��F��v��Ygn�i
7�J�~!8sU�x�m�+�ޗ��}HG�cz����[�ԃ3g��|# �l���E|�ih*W�v*P����B�ݷw~F(��A�8��'^�j��Ёߢ�!�.w��\'E3k�w�H��3Vv�9�ĕI�������&����v�u��Zع�O�4�|���h� �>��$���"�@���n������`
�#_qC%�[���.{v��}�1Z�j�'R�\�i6]{���k�L2/��)s�&��{\I�_j�S���.)b���.��L�a8����I��I��0�F�c��q�M���k�����@$1�z8�ٮ.h��Ϳ�|I����檰cr��+�œ��!�q�J��K1����	�դ~bt첒C6WH��d�ܴ�	B�T+X4D�\�G����MU>N���:�����j8s,�5ݪ�!� #T�5��\e���݆��}X��c
�
Q�p��]CU����zv��u�`�e��az�J�]����B,f����p`�%��YIC/>�q�\&ӣKD�9ԛ(e/��[6+��L���>{,0!a�J�tT��-F3\9���f:p�_�����,�첕���9�՚�ww��h8��ď�b��M��'�>v0ʈ0���K{��Ya�4Pm�ҳ���F�����!y_DM�j����S�\���'=���y�mn��J�3��F08�.	5�Dٞ_�?��Τ4���X�C;;E�i	����Se�>�!�/��G���9z������Qn�3*6����nܠ����&�e�	�/�mY��0�߬m�I�6x�!��m��ԌK�P)\2r�*{>��ۓǈ�e��+���i���2���v2tW�JX�M1����ʃC�#����o��	�\�pd��v$�xD�H�q~nH.��e���_qX�	�~�0��+�,����{ssr��)�� ).�,����@�ᬩ�0��9f��������G{;�״�*�ё�9E�H�JN�m~ѯuu��i�s�֒[Us�wF��c���&����Aj��R(y-J`��Y69j��s/e �c�a�	
ZgZĹ���0P�zE[;����u���cSh'��,��� G���� ����>I2��B
Bv��2�`���b�0~8�;�uy��A����^ұ{A([{��7����Z��=��t��j`�+���. ��o�o��:M�~bhMA�>bGr��+b�8��3�����N ���Jm�O�Ԙ9- ��+��x��3Z�������󿂷%���V؈";B��oC�F5�޵��h��� �6x[N<F�qU"�z��/#���D�F��ħ"J��1������1�on���3�3��M������~љ�5	�>�z1�ͷM?�p���D<+�Q:L�|jl�B9W*�
�)�9�a�f44z1��=��k����E����Y���V�)EZ��+(����FQo�4ܧ�U��f}�_�=o1��O�����M��@�Q``R�"�T'������+(�>r�#����)�Űm��c���a`�w��!3W�	9���_m_�"�,��������.�c�b>.�`���9^	�	��}Ї�_���sᩧwH�1E��9�����Eyc5��L���@����.Y����t �.H��s}���/M�xTMS~@-�ℑG C6�
7띥�� �L�`��C��k�kE��d�Jei2�m]�]Wm����/*�oG��4�1|�>�״MDAf[#/�,	���
�?kI��Ȣd�pƮ�MJ	�1:3�'VUqb�X!X�d\5��&ѹ�U�V��x��G�'y���,3�#<�+@,�o�&�q(Z���7�,w�hA���r|	ц�C�>J�k��eC��Vv�����4�
��-�*g�iN�$�E��ߑ8�y�(����1�@M�ێı��ݡ&Y`�CK}*"85�6�4�)W7����x���f	h�#2��r���8�*oر��W�M�嘗�@Ɲ��<[b_J&`j��Ԕ05�o~+�g�[��
K��tԅ"����z����M/Fl��I�k�9���H9��vG�ף9+��c�0Fa�^�'�Oa.P�ZВs�6U+��+��w!�|k����ɡ�d�RbI�l~����>�v�6��ri��~�\���*�Vc}��O�`��u�T������䰼��i�u�_֣�X��OY�5�q5t���W��V���!�rW����k�E�s���2�_VUѻ:����.�肏c`7�v׋L��mA�P(�
'p����]�A��{����&� }�oȽϋ�Q�����<�U3�/L;��M �
��χI �l�#��'�#��p��e[���VLe���_��t�e;ශ�r�h;S����VG3��\6�0G6A��ݴ��F�	S_Y�"�ډV�бB膫�4?��b����ӱ��9l��|Ƽr{g�&�+$��q&��0���|E�q�Ntŏ#��B����
`atT�$,�.yu7B"tԮ�KN�G���R�[;�������lH� _|c��^����R�z� u�.-L2}E
����x6�9|3���<�&����'~����V:4Jrh5ĕ*+��4ڞ^H|��ؿ��/(=<��1���Dg�|��|y����T��7�ICk���BUT��[���������N���E�f�0��JiI8dv��9�Ϲ����	Mu�#��&�\����^H��-qK�R��L���+��z���1��s61J�_ �W�����67���)ۼ�D�nT�������M�����;�R�t�+����j�Ia�O���BKW S��_�էʰ��/��k�&g��5/h���(����T��Q���{�s}�����{B�]H���<M2�W��Z�:�G`c�DHfjiO����'����ݚ�Y:6��=�r_�^�
�[�]q����Q���.Xt�Ă.z��d��u�G@�����>����ㆰ�7u��� ������ThT���fl���U���'O����t�G��Hb��yL>
�0P"Nԭ�Ke[��{��%�c\��Yt��OC	}�0�f�VW���^i����{������d8li��|�iw{̈́σ�]䱷v��T��RT]'���yˉ�?�����*��0���i��Ag�9����Q�������B6J������'��ua֗ {0�M�鉝�uKC���,��k�幭U�T��� �����0J�xL�,ƘU���?���ChY�A�%�kB*oVO�.Ɂ]F�2[O<fD�\%[���h7r(���E���nZ6���`�\�L�_�U��q�;)�{\��f-��m}�@��;F�+u����KG��j��0��b�ف��L/8�c=�̰6og��׈D����T�Y��c��&��I�>�Ł~q�׷�PV5���V���-�+�����0��y5�4*pǪ�ɘi>&�����~^P)+z�U�L��`�ϥd'1-�m�f��L{Q	e͖���̠ z�����~�(�6�_k�k\嫉T�CK�0���k�Ɠ8cV�-p*��$�
.y�/�tX��I�qwM��fy]mf�n�M|���z�0y�,�s�=���A����m.c ���Q��-��@ﶵ�,���ZO����D�݋��
UŘ�X�-�����-9S�_�o3��̼�Ɨ�	�d���A��x��?��z@��x�<�I�R��D<�������a,�T�&�9�^�:Q��d"����no�U3�V)����r�#�v�����u���+k�Bg�q��I=w���.��5�|�u�(5������u����=����U�'N�X���g��o���Ok��
��V,*r?<wf�q�^�@��O�e�d���L���9�F���GST�:�����:e�u���,�o\���/jܷ���|g�I��^��E#UM^����ѽ{$�m䇌�`zȴ=Ƹ��z��Q��(?��L�֝ag޺��_@A2�F�]�z޸�!ew�=+��z�v�T�ظ]�����d�Cuc���f�$��VgO��t��/ex#,L8t�@ӝm2>.ߒ�����k���r{�\��6xHS��=�M�l�H=��	�z�2�fV�?�=��M�)��2���(4!f�p�N�t���P��f<�!�E�����qm����}h!!�G�<�7{�+n��q,�e��ˤH��+)��}�,��Gz^3?+��<N�r)ȸ:��k{�B�!2�H���ױ��j� ߵE��H��"��sG��;�5Xfki+�Aܒ�[�m7�SN�s��Ji�aB<�s�}GI�$���\Pᑺ��ky�8+'�,��}8��4ڎ�'6��.��<f!4���A�&���8��f�ϛky��{�%�tt�T'���<�Gb�T��j���� �1�x����z�Fr���4Ï�,>d�g��Yh^7{F`ʒ�J�]2���(�ݗ��������{9V�'a"H�&�K�w��W�>��D�*��N�����Ȳ#�c��d�nz+@Øw� ���4�������y����<[J;Z�=��u�z��x�G�Q�Aa.IǾ�-I¾p��{�xy�͞P�Xv�1�f$�, ,���r7Ć�F�����j��v�,����]7,��=\.hs}P�s��c���ǐZD�3=���@u��%H�2Tp��AL�p%S��ɘ�4-m�$Q
y�/��;[;��k��~VQڕd�j���	����vN}MrD}Uײ�iMf {�<��L�:#UeEH
D�$��	�u`XsQ �I��MW�r�b^�5��o��{�}���j�؟ =ɯ�*(��l��m���xڄ.<ܶ�����	�L2��Q�GM��5[4���u"��*v�DRO�]V�S@�%QL#C}�[{=i�2���{fM����O�W#4�[ x�4�1��Tx�	�=���(��T/�V�?��|C{����N6��ާ`�����lwр�#;8��^��������2���:%��(v�q�>��@�pVR.!������D�-�ג���w��p�O����W�L4��|HKkLԦvq汔>���>�o)e&Y�Wq��0�7�Y�88@���!+�8G�s�(�DD��@����\�Sg�뇼�!}�)�j_`�a�}M~us�a<���6hx����8��q����6MAW��<cIɭ�-�UF��0z�s��p&�%��2�J;��k�	����r*�7HQ�,�[�^�9�B3�>MyHd�!D�1�_��=4)��4;5��@2��J`G���v�l�tp�CR�1�j�#<�����sv@ 2)��W����
V.��y}��rs� ���4E����!z���/�d��|�L�?>�Z���� G>ݠ"f����{��8&�$�b�d5�=}y}�Ŝ�Y�c�*E��c�C���<BG�lb)u��(��!�B�Y����X�FTȎ�&�l��r��5}�������شYދ�ß���o�����FAȫD�$���̑���B��lգ�<M�����>�f�V�t=�gs�5������u�s��YmQ��9��KbM��"�!������i����d�k����&Rk��,���`v��9�Ո Q+]w.��sX�R�_�G6J?�n�l^�
�|Y�岮 {%' W�m%D��)�4,Pa箁�hn	�H&50�l�MJ�s��P�һ]������@m����E︟�ٚ��)���t�����&�K5 �C9l)$�	�b�׋�C+�(�M[�P���¶~�ɥ����[������d)�G���˅z`r�(��s{i��c_�N�s����G	5�B��y䦦���HB:C>�
�����8aX����`j����l&!�w�Еlt��sGO�|����M܁o\�sQO�-3���&��w��zo׏���*�)��Z��Euc��
;���K���I�h�G�����@��RX���Q�)m�<e��	6��iu'���f�!ԆF2yIbyv����1�d�3���;���$�9%��Lt	n�5�اޡ�������S����eh]����m*+�&���9KrA����³����
ퟯJy1hh?[��nyg8iS�Hq!�X����G���jKZx������B����N�*y�3���$�ܚ�Vr7�v�.A���ݸ>�]��3��ŰW��4��ā����_?q�X��mt�v�{z�s :u]V@c��ZO��~�C��)�)� �M�ʲ��j��*��r)�$�� �K���u�%yx��-F�8��@��W�Do�&�h��.|�VUc�nsu���z��r���g�W�ۣ�u�1�Z8�P$�0�a��^<K�;��l�6��ƕ�V�`5G��|:�+�D�p��C\�0�O��lmr��D��D?�!J2r�1���?�M)����qN���:�㑤~����!�h�vD{.�2%n�Π���;Ru�+s�OT��ğ\;�����!�ӷnE��,��t��?�BӒ��E7�����yN��i�:�uL�3�U��G/7��*��iS���k��~�,��I3І�]q��w9�^�U�+�p/)���*{>�,OT���Gl��^ ��"�v$�������v�q���,Y3t��m�Î$'��<ݜENRڝ!0�YAK�
R?��c���1'3�*�.�#�7*R.�=	��\��g\�e�#>�4~-�pN�p1Ə�L�ՙ�����uU�K&��3-8}pA����?����@t�/�~��.��fj���'�:IA�f��Qւ���<�����y�̈́�/1�����\� w���n{r���P�CK��$捜~,&��D�ֿ����I��w�vk7&���oj'y� ̣Zv��k\�����U�pF�ฉ�}K����a	k�3��Np0>{\����|6X��ɺ�DI ۃ��:�}{�ah�F�9Ud7�t��*�oε�˶�lz]��s �}!�KDVؤej`�8���k!3�K�0�6�č�H(v��X��J6�����H�t F�@P���a��Ӕ�$�AT��6� C�7L�CZ����i0��R�:�E�H9��n�q���c׋�C�X0��,��A�mE �:���}�Vk��:a)���Q:�wI{+����-�lr)@�x��v��)�:qH��GS.cS��n�/�`�T5��Ǜ��&�F {���E�r߰[�9��#�(��fފU�_R�i��J��"��,-J�{�H�g:�pw��ue���C�Տr� ������TS��:��GU{�0��t�W���k� ���X��?-��SO\7�ꠅ�*$r�N��pH�Hb)��29l�q�?��><���(:Rrg[��<\�:�ă$�8�Q\��i �=c����i�j:CV�O��#����l�b�"JV��^R��I��^���;؎�Fv�ߥ�/�W8ˊ���%�3�Y�,&��@\�Ȱ�ef?�
�x3�D�	�, EqF�0�JP�!J�ڡ]�#:[P�t��G��$1���*^�y0��*����<���pah匈��|Y�@wjWi�q)��}55��\R7��j�;2���P�j���q���2aܱ =`Y�(����ӛ��(&RcC�v�&>	 vLSa�_�ַVMt N���闓��b���Y� 0�ᣃG1� �J��N���%ڜ�h��ۅ҄7�pUA&�ȳ���iy ���!�F4��j���%y�Y^��ڪ$Zv�y�Z�d�h�� �����e��̦(,g'�Er��"A��V����'���N�ug��,!ݟ��,Z8s�[��v����!$��3	 h��-`��Bߟ6EL0�ꚋ�pʰ���q��W����fnd11��ߝy��R�����Y�5q ��?��`'T���-kUKs��9�E#��k��U�e��n�����c�Դ+Q B���2����YDz�m2aF�^r��@�e�N��;t��A㡙D�54��܊K�v��,i?�~,V�p����[ ֜���%�-�?�KSǏ$��!O8c��:U��:g+W���+׻ҥ��q�W��v��+pe�i�nB�L��s�W
������E���dԲ�V���~~|}��9A�u�=ȴ��Yy,2ڛo7ܰ�i���n`��{����Yӹ�T{\iքv��J+�Hֺ�#��GC>=�!��l D.B�\�7�_}#4H�¤�!��W���)��Y����<`��pE������?�D{&c�R�|�|V�s�@���:s'�#�d�a�]Gr��1l���T������_�apD���6�Z�]'L�C� �U:r�پR^2�����?�F�In���C����X��3�v�w�vG5��)�Z��!�d���f�l�z&?;���e-"��+�T&w����)�7DD��UsO�,��R�)�t�,�×��� <��h��a1ڱ��]%�ǱYaRbs��(.�%������Q�@BB�\Г?��A �\�FT�`h���E:]�	tņtHO̴� �c�(ǒ�P�a��CA�h=}L���d!8y�u� 9��r�6@D��q<��%M��j������z���fx��AA�Ȥ�[���5�U�9NW��9�'�^��U7��"��)�u��P�r%���p���*�1�c�46��B)t�J;�{I��a[����Q�jfs&+03�6g�����9#@��o_��������'�%�5U��Ȥ�:��ݧ��֝�f%)�?}����!5�Q����Dġ�܋�[�
�!g~�P\����f'�V^y���E��:�HZ�0E�LH����=��x�5�4TiY��Em��&����I�f��ah�j��V0ۑ�0e�1�Y��|�s��N��g��tᚊFyN��5'�l�2s*�Gh�M2�	��_�>=�$��h�g��0<�'t$�7�B�t��!X-|뇿$on�#�X�I5P������WI�ψ�8�����)`�2���0�u>����IiL�M�?��y&�E5��뫆�h�m��6��yh�ӹMel*�޶l?�}Tb�>�\��2g�bhQ�4�����9�����5�K�eg�ꮷ �[�!�y�?h�/��|Gf6J2q�"ʱ��&�K�`O�S�*�W<��F��Q+��O�~�8�u��$ո��d9)f�)�zb������A�e��>�b��uc4|4��������T�Z��9R�RET˃+Ps��~Ʉ���(v��� �GJc��v5�xҷUx��_�Q�x��]/{}��q�or�jF���`���1nFs���:�e�ѮB�M�R��V��(�z��.5Wτ��JSI�y�w�5��1�������h����.*u�n���,�6yؘؾ���,8c���k��2+�r'�T@�^%� �~�0���)@<�0\*�֘I=f�i{����g�N->���$KQ��M$�;��#�4��-^��}:��1�0�6^��\�؄�ߣj~O0b���i���L-a\����v�{�ԥ�\.*�t�����
0��+
`�E7���~U���Az�_�]ܳ�N�g"���3�n���(�휧��������X}	�;�v��+��X���]Gϭ����o7�o(G$no�gy�D�Pe��������cp�:q��=�,"�{z���ڤ(wYH/<�V�c�����O[D���crڙ��lfwdR$��a0��m��.��)�60��w�0�!�$y=�9#B�ş\��>y��[�F)h�>��O�`�l���?1|�����~���ě�;�Gɞj��MI�@�<��`����K�r�A��+�ႀ��&P�@P�$�����[��k;H��`^¿��K � ?J#���kQg���7��z舞�r����=�5G&�,�S�CZ
Q�0Y��S
gq!O|ZV�i�S�#}ci)��If��B����Z�c�^���z�:|����[N�[��o��7H>�OS\� Pjr����v����r&x�;~����b���p<?=������5tE���~��4��S�����}֐�g��&���j���b�7�l�>΢`_zg�ծ0mOĉnL:;�B�(U���T݃
q��i18)[sUن��k��6s�䙷Bj�DR:�k�����gr(?�x��z���R�7Z����Y�7�r-��R�W� �����f�5l&����A2�rKi�RN�����6E��(	S2�2ɞ�������6�F�J���r���5 �]�W��yN�10[�Ub�Ld��"���?���ݼ>���V���ˆ|;;�
�$��e����3�\���)9�3F��H*4D� ��!�\ji�I��|a��b�31��\>Ìʗ��<�U�J�,Py}���$�E�F���Yc�o;t���]g�2J�|MD���w&���(mx�<Y��5[���>촪rb�?"��wڰ(�3�+��r���X5����tkEr��kf�'�6 �':B���.�1���R�@r̭�?��V��(��w�qR%��"@�$^�W@��^~�;a�@�GN�R��K��$�w5�>�T��{��-T:4��tt��@
�xd�3�V"�-���b�˅�ռ%��I�r�)��!�nb���� �l�}��՗����@W�c��MG�����]cר�o�!��-��"�_y��Տe��#gT�����y�� ���3�8eS2a�ar�:T��1�e��ͳkT�!�p>E ��t�����h�� �6�I�A$��4��{Ezw�����Û��p��� ������z\4̰������I��)�:�?��m%)�	럴���Ѳ@�x#;�v��Z���c#~��3���~dD�j��"���v�	��zU�l3����(>��:�&Z��sR"Q�d�D l>�oY%���Og�U�X��^�yc�	I��x�%b<o Q������c)`\2%:�L�3���=f��;,�
~��� v7���Ƨ�[����0�^"���w#�����XH�"�B*�
vB��=(�y0pz��ܖץ�8(�H��$Q���ˢ ���#�������y#�Uk�|�s��Wy�b#�p�WϪ=�'�m%&��e_��V��`Lu����B�� 1H��p[�ckj�����.*��}煐�)��R���&9�o[�Jp��V��xa�K�$X�
����$֛��?|d���V'qH ���������\��$i,��3zM�/b�#����Q��H8��~��!�E_n`Z�d���1�&�Z��A�H �T>�E�N#���>pV�a��f����+�ɛQ��c�]D��뺾����I?:��ZH[��؛9�x)g���3��Ұ9H�s?)��إ�ABwJ��h�8��<�/XkL79h0���Z���v�ɕg���'����fu�C�s�����6�M�� �ѥ=>�5]�+�]�E�N.��zS}Ĕ��mťQhE��v��G��W0���ޓJV�H$y ���J��<Ԁ��F���)�x� 5�4�������x��U���������Љ�!vDWN?G��ӵ�jEG��S����(�M(������K�n���Э������.	?v����X�8�"q>?�׸)lK����M��rW8N�.1>@��Q>0eK~�2O�$����]�iS�,]��4>Y���Rc��s��I���u&M��t�4��u4�Cԓ�����U�Lmj������р}SG�8el]u5e
��C?���Y�;ڔ!���֧ڙ�"�]c���\�]b"l��Ȼ1�츭g�Y����q=��K�'2������/ϱ��c�8�瞏"�Yu���)*x�p�$+�x�Y��e��
��s�����=ơ���I�p.͘KR�1�����Hʏ��UwҬ��l�[T���$��͖'��`=���*0u+4)������@N�	׬`���
u�h���i`�8���vc��Ⲱj�N=C�s��5T��q������A*�m\�j0��P���y���f5�@C�gH��q�5��B�A[��n-��)p�$�o�W`Ւ8n�_��om�c#�_�D,��ް|y�b���驄�0�W���H�,�.gk�)�-O֚���әpk��b)�a�����A�_sq�x@�����d(�c�C����~n���xI�3M�$F��0P��=`yi��o()�+B�c�n�Z�J�m@�7!��1�O��w�7�]�����
 �
�O�e;:�%;HK�����g&�Hl��k잻��m��-Pc�&�
kn�����P!��&B�����O�F%���Cʆ��:�\��Ó}W�&��G8�Vj+�:a+ޭz��Fl��g� �ȉ| �����>�a���i����[<��0��k٦�[#B��w�3)����_J�N?^eL�ml��gf`?}�A{cR̳,���p��F~d?Ao$F�?����4�hM�ּ� �����ͯ�����
F=c�N���z[��=���}�8���r�;6H�:����6�M���9�����L�3��5e������ə�p!����Owh[>�@��4�h�\��3wV��J'�=���t���r+�r�W�E�$��N9�J�ɱG=����i��S�'�N��R������l���#��y?������ϳ����U�&�����0��Z��P���_*(7\:�Z�7���(^�I��U�\I/ PHM������z}�f�Ol ������Q�}��g,�-^V{.�)װ���0�U�gZ;oB�5������M�V���m�����`}L(�q����^�����O��-�O֫��cK�cz�t��d�THT��1��A�[ ���ڴ�1�jm��'p�����/� k���;���%����H�9�q'z�FPg��owT9�(S��F;sƤ�ff�����,d�,�gx���|�Ʀ�V����̮�#�7<
4���'�ɭM���y"Ys�L�&E<EV��6i^t[���V���3=H�$@>ƣ��6�}.�Z�ݾw��� ƥ/��u,0�]@D�f#�g���6��ZL����^�����=1_�Eõ- c�b�B2l�o�~o1&��r}7�`���Kj�5�J���rFд���*��^_��(�"&�f	�Ĳ<g�3 �u���'׀�\�Ps�N�?�[��⺼��8�Z�;zi��/2Hn��~�`�Զ*8Kr50q�9�x�$�g��
��r7�R���m�Ɇ�+�z���p��8$_ٱ��:,F\U��m
]1�g"�����t0<��ԇ����T����vm��,��3u��Q��L�~�h����>���a���z�͖J �fn�`�͖��>\�'����5�,�lY��2{"����5Ѻ���+"n��ț��9?�e :B��y8��ي�B ���m��Έ�]�b�BZ�} �rTm�Q;H7�
��2&��j���c��E[g�ٽ^�e���$���k'�5��6(�"�2
���|p&��!d�т �U�o�i�sZekTM��MW�Ig&�v�F�?��g��Kc?m&��.O�Z�t�O���*���$9�8Qu&V/���op:��w[]xݸ	�~�'*OQ�U9��_:h^o�$j�Ip�ֲ}�'�
9��(`z��b�th�b�'f`5��W�	𚄞����8�o}�3jh��пM���� 4,Iӓ�c��
�hE6<��Ѭ; �Z�'�3��Ӎ?P z�|�D�Yw� �g�4:7���$�YU�(V�[q�؏��r_�oS�ym4��<*J7�ژ��q���#���U+��3JSUK����I����$���$��w�kzG�-�gp�I�7�RO�Ʈ��y��AlĹ׭J�<�d���W�!�A���k�!-�z�t��zԃX��x�����LY�ڟ-���X���� !)<�ln,
~ �ﱺ��i�
+�ne�BR]m��z!���uy ���C�1��'x>�ּ�;�2�SgYF�\6[_�<(��H~���7
���{V�c��Cn(]?�b�a��җ_�6��9�}}�jN���1C=�I��2=^�t"�=��+�F,�,���x]��˺9��|eR�2}UA���s��r�
�������.p@ǚ�s��z�| d�x��
��b��^��
ɑ�ˠ�.Y�9g�uqê�z$�M���d�G��|U����x������:~�˼?_�Bo��5@�蟐1���;�FwϹ��ZsJ0p��yC:���<���9傕)���T�]�QN��H�t/�<�!`�H�Yev�������'��(62��PC�	�D3���n��=��8L��7)b�"����QZ�ra߶0��aA�g��%�ZQ������dfz��83�b��z���%�2P��kC�p	����HG�4af�ǔ��+E􇺍$��<)���jJu�Y�xD�A#d�w%��ڽI�y��^/��v�r�{ց�6�h}0�B��BH�C�{�	Y8Ȉ���� �E�ˠ���	?!���@�W��p�@|���N��������%|��j�7�.���떹d�ɛ����`�%�`Mun���E_�P��Xl:��1���q�`�?�Vj>��Ks�I�m�������������
>0Adq7�!+X���߈�$+��1�h��o��o]hزٶ�IVʎ����Zk	O�}�:`�[`�څf`�{_oK��dԝy���G�W�<¯
���o &���Ik$��8P?)�y�e2�����XjŌb��!�F�V�i��CQ��%��T��v8C����w�U~ZY���	�E�l ���1�7P?�v�e�E�U�\�@��Q�j�-�Z|9jVfg}��:v��Ý�U��_��1@�~�����=�
��`��Ӵ��x��'��#��[�t͎�/��C�����Ҿ�U��@��r� _	o�ls+��a�AW���
�@��F��r��	gz�bV�����Ӏ$� ��Ki�����Χ�o�6����X��2���TLPK�|9�Iv�:�����:4W��V韲b⃼�`*2�aw��]K-� �:V���0���?ްܿ��@��J_�@��w(7�q��Ȅ��6��6�B}�5V���HO����:GOx7\.�L�ւ��/�2j�y8�/*�3U�Y����-|�U�s��h����T�Πߪ��W�3=S�V���C�+�/2�P���wޗHco�#�AM��M]�H�'ɮK�A��!vߺ����c�׿��b؋61֙Z�>#c�������Mv��'�>��Vة"����:�΋�Yݑ*Z��Ͽ��n��м�#���?��J ~B�֍{ ���\A�ax�]zn@� P8�{��Q)u]����\	qe��퍍�H��f���V�sϾc���	��\�Qd��������!l�E
$�=u»>)��|�?���9u�|��G�L�9�������b�\u��F�)���O�Q>;H'���=�'����z����y��Xl��{
�1Ph�c�O����TEy�dV�d{O�b�/,Z�J���5'�&�q�*9J���o? ɭ'D�7�B�wU|�ӈ�`�4)�&�D�����fĘ��\C�"��)y.o��*��-9B۲��aF��]9W~�VW��I�hg>��j��C\gё��������q����+C V�`�N���$XQ�-�f�A��!��8U�і1�&S~*c���5́���(����
����"�(p����ݎ������CU:��u�,������Z�'���Hr�$]�ۛ����
v�C�Q�X@O4A{s�B>�@K�`/�|�%p��D�ί<R��(����F銘����m�-�Y����2o�����J�������g4�;9KHe�&�_��j��Ua	�Y��Mi[c�V��s��܆3)�R<l���q�1�IE��s�R���������`L ��؛� �*����s ��V�J����ϋ�p� �i:&�/Y1����kp����#�
�#�l���
�L5�'kt#��N��'		z��C�b(��6^t=���ɽm����Q�����}t䇢�,�ӡ�I�O���$|�B���:&U�����oxS�\e��	�|PV�y���EHmT��9�CV�"���*�-����UJ�F�g���I_�7��7��h��U*����f'�?����#c���mC�8@��3P���&������U�	�R#ѥoq'x�X&�rꛝѶ>�$7̤͇��{��*���A�u`��e�.d�yz,#x]�$s��P���lc}q'Ŏ��۵=J�Q�W�&�ԟs��T 4S���dZ�H����Rk���ʘ��yk22
���E>\�M�$W�]��$�W�*E����3��H��ʵl���D��8h��P"���&Q��h50Ɋ&�����=ۡ���U7�dp�ޟU��$ƞ��]J��w�Q!b��S�(�L O'��d�9ezD��lI�Z7@G���k�8K%"�a�(�p�vE�k����7@!�ucg�SsQS�׌�8�Z�J �M![���2��g�x�}�(K��I�rފ��8���8k�"����Ko��\���o�m��kh͇�~�F*q}> g��ek��UA!�36�_��Gz�'�o��Wã����Wbd��S�Ta�e�u�ǷyR�޵�� �p��Z��tV9ғ+��������^~Iw�2s1��#�!^��Cp�oW�1��]�|�Wp n9�O�@��z6 �s5շe/FV��_t�Cw ����d]��cb�;J$kh��ˁ����'�Sk�,�ȶ�L��g�[D���faYۧ�F^��p`u��R��F��&�j�Z�R��KԂܓ�x,��� 4SU=��?���i9�c7�����Jۊ�n��wv�`Qt���X.B��0CJ��S�.ŀr��#p�}�����~��a��{{:�3A���O��.j�w�B��+��s��������ʄ�Q͖��H��;��.��u�ᥣ7�w�i@wN��oM�f��	�}ޝ��J�yg�a"{-���WD�X]�]�����:u4�%�;���ы�\EhM/V�t\V���N�4��IhM�#�$�[�0���v��O��'}�qa�X~��*?�Xufp��.��Ԋ>����x����_"Z�Z�êQ�SWE�,�^��}����GG	j�a\����N�Ñ�;�'�v禁t�؇p1n�IA��u�qLӠp������1����z0^w{r~Qm:W3�Q�t����+��S��v��c�v�� ��4��������P��>hc��X!�|�g�����tߺF�?�ِG�vEp~��o�g(m.D���B~!
��UO��x�=9� �	�Q����<f��U�ny�J�m'lM�I�my�����֐7c.�sEz��S$
��I��a��ߺh4�VX�c\���~s��^T}>�ݟ?פ�0��s�>$���|;��\�n�� L�{ёl���g��s@���/*+RY���Z
����w+���܃&�=~�<��rHD����M][<c��<��}���c0������*.�+ZB��4�������*=�b���������&|UW�ϒ���~�]��!�Y�g�es����ZV�Iy��t�L$U��@_�"t���N��"�KK�YT3�a��
��Ҿt_r�e�	�ӯ\s-<Kjd����k��$�-^��n  3A��I����'h��Z�Ə���)�}Ə�XZ[��ϛ����j�}�$��7:pf�Y3��@]�* .½�P�I��܋V�K�"V�e������`&���,]���9��&�����J��" &6�~]��;Z���t��|�"'ʤ�ೋ�/"eg.&M�b���`l��]�n@^Mi�'�68��Nﲯf�+D^ڟ+s��k��P������O�����9^:L3���5��>F�	�?��F�a�����ނ$bZ?�H�`�/�#�,�Ѝ:=1}��#�V��Ci{���
f�|E�;zsP���ՌZ�ud�:��;V�������D W!$ߒ�F����w��CϷ��,3Z(�N�C{e�4q6^��\��v�U�����V�U��,��ta�rP��7�m���]�^����������$��b�-jh���PA%[�+F��0�����q���҄52%�-�q�ebf�ɻ�z��d$:)J_Μ��Q�u��#7j@)U�Z��E.�E��#�(PW�٨��a.�K,U�n/7�Ĺ:�;v�y4�qZ��@I	��tK�vd�Ț�V��y�)�O�6�RRl�dRXCɼ,�7�w�5ZbRc~-�MI�th��a�6BI�ꞗ-����ߩ�XT3x��W+�V�`���-R�y�mʎ�L���|��.K���C��95-5t�@�����YuiQiT[Þ��#���F(�5��P8]�:�vP�w��+E4ֶ�,�]ߝ_W�?�H���#�Ȱ���cGTF�o��ڒR�*^L�j��U.W��1�x����<��y3	�D�,:�v�2�N"i?��\�>�_x���MR_�[.��@i��A���{y���|o�4�'�7�𒯺�����d؂F�BlrbM��!�+�;�\ݪz�#[]"GX���^�x3�K��ǁ.�A�'� �e:�����j�Lh� ćw�ݸ.�vxS�2n�YSg�U~8q���a��J��Fn�v��啒������=���_�Kiv�S�B��W$����������8��#�ݠ�R�f[x��u��{�)ܥȢ�w��S���|F�[�w5.J7>��f{
���y�u�(:���I�������}�D&I�c�f!��A�\�oۇ3�7}�W��EN�&�X_�S��M�]�L��yy�~�������yט_��uܼ����:L8�x ��CN���`�m��(Q�KT�����~���ԯ��-��F����s�_Ѽ$]v�@ڶ�4�X��.��!$���<71��bH��/Bf6�E�װ,/���O-p!�)ɢb�)�S=��kv�a�Z�z���F�9fK|�= "�U�-���~�G�'ְ���<��o�g�/HB�<��Rf�YZ;���ϛO�m�ƌJ��s\�%��pT!�Q����}ؾ������k7�H�Mx'}m�*w{�q��<M`̢/sW܁�; =_�&��I�FAp������c��X����rV�`�������.���z�ۥ�F���E�c��O�}�6�Ƌ��x������$̣�,�o���f�9��Z<t������5�	��&_��<��P�Ev��J��fF�,�U�&�p�V>��j���.3c^%�|ԏaY�0�\ɵhMYBY5�CY�Onk��ݫ���{��t�oNr��/͎�U3�>���hqf!����o�g�
6�[��9��!
mS։9C}��I�=�5���T!2�H�_wYpe>�	.��gԷ"�$�qۜ�Vg�ݜ�Ӵj��S��V�"x~��o�m@�rMc��>�V�9;�`t�ĽR��Q�7Z��]��=/��l�%��A&n�<�C�$�Þ���h[*��e$�"�8ӷW������P�AL`&� ��p�͘<Idx�O�`;��,lO�}�Խ@cܣ��4�U����2��u�t��O\D����2*Y��C9tE��&���х\q?n�/��f��%u�H�ai�b�7:�������H�;��wE�	sca$�\�63K�j�;���b�:o�=�8�0W[�]�.���Y�de�J��2z�5G�ckYANyo�5@�;aü��Y3����K��T�'9�PY�+1M/%�J�w�dR<Li$��A��#�[�s~�PFg:qR8*�ֱi����»��\"z��#<��#A�`is��;uE�n}TVM��o���ޗ!C�áP�f�e�Q���������4!���������>h�*M*�'/q^�Cn�a��e�X���<�7�I�-5M7�=�L�&Q��y-����[S7�	Q�m�>d.����;��kT�c�LK�(��r4���Z`"Y�ꁬ�V�j���KBeCⷍ�F�4Vn�D.�ݜ���EP�"���RU����,h�dF�t��+nY�=/˿%�aMu-�N
{�пן��)�ѵk)�Y�\X8d=�a�}���)"�Ō2�1�zN��8yC��aS!����v�3�������t�`E�3�� ���q4�
��;Oz���ؔ�L���xF�wQ�~�e�&�ԋHsФ�̨A%Dؔ�oX���&(~��=�4��^%̙	[����C/&$�\�%x(=2[ezܞR$��b ����BWN8��6!��>Һ,�Q�@�
�R��=�Ъ`B��|ȅ)��t��n�q�R��MN�����~���JzlH����YS=Dݙ�yCz?�w�R�<�X��ҎrM��,��6���wD�Vܗ���a��q�O�Y=�K[MJ��_� qz�5�?S��&�y-�}@�vg�揯�c�bdCg[�/�7쑆����A����R�E�a�ߌmԩ1�O��Fn`{ȫ����'��6�ii$�]�[�7��vw߷�d
�>�\n�
b��Y���k��Zp�k��&:}�(f����\`j������́����
_]O.?��0!U�^"���l5Z�QŘ|���v!����|��cƴ��n�7����,�$�}2��V����O]ץ��� �_N�3���*�g�x�d}�3�v_�|�Ix���(��wP5'^��ac ��dBy���T�U|�\��B��R�Ws���������d����������w+@��CY�X ���@��I�&��h��U�R�n&U=V*l�BF��\���@�D<�N��Kޅ4����#o���J,/�9[ULk��ң"��	�f�8����i�7�G�Ns9��n7U���.��{��f�$J�ާB�)�L*{gm:����6�w����z&=��K��B�����Q����9�uՔ��zNܲ&�feHY��w�>.p8<�(±�A۔M�k��Q e��M��֢����N�ۜ�Ip"'E^�_sx
(Ϋf�u?�x֞O9���n���ԏ��bk��E�I*���|YWR��k�i:H+�y��DU�}���-�\P�Y�c�>��B�T��x}Q��KX:����-|�R�R� �g2�]*~��J��p��-G6n��B��K�D�MB�r�,�\ď��gæ��<�IO��L��nJZ������BM� A����2�K�Xp�w�b����;П��VMP�Z�ma>ٟ���Q�8�_u�	�]j��j��K$J����#��L���_�T2x�2W)(�Ά:�>^����"e��_�����v���2��K���B�Ho��x^k��3h>�[�Z�ȗa���kK�kF����uk���4��<J�%������V���?j��q��k�_�K�m!�PAj���t�p`bGq,zYpU7H������`G|L�v�sB�qljk�T�y0�{�Z�
N�2����6^1�P�GU���\�79��9��}�o��7��#�.ǻs��uH�d���RN��o��
 �A�O?,��������:#�p�U�gY�����=���T!j�L�]�`+I��t��?���F�"m������@���=�tNYI�
���׏;RG�C�J|\ � �z3��U����� �f�_3�s}!�k<�M$�K�Gշ:ՂM���c�Y���H����R_�Kx�k�����c������G���fZ�@'�p��Ʊã������g�t�=%E��Ji�ll��?����q�5^�K�/�2}�Ƥ�K\AT�eF'"��:�r�%o����>�kbβ�)ۛ���)�V��J\�y�1BjJI��A���(�Af��k���77#�u%�V�z��K1JB3,_�4�G�^ �1v�E�Z��o�O�L��񟼉XFʯ���
G��L��JA"�cɎ�@�Ebm�@�K��3E9`�|����`L�݃f��+\-7����<`�S��������._T�$V
 �\{�]�不�BpH�F˞�oAM�`����m�J�#5��$�,�/��=��)�PD_�7J~�Y>/��ɟZ��r;��z*�يvp�wK]7+�L����TK�η����W��!*j	T�2s�U�������4���l%Iz��݀c"�su��q�y*>ٳ�'�u�fdU�"����9sZe��י&� �T�Т>�K1D�g���s�M�Q��^-��
���HK����:��:���g��G�\[D���4��[�x�1zn�Db%�J�������M��|�Vhi>�h�_�w���x�J].��͔�|�	Ͻ襍N6�h��h���@���HFR�IB��� VV�t���|�oy�뇼���2jSp�
-PW�Z��ȉ���ÜI͜��?�	�(Nr��5|͖���eW>�s����{�����K; �>���d�����s��V?���dQ,�ݚ�u��f�/ʘ$�j5���0���?���:��a5��m�$��c�H���Y �W����t��P;���j2���q�����K罇�s\����.C��{+D6Sz�-���o5	�����x #��H��*�]p-���w��YQ\d>��O�m���}V{����%J�����ݘ���a_
 5�3N���U�����OD���؈���ψE��LYҮ��m;0n��}^�����H��,��g��36G�i��B%��J4vB��
8(�5`�.Z�34\Uf�1ꥸ�}|mt�G>��`���ٔ�;(~���%Ұ�>`�i�&�Љw���R�9�Y`�S=TJz�Vq�K���/$�%��f�;�c���.-����)w;��m��h�@W��T���-v��<�M��aR&m����U�HURN>���@�cmUrI{�2����z
��&��s@N�)�	�����w�g*r��X��eI[OK7�0��U�!�M���z2)^Yc
X,ū�G#�X��/�v�[�Vc��X�J-��Qؖ����k���_��P�G�;�8�;��h��(A �K�HD�o*�i���r ���r<�䅾�>�Z
h����!N_���+#\v)i���'�8E�g�$�?���Db�&"e䃕�NH����އ?S
�<�A+�^�������'>�A�_������M�{��b�YM��&ZC�V�u����N)�j7�D��|&�[%����ib��/<u(3�0�G�~��	���8��YZ���И9]��ǅ�#ѐ̞t#�˟96�Bl����
5�_����K�_���W��ǄKU��ta�Q����6Hӕ���������f���kO�y�a�յ������4�J�r��x���`��vH������gB�iF�^4|�=cə��,<���?�-�#��,%s(�C�'t}�W7���@Y�UTP�Ht��^�w�a�����Վ8,�C͹Qf���C�%�z R	�BЧ�r��˲a����`��ڟ!���{IK��p�����Zw��]�9��D�N�T൞�������#Ul�l^�����������sˠ�\A�Oɾ-�a-�@Dy��1I��s���t_hs�~F��K3�A��x����k�fS�L*]_�=9$�ݙa�kc���(2������+8~��o���������&茊�'�'����6mEC�ڔ�|�6�^J#����'���:�9J�P�O#�'�<A�����63.̕�[�{O�s�Ko��u|D���ʛ���T=��k������q���M��� �F���;�`�]��:��Dp�
|Q1�Syd��]圛�f^,�<�H6<�n�H1�:b�Bh�O�8�-;�?�}Ż���Q�q�~�0*X���Ӫ�Z\��ҙf/�[����u� B}��<D���O@` ��1��c��Z�oV�+5l:���v榍�	2��_z�ub��A!6�I��F��(�=�l�ڵ� I_'��Rc�J�������~Rp1�i5mS�z�#$�U#[Gs�b͐��������=��A�ݔ��Z���GU�S���z�UЙ���w�I�>Ϝ(��8�Xخ"Ы�����*��x�U�1��-!�P
�E����PVF�X��7Z�Rpo�RH)J���%򒒉CF�ڗ�<N��|@���XZ\R�'j�/����]�7Q��bzZ~�yq�-�CM�;��?�a�t��&6�Ƅ�Vs߷=n��i����a��uܘ�����%�.hcn��j�(�Ư���.(�*2]��s&�@�t2��Sd
��59���Cf~�p�~���:�]_��%!B;g�c�̌J1�ơ~i�D๾%�D��4T��[�D�����_f��P������eZ +�,Hy�ʯ�dTxl�^�5Q�t`�к��b;a�.1ޗtq��ki��`���֡�˔E�z)U^�]$~Bӯ�ei�Ӗ�]�1�a ߷�6$��1�x_��o��˃qT�~t��@�>~��Ⱥ�1*l����k�[aYƣ,�M��peK^��gҴ/�I�g�zQ\���oE��#≾9]%�i�P}�AϭA?o�&!�6����7}k�t+��r4� ���77��~�����*$?�K2�O�3���N�h��%����A[�V�_Z���"5@p��r����[��*����P����L���@3)�Y�����e�(,�Z�jbTየ��$o�'BKBp�xx�}��3�_j�#��n	T2a@��k�|��oJ ⳨`�<�S�z��D��fN�h��LO��I�Z���S�.�4�y0K:�{C�p�ۥ�����W1r�r{A]+݆R�op�{�q�&��j���w�>
B�e��\6͹3!B�bU�T�ߣ��(�phRX_\xBCc�E�yc�Ei4��d���:�3_x(|=�<}��2,��J����(b��WIoPg��E�[��1��lX�p��}�Bg��؀	���+�D���]�����%�;R{���28�8��Xs~�2�z�Z�Z��R�	��ܷ�p�N��<�I7����t���P�{��/��`��'U�Fl!�$~���v�!���	����sad�qK�LA�:pX���}����f��xtZ�U9�m��W��WZ�
X�HK�zvV7����@SG����������W������}N�ф�,e���ve�*�	���
���{]��T$��UC�%�3�GA��XiQǣ�N�9ӡ�J�<�Ƒ�}�~�ɎSO�,�,3SUG�m��bsZ&̛�p:���g�B��=7�x'"�px�[�d0���\7��G��>��p����蓳-
�@�B'9��Q�7!HQ
��QZ��9<�˸r�.Bf�a�lƷi�����.�U�����T9H]�5Jd�鈠�c���:��֢��k%,���]�,��&螉ٔ"��ߍ��X<*��x'�;Dl2,}5���ZC�k�9�S�x��=b�i|�P^�i�Q� e��|p���GG�`�*�H?�����"y1�5��kL��_�6��AT��/N��'�;��×�jX>8�Q�Y�R�h����m((π����5�
���,��{��kY���z�p�_z��𐛉�Am�;�A�|�P�������y���;�v�_ط�&��-aY��~�yDi_�Jp���YO	]��o.sgћ�����X��d�XnU��j2����o�o�W�>fro����G��KW#�d�Ll�-[m0��4�gk..��ܷ,g˂��X��K���9aLR����M�OX�UX�L��mӮW1�T*�kNO��Y_��]�ݯ�#ݲ	�P{哻�B��r��
���p�Xc�D=�pfe�hT�ċ�3�N$%�i4�c�hg���Ô�'d!���3@V7�X����5\l��~�5�\8Q?Ya�7є�(���ޭ����o����rםMc]�P���@����Uh<5
�<*�Tv�*H3�+x��R1~!َf�)��	�[������NX�!.<����S�5#�]��ǰq HG��(ՠ%-FYќ���z�Q��&�dl�mf�*֨A(�wD�x��N�h�F"z(<�|�UC��|ɳ#k^�OYC��v�G��0�o�U�C֗X�e�k��� {�?&�db�z�>��|Z$HG�$y�oۏ��Fky�I�v�DU5t1R��,�o>fS�{3��#k2&�gZe$CA۪$��ܻ�9�v2Ї�}��j3�o/��.w����s��8� ?QD���#�Oi�y���~J=��:��|=�-sv�	��2�c�`�q���tv!s+�037t�.��A`�s�).��bc`����Rn�����-���d'\r!*B��}3^�l�g?����hꦤe(y�����pyl�5�Y��[ER��G�g���g��l�ۭz�4Fν?����!Z�;�M[�^��[���D�O��^��.|Lp0��)rqc���'��p3B��?��j( ���������WZ�{�{>,�q|qqxz��`���OC�l���iW�x�;�-*pK��˓ ��dP��r����
JYZ�=����*|Xܻq	�6��v�Z�k�+N�/�潽��Uj��3�A���3�
.�o�?6�M|�7`^ȤI�ɘ�+�w]��e�]5�� ��������5�NI}�֥�rC[�+>��l�DAqR�5�`S���]|t_@g�����*�
4Ia{LXV��P�.�BD�����U}9���@ڬG�E���"���8�3B�YpID��)ҩ�<M�9�a	*�A7:���E�b����N^���ĥ�6N��z��}R�i�7��d{��5�F��WQ�'T{0ak��g��Qp���ڇ ѣ׸�Z�kd������$����Y�a �(D6J�S����������y�C�B!)g��ܩVd��Ց2��9����yhQ����s�$�c)������J� �'"��d�&��vLr`8l����U�Z�u�?C�$��̖-{�"
����N�'|���G�P�q�w�Ĩ����9��"LZ��%ع��H��6h6KA���	�z�Q�O�b��1�>k��F��{u�[x���o��g#���94B%���W���hVћ�x���&
�x�c�{
�#N2N�5x�Y0a
K����#��{����d%H����D�]��VUT��u!��PsPl�����^�V�������)i�.*���,u�����f�4*�!9�����^����rD���j����r/X�8�#���3�S�)�����EBp�p�گ1�~���:S>A���_q6g�`�pxe�L#Q9V|�k��9�++ �AW��Y�P�w��lem�RX��P��[��������D	L3�ǯf5V�:tS�߄r9����TFEܣ'�ぞ��of^Ի��V6L�W&�7���e��Az�����M	�+(��.�B�ЄЄ����O��B|�hs+H%��j�zf�C˓���p7N��4��e�y��_�����%�w��k^E�y���2��.�N��0�fn�a>�N<�O���T^�P����z�>up=Ԩ��:�CRTh����kP��w��?'����E���@>�FsYN��o�^:F�P_Y�y�ĵiU��1Z����>�.H�����Y3~ִ�*��ޫb�>p��<F�a�/͜����3�t�M��dQy��&�&=	���X���y�0�PQ%sG;����������������� &Hy���X���^V��/(&T�D݋�q�p��Is�Q��/���Kb�|�#]�f�E��8�?w�i��RQ��Ӆ%]����(+��m���D��xM~ Dc�*KC�& rפ䜰��,<��+	2�N?2��^��!��~���ˋ ?��GE� A�-2��4Ϟ�d'D]*\����ݤ��Ǵ��)Zk�V�8/Z�}����,y��_ ;��7{��𫢛�|>���U�b�}�xM��c����o%�.l���~��̒�2`�B��c����$cw%%Sʚ�^/=����C�Y�=��zb��g��]G�Ct�+*�[΃�:�6�\��Yo���c�ڗΘ�-�lu>m�=v')<���e�UJ��p��}��y��+��s(+X�v�����f!(�ݺ�շhm.y33D�G��#\\1z�a����i��+�"��0q�1�*�ƪ��BGƳ|i�Q�Nq�-� C��#�|^zdK�2|���:�����
5��������1�Iߊ�����?��f��%�JH��<@��э�����H��Xr���.�d��ePA}������I%��E`��j�����t��V%"��a\�N�#��Vk�8~&Ϡ�b���n�I�U��d�oY2�:1?9_(q�zq_Yz��v�Gu�x7�i�S�Ì����X�F�41�/z��4:�P���SRG��ΟPr�ƮXq����E��M�厖g=���F����R��V�t.N��]��y�%�5ำX�@(�}R��[�N����%��`m�/�ao��	��H�~�:���blE��9���'{j���G�����|7tT���'�����<�`��D2n��}b�kkk���  ��m�Y�n9�pCI^=V1��|aê2�^���ܚF�с=oM�-s*	,z�J�n>�y�����ً����9���a�׀Ik82b�m��;�����J{�{0�̸�L��� w�B�S�߽�P�Ҷ�%����f�u;���>GF�r���:(���R��9�L:	{�YW7X���[��k��4��<�;{��0����>
fz�4���9S=~H7�? )�A��!gO.�p���D���a������m�
�7ȫ91L�[w�q�µ2<5k��k{���~^3�.@�
lxD���"\���3��Qxs���*�G�xyPd�5R	(��M�1pÈ")y�!�h�����]8���M�ϭ��-V���N�K1ё�|6�\�U�@` ����>�ko�K=�"�Vv��r�c���XofuD��}�R�=���Nk���=K���¼V"�/��k,{}��.S��݌F�r/��j��<�B��e��ć ��s��Ȭ�M_p��Q~7 �v+<�� �9��U&���`��=Lךyx��_����0Ğ��Ժ+��R�మڡM�6����U�w�F}G�����P��>{�M�6Pe�r��^�����6��s��cH+�t�]�3�e<"�x��h�.QB�<�_G�̾'Om�%?�;�N�Ln�m�5ޞ���Ӿ�W�ac֫���U�0 ��k����w'T8�@��"��tIs-�kU�� c� �Oos.r��w6W�GC�����Q�}G��'�jd��
�8�����Ѣv��Ho ���$@��c�@��=�ء�n��Rk-�n��~��ew���+j���`��]�W0����QI��d�{�J��e�$��
�i�׃�w��-���R�C6ѝM�kysf��lL�HX���AFyV݉���i/����A�eJ��Wߝ5�?�aӒhÔ���$2x��#���>\־�}̼��m����Jn�����m���o�8��@�տ~�/CmƝ?���Q���P�PX"�V|���ༀ[C�`q�q�C��.W��}�;�����~8/a�0ATqa ����N�"�w��y-o-����/�:�kq*
����Ii�b���"tAKweO���Gouå%g�ݰ������%Y�wY�K���H�MEx*AA���p�� WI?e�	��9��Ӭ�Wz�4_��Q�$x��p�ɦ��7b]��~�)��X:Ϡ�����p�eۛ���Qm�W~[�lIg�6��#zrV�s��M�e�2���0��1���X�7�����6N�R�U�2�ӡx����Y�![^B�B��v�^7ʂ/���;�:F���?�ʾ���'!0���~e]�Z��p{�\9ʤ��ɢ��.D
eN&��L��t��)p!�$% �<��x�l�1�:�B�+s�3p3*%7Iϱ���U[ �k7p�g�&P�r�M�4b���#�����՛	�q�2W��E��i�����{aS^r}�<9KU��FH���A��
�R����u�-L,ORKͨ�Qޜ[{�1B0�qv렜���!���V����v�٥��r4N����0�ux=p�޽���e*'uE������������h����:�i�[��rq����4_�(�D1��8����Swۻ_�Cv�G��<>�E8$d��_��jJ�vD� �֜���A)���h��~���F������K�\@qe"C]��5K��{�7%�(����A�_�"m;��	s8���!_�x&z�(����b%�k�Ib��y4��I{��$���U��̣G���,˨�C���Зg��CGf�f��-��d�,��/���h�I\���IY��>�]؃˅Q���6xS(rJ�_R���6%y
��E67�l�gY�ی,���ծ����	a��������X�"��D6��	n�lQ��X�w��.t��0چ�d�I�k�hFH�![�`R�����')�(c�)�o��njg�y�v��gh�:q���1�~Hy���^[��� 5sy<}_�IW.J��7l/\#�i�(:vUx�u���>��S1�f��3F��v~��y�͸s�#S�,���T�=���H	�� �������9��k.�[��ǷЋ�Y{}�3?t�EBZ۝�M�Pd+�u� �Of�� /��{�4!�u�V�H��x�e��9�����/S-;UV�ű;����n�sV@���G��Ҟ��Ɍ�J�4��3Z�C��/$?�f��B=<�ۑ�</�D�/��� 9�K��^{�e��j��!|����se5��� �$o\�������o#7[Y�]���6�5���U! R����r��}�H\��;�R����"J��w7���]n7.L���<��|����;��ck,͟��C�թ�3��<c��LK��>�$����̾LI2JV���:>�VB�l�+�/��~�G��g>cDV׮s=ٙ����[�/�Ef��HfQ��l�,}�Yq5���1-xb�~U�ق ?��.cI��� r�Y�Q�Q��G�ux 9�Y]|@�P_�"ikI��6F8>�r�s���u���QA"Fwi �cf�8��L�ކ��0qI�9�4\/�E�SV�U��f�JN��UA�Ą�x������dY��)�鳳�t鲯S&Ɩ���l�2�b<X�f�kX�:���Jl�4��+֏>����5���^H+��0B}}��[g ��j�,�,��:o��i`&<�n�ɦ���<F���%�&$Ʒ==�[ �%�,��(���Z�p".���z��ꤰ�F£þ��#�o?�T/�������,l�O�4d?V�.G+|�o�I�C�_ܒ7H����26C��Ne�����B=Gb�}��+�j�J��q��Zh�s$�}mW���-���>��R��Q�����SIo8GR�.�}�i��o����^֍@V��>�x4��t�J�$�"���M�_�P��?%�tO�o�i��@M7�?: �KX7� ��q5���W��AT<��2���i����b�f�������+>h�-H�zj��������Ż/��Ŏn��O���XmxU�X0�:ƐU,7�S����x:(��'���{O �c���ﾞf|ya�k��z��E�:�2��#��4'hp��K����q�J�j�C`#9\j�Xo��I�mP�Ԑ����hQ�zU)70�e�߀��[��of�9�#<s��a�����|���l��T�h)A���1yk�o�᝭۰
y/�,��bΕ�y��x~��҉U��~��_��2�F4فX��-�����`�;m6K SJ�$'<�Dٯ������*z��_�1d�#�w��U��UF�����V�_� 2��i�'�� �Q N���YɜBR�,$�<��ƅ�i���.{��j����n�#{��XEt\?�@pk�2�$T߉�E�ɶn�M�Fxuă��A�f �6�pc�q��O�S��э��O�r��&��6EMx��� F�F$e��#|�ߠ�M~+PD�R /�[R�53d�<��wN2�5�WY�� ��s�y��+�߭�^)/N�p�����1U鳽BP��*�}��y.΃��Ϧ�bWM�l�ARW#$t˝R� ���z�j�����c�rq�|��@�6d���|K	�{8*����Z��Mk��c�<�T /�2��#K�bR|�F���"hT���4Y���Al:T�Cx�I8D��J�I��c�S�$Zy����3ɗ��O�6���h��W^��QY�2)�X�j&�\R0=�켺�T<��`�碄�i��H
�sJ����lm]�\T�/7��v܈��hA}K1��*˼Hj�{���$TQT7w�� >�ӃW��h�|���!U�yDc�w��#�u{I���f �����7�B�
Hʳ�2��L��bGP�3�� 5�M���3��qVd�����;�5�T#�h֢%�bI�~�F����t	Q@�@��}<�$������Ջ���=���*�BףN������~���w��di;����:8ymKg*��X�bHҳnop���P�<z��"������Y�h�㚜Y\��İ��P-h�Pt�E�#�����"a��8��2�p��?��|=GUN������W�C��c�o|���",�ŧ�]Oʎ_�A�*O�\;���+[A�k��A�F�o�HNT��XE��LHLpS��&� ��a �H�S�����:7��$Y�!J�|y��~����R��L5�,g�նp.��F�U@	{S���o���i�?/r�e�Q(����b|��x�(�F���iJ;e�ۯ��dq褽Ŋk�Q�đ����c�]$] 8�?¥˄u���>E ���6��B�$�;�����r��8|1\Ƞ�����⬜� @;AT]��#
R�Of�T��Eò&��W"�ݭrMO>z]� P��-c� �M?O�3o/��qem��9�I���j�a~0bp��\�p��<U��n�.D�����V��ޯ&�;����"h��=�E��,)�M{z�ƏF���k�.��ھET��LL�t�n^����*V���$ĥ��ZoB�~z;1t����'�[�{�$yZ!��Eb����|;0�a�cC�B����V�U��O�:L�Ϻ���{R��(d<�עk\�rUީ�j��bX�Q짣��_�]��@PU[�� �Ҿ}�9���t���]ҭX�Ds�*^�]gsV��B=�փ������J�yL0�49:���}���X��Vhf�_��_l���4If���Z���ɻ���dc�F,��{`���0	K��������1U�<F[H��Sx:N�~�l�y�W��oCJ�K��O#;m�$���"��8�m U�v�e��ڛ��w��~�|�Z�ա��[[ �q�hhǘO�[C���� ״aA�Ȭ�q��A6!����o��"Z��q�Z�6]���B�D� lXF�Ui��BF�V���<�	vBVe�o̡&����,��Sf.愍m�S��S�w���[V�Q�K�X M`]2όqR[�!���1r6 �2r�-��tp����W?d"�%��Ā����*q�m4Dx�/lrB?��Ȍxw����d���73��}�|V!VC*��U��k��[�� �4&��-�s�䳉�cB�I6�r����C��g�x6	R�eP���ɑ$���f�L*��J��+ޟ��Q;��`�c'+��?*��gᇟ)�qu��{�{P���}%	���^��;@�3.��Ao�Ƀ�/,p˟K�*=�׳:�+)
Ɉg�@|�L�∛c��h�;C����\�	�x�w�B\6;@��l�$�����`t�8�����M�z �u���F
��y��M��p��rGVr|3ohr�\oȑV�H!u@1�������ȔI�霱�xU�8�Hx���%�C,@�0���뇝����0����*�w\���y�����>VUE�,"g��}h����T��5<S�f����ֿ�>UQ +��T�1 �̀��e�I"��$����d��*��\$c��l�kĖ��^��� �B����r�B���K]{5�J���R{z*����W������]�9�-�����3����t��O�+x��Z����K�az�ߦ�k�_��N�-|a!�~���p�z=3���"����O����qE|��Ք�J�uŽh��:��*����E��.7k��{)�%��6lX���l�3�Ы��Z�}i���d�DK�:�D��75@g�[9��][��F�M��,gv|��V�ܣ�����7��Z�E���	Թ����цr³�ӱ�?B5��_���@MT-��/�Ҩ(�e�%�v����t��:�n�{�,�u.lƪ��Fkt�Q�jPMDh�N֞�_	\m���Y�V/�iz�D=���uRn����Fs�'�hR��EӴ���>F Kz펛*$.�ϧv�����[V
ږ���ʼ�*�4Z㶁Gr���0��xW���A��kP�M��n*1R@X9F�ĘU�u���r��"����ޕ`�h�:A���7*Y���.͈�/�����U�9w	3,bV
#�����7u�'�Q�����U�y�&~Ծ�܀�9��	��g�s���W[q;��Y9�ƾ����)�F�Gm���;�9��.5<���n�QYY�99�׈�Ʊ�*.���L~t��vB�`Q5.������K\qI��Y�F�ׂ�yg8v��~�Uqz�D�7�ؤ�_/�í79���8�{�s��~�~%�ŉ+��s=mS�:��H�20�+�N�����>�@���oYv;�\4{K}��մ�&o��1i�ف�bGbqsO�?u�l�V�F��t���׵Z��m�6�$��;�g���2H��E���+e�PH�4��R�|0�S,eݧ|������Ǖ6O2���E�2����^��~���T4�+52�F�oU�b�^���#�?��5��ī��!�]����ozJ����g�b�f���	�#�c%��@`\�ƈ�_��{;O��\�_r�b�sitʴ���D}�kD�|�K"��.���Ԙ\PV&|'I�[���K���B|�	��[.ǳ����ۂ�Y�Gݻ�z��C�hWu�rix�]_?a�T�,��
:�͐�����$��'	?XF�l{��|���'��؊�~�!�m�cU
�Q�R�$�x����I��B���K�j�%oQ�T���;����k�/̖�Z�b� �'��d&H�M�e��H��KM�f���w����\�&PER6@3�,;�%%:�W�g54�ȧ�-h�~M���Ľ���e�>��#����ʴ�x��j�E�
����&�t�|Ѻ-�2:B')N�Ԣ�d���{G�Z��ËNi;A���=Vb�ڥh�;�e�o&�eQ[C�e��3�%�V��
�g���y���D��-f_ m��1���l�^�Shzj��/��HA�Q�/!�� ���ڇ�ۓY�����^�_�5���2]h������'�?�¶U�(RO��}M�8=ڧBt)H�.������Iy�{��d���@%[��H�ƺ���S!�]���	s�ƶ�����ߟP$�0w�Zɥ`X�&��t�E�j�˙�J�9Hg�(�!/�]_���9����6OKqŢ0_��Ȉr<}o���~zfJF�ֺ]�	�7�"�#ې���y���Q�u�V�f�	g�W>�շ5q�X{�N$4��;T��,��+,$��+KHJ�y���o��𙃤��L2n��z�m_^���ߏ���0��F�2=���jM��9k�K��?_���j@�A�e��8d낙4�������N^w9�L�wޢ�A� X�����Oʽzk��Xx^��G�S0�K��Bpw����n$>YZ�D5�2ǫXeWSa� st�ŏ耭S�h6��[�d_aJ����傘��ڣY�S^��՚_/����׹������ Z�L(p����8D2��][�%� ���>��7��'\2�@ՇZ���k��Y��Aс�~]m��@r�J� ��D�M��"��E)2�I 	0,}��G��Q�|�!��dJ.��oL
�L�xX�j�QZ��I> IZYV��t�;(��@�8��w���&�c�B�^�~F�/Z��P֕����%��"�b^�"��м{tG�����֊���F�y~�髃=��U`�"�$3J���\�'���1s��
��#�*�2�S���B��ނ�8q=P��b�T�~C;��~g�i�����v4٦0f�w�dob��H��e�-I�t0��g��/{��9����*;���b�C\�kd�Z�����ҒNv,�**B���M�cvٲ�
��l��j3ۙe����-&�4w�����8ܕ(�Z�˰�g�>�9 �L%EC��ݱv�Zj%MU<�Io�X��﬍c޶��idx'{���]� �����o�H}³����F����g �b�0#"|H�n`�����-��=ӹN�����}���6����K~�$��
/8ߏ�<�U��	���H�ݿz$Q&�&�j_uð�F�� ��LI�!�u�2��t�l �JJ��S���(�TJ0�}E�����mh���ba���� eesO!S%9�,�E;�����������
f��}w�㯮���@���Lf*�/X��~��1�+B���M�ɟ�ikh@��7��9s*q�]��0�6��*5��=Z��m$�"鲈�*�~�|>�G�{����)`O�ِk����~R�{I�������SB�4?ۏ��z�y���dNY��]>%k0thd���7T���gH�nl>����Ehjz����	E �CF>=i��7�B����Ί��t�m���C����џ��y ��Cߖ�p��h\���|\���L�i��]�&��[�䕟������`���t�㦰�#ǓC��/�L�ʦ6����?���|������4����++}R�Q��o�$�o�s ��ݡdd�c(�H�i-������,�kw���B��B�j֥��($W����<J��6��dfs�D�*Cd��k���j^���@�gr2ޗ��X7.M�N��X1/E����\oz����.�Uep
>���XC�l ��]�Ȁ��;X��v�4�q����b�C�5rv�j�i����4\���vAӰa`��h2�'�TP�s-Mu�e�9ҙ�j+TV�rUϗe�=���K�i�nz�p$֧��o$�~�M�}D��^��]a���dg���K^Ў/ޫ"�_?���(a����S|�z�.�ˌ`�'�����3dr��_I�"lgW\>^=��ܯ��D7w��\�~s/VM���f�r(9�?�S�AuϺ�`��~�R7l����SA)��1��v���� �rLn&I�����f9��?���R�JL{�,�}�2�"�2E��|ՙ��wi��m�����U���a����D�Ζ����X���vS���rG*r�U���_���~���x���Ê����](BWxqt��?}j2x;����Y��/L�Z(�'�˄���w�ӽaO�+����X��=����}�a����h���g-IbN�3cx��z�@a�Zz��~���	�H�r��O�5��Ҍ[�!ʕ��]p�^�;���=�g˼&l�#���fq�e�%r���x"����Hm�r�8ħ�V_z\>���D�Yݐ�䚉�<E�B�2�07�(�EJU�B�������|T,��������9|����JÙ��=1�w���M)�R��eK�Fi<��?ZP�l_l�p>�0Z����2� v���b���JF��Z�L���Ǻ�y�N�GՉٸ~x��g �X�+��9�/��F�{g]f��/�!ݏ7��Z/���߈=��|�Ҫ���U�^��������1�����@��U�����$PĠ>�Q�	q=��Ų6nQ!�.!�A{�Rؿ��T���?��~J����)�";���GP/��[+���%�������U�ڔ�|��kFI�xkf٣g3S�}� �)_C`<]L�-��W�\�b8� �&��"3��P��UqE�#�jvf�u�/z٪���7���ս]���o�Oq����V������l���f�~�2�(�]����Kr�C�j���v�yJ�< O��N`��>�A�s��/���L?��/�<x�2�Z����ǆ�,���cbC2+������PH���
˽�v5�i5��}����aJe�M�,<��h:ԢGځ����#��cЊ��%8��<����#΍�Y�Uk�O��|�(�z�7�p�F�l�-�R���IvM2*!G�}�9�&3b�����ֹ���6&�c1���٦M]L6J��%&Y����o.�	�E��щ���T,F's��c��_�&��Z�B:�h$�kP?�a��I�Mf�ʓj^{�5~�_��iI���0: )�e�,f�+�Ble�>�\b1yI-���]�����]� Q��%���,?p�Dq����#2�`~R�����i��XA(�Wyx:VEp}ē������!��T�r@�ɔ7����w�K��'TI�_`����<���P��>&�P7}�����'�+X�p!\�9Q��X�v�a�g<�iАN��I7!(���>"��c�}-&�c��be6M��p>��E��={� �X*/r˻s��?a���Fʗ��pm���'2�����.W��+c�+ 7Z��L�����n%Th�e��_C~Ձd�ˋwZ�2C\�?�w��lݍ�d�S��k$��2IH7�]I��I]6Wkd3�`k��M�8�O���N���[�����չ��X�7V4rb���q@&耱.W���!Fw{B�Uɚ��p��I+��Lw��K��%��e�VV7��$B3x�D�k�"���H��� ���W�,��2~Yq/β@(����gz۱{ɳ)r��慭�fxٳ�7��)�h����[�z��g�%+���vy<Ћ����j�v�Ӣ�M����UfM	��v�J�w����	p�@��In��U`���?u���%v_�0�A�V$��8I�����p]'Vk�B�r���):���QΪ@J�>1�6�� 7�
���k�`��Ѧ�3a�w�[���<���W+/��x�b(�8;�_k��d�l���Sh#�]�zh�*D�zvs`�����Y��=���aRJJ2c]U!�$�_��k���MXEF���=�h��1t��I�Ya��/�Gq3Q�v]�&k�� Y{,�D|��8OşHc���.^�z�+�L��_ʯxh`��;�Of�$��������?�I��y��hF���L�E���M��b2���Q6�o�@��m�w�{#Ld	{��b��<Q��p�}7V^��P˨��i���B��b�BL�ӈ�i<Mb[��%R�s�w:�Q��J��S��X�|���YmH�&�ȎmUh\6u�Y��rg�5���z�w����z	����2��n�~OVY!%\&����6��He1���u�H��lE�����̚�����#k>:# �iD���s=�9ɣ&�(�����L��ݏT:�R8yu*��P��D/���z�8��A�X�3����ti(Ó˕�?��uO^�}(�Ը4Їr)��|��ػ�~�oD�CBYiB����6"0��5�a��HZ���?3�b��z6Tip�09�quc��_�$���WDS�}A����A�k�n)lCL�;����LZFk��Q9m���|�����>j Y�`)(������q��Tf��u���d˛x�������?K�o�l�}��av(��r����۲���C�>&�*��h_=��&��>�b 8��	�E�������
FT�(��n��!��},/�������)<m��-�8���k��=;ov�'�S���pd*�s�)7�j���[1_@�� '&>�"���v��P�親���-��VH�f5�<G$�rƊ
��l2C�_ɘíg�|�F%�kq�:�Í}����c��J�,t_�/Ӂ���[��lYϯ`��Ɣ�.��q��ʓ�#�S��� �v��L�n�X�L�b��yw�4�X��)����7W`�pQ�[~���O��HBfYCV�q��d3Sb+��'7��~�.my,!��~�a��¦YP���=`6�wLU�����m�#o�ҹ�\�Y�z,����	�Qqĝ��[艌�����v��7P��t�t�ka��Wk�U�4�����5ga%��"Iq�	�i �l��;d�+< ��{�ޤ`��Xs5�=(u��.V����r����cOÖ1 ͅi�.���5*� Oo?M��f�I|�A
DF����[9�Ċx�pj���*�>����P�v�I;�D͆��r��k�QQtN�`]�L)���`%q&T�ҙ��P;��Y�M��T�<͈(I1%r�5
�M���,eCX|�,��Yԥ|��C��#���֎{�RyG����gP�w�\��[��ׄ|v}J0�A�c�I�����
,{R8��oB`#c�C�t�c�CJG���N�"	[���;�o�)�f�f����H��&:5ͽ$�tS�Q���
0Kea�  �踓�=��>3a�����9o�+���l�|z���ƘHZ�1`Q��?�ม�bIf�T���MZf�4s(�rE�"9�4�W�]��{�x9���m��n�4���aJ�2�s	��V�W�?�7�3Q�E��M���ӕ�{t<�o����׶8�L�^�ē�`o�����,ժ��l��f�>�[���gxz�h�0m�ԓ�]BW�z���E8�X���/}{`ߜ�����K�7���zf)�m4��9����.�G���r��^I�(��mg�;��7���
RE�6=�����1��NDn����24��ҹ�=�= 7�|��P`��ve	�<��߶+V����a'�s�'�ʝr��1 ����-�ٿ/��c43��ϮGa8T��I��K���?���bi��#�n�*O"�ˌ<։�
!|[��k��|P��+�y�Tg�|A�+زK86��JpP� �J��O�`pY~&�qa%�I�l��WG.�=]�n�ʭ.*��d"q� ��E� ���:ɸ��Os��F�����l �<�` h���5�A�1]��G{:�n��������Z���� �y��9��1h��!c�n���H觭��U����O�P���2c<pIo���=�mQ���2���d��\`;��o��C����N���%W�KV�tLx�ŋϬ�V�����IN�x��)m��A%䈀4I�(*�p٨���6�-څ@��=�)��>�j��\��pŀl��������łB����u
�[cТ�,Fa��E�B ֘��o@]q,����z�����;�$Ѿ�u�4Z�Wճe�]@*q6:SNsTs����LǕD�r���i�YH&3��q�9Y�+������%����� ��;:�d��v�(`>�l$�V�3C��������<'�r��9.�C'�jmg��&���+_��@���M�Mԓ�l�D}����"T��LsA�����x7c[Tz��ݘ_ӏu"�y����ٝ�ǲA1%1I� �Ș^p�@���kH�:�/mLPT�e�M��?g���]]xT����}�p������ ��2"��QM:~����Y~����S}�yK�6�
n�!+���Ĉ|<�	J�d�+����+x ���
k�Ǹ�cK$h�����ۧ3$A�*[R�� ϭӟZ@e��@��)(vn�N��R��P<����&U K�+XϠ����0��E�KŌ�28�[f��Z#�_ʙ�+��X��V�9c�̂i+J��WحҬH�[�a�ڮd����"�.��j���Ο.D�X��g@*J��oGW�yC.;�U5����H!f�v���A#9����ױ�!)
��\T�G&���`���𓎖��B?�����T�����!���;o�D�1��qp�>�j������E��|������d<�Q���Iߒ��w��ϻ���̘�Ը�cq��\+s&�"�5ȁ}�[f]��+��J�_���ٞ���=!-?<O�o���7��9MGW3&�P�giO��+��Z��k��1u}�M�mC^2���O��J� ǰM+���ǫ���)O��J�<J��b�B���_����Q5#K}^���ߖ�k3�G�:dY>��&�4�υ!�U�(hϛ�)�^zH�Җu�k��c���C����}d�y!.[0��=��6�x�����{FM5����j�����Ao9��OR�[.=��E�8�m1�\�{c�W��i�(��\��㜭P����&��X|�E��Tm`�tUe��
)(+2��g}�Ǒ�m�p���������3��_Rr�%)[A�*g>_�`������(�(�n9Q�e��]96�*v�y ���˸��f�$�E�Y*�ޛ~�I< �w#���:��$5ѕ����e�cD�L�,>v�fC<�=���(Y$!4h�G��� �J������_��w��k͛Ei01|�ru�KBF��`q��;�b'"Z�����L� ";m�<Ϸ/'�z?�isʄ�q���\�:����<��.�"t3�5�bg��]u8����đ��heq	�䡬&�5[7	Ћ������?gS�Xz��@�p��G��s�8F����nK��*��U�h�&Bs���t�Pg���5R̕�6�=��\�����!�#��+G���J�ϋ����XP
#�,~((�k�UQzD��Q��O�'Y�Lk�������;�j����ʈ6�h�r����W�mmό�_#?�s�Y*�:l�"z�-�t������k;�r�8� ����rJ*f�,Y��\Op�iN�D5O�x�"U:/��r\��*/�K�tz�)�� P����,�3D<Ƶ_t�3���F�a��R߇�Ŭ$�M�v��h2yK�%o��N4�7�Ljۘ�
�`�3�ᠸ��2B_a�������U�h������9Kc�%n'���S��F��O �_�q`P��+  ��v������r��yZ}��\�G�����2*�R`��AE=������_���\�MƜ�!�O�{ە��-�-d�w�,[̂�"�zl�3RV]�,6ZRsŪ\���v{���i�'��i��*� ��uu���?!78[2�gVf���e�wU�j�F�̐�w�#�:�\`� 'Y�v�M���M�@�v�j �����A�<�M��l��3Pʸ]b1�����l}*��}£��2f޷�)��7ߏS"��o���h�UBX@b�)��}�)|>,�N�QQ�79x]�Ļ�|t��x�m�𡻰�.tZS,@�� �M�/���>��DI�0��N&h�C5��$���_�'~�OwI)�SB���9@/s�JPW��#F%iն y�͒F�&�Õ+�i_� �y�ȘD��Z��ƣ�׽i��?�Iw�,	`�'�d��v�����$!gYI��!g��D��H*���J��qKAR��� �E����:,fh�k�xՠw��"��\L��D�;��{��� f�!k�xR�{"Z��~�A�*7q��E��|�����
SE�v~�4@lJُ=�i!]���g��A�1*�E5��A�O{���P?T��i�R�E�h�DP�ȷ�@�)�+&uu=I�p	�Q�kU�؂՜�,kN��_[sj�`샎�AMH���ܔ>={^a�Zf���P[��z�c�L�jVv�>�3@�-|�'5��rq��
C��b�X��%�ɻd
�0-����z{r���3�Ē����a�����"�.M��y��u�*?Pdw� 쪧�x����	�P��HQCd��w�%pYʔ��������f���v)!�
Ȇ�m;����'+;�T��JX���M����Pm$�զ ����O �AR[�7�0����B�s��=�]b�������z����w
���2:�@V���Hƺ�`}�� ���y ��3Z4qt���T��~�%�+M����}�8bE�k�f���%s[��c�+��h��3��=�XD�e_�Q����Lp�L��d�Κ���A85�_�r����h��婉$�"|;�&I�v�0��Ud�+��Q���8'�����ǂ��j*Ss�$�P��2����0��v(dl� l"`��r����z^�N�A���^}.w�㬞0��(jQ��&=>	��,��l��sg'��Vh�H?�y�&���,T�{��������b��?*�T�e���@���U��F�}?#���3g��[�y-	-}���uw���Z��d^��:m�X��H���s^�l�����I�{?e{x���������`0���4i�hau�^qʇ�^, C�j|�P��BUd������j�֮�{3��1b~r��m�N{�k��E]�(�p�����ƶ�e���'���2��-��=%���]��Ѧs�b�������ʞ���}�H�4�ݿ���� �G�E6�e�����<���s[�cO��eĀ����X�o����P�#F�۵e�R����CAG�	�ZO����I�)>���Z�Q�4�_)��o��)� ^��R��zj���t��*.�|A���1�y,2ew�F(�;t����\Qg�9��Q���(%9���U�<B|�1G������2X�һ���i��4N�a�)�Z%�k��Xz���FV�F�ĭ#f����D��q��.��?�HZ�0�U�i�3�r�ԧ��+���
�s7�N	��NPE��o��I��ǭ��'TG���϶J�� �x�K�p���п��������e��li��J۠K5ہ�q�}2�+IU��j�O�]a%�z�-U�u�|�>�)�=�:�q���٭�O�)�y}YQ�s��
;�9����$��L��g|�W�����ݚ3,z��,��v(�8U��5S��� ��"��q�Ge._���)��>��rQ���>ޠ�/����O���+�v�Ʒ�k>J���3���''������G���
!YM���*K�X�E$3���5=2?���'�) &P���{��& ���I�s�*n�J_��:D}�r��䈐~�j�˪}çiA�+� }�Բ7�H��l�p��¯	���6��v�X�N�"1�t��ra�~�� VyĄ.4V��A�����UZ�8�5�<�
Bf�[$j��M�K�i�o���� x�jq�J/e��q}z�O+cTM�M#$1v�F��,[�w�S@�$�h���U��׶��p�j�-��&��qk�
̃yw}�_���(}�ibRe㣦/\�2�Ɖ�uTM��.xXn`ᛐ��F�.�� ���	#?�3dVo��PIU�|�d��2�>}k���>�ƍO�S�BV�A��Wpf���/�!J��]��IZ���y��C�G��P���w[ x�,�!l�3�l��ƽ�a�� ���\X=">���E����pSN(z5�o�&|�T������f}�����
0��/�ݜ���;�c�00�E�AX�|��
�,Q�!��F���l
)��T������JtQ�����F ��Ie/d�n���~��ߩ.b�*i}���81ۻ��cR �����@��1�����O�5
��7��ӜJa��C����E-T��W��sO1�ā`o�OT�"-*<ih,Gp�Pz��и���`e-����#,�B���˜�
|�.\j�O��TМTz�@p�V�tt0�,�bg^w�3�ܮ�_��r&��žs�o��%�q��pe��J6%���.��ߪݪ4���]}.���T?��J�p�o؜x9�vO�FU�;������prǛ�,I�@�[�'�"Ox�  ����X��EnVH8q�����8�5�4��zmT��%K���� ���$F�#e�}K(��`M� ܥ�#�o�d��U�;e�����[����F	�xK��u@Py�r�ohp^�6��ۥ$�K��}|��RI=�0��6�(���l܈�FPϸ�K���x(�)����'FҪ_9Gk�<!��\a��C�I�W��n�(%��?q��>x�����S�zOܤ�pZ�\d
�E����2�����{������7��o�j�kv(Y�Z�a��+	�|J�e��g\��b����d�T���?��iEV"W/�!�J1No�YCU��Ob1B4lM���G�����S�jØjh7��-�>_'/E��^��̷,��p??�쵗JsԪ"�����5�foUw�P�t|���"�툨��e��ȳI��}wg_P�I�WF�-��(pa ��$��8�	�0x֔e�]	�Cc�����q����΁�i�(qb�V��5�w�u��N_fTL���»���s��d@;>���1Md*\�[9|�s�T�/�F ��m�X��R&�
���b��l-�~�Akn�ϏJ��;(�h��x �2 �
��k����ּ�9P����鶃�4L�&��y�d���	��c��\�c�M~���kY"���G��h�/K�X��#�ꌻ<Wy�<��P��l����θzj��4�[��3U�}�l7�@=�}ND`�f�d�Hxꅓ�vFH'!���0/���5F��~���֥���D�3}k8� :q�!]�G�D	@;�9GEg�̢ew�*���ίz:
<cΨ����,](�e	���̞�RPa��t�e���e��?��F���"=��{ř_��4t����+�)�:�01�/�r��t�[��p�dB
?WfE�&�q����Ѽ̰��݉9�%9"�2�E�S&�ޘj�e3�o��O$:+>��Eqy�A1:��^r�)c��oC^�����Rs�ظ
?/�{�Dt4�g�)�(������!��I}���A�c?��nTp܀2PR��1d��-��ȸ7���=Z�b�[�S#7��j�/}��fX��B%F��Yt�Xz���c*�{�Y��u�O/��9�[&�`�w���帤���.S�����W�����S=5����0^��[
�%"���#tV0��/E�*�p��>�?[%�<Pԡ��2���������L�T�Y$8Y�6�SRǻi@[�@��©RP�e�N~)(�UZ�cu�JZ?K����JE����r���؆x�9@E�4 Q�"4������\�qT={j�nX{.!��[&4�M��ر������6~S�R�a^��#\�0]قI��7�"a�|x�`�纩V�	7����+���q��/v ����
��&sd� �u�7���Si+Z
χIMT'�f����2P�=�5�6��y	rx26{i�W�U�9�I2��Ag�{R�v|{�)��A���e}��4�J/��A�!/-��U@����v�˔����;������� ��
��fwDջ0,�p�̪&~�s�J=�d	����?~p8Y�eU�I�>�0U�� �NK�U���q��w��I]7 -'>BP��@Q�рIC>����C�� [lK�f�������u>2%��!����5��G���H�H��A(t�BX�[��ˇ��л�A<{�v!V�����5fw���y�ft~7yuUzg�Xw�L͋�b/��O��P���Ў[E! ���K,W&[�Ox�
����o&v=�g3ԉSes�M��7G��A1q\����(dj�0".�E�Y%�F����'���NO/ �m��Y>
�i�lM�]ظ�܉t"�a}=ɒO��5j�B�Z��z���:X[���Tk8�n��j\���r�� �ܱȬ�_A�se��1���WG��_\��C*����(�����'/�5�??�ڪ�㗉CӐ�R:}��^�9�!]`f��ݯ�	k��.����y.��f��&j��w(��Az��q��n4��S�f�dO���P'�   sUpƖ�/ ��ª1b�����@��2���Y��#?�F��"��4k�ӈo��$#L,EK�:\�(�H(��� =�%K��ZL�p.l���>�T1��a�B�	nl�S��E�����p����U3Ye3l,]�Z��I�_��v$��9�������p,�ڂ��{C��p���R�c��㍃��y��F`/�N�K�pȨ	�ȋV�"M)�[� $	Q�7��9D��u�*�����>�W裛�"EY���p��`��Ȯ�7�+w���P�V����÷�=�F�q��0}�7lUk.l�����1ݸ��·C��ϣ��,U%=�uXY_	�^	�m���nWw=ji�U,���,eI����������m��ǣ�r�Ό2th���e���H�`|�/HO�#��#	��v���a�c��GT���UӶ�?'?x��~5����&�1�'�WL����6Y�w�(*a�b|h�H��&����i$F��e5Bb�Ui�ʽz���6��e�[�o �{6'+]�D���W�K��	�U"�դC&Z����zT�ٺ�f�����*{+����#C���^� ��Ƌ��Lޙ�ڢ���T��������\H��`C���3��/ab�k����� �z���\��~u [�;��`�S=:��9m��1�.X�rN���岀uqے�+^���:h�&4u;Y��:����=�Ug�d�a���yW����ۙ�����A����p?��S��._H�D��������G��a�j����ܩ�O���x�6����SےYye�s=���s�Bq����'>Q·�j^�����qG��6���J{�.?��Us�:U�E>�%�=�����r�X��'`6I�i�ҶsW�!�J�87�
��Z�h0M���uU(����<v:�i���s(럱��$���h�<jB$	�hi�t\�_
>���tٵ��������u�bŧ����.���|�$c��_�-j;��}wȔQ}�q�hY�֩R����5�$�+�1�d�ԧwV���J�S��Ҽcr�yc<�]ٚ3q͒��fM~n��t�y�f�I3�Smf� Z���#+`E�t<jU�"d�����A�����������'}H �k�+ �A<J)��^�aNg�g�w�A��ߒ%���}l�n��H��؟�|s�w���2�E�x[B�g��s�;;(��f,��DxdH�Pc�q�,;��^�˩�X�M�E�Y�?�̭��x��ˁ� `���8Ť	�I���-�]���x/�*�y�^�O����*C��P�;q�Z:sd�U��{����k#�����Y�GnP7ݪӹ���������P��K��.+?���Љ���蓝r��A���S����k��"�U�~���Oh*���5��ss�C����k��c�%?Ȼu3���w9G�X#��Y��bb)�֯�r����:����碌i:�Ogb�� o���o�P���w����F������Ps�����6|1�#�"Z�:�C�$'���>�$��+��ݺw��5E��+o��zh�ꁜ� �1s�/S�G	��B\��_1�-|j��,�Ha��o�Q��iTXJ���V`C�w�e~��J�Sʪ-�g�\Iݔ��oa�f��c,-L�{�:�$��0�).ad���q�d7ax>��E�1-�z�@�۰+ZԸB-��r�Ku��r8SH�\.��w}#�I%l��W��ez�TMs��Alۜp�Dʋ�s�w���؟�ڳ�%[ß�E�����̢��ZJQ�=IER�3%��GWQ@Nw+�S��'����첏)�ְ��b-�PF|�k�c-���$�o�dE�l�2|�G�Uݥ�Z�'^[�4a�{��}�!���l3�J��?��q��vF���	��F�]��\�(�CF0􂃍������b3H}�e�NC��xW+�����v��w6H)���U�f�Ez!��.K9�d에Q�]�l�@ �g�_r#)I�ւ��^*�9¹nʴ�2ܸ`D����	���L��Km�AO��%٦���qe����(�9��.i�]Ў��3瞸�v��8�߀k�k��!����d5�9)�DD,�{�S֕!�S��qG��vëh/�.l!)�G���z���)�g�.Eȅw�����.+	5�&�����#b=�.v�~�P��'������7+�� Z�s��/� ��N����w'�x��0h��S��2y��)�r���4~��p�;�权 ݟ�(����@��_�cEMu���g�X��A�]���'|b-.� �������bh('�x��7�+������L�@�����kqx��zX��cY�c%�8# =.^yp>���7�����!�eW!l�Sw�q�d��$�3 �K��j�iM�ɠ���$���O�,Ip��Q�
*�_t J(t���Gi���L��=�P�������}���W҃{��޴O�J���
��X:�G�GD�\���T���ݼ�J�-%Ѧ��7�L�2�r8���X���J�N���S�IVRD�X��!r˔���#�ղe�O�ut��{:�@VC���3��@#10�hδ�� όA� j"��*�N󺯚��_�K�1�x=�QO�[|;(���Ll�Ð!�8���W�/��l��J,>
��e���	)��C���Z���dg���+�a-J���5[��Z����D�"  ڬH���k^�^��i?Рm$�p�$�K0���3�|�ŋ b;�=����2�����B�!��C^���/��a�ɇ�8C��=V.$~���e�8yi$y�:�,"!Q�t�So��o`�D�?��0�5E�A�h���i?�Mb��/�y�ַ�gsoӕ<\p��]j�h�}�Dl�-v��'Be'�mr!����c0��^3�(T3WWai�y��ͦ_hAIε�r"��$֯�PDUh.������qL���fͣ�����q�e��`G�x���"Q-���,�N;!�}�B���xN���<z!	�����	���KD�qy��8B@���fI��j���S�l��	d69 �Gg6�#�W�ծ��?�,�n�F�:��+��?�`��t�9a�N���#�U���IKe``�����k�S![&������]I�	�ghM��})y�ТV�yXψ��b� o,C��e�*��?B�쒀h��TEs����A�xk�_�g׌q�D�ٴo<B��7���ܯ�d�3�nĭ�MO��a��\.�2�tWtIN�2��f���ז���4����!��F���~�Ì�jhvaGH�^D��tSʧ��,��s�Vr)�0���A�3{�(s!W�O��eYɋ�B������x��t�����kt�-\��ْmGH�?��8��W��/��+��9�D����J��s�,M[��"walf��hgD���b��*?E�^dXg�X�0AhJO��o�tm
if���8U�S��������+���{��PI��'�zl�����2������X�`���I�)bX� ���R��}�cz��8�{)�ꨠJ��@��!(s�j������A@?��^�1B�������׆W�$F^0�T��U��-nu��c�%f�UWٙ�u��O5��0H�k�/����]X��Ý)OAK~ ·H	�D�r[���VΒϰ}1}����_�B�������e���Q!��g�"+�	e;��Z�� ���(�0q/�)����'�Z�q�r}އ���a&?va|�.e��(�&�B��:#�����S]�?wea���� `��B:�S.g�
��"�l`G�(�[8^�\�n�T���r�ʭc��gc�&�Ku؝#8Į��.o�P2���E�9R�Vr�?/)XS��� ^58\p}!�	Qs��;�q�\�3�X��6�< XH��ޗ<@#TgU7�N ��S(1����{��P7���gy�ͅo��v����4�!�Ŗ8�P3�dQr%T*I�p��ڨ���G�l��HivL���r;2}*j�1 M��R�������&�k��9��BY�u=?��O��m�����k 7�l�����d�;�U!�p�y�G+R�1�zn���_oH�&��͗]�SW5�����epR��C_��x���	mÊ'K�㥦���@^��G�":1�Q�:ہ�`C:��11�rC�"�U���v)�b�j���RW�g� �Y�R'=���%�]�����#�?Y,��1;�E]W�!��"W��"��:����qQ@����R����j�y"���&g��$R=�]I&��V�<�&�i������ �ɷ���rP�I�����>��х�ğ����@O>���F�{�b%���B�7j�c��a6�{��}���1J\)^��=��4�'�騛�و/+| ��+�j`����_������ٺO��^�u<�=��*ڱ3����T3S�9y���D7���#�a�E�Au��"�.��Q����y������r�ǡ���n�!Z�]ccbN�������X��Z��L��v�d���(52J!�z�Z�}�������tV�{5�g�Kp���\�gY_S$�>�$ڗ�����%��0aK�OT��RT��F�(��Z�6�G�g��0��B&�>.�ѷt�?����Y4�xn�8 �=��4��{���>s,�R:[ ��[ԡ�@,��	��5

������D���?�6��Js߯��ʗ�i���BG�z�<S���5܄�u嚵�Ew;���ؓ��ۀ��Þ#F��q��2�*T�׸LM��b�����՜�ƏFf�Y!�78��Q�\�{<���Lq�j�U�^�b�Ҩ 6���/ȓ{��7�($lw)ŕ&�٣GG������g8��P#+�{z� �6�t����d��F���QX� :�M!KF��� �`v�Ig^]����x}��sv_�^�W�עf �K�Pw����Q����|#�$�G��Q��M���m��ޓ�n��&�~3e�d�8Zp�vW�N~X�Y{�7�#V��sa�Ul��e�wՕ�O]�Gv����<�N����_�ă��b�Q�M<��{>r�7P&L���+s�q�<O�E֔wB�3�M'�r��i5b��G���:C4�m�Z4��6��.�n�B+��8�!2�-���]]xQyrf}���N0�:�2c�t����=��������,�/r���v'�˖�~�UH<�l��V!�&�~��ʎp�=q�6�}�iH�&�6i���j��Ƣm6~1L�ҟA��M����3�uE���K�M �#l�(��K����P�=�8,$��o�%z���,�Ou���̺F�Q�Z��_L��;��:�,��x5,��
���-���qUz�G1����i�ܵ�L|u�t����x��$�!j,ʃ�w{��R]r��4F^1꜊,b��l1<1��]~(p�*VIv�$�����x�d�r��h�0�i�:0��P��ٞ���AE��9.�䤖S�2p-����[�E�(ə�8�N�XY��-�ڔ�&e��)��i��*x1��eX
���J�6����P[�c�s8��m�~�:�2&�p(�/ִ�To�wT�k�3E���q���Y��'���\R9�t��ۗ���:�� �C
����Un@����v������T�ñw�h��d�������%���.~-���&��>���i]DL�6�S5��ձ�G	,�n�#Z}����Ų�D���\*�27�����;糆��j�:"�ucu-��{��ض �\�AO�R�����{cQ�����}Wo���ԧ쪜Bn�+� �#��H��]v�7�-��<�;`2'�����p7�e�� �&�q��Ķ�bg�.��_+k͠���i�{e3�a�[@B���Z�U*�`�&�8G�=tU��r
�;d�s���A2���#!��w�\�сP�;��X�"���hPG����2�L��ʆhi5���)O�[V���N�&�t�ZGJ,���k��h� �3˪&��`iNp$�5�[	󐼗��w"�M�rۇ�,C=��Oi��U��Y�� E����/O�r����M��]�m����rO���(�7�XQl��f��,�7�w��0��)b�A���M�ғ���vH�1���"��N�	d�����ea���{Yu�� 6��=�9��-.�>I]̋�Aé�K�m|x/�D�-��"�X�(-�T&�O�Ԩ;6�PXH��pW�C}|D�f��<y��E
O�BH����w.��^II;���B�ɼ^��i�;�c�3]rJ�g���Җ��*9��� ���,̍wf�*����)��a��ݠ�fd�J�#�b�����K%R�¬�����ٞ�s��R�9#�7�n�	 A��F���s����V�	��ī��H�x�ivwd��c��5b!\�@�����5&;S���S�8+�p�qI����9i��l��\,MÞ4��Y6�q#��O�J�V�1k>jf"��P�ϩ�4����1U�K:��Z����Kk����ͣ#�A��K+�Ip��n�{&K4 �A��!�$@�Z���O/�+���5����a�!�v����G�� _���u�A� RW���+�G@ê��������[<��\����i���}�Y�Ĺ�����,��a��`1o*�kE-��`=�Nd��pS�he��@}҄` ����0�1�	L?��
��(�_��hR��G������H)���)�7�y'(��w$�x8�w�"N��\�o��ęY�>��V��%S�sV�a�e�'g���8����
���^mĘ?��`��k�!H~y��mO���>>u�p��f*\/ǫdP�aM�x[\��2x�n���������(���N���u�`�5�[~ ��.X������͎]%�ц��/�5t��_��6���O ͑��������M����8?6ԳP�9"�t�c���['�3�����
{�zN��ƺ{�{tnE~A[��ir�4���/�4C�S�.� �f�/�L[Ԩ<�!G�AB9���ү���x4O$� sKl�����al�AR[@"�V�¯�p�0�?P�(:H�������IeF�-�f�)���ҒC9gk(�2�x�Y�m����̆:��m�g��hr�	oZw9����ktd`O��e��Ve�8m���o���ᱹt�dNy� �r�n#����Z���=�ĉW��u�y]ϗܢY�;��+jq�,G8%wI$�B�L[nG���8���j��O�RgH2l��Զt�����c��[$��F�E�ZT��pr�M\2�M��.�陼/�X��:����gY���_����Ώ�6�,��?��:� �:EW޺Y2�2��.h����Pm7A��g��f{yH"�v�4K�)[A�,�RA�w�|c;ȵ�����3��-4�7�ܢ,AHI�`�9 ������7<3��-�9s��x�p&����vN�z!����!�$3��y�G%}�x\x�<j��Z��tyIY�a��K�P�5~���{���`�Q�e�ҙHs՛� ��|Т����qbhʠ8(���T�yO������_jψ���i%Kd��Eo�j�{!NՔ2N��a]���s�Z9�ֿ�T/H[�^�ߜ\43�3#-�����2"o����}|��Ը:�/_��³Wq@����,�ur�_��-S�V���HL��l��+gKs'=�F-�]d*���1�h>���F��]z�-[��Z.��ڢf}��3��M ���AO��i�.G4�;6O'� 82�(��L����\# ٸ�ḳ����?+���X�3sr��J�(�Y%�߱5WǤ��V�sHC�v��${`�[�zჷG����et
ao<��!��ǗyMw�>�����;�>�J=//�Z�Kr���
I���XГ�,4S%Q�^�W���-�ć��W�N��������1�j���(���ޞK�Hj������0�E�񤉄��0�v�U"�k�R�^(-��{� Ai�P��G�zN�`��\r�W��֬������ʿ[��k#^���}�2���Rn�
̚��eڃf�q:���k=^U B�[�D�GG�^���T���{xX���،Ĵ�<1ky�������w�w�y~�i��<��m��'a�5�F���l�^���!��vc,�޷\>4!�
�U,l
��K��/N�=NcW�O�y�HT��!���]��%�`K � h5��8��3�ȪED��J���<�+1T�)��L"Q��R�����E�/gZ9�r�p�����<�$�JB7^ RU�Q�
#Kb��f	�6�c�R����N�DPzTE�������Ժ� �+�U�\�Kc��{�t�K�X��A"\�-lXbf��E��X/Z� N 7�s�j���:&��!�ʭ/���~U�6UO���w�
�8�}��=<x畅�b's7�����jb����4�t��Ӣ[���L�Y�#�)np{y�{ġ���{��X�����>d�����\�ɺ�xB/	`�������vQ���,��T�������y�}�i�i���q$?���6��n	f�#����<c���MV�$�����&�%�<��>��j@Y�MB�s��,�2J�N�D��;C'��In�o0��jo�zВ���>�v��\���cc}�����F���B+e��_�%k�#���z��"�!sE�p�d�*�f� iD��<��V�].g�����jB(-3?�/��Z͛{q���mf�o���ŸS�,��CE�be��,'���~H0!R3�%�R�A�-�8�f-4�)�����Q��y�֬�������-˰���:>vS�?��OF,f~����9q��i7��N�)'Elr���s�I!��~��W�H"t`�Z+��'_b�n���Ԁ���/87�&�@��(35h˨�,��(�!�i�[n�����[D����e]%҈�oÖOx2dc��b�Կ��� �Gc}9��%�	gT4kFe��݃�dM��anăB�[ݶ���::��z��ǽ�:�z ��6aIV�?�櫬��
�� ]�T�dy(!����"��$%��J�$쇑v|z�'=tk�j*-w�N�>��~��d �#�/�/ȶbjBY���/sD7���6y�a��������]֖��[�C@B3�f����u���v0pƕ��`ЧQH���w.�j4)BI:��yeǻ!������0Y�VpJ�k�h�|�N�&�_n�C#�msjy
������>XC%�N��?�n�=�/j�L����p")�-�Q1�yXu�F^���^hq�6*H�6u���ww`e�9\��8�d��̩�d{S�1��M���HݑQ��f7��_ZK|�h���|f^�8���v���t��b�Ǳo�jM3Y����B��Sw7�
@��(B�í���,\Agq�0���g޿93Y�]��xg	[�G��?*�Qˣ�Ό�tl�ov��kv-+��ǻ���2-�g�aC��Cx�^,��h L�4v@�=X����ru��R�@ّ����;<�kţ}+�����e�<@��f�M۴��]z���z.G�iϏ���MCq8܊I��)�X��;0��'�O���S�*ĳ��N����#~{
�j�7?�F��G
0�ݨ����b��D4��2i�l�����9��iߜa�+֙��^R��_섦9��T$�~Z�11��r4�����r�&Hq�$:�3�M���W�p*�]�fp�~6�v�I�sx��&��
/�L.l�� &`s0��z�w��&���X��ڪ�Ctޕ��繾�@�[P~�~�$�Ƽc���rq��ur���3����sn*�4�摿�᫴�D���'$%��8&T]�؜��E@�����9N�&Vp�ZKg/���N��%�ݱ*�30�q	�k�n����-��a�H�/�<�e�h���b�[�
م���(����dk̻�r��	��s��e}K�-���|�q9%,��}-�kmJ��Qd�(l��%i�S	k��	6����䳑_��+#j�3�'��=���K�n����TAe���5k�{*I��~�Ny��c���⵱�f�b/��+�O~_T���M}��9�G$��u�-���R� ]�5��������so���Q�C��i�ͅV�O�&B��>�����P���IMH�I������(,mM��Ҷ^�����G��о�3F�1\rÎ�X���������C�v�m���A�U?�!xhl�]\�dN~e"�Gc��b^���&x�3�E�m�yHgrJ�z��DӢ�e����댝E�4`�-%�V��D���j�ŔR6?�NӺ����
I�������K?V!2��,�v &9!d��A�cxy �p5ZM��P�{?MO��zu��F��K>��m�<ͼ@2W@^y���������is
�ѥ�nq��T��$�1=1�bP1�l�%�ÝFpE��ǈ��5���E�m���i��{�elh�>(��P�9Rx�w�$e���hW	pI��4�H�a�2��FH/�f���!�	_���2�:$� ����N�.q(_*��
rE�d�5�ޔ�_����:�n�rC�7W�)3�{$+��_Cm̞a�ey����Bd�5%��j��m�L�{q�V/�{W��}��6��;A���T9E4_��2`���v���,' �3��:���9��;T��ݣ=�>������P��.2� �%���ؤU�3ܰt[|
���R)漊J��S儰^#$b����c�v~�;<�X�#�K�v�h�҈o�:�#�,�Ă�z�����G����R<��Q��Ao��[F��hW�����(�Sk䍰�E�;����97=�Qq�Y#���b���*�:$!|�L.T��\y�O2�ݥ�传a���8aDRhY��I]���7�S<N�����͟��`��t�]n��_��c��9RL�cΊ������`�A�CH���^���4��NB\������o��@n�E���a�l�D4����zlq�>x�|%�2�6��6w��3Bi��#r*�D0N��
��~���P��m�*]���;jaC�6���n�Ul�����+h�T�yt�|�Ҙ��U)��r?a�+M��\ҟ���n�3}S?(Ȋ��U�G��e�n<a@���ڊ������u���^�F�J��!?��G~��!X��9�G�|s�21G�M^��=r�է�CV�����5�L�����x���I8_[V5���/D�&��N^�TKzc��eH�ãz��n��B#~ܸ��<Qz|��?�0^�E��Hx"����DM����C8�;��ą"$�\�$�H"�d�7�e�pe-�Ǳ����*�Q�n=��7wI����XT�]��C����#��`��UȳZt2��:qZ�3��������Z� jS��������}\�N�xj$�{����s���<��Mr^�Ici��p@��p���["@ig���]�6�4���[Q���������T�*7��+�N�JnW�c�I�T`�����aG��m��P��EB���a�ʲ�X�WA��,�w�\�/��ʭ�vc%�Tx)c�4�b��`6&��a�Z��UH��έ\��YWA*������\�n|���r�mW����ڱ{U�w�w�,�d��\pi	�H��,|�c" ���&�p`5c�=����o��Ӄ�r:.�_>Α��F���.��� ��h��ޡ!}�+�ןd��VcGF�|���5��Ql1l�x#��9P@n��z��*8�C���7�貸%���Ji;��D<�2�و����V�5V$�=;�цN;���|�� W�:���f/��,hv%Bm#����v2e/��;t"�q�@�S�Dn9(���<ޖM(��q�Y�G��&�Y~��+��.%����qǦ��K�f��|(Qc띕I��o(��i��>Jf��G7!��G=���?\gmCf�i�X��C�m� =R���0tc�"��9�+���F�9���S�1�f&R���.�m� �5���"Y݌�]�/jN�S@��q�UF��7�Ψ����C�Yn�̰Px: +z����P!h�sr�� ��vR�}��aKR$�a�8�x�F��s}@����B�Ʌ�/��7k{?�8$��R/%W)?ta��px*;����N�
��'Y���|��~�@�f��~�{Q��RB1W��-�&���B������/�G��߭d�N��nG��NIa�9݌d;��R>�>��e�i�)w��	�n�]C^��[a��37��[eH���TnU0]�����T�/�q#�">K��d��\~�������
��F/�6�ZޡU~�:�S+n9����n0c��p#�l�ʨ�*=�!@�F(�����)y$�Q|F~cˏ�5�W�7���&�_DwӔ,&US�/c�(t���;L�\�+��$[4�"�E7=�3�P��era7�w	2xh�$9�دh���s{`�@9Ap� �����Ɓ�����σ��W���r��D�u��;c��>���jW)/X���l���.%}��%��L��<~��u�^�skln��B�l���Msʢ��C����8}8HF[����CT�� �:�ECr�(K	9 ~�}�h�����f��hM�X`���W�$�rpo������*NL~���]�L�d2��g~��`�z�Mݳt.�V�0�?�g��7nq�]�1�����'����dD�'=\	�9d���b�,��\��A�W����5OC�n��çVW��n&	�.�zJ���w?�
�#2#��Abc��,;+���H�B�Z�o �_=s]�E���.=�E�}<��F�ʣ9?(��-0�8:��Z����4Z>�G�H��D�==�:]�EYp�=�y1�K�'7���$�E��n�?2�ā�E؞�!�l�񸇊���Sܻd���a����<$(ѳ����n�+A�=���^��vF�P&7������?V���<�;R%�1��骍a��mӯΈ�)�޽�yG�=8��Ea�א'��~إF]��HS���?�{rAn�~.��G���*GAǮ�l�}�%��?�TBQ��( Ѽ,wX#Z������ϫl���,cf�����ƺ�8h\�i���o���"#�أ��`(D��3��6s��Y���(��3~�`�ǀ݈���?��ǈ>a,O�{[^�O愮!�8/hN��.`�Z!<�?��p�*��)g��-�ɢ�G�4.���2%Ȩ�t�U���B��]�#(��!q��lX�/ҁ��Z�X��PD�T���.�g��(-Z,�i|�>?'I�܃���5�	,IP��6�o9�z����Z�8��d��_�Rۤ�����d�h�_aF����f\���A&�T�r^y&�F]��Ж-U��\�$����@	� �W�r���,@��'܌��J�s���� ������]��y�,�$�8^eM�����Z��ww���U&i�x��+�f�ф���g��5_b���x$b|{j
�W}��K�d����to �5T�]��C���Ղp& CRg�k>�ZH�\>3����O�:]��$
U�gK\j6S�y�zL;_f#+�_�z=T�J�͝��z�Mδ$^�CQQ�Hp�Ow��F��k�W�eE�&�/ *V]x�t&5�x�}�Ĝ�9f��b�"���¿ᄭ�ӷ�w=,��Rw8Zh����"e�� {�ďL��t�C9�!��j�E���:�+8Z�E��M3�g�@�qW�N�l4�ȝ^|�46���sR�O �Y]�G�/�,��=�8��'�[*�m�h-fj�l�@m�Z��=8��(y���-8�$��q���#ƛ75��⤰hS��`Ù������O:HV�M���E�W"N��'+�%˟[۴ge�m��s�0��v�~i����7E�� �0}����L��xo����cZ��d�\!��/�(x�H�e�1\���m��=(��y��Z`;�`�y-[�d+�i�"�u�e��]���t���0�~=1�#��_��훾"HQ(�}#j5�ό2.��mDd ��.Z"�Џ<��`�.�A�D�u�auA��eQ�o�|�����=��frdG՚��(���~L_$��G|�kZ︺���pK�X�M�7�Pid�׆�MF���7�rF�zڠU������</���G'I(Δ�6�1WBbL'_�=l�cI&k(B-�4�-]�j��$� ǣU;�/;-o�����%����_�tq�<s,7�.K5WcYHoK	Y�%DZ^#��ַ�}�'a���9ȔC��SK�:G\����)���� ��&�S��)�9�f�@�$1�*��~�c����[/�>r�-��T�=޵�
fI���R�dD�H{p�!AҰ�f�;m��n��)P��!U�m�Ԫ�����q�)��a�Ё��9[nD�n\�E W=D��s���1f�=�����?�>jx�8<��K0:�C%nP8~����[�+JʜR��Ё>��s����~�k�l:X|��&�М�:�W;�EAj��I�_m�]�����.��{lwe�T����ت�qu���DY05��~]�!�Yx$��?b΅L�NgKd72l�9 �
K61D�[�.�e!���c,�?ؑ�jk¨����\�� ���b;���KO&bA�q�; rn�O<�{T�c�o0�或l��1�Y�S�O�t�
�fg	1�X;j�qY���݌�h�Tr�Mֈ^�ecѡk�f�Wb�8~�W(Q���U�y�y0rzu�i�kd C-ҟq��xX�6�"��7��'��������xts�
v}���,V5�G)�bWW���ӗ�4�^���)��L���ߵu+#0z�B���j�l1<I���H^�>d(���F-�D�-�	7���vc-E��zfvr��we8���4��o=&x�,�-IG�0��x����?l[�r�I�������k�ݸ�7�0���F�
��@�w���@�u��i�kY��7G��u�vh��"��R
��Q��dz�@�����_2�����,i�"����x�z��3�{ڀ�	2T��3 �@�V݈IJvS��5�Qf?uq���T�j4k��/����;=��v��>��2N��-Y{���"�1�^�=<�\���L醙��Y6�y�U5ΓQ�u�܏Y��ty��|]҂�����뙀;q�7�p�)�*����8R���;�$��+-O�d}_��EE�,A�VY�+��u�! �eZ�e�Nr�iS��1�Թf��=���I���[nG�B�|5�S�?�g�8�L(���/�,H���������NN�ˎmW?[��b(*�=91岕�����m��En5H?�C���_�G>4��]��@x��&��	2-���1O����`��f쑡���P���<_<_�m��?拓��а~a�q�D+7C�q}]-<��p|o��@�h��<&�J�ݭ8l,���=�ˎb�,㶠q&��Fr����hDq�.���r�Pn_I�H���|3�:ԥ�-�kџ9�Rr"chsG���ۨV^O�6��%��W�����q�_T�Ó�� ��Bx�r��0,�0.=Y�Q�k\��;@�ˡV���Z.�H�꾟+�r0���ho�!���{��K��)�Q�H^����a�-��k}ؙ
� 3��1�<i"�z��`O M0�m���n����lz��7��hk�L�!ڤO�Th�y���& [��G"Ou���gQ�^m��^�W�TU���D�Vj�$�p�p��� ��<����))z|��3�'����-<����Pų�ڸe�Q�QG��"s��_c? �\��&c�g����ס�S�ZJfXt~o"`@����e
Y�V�"�6�����V��e��i�PH�������-w�(����S~�]�/(�R
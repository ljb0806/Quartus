-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nFDiSVnA7RDpzXgWQRI0pZyDuBeJdYO/OPQ7rmaSwEGIdiMNkK+Tl2xD5gZCvRoZ86ovw2gjJbEQ
zWG43BiA5GQ2+yDHJsS0KoDD0mksgkke64H7C9EdtkxfOt9OYpjYvoEpJbdr/7Za2USoBL52NH5E
i3fof9961fjhPUmvyxH3VMFLCV/YXjNJ9JvWJ9IyOPSMGDDXTcCqZRvzumjACoTnthITd8xa670D
jJVaJ60qi3MFaUGkbJQv+yGfihTh7+4RDNvXO07sIdTjKzJRZNnp8LSt6ei5gf4w09Zl9YT5r76a
lk7IbqPj+qD6b9Zu1KhBDH+1RLdbqYYIjrVcPA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12960)
`protect data_block
ovkWPM7t1D6ITG3Vh6O5VbzVLbGKgEekOZNzzo2kFeJHWxOVx5w8mHdEpUWwJTmMDhmnQi6jnqHR
BVw2puEN267cpC1azoBgAZssZJf8yx5Sdh2v3boI0m2hEw9OjhQSRyjqfCQBpcdv/4sDt2JsZuOO
qO5FNJAIb7l0dYaXft5jODlAu/D1N1Yhu+IYv7SzKZ+GIbJMElSOaGcwnaPeLnF//w3wCAvF4KNM
uxYHAz3lqtWcLdjRVwqzDJE7prbyMUXcJ8M7/ZiSb3TIjNIDtRBwBh9y06gNrVAyPxXEs5XNok9C
VbHobH5Bux5nSbiDOC8QrRGKU+kUilu5YLZT9GhUSOwCZ0Ti91KpfA8oH3Xb0rd7gBn+kYW0rJZL
kCY20s5eMEp2+xiNf1XBcPfapJ++wO/hcSnqaor61KvDkvHnVomlnl/2JJoxEBmYN/WJzsw+iU+2
DhwnEibvohle5qhB67sQxx19HdYTeBgfVtAf3Z8b3LMlts8pQb2oOrhbFrJtsMRtYOZ2V14RqWok
vh7ep+pn9OSiYmtjph67Amxflg5ZjDPNFnLVoqvdkXI6roEYdEnBxXqaR7rKgOoPlXmV2uHOn9KA
sP3j+uNwYvUN6mGdXIP/dX1fPRGN2N8/xQ4epVty4wbbWhVL5LM4bJmtoqyWyNQXYRysIOkGq7C+
jUbM/P6kWN2lOt2KPcLm/iv0ra1329hXczFCUr8THwWNOnK1BT22kI/v7x+4Frt025NSxCFCSYuc
nVBc1qg3v1SSGevjxB2/TZDDgYnd/Wg4L4hZgNt130GcQ0whXSLSfAjLIU/e+mkNsHDUd7FY4uIl
9BskwZTZwLKT66SF5OZaF0I9BTSSiU9nEEKA2v9+KWuQPDT3jPUpLQX0JVoVebQW/ef8l7YIfq+O
FX+QfMck2wJ++o0XZ+BsN+poiSV4B7CQdrn9hbyA/fqf3eCDJqt1AyzFiBU6gTza2oH/spBTYJ2V
NiLZj70gjfvfMW0UXbhraPbxaW8O6poUvhSJwTWUznTFpT6VqImTJIfSt9cghwJKENQBOOno+TA2
ClJv89gK+Gpv62I+DvFQC8eiG45n8gxAOid/JaI+tEHD9XCDSMfLG87Ilc4zhXEgyi/l9NBT2dY7
OxUOYQYW7fZHDoOoLVsSyKz5fMV10u3DSLg3wn3szHyELo026eC4gYTlFCKEtyaPW8IYulz0gGp8
Gw2btdT+wc6rZF9PHz+MMR85yFWcspEm5Eac4HnIgekY2M+Ve6Enq2IycyhCkF6JV1brICk6Rvdv
ODkahHwnlSc3YhLzhJzAYO8FfsJj/DUwCjVi7G1lK+SnSiYmvhnoLRAwy/mvHNQxhrF7U4GDijD5
QNHznthefZONssRqJ5SFNkepolt6ISG8gkWReNgumkHldILgT1JN6X7B6mAgf8Dqr60epQgN01vU
042VF4isl9eL7uazQscwgpaXpkuXAkJMgQIa8ISazdaM6MTUfuWt2o4k7lyAiJQOKaCr4MKm5zR3
AykhaTDaMwNVfZVGgvGpNhzBzRASbdPq0mAR8CPwzLm1jS7NOrZQP2PX4hIHgLOkcv3MuU4sE/39
YIH5Coc4YvfYlUNggvMNykmKYXV9gBhUXh6jSMZOe9oHFkV57opKek/ZPFumjCUqFnhx4C+mLYrX
kPgYvOOGfGuB8ZfxsnKRvauh18kRSs+hWqqseAGD6/V/tsoHal2CUBd7fU7SdEcqPDAmzVEMvuVu
c4nEOZW9TfSvVEI1zxpViyEDbuJ7jGWpnFvWZgHeP9O46H6imrTLTEapSPryk/RnoHewSS9FS/v2
Yzhod5Z04O7Fkxj/HUsnc74wqu/Q2ewWH+s6MFs8SXgetnD3u2x68jgEuXT4Vy9OawZGq3tFGHju
akISjfQKTHPIlOOXaKOWaKMiDBUzdmv5ehOKhsLw9/ueR+ESmlRjYrRVNSoVt3htQ7bGyNwcej7p
ty75sqX4vZ0qXPicrvA2gLH9NOHaQ6bVrw4RxIi42u3vWw+o8XGXaNA8syKRZ71/kIeWVmQjYeQs
YbGZ/8RBfdretqXRq4hmrZPwxYIN1c3ExErob5SnE6ZBM8Ch1OZZO1e8DeLBnjvbo97V6c8F9xHw
N//blZBzahjQFOLwXiWURhumBb2/RNWmvFL8jstdT1gG3EwHIZokaPg+skqKtoVa3tNmCXKN6/jx
Bx4cHboJL9xdz9lj39yTQkLOgYiSDsT42/AbTdDbuXn/954xhuB/3RNUs8kYDhH64cknNXXnG+ov
8SbXdQm7r1iaIX6rKA6num8eiKiaGv1CPMjiME36jPDRuqZbxxQEX4FA/tSzNFxp931pktS8Gsxj
CLG7zBO2RUz+kBA0tC1wEQKSh4L/FN+a2YypiMogEzWnJQCNlsWkyHQmNo6cAeG1oGwZLT0/7x4u
4nhU251HLYV2HpkBP1Ymo71r7J2c2GIF6JRXlmorAJxXLqOwk9/uFznqJriNWiBCnW21h+WvvY9G
nKph+eoPKeTwRpNXM1sKBkwCo7G3AWIaSJOdTtB8DgVbZ9NuN3YYqLZiCGu7CLHlSel0RCi2AyJi
g8PWxPzfmNsTKOJ01rdytXpDVIjKSr2XlWXCoGfQo2aOERSWss/2BoufYsSGhtd8jL47IniPqFr6
xgmLMVp2cwkGiEXP1Pn/x976LlbB3JCeALIGX4DHq8sUBN3WTgjyAvUN/xE1CIW/fQ6A0aGH+48q
S9okNXmYaEP8UPriKrOmCvSo6QWTllC+pi7pBvo9K+5oNmn1JCyeItvArZnDlvRJtdayU+mfmUtS
oj4HURzkUra1qwVEnp7h6udvQVCe8FgSlfj94O9ud0F414ft15T37ejp7Pm/HJgvkrhco91+esBn
FVL7UOEyizbxmmplWeVHpYtyPbaK5sM/YfcdqXw1HyGwomVuEIg9DCd468qFoKOsWBN2xEMotxl/
Onx1PKUWrumFIFjewJHnQZK12bQx8euWUdTyQJqEVsDd8jI/dEDoXPOHtxJzpjn5Jas9PnuxUByT
4ijafTh1KrJui3pmYCAslBwn4KGhkNtQFgF3HlorTB+cFmtNE5wudaIGzP/prgW/QmvCw7nmbOSm
DwbbysjbHpJkaw3HDYE/9FrDV25U7rJtNrvatUA+pDORVZlaaoKOc1fV8xZ6iAp5bVsItlt4BY1h
wGQNKfIrHHVXudBAFqQC5jeQ+3o14Er+Bc2O6EyJgrpvh7gkIFS8YBOnchovYJs5vdK8agEgsOJK
EzdoOE4/f6QpX55GR6+VWeE+U3KPgXU6eR6gM4sxuVloWWEr9+Hr25vDsug0sdKduErnRygpxgIV
vj5RWYJH6Oja0jFC0OwbomAiPVDrNkUDOQteJ40cTCtz+MY61qJQYlJKlXRZIqX2k55IkkLLswah
pTJsYg5p308Gxn16QvoURpFpOBPgXQccS4T2OOU9Um7g6MokYtqJbNTj4GgFPG39tbhXOTgk5fP4
jsVjVIO87Emhjb07vXZ3ozKsQdppM7BagS84CueM7HoUTLJZuZWeywuKYmkNleCb6lcF0HSuUKbZ
tPephU9Cs4ygmukp9H9v1qQpdukeEc/j65+KbEmkBeS6ijFQgyAZte5ESdikGN96RPC8JM2ZhB0Q
iQmniiMJc50FRMoIPksBT9W6aDOggn5cR98JSXeJ3wx/WPKH1s5YvBWzxfaDLnN9lDKAR4wmq3uV
npjgfuy98uA2X5lxflk8vuhaTyv8CpWZ0H+pu/GTC6fsaEGd/SHrzlZeKzD1M9AOLQXEa2sM06Xc
/p8JavvQTb8kuyEmXjpk66PoZpUjhMMC3OsKxRFaex3gGS6Uv1Nu9ehoMbsmuzycOYzcbZqdn5Qi
j2TZLe1mFFhxP4QrLxDU7HXd2/80r8ed66qPf4SGfQ/HOm1mcok+kPfdoBJylKfizEl0szTCmMGC
584lYL+53ZipkEhLCyeVyCL5FquJbhW42V9OTvAgaGnWFEr3LFa1QCaSGQJI2weihCXRftKWrQ+o
7dyDMGIYBAra15aHtKdlHv80Ka9df6FQxvnqqX3i9j8/e1UScVGHMWPJA+6+s+/kazXej7Jc76jJ
zw2E+tIPlw465dePPRrYESgGzpH/Kkd2nNwwWuyOhmvnj1wKW5hZ1N/9a9lI67NxF7AjdXdNzFWX
pAvsgZqWtv6KyiYf7E+1uWsaKDkJjs356NVB5zE+/1ePV9wc0CTRQB+pXMHZS/UX4jAWAwnxo5PR
SiaPdHpPQ/Vp5CZtS4tmvIwvYaG9JPUhuTCeoiTKwhbgBxkWP6qP0k1OEYLBsFzERYS6b6gD+eHJ
Ltw5KSMOibVRYJVA3FeMFSH0NmMyW6tNiEKpu3jfimhFCVNNmNKnom1ziOwYA3YBAVwNMYPzjSTS
2jCJodZ/n9rE4HokgZj6DZsmW3sDt32PxbpHk/tYb63pRgVpaaZfyAAr3kPmkvIblXow/VeGu/Zw
VAQezpG3d1QM1d8+kUWVi6E6lxMYMwdBbqCj9wXHg2Kqa3B5Q096Jduvs6cSSz7mCYYkvCXEFKs7
ou5F7dEeAMNAXbvlGnodzK05JigD8YZxzvWQp2ero1nI4BRDFcE9sr2PMM6xY9PCfAqb4bZ32Dmm
u+pKmXAjzat6tnpOYBOePdMzxPvmNDKPI2Wq19Crfxe4pdtCnq9r97PKHHiW1leVGZjeh5wULwsG
U4cJ5mfY1FqrMkgSUaC8u1/WRdH2CM0djnX+Tci+QhwC6YFytOZtp0TQ8aHettdQ1uzMvkS5pYT7
n3eeFKMJ4/uIhE6Z+31cQOyr5XzWQtXVAkXh4NG2z7CVFZO3rV3tqv2C5ndyMFILcvfQuT2J0ZZG
I3yA41s2pR8DQcnxUVYp9XWiPeDjn/bF4M6Xt8ishVlxJeTdkpMFgJHOXV6xtNBjRv2EqwK5z2yK
1rQVuGjto5Gswtu7qO6kyRsbPHdRf8L9zf6Kl505FnDwnmkzvmkU4s2YzvS4vzZSDZNt2mE5U2Zh
FxHR6gmBQAOmnsDtCjKj7ixFX1BgZO7fMUcpn4dbnAbtvcWW9hn6myt74ErY6L7dkZjITdfcmGiQ
Kf+jHJr3DFSyCbvDS/gBowq1DnpFMY4+X+J36SX6dPQB4mehcOhxNTT7v4Ux4TSb3rqaKpVOi3FI
L6i633ihLpxMZoSQ0DKj0FrQQzSQeVS1areaLHwD+KMXCWYe0suM7BVi5ov3+kj3W38sAl2IqHlg
EbBYe/idUL6g9ndHyqbbOzjNYtPrajmmJriHq6IYKLj2KU+ZJbknrzmvGKFCG60got1TuswQYHky
INLLYWNCj3SSPY9fBavD897iqF3aiUkvD/TDX9F0ghoHRu39T3sqmMB98IUR01nZc4k5r1Yass9y
Cnopyh1S5drzgkfec7kPI375qU5xODCdNO9a1oabeKqkkWPR2GvFPQ22SDQ6H6s3cdR7cFUgc+Ri
CQEX7CL/Baq/L2sMb21hOyBYNIBBuRAyT5oj7ntYZzYQ0e11mtGRwKDKUmgAlsiMwHXsmSv90SW4
sl4vNzDv/9vHNKJCHCdKbsvEb17upM1sN2mIM6qqXeoh3W4JvFRQX/kN8E2IrjxMQPt6jceSanGi
DMJ2CdckWcMPPF0sJvKJVc164a4/X4fK5a9TZIQxfo3An2KFqLOKW54sFMqAsW7BkpQsitodP9uy
3SedMffMrOau6aXsMIE7k0LpBl0X8s9pnxmgqAuIEV/A2731FyDLWxWvwVMBROlokvMISmzeEids
kdIYbjs7/sPAVF4yqpej9GvhWFt1K0+I5VFwhcy6v+E8w+aXTJfvXXu8sSEVdGZUGX4n45J4wazT
nsqzGso1TbRmo8//nLHeyFYKT/dCCqdQdorNVwhoDD1JVVzgifVfOntAYrVU967eaF532QR6lBVc
7PU0r3j0wCWVazwrrlCaqtkxPZyJGroTZoeygFLdSDrveAxZAVVTFUJjApv1wXDTS8sLxjMFj8GN
8L7XDoMcPspwq27cYaVMO9ZrEULKJzYzew2Hb5HskNorrmdlINbPOjCJM0KzHEGiEej4GBu1Ol+u
xkiLjA9t+SeRzJpZSsER26DRh7b/0XuUwLIN1rRkqV62C3fBKvTiHCkw13c+A3dj9V4F63nwc4E8
mY1UY81XjOZMS5lXzHLJjelaJZ3S+ZnUhrwrNng85TGTehflKp+ZuPYfgxUs5GwjMmoi3kZY4LRW
2VdrAJsJO+eSBuqGFxGJeuzZ7UOcifoYeFF+W+wKDtZhYd+q4xmjacsWeWlc80sw/s4XOa05UyGH
RYKQrNJ0uKloKhHB/xQI2G4bXOM2MLAlqpAgSkwqnDFIabVtDgGEmlujM8vtiA/jiKT30YSh60q7
5uSRTl2hO6uNYQi2UNBC41CTA3v8DmLAVZmH1ejiakDlrUvH8gyl8MHsXgWOR1I+V38yVX1z3JyU
MO9F0N6LTapqL6RunyUkv73MRArRudSfeWom/u3uOH46pq6vxJzirOD7JzeMYnBT1VDP3XtW36nU
3oC3rWOtGE5QIICdZHTEyeR8IVN9RyiVNGaVVIlnFd0HbZqeFeD20WeAucJRjUcR8uKlHP51zRp0
1hREAjzlQPnYtJ2W/3r3FGH0ckeRfpdXdal2eKGap0jC7gtTHEviqoGIYV3506X3+EXdqxIImdA0
9rQyRDc0ZbvsxnJWHA3A/c+bAZv1jI3Sp7O4yFWk188vMG6MmaAY2SpRgsvUJ8H4L2FaUKrILctB
WwYkGXiv9dUfDxhHBcLX2qh9kIah78V4JUwWYnB07EMnQmPjoeZwfQ/ZvPCDUfDceCPGtteMdSrg
d0KyAeLUH3odwGsgPQnCweTCu+dSksGpkwEkqfwHQWbFBOMBZm7bPbCXxB6cFGN4e2SdfdOFvMwM
lubtHKly7AKAsx1iBPhtvv25aV2Yf/JsEDzeTcivKDCsqw03fobwLZulj8Q3SqrDHknn8utIrHO0
fjSy2ms8ahNRF+lqxcmmzPrk4HYhwln+O2zj0ZvM6J7ITo9HwLtY94hJh+pOknOJyoRWh8UcaS2F
z3N5obZ1MrXsk5RZ4riuGri5SWiWCDZZ1JLT3rewWtiVXavXbp1zNLnZjAV0N2c/IuPgrN6S9eBd
93+bC3vCRIi599dAXXeMRXyG7QVADVxne5LCN+wFWp7RadJxkgoNWn0hOhP60Bs+sAE6jYsJOYA7
x3izhHAUjcoLnFydXUMTq+ztFjMSgy/vKhipZUM5WQ7kH1IZhDd6dPy5CpCDFj6DvZUo8sg1VI/w
dh2pInWXD6+usewr1K4au46LeW8G4C/H6ILUVDLBq/2Wa42lqfGaeQbO4O+5lTMuqI0lOXvxv50A
dCd5DL04f8uxIEKHadfMzlAK4Fe7fOROnOeCf6WFNjF8sxGP6e3GiQSudCdTNyyBfJndM8HV0tGa
RoCFltourb+3G+HR1DdL31B75H9z0fI/s2r3J1riYwOJz1gbVVqVbs9dq99YKv+vwR2lA6NqOzmX
TgMZq6oepPZJzVJT2pVjFIdIA7n4r5zohUs0pJCQUhSt1PVIcaA4kJZh2lLbQyx5jovtivsD9zbb
Q3wv86RVVjSO8Tl/39Zi1LKxM//qCMhpoQL+SQl1GOy7G8+z/hXX7fy79LkSgy4EPl7AVULX7uvN
58l5vewNgazkFm/8EnLliP70TCuCd+XvnsCd0pMZQtLBKXVRtNLu52M5xZkgvQlGf2MWG+nCIEvU
6AcLD9n24WS2DZyZCNGVYfkxR/n2ogrOI08xwB8jwPFN45Vjd4T5aY8VfOr7aNtc5GzqUz2QQDPK
mSlLt8qX30VRYYF7EcjzQ/3rYbD2ym6sczOBUztL4wP3hU9eEKSzcvPwGAlF3CNQnrjx47lyjzNf
5nRDuuoYeclxLo0epTEirldVd+z2dgA4MjT2cxsbsnarsu95oWS9kahT06kO5G70qjh9yAYzdUq+
IJvRkaHVox7xVLY/3DdO3fAkBJYe3vwpZm4hQqcaXWP0anPZCpZ8yDy/jyn3bgCYv8dSoGO1M1Wv
sjz7ZnoTVlfKCE5PHpTVs/6tnpNvHM/mYwp+fphbM0VCvPtkSSn0Klo/aBGRAfqR53BH4EyuQu5J
uekhulBbU6fa8c1ZgkrPxBnazgaISNIfRuk5bnyoI27BPdXbrG2TrhR/NN6Pabp+gI86JRug9LCU
ghLIPS/KhgwVNxlUi+YJxxnBlv9ocZFjg+0TU7gFIIo8xjiACYT7h/yXrODJJLtIWolTIVOo70qe
Un+Dk3qvBaiMIroQQ8LL6q0S+WkbCu3GHn+y55g78U242XbsdtnaBJNWIezSk8NaCUSUYsGnx3cZ
IBJgtOxXkupI2ETOtITAeei2Uy1bOSkY3tSvc03YwnpJiiT+qmDJBJ5HzWxUYYgEpbWaV45EmISu
NbAMiONREg7poFBs0VnO+i2FEiZnDqjaeqXXkSYLdHgKXl0/stjFOl/kdADMrYq5iPxCOe4YSuE5
o1ObJ9bMJ+Gyp4C12WLNqts2GpV2Od+3VR9F1fdYUpkZ6pcg7KsH8Tgwo0E0A+WZVtHAmGc0Hsis
pZg4CqL39yzU9iasIFrV3LjCPdmVHtSIXBj9CZenHf4LVMvJGi0hlkKUhwuRDYkyHdk5BN/Wh8Zc
CoK9mOdhN7g5HXCncMggTOZoZ8Zkb9ChG/2tPhN7zOgH350MTLAz+v96eypJWP8AdjTHxNBCMfKg
DaTr+uUI2D/TGTI3pPNKzII+SaL4273lXdccxrrw6JxyS5u6sU+jFsY+L98hLKabCqMVQnwZs8k9
MaiRrUbq5ridDz1ntaGatQOkLqCBpW6p/S9ZbaMYZn2ECIhEEY+cGC9zEhjaRXUQ7RcZLNzvfcfe
MRbzoX1mk6a/nnHegywgTMnSm/9YdnOFgeogK7BtFWSrLQ/+01Qx33Fa9i6JJcET0bvb5SsoPnn5
F3SrdZc0WotV7EMhfKDh7oOQ+GId16pNj38mcXneRd4uA+3kRgpqo7dXvQWJ3MvcYbf4Jyujr0FF
zHAJvHi1ZfKDof0SJkiK1oF2XQYsQSkh8qJXDVsDlu7SERBIgBQKF0Iu1mc/1njPCeQePFuehkY7
vispD/1OwiRKR3sQetTb2a9uKPQcCNUug+sucQJcKzuxOPgAG5AbGwUUJ4af6QuQXSsmdfoFqbWU
226yOLZCo0fy3EnTbHUShSnfrREoiynkmJRC70RHevfrybVy4WOIituIK83rH4/7lNWJj7f3cNlA
uStZQI8tJ3T8kcWZnzUnrChsV5iCqzNSklKUZyUOzvtLKPePeWeedK2VLkMVbE8XgP7VFglff1fe
TQTKaoka0g7FzVdEnDR0Gji1XrAmSCBdGw1LkkObOzYJUskj3x4D/UOg1EPSVIObcdxdf44S8lsI
+RQBLeP62yo2X/QE/QiPTzwk57tRR7xUiUPquQEL0LqswOvvluoFJJYlhuyQgf5M/7I3HhLD9qEC
tIm1fEIKzxv4czi2vN8ktVYPoNZTajEfNVGfm2Ttj2NkdwkYBhk9eEDH6NGlbzMUr5G6JHyW7YVX
crMX+lSPL3kRPnhxTg0PEvjGClc8H5EJkAK7lFln/O76owizHXl/0Re3fK9W5gvSrmtOe81lR+aX
1JfELhKEFQMDgPEm03I54fQ9WsAfuitnd++4FhJuMzgTe7OfendMKXrzn6cN3EZWEYMNO+6RAtYL
3rHNV6X6VdDBW3iIpTT9mGBKh/Mkfxtqx6nf1n52CsnAxhVVGF+QZ2vtRxTc+s+4aH7wsmIQ+SXT
X7MzX6ilwwDZ5X5ib+XdwPopaWSduccT52/h5ooLjry0NFGkyazsyKObICrkMZXes/SL3Iwkb2nX
X7ZJc6hs2O6yZm3W8OZY88i1Av3XcLJ22A5B+DRfeCoRiswfhw1CZUkF3gjs1cR2wXfUFyM1HOI/
WenzymygyQgxin2sQ0dPdzudm/B/+oC00NEIgNLyUvXVT7dn7JB5jCHOmIUAtcFBmF45pIFKIYle
NXZTdUfmQ6F9NgXrSWODMYpkl0u0sSRh6daa97ymGWUDw8fvhYQAdrKFm91a0pyvYsusboXASyaY
AscVQh5Sq41NBpZbfVjhRXMhsnPNBpAjWW203i9BEwDFO6cXZym32epaDS9RcmLqfPEwOI+cVwLt
LZ/2Ltgt088gfRoXV7pLFwST7geg/7ZLgMkXr/ni4BNHTU9aHG/qUOKyM2KQ6HNoS8TK4nkjEUvm
bO1ZndBjZKzg6UuMKAwxw4IHKOvqB6odnmm/b0HizQr/9WoMQenoMoytCxfeYiwDIqrc93ncig02
kHGN96LepEJbiWpGZRLf4ckIy8JcJcph1VipJeTWleHoB38q67X6jqppNI/yoGtmjDr4DhhJxOVX
J7fyptzwX9Lu6kkPQdmhn7DAsaNdb6s65w1aNK8wWa/+MSIA35miwX8yp8iHj75BrxjOQwX+ife+
rvOS2DLYPU2zwNfAMPe15RQC+fdQJYBlUlwJBCaP1yRxDRg+KXEA7/PmBLgGKljPG4CnGfBV48/6
DeWY+EjlKELqi8akGnnV8VP8hYYSHmtarHd6DRV4JKG+aPxWbe160Vo5PIZ4bgFLCh6yyP4Txdpj
6PSy5fPs32756PlUkB66jzfzR2Y631yuYqpGJoQwv6r6XQpyzG9fKkGxNEgnZXCYIJ9pS/Jnfc3l
hVSShCIXw+KOuGmquxd5tAdRNPzmv18yCvp4Gkp7ZRgI/gAT81+dZ77PvwClcp6ea+9WhKyUpd7D
3NHYdcLx0qhUjfQ6Yk6fGiSMdrjyCN4rl3XJMR/ucgTFTQFwIeF59IEAJMT2UoJ9kRdc03u6b6+J
5+Z6D/Af91LrkabjIN6SEPZMdxurTwF1D5PR3wMYfvNocBpDY+khI4pA+mCSnayipfe3oHnQc0ic
EPJFoB/YHwINrvnI01uX2GCT8unQXnFBBRFEWsZOJIiI10h6DUYAf6fw3q/rM8yBRDuN1aouAqxq
Rdn8VWL6hCLpyBrb0egFEplEPbSXBzZSS0klmSkhIbTx7DXzLRcS/9sVZmzClUuGTWzA2KdJ7OTA
vb+90Mzg0vqv06w5xIaz5XxxuSBW6NuVRVlK9jPwkO1ehnX/buJw4GsUz8X3NIiy+pJX9w5ktNae
93SGcJT8hsSgtBMTQdU7voTJ24DhcxpuxpS1VACGkphU8XHN8RzKgPXxR9jizQ9HGhfchfqn9S92
kzfA/RCeKRWwqG/b3LZQVEAs+aksukZXKBxxueeCkF8S7bWLAuKSBxPUYkBZrf0S+UT54to5xtZa
POI4bFaZeU3MncXTaTU7snfANjibXBj0oA2FWNaie4s19mFca0MGerwyZvjzjJMWRDzztf1DPW0h
BacBkpzydIKt30/arJxhndnadM+DvOLyXtjy8vYt6cZc8D4wayk1ltTKf1ANmPYDj0kS8apSUzvo
iVuZAuQoCUb1q3DuEm229bcPxkTodPMJa8/MtaU7svhVZZFZjHGGy1h5+sh2I/McITZRHfS1KDeX
RE0zuYVyt8T06vEKmZV/q7zkY5WYe6E9b/Keuaq7YtUpYGAr3/Q+7Cb2Yuh7l+kzyIDL1P/kgjJh
x5Cno6X0Jj9PZrvwxtdVlTO3fhjo6MNQeZ7Z505+RvpYB+/O4xefgKlNh6pu+L8WEbOGBhuLW962
h8VxNRskTBh0SpCtinAuCPXNfTLt6Rra7pNQViLqPOoHmfCk7im9nQ543nG+4kH8P8j/fzv0i8EZ
JOII4kSZkgk8brqIq1Wql+JRmftKNZ38a9zBPoJb9EJx2dktFKdJvs0pi4J5vMRvVzpfxg60S8vC
7DnX9P4M0oQ3hwJNscQbunueG3yDM/i28D/yDYRfpd4coQ1g6yTp+9bNW6k8+MgMVsoM95vnmcg3
IZ3y7ixeUMKwoLzIwgH14YbEQb6Z9Vpqpn2rRzTIIc58PBP0B53OHTGj31qVGamS52PATNg5JlHv
BXRwuRP0m1u/A6vAy1wf10COiozK6igIROD2H8CHtfcX/RTkL2AKJXkks2BlKW/fe1Xs1gtIH1d0
/TRQqpYDUBN/FFzUpJOBujoayk/dkIb9mmlqpZmmHFAz7kZ6hegXtGGoMUMCDZlWZYdBaGtUJAhr
8XLN9Zcxx/IDgu1T6dZWvj4bWUFOM/Qyrs4ygIxyN7s2KVm36ZMAWsNXbkdWW66H+p4AVquuEnI1
nDliECrjc8aOdrDMtzMfc96v0SmzSyIX3tXa83czOruwgAn+2/Ke+YWzavsxuNAdwPhn3Cur8xwI
aBPjMT2ojAJPk0wIJ0hY8tZ/hnLeKC+Jw934356tQ3QXANPyhmhPqElKk9sRJH5J1KcebfLFYSan
D0Rjm6/ooAqND3Cwi1Ghkofxa05z8OPrOWdzFK9tR2B/PBapB+53Ptmd/W3TVTUcfcwnouWMd9WM
rIFbHjy9ob1+U8KXi/VWsGjMMyz0XBOGMvVoEWaeminTEbX40a8yCboNLrRBQBhyYCEZeoeQvDvT
n+7tDDuzgwS3p1eyHxHmujUQ5hT/DHTAUvEZwAiaFWt1v1ggSp/GnCuwxkCj2pCiPuXd0MIADEem
P8xdMzrt1GAQfpBkbAu1kvFyRvwHjUSdKCDGpPUZhj/MBTclmO0hf2vx+MG+ytRTm3ftDBCZ+dCa
yEJQVkTWSHmjzLSmhb3PpXWzLjpW01eOLNGtfKXgcitOa7LRYShFMiSTOKs2mYo9vJsHaZK+Vcb4
phtLO0FY2hwVyjHtF/xsn6U3daJ0JqZ5lw7ex8Y90E4pMMuv5RekKmMipsIk7J4+TDSySmuVNn5f
Wd7W2MXMFPur2BZ1IjwZIOchTWSE7jACeKNCMe2sG6Oy3TeKWDCSJBxtNFQnTzowgRP8k/UudzcB
GqGEIH9YG5dirkfAys/uFHQ6J+jT8F/oRIqN15fHMWeWNvHc/lmoqVYRbg1ojuTqx2Qh36e3uZqL
XlLXboLdI7NXP5NgvschKM0Fxi9dH9NkM5BBsd6Czrg7VkAUOXXpospGqZxUrqaj1EB79/sGn9zL
CTqss+a/3m+qWx/irqGANTRAfYa3+YWaI9PgUB+3g8Y7x8p0E0suonFCDKJYDyUDc9UFmuI5N4PU
aV+E82yRVqCbiRU3y865ZW99BhtS4K4kUrmG/V3xdrlol2en47b5G/D1zDau3JCIIXgqiGwFeIF/
v2lsbXqsCacYwK0hwmXV/XWzuwubakqcB09M7IuFDTTemaQtslpgSeW6fZ3GJq2cusTcZK4kO5st
0rHrG0sfBs+WVDiMhB1NE9OiIzGm/ydEoPzAsizYoZ4ZSTtZxKksoM4lJ/G28UVlZ+d9Sqd0KOvF
NwuC5Z+Mlr0usK0LPhgrOfRsgv8jUZYTuBK71W16oiAxFj5XncDfCK1dGqXBbJ5Z28+7rOHOVYdt
Y/Ou0SDaBPtj23fZFoPsEPbOe3zb8UDAox8NTXn4GeedsAGoWMcTT12oPY5c2LpjHOWoQ47E/rQr
xAhqGIbQQagy7PiuFl4tI6Q+h/NdjFxn25tW68vMWW+Bp8Q/hjoGF13WyScmOyemVmrihYPUj7CI
6pfgwa8l5fwYn2S0exLm/kc+ZT4EK8otIzNGLiIdZuTLOiePrn73kz3lk4T6EC2bMuw2AzseX+cQ
UYpBrIRyxr4xrbvo0p6UhHfNcC0Oi1HGluMXN0W3jYjxtjr0jZv8H6EJAZ1mUa6HqZ0BKf0PlE6M
agl5zxxAi0ixZkk24KP43OtvSbQG1Y0IyjHFO9lFgRHwBO8okNe7/oU+tXgPd7s45Nx6XfUaf7/1
Oi4J9Bw9yQQ9XtqB12ybGUdKHzwm1Tjc/MOVUZmpINQJcS7JU0JOKK4NeeCDHo+OZGXcU1BkMLV0
skHRobwdKO+3FPeMIb5Le5Zl4NNqXZ6HsGhy1qTBCto6Aj9eiuaDJ/nxBJuAw7UYEDfdNI/bzDi0
EgqY45rB1E6AFQoGznt9yJi5JWv2n3Ixt7t2elLjIORhxMCx5OfPSbAMFv7CqxRHeNv+9zdNrHBC
PAsyMYVw48LhwIt7peVuTL5HPPj+DdJNdyLUCOTaR//LCLYaxC3CScgdVpRG4f+ePi1rjAYmxYa6
vQQN+5DUDQdtufJwesOH9e+lqY0u2uEAji90C47uh/S9NTafgzOw6KK3Wo77B6tLCQ8LDugwUPcA
X/B4K4JTUnRDTqmDWet2NgpszFRo3UEE/54t52yVlqBBjNBjn0dgQHImqNdhdqVA+/r9spjrWpTs
4e7zUg5DfLd1znqgzIIic7ig9H5iItTMT8uacAjiV52GcrfvzOljoKxoymdFWdVragFpK2cec1uS
ClT8Aut1iqUO6OpO0UjC6+44ajV3wQlWrQU3X8+drCRdh2AJgGgj+cNKxybMyK4Xl38ikG+NQe9l
EEPOiiGw1YFAVB62bhO0XY9wPtZnHhxKrofvjQc9nNFEifmB9+TCQhaYR81yDu5XR4pVZOWeDFjX
sYs3xG+LInmD4UhJAIQx4U6OfSTHVBFQonk+NbvAmV0CltSc898mbXAW4hKt8BP+1YnbTK4o01EX
t9GKFVBd62vEe6SAv0Dzab93ovSiXkoX8Yw8OV0iixVnVOaiW3aGzlbLP3OWmnSM6FYNsKvxovEI
62sHFEA1ThgeJvT5KncvZl0+L4aih4j9z7DU3wOwURkyRENKGd4yjQ6vJ1LDREZG7BMOK2P0MJEy
Ssrvb0N/ZxbeIw15zGtZwbxBAnju4zCmacMdgfO6GjitK0ngSCMVg6oTNhbl11Yp9/MZmUeQFU9N
QaHPPkGcqx1TBtcM5Yqk61CljAfmnHFQjwCtkaxKzYm3ifI3+OsxweRLMJF5+4zufCVDo0ibc+2+
nAz/mqEFi4HsVXYAhpzb+DmEKSk+k15TZi3gi7kPUZd1O3I4Y5mfQLjpqsOS8nj1Y5nanuMU9xwk
N1mZDQoIEU0bFqwz2T1+49fyDOnsr/qAcE/sKwVXtINHsni6PQNXhIRZJLMG8RAgrYdoyUlJpqvX
0BajRdQp9YWgGbrcEHXP0G3ffKO1jo+y39ZrAF9tUoMB8S/tPbcX4kW/iX6YyAjEpiDJTGutTkkc
OEdH3kCpmor7DrsZBS3hzwUP1H6vDg5r/kkHVCQR1wSTXRq3UOw0WhFm+KoMLw3zkWHkMiom3UYL
0U30dtQot2fOke48Mr0I2k5y54yY9VPJctpuAU5H1n4Yzwg33j03O0MLCxZOSamhtuE0xlhAQHua
uZsJM2zH32dE/NbKbGmHSJhwxuD6wh7ZOt/AARq0kM8RGodJeISjU0y4PqmWKX/gpP3209ZogMFE
B/Nd3JJvFwMBY/ke3e9lcSO8c3Y0xj0GUiZmAx8nEeIfyNmeK5FSNn26eFImRRxbrRnR1oe3uK3C
x81j7xXk5ndr43CjEckZRqePaXdQZLx/maq/MTETuktxj/s22cs+Z6R9kg4wQwssXEuoeZ/2b6C6
C/ZRye4D4FoUz9GbJRwEMiIzWkoKxESH/gAKt8heVuogSdBa4M4e4kLtUrnxYb1IsssiAGSIZpRZ
g4mVFASULrKONkdxuy0oFiZj3Oh197tCJhsu5i3o6uYKPGMUp04EZTmUALLQsQKnb+UfQCfdfOvK
UYOl4XQgRaXp176EUYBzCpR/dLiMn6Mbt3hKCTB6OfhVSSRSgkqkxfQY+jj9hkxGF9+e2Fg3FzHx
tlQ+syhxSRZCwoO1WfVkjqMj2SKFDR2h7nQMcaxlIzuyPU3B3MqsdwDx8d1f3E9qCI4HDhexT5AB
aG8NtdzM55sTkBuKhzDxo+yR2zBZ5DHGc0EUTnQNqYuPovzb/wfiJJXntIQfVNrDJhqGwBgiA6i5
iGambm+WUS19ivuoCVhtUTLQYPYifLP/QpxuUx9iPmn0XMpIBqEWNyxjKW4Lh5gDpmOB2xLXA3f3
vbPad11h76gs10f2ekhZAFUOOQOTpYP5W6h3yiAAjBKYKzApL/yyRGKyTjEr/uiGlhgnFJDUt/W/
Z0OFkMG6JCp7emCLfG3F7WDgOK/OS8P941N5wUNGzGfHmVJB05Hm7kF0cJlTLDKRs9Rz5YaRobSO
Bykgs5NpHuHPobmZ2gcDmSF6XB6e5Gnq3MpC9ZEJaG7WdRa2sPDb4AppwTXkS1b5MU56wwVDQ2rb
tz8fN4GOhe/rBPUL5nyRvtJPXaiRso34G/hdWIP5i40FXIoCViCFkVJl13Il0ryZpR4cteGSGNal
Of2cZuAWQuEWKYtvlS4kQjQ4qBOQIrkwuHKR9SlWE6LBcpyE/UNiC2j6ob6gw4GH8zb5TRSsN3GH
9/fpnXbzzBf1qsKNN5F5TdVMOWiWrUArdeRllGC0KfF17nehVfJ/eGYM/kowZ8CLjI/GcMPh36H8
vKdUVJEkB+4jeYZXcN1N9XEN7p0Y6xr+L2x50ncTVzw5vEJahnsHJJjZgjGk2XvHdQdZ4yFsLxNc
Lfv1xC8vMOvIFTnxmFVYsQFcesqEIGN9naYz4ut1RfmEZZyIhyZhax8i3hmdVu1Yb1a51pHwyocO
6ECZacifLOgRwLqvr8OqQ1zs2TYkpFo0Cx9H/5JDtekoCgWwV9VbtMbGbMOAqVgGSjhHNjAi0PyO
At0aNGAJk5Xg+h96XVgCRTVlugPvIONuTZeison+mKLTpSQ2o434WDmC0bqmSNrCijshoh1FDGlE
fsCiplmBadE+rMpNG/wVBdaD1pc4dwbZQ1k1SgioKDFwVR9XkcAdCNpOHGDifP2X9B8D760t2y9E
ejFd2A+DNb/EHPagm7iII+xZ0UxAsTA8y1QhJveIYlUNwbNo7lJKlo1mNARd8STXUoTfc0dHOOkZ
cLdCWHLLFmKOhLw31uY+3dZttQglzVmDEtWDM7qJOum/44KSTpkkz76VUK2nN6JDUiq7+GrAojry
MiTZDivs/z9N3CIsgVdup6bBAiq00ScdrK6u42o4AMcK7kLy2d+CkkwKUTu+WdlRSYSo42lquc9Y
BN0O2orF8XMdU0CeRYpMA1krEirFfIHsaaI13xXaIjC0KjeLNviXMdoYEmcnrdeMx1Pd91GjLmAI
XGMMBzDNbXhuPqRL388W3m0Ms5qsTyeV/weh+tAdkNg9fMFmX7EuWVw5y261bjHQwXTaWMLx+WIg
xQzFsAqY66vq6VM1UQ0V+6+pDCGcxXvVZf3TGmcseTEbTYX0q5AuVPZ11f6BOkx+K89u1MO00yAK
9xfaGhJOGXwrzteEXwPPXNWvziqS
`protect end_protected

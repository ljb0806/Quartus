��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7�����������	$��BR/�`�f����=|o�hN�<Q��^0Fx{!o �<v��	 �[���y1�E�Tڅ7I'��7�'^#��́��y�'�a�� O�KEʇ�m����@��=P%#3��(M8���p'����U*9�����J��Zm�;�}j8X)��Ӗ]?yMm����mN.������j��p�]�H��%Xg5Ԥ*�X���9y�J���\���7{�f���]V���^+�F��6��?k	5�H��9�<���w�at��a�oA[3�r�QA���R'�`R�^�鷃07���)ص2����d�\�跮�:�˄�	
���A�6�o3��/�i�"4@��{�?a��s�OMXvH�-�ϊw���՚��r�4���<�N�-�>$�_v���<ƥ�3m��^kZ�r�7�H�m��(�l��9tz~���nL��gT�E�G��)���mSG�8F�	�����uG�l.W1��x����z��P9��Y���䚚���BIq��JW�(Et/ޮY����(��s��^O�B�G�M��-O1W��K��/�6h)Uc���7���T�Te�n����]���G���Mר�;��o���M~ ��6�8p�^�n��v3����yA��r�d2
�bU!ɣG��Q�����B�
�e�<t}J))=���3Q>�ǜ��Ε�$�6(-����y	����gB�Y�������֛ĢdJ����8q��c��je�a���UtaZ#��>9
O�])&?�g�4�7��.�5�Pu�C���n��46x�N25%�!���'�Fc�uf����	w��(��W:\K7�
��-��Ό���Z>A��9�:yf�Dxe�d��#�#��l��𖀤)=|FŜ�3����]\6�-s�A1�ת7������ņH��ǁ)͔����L�s�3���po�#���8��TC�!��	�N����|>[�pX1G9�e�c]�i5K �;�9����Ij�#%��E�3ts���9[M���-ɬ�q0)�6{��6P	��=O��rHdƣi㋽��i�d�4�S�(���ӱ`�3��Y��Nn��Eg���ۊԌ�̿���Q� ��ޝ�vF�x�!	��JIO�t�=>c��k�-[X�3h�^�YX��T��t�s�u]R���i$j�����c� VK�b�.e���~&�F,�o	:~B���:�Ar��8��*�n	)�ĀZSy��pI�|���n`�V.ûQ����������E�@ѩuU��V�uw\q/�d�����	�������LV�ïs�
LSuo@y���l2K 2�j<ք�����J�����V�p'ΰ�_>t-5�"d0��߱k(,y{'%�~�He��y��bz����{=�
�,�3˝\]��i� @�d��82$�J$zQ��\�[�����O����O�ƍ-�1����@��.(�M� x�s#�{E�mgW����	Ix�����o�}�њ�T E wzښ��DmˁyEN�. �IJ-a@`��"�V����]��Z���r��2�}�͌&a��g9����A$���c6�-	�G�(c�S��
b&NوP+1
2�E�!@����ӫ'DQ�G��.�
�a�z��!�vi2�s���6Z�)ϴz7��B|�ypn!u�Mn-�ǹ�2T�E�CqMm�SP�Y�����<�@�Oܮ�D�o����Ms�u0��0r�� -�4Z� �'/qQY2��3���I>C��1�Xl�u4�!u��E'���8��Ĝ)O4^�8Б����}M����e�ۙ(��������<�C��٣����@z�A�x�s�1o ��Q���<"B>��=)�`��9���7�[��-�`����i6?�.β4/��e&���`���bU�U�l*����? "U���O��^��uf��Pߠ�=V­�����Mj��(ə#e�IѬ�
6�N��jP���4#@ ���˽��;�ܟ�r�3�a���r
P�ŢK�s=���$�c@��4�	�p:�~i�����@I I��Wsg-ֈ̸��������s+q>��Ǥ���O�D���H�K�K~LJ.&Jp���PEK2l�X��ᡮ�|? O�+��Zǵ�fY�G�ǹJ# {ϕ���������m���6�ã�,����xX���wإ�<T���R������\m,�
����ȾF�*/�<4���,��VX�C�M��6<DW�L�F�~�d�(;v���3��$�* �u�l�&���|95��Ba�CJpL�r0�o�Z�:Z�ę�O^�S|��ǈ��ΝBr�Ys�?��3�Q�0n�5j/���Է�.ZQՆV'���jA��^8�v�
�2X��DS�asM ������gVJ[���¾z�;�-�\2)q~�4[�?bWk�	Ζ��L�[B�
�Ҁ��܌�h����ni�Qx�J%��#p0q�2�;賚��v�߸��;��Q�`G5�$�œd�Ip,u}��������T���?�3�/�2��g-�u�گb����=r!�q�]���X1*�P�B�ϊ�T�����<<~z��Qj+	o��
��سEŷZ[q�����lY�LOc�Rc�B�-w��x̚�M�H�\���T��/!�Pj,8�Q��y��r!^�+.|3���:����Ǒ�(Y�JJ�\ �.����}��$�e�M3r�N<gÁ��+�s\ک�s��U��y�u��Ǯ"�O��N��5/�8���5��V�a��^$}).�w@5I@-�_���7�!B����j���C{ʹ�R����ȥ{FH�Po�Y5�'�`��E�V������	"*�k��4���ѸB��- ėG�ec���ǇpS�>���Y䴋�Bxԙ{����B5ef�r��@�����3*��G�l=�G�+?x�̺)�o�ƛ�!��S=&�
^�sw�y�.{���RNg��7�ڐ(�_h�V0Hɦ��,�P �Ne�ќnR�<[k�8X����7�Y-@���e+O���|B���Ϭ&��~o�W�����!b�w���񸐖�%ך��I���<�D2/% &�_�R�g�,@o��L���A©P�6�F�ua�ɍ!�}�vGX@��Ez��1�6�|�=���r��C�@L�{�Uc��&�zc�!a`3+���G��|�y��}�5�J���[�����<4�^Y���k.�3�G��t�h�1���ߦ��*�W��R��;�+`pl�"�I�5�1y_�7c�˅��H��y� *!��!�, �7ýC��E&mj/�����T����P���p960#�ᑹ�+�NrB �ȡq"�m56rtN�r0),��2 yzGjMvn$�K�5?���{�
+�Y	Xk�S����W�0�z�Cd��� �G1�W��)��O��_Pփ������TϹOu�O��#�?<�����S����%[�6Ya ��&M*�j9aK@��^ibU���,5�x�8�bkU@�C��[j��o�c��˖�AɈ/��Jấu������dfI���e?N-�����u0���g��t���4s�v+B���4T)�U�
���9Л�{殰��ҍ�55y��qV��Ц�b�c�5����(lMAHp�T[��1��)ؠ���Z�h��2��ߢ犓X��f���[�=�? ��.��E�&��o�}uC�W�V�� �ս�ˇ�V���&!��U�ϸ�_��v�I ��YRE�H�ۉ�B��,�2�-,�n,�"?��.��k��c�DaTڞ'��0^���ΰ'��M���-�R:n�=��@ �6>��>��ٶ�C�r�K�ʫ�Es�3M��D�60L��9r�M����ѝ *q�l\��|���E�:{=��b�dZ�v�EJ�RM�tu���k ��M ��#D�TR�~�w1R�5\����� �g��jr���hF��w�=�kP�'�8��>�I��Jᇼm��0$���|��WE�ƚ���D������,'ʤM�b�9�y.�L���@����%|:���z%�/F~(uZ0>�'��������ژΌ��̊���v{�$|��b8+�l3�`�%�۵n�p�a�9 ]+:ǀ�0�
����F���P']mf�t}�A4$��+�旕^������t�֗���L���NJH�&l��+�����)}�X�|≇.�"��(>z��'kAr[�����{\�^�p����!�;16�i�Ѵ��b����,�?C�����;�b��#}��>�w�zQ�!�(NG�5�)!�sq���"y��?u7�Z��Z�|��A�D����E�:���l��i��ܻDA7�j�6�'|��q�^�+��=E�^�n��3 �f؀P��ǉ��/���Q����g��c��԰�<Ș*p�/��^?�Q���Pܮ_W=a���RG�5�j1h�b���)�0n��b|L+�bL��Zc��_I!wȳ|N)�=��ǈuN�?�wa���	.�Js~��ji����Y[�&I6.Lc�*�8�q���fuӷ��.�7�X�͸갼,�Em0�/�-��d�Tu����'��G�q%��&������h1��D���%f�`�pL���N�(����F�CA)#ت
���r����LJ��)��ۼ��W٪ȸ@�W�����ӧ��$��)R�L���̝��(k����T^1�$Ư_~�]t�U�F��A�N����A��hh�`CM�m�[w=ի�V>ܔ}�na����D9,ǸSJ	'�U!�㕋���V�eW
�F�b����)�����z=��Ea�cqML���xa�ߊ �Y������?�b d�#��{qqyJ��:iG��ڡ���T(��C� d�!�� ��mܱ/l�\,m��C����������i�\�5�h��r���N���  �����X�b�U\�7���s)S���`��W�%�@�Ȩ$+3�vԕW����W�I''���{Z��+<�?�D��S��6��/d��a���F�x0m/=h}in������<�E��ƘĂ$�W�4������#0��D�ۚXӕf���}׀�ߌ�\U���R*4�u�!������������P���J���?LO�m��Fm!|�or�~3dKa���d�םc=491j��@uZ�7!p<��m�+�.VHV��g�s}�ݸ�|މ�37>sV�)ٴ[!�[�(ߵ��d#���=�����;%w�K5&`�>�Mx�(���PQ�*c~A�6��ɩ5�DOvNy���7�t�y��GܡPu�ߢۯ�0��RpG��%�JU��l�\���N��t��I�P{OK�QY]��ӡ3�?p(���2�8h�Ԫ�1Q#�yд�v����z~Rs֊��d��C�M���1sG����ֶBl�[5���	ݮ��1"�1K�J�0�gS�IQPR�1��I����o����I�Wwi@wEY�V1.�)��QPEl��Ǭ�ms��:?�lN�x��^wEҁi�Ԡ�M��MiC��br�;j=�2�k��Օ���ޗ���@z��
p�1�P�`J�s����8�*B��0����Ż	~��{��c��}Ķ �;9IۈikŽV�j���K���؛�ƫ���m��r�@�3A�Nq��,�ߘ~�"���T��;� ���8��6��ע�f���S~*i�c���z��Dr�[��D�p�l��u�Krm����11�>�i��:x���]H*P�._EA��uH�`tΕT'"5שg��fF]���ggS'��f��3�Z���N��u�|+1�����{�M��Ȅ��3}���T�����(ϫ�H��	��|�(�N��a�nR��`�|YʩP�D�)�Q�V�0����������KA�^����!�[�]d��k�L+����o�����/,����C�D�������G/+�Yw�C��e��ɂ���7rBu�M�z��r4���}�څ��h�>�K��UJ!����c�A_W����n�	��4.���� �l��uBQ81t�؅a���|¡OL�F@�-
Nuޯ?6�~_���y��Җ��n��Z)[A> ��'�5�<��W�s� �
L���Ȭ"`�6#���?�N���(Q�7��p�}���i����?xy!��ȯHR4�`�x�9���=�ckQ��,�f� :v�a���;���u
nL� Y�a���gt���\��#��i��97_�&i˧�w�!�����Ha2�,`kTT��A�qZ�ĸ�{���-|�]��^�Z�y2�HQ���;,2�h!Ɗ���T_{���3+hn(�56���&b�{N,��C�m��ɝ�9pA��<.Kt���u���Z�^6�)H��n�x1(��Ȯw�T�@�p���P�W+�<�9��E������P[���}�Y��܁ �P,cR6 ��L�XE}=P|(�Z-Y��z	:�0��	 �2�{*	�z���4�Nb3�yA��s��Z����c@�T��`����~�x؅����0g��g����nbI� ��p��O�����CE�)�"ԉY�pܻ�@n/�ݙ��G��}�٩���Y\�aSJ�.8^#9٘�'s#���0�k��f^��G�|#����Ki��)=�o���?5e��r��f�n������Y����Qf�;�0;Ѹ��7)��J���6�}�-��$��g�ɘ7�(�]���TTU��1��!O�k������ܵ�*��~��ng�GCF���`�K2��m�B}�j�>R`j�k��l��(�[�S�IŊ���8�CPJҌ�̦��̻����p@�6�� �{!KRA8Vp��l�%9�p+�v����9��Ӟ����TF���]Y76�����s�K})�qF��F�ꍋ�a�KpT�g��:�ۊDl�|,^�GO���׊BK\:��6��^(	4��o^��,���@P���'�䴹���A�~��۲� �q�@ 쥄z�y�����Q t��>�ͱ��^��R��8RfSZ�����;s4��
����yYIRg�I2��J6٫��kBb���pX?�K��7��7q��%�T ۠A�r���zO!ڸ�sǀN@�I�w�t&C�F���}���,�u��|ܪHSA�W!v�#&�N�=yDF\�^Jz��DU�L��+�y&SKI���^��p)���(u]*lތת9�8Z����Zq"�
O\T�zGgˬ`���(�* G-�����Jr���o2�J�Eb�`��.Ʊ5�\���x���<�I�"�7��Cz��L�(�bG{��?��ApHc��@x�f�z�[�K�;"'1 7��f{�.L/��|�9H>�w�k��W}��9�^�A�O���&M�����4��<c��/fS�T�D<���_p���T�tc��\i^��s����)#�@��dw���Dm��œU0�7h�m�U�);�-�G��m*i^��d��lNZ,
)W�h.�,��7�8��e�U�5`�y)��7�-T����G�]&&mx��ј�n.�9ļ��$D��d߉�����8n�u����"�$���EUs�at+���k\��T��@
ɯJ��`@���ޫ���4)Y�RVk�y�W��1ϵ��+�%�� ��sK_�F	c�$��G��������ckb�a�3��Qe��:_^��S���h���� H�k����K�������}�e72S��1�f{�!�V�􅤄��I_��C�J�B^)�,��X+�5^����N���.[�T��\�B=�y��a�q���}%ޥ�x�Gv���V���M;�!9��Ɨ�0&�w�|O���)�
��Š�4'}ڢ�7ǿZ����kp		��\�F�}�M#S��"z�>�2�h���v�3D3n���gJ�a�W���~�_g1��h�(Bvj�[�E�a���G�hD��S�|�2���w��������pٛ�׆q=��}2E4�\������$�d��|���|^`Q��7z��
۹Q�*������̕�M p��^V@�z�z�-�E@���6��i�3U��LI�K�Đ���T}�q�l��5 Pײ�����'���3	U��%-��6(���I�������۸��,]#?7R���@��\�WN��<���FW	�Wg)���Y���"�v4 T&��SdߣA��(�P��S��Fnb�pI,FZ|�˯�q]����|��d�C
���N���$ ���8���O�V��Xe�E]�kɈ�`Dv|��ض�I���H��AQH�s�D���l?�Hɫ�$H���� �{j�q;���9��:�&[*J�=1�Î�>�v���6�=��� j�rNƞ�����
���qK]��M����9��ɋ
�I�7���^�'0����r(:F��&ϴkv�)e�Z�`����ae)����l��a��g�հ��1��@�Ш1~V�r�����=�R�z�ba[2�����~N�\��,l�m��:�ul�R�2��6�RO����V	�KIk�񥎓`��[�L�B����?	�y[[ճ R/=v#G���Ҕ�1����O2�A�*"O�saQ%�H�P��b쐾M>?h�zxa��d�����w�T?pt�S��iukF	�kS�+�^K�,Vx]�[��=L��������Ď@�%@�25���o����T\@��!�� p�/d퓝��u�}��R�9���
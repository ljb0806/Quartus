��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��$��~n�8�وr�����T��Yʯ�aQ1JO�J3٣�$�d9�J:����`ȉ|D��)I���{����>s=ˍQ06CRխ��7�sjLa0������/���	N�ע�����S�;u�����`��HwLT�?�1�J�s)��*�����Av�2E�9a��мA��r/P	&�!h�-y�!�����$a�Dx$h���,	�+MӍ�Mߕ�W갫��bf�ԀG�|�X'�6T�q�1��=�I�����p	����$�\�s����n����P���?8���$��H
�b��̸�x�tvz�=�s�''sj�մӓyޟ�\Iߘ�C��\7��P���l�x�n�iO����qGt�xŨ��؟{{��J�$�艛!'#�fy>(�3R�O�a��^e,��:d�,����*�����Y
�R��j�xPb�:���2;�ٴ�D���E�	�6��f/��:9_~8��Ҫ��@�2������<u=���5�f) ��LO���a�e�i�v&P��}���o�U�9�Ee[�hK���	�ߥf���<���:=(6�>��Ώc���e*�4]�r����$�\U��jN�	�T3x�0 K�5�_��[V�>�&��`e�¾��Ъ��6�`�P�G�������X��7:h��`s��b�͘T�7�7sw=�g:�[��Ή�	��'��A}�8B�����,�ũTwa�s��tq�m ��8�!$R�ɎJ��K\D�+,�mI��qLɅ]�
O�}ߗ�H�
LF��^�袨�׸#;P∕�H2��+�W�{6ZM�M����@���� �&�����a~H��pދD�iĘ��0og���E��+{?<O�^�w�҇#�e�X89aq���He����i�b�_�O�b.��1~W�5����.'�;c�l
��c�E�&���E7rVL��i�7=p��?��2�(2HE�-`4���M,9�]�T4�̃��S�.��є��U���l��h&��"�%]���kVb���`��N���ޝt�D鍹k�h�g�5�����%�NşG�~F9s���Fa�mXt�(;4��K����͉jɣo�@�]S�܍�Ԡ!�ۧY��_��������,) �xHT��>��d�c�v�g��/��Z�W���	ֆ/PqAI(���󥺭+|�zz5�:�}0K	��gQE�*W�D��}�Y"ͪS<Tm-�ޞʊԌ8�y?2m��8�\��
R���;��p .��K�óN�o���w��?�S#tjTv��ܽ���:�~�Sv|�&��Qe�K1��q��Lze�W ��%��8��R*�y��5�C��o��AX��� �5
G�L���~�O���������a1�B�u<��U�ݪ� �mx�!aD /EK���|�3��������(��$��������ú*r��<]��J��'ь���<MsΗ��IZY��O����n��2�+����u��]xvœ�;�����r
�nj�C!��)	������
��V=����,{�#ڎ%E�y���E��W��+D�sǩ�1fe��!ƜT���,a1��_� oxu]9���.�egǺ*��#y�	��|�y��K�	Q`M;k���M�/���}������)di���<ez"��S>����Ìв.F��/qv�ӈ��w(���QqP/�4#]��%�"����r'�;Ku����2�&�4�`L��[�{s$�3���N�쪆Zg@�b8��S����P�&ƫ"�NI݄�_PB�[�6鑌����Q�D������tg�������hsq�/_E�O���Z�T����� |D��y���PZ��4�o:V{��~�rS�,�DpZ'8�ZY��hڍ�%.=����1��a$�Z��V�\�\���ԧ�>�v������]
`44k&��i��+3����M�vߟ7W��w��ٙX�H�A��t�T=�K{PF���~qC��ϓ�_�O˜�޼y�if9������)8D�sES�"��BS���r�kh&�+�M����t����f�pӲ�v\������Jw�?l�#����=:��K�"�
i%�O�3�8s��]��D�9P�U1\[�����O�e
�l;��p���D�zD��=�FL>������'+�����#<�{�nβ��Md��#$q�o���d� �l������@闳ҍ9n0��G���̽y�,�� �bkJ}�==�Rd0ˣ�羃�5���������p���C_ ��ˌ>O�n��__�iɁ=Y�\��s�K�!3�!���IK���a�k�hu��0��Z*�r_	����s;���7Qg���=��Ұ��m'+��JQs7��D&���|�gӡ�t����˼�2u'��o����$�K�ʕ~���0e/��v�n�;�W��Z�H��yX��Y=�h�"��Y�W>�]8*_?h�ԁ�7�"I��5�Y�ѷ�����?���w�ʉ/+�-!3�h��)7�]�3���B	B�:�1��0���^_��94쮥M׵ɥlmv'�E=�jY��~���r㈳lOMA���͖&�����5"
��i�_T�&0�9���W�8I�ۘ����=�W6��A�|�Q�2��L��f�A�&�C��%�IO�/����-�����/��:N�m�a�=^`����G`q�:�$����[�e�	��I���˘:�?�l�'{��
��X6̻b�n!��}'.'�j�Ζ�����k8/W��v,<u2���u��%��f�u&�i]D�d�V���#L���i0�W�#O�5���R�G�P�+�#�J��y����i#ej�(��dpp��e���y{�Q
�؟���ʎ^d��?͠b�8Z��!������b;"v����J������������В������}�@:ਜ਼����h����[����=�?�yB��=v�P�}1�����';i��\��yIH~C�'�ԏ����yIh4�Nm�����2Ж-�&�ߠ���B�؊q�c�W�� �b������0����!k��X@��j������wwy,gq��Rc������p@C�z�E�Ѯ0����������#���ᣐ�,�6�gc?��0�4��A^�Џ>��P��=�*vɃ�
8�n�����=:�h��F����qp���aeDj���A�)O����T��<4{�!<
U$2��a�¬i5�Ml�LL7�����|�)L��� ]JDef����+�)��k����z�8��^�M�����V�����N����x �������X��g��LU��o��������щ�T��|QQ?�G� ��3�~���Pebh���3�-p;�%�s@� �m�ý�Z��D�H#��Ky��j�˲��)�$�;ٔK$C��۳t�u�K4JD���L'���4@��&q(2�MA�ͳi�P�;�#;�G�(<���ğ��C���f����ZU��k۾P����q�aQ��vX.�#%3=��P����ŝ�,U�3��(����X͉p�����f>��y��!�nղ,��*��Ta�(��m��(|��L��E,{�b����\ePL�na�J�%�H�G����J����fI�leT���7����"�0+������̘�:!8u�e�Jz"��ip~��s6G�jH��K�'Z#����Ib3���:V�s3�/~�.�r01q�G���!쁕u�_~>�I.t�+|���$�g��:��sW��Jљ��2u��N�A��m� �^J�eF�V�R�NW)����>x׾��5��o�����Ws�h��y��ݺ��
�"��P�����q?5Zz
��~���l;���P,�v� �������n���0��vy��΁�N@��Vuw�bZw��_Q����[�����s���D�\�ce.T֬�cmؽl 3�ү#M�U�<{�G*F��D��n�Me� (����by�S��زp�n�0'�u�1U`�؎i�� ;�O"�S��>o���jޛ��N���@W�Xp� ���8��-���Ǟ8��a�!�s1@6JV/:N�ȅ@h���/����p�I��u_)�����T�z�V�|u��X��w��oXB����V���G.�C%��:����Ґը�����-gvΑAYW����2/uM�Ѱ�Z�OYR�֜����ϑT�QA��R�fK$����yL�j���(+�N�6��V'�?�%?{������Ը�W�8�����_*�����+į�����Z
S��1r_8Ml"Kߨ�I�q�&4n+.u��H�&2H"�do$�K�r�ˆ��Ζ����k՘44&"C~�rX��3 �����B��b���y���zC�Y�&��$ZG�F�\@~���	��&�;����hĘ��l���z���M�Jf|^������RR����qqX�K�^֟01�����FM3�Y���3fb� $��V�rW�A��n�l�)X��>-���q�/�վ��YeL��;Q5��"�üHk�0�l
`��ћC�ǿ���}�c|��RSs|����;�]
>��#�cr��B��Ⱦ�كaб���}�� +:D��w4�s`lfk��j�ѣ���h��F�\[�>�(`f��ψ�������`��$��xd����:����7���@[o4��F�,����GŎ�֗�J{P4!��A��G|$ٗ�Y��d���+���dR��(x�k�e���cz��ک�(��=F.P.f����D3hOw+��͏y�F�|V#hҝ��L>��I����1A�$�6��y��AXu�QƂ�3���"3���^��<�c�k���Ƴw�7g ��Tcc8F-��n�g�]�����4��)�ӳń�+�'ɡf���񎮜4��T�V�Xk%�����f�C��}Rv-Z�&l�098�E�ɯ(,H���z֙�滁IE�?����:Y���wg�d�w�&7rv���(Y-�)"s0�+�ј;X0ד�����;�OA/��9dA𴁳|�q�	�L�� ����\�MD+��0��	��t1��!K�ً���C�}�d�tW���'v�$w���^7��7�������Z�wf�t$Ǡ�� 9F4��r�?31򬤵�'y�NBL��)��f
HO��{�&���(R_̈́)�����"5�[���8�xJ�u�a7��W��|����H�w�:O�B!Ϩ��kE���?�#� y�-�(���z< ��E��Q� ����x[xH�!s�\E[q����&)�%�Z�/緒��[�$ħ^���|����{�A��ML�	���XX�<<�;fz?�	n��'f���_����#��G+
����ϧėT�5�h.仰W�ز:*�h�h���j�_����uOW?Q�~�D��.5�$9Հ�����2�m�6�/���j��/�^�oQ��*|�"���!�	�%c&������Ӂ��C*�����Z��@�&(A�F�L��K��9��|y)��4{���jq]�H���k�oY�o$C�J<҅,GϨ�n�͌C1�&u�(�oy�+���pkq���&�f��-(�Jl�X��i=J�C�;�n�b�b��2c�u������)�I�:������ހ��Oj�������> =E��Z�`��-�!�cw����P���0�t��)F�o��_د������}ص=�NX��-$�Tϼ���c^��]�^$ꢖ�X��Mau�%����R�69��/�[z?nI�v?(u�+����N�p��Ra�īh�C�P�7����aa45dS0��NK"3S��Koe�l?�m�8r!���?�ھ"ϻ!��r`Z�����Ku�(zQpmm�Ӳ9�nb���|����I��Ŕ��($�3m����{L����$���@������s�����]*2i���JZ��9
�s �V�~c}	�"4�'�r������νXQ��E�ʁ���0'�+��B��+��:)�!�'K�N����'$7����F(o
X�/��&�	�&�N�*gAJ^��7��$���v�K�c�x��.r�﯑�̂����\	�H��P��彐1omc��B.K�v?�7e�g�t��o�Nxʜ�:��2@�H�����\��a���Pu�����\z�ҕ�c��mںXTV'ld{ⴞk1WǒH��' �G�_j�~4��H:���fʄy/���m9�ى���)~�ЍHa5�XǏ|�^��������8Wb>��t�&�ni��h*�W+#r'z'j��A�@��&X!!Z����d�?��0�u���{�8����%��������-1�ɪ��E���aK$�3�ZzI˸A_���z�dJ�[�~rV�*��A����d����q�8S�A�}��'�4�M�|	Y����nPaA<�So�k�B�yV�ܭ��O�.�Fn
���n�����[}wp|2� ��?9��^�3겺�pƍ�}ӿ��!��4m�	��@ۦ�j8B(/��} �o~�i��޳Yh~4��L���'��QZ�VjI��N�E�^7�O�TV���)�mki��p�5�Q���0k7���Ֆ�1����f�xj3����HhOʺb�� ��3����멶j��@^D2c���4��b�XFPOAV~>�d:��@E3���'�����|d�%��8�w�3�	�Z�ar�z��+#����K��=�=�����D����J�2\Z��Vӳ͞Aft��Z4s�6M98믱��U����x�m+��n_EƝ
C������$ԧ���s�9T/Q����� 9UWZ�3���{�B�(@�X#��)�h��3��8����M��Ȼ�M����z����*�1(�����
GDrnJI�r@���R���4�G�H�c7IIA�NTn�.��{C��ƪ�c�[�'@�Aj�z�fj�Atv]�C��F��2`�Â��3[��B��ug��E�R&�z���.zG��#��hH���w%!���V>r_)�F�}�;5�k`礧����.���l��'��-;r�2`B"�<KN���l�蛝d����������.��&�A��h0�V"���7���KΙp�lYwe��t�Xf�4��]Ԯ53�% |�]����Qo`�ↄ<FWoR��8/q����dZ�1�FYe�R��;�ks,%�Ì�b� 1�V���́r:���j�&b���\�z��~J�7#?y��^���?x�ܤ��Ђ��Q�	u-����|A��dN(zLa�]��d��E�s���+������Z�ow�v�A}�l��.���Z�2��^�/�5\��6e��qk
8�I�TŽA��Ү�S�8ʸ~�u�}�mh;�h� �1|�I+ѩc2��UK��]����|փ����&]���`v���"���Y�NF'�=��a0��[Z�۬k�-�Y�Z-Ao,�)WX�����1"��Ó;=��p=wVԣ����J�i���)2���9;�P~؏Y)���7q�-ݢo*����^w|�~�ã��AW���w�L��c�>xb5<@���T�d��w���Z';�O+C�oC���/�Uߕ���Ȗ�ɧ-�g$���W�B�#�\�V�է��ML�j����>k-�����w�:���J��=h�J ���������T_��� `�z~�r6'���ϳS�T\�w�i��٫,��]�	 ��0BV����_����
	�ٟ�L�W����=�z��t�����@���/���?"��ʯ��� ��0y��O�r#����<1;;���\����˝M���/�#�i�cн$���n�4%|ݙ�k�����w��)��6��+u^�?A�Q{��O�,�l�Ll��żٚ���Jb��%{
�9"{�3OSh��"�G��������$c���ǳ_�I �L�(5��"�cH�@C1���=I��.����?֬:���:�	B&��g�5�C�)܌����O�g@���\�1Ӎ��k�q��tMXх��M�nx�#8nă9X@P~�p=������|�:��PPO'�v;�<2$^�W-��Z�l��;��-#>x���[����
�p�lK�9�]FOV�)T��v^Rd?o�7~u65��#��D��x�\Xa�z��`�c̣"��kn��WO����qUeȡ�#̨d�J��pܦ)7���ځ�؞1��w^/ɂ]��(�~�!��4 $����1�b>���L�]�2�������.��p"1c����BAη�3?xP8�ʇ�	m}�TP�y�5�`EG�X�#6϶<�T�t(H��D�f�D���K���p|�{m�6���&���f��Z��wH��<q����OGTs$9~�)q�ԊgQ�$�9<fcp��tU��iB��\�0��V|��s������*Ϧ|�"2 u΅E�g��J5!c��)}��0�0Ĵz3(-}T��Km�&���+�fsK�b�!�snr8�6CY����'����>��Ǐ�a�{n[��!��7� [D�
J�#��?��P�+(̹���$ o0AQ�ۖH}(�WE'?�t�:]w�3k���(�|��^Fw�)ZFN�nwz@�����{��XS'.&,0���ӄ��y^���g��U�2Z�
����aY�V?\��o��;0��6�>@"V��~�<�u�m�R�R����M4�D�FS��������$-��8U��߲���&;N�e� J�V��O���ȼ�n̻��0�Z2Sr���ͣ��?zɋ���)�ӺT����U�٭TKh��xK�
��x�M��L����� m��{셝 ��*���t_DΝk�|���t��b/[ ��p�T �h���1��|F�V:�R�$�-�C�*�:F|���s�����L ٟp�����i�q�bQ3��Enb�a��q-�6�3����1ď�o�(#��~�aW	��"��<u8h
��t��Ud�f@|6��SH�i��I@�73݅,�K���=v��WSJ'B5�T���u�L�|�2� w��,b[���-zN�L��Z/g��O:H��Bέ�0�����y��^D���.�9�o��	L$��8Nf��T���Y�1KH�4u/���i�t��-w�*�X���*�{S�`�*��f�^w��눭���,p��G�<ͲLQ��f�>]U��o��@��<LdkS	�s�E���(�D�n<3�1��@m{��3��C+hy@L=�*���EOo�FK�Jq�)�3���CTJ��t�l��}S�u�����Yn����ͳ�������>�q�ܣ�1	;���s(g�G�lB���j���D�e�����2����յek���n��o!�YCG]�@,�_��|�yҎ������ekS��=Mf��lf�uH������'����q
�=9@��c� '?�jl�J ϽO�z�s~�f�I�T~��4$�:Ju�R9�����'���1��� �������3�_>pR����BP�fR�H�:���Q8�.1]�����?z.�Ꝛ^���0I&���8�|����ip�>��qC<���j���6�)(R���!�N�6:�f����0���~Z�N	�'���u��������,7s=p��$K�Y�X�vG��4+���
����/�ؚ@#��UM��;fh �y���Z�b������$H ����m���\5�Խi���l?�2�oFU8���Фl�����1���9�tv�8���1�]�c��'h�j�
+L����~��#<�~)o1�,��bvuzg��E�˕�Vd��~_-[��@�G�M���R��I͐{�Ƌ�^c;�P�
��-����oΞ_?7�Z���e��/���9Gx��k�r)w���6yה�;Mй�#�xoܥ�����)����S��kԕ��\9� Y���O!��99
��4��캌���6���״����]���);�i@��-Ũ�/���<z�E�����sq���3�e�`ٲ��/�54g���4�����&/T��'�����"��7��)��1�^8���ө��:���6�2CF^\0ԏ��U];}��Bd���>����o�$@�J��Um�_/)�s��a?��,��|x�d6u�:����K�ˣ�Cjӆ��1\��n��~~��Cy�zp�3K��h�u��ໟ������j�Pwħ`;;��x�#x��sEY�Μ�0�p�lؐ�totM��6�[�����Q���	ʬ
�}���O��.���fu��u�R�N|�-��WJťw���i���+� �[�X�4�-��ҳN���Wu�o��Ą��G��*���>��<���4໰����4�֯\�x��7�����Sz���A�BP����hB�'��f,�T�A�����x
�5�͐޲ߦm廥���� <�!���T$-0��Ȩ�@���/kcӰLoi��o0lғ�l�~�}�Ϳ��6�78�*T�I�ǎ�wƓ�S;Ot0�3�)b(��ݳ�\牗L�r���c�R�>���l[Ҟ��HfBu��SB��4�bj,�m�]DɈ�� q�hl^_r�'B}��)P+lr�Z�d�\鋐�kL�ۏ��D̋c�j�y��{���P�F��Hf���'Q�*�sz����O<�<@���2N��ݺq#�"�Z�_&�1�i.�H��8����$�7�H<� ï���[f�JWZ��tp�y�{j��t�e:������r��~�-�n����pf�	�_� !ꝺ���]�(����x��'�n1鵽WN�ی.Ox��#:���X�Y�H����k���t`Y����&n���������Ί+��]{:y�;Nq���/)�xrZ��*p(q"�m�k. �hM�X'���:����t5ql+FyƉ)�zm�n�xH�X���;3��+.����+z�\��D��G���B)7t��F���4��V�������a�h�i���!g�C�����ñE��T�%��Dg��!�2��c�82���x�9_�G�8���������c��*q%\J��n|(����EN��-�&�i4��s�'X��[8ڤ�Z��oM+��~,о.z�2D%�;q��>�����I�^�����&kc���A�jd�v�P�Q��LGyʰ��<�҇G��	�~�Q�@W9,pu��,pĉ�|�3�Rܰ�98%	{�А�	2\ybTRJ�l)�]»#֌Z��8!e�X�S��Ds�5�IN=04�7O�c�:bDZu��Fb�}ْ\<��0x>4�g4�N�ԻPͱﭥ=C4]������j���埿5��Z;��H��Z�O?��G̊,y��[�!�i���D a?�1y;��Ze��JJctR
����1S�4Y��6{`��~q�5�Gx#_�:�J��}2��4s#���i4�:e/�;8N>��u�	g!|WF��8ߦ,�e��\�ۚz���=��L��J:+��lqO�T��n���x�U�}/�<h���yTg8��%3R�A�T��Vb��n����F����At�En��-��>	
1w�s�@e�ɠ��M�6X0� 7�Vl�����I&�'.���gF�H��/�N�b*ڨ��g��	P�H�(�֖W�&.տOS�G���Ad���CF�4�	X��]��t4���^zY�g:2���2��26`24�օ�������`U�Ϸ��}�][:�:���T�?P`|H,��jn[���Uu���-�����e���^c�G�/��?�r��Mf�d�
�&�i�X�������ѧ��a�"�s$z��)q�L[�Zq#�-�G|X-e��/F��ߗ���V�o.�Yb��8V�XK*�'i���2��D#�܈%�Z�~]z�H{y��Un4N�aTi�U�_�e�=r8}�_��E�"��m/K�Z,������H/�k�Q�oR��.��j*&R�_Яmwc��>SV*�k	+Fz[m�R��~����J�ꉱ��}��}&5�Xm�'<!z����BB�`�.�P
��ѝj:��ީ׵QI�3����@V�Q���+�`b�$	|ܩ��������LE<��_<k2bJ�ƬEZ8O�q�_�!;���-��'�yD�8G�i49G��,Yws�7s)DA[N���K��E�!�b�w��{�
i��@
���LYT=�կδ� �~��*�[�5���X�Ws��'��&���e�}��� ��Sv���1�:j`0��Ɍ�U)��>>su�m�.T;���_�6"
%=-���̒�Ό�i����c�Gy��!t�����j����+�~��ѽ��Td�fѤ;��7R���ca������۪����z�E?_��h_��.��8���(���Ke�RQ=,\�
��� ��OS����e�g�.������d����q���>Z���A��UҨ.C%���B�E�d�K���~c)��6��:���u�|3�"Lu��v�t�x����	�
�v��
Y�A�Jz�| 0���:uUg*�3,)Ɯ@�ۇ!�H�{d��$T|^�L�]^vվ��Hu��������74����X�}�~��'��:&zt�����2䨸�'�G(o(����6�qxz9n�M���&5ā��a���.��#p) �����E"9,vn��������ٶ��.�Zw����r��Gl�ۨ4n�k[�i�^lwv�_�7^���w�w�Bޝ.��4�+���]>��/1n������O�R���`ߜ���G��3�ߎ�QyQ^L����c�?�������d?�Q&ټ@���������eS���gM��b�3O�&i�8$ïx-��,�G��ыUB���6�5?lќD����N�v�"���&�zxl2s�	H����Q��M(s1��^��.ڹ�ź�9#�[�יp�����ʷ-�د�� v�"�����J���ڢ��i	�R"Y�a�=>f �;��&C��݀���ث<>��i��A���H���D6�Yr�p���5t��ԇ�D�(,�V�L\,�Z_�§y��:�-%P�K����C�{6ƪ w֪�Ձf%ބ�Tzdd8����J3���
��l���ڙ�v����Mo�K�.��<C���ؼ��C����cn���u=��<ে��(�,Ks�ĉ�	y��A����T�}u�:���)8��E�L]�,���Ќ��2(�V���<�MY�;�fD �Z&%|#N&۽�M���1'q��m�+����=�~�&D����/�~�p�L%Vnt��7�_L�?j�8h��Yxң ��+^���J^b�;=���Y�E�ʹʶK�-V���{]�M\|z��G�������T��-��{��&y�MT_U̠��ڣ���~��/�� �+��j��e�<2��JhT�7rp�#OP�4]�<��s���Yb����Sn�\,��E�q���͗8��������f%�ܩ������{I��ͪ������~�kّ��mTN�e�h�����U�H�֐jjE~��,�:Td疋	��?���hjS�>�W�V��y4�;������À%�oӪ��(Il��!}�5����=w�Z�arH��y*�G]Pr��|��z��?B���uS�rm��f�wR���V�1�0��=*M����Y���%�k��ڽ�}�{����2F���7��!�=9�ҋ�������a4o.6	@U:�"��~
��T��eՂ�`z
��S9�Q%��,�a���yȕ��q^x�ɡt)6�̛����z̊���9J�4�ae�<s��L��*�;ˤ�gZ�Fj `�d*�p�$G"�@�J\�:�<}Z�f�l�-�&�7�}ѿyN�<���/H�5s؄���n\Ȳ�u��kq�$)�C�-*�Cv��4�=� b�atZ@S�:����{%-OK���ޢ�ǡ
�bAR�C�5��;G�
�NN7���t�q�?����	[�-;[����OK�#���O �̊����ڟ )~L�y�%'Y�Qs-\�f�㮴@G�΂L|���8O֮�a�4w���� ���;�5�|�a��?~���k�%����܍ �9��2�F�f���D��[�D���\"(~￲�?�i�)厥�b���_L�i�-���S���E_��Y;D�i̖��>X��ܫ�ٙ�Z*��6�ִ�)��F3�XI������m�O���R��G�[�X�d�l
�頊3Y-�+�_ dM�$�U-�g?�V�TC�6�q�u���6*ܨ�����@>�9�W�ҥ�ܤx�/C���M䙁|���Z1��=��u@%�3�ȵ�zZ^�A\Jx
�P%����QB��l��
>��r6Ge����$�IdiZ08X���sd�p�g���ҳL�\����+��V뻆G*�&����u>�䥼�!1�u�s��u�Q���,P�w4�u�`,��8�K��0�J��q�,�pT��;��=���+�nAᑪ���9��w�L7�f�r�#�^����(���1&&��z�%m.�9rZ`��l��B�^�ݐ�3%�L��p��n�s9%�O�d���?����M�����^���%`a2S�D?5�OL�p����^�v�$��?u�-	�0W�|l�#�Ji�I���x�F&҆\'�0��V�ԃ7<������󀗪��y~*��������M�_��Vz�������1p?!��G��S��PI��%�f�jx�&E���<�"-\�Ԃ��i���Ҋz	
���_�X�p����f�OC�iܤ�8Ķ����U��Wv�#
X�j�M�sĴ�0���4�t��~��~B%���z���b�p�g��ϔ��k��K�L��|Eo`�ԝ���O�L@�g��|�I.�,��/�^&�
՞#�ǣ��x�p�S�e��_���?Z_��9O��2Y�k wa��溊�=r��(�qºb9��|ch$�ϥ��E%�~L�;~*�Bn@<o�������3B�\��Y��L4z��sWb���>i����]�<қ�I9i������>H]��Rؔ�qLbS��zګǝ;#��qp,�������cЇ��Z!%|�s��$��ї�d=�����@�l�C1As\�=�:�-k��Q�^�tuz�P�K�+2�X��+� 3y@ʁ���M��$L��CZ�OH<e��E�v�ʀ~��.�K�_���̇�S?k��v��_L�m��۶�v�G�I6�'u�^�1��%�N�R�o�	���C��3�k+�4�G�t �u�xqُ�7~�D"�	��0y~JB�@�l���D"�2�>a��?��w.��7]�@�]��y�׈Iv8�R�q���(ƦO����PR�Q**6��j#l7�!��(��TJqJ��,���fŜހ��?�o�{�6E�?��u7����[�1A�D����@���6J�3�^Dj���2[H\^�䌜D�p/��Z��Zˁ��qwPwk�K�d�;D��$E;l"���t}��ow�����]�J�q�Q�E��}ʿ�a�����uʸp��w�2���	�3+�gU�y����k��PrSw��D��^C'y�e���*lk��H�%+�ԩAT�"�(Qϱ*�P�NB�~7%�k������.��՞ 
xM����Q/	͐q�=A�H�Vu��~k�6�@���2<���QJ�m9z����d"� �B�p�!�Нt&�mӺ��;g���3��`�U�u�p�����	#���a'˄��'��قuc��tN�M���B��NQ��gQ��v�5g�~RN�f14���d�����S�$��v��'6u�� "��̮s_U1�t����ɩA��h�j��7���%�)��W~�\.�s%ޢ9%MVTY�m�����1c�_X���K�?�a��?U�ì��!̰�|���P��P|\��S�r����#m~`��/���nC�Q�K9ע�>�Cs�H@b�MAX��[�g<W��?J�}G�p60a�OY�E^�Єq��4,���AՖCMr���'��o�?�BK�����no�	u�.�����CĽ[�9X�[P�tC{��d5sJF`tqJ�`#&����5�cw��E�_Hy�F���	�Ww�*tT����Np
q'�4d��"7���Y_Ox���=�	��j
'<L񲜐�]���z�'Pp���Ak,�91�:�8CS��ayt�*� "���o�_j�a��5B*�{ �"�0�>(D2�ط��T�F!� �ӣyf�-�=N�)nܵO�C֮���Y��9�� �+����$*U���z'�1��X����T�G"�F��UM�hRR^x��*�x<B�:4��/!h5݀�p�v�<�/>ؖy�/�����34P2���4�(#^֧W`�0&W�$oĢI�uq凿`�H��-)���l!���z�A,$g�nى� �Ƶ��.ӕ?����\YV�N�L5��1�c�GOCZ3���gt����F���������i�d�5F��0������f���ٽ��<��.s��g������OCPh�3�yL���Kܻ)����.iʆZ�%k��@sz���}�nf����@X��m]�y�G\�&��m�RfpS�u#[>Ge�m6�yo�����cL%��$>-�].�ʁIѹ�N -#�X�e���)�ת?�M�V�4��Z�7���a�F�p����f)iJ<�Гӧ�D������Z���YH?��)�r�G�LR�#�q�tj�,w��>�|��2q���TO}�{��1��T$�7'DcuR�&��\,^G�a�R�9��A������ͨI$*���1��p�"��wT��z��|���:��HZ�.-Q�P�`�1�l���l��h �z."�@��vd��!s{� �*��;���(���<��h�R` 	%6�$��<S8n���H$���X�ش����3^�"���>�D���i,��e�����=�yk�]��� {i}��ůA)�`���T��j��޳��H����.��G�>��l�M}\7� ����f_�8R-���`��2�χ��vN@`0{��I���I�+���عۂH
O��'t�B��N���;3ayߧ�B�$_�y���1\�zV�\�)O�[�"�hknA�ҨG���Fd���ђ�;T�bOG�n�D!���z6u��@g�Ps���7`��%7�������k���D���1�yZ#��]+�REӒ�s��v���@��[h�oU�L��(� 
�4���#F��CC:Ez��x��JN��*,�(��O[�Q�h�Qs'��A*z7�t�`��i�Z	ө���	<�]ݞ�}Ы�ל����?�Ot��1�]A!`$�������L����21��}q\�m��!�$��5�I�g�LF����
I{��F�.�a����y�mEu�t�!-݈bhj�dY���h��d�N�k{�+m0D����;R!���&jk[P�@�a6���E�
�豤5$j9��E�cO�oO��V��Ft�`� P��f��̗�(�l�U˔b��u���P���G8����eo%=9�z�Eq�,���	���úa�ɗ�ܚH_��A�����~\����I���&�e̵�3ǜ�l�o!Gz��oC�>c����! ^���}7Y�hq)�~73F�Q	����*n�V�a��fkY�� �\��Ŵ��|�@���r� ��E
!IYS?�N�5L/wR*�>�ʯ�V6�p�v�Fe1�&�@��Z&�X� �#g��rZ����P�yv�����N#��{E�Ni�׭>�7���#���8���59^4ǰx^�A�x߳>0��7g�1���V���G�w沅D��g��͎.�GL�ƠQA�W�ٷ��M�RڶS�X��:�8I_S��։�|�$]b8��;��4-��]9?�C�H捸0G7�81��8a΁�,%A$0P�ަЫQP�"bΧ,�	9���-��"n��-`�M^0��Pg�3�,�������R��b��r\]g17�5��Ⱥn��@k��Ec����C��`�9�O�nh�o�Ӱ��"R���>���7��tU�N��㴪�۵Ǯ�	]��4����։T��Z����K\kT�������hTڜ;)\�ETv�E��ƼU	d�DJÍ����5#s_,�y��S���X��i��WG_���C���@F�k�!��"�ۄ��STf>������e-Gr}k:�t�3%I�K{MS9��8��v3r�ٌ���Z!ѷ8y,۠�!߼^;��6��2�
,�ܡ�Zu�?�G�tE<��)B�'�y�^yg���=iǼ��]��Ffn�][��7p�*��g��0_��w�b7O��Pk���V1~������Wm��x{=;���O^�w,�K��?@v�|.Đ� �TW�Ǜ�@�Ҽ�᭲ej,��\Y�k��$u=s�Q��T1�������i�'��dK��ԁ6��x�T���5� ;�tD����Eǂ�}i�Ks��)<�&�r�=�3��'�v#�_�c�����8���� ׄ��fF$11\�
(V�P0&Q�Ճ�/GY�G���8E*8�o$�i���N��*v��i�ql�S4�<�L��_��-6�S���,s�)��s��~�Y>��	��4E�U��`�"�y��VR���Şbw�Q�c�����~�Q>	{�����\+-=m���Ʊ_�rZ[p���D�j�B������|%���:�g��
�"uŴ`�:��)G׎��i�W�,k��q��X���nz��Y���D�y����^�y������#Ńd}g$]��NY���-��@+_�!�P��E��}~����Nf����1��:�a*�q*<~��23�lp��G�r��܁W����"HDA��dm�<`��=�;�B�quw��� =qW�L�P�����P<�v�rA��fP�P�!��Xڪt���p�׿��u �:��GV�$�t�o4��X�n�P�Q�(���$�!��ڂ(�w}��0/�3#3֎c��L@�bV�>k��K�%�#�ߏ��.�`�YA��h"��t��ҿoOAm�$x=q�>��/ذ�V��G�0��e����>t�{]��i^Na�
3�a䁜�[���k�F�T�����r�K	�B�uP�2��ao��>��ڭ��G�r݃?��|\'C��#����d��=�t;ͮ@�T������al��])}��)�>��2]|�
!i��@P��Wp}�Q1�_Ƈ�����p/jF�5�:� �x�R� �w�jdc1K^g��������u{y�d@��>*��ӏu�S8��V˫zC��'�B:@
lV	���@����2� �u�=���	�W�:>D�$��J�����r!��v_8����1�N��.t̾�|�h��O��	[���e�>��o��oς<�^�0Omi#>����d�Hw�X9�Q�д�SG�(����Q-I9zQKkU��+V��nhZ Md��k���r�����7�R�X���)�4�,�84G�Dt#U�J,����Qq�����B])wh �q^�U�t[�-�?VĿ��Mޯ ��Q\�<���Ë�g���78pk�o8+2W�J�OA�@`B���D�X<�]-5���蠄�j��،�)�1�q�9-W�|$��d��05��F�"a�8�\�S����N0_`�?��: ����j�^9_����a�� )6�4G-*������dq�s�#a>���ì��myh�b8v�+�E����]��^Wq���˙������ɟ[�t�5�iQ��D�HQٸԅ��L^��H�@(�8�ǲnK��&Y�|��Qu�jVr�/���_�`z�%�T@w��8W���1I�uf�}�қcK�NZ��oQ�,�^�&j�8Oe�^��4{�����Yl�B�C|�rq+���9�*�C"�=�;9q)��D@��gmse?�]z�v� {g�ŗJN�Uq���$N
�p��&>.�y��Mw��DUG^��!i��ñE���;V�����e-;SWK�������~��(�L�5rE>,���^@�hPf�%_eҴ��k2�MQ�3wV���e�E��Wf�04'~h���4Cόn�(��g;?i#?at@�R�Xm�'���U(؛�,6z����@d�Ms7h���D��]*�y�A�X�g7�<�����y����w�}*���k�0i
@K� ���d03L�^b�(����l�s)�?���e���<�n��-8Q�}2t��f�W�&��h<@��Ps��(k�ԅq��i�l������%s�31$��ҥ�#�J�W��^��䖳W^�Y&�ZnY�#v~�\~Gg�ǼH�ѓ�^Ǎ�_�"��J.E�<7����	��e��=Y�?��"���Ѿ	�x�i�f���,j���7���x�i�ƨ�b֔c���P����Z�عq�,��	�;.;����	�g��םN���p�U��5�u7�gw ���;��7Q0��W�{�zwl/6Ӎ��Z@�iV�p���O%��n�0�L�:�؞}�.�i\���i#W"�]��Zɟ�ܤiK�r������_���0�reX��ٮ��(�S���ϴIy��:�\f2���kT��N[�L��z�䦨	\j�)�2������_��23�S��?},��4�*���3I��Rq�u���+5�j�,�!�>�fL[g
��y*��=�z�k��[��\m$OyW�\h�{K����TǅN����m%7����z��,7�[D�����~R�d�5�T��ؼ�>�	6��~)>��4�HZ����j����ˇC1�'Tn���zM:Z�(m�""4�眐_oԭ�A|��\��ʹ�*�L���9ǜ���Ī�_�	���2^�����cm�޼������k��oA(L�vᆽ��i���׵�����o���W���dNIk2���=c�\�y�Dr�Ӹ� 6��<���UGTRR�Mec���|	٤W�Y)����Ȍ�������\�YJ����W�(���}�uT�k%�#���7�Pչ#k�z�mb�N�xRj���Ȑ��b�	��J�c�yI(eQc��R�ɸ�����`��/e0���������!|�4 z�A b)&��q�b�|pg����AS���_�"^_�6C|�.�w�U�����wdޗ���`�@�n�y#Q�y,<�eX�"1���2�p�ޣ�	l�;��_G,�����i �p��2`��42[����~�ԨH��ٸ��;%%�-2ļt�*P	o�e?UM�/��8܋��ȐpV7V�j^�oD!�?&����Ļ͔��
֠���f�a�����,֯�EmX� P~���vش���v�r�xZ����^���5�z������>��]_����4��;��t]����Ao,���L �X�2`��h{h��׼^�Z�7KZ�$������:��b%�_9��U��BQ3T���1r�u_��<�����*� �b�y���.E緸V��@��)��Bǌ� �Y�5�!nDT*u %�c�֭�+�Y��@��Sd>LڍX��h��\3�X��%T���&�n�H��_(ހb�^�i�"�m�%��
=a��]х	����DRY���{�u�$����5$_�}��cs��)6B	͆1��6D��p�m���`>1�	���CP���4��:o[�S�8�gP�z;."�ޙ�d1f�tQq{r��s�MO;����K%��{����౜����Sg|ʖ�H0�gIi���J�wN� �hP��¦�C��Ց�Xq�]�8�Dl�bN`�i���e��R����6@۞�i�5�!�V��|�p�v�!���'�/T�'LY�+�gV/i����2�]�����,oa�{��$�y�4T���H�Q��2~�h�O���=�G��ĸ^(t(�ĝl|��p�����`�k�L|�V_�¶. ����U�1���r�4ʫP�i-�t�l[�$��ڋ�ޞ1��l�E��?Kt���_�]3��@`��]��6��y|�[����KB&�x�-޵��n4Z���Z-�$;�U�s}�J0Ӗ4:�2��3����K_��V-����9j���>�RX�����r���_xL�����!(z)p����P9��E�;Իf�tV�m�����m��R�
C|K�9��2�)>�	W��=]ϯrHןd�=_����{���}"�]��k��X"*��cδq�cre�E8������6]���u�^�e7�m�ڋ|���!b��\�y���2��H��H�=dϯ{(�-�E����Wԗ�qaړv=9�*��Gk쥢ae�?q-�o��<�;n__�JPV��M�$e�9� T$���䛝�+���y�=�9�6%g?����8seB����B�D�Gc��t��8j�"[#셆�D�B.��h�Ž���|,�FE��$ "0Ayğ%QȬ��Y%d#G.8���Ľ@�c��j>�� [��8A��֢�[����+���	���0��iH�G����-�2tz��K��ͻF���G��^ŉH��������Ͻ��	����3�Z���W�u�I���hV_���/��PF)�s=��f����u��mh�����Z<׹.p�(�𓏠��ҭ��0���{��IT�+��sT�A	�#���ܘ��ߠ��3��z18�.���f�D-��d_e����$��{�c���,*_f`�����ą�.����-������k��[��p��M9سn�%�S�6�H�\dL3��^6ܝ��H" �e�0�r>=y�cv:`�;�#C�ߪ#X�U���������7ⲝBd���H�p�x=��M�v�\_��Q��}��ǌf
�MnY�%J�}��UOP(_gJ��HƁǔ	->�%nS�=�N��
3��)���q�H�źP���!N�h	���:�Y蛶��x��@U�0���")(xM��Zư$���;�$W������H�<S�Zb�����k��̫-5�!|�ɄJ`��2B��ZGro7���J}V3��`&�wC�{<�ɮ�8Y!77�Oǈʐ��{�iJg���| 1��9���f�u�V��D��C���wlM�f
?� O����,w��V�ߩK���=팽�e�:������S�*|`jj"�(u���	�ԟ��[5E�4K�)�U_��I#d�;?_�.�޿5=L|�ĳs���?v�v��mx�y��UL��E������W�CKO��S@�`��;_��A�e	����'�����=uT/}�eΰ�u��&D�n�͔i�ܠQh4�����	�t����\[������
�B�gTvs�XFE�V��U�$�X��;;Z0y �AY[�{�z\=���ƛ�-j�ٻ/�o��=Q�N���5q���g��MD��.p�@�O*E�����DO n����%5_�s���zt&�0�~m�IA�	�^�p����Y��Ǆ�^�z-\g�F-L�X(9ӂ�j`����$9�@h��O���J����8�F�I��-�%6\W����/���1r�����]�je#��O���ݕ|����{�E{��v��3`57���gL8�-jA<���̮����z��mP ,`��qBi,��(Z�'7�(�/�|jr�4+2����Dύ�y�T��<��S�X6�q�:17�;*�߽�������25O�K��S �����#��փ%�f	�Eŉ*�c�w���cj���B�ݵ�}�TS_a�H;�i 2�,�$v
�I���b�M=��`�L���Q�� U��_̜�r�/Z�Õ2�E�͌~N�i"�*,�{�����}��!a�V�s9��P{�����;�C�-T-?9����U�c����g��'���}d�����W�a�
�����@3�093�6�:"q�v�̤vcw��ʰ
���F�'��T�t+���:2>�d��>���̈́����I��q3��Qx�	�tE	��éos{,JL��Eg�	,����6~@y�P��_����)j`\�֔.�R%N{+;t̕����ĵ�4���fJ�T#*x9��{��9�����ݕƝ���܀��w�y+'�3p�5٩�A����v~��c�"%Q7�Rs��	4ka�T�zI�|�3�aB�v�iWS�v���6��g�B;&U'	l��(�a�kٓ[	����\��ɞ<y�H������u�x���ǿjS��q&mA�bO������{�$&�΀v��^8 g�i�R����¾S��tBP�&��=�ڮ����7���[Q�-���-%>8K-�۸� G&Q_nXo_�C]�4h�+��>�Lcl1�i�`��Th6�2�'7���f�5�	���j}�j��dVx�Yg����Z>��?	�����3׆����Z2����0i�`"W~	r|���]�3B�2��?W���N��rb�?���#��+p��?+-Lg�&�%�h �D�X|��#�����?"��I��EW61�FxS�-��~��Ej\���^��3��Q��}GD����&.��2���@Aq*���,z�M��k����^S�e�[P�l�f`�hC�Mq�y���	r$�׆�KA_�����l�.�1�V)��~��S�9�nq r
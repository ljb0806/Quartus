��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��YOf��������Y��gP&M<>Q��R��:�d�y�.0t���/����K�����)w�H��D��]��v��ԅ
aJ��X��w*������OI"����P��ʗ!�������M��i�4	��M�>���C�Qy����qs_�Zy�͑�|Y�7f��T6�7���J�]�C�
p���ϭtV��k����1EE�ţ�wT��|�:s!�K�=��͎6)����%h����|��+�`���j?Qf��k����F��jRh�ߐ�{�
F����\<�L=q�^݌\%���m�ԌIZO�*|���V�j`i�~5#þ�CO#p�sp��z��~:��NZX��6@�&�y�}&���6^w�cBYg�+M0���NA�{�%�Z�^�{{x���T_o��%}��tu��l��w�=}�S��4qx������_���F���J?[+m�d��0i�{k���/?��|A)�wdV�u��c>*�,]��^E����@��uX����&��xn���/���"�%����&!����r\��A�du�`�Րnx1�� ��O��sH@:�[]��S�(�c(��Fc��B�̜{f�f�u��+��3a��^-��F�T�b����)}Q{<|�<6��fcp_��
4G#��!@��Mmx�����vH�ۭ��m�*������v&�òc��*��X���*(hco�6�jl;�Lm6Ө<����<Q��B�E�
]]�.&���*hE���:�.o��z�ʕ7��'mt�߻0��'�������6�k�~D�[��j������A��W�Cl26-���M��	$��a �W�Bz�y��~�ԣ5V+��2�]��}�V��S�<6�Tt���
"KA����=�E�S����G��F���bl����I�Q	q0H4�̿w��_���8]Pj��ʢZR؍5.�d{�{�3r�5�QvEm"RuH�"���%�T��� ��қ�g�	�'v��CTU��u��3�$���Ew2��K#*o�9�L
�e��]�I��Ķ��ƊJ�ҡ���;�̂�r���ѪO�ˁ,�*�;�� L4-�8e*�H�!���n\�ʡ�2Q���zs=3_J�mW@�k����#�aQV#�s�q�8च�H�DA1 EuJÆ��d mI�;�����.X�w�=ϻ��>Ȣ�ƛ��B/n��>�~z��M��"�x*sAZ8E����>h�>u����`Y��`M�W�"/���l>��Ʊ{�F�x("�5z+��ď� ��n,1Ӗ ���Ep�x��㹬6����j'����l�?�=�l"��G��g�"� >@��hsd9�"������MO��B���V{�	�ANi����P7s2�2C>2�G���o����>6�R[�o��*V�,���$�7d� �@*�#�C(Q�x
D�X�C0��Ț�O�!��h����wo<:tz7��8F`!�D5���
D�l�`�!wvR�Y/^�Nǈ�/� ����xhc��|B~�X1¹t|r:�ֈ�3\���/��9���{"���������w�w��l=���dn��M�ɩif�3�ȳ ����BC)�D�{W�m<o��i����O��l�<��vf�pA����~��@�Ek	�����q�?d���ߡ΅��
��
����Bz��U���h��wF��)�����ɹ�t�.ے�"58�2Un����*��V~�f�Qڐ3��=�e�Jl)�CB�y��F����x���{�9����0�IpLM}�AE(p/\��(�DX�"���cmfe��{�0�Ք��!E����
+8�~��t���V3X�}ؽ�S�1{.8�#�l�Kg�	E��Rf���l!�Z���޺믱v6�X�2��Fqs�4��t���
%*�]n��2׈/�Fm�
�$��A��*�U�\��|O\��ݛK�����	c[�*}�a�J�7#>-,�NCE���C�
-(��d-�d�Z�	ܯF^!��{¨za�K���cr/(������ �p�?й�B0��W5�¸��>L�rł������!y��l]ύBs;�d�4:�ɱԕ�#��Hd&X^�v��`�Og�砿Q��T5M�������o`�PI�8�L��,�Nxj�M!�u.��X��.:0s<[�zDb�h������x6�5�fDj�&�H���uQ�=(�C��rz���F��%�Ag�p���a����S�y������K���%T�	
7��V�|^���ǮNrQ7s6ϠG>�(��xā��ɜ�9Y�ZFs���������0�M�f��IX�-���]����k5��Q�{n��K�P�����#7b���K�?#���~&/:���8gN�mX���Q�,�	������ �30O�Ȅ��;LT#9k�q���8d �c3���k��;0� ����Ce��$�qv|?����t�\P�2))���k��bg�R��/�1���F�J	!Y�v�h�K�[�E~���|ū�2���gG7kCF/��$�"�*��%(��.Z|\��T��a&I#��YƆ�D� ��t-悴��������T%a��/Wٿ��#�X�_��������?V���9�&���+_�I!{9M���f��±� �')ڂ����+;�����|,���#��7pq��d�R\Z���é�ZȮ�S��t�۱�q�n�����{��ل��S� �Ymˠq`;��}�xZaK���8�)�wӟh]�.Rb��j�+i;B�3��Ë-&_�����
�<�!�����d��S�и�p�8��O��Ȕ�bO/�/MJ�33���������S	��AK��H~����-8��k[R���֕�ޖ�+](4��,Ӫ+��_����Y�;��ƼJ�m�L�������8�*�n�@o"K��f[IK�}�fo�nL{�����t���|� j�pʰ�X�R^����ҁ�@��55���,���&��uրo�6t [�^

���dJJ��C�U��Su����������������#��ؕ2���u�h��-#��:
��&���+����X�(����nJ�CBs����L�W�s+K�1��vK����V�m@l�,�Uo��#�Hղ���Ou%bB�J��x4�2wE����	��A%�z�{ /�����vY~K��3�dL$���taz-������P�Ӿ��5.N@uǇ1�t���;At��irܢz��Y�)�Q������Vy��k�5Bf	̈́�ز�+��Iy
w�G1��;�]�u�i�-3)r'FP����7�^Y�̯o(�5���r�l�*g��+���i��3��^-�a
��T1�鮲5w�t�N��ϙ�/C��U�$MI_�%��pNP�̠��d�c���z�Q뾪��JZ�]��,�F��ؾ\ҹ��ΠQ����9��pQD-�C�$�T���Zo���}�ɦ�䭣+���cɄGĿb*'��i.����i�tPzv�qKFY�,:9v�7��L&$6�C��W�u����vP�\��#����C��T���lM��>n�d�>6�qZy���+uK�f�
#�A�:�u�����W,[�N�#�(��]���2�`����/�q���;�丅vK�D������[a���s���N}���G��}����]Y�A��]0��I��6������,��,d��ln�����  P�D�B�0Y��E���Y|�J	5�x�T�
�c��uS0.B/�)����,�x��w���b��[Q^�r ��y�8��������>�M�W+����HD��x��n򯻱&��q^�]������J�$	�;ǐ�O0��%��}@���\j�C\
�����9���C���?����{MQqO�-��,�7�5��g:%ˇY����SQ�T	]Ο��*'��>�I��p��з,�^�3���}�.3���9}���o�q�g��B�xB�$�0&KnO���$}Ւ���nYT tQ��7#�fo�*������4�Եw�*C:�y_΢�M�|\sZ��&/A<�e�@�Ojny�swGdC�ܐS^��e�����i���=)4JI�g� sl����"���� }D-���P�zv�T�A{jH�5���Q+�TS35�
e��:����	bp���J��BF$a�_̜�1�Me( ��:5�-.�5�� n���;��I�^Cl�h@9���'����Z��(o�(��D�xf2��0��怕H�R�=�'=V�M��6���˪�yS4M�F���JAf��,Vu�Tk���p��Pe|�g<�άt�ܩց%FڛY�ǋ9�>Ry�a���@O���~=#Û��yt�0�����J�qx0 z��.ꯟ��t��fSx�z����n$�ϕ���*�J�/N�hV2qRx�����'HT�,Kק�J���N�0P�:����cҎk���K��Ѥ|HzE.�I�jɟ\�(ǳ_Q�ᝅ�e4`��")F?�W�l�r1OI�t�10�
���u�ğd�З�?�HXS���U$��%?G�KEe�9�a��9�zVM�^��-�[	�� w�W��n�	�t	#(R�����,��v|�^��>�{�O�/+��x M��"�B ~.�%��	��T_DYT��l�if�[Ӂ҂�~�c+ᙋ�M��@w�ޕ��i�A�ݤ��VE�V���(jv�f��
W_���F";fu��-�|+RKя=Kp�������ȃ�|��<�+7wm縊Ů�b��L�X�?kk�5ύ
�Un�JZX�F�\�c$�^�	�}wjA��}R����s<��t��SJ��3VN�6!�Ŷ-.�.HZ`�ā}�⡊����hJ�j5��g](`i'�hɳ]��>��B1�:�7(%l�'bD~Y�Qk�P�f!%eٙ��{8���o�}�^��P|ϲ�Ȧ�l ��@"�E/#R� 4�����9����@��e5%��c�����$З�d�>� g�b��W��XEZ�0'P%l~s��
�8���T\��Ld��S���-�19\�=�W�%e�h�nf���9� f>�c�S�]4X*�\���|*���Ǧe�]��D�O-�
��م�#)��H7���&�1i�?��VË�����V]���,�Z��;��f�C��´�h���������;�s�F��p��T`��"%��H��%*@��4��0�VGZ���l7�j�CD!҃��Q�2��}D�3��HB�z� *���f-zl@�lo���w�S
rm�$3�ڸ�Z�5
��R���FI�4�{��!(G%�z���j�-�ߐ?��z�ؠ-7$B��Ȓ��7a�$������2y���ҟ����ʖxS;���k���u!�s��'��J�$%(lv���DCY"��LR�-?@<�Tm���o5�V~pY!�Jȵ7Np�6����qj��~Rۻs��dC�w��.���C�tD���5���Ԉ�S�"v@(6�@&�F3�ٹ����~����ة�I�t��O� �U��j�� ���K(���+#lRSvj�K�����@G�}E��>�kő��ӕ�f�:R�}-�����y���0>37�6��r�ǘ�څ?2��\�ݧ��5���c�J�+���7��'vT���7����s��IG��5�!w���\�94�f	\ ����(��]��&�*� �@-�;���+Q>���Vm���IXn�%iY�%��
��֒V�B&�}k����I��
!$u�����$�X�D��s ���6 RZ��7�w��~�EL�s��o�fڪk�T���z�5�35e��O�A�z��ˠ�r��1���<�E�Ъ��ꪸ��pA r� 쓸؝��P2��~�+����C0�L����|�|6�:��Zm�J�Vq�4q�ZN��>��A�q-�>�r
'\'�g�����$��?�N�F~�I��d�]��KdUj�^�q/; �Y�a��y{�<<�t�։��R�W���~9Fm�掓-��� ��ߊ>����~����^Z�up#"#�r�Tѳl<��nHX�SO��T��aqX#�u	�Լ�͞*"^�[`v-#��D6�õ�/��Qﾙ�wS�WzH��Pt�R'�E��Iw̳ /Ce2�E%���!�VfRRbhܵ����'�8B��"��6[��3��î�""�%"�M��]L���rތJh�	,<��X����CѼB�#v7 �7'�[O��nY���4��wty�?�F��0#�9��8C��m����h[A��;�G�kh�E(�X��
Uz��c�df-і	m�W��LRM��Z���m����%�ك}�;<�oeg�rR㥡�A��-6�y'��xC�*�=`��V�������@Y�~��?����8�跄��3i�)Ⲯ^�ݩox��cxyT��	��5��e���$8�ֹ�U�i��OT@�C�$�[s;��Cqa�2��Ј
aƴʱn�������$�Y�#��\�K��2��e�j�Ԉ~��.�}����/�8VM�)�����gU��%�*q���u��>Q��@p�r ڈҔ�R���}�nT���/bu� ���Dl����1p,9ua��+B����5:���weˏ��3m�$���[Siy���� ��2�`�V5�����{��щ<L�(�yl��7am��^mx17�ZZ����0ҺP��Z�'��vz�p��wi�ҳ�A]W���I�gEح��&w�2��@�\��z��Ф�ؼ@��#��y�&�ޡ����.��-�S� ø�8a�fpB��"Y�h�C�<�p�7���[�1�X�������M����tˁF ���g����({gO�P�\S�nm���̻��+��Z�d8�yA�%�2\��q���eң~&���#�ˇkČ�t�V�R��w��!��v��j���q(���M��ǧ���źcۼ���E�q�)�|�Z�Z�"��=_k��F�f�.~����u�=t���*6M��|����Fp��!ӉWr����*T=�3���3��m��dz��X�F��ry���PF���h�h�f�ǣ��oZ4/�l�v��H\K�;��Y��Jf+� �r������dP&r7����(��7s�g�}�j�mz���;~��4�� eV�r�׏ۀ,T%�U�C"�y���,5�Z�-�F�a�ܨcѥ;�Q	��o�nF*-��լ��"r�5��qu�JtS%�Ӝ�L�q[�Aa!�M�����h%}T�|�j��R+s�C'����6Pɍ҉�� ����Ԛ�+E�a��b��qJ#������A^0֕3oʍ#hM�%E��1 �غD|�ر���4�,���k��S<����+�@��'���z�mf�֧j���V������_�5"�W����W
�l8�}�=`�Ēh=�h��Ȫ�(�<a�x�_Leu��h�ᙾ xd}D�����O�ɿ4�(^ ��Z��������lWC_z�R͔�u $S�y ��kؑN5�
������Sd�&���T�w9�LW���_z<V���T$B$ l����:����d�ƛ�k2(|�	�О������ti�<��ع�|戤T��a}�5�z��W���FM�Z��wT�, j�ۚ^���yW�_��"km)H,�QSʟ��<a�]��� ݌~�񾡃��+��nZ�iN2��6�[9VȤ9N5��-��X+��p�~�`�p�� �}
���ZZ�� 
T��\�IOI����X߹r	�Z����1����*�9Yj�Ī)y��n���*C�����Y�ԉ�FI-_����x����F��D�ݺ��D���=%�.��&����*&��π��?7j��{��Ft�Y��d~g���s��G����o҂Ɗ3����K����l�0�Y52��דL��)(dMg�!P^W5v"@#�H;Է܍!6RW�U
����6�zό��������
 ��:�r�O�/ ���z��1��p�,�4PtD���X���U>掾�35��X��=;����G��"��L�a����s�	�k^�dj�ُ̞B��  ��� 讒�,�V�D�������N˼�0�;L����H�ݵ�`�>*|p�L��F���ԡ�.���I����m�(�z�����љ�Cm9'�>8�S[��&���l�C���
�wm]�9"���Շ˘6洴VkUԟ��-CS^�'�6�h;����)��k��<*��uY��p�s�+9��ti�͒A7��7ڪ�cX~g��i�KC��2Aމض�� ��<㖯:Փ��ڥ���ʳ��0}�%T�IʋX��m4�(�KL%�˦�?@��9�싅٭q/���A�I>'�s�[�'���yF`��	�fz�+9q�3Qg��~I��f�˖�	J���3���J6,�Q�#�&�˖��HN^�u=�	_��ƿ�FF�@��(KH�2ء���W������nRm��3�|Hgu������a�/%��Itֶ���:. �9��ߥ���t����� �����0���#k��fhww"�+Y�P^��a3H�a�J��_�R��)����rN���j��\�CQ[��^�35@��BN�^M�}�N�V��f�����)a�<�E�sR%���� O_f
=�K�7Ь��B�R��O!�������@��6�r��1IX��C�)�v���>AN����23/CA6��-,�?�������D��5����onj�N5�[g. Mj P�W4�"o\M�O�P;�~�3�\�d�d�g�'�E�!� �-�J�_����^!_E�s�/��o%���#W��'�j /X�)��hJ�+�TF�����(�K`4"^"iGl��%HP�iU&r��b�G��t��׃d�F�m:�-���MN̒�EB���-�ٰ����O�R$4���Lv�8��ژ~;��MW�O���c�v�^�5�v�mI�؋�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��N�BC>4��������O�~B�R��j���1.&��%L�`�+4�-z��K�˹�֒C�@����<�;���W`��u���O*\u���D��~�WZ������3��.�ik83�~x��,i�Yu��8���sz�9V��X����/K@6���Y�D8S��n&H�Y�z�/���M(I3�K�r����L����保JE��r�G���h��~���hkz����ϸF���qN���3j�ض?T���o�Җ�*�-��jo�')������g,��������ۖ]� �B�e ��e����VE���o�\R׉���8 o�4=��ėG�xhܹ�qs��w����Q����W�_��ϐ��6t*�w�v��Y��Y�H�EobJ
Vԁ���j�Ɏ���U@��r�\�'mc5eF�֢PFV�B	��N���f��[��-��o��Dk�XE�v�����7�Z��qk�\|��H���:!�.81$�G)��r��Vf��]�DE�8_j	����ȋ��lo�`nH�|Hډ�2K�y]dRE��)���+(˛�a'��Pĩ���\�H�����1��ʽl�cXE��W��l=���ڍ��\�T�x�(ĠgmZ��� ��	��m��xW^hq��,⪤��A��>Pv뭾�l��
�5�;�^}�"��o���\����Ҍ���}��dize	�2.� ��Z���S(�В������uR+���� xg��p^ �^^��# NC�#�g�Y�;!S֨Nkg���a4z���Z���iuu�Mbd��q��/�Q�P�H��O�[�ҏ��&7�uS�U.W��]8(�k���/Yhzm�������ޣC �8��������c�IQ��{%.��`S(B�V��`�Ĭ�>Qr%�q����]�!(WM[�/H3�mK���L0idh}��Nۉ�q�Gʂ���϶�'��i������^� �z<ߠ򊞞���U2��3 p?$D���y/���#nEC2�|٧�`6F��A��ʧ�����؂RR�����S�p"5�J��g˿HRY�{��4��Έ��үA(�;^є⍟�7�]���j��٤wJ�GZ�+3;��U���X�9/a4�+K>V����%�c��ѫ��(��������o�-��rW.������Wݓ��b�TP#��v^�n����
߶u�o����xoH�<��M�7G_���˚�����>�R�����G��נ��������r��������� G�t�	�#�f"�A��	bb�N�&\O�(6�t=��tfW�e��0FX��ľ �_l���G��)>�h������Z���z'�����إ{Eܿ �26�\�"	����E�.=p��_�_����G��D�Q�;�'F�glz�f�3{kL�.����q��I�)��H>r���Jt��D 2���ӆ�,%�Wrn*��!�X��ٙ,�� �dUde-�2���ᰱ��W���ڞ�=�5��Z�8�����L��0��5ȣ�����Ho�&�1~؀��R|P+)�1a?-ʬ�	�M�ĻG�L��^$o-���L9�J��ԋWh!{��,�(8�?"q�^�3%'/x��4++�k=$�>��U���2�N�T�B!Ba==3����ɰ��L,3,����+&D/5'��B?��*��2�a��&���3���0��}<t/oy/�2>����C,&wŌp�d?(v<�� �l�~��$�R7>!�c��Y��'��w�'W���̞�ŽCۖk��b��1��XmS3<q!�ż��^ؠ�]�4�� ��z9�ً��H�T��8���d��O��%�wz�ZT��~oڪ�5�u5)��|u���::�������K��]���2ڲ����Q_A��F�2᫫$ߝ��P�M7��*!Cw�Xҭ.�*�?.��āGʮb�v��~?/���g�t5`�i�:��>WL�:�������H/]%��(J�4�J����~0��(l+Ҭh���êPF������кJl�+x֡S��Ů�5=y����E��4v����[�fd&�m��8'�?�Bl�:S��-�_��Zh,�"�}K�S��g�/�<ç��
�%*Gf�o��R�Ƃe]ګX�@8�Sw�-@�>����]�Ĩr��:Y����^o������+Di$P�_����6�59�8A��db��T��9�,E�a��w����q�P��VZJ�8�F�l��P#��|��
��urO
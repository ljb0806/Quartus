��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB���šp(&�e�
-(&d��R�ӆ�_������^G��xs��`��u�]�pȿi�����ps�<�#'oV�������Z*�C�*�' �8d��{��&0�P��ǠT�M�D�h" x���0�}��F`���̇�n��]QZ`X�:���?��I��O���E�P�yed�lHI��&^q�X2'_��������"����|�*��ix�O,�������L%��Jp �Y�"��'8co��.��<�R��֪����-��L�Uʚ7;����8eV��e�c��$�p3�a�^��$�Gk$I=q/u��ٹ�9�yA���	�@f������J�""��@0��	1�*�*��B&��GR7��� ����-u�VDQ���Yj6��e�D���pi�̰5"t���8���}_y������JːV��݈�_�țK���Hʿ&����-�͗xR��vۢ��Ǟ���.��]�)�I4�Q���Jm�����K/-�'l�8�B`|ı�&����;�0�ڔ�(�W���:�`�ӌ�?Ei�u�$���^�q"�7�#������|a;�uO�{@�	�#;�F����)��WL:�W	v�#��S۠��$����eߗ���z8;4�^�Tȍ<����L���T�3�G�UK���O�PՐ��Q=GV�AM�=��c�}��S�|T-z���W/vhs���J�xG�J��b�y��:�}B$�F@��iB>L9C�c���g<����G{�P��|������>|;vj���ٸ�`>sa�db:U�l��zM��iK�p��iK�[J�4,�CJHo{�{8�$�ɔ	� �`���d���%�&����siع���N�U׈fGx���X�j��4�p� �e&ޮٴ�9����Z���|���NY�/@�aGQ�!/��3[:)�5�yh/g��@�g���=���3M�
���p�OܥC�m�'�|�I�O�w���ED�l�GY�u6��F݊�X������]��r�Q�� ���P6��Jp�=�(������|����4E��-�Γ3� �Sv����+��]�l�������ըĺ�Ϧ1~#�]A���4Xhb���ŧ��£��0����ud:y��PD�k�-��{�+��;mJX�5,��w���z\&�E+���&���,И�N�h<��I-_�v�r٘���LR�ʞݚs�}rC�Tt^�GEe{k� �b�\� �n�3_ۂ�r�cW�V�����l�Ӧ��>o�6֦����vx�m�䈁=h��ީ�j�6,\K�~Tu���`��˾�3I�Sc.M�˗Ǽc�彤l��fy��tw�t��?�BF��0N �Q	��Y�5ة�[�d%�u��3�N���:'?�������������+�9��)X)�N\0?�A�g�6ɕ\[� ��/�|gxsgn�(��Hd���SX�劤�Q�=�L�o*�"c^�	�(Z���	"���P�ļ�����a�T"��~���g��	��&g�X �&�+DYc�9O/��P0�Mꍳ��@��ș���v���'y2�_ ����F��U=I��3Ye�ѝ�8����ކ��!���F�1���{ؽ��'��P�>���Q�{#f��ɢZ��mJ�}GHy�X&��z~�x�[��ީv��:�k�ZF�s�f�Ŷ�e���&Ln�,��W����l*��V�fx�ī��ҴU����i�RC��m������Z��c����+��I��
��:�	�g��&첖1��e�:�oȕ�{nz4�,K�v�(�B�9ꚮ�,�W���� ����#s�Y�^���e���/�;S�L쿋yf������z	ހ=�0�����zD%Q�~�w�To�1����lq<����8J�[}���Ѡ��mr���86@�/�qcS�,y�d}�������>
G;o��s���1G�i����Z�(M�����9����3�H��l��Ie/k�eԩ8���J�749��3Z������Ϟn� �-�3����ژNP޶�${t�m%�Y8������������Gr��A��Vf�7�"T&�&L��l����A����}�آ�7]|l�Y��_hoH0�)KY���nZ�3` �*
���%Gp����K�S��>m��ʌ�Ĭ�7���y��#�wؼ��5n5Ӊ
h�Q���B˅[�K�
��f�D���er���/�b�����F[W�GH��_�<:�)��0O�z��J���t���sfw�?:nu�v�ò����aq�Ì�&4�8�����sD�M{���^�E5�%U�Rz���*�n1��/���
�f��ڣ5NVG:����u�K
&� �R+�������Øp�m2����A;P��2��?�!S	�,T:���t��u\����!������_Z�K�N�E�G$^r��.{�o�h�j@j�LH�ֆr2~�c��FRsiޗ[��]>��wr�kt�jIk��3 ���$��Fֽ���4��kȖ�8��}�M��K��(���3Ftrr1Z����������E�j�6Xc�
D��"����H��
��Z�HN��A�g'�
Lw�נּ=#/���o[�"@�� �1�c������	j�y'��[(%��T�8�?B�RY�׷k�+��Z�|9�R��9�㜪�W��j��,Q�mfX��ח�Bkɫ�������I��aS��'D�^�mg����/*@2[$L��#-:� TtBљ��6�2�o^."����?<���@�f���:�Ca�Fnp0��Z���؅����q[Z�9���m�Oc0D:w2:�ZKD�B�!���V�4p9�.�q<e/�0 ��D�j����U԰++�� �.���Jv����^-͔-i	���C���a:�r�qi;�_(�-�t"�NI��.C,|�:���	1l�+��E��$�� ���ʦ?�Ob��]p߬p������uT.��|dtȒB	����q��m�ɮ,w�Ivy�f���% �D��hZ���h��m����h����¶g��jk[x9���c~I�.���¹�1I�(Y��<�Q�|�ң�<N��b9��߶��BV�f
B�D��^^h��6,�@Ц}۪�����Ü2b�t��to�4*��D{�^�f���o�&�V����DQ�$zoY�|�sԻ'u���Bu��ǋ���7�t;Y�L�9��\E~$WU���ޙ�}���p�9���⇭Ε����Yo���i��w�/B]��]em�M[)�b4a����1Ea��$�.�o䱔~)3[QLoy�6T�j��ߕGu�Z3�g:)�"�����3�`�I�9,�ߓ~��yr��4t���c045����Uv�H�h�.�4�@��
��➲(�H�ʘ �ڪ��B�m�|�  ��$d��!�^W��q?��c��Qۜa���F����`�σ6:[18�~]��-9RJ$�
�=G��o��9d���/'|H4J�(_��#(����n�G/'�Q��C�����1�Hv^���ʝVV�:!��oW�mi�&�(`d���lŅ��) n�Ֆb��d�2`T �5vf�I�7�kM��|Ԉ��'�˦��k�.���Xۺ_!��ں�B��lx���r��8-2A�qə�N�I�cɸQ	���6��z�X��<���{�����mS��պ�|�%��Ě�i�R#>T�+S��>f-�ڙ�Q�}b饵�\�]\Z��4��C���YP��B�ʉ��F���YE�;)"ּ�BQJ��[�9���(�vF��P�C6��P*P�ݻ�
W����Y/��e3ە<�\W���¿1lY�ٱ�${ƅ�[�@��P*L�ʺ�^1B�B��χ�3~�h�
�B���,�n��8٬�#=��OaL������"��y�A8�@��t��Z�]U�1"�^�y�Ef졖���S��P�4��!f�"�6X�!w��x
�@d2�<��O��&v��Pp�����*���H���7�s����i�p�@*�XZB��u.M1l���V<.	ׁ������w��s-�0��j\_3�ݜL��o/E�Q�|��v�>���T�W���g���ޖ�*�@r;e�Jc��t���8��9+�����9��c�9�8V|J��J�m��a��-��T<�j��/E��TL���^�)�<&
�06���0<KS���_*���%R�ފ���h�%���S��\�eM�h0��./g��%�
�O��_�G��-jx=��y�����m�C��Z
���|{�p}f	�����2���f'�@��M>�33���eJo��1)��E�vn�_�Q�5�W���'��qg�%��J|���eZ��4;wGEtMo��N�,Ji��̸`�1��I�0~����:;r�˫x��=Q	�$���� O�v&��p.���|�W���t��E+�m��$B��I#�]��Sk��<���)�j����_ �����=�72��\�� �Do�\yp︟}�u�0&ݺ{��j�>s��~�+�X�Q	b�<��d3!F\���#�
Vbn���wc* 'r�J$���+x7�;[�̅��a�.*)����D.@	���T�|����9>I�������9�  �`xUS���	������]���o/�ߚ#��#\�>��{X��^��CY	����沚��b;��l
=K��o;�6�d�*1k�s"�q� �t����5 ^?�,��Q�"j޲�W�w�i��!(׻w����nbU�A�q�cS����m[WH�
l]>��~��$�iT��6]�=�֠f���T]\J�Ɍ�ד��p	���а�����L���>97�ޅw�RE�kiq�_�]>��T���*N�PJ���~�/�������h;�`���y�1k]Ky�q"1L	B����Q���T��ԏ��|�t� �HH�u���@��y��.P�����$E���?Я�J��m��VAI�l.l�X�#��y)F�8z��5)&\���*���Z������\ q*�&���	y����k2̣���Ft�+e:������QK����XN�)b29�����NGCԄ�1<52�W+x�.S4t���Y�3��1n������(J�C��z&c����ҳ�m��"1��:5��'^�P��O:��K'�E4��y�o(����e+q1)ԓ��ԝ��n�X�k dژΕ�E�0�`w�"}�Y0h~c��6��I�R��⩟����ᦰ��	��s�aӁ���`s^�RlUۧ�tV��o���X�h�4%�*�Yx7 �e�Y�3�AaFP�#����MKl,�
�� .�dg�Xom�� ����K����Ǫ���w#�� ��1��Nu>q(j�G�&�
&Sj~#����\�]gl�p?�0ɀ��Z�G�ބ%Fu}�2s�R
5��~Dŭo��K�)+锊�q���Ԏ�~[�)��sՂ��cʜ`I�>+���|ǳ��3��l�kT�=�-?��/�O�#9u1���X��1Vm��/L�G�F#�<:�F�M"fi*��B}�Ak�ds��=:�$�'��o��8� '�Ԝ�ð⌂H�����S@��̹���z��k.����!��u�7������{�
�q �fH���f6.1KX��y��eϿ�Աv
FZ��W!���%�=�Y׶��k9���{Ng�#zn%��F�B\�ī������X���4�Í�gU]�C�
�G,Ѳ=����b�Ӿ̸�w�q���Q�Ѐq�37�3#;�H8\>����W���s����2�-J�	s�P�L��đ8+?�(��\/4�X�M�zPxg���(vޠ��%�f�3���
h�>�Ld�=�3�[
4q���IԚ�~� 6��t��(��H�D��:�n�<����W&'e��S,�rA1+�K���c��uk?e,���ft\jD���k���;0� ��s�#7i���Ƥ��i�씊Ȧv��z��Hn m�<-0��@���O��F�{�~o[|��������c�O��;���3 YRp| ���UEY�$�Z-�ƨ�k
1��r3L����U��6�4-|t�%Dm$��������@U���PW���XF3�[)�B᥅�N�L�����U�Id"�3&8F��Ρ689��g�"Ðil�5���I�����v��|��4�ȣ�v�C5HZ�D�%ϴ���%��V�։rM��������UD�WF/��+]�Wj~����#pq��tH��m�<�lE5l�����/�̇��7
����v&x�O<�!
�l��?(�L�u��%!�r��2w28I���Hs}�ǆ{����W�"�f�Ԣc!變g�LR%��Ğ�}�k���E�
�곱��M��T����B�����e����O}�Go�/Ļ�6��Q+�]gb�"f$*a�<�Uf��v�rGIj0ɶ����ag�,��2�ΐ�>b*�[�O��K����Q>Ƌ�/M�E��$�M�߫��!���JW��۱^#�b�<F�zV��X�(��5ڴgٛ5F�%��Ջƛ���l!\�INKp��x,�S��}�9�ʋ_-Â-�������o�~7"GqKR7��t��[�,oq ��I�ۃ�D��S�8������>���d/��eّ\۸cb�Bu��R(S�3�#��J�DĬg}R�$H\�TX����fQ��r�@����`���^-�oy�V�S�m��}lۇc��лZ�t�E�eȂ��'ŝ���q�&��D_���	�Nޖ�l����Ũ��11)���g�oSr�:^?���������<��I����d��8�X�0�F~̱������tq%BTDLl|[Ś-d�j��\���UI�p�(VM�R�5�E���5/`�Z`�m�j��9m�[^�,L?�s��9�����U	t�p�{��_���q7�� �V'�ji�_}�|p�����Z�d? 4�yGS�{[�w��X�$qs ��d��}{��I�6��=/>�ȕb���_�[8� q=��@�w��-*!˱?��e��p��e��xD����� (��3�9��(/3��7�I�wk8��_�=L��� ����,�	�w����ݷ�`=3��╙7s��
s��x�Tԃ�!�s�&�! l����M>��d��k���CB�a�*�V
!q��R?o���}0�Ag�Aݡ���vV�D�Qo3,I���&
هi%��nBcN�U_��ޕ(RO�/X�n5��U1 ����447D�5�e l� U9"u</��u�A �����u�9
F+i~�}��Z����ŷX��t��a{#�������1;5���(^��"b���٥�҆�P*�ԏ�KNh���M�|~6�$�=՘K�g���Q����VM~4�/�(���|ގ;*lL)ɯ���m�hLǄ��G��R��et��3��
��u����\�*��rL����7s��r�[Up�9���Z�pd	k�� =�+�y����3Ệ��eD[�0:�Ē��[��eI�ؽ |Ȑz��n3�U���̍,����� ���]�('�Y56ɡ���,D$��LU�?���h>g_�ja�����à��HG�c #
G*%�𻗩�#�-��{b����<�h?��{	h���|�AV�0M����O��o���.6�
'��$u�.A\(^��7�[���0E�m���|�>�ϼ�� w�aq�L����ɦ�{ų9��a�CLbM����%��#[ͽ�����z}�rf�6 <l�1"��좕�>�Yk��P�7���WC����5�m�\�w�����ڇ�E-�בoM�>���h�y�n��Y큘���U��V�dcF�5PD���z`��R�G
,���$�p �shL�|����j��R��9$��y<�B���#|�D���X�G�p��:i�s�Oj� 	W�:�>�_��\��'!ͤh�ܼ\}��a�E�7�Ĳ=^2Hb��y��6ް��6)�J%)Á���!O�)�X'���F�L^c�b^��[��q"�=���q���	�$��o�Ue�#��yװ�b�̃Zu��a�#��� c`e�5�XA�<� �e62�?��wā�]<�v���~��I!p.q�?�I��k�`��NBW���nĴ�1�KU��.N�`W�/F��&��J1�U�\I�r��{�ԭ��0U�Ex�������"��t��L�"_nؗ�ޠ'���b'l��. [t�&Dc�?�Ȕ��{+�BA�N�����ec�q�_���i�޵�/-.u7��{�(�`=�t0�}_�[))?N���T2~(Դόq$!u׭n��$�}E��_Đo�l�lu����,wv��?�6�|&��G��������/<#��8D�=�Ӿ�o�7��6��z�rR0��pָ�g��0�9QH�|��ş�,.��*�C0�|��\H(#�k����H�z�%��b���C�^g�u����Ze��3=*t^s�Vaǡf`���d��)��PE��؎��Ń�\1���#ۜd���R��'�9�����h:��n�����58����p���?���}�ﳎ��P��=L�@�`���ɊDmϖ2e|dR��X��%��<)ٯ����S/��n�|�{�����cW�x��(ós�Y�7�G���kۯu����#�>�7��ԻW�<h�_��VoK�]328��} �ʱ��4�����s������u�(8��/^�SC$�'s�I5)5s+��H�'d�������W.�1�����f�H�Nqv��A}K�N��+��Q���c{��s��r������py��Eb�D@��;A�������>n{�[d��=EGcI\�	��!�����y����3g�� �q����𱆝��F;��o��+�?-0��WKѾ/<~���.�$�Dj6������#����Srsĩ]���r��Wn:�p]���Q�#���i��s��uu�C+<~��:�A5:>"k6J���3�At);��j$4��b=�� �|�p������;�,-���P�����
�q-)`.�!: ��DF�D�Ă65���{��O�`��C5HG�� �-��� �mn � 2��5{XP�cb��r��׊Y֘e�԰�)�!��'�?���~�MBz��0% J������1Dc;�o�W�V��֚�,���>n3y����G��+�k�m:�u�9�)�e�Y<��}��W �R�}��b����\�e:�&m����m����Pf���Ph��vP�+�c;��9��,0DS����(.�e�h���_����7�[HGT��~_�Z�c�˞�GQ#�z�_YS�/�c�o�+^��_���(wJ!�!Q�FrnSC�yE�����\vf򚁢�T��{z����ΠT��12Pf�+�Ch~`�����yLҟs��)�@��ǻ�@��^�3�zQ����I��i�0A�h�.����=�a�;t@�_��_��%!�d�������ͺ��6ܳx�H�XQ7)��u����wa�Dȝ�T�2�������l��
�,���"��d/�x�䓈���
0�,c��oGL��&p�i��:f�D=>)��ې}|�@��+�)E��;u9NJ��*��4��u\���=5#��#7�@��S?ўSW��T4�D����uB��K�}�W.`��S�
R"�����2Eed%ISz��f��(�%}ok��R����+��t���)ǖ���]Ɲl��|�����S��=��8���U'ƀ�c���l݁�����.�Vd2ۦ�;A�T��(aqS�?��2%Se3ǆ��J�*��q&m�ZX�1��"��V�ũ��v��������iz�1�o8��^}E�Ρ�i�Z��/K��7�A�5'� k値�I'.����d��T���u�T�0���9��������?��! c;�r��9VB�{���#�al�7�y�'�߄��9੖��,Y
uX�D��w�+a����ԁ�é`�.�j>�+y}l��Z^��%oUQ,�~��>� �����L����ڋ�X]�F�k�xۥ�n��;C!p��:d��H��T��p�lj�3;�s��K��4��<������*����;���0Fށ/߬�g�C��Y�Tl�r���xۯ'.SK����66�k7M��ڕ��O��:`*�����0�'*\���N�N�N��ゆ:�fe�S��m�T@�lw �$V����(�X��b$�@,� S��ߡL�k���]|��9�ݎ��Ǎ���S���J�)�&�"@til����x�F���2/�w�/���Re���zb�|Ei�G�1.+�8�!�H1�C����*-Y�#�3���R��^gC�)����6D�jܓ���3$u�x_�Iy.*�M%�n*�=I����Û�9�ې��<.T �˾jc�_����4�7�0h R����Z��T6Ҳ{�D$=tA��w�p��I♣k�Wՙ�?kX���*��������	00ʝ7L�����ҍ�E�<��U8r����V�5	ډ��ә'��s�O`g�\^r*�!7� ga|��t C�r�ex�E���S$r��Ⱥe�������砼��!�Z[�{x��''���X����ڇ]g:֐0�Sfb�p\F��ɷ1�k�F�B6=m_��o�V�8$�Ul'�L�,�J��AKb��-D*���D)���+H&��T�3�ʶ(�kV�\��E��A�=�J3��~R�6�|̆�[Q�,��ū����Clwg����\Ϡ�d+���p���XG( 5����4lJ�(���}5x���-(y̦j!b"��|�\�UP(J۰`S ��|(ឣ��bl��T�)�1Q/ܻ���V3pZ���ǽ�+{�\B��Xx����p-��{:u��A6`g��k�u�?�o1��Wvꌩ&8^]4�W$P:��IO�k����ؓ�Q�p�����K`/�^�6����u�]����mU�blMh��
nv�6�#���m�1#�Mk�4VN�䈫}�vg��_�ե�[=��y%���:O�&�a��I��,��7��-���䰓L]�!��6ݭ<6�׊���xBU�:��q������-0��$��=�a�ȟdd��\Jk:�T��,�O�е��i�^/���8�Zv�n�"�f-[Ʋ�j���ԕ�/�b��uj�o �H�6Q��-A���=���;���D����pa$$Cc�-������#FIV�.�ZV;�v�	�V{�'Z����8���l�WFL����/�VJ�@�TX��&�24�`��J�p:I���b�s��3�M�"�ǜ�&:7����l��"u6�x>֥A��E�*6�7���@��p�=�Mm�b][��{�4p�󗈭<zD���(��DUS��$��]W8�}y�k���Kn�I!	�s;cƠ��D#e��ʗ� 曍��V7yێd�z`<�&�K�F��x��:%	���P2���L�J�櫓e�NH�G��΋�<|�g��yrz+m�qS��#~�8��&c�}`��O��%tZ�'��_%�5�1��Q���߹&	����Եš���A��5��>�\��܏���W�`p0��&3��,��!<^�A�Jޣ�s�L���Fq�X�%�rѶZ�YvN�_��t̀ԗ����*�����X�`���hC��s����Z�3x��6��>�?�0{�$�T9t��G������9�
�� ��[��]��#�K!�_�v� "�W��/����A+Ev�)ѩ!~��Y�=��p�9�X挻:����K���v�͢%���:' ���$�ͫ��&�Y/�SrS Q�[���y �SO��ӝ)\E�ϢK_1n��e��J���j����T+�Cj�1�*�pPK�Ǥ�5��Nf��M�z�~q�y�Ia�̄L�c��n�s/x	�Epi�cә璉SJAHy7��.D>j�A�?������ӗ��gj�)t�.���z����j�ۅ���%�>8�Gq,�4��K�[��tn�̿°������>/bh��fE,�f1�����}72�w���4Q�)�E�W+[~�Pk��{w�8�C�\ʂv�݋��HeV�.KwP��9{c���rڮ~��2c\:������ᘍ-�����(Q<�<��;]'F�VpN����n��EK��V�dѵ�݌j�x��rx�s���W�y[R�3�>� кݮ���
J�C/%FP��L�L޸�ŧ�,�u�ؠ7��Y��	�䨹c�ҿft���Nb�_G�>n��,�*���8t���{t��	$��aP��0��T��i��<=����[p�ә�C?�51~�!Q�e�ST��y�iUE`gj��Ն*�m\{��� �	����'�)����2���'��M0t�<)�O4:$̌�$�$L5ub��ҝԩL܏'jN�Se.�]�G�����L�E���&"�Z��;�N'Cb���b�|��_v�S|\���*lD�����(  �x��YW�ms�WQ������,Փ�c!~<���d��aφ'u
�ͺ��σ���*����.�#<H� �r&
}g�����<>s9^Z�1[-�Ovjs=^|K+&��y��%���*��K�v�Ί�ٛ4E�!G4�Y�̇�R���}��^ν%�05v�;��430]�%�+ ���(�Cք���2�(�m�������z����J���9�<G�;(�p\��Hۍh�k&���&�	�O��P�
O'#�Mx!���P���\�CVyJ��_��d�����8�X��t��O�"P�S�̈Fe:2�����Sv(�Z���/+i�Qt�:��q�=�ϳ���e)z2W/��l�,��n1�q�r�c�^~.R�r��]󀁯o���=^��d���O��`ꕾ�U�Q����ӵj�ur3n�����Sf�-m}ɣ`���H|6Oq+�܂���:{�'�@���<�&pf*��t�����C^���ۜ���=�M��,G�.���ct�{&,5���a�^�5���f^��1j��25�������X�Z�����C��24����[�,�Q�J4��*sV���Fj&ղ~��yN��SA��Ьڝf�N𠆦U\����R�#p��^Ɯ�찠5b���g�[���(��Q[�j�R��� 銢?Q���(�����J�:�(/��Bd�r�v�q��p˃'d�?m
Z�x(݄���/�hAgT�U��8�
��-˝�0����G��ٵ � m��W�t�]�����e�����cO2���E32�t��$28�Nk��������0��N�A��`EBsüxT(p���^��'ٗcR`�xu�[%��N^T㆛{lG�O��>���n(�o�cҁnY�K��'��<����s�p�# ��"���V�ʅn%]�>U�2���IWӭaeѦDd����;�}���ǧ�� �"!�'d��7-1'��%��ٺ
������<ڠ�@4m��"lM��}��_C��O�t4P��R�|0x����3LX����f��?�S�@�%�1v)=MyGe|X<��FF�8��S9,)+�~��f��we|b/e�آ�k�})&X�v���٘X�u��g�@��j>��\[��tڪ��¢*�4����{3��\|�>N��bB뫗>�,'��h��*=,1Ǡ��Jdz��p ��D��\��2���@q*՜�X�i�������Bm��y���3���
��&x���AΏ�Ko�����a��o�ް�݂�7�g�R(?� �ڤ�T�p��_�' OѣU��Pu�</:̧�8����_��'!��8��3��v`I���g�
sį�'_|��JnilP��{9Ba������Hv�G@�����f�e�Վ��P�J��T�}��R����Dӟ�Ѡ�&l�@o�E>�4Sd�S��#E��@�r���f�t��~a����#�ޒ\�"ʿ����R�3��$h~��h�A�[�L���h��b�8�\~��'Wi6���noء;�,�mT�eK��V���H�1~P�J&�gPa둞��~����= ��M���Z?|���VG|ũt�)R7����=�����𣚵�]9����DC�Ô��3~�1����f�\k'b3Y��(K��Xm�3W�eaZ�ZT,r��^6����O������ޘ腕�>e���m�p�vi����݅��������t�I}�����eOz�T���l�¬�k���D������V�S�d�8��/���&�h��\g�`���i�<�'g�?��K&5��u�Z��W��l��$���W 
�R��d�=X��t8�k�K�7��_�&6��ZL�_=�px����K��G����=I!�0��UWg
v��o c�B@	�+l�K�dF����J
���2�,�Y��O:8 c[;L<�q
�)|����,�D#��>�j�6�����I�����e�S�6�]7����h����ɸ�:�)t&�M��
��s���";"��>fYt�mu]7���g�O�����>e�l�b!zz��9���D�8�(���N�5�zcϳ��6����Z�W�m�s���ǧ����n��V����D������r��v�����\����0����-rmm���I�c��)�(l���̪�@����s,�W�A�c��u^r�qnSO'aC��\�16�|��:�2�k�6W*�#!}�ڞ�?U�i"Q.��k��U����!�a,Z΢�L(���u��Ƌ�����#T>��A)9���!�cZ��O;k�ӿ��u����d�9�ט��)����hH~���R ��BWO8x��]�N0��=$� ���K]�a,�!Vg���Aʥ�ʩ������T�������)�5\�څ�5-�V��a|�\�Bd
z���:1c)�`h��)@��g���=�	ӊ��H#7)d��I��cج��1s&��N����Gz�� O��a���p{лN�9L�4���_#�l�c�E��hP!Tl҃r'[ܩ��i:s�4Y�.���.�䡥fNL�"0'K���Z�f	�0qV�Pz��}!��ݴ�mXa�����3:]���G (�8vC��H�!j8R���^��M僼���3�/�ʛ��X5��dⳖC���X����y���*��x�g��9�kC�y���L[�t����5~�Q����S����ֹ�΅)��� f�W9VL���A���yM��6,�t�%Qp@�$��}�aZ�=��\U�!��Qg���2��L�;Ac�ÿqJ���^0#�H�H���RH8 |�i�PR�N��yMZ��/7�~��2��L-g�J��=�20�|��$~B���OQ���X�m�94A��@X��/�<dU����Cc���{+V�()N����l�Y���AY�pF$R�ι�x ����ăB��øмۘY�.�vwd��rW\v��+A�(�/mW��˃�ʨ3S�69Qe��V�??$�Ӏ�s�tq�)ER�,��5p(1�8��g��*�t>i[�*|�њ�"]ᮒѝ�gw���=w�L���ê;>����j��Yv�w�9NT�+�*i�Ԋ�ᶛ��SP�ڃV�"wt���s�:�H�Z'+Z5�֑ $nk���m���d,�<��_��m��0��$N���yb�bڈ�Z^uDB�/*�EpK�Q��/u�-����4V*Mv���8�U껕�!����&>hT�,<M��#Q���O�?�QާR�ļC��Z+� 	uG��#��;.�#AإV� �iޗ\y�\R�$D�M&�k�%7� ��mR�ǳz)���ب�DG��pe�a�d�
,UYl���y���D�? �`�,�`�
�������Q��*�.;�������4����0�᪲e��Д�_!�G��}v�v��.�l�P�۝��OH�`�/Z��2+����wJ��ݏ	a���%��@L�	(���y����`�hG��V��� Fy�y�=
�E�7�iK���T]���甸��o���B�!�h;��� � u�&ܚ7�~7/W��r�-
�Y^hK�ߣ]��{�6����C5����%B��f9�ȵ_!��`�9��<��F��S�@"���P�"��ì��Jv�iő{q�r�~rc����{8�؀Y�]���B-�����f"��#�LR䰈T�CDH�iq#�B!r&���$���g���:5\wM��3�f�]�o*�Kp/�/�`ܤ�{�̢���^M��������O�T�<�$ 5ݦӸ����Pu�9NO�bK=�����DW7{Q�0S ��{]:���Վ�U��%w�F�w�����o>&�E#<%�&=��a�1)��K���˥N�a��gZA��6�ʈ�>�m�-0�V���k�T�L�U!��[����
��D��\�����O�fRP�+���]��8�
�O�X�|�$�	�����	���=�|�v���xq	(2�m�f+�l����`����j?��9C�� ޿脽}i}a{g�������
~e�N�uLK�7�@=��I�+���_y��;~��xb�-����M'O8E�7h��=�B��Tp{`���/�	��=3.�l�i��EK��V�w����q�k��=@�&�
ě0��T��F��F۝p����0�8����&\���F6���sf��vOڐ<�����a�U��С��($��]@���x@c,��Nf���:ܺJ�V�(���Ó��ė���q�}'��c;��ǅ�+Az�kոVX�9�6<Z�m����Z[;Uk��5U�R=��;p��H��J�#⩾�v���C��}��
G�1���Ӻka0��MF߃_q��I�� �b�LGw����MF��u@�̭��5��~@��$�� �����߷�"*��[.IT��F��q�x�_���υ��F�B\��S���&�ǻ�w������q@K�%צ�L�ֳPp�5�!^��Q�� ��rkCv��[��j%���̖l�O�c.{��Gw��r�|u- D	2I5��W�3+�}J��T�"~U�S|_��>�`�]��}��#�@l�!��<+���Ԃ"��f^ZN$bڂ�F����j#LЧi������.�|>9΢��S�Ӊ�Ƈ%n������AqPR-���.������3�ܫ�+�s��S&�v�ԙ�%]���#��}����"<��*:��J�	d���M���qےJ��o�u��:
.N��W4SO� ȏ+M�2���X����Ԙsi�Î�7��Q��vT4b�M���"$��;ym:b7.���RP����T��H�DIi����'Z!���ǿd� T����`>�z�˛�
�C*�;<�ߊ�!tLAE��ŠZ�tm02doW���r8ӟ8j1�є��.C���W�v}��d/�
�]�L+���q��,�;���&ݰ\Ɂ#w���I1����_*��F7GkD���TT��c��b>}�uF��1!#�[]�i��,���M0��bpbV���e7,B�z̸7�>lZ�ծ�
(��G[o6��A��wǣ-:

��Ǻ�$�p�y��B�vL���L������HX��$���-�a)�����5]��]x���1~�������=a���\0���:�+~�X)i��ϼ<a��~����r���<Z^*�Ob��w^�!@�G5zP[1�����8�|��*,i�˖���^}�L� ���=�Ie��D#n� N�2RI׮��j;�k"mZ��8��j%vA׃�8W%��=^�;Nr����TF��hd�Zc��-R�Ɯ�*_4�f����&;ZB%�p�1�3?5���{�<�����B(��x�>�鑢��\���ՙ3-�z`��>n\#EN�b��8�r�U�(�?L�b�|��}�D(���=0�{Co+���S�<qc�]�1�5��#�޽-@UR�XШuh�������n����=�ˎ_|ѯ��K��MY�bz���=���Ն��M[� i�����ҵs�Z(�H~�®i��|b@��W�SP��*'�tL�o��f��Q���������Zώ�=������VR_��}t9�El��D�D��Q˖��2e��*����qw��	������Y!�|�����~�J}��+�b�U~&$D�C��-�/'j���w��Y��7R8^��= ����
�4h��Tr��	��>���tǇ9�/��v�����s�%�4��D��s�%z�b	z��M��G�nZ�v��n�Еե'�B�1��u6<}�)��aN,����V<�	{�\�{�?�"�Hr�������Q�T���sm af֋�; �:�Eg��yQ��P��:�BGU�z�5���2�U�Ƹ(��P���XX�q' z���g���a�&9)���^�ZH|O�
�� �Iz)��M�g���Q���hF.��7M��o� S�.�A_���HH���dk^�ע��"Ch;ք�Zv�n0�ag,Ḽd��V�i~��A���Ib��Q���'I���\ې��?yo:�G��/���d�΋1�5^�:c�o�t"�ΰq�;!��BWQ��P�tu-� ������k�b��a�	���?�C&�a�8�ޘEi;�}ݍHH~�����"�,����5���}����*���0��6�����pZC6H�&h�)h.ڶ.�fsIT��@��!�����?�mB�;�\m�r>�a?cJ�:��������#�a{�tw�M�9���g����p}ܤ(�m�Ƭ.v͑�sD>IA���D�	���e�cJl˅�RL�6$3N��#�n��Dl�����D��%ۑA9[gE��0�b�v�m�@�kݱW̄O��Z���������?X�%�݇7��Gj��֥�'idt���ϟ\���OsgC�P�����|Nm�!m'ZҿD���궜S��١ːmru���O��duq3��ŋ��z�۾�C_Kݯ?`�Y�u')�ԡ}6�A��n��#����Gmm����-O�M��}�d�H#��l	�~������{�I
��3���1>��[��' ��D��!X�2)��m�ѕ�=u1j�������9�1b�bKP�	��`��U4F^]�+�}�RRw�����o� gC����cX>w9��")�&%l�M��;[��p�n�����^��ʧO
'9DB\eM�8�J�S�֊U\O��@����2���_8�Sٺ��9؏��$�WE� �����5xl�u`�D�v Q�&�p�=<�@�fj	�N�gC��!���z��|�Ԣ?�z�$�v>!S���-���^�(3�#�BdU&�H��]5��!`v��76<Ͼ�c'E�k&pc�d/6���1hc��oH)�i�V3H�CTu�q�+��#�ps
B�t�* �_�Z�6�]�!��z���0'#���.~[7b{�ۤt�(3X!K�� d8[����C����h:Hٳuc��ƹ�2N�/z�j�oB�}8鷈z�b:ޤ�)y஝>mn
5��C$���H�H�v!Kb�����6#�'1���-eƉN�W�C;�(��@!M������t�Q�,lт5c�E�ޮ*�ߗ������}Ȃ>�vbK�YA���N�ou�a l���^�ώ:�V�pܧ��W�S=B�ҽ��cb�FFcD"�����nG,��oK�{d�)ڱ����A�WҠ����Ym?��,)�Z7R��3�ʨ����(W���b���-��k��2�y �ה�0�*�c�E��B�JH��01�?JǍK�����d́�փ���2"��qd~y�-���Np�.J��0b3��N]�����z�F��&�Nee��wz���#g{��j��[�:),.b^Y�%˶���Sd
NI��{6��Cg�&$�$j���H^'`=�{q�'��#�������}�1�y��zLk^�}V�����Xh����K��g�Y�A��&�����X .���� 	��y=Fgk�n(���|�(}�'�ˉ�eA\f~2�oИ�@XM��k���%4�]��3-P��=.D>��&
}Ŭ�{p�
���aH��� 0DҘ�����3���=������(|x��E��u^�m��5Z8h=&��1��H�ҵ���j.�]�<-�X�ϦF�;.ԫ�^�wz�{|�\�4'\�Υ�R�K>�Ţ����7W�3g��h�`��3�[MŸ�#��\?��c�'�ߜ������Vs��Px˒	1IK��V� *�?竹BlV$N<�����T2 @�����-0�[z��H�)��Z��#��ڲ�<΢���^?Z�j�1^���#�WG�,�[%E�f�p���<�X=c}r��%�@`������i���"U�D�w ף7�[$�K������}��u����|`ICW�8��g��\T,��b`���Ztl��������8�>�ɯ�ܑ���&$�����q�m��y�|��#�{lЂ�CGȶ����a��`�>Me�y�"a(�5�d[�=x�R
1qED�����(u�n��7�˼=W�/56f���+���9�3��(�wd������՜��򅮟oL�6�a��]��ҫ/-C��
%S�E���'(����C�6]���(P]�6`�:Pi����	�z��2�.#jX�v���V��w~��z�ȣm��;��Z7�����o��U�b�[d��1�iX;������Kazڠ~�+�o���VN��t����AA�r��\�}��bMWɌYU�V��y����?"-7�!i��QE���6Z�0?�*ur�@�lE�I �����*l�:�գ+fh9�-���RE���Aq��[+�S,2�[mf���/�%�$U���w�ZP��qN�H#��X�X��g���-��	�,{N����X������姕M��V(]���A��͸廫|[�4�($�SN�m��G��lP�u��Ք�I3q�*�Z����ýݿbn� �1)��{N
��WM�p����J���2�HNJ
���*H�r;�v��p�W�,;�SQ�ʂ!Y}����
�z#Tx�䵗<&K�p���Z��+y,(V71�Y7P��E����u/x7��VBb%P�݃nI(�ڗ��; w��j�r��H0�x���Pd`x��7|#p�ѕh�]گ����x��`���w�ᬧϒd���L|���D
���;/��
�t)5�#�#�4&���[��o�$h�g����N����A�����w6�I��CD���H� �[^dY�o,g�gDxoȁz�^���.� �,0w|�Tj��ݘr �j�1�3zc���r�F{�ڻ����z	�A���|��:2ңj�I��#��O�7��/yi��>Xz�lk2w��Y�| �K��ؾ�����c���9ue�w�H*�2�I���Fz�@	�h�F�'��DJ�+υ$cs?-I����[͐Ӯ�D:kF��Pc[��!�h�o�Dy,g��*s���}��,W�S-n�n4�Y�%�:�@r3k[�x���l�͞���`�/ޣ!�C�YzNu�����`K�L����C�6z�mTc�y�V��dud��z��o��fC������15W�|'��)>ǭl�qm�A���I���,��:1rp����'������-��|<1A�Czu����}�%lP�o��rX�h7�^O�REm;Ɔ�5�M=�	�S[�-vV�Qכ1_;P6>�5%W��M\Y՞4�dD�M��4�G~���$��jo���;Rś�ڃ]�E����#�a���
���ѠG#0���'�tl	����ӻ���Z{��7�ٷc���̒w���@���d����t�b��-�Q��UH�I�rx��/�=*�~�54{ҿw�1~&����;��r��U�η°5�{�E�³��̪��wW-�`��. � M<LV��*@��;�n[`�䰴Ǿ,0<Ħм�NJ��[v�"�S�<%Ǳ��e,�ض��������l(��H�$��NG*r
`�w���}4*�W.��QȔ"�`��C��tO4�(Q���cT�P��]݇�=�8���x �!>��� L���h��o��I�ì_���7y��0����FF�>ݨ��y���8�
t�WQ���K/2 Ɂ/N���H$j�~��U��N�)�.N���Q��?O}/�J��p�+ғ��'z ��Z���z>�}�[���Ă0��~0ݳ���UW�Q6�x c�>w7u~��J��l����ҥ�(�(QRj���#�<�	�.�㔰_f����j򞒢�_J��9 t������F�z�٬ҡD`t����W�4����"Mm����"D�.�%��ˊ)_�DuEa�J줩X��H�at +��+x!q�hh !��(��0EtS@5�F��miH>Zΐ�Z��uC���ݖ�m�"B�J_�����H���Db�rk��J� ��5m�fb�+��M)X�`���]�v��I|T�`��v#��g��Vu�c��!5B5��Z{8 �T����"G~��VzGuosdֲ�*��g���u��:2�J7����h��Š�//�3V6&��w!����=BrTġ���b�J�K��"��~Cb8��Gd�;U����6���������U�����`|��m�4�adn.��
S��Ǿ�4��@g�JJ.��g�юMK {���*x�V7�*lʶ��)�3<^��yE4�g
K�ƲF6w�%c�Z�G��Ƨ���=`d���fyv|]o��e�ǫNk
�f������['[	tvц�F�T������mi�ܙ�Ϩ�B��0��n�50}-�ԣ���[���1ݫ���(ns��U_�׫Q�s��-CUM�s?�l�R������H��Of�HI�PAI���@�n��Vi+(������$?��=�dA�(X.��js�ڨ�U�[�גc�eV���V��a̕����dI}�O��w�m��{)�Rn�K?��z�(�H	W<3]g���;kZ	�c0XF� ���D��;�p7�ya���&4X4U��]�:q��|s�p:����"�Z�\|������ܺ{I��澋0цQ�� 0�i�B�F������5��	���͚+TmM�����ք��Dco�" X�Q�K�kޚD���7Ȗ�s�v0��N���v���L��e��Be5��7é
X�"��m�C�~w�udD�Η,d���L-<:��OUZ�����u�^���YٶI(6�!���.h���i�E�=�F-�؎&�x=յɥ��T�k½*��%�F]�	�e-��uo�{p���y�� �ǽ)#�c�^��؎��4T2<A  ī�9������~��o��8���7�wtYr��G�R|B���n~t���I���:��(,ug�>�#���Y��YmT^�����d���ȶ�X6�ƥX,����j2��5�Ⰻt��<<�k$>���d!����-Xzh
��l� q0���9zC��8�|"�����Xuo�V�(��ⴶ"���Ƈ⢕�����dB�e��"��3D���N���{��O�7nt��:K����:�9�F��3)��>��"D����
Ǻ�����tl'ec�9.��QБ&�q[��%���.f��о<��mH���p�,R�$�ܛ*�0��e���C1M���b�3��j.���̓@1�:�{���ArK�%�Q(-��V*s�����)�8�dQb#��*�?�B�� Z�?�6���=�XR5>Vf�?��U�\���L~��F��	�#|<���$T`����Ol��\��_���߆G5�j�״�m�a1��������4�����_��3i�޸�N�2�Yi��]C�bΨ��1n��ug���&9~�"tZ�S߳��v"kWO�ڏ��
w+�V��^˸'���p{�;��Eg�o�����-ej�3�����ٝ��uWK�@6����)��GRV�<�x��7�g�kF��ܿN�;W<��1 �IJ��Cۅ��ٺ�,N����Q���**l�x�%�U��&��u�`���<^	�[sVt׈Ñ�����_.X�N!���\��>�ҳ�������6����Z�q�(O��R��v���`g�7�s�3r�����,Ы��s����KY㦯d���Kv��%[bdĳ�BY�ܚ(��j�)Hy8AJ�dR/8�_$��m���U��G)iT��h%�r������?ץ�A�;�y���7	ղi�Ug����������ӭ���$6��^��VE�'�Q2~Z5�_֙��r�;��.g̗'DM�
��E�ȇ��gxf6&�Ěfr���c����ww0��l��N�i[��ʣ��2X�1�$��K}��(
4ÃW��y�]��ln��;/�c9/<��G�~?���*V$5�5��MFg��m��Y=��}5+��/��5|�,��;��8����jj����3i�݄qWA�&'���l�25ql��.k(O>=�ـ@>N1���@P��Կ��#��hl���V4jR�*D��� p#�Վ��;��3�"7�^W�>^�I!��L-g�zc����c ���3-e�e�j�P��hWB�����<��ԶVŊr�8�k���[���{1&������Νٷ�2�nڻ'lD��Aw+���z���������'!}E�[a:Ȕ�\;`/:@�+Њ�t�{�: H�D��u֫�a��On[�C,��O�ѻ	�Mt�>H�/,��6�Y���aC�|��mX�����]�i6���L�ߝ�����	��o�]<�EA��Q+�&��s�1F���Bjc��e5{z���U����ƶ�q�TS�"�x����)�D^�m1�j|�)�2��U��j�i�� @���y
o"W��9���:�aza����o�[���ehP��A�(K��3�.O�	u.7�$L=���9sVh��``���_�f��6�+?��慼W�r��i���n4�D�?�� ľB8#b�=[�:+ R!}s�3�g%��T�p=�}Å�0��5��,�c%|���S�v��́�F"��O�֒p�nK��b p?=W�eP;�5�5t����Y���֘�C�a
��D.��Hy�VA3�[8�؋;$�o��U��V�[R�~{B�M]C�z�P�ͫ2�mL���4�Q��*����R��PB��R��/k�L����S=>2�b6k��)��ض�<W9�ݜ�G�?
�GE\�5@��0:��X�/Nķ��6�kǟ?x�Uɨ�8v�'jA�+�(|qN|���/��b�|q�ؐZ�.����+=��e�ӱ ��i���[����}�荹qd���Uf.�xaݥ�%�K���*�$�وI2Rr@�Q%��a����G���M𕋣Ҁ��e�y�s���	k��swS�+=�F���3�3o_2aB<=#W��P6�U���b�o�����),Vɐ]�5�aT7Qv�r �\�	�n�+}-^,�fnc���b�`�Zռ���eV��1�>�i;��pc��&EJ���4m r�^��}���,�?�=R��E���9���kVQ�lO
��J��V�JY(�����^z,����G�2js�QH��W��`=p0f*W;��o�����1s�QY5�1�_	�h�z֕h�J� M닝��3�|QPc��h\G��'e��'T'	�x�w�Q�h�A�@���_��gp��.]`��O)����+�$ê�z�Y��z0�r�p|���D�x<H�IK�x8��~�}UDK&�8h�|w�IM[O��W����"?|(iW��	U���0� 9����jߤ	��c��Kf�����)�?�X�,�� �ft3u��<>�j�g� �b��8T�z�a�J���G�1ޱ�˜�U�t�Z����ͱ�0�I�Ż��c�wg+,����fM���F|B?�Oa]Y��kpʵ��]`�9q*3�Tmΐ���/�xGr�4�.���Nѳ!d�<�o���m�����6��MSfU����ʏB�u�J�~�#�x�bC��c�"?�T q|A��->���b��~������Lm�A��>��@��W�C8L���&�uI�,��X��A���F��P��hX���\.�Ǣ�`U��x���w�OAn�(
�>�(�fP���VW?&�N`:�unG�D#4��F��CT�g��D���Crɮ#���z)b��xt��G�4����0��wQ�wyĞ��R�d��S��`Yp�ߛ�Ǖ�T[�ر_a��g��ΞV3T,���eA�l �h?y�&5��R|�DW�����Γ���q�I,jX
�*�Uvl ��k�w��(7�3 >� ����M�0��aϐ�q�vW�i.�r�mu�0��j6q��]��X���jfA��N��M��Q��8gDH���w���Mn ��<����?(#�cr�)�����"�C��	^0]���M����'�Ӕ�Zj!R�"c㨀�q�Ya8v�[ߔB�r~��t�-�Ҳn��Y�<p��Xm�r�p��W��Qw��kȝ�*�8�nz�A�eT�1�	�]_�Z���p�|eK*���J�����a璺�]��M�qìQI�����~c#��P���^d��:P���׸u�Q5��3�B�2b���}��d�����Q��4�4P�W�;�X;6��x�,_h�('��r�c&^�m��J
�$W��͚��V�<���%�����h��s5�\'��*�\|^�f��.��3�>��8�-�d�n�����Nd���}�/�(��~�`��s.[s�����z����5�M^�ٛz�=k�>���G�
r��jG�U�59�@�ٸ�xPF��tȖ=K�v)�󮦵Z�К�-|�Ǽԩ�΁ȅ��y?!�`���[����_��s�,���z����ܹ$Q6s���� ��؊Ne�̣�/�P,P���-����5����s*ei֏D�%���ΑnQ&�M0u�/�H������נGL����[G���a*��J׃ur-ۃf5���G��r��)�a����Fn�Ҿ!���
o&���U���EC�x��3������� W*�"��/l�$�cR�Q2+D^%My����?�v<�s3&H���*N������jqB����� |=��:�QYtU2#_�{{f=F� F���l�n16��ňh"$�vHѨ2����Ċ��X�U6��縖 b���ߢbg9�ib T'|��Ӧj�e�ᱼT-��q�ap�����B��DN�72�KB��FYI��L��� F|��>�wEp@�(e!s���o7 ��9���%ɚ�+A|�RRĚ�w��v������P�S�*�M��g@Lm���BDQrW(˵q��Uv��T��|pg�WnʧFԥ?rM�L>�S�dݙbG�B������TRZ��ڿ��,�^%I��&b����^��%��O�~����V�߅^"?���C�Bur/B�H5�"���8gC$&�r��J��Q�X�۱��݋E��������>�!�#�D��4}0����χ�_f��_:z<�8�l�ƶ�Z�.�����O�kr�ޟ���'������~����)��u_5}O�rF?�g���;��7�g�bt˃Q�{Qƽ��n�p<.��P���^���m>;��#Z�M @w(w�B;Ny��B,��4i!;�r�\޽��F�i0�|�<��(N��#����-�V"7a���@��\�v�A�*9����}} Z2e0p�Jܰ88vs��y�v>�t�٢O�H:k��Ɇn�īʔ%�(v@�zZ`��(�@N..M�n/tB|%�����])��A����׃�x%�xyp?1(�Ө��zT�����dlss�zw�E��ncq�������l�<F=a�-ܯͧN��P�1au:�H�8(pCo�e��(����,����W}+)@�.g�s7���|�ZD�$����W��b)�$�B/9 k(u�Z��V�_SX��Ŗ��)('��Qٲ3��!DJ�G�0��5��#7ΧM ���W�Ao ��MS�2�M��V�`7V��ʚ���#���N\=���g/jVK����}�K�ˮ���ws"P��G���xT-/�K��8�N�H.�*�B�y��b
gA���K7���ɭ�7��F���$��k��g�S8,:���y�H��m4$���m+���]�m��.<u�	
�Dbs����w�=<:�����(*�����/�6j��XӅ|�ĔO�'[4��(�6s�>��,�]����8����Eg�;��>�[}�t�}i��2�������̲o+���}�/S{J��Q2�R��I7S1���7����,�;��8���TU�I�r ������O0�$L�W��7l0��K�H"QU�]{)t���2���0�E�m�S�:�L���V0T>�myx���2�6Ug2~jϝ���n��h�21��
���;���\	௠(Y>�\$Cp� ,O˴���e������K���i$��T�Ϣ�,L6���iȮ{�\��6.{�ܴ���E<%�<?�*&/�����|O67f*;ܶ	�
�1B͖yЧ�Q=��3*��������e=�����B��mͧ	����.��Uz�X�+[AYv-���n�	�* \0JMۍ��nU�I������GM�*�����^�c(Ҽ�()f�m90ޚ?��ն�.�9:(T�����s����Tނ��p=j�����>����ԡ�]6�7P_i�RS�Zld��´��V�/�/�L��Rt��h�W�F����M���A�Dr����X���e��)!��fg�|�*�E�(��et����p�J���_�r�s��y쀴8�@�L�(��o�ʝ	{AÅd�&]1�4rK^�:/�t4q�}iCy+_6}+�Rj��*�>V�
� �����X�3K2
G���_R�KC�xn���3ϼ�E�h<�>�'��h�k��]�m�'�j�Z�+D�"4w�D��d׳jH@���"�6Fq�yW�uv��������H��"0=��Z�_�OT�8�� |_�4�C1�y�P�����\�1$,�9c���(��7 ²bɪ��ӹ�$��GR1�vd�Y�)�.�+�y�SKQO��~���ew3m4op�[��8�Rg�d+5��s��jN q�S~��\��
5rݟ�B���z�ޠ8�le��Ҝ�SY���3� wp��"iX޵�\�Bsm�D��k����gj �)��vqU��eiO�I]�.$���(��{^�M2-�$��M`��	��m�����mɃ|T�n%��2^��Eә5;��i�af�x���J��;D������S���~�T��"U�-*����jb��~KNu���9�%,,��k�y��(�s� th�60mjl�n�Z���A�=�B%�{�ⵒ�#���x�L���6�[���q�
�M/`�����.�Vۙgi�-�9���x�4�<������;M����_Pl�E�(!։��T�ʢ�cA�	�������O˧"�5���8P�/�6Zϒ]\u��iV�cEϏ����.Ct�f�<I6���f�{�����6�A8�iNE{�C��B���"��֥Y�@�f���ે�+9r��lb5V�����Ig
M�������"����t�f,b��U�-��im�������S�и�]���5�F!'G>Z�$�/�&�(�`�8C��M�cƉ�~��~��+=�z����d3�UXab)s�{��I�
v�%}�0`�c�o˻	�B�� 	����t�[��h�A��p�����"����~F��ݥI��?!ղ�����5�&$vb��b���t�l��`f�=�1��6{�]����JGh�j�iL�G��!� ���0C���t�yi��cNc	�p�he�ſ����K�#�����~%�
���0�f]O���p�¢�.LN�ơ\�����X����ii��Zl���P����]N-��P!^���W0m��C�|F�C����d2wp��X����zt�%�I��PEV���=�OoW��P^G�h�c�����I(�VI ���B�J٘����c��X*[v�i;�?�<0()���ռ�_���F�4>�S��)]�ŚQ���7�� �b�?�Ԝ�����iߜ*gӁ"���IF>bb^[R�M��WK��S+\�dhBɯ�x��I�Q��i�X����3�4�f�R���b/x���gLK��*z`���'B_m>�
Q������A��%� Ef����.!��cZ{��/����ͬ�i#���V&L�`��Wz5Yv�G-�$	�U���8e8��6-��o��0�U��7���U��3`�@��㶯�c�fS�9�'���}��_It�HhWx,vU���/c�C�g�-/>���w��-�t�~C�ƒ��EG�y)�u��59n�ǥ�<��k�3�^ͻ8��4�A]'TG���Es����m��*e�nAK��;߼�1�5��.�����]�ܚ�GnZ11�^!N��x��������}Q�%B�E'��{��Z�5@�d�^�F_�2&8�x�gٰ�ރ[Џv�e�z?��E�Ad�9�����@� ��?=�s�鎨�O'`�ߧ��?KC*|�b��/$g���0�m�/u�BמC>%�#&0�G9ӻ/)i<"�e{}�1=�N-:�� %]me�q��y���"�AdlH�uMO� "q��m�����v�R~c����q��߽� 6{%�I<`v��� �SP���`2�%T#��a3"���s�q�	f��sU�Y�m��/� F\,9��P����djR� |��x_����xN+v�g�p��ߨw�"��G�(�
�ōՀ��Ţ�'��Dui����uZ��d�.s��&�*�X�Tg�ׄ��dS���K~������L7��4m�5̢�ip�2�ۥ$�+p���;$�FE]�t����V��y�\jr��%�!�������
[�B
���[%1� (�Qc�v9��P�d��uM�`��z����;�$��q �`�=�;��6E��q*��o��FZ~7xa�9�A� �����Ӎ+�{��ib�w��&��hu��j�+��aC�z��b�[�X�N�QP��$�c�"�j�h�t������q�:\^y]�Ѳ���S�bG@]Wƣ3'����	r�%#W@�b��A�`�&EGҽ�)��#�ŀ���sg��D��:����	����j^]�z��j^��+��7�����'�C��߷Q�d�
�-ˀ/	�oԤ�<��9�8��Z\��aǙg���<4=����3�#���y�rB�����7:W����܀y:3Q�u�Kh�,_]v���Z#�H�"��9~�2e7���CX�O���C wa��4t�C�賝�$�_��ᕬf+�-Qg�S��4��Sp�QJ���8h��O�����~7�J��-��������?*�'
�o���_�ڥ�%�9��4����[�$$ր=�M^���,��'����f�mI���a�30M���O��H�$�H�[�8�ߋQ<�*�^:*>�������� d/���I'S�Iw_k��ut��Kx���>�ӕ\�t��5�,s�%�WfZu�o�[�v��9��2n3��yKa��V����|U��n%��B�3���X,��Q��3��*�15�M��D�埰�����G�==[�q�?M/�D�̂�gS$�.Դ���� �%pS �w�n qw7_����L��ͅ�H�ւ�N��W�qn_��1] �wJ���o���`�5c�P�5�P�@^���P�e�v��7�����L5s��[�g�Pu�{�P@��1"'�+�I:�w�;�v�����#�1s�>���#�v�o���;�vP���S��+��z�����Q/�zW� �����vt��mxL}��W-z�V\�P����Ȧ��`GU-O��I����������Y��n��z��R�0+�Cm��E@�@!پ?W_�1]�����8x2k���������V��r�����v,^Z����7�פ̈́�LTS�<p��r�2f����	���K?(� \��Y�wR�9d�۟�ۆ��>�m3���(��2s��<�rx��IHR��"qX�(�`N�c�.�dL�9�eb�_ �+]$��w�R�����V����E�}Z������~vڔ0�·q�5���.qZ.v!,�D�9'-���_����F �,� �}g��u���˜����X˺ �1��^z3��W��^!:���5DfU��ľ�K ����B�ie4u'C�&2����B��gt%���+i�ũ��X�3�[�q���\ �	E۞�MOC�!0[?�`�׫���_��ty/��޴�^A���/��I5��.&�x䴁rvS�_qV=$�c��f4���e6�w�v�IO�< �I��6�p��&�Nn�e���>�0s��@����o�5�u�V����k��n�V^��m+��CP��[�v��"v'���������+��X�G�).6XZ"PU�(�g��/h�=��3	��a7�[-�T��y�Q������߁�b���T�v� 2$����;�aSa���dg��eϛ�d�O�%Tu��K�h��o��#E�U����?����P-j%�(��J%=O}DV��3�_ƀ4����DS��~�M��Q��E�Bq~���c�c�&s��tPWXn2�X�%��^.0%1N���.�7W�0��Z�t�|���HSy�%L������ݥO��MĖRj�ǁ�rM��c�kNjF�Ф��Y}�xˠ�>s ���t�]���xov>�����RM<�Za���˃���nj���������?�}��.%.�I�3��7�n������b�_�C7�>(��<�r�UP"H7�t�I�[�U���7��+�|p^W)�`~[�x�+o��!��f��q�l�AZ�̈́N�u�0��Z����S���R�vG ��4���*ƴ��/[_��.cjǄ�O_�eM.2�*�-Cx��e	��ڜ	����?�E��utEc:=��hѴ���� L���r�� �p�ȏC3�6?n�h6����! T�x�_tof��R����*sO
�_T�%�y�D+����Z��|�e}�p�tm�� }�g��t�2�6(L8|�Tm�We|�8۰�<2��&���t�@��5�S��N��o������
���30a��a;�/1t�kx�Y���5���5�֔?B����q+��D�e{�����������++�͕g���a�G��3�ҧ[���_��C����S�ԉ�_Ded�۸�I���8��ћ}9m{F��f�;�A�i��:��h�nT:�0��`~�(Y�������h�=Hv,�)�	y����G�8���'����[���~�蝴aV����Ud�)�����%7�l��R�h��6�3ʢ��L�B��!;��1% �Z��ġ_�m�@R-�����X��-�bLR�����6?��TJ(�!t��܀L����z|��~vG�V<��Ae�N�($���G�c4���)n����#�	��unԳ�����9��{�������t�
�U�+����0�����MӲz�8):^�9̒>�J�SI���-��l)�l��ò2�VEw��p����E�C
$�YUm�a�g�EnJ}�u�ԅ_�x�Z��s�������~�*��¬3L�ZT�r�r@���2�}|O4����$	�����r̺]D�fj���4���t�b#�<�n��2���G�p�ʵ�eѦ�2�������4��a.Zg��(���ͻ�7|��쮍sz��Φ�#������D����ef��DqZ�9Eu�>|{�;��&ߡY�>���
��ͭ	'x��<$����u��LƄ��X�@ld�OJKV�PG?���BR�[sN�����^��%9�n͈;EX��Z�#�2�b����v��}M����Ä�@��c�j�Ƞ@����9��GbSWx��+
/'��3α;���}���I`��ϭ�wV��ɞ��vS����ǅ��e�zY�̼���V�]BvO�O�B1���q�Sk�?NtS��a}:zG��>7(�f�᝸K|q�Hɛ��6��4�c�P�I� �o�,�<T�Y�&�!��y�p��X1-�7���7~�i��N��(%U�&��t�ec⁹����<�|���)0~��R6b�?_8e�m^{�&&t���l ͡;���ЇMI�W8�8�)�0�r�9� 9��|��:��� �0���������I��k�a�*.�²{ҵ�6�qef��r�����=�yMY��J���M��$z��h�9_}�)��kq1�Nѡ����-Ĝѹ&�=fh��ͣi�i|�a�d��ޓ�Je�]hA�z�A��Pơ} �Vׁ�3Iqy	��	T�>gu��*)���,5�|N�斄EJݲ��+4�|�q�0��)*$��иxYcw����!�s�yg��U�SP\"��8sD�o�������ߣ&�Ŗ��0�6Z�u�=�Ѡ�����=�K��$��f��R��U�
7;�J���������)#Ǜb��S�ݦύ�L�0��XW��8��+��`f���C�MZB��A�2���+���ha�ݹ4_,��i֏�I��f��NH�����Ư��=����2$��𚤽��`[:�y�8�)[�s�1WT��$N�w�M$X,]�Nhk"t��;���E,e�D�AtI��O����y�Ţ.��_���C#���#�ܖ���#��~�q>� �ސ)@{Û�yN'�O?�!k�E}7�j�q��ETg�H��5��Y�;CԀ�1IZS���1���$R/O;1*��rA��P(ߍʆP��s %7=��:�|�qEB,m�ܓ�Ҿ�V��=q���b��uf��I�vJ7�R�V��}EӚI����K�|�|IM1��O�ԥ��3���I&����+급�76��\H��0����(����D��� �g;Y���4$����C<Tn%�*)jEi�'����� �$��۩��ky��O6�ǎ����� �ˬ�(ޅ=��c���/ހ��X���yeX�EG��۟O�gv��ե�g�{ɍ������f�pmv�N���Q���m��d�s��[�͠��m�7A����n�V�����zF�h����Jd;�U	*�n6�zx ��q��b'2���LD��t�������gXD[ ���*���aUo
I�X�+ҧ�;�b@r#p�����om�����ӗ�XO{AE2Ϸ]*j΄�+.x���?1���,��?��P�:����(���1󢐷�m߷rTM
ކ$��"u��6=Q]}?>����D��n"/h�:J��&��54�y��g��M���h�OK)rC|i����:�9]
���|⿺~���NU�&ٖt4GFFC�/g̰�WRs\��GX�vZ���-v/��C�jH�t	�����b�P���i������gˢ7>�E���h�=���s�:�_\��/��1�¬f�L~���yJ�ouX5���4Y�enM'mM�� U�;���Q��va����N5*N�����MX��t�0#�J<f�n��$���cl	�[-�Mƫ�bq�
�r�:C�vV	���$?C�����d�Q)[�m��6B]��P�G� ��f9K�r�_�M�fY�� =�CG�s�h� ��t]?+�����;�\0o[�'t�����>a^@�Tأ�P��"$/�S�������u�cʈHP ��0�U6��I;�a{.�?j7ݗ��Y���[M���.ll�E��5"��VB�x��X������^���	�d��(���,������t�0�%�m���g�C�� �W��RZ����E�0�}mb��A�H�+h�O���������O/7�h;��AtM��)���k��
��*af��48�9@�\k�M�r�Sy_).^q�-��5�\qe₪���hQ15���� V0%�9 jk�g�0����u7A�c>Χ�<�v���K����ޮ9�gOkPi�~$Nf��u��_�/�|�x䯤�.a8t+����
�͇R�˒�（�E�G O�c;��I�b/�4����hu�&�#�@05�S9.1��X��1��k*]�M/ݤ��r����?��xy9,�[�j���N��d�32�2{��y׹���"y|2ͨ�_�5��<���8��$�1��1�9T=�)t[SX�Q师u��A��n��.� I/�8���~�_�g��
4�-�#2x��@������!w4Ь���d��i���5�����&R}XD�t�t��p��X@1_���li
2��)^w
��W�������]Y1�.�p7�M�A��k�:�bد�� ᳴�^-E��=�ᗿ��.~Y`P{��2�D��A��B/���HJ�?���{�5qhx���>FS�~�܊���>TSV�AQ�kY�CD�˗�5���0�hg1�H@�f�̯�a���1"�~�.?nc3���=�+�#EIjjat7O��Xt ��������W��")h���&N���٦��	��~=]u���`TH�FPZ3|c�;��/�K�!�� Řg��K,���u������_�5�ϫ�L�}��E1+r	}J?&��q�u�Xc��k���P���<f�(�l�!�x��6&�(�yQ�*{�c�3��OxI�����Om<D�u;��`��$���H��vY���-�l�1RZ�rsI{3�d�8d�"��'����+ �m���@͑��h�^��y���:�+�O\��ql�X��K��, .\�Q���y��`�+����:a��iLֈS�BέEb
n{�o{�^��v�,�1�W�2�s�n��L}n�ۥ�"���u*D?Yd�s�H�۹��)����R�>v��F��z��Ej8KЕL�����8*q&��@x�5Y��)HJ?��l�9�;��-��'�a��"u0S�y8�ir"R�	�s�i��bGS�QZRo'�R$� r�[}(��J�=`3ɷ���u|����r~P*���R2�D= ���d)��~�^c�	+��/��E���Β�M[�Z9y��J����+w�S��k��\��_�cM�-�7aW�z0q�L�F?� ��O��u�t��L��B��a��2��=Xl��<V�N��Ij�� q>bd��x�B��2����ʥ��<(a��F�_�߽��Z܄�� �)k3mf�K��_���Ns�-6�!��=��wx�=��*����������#���+j�)��Mv�w=y>�4vsQ��z|�Z"me��cI��#�Kg7�M7�ܧл8��K���������/O�z�\c����ޖF_�hP�d��L1���Y�+xm�{��FEC5X�t&l��;���-�:�Z)-��$v�c4�k�|�MPr�L���Ϋ�'=���P[���ј�c� �k�������J�t!ت��5;L��k��'��G�7�Y�ҋJ�2���Z<����%���+6XW�Xe��Lui�p*`�w���a�l���Sk�Y`Zl�Xz5E"��9�92DX�9������ �
��Э�=��< aY��Zl*F�k�8�:]�ß�e/j�{����7F���������2:9���>O�C4`k����̣�Ѿ��O7�r|��XS�Y��i�B�t�⒉-��@%��ȶ�԰iK��n�Ҹ���*�����䢕�14�6B(��0�o:s�^^�1�2#�q[�����/T��X��`֢4�Ȼy��K�5�����ZqQV�ִ����.,Z���݌�� �E4���]�S�
���M+WQ69dP�ŵ�T��{��#����#;镊�i�fw��f�7�$�,���ZW�޾`��N�R�Ί���R�yA��B+����Bܨ�c�@����,c��e���8c�e�Α�ܛ������}�~%��9�N4���5X-�:Ff����x�&KPn�	)����Ɏ���cs�M�� ���Nx.�,r>n����Id��x�.��~9��<U��ǊY=�����ň��o��@g8�ٕ�#�Oa��1--+&��*�� �<D�s��J��aǀ�f�D_ݾݘ�.�A�{e~BB�fԅ�bI�*f�4:n�M�Z���c҅e�� ���'��R�Ʈ�6Ǹ8)&`�ES��`?7I�姡:�.���m�0f�Ob�oK���W/������-E�g�>F���	^��g,�5���k���`��3J��YE�U���(�,ӱ/]RM,*,+��0LPՂ�:����!~G�%ʘL�2��"���thaƪ�|�%~L5
P�E ���Za�w^^���|+��X�a�1���C_c�2Z�K4Q	oa�Z�?�Gd���`E	��8
*����c�ݝ��^���,t���tp�CF��AMQVUR�p�MiKF��U8�'�J�XD�NU`�=�2��PW�%v>;Ȫ�#!�y����vHPG�_�dq7#D�Th�'b�ar��`���m}�T��'�����^�:����򺯢����L�h�����pl�F�;���^$��� �[�7�s�y�酊hA�m������=�9��(�8�9,|������G������UO\s
����c�7L�nU&oR����t���r��+���8��|HX�f��p�@���;v�^��ʬ`^�57sF}(�
'��ߒx��+EA�5�H��<�G�$Ɲ�������ڇ5�5�X�^�Qu=f.�S�������4���T.�~}'�<tU �o��>��f��vO�/nʇo��c�|ɨW�	��\�����8\��ԕ�16�X]��w��?CХ��q�F%����(_ҫ�*����3� �� B��p���A��t��Z����ş���������;�F	��aUl����>D�'��X�I�3 =��}����k�H��܄�0���
�>�s��j����� �mxN����ogi�<dg�4N�iޔ~�&�����H���?�1�z��Ҙ��%��' �'��S�1pW�n�|���������H�xu1���|/�O�Q���z��{���Y��|qc]��δ=(�B�|%��N�(�c\� �v�b�A���(�>�D�������[�y�b�o��j��2_o#Ù��v��Xv6��8U�\dI삃,�@_��83Z� ��f�����^�Y6<Œ�cW<��v��du=pXؑ������QuV?**�dܔ� ާdB���:�7xCYTn� ����D�. }�5�n}8�n)K��e1d���I4��)2����4N��`�^_�E�qP��	4|�����~9�Wn�S&�o^��Ex���L�D$��j|k�v�眬(�������y���Q)�Ʈ�Ƶ�Q�7��˿��-}F	�X��P~է 9�@�)!
�=��&'Gc�9FΒv�:E7���C�_���+^	�WF'A�=���=9���s��!��&o�����=<��]n�Vy�*,!�oGO��Q�����	������!L@B�C���+ڧ�jj�$K]^�N�_UtK���⤫9���S$T�>�L*���$eY�[���� a��i�`�̓����>��cKD޻����/��m0��R��'��|>/0k&�2��[�������u�m0.���Qk!5a0n��% ܯ䚻�n�唒�t�G1?Т�9���Q�l��)M��yYK͵	���Ł t-��4|��c�9�W�f���*W+P
�!s1%�S����#�[��=�Cgu"�*��(&@��(�@[uqk�PN ��9;�E6�m��+�n����I��%�?�Xf��%�,R �}D���u��63��s����_��jA�l6,�nL��f'8wt�gW�O)��s�N�v��U6�:cA�2���� c��'u.�&�#�b�g�R}��:�9�p��3�G1��5(�J�4���YkCaO�k��%{,�_����Ƒ@��4���gӔ,U0��*`���I=L(c�(DI=D�nqb�@�x�&�WT���VVUZs<���W�4<�B�A*gT
�_Ab��c�:�%�޾��'BѪ�e5"�@���SL-��oB�T9��(!
���)�r �� ��@�}���.�1U7���"!���#�V�l�6P���%q�mH�S�v��>j5����#�m��Ow����&�~��ل%���=?5�7SV*w���
T�`m%m��[� ��V�%čh�p��e��Qy��\���L�D
���NZ-��<�"�ם=��k?%悑-u	؅@e�j�>YP:�R.x�f�)���,�<^�þ }
D��0�᯦e6b��s`n����+��\
��'���{_x���1'���"R/��
Pw���bm�K�a�a��8'�P8�@�q�nw���$�E(t2f֐uTO�c�;�9��ٛ"��J���XO�a�](�f `M\j�`��1Y�������i�4��/EL��Xvr�_h��@�����s��M���Aj:᝽���n��i�n��߰K*��(=��F�����j�@�"�PL�A����y2足�\GL����;?U#��0���ne^��R���f�y�r�`T=f���ȷG�X�v*� sM��U�YRm03�@�H k��vc��Y��uIo�4&8ބ'�86D�\���LdT���|ܫS*��ݝ/J���|��� 6���ސ&oiP�|ݱQnUy�>�q�?B�˳!��OL?�li6j�	F\�����`?d *�yܡ�#�W"�_F�p�#f%;¬��r߇-�\��T2��݌}W	AH��'+��%ބ�٠s��V����0W�,/�y��6�W5Ov�ag������ZD��o�[�m�K���4Ҧ��~/�E;7g�a�
������Z�_�z��YDR[�y�(�NWF�$��D�/�7�Ք�(]gC���.�'~Z�����ڟ����D��*�rz� ���媟*U�7�����Aw�F�rM��i�Q#&�I��.i8�G=��|>G���ÅwXi$r[dG2S?R�Q�ZR��M"y�O ��Y:1���s�c�C/�a�C�>g�En�ϻ�oȓ���i��d�Č�%^�~�nz|]��z�H!�U�V9{0��+�'_���ZUɥ=`����%�� I@���pi����MD�.�eE~����Ĕ��ѵp&��Y�=p5b����)�%B�/�ƁENwϜț���Ϻ�"�L�5ad�s�w9�}�/Ň~B�o�3��mH�Y�=��n�X�B��.�}"�I(OX����?�GЕ��M`B֟^�|(����\�\ M;����`驴�왮�a�젼���0��h�9������X�n�Md�ݧP���W�l�PM�'��,$@��ڸ�jbmG�\7��9oj�?;1�'Wɔ
�L�q�;��d���u[줺|���X�շ�棤�,?G��Qٛ�j�G�t=�
 ����ߍ��ʠ��{��޾�H�m.DP�C�?xxi��Y:�;��>� �_��C�T��~�4���67o�BD5�"Kq�D�L�,��"�fq2�G��~!�k�0H#h[{�U[�z�VZ�]l�6��ᜒB�1QQ�~<5!&T��{��M�ݷ8��i(r�^�m!y�\|�Y�}x���F�הl4��/����u��(Z�����c�
�E�u����z�u�U'�-�ũy�����Є���@�W��9A�o��pp-���8���{&H\yM؇ӽ��]�����}�.�����U�KE=����V��D���ꯎu�q�U�0�dV�j���m�� �,���mB�/�� 5.��,����iË*�~K��[�'��2�cB�q����;AY�Vf~O7��A
AR}�]o�%�8V�q�.S3����+�!� �� �[4[�����h��N��^��j�t��-���nٿ&�Az���A�*Ɍ�{d�'���Y�p	��	<��Ġ�	�[:��Qҽs�h����Ġ��M�����wς�XܕĪ�[��!�ܝ?�WU�����H��@�y�m6&�p�+YUi���6������9�4��sD"�o�>O��˰ri6�.a ����#��V�ֆX��9I6�iB���t��!Z2<�|�m�W�&ف=���	6��RǉU�+ߡf���ocԨ����,>��A��Ҳ_1�X����� ;(`o+��M��L��W��o��3���sLn3b���b����C�W�&���=U�+��=[�%���E����)� KǂT�=#Ѯ��t�Z��O�h�$�����e�	�hS�fY /�0�\}0u��*1y�
�C�afTn����`� �x�a�-F��L���K6Sx:+��u��t�Zt�_B�S�i�"����;�DׂSɦ�ϑ������\�>��i*�7@U���_`��ق�~�YJ�*e�(unב�mo#�������ݝ�Pn���@��z?�$��v���H]�g<���%�c]�4qj���?����,}X�k���p~8����Q���e���q���;%8�rY�7�;en��}ao��'�鷯On�7����i��A
�����(cB/O߲���n�ZU1g��ѻ�`|��ƙmF��G�ٷJ�m���*R���:��|6ei0��{���>����k84���̀dlєB�A�?.�c��y��kT�
+��ґ9w'e/�<�~�{���Iև��nˌ�������I��O�*��<��|�( M�AS���2(}��o�n����o�&#�Y�[I���Mg��kE�͇"���kO躋j%
 d�
�HB��$^൱Xc�R�i��$*��X���m,���ޟE�^��v��Ə��I�X����H���t�r'#݌i>F8��X�����*K͋�ـc�{���#y�Q@(GƸpZl׼��y�[��#N�h^=M���_�G�M�Aɵ���Z4v�H/�"e��c��;��dH?*O�0��oZ&��Gp:�S12ONz�:vL_���O�q������3�at*�O���6�w!��n�9ù�(h,؃А#�������иz*�#���q)�lsR��-�(y������D��g�/ڎIFW�G����	�	�l&�QP	MT�h��j^���zou_���1
:f�H!�+��V�{�%J�A!�e@��ƫ�yWޡZ��5����n7�ψx:0.r"x��ݣ8�	;���03��Tc�9���]"4��)�I@�K�%��&�bq E�E�|�vՃ�?4
n�R'~T6l^k�u ǭ)��roc�ť[������E�K��;�W�'W�-~Qo]�ft=�w�Z�$���M]�� �q��LO���0q5�`�T�w��cnG-�ڧ.�Y�G�V�a�Π��<�W�>�����<� ,W��
�M=��UcZ-X�}�_�{W���#C�|}��\im�S됼�����*b�]ٱ;b�ƺ OW{��^����:�K��4���IѦ�${]��2������M�6��s�:��;�c2?x�����Q�,��J��%)�;RI�W�	�"���U;X�53sՀ���^������QE������6�Cl�4�X�[���\�{��Lvy�R_�֊U�+�
�]4PT0%�]����_\cWiG�x��P���"ge�+d�j�5��}|R�.ioo�ͧu+�F� /E	�5����1��$�pq-�Z=��V�}�/��cB�=����R\W�4
��������*���(4��%�p)�c�/�-���S��5p���7�[`d��Փ�?��g0��Og�d,�9o�&��&�MhN`��)������o&��ڈq�'~[���^���U`��놀`��t����N�¾J���p��l�X�<����7�M��zb���}2yhoW��g���c�l�0I`��=�6�5���-zz8-�D$Ƃ'�>��ڒW�����U�X�%��۽�%�7�r)r���˓0�|�|��]5��7uI8?��C�R
��!3�����[�1�":%�L4t�ˇ�:D0�Z��-l+���z���sKBV�ͩn��D��Ŷ�l��oS�U�\���7��	���{�g��B�>������K)�g��9��&��J�KI)�/��6��v�m�n�����4����e�����jU�a� �a�]��>�oz�~�^NΔ�Y�
�K�Ұr��۩�B�����uPsCB�3��/���Cr'gV��Q���#iA���"��```��\�Jt�wa���x�A�y���<QT�r�I5fnL*����H���t_[�nH%�'�a�N[?,#ؘ'�J7�G�(t,��UŌ�1;�T���T�M�O
��lϹ/�>�bM��u��5�(CʆLTab��=���F`��S�4���Xs������[���yn�u}tٚ�b7�E��m9���@G"(���q�9��Q�=����T��a#.دϰ����S�H��LQ�0��L�(���{��\����U�NZ=��X����S|R�'����+�_�w$��f������Ⱦ~[ۻ�$O����:X������WUz���1��� I��g2���xй�̘>�k�"�?]�.|EKtn����iQ�*��K�b�v�sʾl�dd��ℇ�f*�:>}J'p���*,�3qǷV-�z7)�m����+j����D�|w�H��x���nT'ĒqQ|c%Ƥ��:������$͒�=<:�	���4�BpIi= �������� ��i�gޘ�*������J.�~?u6I�S,�R�yh��\����=]?�z�!��r*,���I1N���:x�X��2��7W��U�h�1D[���<x�жBȃ9AaY�����V����{�`A�#��5��w��a��|&ȯ�q�^U�o_�-u0̡��?t�eHbڠ� =�꥟3�Mֳ>��D�NQ�\�A�`Y�:}�F��p�3��;l����D?+��m}_&{�S�ǚX;�CKAΔ}"3W8��Jg�.ۣ8��w�\cS_IV�cK!uJJ���1�vצ��j+�!����$aH�?β+�_YnVI:���k��Uc0/`�������؜�U]������yc�.��־)������,��Q�h(�E��n����qS��Fz�g�Ŧy8�Y�KDԽ��䨨`R��M�wT��Pg��<^C}T�s!|�Mք�F���e7̸8@�&ح��Ĝ1�b8�pv��X(��%r~�c��Z�2w!����D[�>f�<Д��� ��jP�/ �d�t�Z��|^��#r���j�8An�r��|WW���z�=xނ�[�B5�W���3�����C��O� &c^������3Q�n��b��~V��&�8W�	��	����/�-����."���0���M���.9K�A0�չ��d�攨��ę�i�u�}�cW�}�`���xiM�y֜���
g^�J�s �����_1�#���<io��F��Џ)����R��=	E�ɫ��_�j����!r2Vv_^��&��q��.���̻�S����A'?<�Ċ�� ��d�I�V�u���<�s��M�$̫����$�J<�Yx-v.�}5�8��T9�>n��
�:R��
s�I�b�8?��@��9��ޤ��Z�/�V�je��L�_�~/φ������0&��hG�ie���,H9Je�ݿx'��Y�,�@nj��B�¥OC�'�C9 �X{��F����ʲ}YVe�g���<�Qe�p��E��i�)���N�F�<>�=��С�O�K�̥��?Z�f�(���{�Ž0с���ӹKG�����"y; �7���7������x��?�6Z��`���g�lHdC :�zә��.ޞ����FJe��7�����!����_�qݟ�7܇P�2�xc���a�����oP�1DŚvd��Q�%����dYdvg�kFU�����>ɇ.�#�i����jtoxkvŜ+�k�΍rۢ���J6�O��h|�J�/P���87ɜ�&`A��zX�W?jF�I�����`�>o�RV�a�`1h���4-���p�V�p�ςJ��oF���PGt=����E�,��Z�)�ZW�]}��u�oL�$7��.;�J��Á���!���n�`�`t2%p!)�P�QFY��1�nf�p؇Km�M'�5�Go���3����n2�6v�q��q��p-�F-���S/���9�,�$�0)_��
��p~�@����)��u~��~��8��/4������L 5/E��4�i�]Uب��5�=Skr�`
�R��D��4���+(<�=_k�D;���R��׃~R��#W�tl�K�=U�h�$��皹^ot�$���-�
8��;!�_��Q�{����bfXGKߵ�aEНO�;c �|�EbF��fh� ��[�?aB��h�5�����S!]�z�%�w9����)|�m��E��J�ʁ3IT�N\����Fk�z硴�Z��C��z
M��M�Ye��*_�6���?�cς��0�����[띇��w`�"���2����~�������e]�d���R���t��!���f�p��J���^�k��u0"A�t��A���ixwe.��@)�Q���(>W:|��|�(Z�|~��)�p%'���4�$B!d��x���j��||-�?n�
Di���=�B�x
��
�D��>s���X᷽�ME쀋����{1GD/	����k��v�l���ܦ�@8FJ�f��1f�5�j����]}*	�F�]O�@�[����	��||h�|�_��dP0�虏�"K[$��d�whr��!?���̋�C���Ү���p��ho~;=�wį`����_��D��Gu>���~����f��AlT,7N�3��.��M���'��_iD�����ض�"�6�����ٹ
N~���s3y���i.��#]gGLJ���ڜ�g��eF��I�4iM��=j�Ch�h)2Fl�8Uz�4�B�;/���m�"]}xub��_?��NL��������h��iQ�R��o>����4OҲZp�z�㢤H�ʖ
}}pv���!��s(3,E ��.K����륁+��3��i��;\�����.�&P���=$�����U���Fݯ��3�:�ܯ�l<3sx0>>>!���(�~�D[�c�c��$���e��"���Hxc�tV�{dN�QD��شs����=�7��领Ύ����=��WnAdd��I���"���Ȅs���9f����O�X͢�ʈY�hB2���s;Z{��ۊ��X1����ZO���'��y�ɅoMv6��DN�da�չ��4�]E���=���cVx���;}�=7��4:�&�>'W�o]���$<�U���,P�-��Rơ�c�%	���.[q��w�sߋ|]7;�r�|�9{�&[�mekW򿁞�N~�_�W�i{��q��f}�e8��O�<R����?щ!�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_dM:Y|����Sp8�<�@��N��Bp�^F�Ο?a��z̵X��D9�����$H��!��=���3���0_Xo�U���r\u�
PCu��
$W;�H��b%`uU�XE(m[��7����������@�)V���d��`��������xB�YA��?����W�^�D�����ڳ*x MW�w��<���vL��rnO��ħ�`�4�&E��M��r�=���ċ�=����_3�������O����L�����E�M����dnL��5J����6�,F%{��;��� ��z���E^6���{35�C��3T.-���3��ǡi�i
�XEJ�V��ّ��c@,k���E����
Z]p֍���2:-s~g5���^q)Q8�T�F�*�~���7zNDb�a=mը��&��-=Vy���ǃnn�o��P�t�Ƨ8�����M���`�Vx�;ix�څ}l����4� ���8a6�ZUp��h�{�Br�u×���O��f��ڨ;@�^bB�i�Q�[UQ�l�r��TD��~6��Z����]����F&'�<кͫBgV���f�V��ߦ~����8p��b�$K��J�|�^�[`g�BK��}��H�|��w6@+8Ұ��$2�Y=��v<�k�x���v�C# ����6��	�)ߎ�-��z"�7�+�C?1`u!(d�(}��T�[_n������gaN�rx�f�Kf]w?]���uF�Vv�t�"�M��x����ǫ��#�{�#_���8|�ߑ�[v����6��΋:�
��Yo�7� �	C�3t<��G�.�O^�p�����=�� �WMo:�Go����P���vEV��~e��Ɯb�/&ҁ��H4�����1?t�v�¾��ݑ��y6	� ���Q����c�=_b�;a9Dyv��� �p.�^<-P�ts��h|n�t�:z�i �dT�yM�E�	��;(�`��d?��'g�Sv��.d�J~l�=e~h�+ ��~D�]�7v�k��<6�s�bV����� � �s����i�Y.��:y�B��?¯4\M�D^�1�� �kbx)Ƒ�+��V97>�|ř�:_R�F�χαO������v�Xx9���nJ,�3l��[J�����DiiKo/��BR�~��	�I:[��rǔ�������r�G�L2'�t�V�]�mO�hgq���"
���7AN`H1N�\�,:L��Կ��e1�&�s�P��԰��Ƶ��hZ�ǜ�ܞ���Ð�s�(���Q��@kP)a�����@=Դ���&���Y;��g�]�D&���[���EfO�������#(���_|GY��E�9����󃿐vN+�Ttu>��ז�ߖ���.��!����88����ܒv��	�����*~��lO�A�2�Y�eX/�PM��pp��qn���y��k��73;4�>u{9�xa�7��e�N��6^j�13W��-]9[�s��6��H�T�l1�{�+�3���9%�a��[2s���S��i��kZ< }�o�-5��LO�S��n��2IDֹ>l��J`g�&�Ch����׸3��d�_Q5��c�@����)m9�L?I|Ͳ�y�.��=$U��.F|ᠽ���.{����Tߩ6��V�#��.wt ���J��]�B�����ך�W��h�x[�%��"�;��-�-3� w�^���e�H��I4��k��ӕ^�J�P8��6�����7a�s�/��=�T\����ZQ��I��*x�]��g3R�[�?�}��&��R%��������d�KH�HvK�M"KVΉ�p�"G�R�d��������n8���%�c���jr��5�ɛ_�У���2e��f�+��=>�6�ml�)� &�N5紏Z�J���W�ѣw2��הA~'-xU�3s�	l��3�y�VV��F��-~{>Qld� �%��hI`>�l�@H�I��~$�r�O�K6֠.J�5�	"��������m<�z�x��PfIP��0=t�k��r؝4�3�a�v�zK*H��p�%���t�M[P1B��������J��Sj ?y��C0d/�/;����ԥ��c�&�_(��i� d��T/�
��+�ڲ0����t��tK� �O�ɨ�FF;u*'}����?:.$��'w�tGi�䍰CY�����Ńn6it�u��|��͝���V�ڮ�"u�E �K�j^��p��� u��a�n����~�ߋ+�i�{�*�/�w
�:��EА9��O��'P���*�΋W��%���{7�V�Q�v�HP �vf���1��`����L���7��f���.	��G�l�I<�?�]��q�q�9�Lm�e����v��Q-��`C������׫��4o��MA���#ܗA'��_���2a�q(hGn[�||L1��aiOU�":2��
��AFȗc���#Jh�BhY�vn��4��,or��07�h��eWtH��y�r�!d5�皣%������k"��l?Q�z]�����N�*��J������R���l��pb�A�9�Q�"�D���e݉�
��*
��e�aP0(��{����������]Ŀ��!�_�$�rg*Eѽ'Ѐ^��g� i�OK\�O��u%
.H��_b惠竸Ѷ�Sh�1l��x��ˍZZ�|A�7�),e�P�}���I�a�5$�o����8/��1٣�����b"j;��a�vRf��"��/���v��Q)�|����o�ф�U�=�,m�,���{dD֗�4$�Ui���)�T=<9c_��V�8���(�\Q�g�0n��G��4tg
c�X���F�6����u�g~W��bh�u��|��-�Z jT��C���l!�J�����8�;��la�g"��}͕����)���!@�e6h�~p=�Z=U��I(�����C���s�B}}u)!�yN��{�z��6aU�'�8�ˍ����M0m�8����Y,�� m�{�͘i�"l�-�:�����͕�E�c`W1doL�,3�c��	v���5��ya]�x\���H���,���t,A��m��Eu��젤¤sѫ�o�f��[��;���T����^![S9�<E��g}#9�y�wY���t�]��}��7�o�q#D$�}O\�)��$5��s��i��$���j���SG@�Ss-�K䊯!B�"N�Ul�r6�K��l:ݎ�$�eE�Y�P-�۵���T8����/Լ;��{�#����|}�`�9��d�`l����
�q�f�Ǩ@����
�|�2%/��Y-��xb�r��u;�˵[�=�l�Ya�uÁ�X]���P���A[�f��<�P
x�k��UM��\���,�'u�5����'����	�B�ʌ�L.HWB�x�|�Yd[�!途��
D#a8$yŰ�9&����l�Q�i�3�nZ�lC�Tn�Wq}�X0n�����(�tGo���"9��Z��8Iw?��Q	p��-��R�����55;�9�����5�ƍ�8I�Mj�*�I�4�7X��y�9;{[����+�&���v"�#����޾[�r��d�����m�U��%�HI�G/��cg})P���2Ihc��~p��@�x�|�����,���i�xB�$��}� �k��^)%,\Mi��	иL�J��j����lx����9��M����Ld!7Ν�)��Ƹ� �3�'R Q�g%��
������\���Ǹ���]=�P�N㽏B�,��6��}$�.�<�Ҧ<�8~�1|�
�Q-	��Lۦ?K�b|�Pr=�C�F��{�"����F�T���M�3�<	�+@z�9O[8ڻ!ȴ��$ۭT�R�rIJ�{�I��?p��Fc�F��]��?z�	�P�W�d�\%��٧O����o� ��QxM\�@�
���V�
������>�8k �"3ֱ�bƛk�ןG�s^p��n0��H0>`�x{y�	09�|��M��|a�>���i8��f1���^(�B���R}D8�=4`�YZp��(��{���%׮ )?��G����)�8b�#�dpӖI��p!n!��O���.�Vчc!	A9"³!3�X��_ ���`��HS澔]CV�7��R҇9�����u�ag?�5�r���R�f�a���'��)�]y���}��O6[�o��4�NJ�����$F�z�,[��I���d���Jy!{�����|`�P;fs�/�g�"f�R��ؚMg{/�_8�N"6�\Y�LxN�:���!U�X�fayU^�<Ç����Bێ�ky�@dK��v����ΐ���|eg�쇗������8�I��LZR��Q�)��`��������eC�1�H�	����s�FS���+ݳ��s����y���DA���7y��o�Cg&� ��̎��[��q�������%�F����{ZD�kq�h�1[vF}'�?I�C\zWW���������I���;hLe�nͧ�ͩ���\f�zhR��#D�t6��&{<~a�N�W����v�wn���c����S
.یD�^I��j$��ڃ�I�:&[Zߡ-��Z.�D�����ˈe���;~ �6))P|�J���`�zH�
����I��l�J֍�!
B�M�5�����dbPv�L|�*����g�c��R���K���O��i��ɢD�z��U"{�s�|2}��ͯzl�^(�h/&h��6����� rߤ�m�	�	�eq�к�q2\3|���q$�5D'����<u�V�Kf�=y!D�E����Nh�Y����%A�ǉK�B2���%��N���S�G#�!`�[{�J퇨񽑏�PZY�iG�?&K���d��Y[ڗXA�, �@�����|Ŋ��v�=:ynk�����t��:MQ&(AbD}g�d��27��T�M�D�/SO������=&d���zg���p�Rh�b� [��I�%�L>�/6��&��|�Ϧ�=�N�K,�J*=��!W6�4	e�Q8��L���l�"`}�/vR���5M~h�O�8L�4usW����]��sޠ�4����'	"w�z���X��1�>2���Œ�k���ب��ׅHyӐOh��vߊ��eº��4�5u��9(�㽑z]�<�Ǹ6�&�)HkӪ"5E�%tb2H=��)������mJ��.�?b�d9����#["#��%lw�~��Q�c�1��|��@��:fK�|��4� L��ۈ���4����/J��.�k�l��h�eM.sS�d�7���3���6b!8htehk-�L�Y.��ƸV�e uR���\���eU]��h��"��<���{W�<���_P����īMf��vSY�i�I}���ڍ���$��fv���ē��
��bX�} [�Tr8���9[�g���!
���<{2e�Bmݶ�^��sȺa��� ��f[�%��0�#��s|<���:5�Ū�R��Ҡ����{w��v�v5OZn�x��*q���}eKqak�P�(�W��R�:��w��E)��iғD�7���`�ax2���4_f��za��W��^��Ϸ�
�
��
�$ؙ`{��rao^+/E���e�]�¦�$Q�eK�B�23 ����h �1�͟���ڨ-q
2�.��i{y]pT(אw��{��/n�AE5������<��Dt���&'��� O�U��9�>QYxE�E{B��Spb�+&��`���ʋU;_�pS3t����9�ԧq�d �$����<{��Bİo�{K�0������֏�<hn�Q��N��V9�@H��~M��gp��y�z�i,�寧H�9z�O�*����B���o�$�+�-:�[���7N���6]�d��:Iy"��@����|��˿60@%H�i1� ��"uzS�<�^�PZ�~��D�+T֚�ΆO�pe�
<5�4V����cxs?9�̆h4�d=�X�!D;d��a,hp�?Ř<�:��maD_q�<���d�:�ݲ�W7�$�
���6��g`�n��XV�7��$�S���[i�7�:I}�T-/�}�'듄eC���􆣷}47��x\B��e��IrprD�[3�|i�M
�>��� �������l�u.�D��yVc/:�d�4�T���dkLS�8�毻5j�)!�+	$�ࣳ����c/��H�Y�1�C������Ҩ�n��oDl�	��s�J��&	�>Xo^
Ѫ�W�
��w����|ɯ��W���b��s���M�@�<�`�&�}�xa{��"�kt��6A� �4l���
�2jڮ&��Qן��^V���
:B�1���9�M�X
!��1d� K�d�GbV��.���5�kF'1=���f�J Q V�(r u�u��mA�xh��mN�۬�rO=�?��LJe��o�܋�/�-�إ1\>دLc!il��*/s���UNް�ukm���K�OR���3��B�tf�>�p� ���PM��7\A��㴳"�*�$:������+��+mp���a�C�K	X����&�M�2s�?����1j���.���Q+���d�.�͉+e�/+������@)E)�	�|*�b'�GH�yh����Bv�2��{#`,l�lC�}��'��=�/�v�ƽ���S"�6��� CBE�8�i(�dHmU@J�Vsנ;��k�]��bE��ɵ�ƒ��|�h�q��j�QGE*t�aAc��fq��Ϧ<�Ҿ�>�y(~�˓7��&Rt|�t��2�2c�	3qu^!:����-R�I0��E7s�D�K�g.��eKt��ZbOi��2}����t{u|oZL�$�"���+S�2tqb)���4I�yf\]�^Q����<����Ny�E�Q˃J��l;֕��8�r�/,o�]�q1
~��U���=K��љS���ʚK��kA`�{|ZkgT�iG��r@{���y�}�֔�tj�};-Z`�OOlO�Lf����҄@��?���=yC�=M�����o��^��Lv-�Bx ������!�7��.wz8�h/��xV�AB��A�?�XG'�b��M�[�k�`���N3���C���D�V<?���
��:���ݚoM��Ho@����^��i� ��$�	������4;�!d<K�"1(��X�S�>J'�K��05���Bإu�E��@V�0OG�z�a������Y�Y�����f�>�X��9ˊ.�v���n��(��Elo��W�>��:m��*��TFB ��=��n���n`�f����*ۧ-��5U*� �=xK��h�A�w;G0�i���,e�*�B
�v��8�Ć��-�zN�VΗ�@�f+���q� 
���B��=G���m?��Y�K�&�:�9�3[=V ��r���cJ�tc̻ �����=���O�h��4���K��{\Rj�m��,��T7�|W��N�Ҧ��5�H?��86�u�t�?���G[�X Z����\�EV�@�FC�G�=ΈEC�{7h�;];�=I>b����x_Ag�ج��! ��ԵG~���	S��	R)��X�Y�:�g/!cNfRx� X�-�	��m�X\�#I������FJ.ґxDf�����Ʌ`�ǎ�q;�}1,?��p���C��0�p+�m���#����8Z*J�]�x�|B�o젧[zh����B����l1D��Og�η�I*T�*iʛx^�?� 0��s�Je���W�����(n�!V���0vN��2[��wyx��8&�������k�Q���')u[�A������w�o�jŴ9Ŗ��FT%X� -�f[�kԈ�����^ ���>���5y4m�S0X��e��l��\R,����_!�=@XU؟��+���ī��J. >v1��= ���hI���%=<7��FB:�O����q=!�2���@�8Mo$�J���ݶ�{�X�L��Y�����&��]��gQ9�3��ڻk[>�A@��u����@���_PK�L��Z����gR��Q58G:�s�7���s7a2cby��V�tޝ4�<��$<��(����!�("$�
�)�q+9q��N4q�bwwk/<�( ):1��-Aj�Qv��~]Z^HA�"�^~Y���+� t	�mQ/iN�pG��ښ��*���0C}*�z?t��Pȝ�4�`4	jk��lM�Q��	LM�$m����VH�ɴt���/	�����r��|�Å�F��t�Ub<u���K�A;Gx^���8Gߩ=;5�;�j`�����Hܙ�LV����mM����p���@�ܥ�ŗa�'a��يS؎��]�i2��O�����)��(�է%���6'*<�J��bm@U��}HH!��`�gm7o�ȟ�� �s��	�,�hه���/ƥ.���O�t�G��)<3Cs��Ȕ{zs�O���@K,k����~])U���_�s���6�,�e/AL�{Eu�����//�J_0�؝����lI��f��@�HOk��ΕX�� �$���^*��7@f��R>fծ2%��.md7��c.R\�䕶�����6�7=_yߌ��`��7�o#�����߇{���#�ML�`�u������p���>��T�m����!���g���s��r����$�X^��5ogsw�	p�҆�s�L?O���2xb�;�މ˧�MI|Ա�D=��w�7{��/�F���*��*������C�J�����1�k���c��o����2�v'VK�\�&ߓ~��2&��8��v7Eiɍ�_�L��}��y9�~�����T��&���R\�]�wl�>�!���k��$(�����~�25Np���S�k�#��1�A�JJ�U��㬗�l�Q��٩�V�\��zD�9lC{��*,g�pNx���2���T�NX~�QuUq<���H}+��σ�n;<���n��#y:��͆�i�d�n	{@�>L�S6�m�L�{��(b5���ѹ�'��@�T��_�aU#cC(Z|����"��c��r�y���ˌ�_q�5%z��w|���+~&�Wc���1��Q��݂:l�~�[����ZxE��y(��H��ŝ�<E��譙��B�Eh�:|�s��*_^��������i��R��Ȑ(�A�5O��f´���A��'��7X���<�?k���zc[�T��Q�����\|�����G����I��n[�K�JQ�H�g����gkd���v62,��e#����Fb nO��˦x�d@����?����緧r5��ghH�O��m�?PY���r6�.Epi�z?�_����J`�\(��Do�؍^7s�R��#���J�^@p�c�`��}s6��Ih%pͨA����u�ۆ��|�d�L�nl�.KkP̰�0��H�9r�_2De��K ��0듃Z�+>z���8���!ϐ�	���a�:��0��&͘2Ve��lWt,8���$�G�'�;�
�-4��)�T>}T=�nlIb�'��,"��3d���V[VY"�Ѷ�&[v虇��adk�@�m�c�� T�4���ȩM�)B5��/�6���o[�Xr'�'�r�1�����`[6�/�܍�,\8�z|�}((9ڧ�5�s�smp�_��ɻiA?w��J7����������;���Te"mx%�1m���4\���_��K~��/SU�S���e3��O��P�r	�^���H?�XB`a�g���D�h��o�?�'o�]��%�k�R����D*���%�Oi�pK�	�e����%h�1(����z+��@'�{M0�m�Q��)�>��������x<]��4��З�(z��hD���1nh��{,�-@!r������." ��-�AW������eg��d���e:��#% ]W�����&h�<�A?.U�`a���=}�3��H�H�am4v[ߙ)D̸��H�f�Ӊ���(�	�"[��1�e�Y\-K�ņ�o�� ���5wp���z"�F:��w��r~�-��wN�rzb8A5�q]淄$��5���T3��[LX�&��[��A@�]ez�J�:�V������2���G_���� ��[܋/�/P�
��݅��ǚ�0X
c�d�P� �����TEҙ܍��P"߹9Xp��;p@��g��)7f �2@c�C�Yj��`�nۃ��a���9�5"�PB�-����G��P��l=�6��2�h:�F����F��S
����8x ����f��ĭ��� ���Жv���̪vBZ�SJGw�'��+
-�<��|�|���T��p�宋�� �e��S�	��X��{h��w�:�͖	^C3`w��K�Q�����6�H�FƯ�4z��j����uN%a�v/U%�% �bd�r���z���`^�s�/?�q��c��y���քel�:���iU朰��@��(q�X��7��d��Ft�`�2�;��_��-T�h��zϜ%��x�</g$���S����a��,XXRl��I�2��H�A/�4��(�|�G0�!���T�}ľ7:0�z��e�6EF��f&�����	=E⑍��]��-��p�+��g��8�VŽ���fC���}e�y���*�����oU]6��-`��3#x���>3(bk���F�Wێ�֭u�eɎ�te$	����Oޛ���[͠�-�2��ai��¸����4�y�bλ�(=�*�H]6t��o��0W�u<�����(��D�_���J��>���ǰ��0��%�5�t�i��5�V�/�N�m� �]7/W���<������G�\�^�\�O�7���R���N�ȃ�:����Qj"+�K%��UP ��Ŕ�:o�w}7
���U��:��2^�A�|�Zw���¥�mh"uv�ļ�!Q���-W�+w�$
�H�~.� a>����
�c�j)�IVE�$�N��*S��;~�w��6���ɽ��(��[���� G�GtZR�R�syXI�P���.3�����V��O�O:�)K�V����*�x,���7�e�ʫ���a��[�W�����&O%me7ߖ���=�5|���8�����=YL���ÈY���۱��=D��O\�bx����(Sol!��A���;�}RH������<���UԳ��X��}h��`�dc 	�K)!�n�6R"1�hb_��h��~/�DY=8���k�[�O�E8SL�2�	51�זr�cV.��}6z	�*A�9�#�d��CL���Q�Ÿ+�X��z��1�Y�C��uJ��Yk%_f6��t�X�	5_~N��6�5��%J9��t�㚇j��!wy����nr��\c$�tB�t��/���˜-~G+�2��9��8P�&>Dl�m��q�l��,�Hk&$�z�E��Ws`���.�uF˵K��0/�Y-&���_��~/�È�%d�8T��J�y�%��Jsi�}�ہG�;��ݶ72t�VGq�u�P�*o�"w;�>u>�p��Da�3�!s8c�&�x*ܐp3B^5�J ����Ld=��~0�w1@�=:�_��2��L������q"?�ץpO=�a)8�?ri����(�:���)�DJ��I �2Q�<��G�+ M>z5�~/��XC�T�%�ҿ*o�㊃�����Ҍp�+ْ����v�6�~�tBN��D�������b�&
��z0PN
�	GMύ��0"���������n�$c�Y�s�w�v�K4�I�E���j7�=6����Ќ7��p���8�~����rH��V��D�ف�d�<�x��DO}�~��bQ�v�����"�f�U�T�2�!y&�1!\���uX���h���-"�@�z��к�|4$E��ĭhU��pWS�zݎ��I7*�?�:	�9�����v����DQa�$��SU�t�}7)2)Y�
(��!�hag�T���3�Q�Z�H�06y%�����\����+Ŷߘj�5B��,��R?w��Q�o�1�BU_%l������S��,���|��E������;�^�9��X��ڢQ�>�dy�.�W@��{�:�\�]N�K�r����ԡ��w�� ��k�w�����Z@]��^�:��~O�s�z�}��d|!}�.Y��0�)	fƆ�d`�M=��6�߆���j�b0I%w_��w�@(����e~�ډzĦ��P��:�	�Lawx"�cԑ��쥉|l탍g*� ���ݯ@Y,�'���9C�!�Bf����Cѝ�g;�ĉ5L�~/��eTW���)�d.8���Uj�I@{�(�,T��F{��/�JQ]nr�4٢�8o� ���渀&X"����������rj2t�9�4M��/�X��qƬ,-6��zaV�B�`,�b|B�15�A�}��-T���N�M��>9p,����&B�@#��C0��R�G��f�$z>�!����\���H|{z�������ѕ�;�*��N���.�p66-�KZj����3u)uBr[z�G�J.�x�����Z���޽�����DLEfDr'�q�Ў�	���Ԗ��4vRw��2��h2���:]�k������*��WK�<�^3U	�i�!<_TPn��#G�Nq�8�/��{��Պj����G&A�i|whD!�֌�G6S�O�;^l�N�h�8��<I��E<{K��Ǚ�7�7կ��{!dM���55K�@��Z���pƎ$,3ݶ }�r�:�
��5���	*��"o ����
��o�A�E>b��A~�K�f26����t7w7.�z�Ð��,�I�q�N8��D>�?'�X<�?݊�J&g��Sʕ�p���K������_�nь<X ����֋s�d�p	���-�]��EΑ��o���L�s����i�6_qb�F�e7ߕ�����{U�v���Y��~l�A�HVC:YE�2�O`��F��~�a��ԫ�j�� �zk} �u/%BT���XU9����#�&6�7�I�O�a~��;9�0e����=P����=D�3�cح��4e�6��W�ފ�B��2&ַ��ᗘ�L�С�o�g�Ο�&b��8�@e;,ٽGJs+ �g�L8j�*��~3����{GКO{��!"�M�?�Q�#Y:���Q>r�S�ߒ��`���nƂ]î� NX�-}��"�;���R�}�����Q)��~�Gj]��(!�G�B�g���g���X}��p\�fY�5"��HI3~v+M,+rmNY��N.�e�~��<x�0�L:���ZS0�NF��U��`�!��ᘽ(���mV[��~�AR���Z�WN�PI�N�,�1�FC3@<�����af��`�8��v������L��������E g*���B��Ad2K���+]��ғJ ���S�n���xAê�$V��|]"�ޡ��7lg`�ͻ+�뛶o�0 ~0��9f��J�� j��-,���!�߸@M�ʗl�._��MN,+���$�9D������(��䎬~�fK�Ɨ�s�\[�i]2۷0p�.�I��mqZ��"�����5#`ͶV�4_�CS����xp&d�`Ӏv)D�UJ�v������H��u�G8�H���iZ�Z!ᚬ�-$O�s��/Xv"�b�ɸD�Qrw�(�� }_l������Ao�84�G��Ԍ�V n� Ԑj��|���1�j/��+��?�xR�����1/��q���ҹ��B"���6`�w(pM�'�(r��;.\��Sq�%�?��
K�Ɲr��˦���h����ӅUu����=�b)Y�k�P��F�^��Y�K�K�YJ�KKx0�|L���}j>�zlX���$��ڪ@�Q���-Xiz��i����ِݦ�j�����,O�(F|�
Xy�� ��$��6W.4$t�E7O�J�6�V��΅9cYj*4V�!��o*��FK�UNmx�Ԃ<��Z�\'�?xG���Z{d���u�<�i���BN��|2��S�6��[@�w�Qfr��ZV�IK�J�-
P�S�V@����cP^jc4-�e޷����rc���ǇK�qIW0�;�t��7�\r'�|�(T5M_t��y�6-1#��6�LŐW�8�y���4�T�YV�2���J��B�&�;z��9�qVIs3:q^�#ܼ�^E0_E5S_
�띵���(V&	ǩ�u�|Uw���9�)�bMx]$�R5c|�!���V�qw��	������.q>��L��l���J3��ǈeO�Ѐ�x!���.��ц�Ҽ�4MY~�$Yo�c�ܫ�����C�ꁍ��$�&"ϝ�:i6L�(Xc)�+ �d��M����s���;��4_U!��U�>�y�*�͇��w�iI�� '~.�"�kM�D `���h_i����[a��U(ƋD/�=�����F���%|��W�u�!���������v�m��M���F�8�����t|� Ї���|N�����Eg����q�$̲��?���oJ�=�"J�_QDKd�*�HF���� K��>�
���wQvfD���P�L�%<tX�C�+m�F�-�&��;�+���,Z�`�2%FI��q.���e�]ӝ�oR����3ß�%�6��@�W85 Ɖ�nۚ��e: :��z������gnu��^LQf�<զ��bk�{4��uH�2�C�G�h`��#�i�; �H��Oh3"�MA_w��/F�4�xt�S���pv�#�Z����ۼrU�y2�>� �U.�� ��bI�Є�e�FRC��e�<��M�(����W��:�-�<�%Ǹ�?ʵ����4���'πF�fw�ma�ua�y�(Y.D���S��~�{�`� �d|����%�u�|���ESQ���	sh�?VO*�ɍ��D�m�#hPf�y�3uB�����ӓ�CV���W�_�ZDD̮n���^���^�� ���x���=e�N8��(˓l����7P�@��M�\fC$�GnV&����(
d��3suߎ�k}���$��Wy��W�\�e�@����A��U��/�<@�A�Hb�OV{iK �
�B��K*���XU1g����x�V�jf])#�`�����G���o�\��%F"�J��!y����W�_OR^M8��l��d\C�C�y�@���@$�b΄֥�Z��^�n��͡7��%o������$���3R�`��c��#^��_/�L��^`Bf�:#?9�J�i�Z�m��6T_���pZ�u�g�p�˖u��8-o�pinݚSb�ͅI����-���L����L%E�ySuk3�ՙ������LDB5h�`.��k_���}]�"(�=)�;6�E�fs��M�a����L�a?v7x���xˊ(�0g�ZNԵ�Pl9�l��.^/��=2?$z<��������r3�Zo���E�(��?�s���ވ�������f5m4yer���O^Zt��
��,�+��A-���@����X��z9���Z� Ċ�pl�Q�7[��\���wI�%X��IYN�6J�J��j�л�|>b�j����_J��?;���=����jvU���p�J�L���e`ۅRɾ/�5������>էa�o5�9̱��͠i���˗]�̤�!�<�_"��H!��&���b��������`*��D���ߎ;�5���T	�sM�#��6�L��q�T��?�W���x�Z��Å����U���Ϲ��\�+��ɂ|g���tbK"s}�g�XM	�'B�-�e�1͠�a��A�pri��I~�y��*���A�c͵����/���<�(}P����Nvi�x zH#{��v�J���/FCn�����8���oêaZ�j!��S�]��x��;�X.���6X9L8�-�ZfC��HB&Mܽ��6݀��48�it�+}C�0G�3� }�@`s&IY�u�,�n��\��r������h��̓U�Mli���4�	�B�	�ԓUV�"lwa?�W�"��)��ɨ��&�u2��_�RO�J��t�q�]�����'	�1S������X����-���a;(r^ q1g�K�Ԗ~������Jd���{a���PXO_�Gb�"���
O�^T?�"p��4ںBe}�Y�"���^�e{x��%Oп�`-��G��r|���h���ý��U?颉ꖎ�N�RpC�ɦ�vBb���:��XOJ$��v:�u�gY\��4{���l�m�����tn=W��O#�<��v�"���;� P�縌�C_|�����ez�u�+.ǆ�C��R�F-D��!O��1 ��X������J�Th;Hd�`^��.I��%�u'&��RT�w��e���g/ȝ��U���ړg�Ս����/���H>`=��VI���OG� �,u:���۫�N��v$:Ç� �C}��L=�}�h��!����2!Kw�EU{�2�u�L�@�o%� �U!�A�xnkO׍��p$P><��I�O��^�?c�J��цU�-�� /�
�7	q�NA�"�p��͇Q��=�/��	\��{?�=����l��S�HH�#n�#���j��ݭI�Y$���0�8�dS�3J������U1����x����A-���{>q*;��|pOѸ}�hU�|q��3�nb4a��tj��4���Y.D��,-��jZ��NE���>��b�,|e�Sv��R5�E���q>���<�s���w�cw�,�7���xKȫm:�Jv<'��꘴�`ieغ��U�����Fq;�)�V&*�����?ɤӑH�}�mo��n��G�'�̅>���P��>�,YCÈN�o hN+:�����劤���9��\��2RWFBb`��e
I����EQ�W�;5�P@����6���9�W0��,_ ���H�i�ʁ\m�ͤ�\T��X�=������OLFy �1�>Sq�ڕ4 �H��T��Ė��1��__�_�)&1�{� k9f.�ѧ�-�?��0K%�:,f �3�zpd�6�Q�Xwrݗ�*�(?I����{�	��OP74'�e���~'�y���eA%�Dk�,���t����'��"�'!��;����^G��E���d(̥�:��j�)Ң�"�����R��N�+Z��� j�M�LXFa+�%���]
���@u��Hĸ�	ڔ�2��e��Ğ~�G�]��C��R[�>�P8�8V�%�O ��ݢ�4�/�&-.�}�'�Ӻ
G%��p�=E���eK�J����c����8�f���"�U�<���]�.G�v7h�no9'�ا����1����W6H�F.��PZ��T��U�Zh<�-���
�ω��a՜���  ~�2��j�j�^��&0]�y����l�Z 4�M���V�q&��U8Ȥ=�c������|�9��r.�a.-il���;_m'c����LrC�/�ӱy�� �m�a�-.?���|q����>�S���d(ݞ\�y��*�����˱U�����$.*�0O>�;�<���H>_��Фs�?=<�; !�f9�i��7יp U�$>������L�|�O�J�5o�����3���$kw"���*Ti؋��H����)^J^����鸉Ym�5��*��k9�$�k̀Ӊ�L�R�"�i������l�#< �� ��]`'��^΃ig5lIY�b� �9ՄR6h�C&B@b���C��l�) �g~*n[;��	����\;�z<���j��s@�Io�q��'�=+�m����Ky\�@��ٖ�^c8�u�!����c�ߏ8q���a+6��QWg��4�<��p���,N7�Q����U����(�u���4��!B4^,���}�Ұ�^��]Dv��lG��GSZ ��{�0vr%R�w�$?����J?!TU5]�?��k^�u�J�H�Uֹ[���=�|�X��b|���Bv�"wK�:�*f��N��7�2<S��' �A�Ѓ���/
��,f�F��\�:�EFv��@��j��vn���&U���˟�ވe�K�^��;Q�4S�n<�='��|�̗g���TzG1���#��Ƿ@%�T~F�7� ��6w4�_�)I��5�n�k%��]�v�^Aܾ��Z�r�Cq)��&o*\��� wGK��a�X��*�(!R�[r����%o�"z�����]���3��(f�aUYQ�濢*S�^t�ꊐ���{&�⸚Y�:pS7?�pige����!���)�64U:6�m}��y�+�p��x�Oc�b�c�,xg��N�??6}0�T��m�rC]Ma}�)��˟F��J�NcV�_2)�v�X�-�D^u�N����-C?�Na�(�O���P�w���k�y)����s�	��#��~�`�v�%��+n���u���+#�x�ʶï�����"�hrh]� �I����q���d�[Q*�&%�����la�$��c٘���6�.�<����&��a~�&�a���>Iys�r��c��=��^!_7I<���K��xR#q64M�k����haE䌺���PޱV^8�v�B����3R9���V�vL�#��y�b�sGxm� �h���� ��?,�����-(�� d��q�lө��u����;�C�>rh��z��BZ�Ђ��Q�c�{�D�h����8n5�&Q���9���ϱ�"��0��7l�ʼw�\�1v��`�xV��P��܊����9h�@��P��Ջ<!bŐ$���`�ٯ��Y�"��l����Ul�.|X��$���fĭ�����V���^b��Ű~n�߷vi�%T��z\�*�-m���o���$�^ 0��;��I��w���	��$��^끋�K������z�E����.�{�[�I���_� �Z�tK�1��SՍHz��2-x7oT�n�f�:G1�l�(��93�#���3pp������~h�C߃��J<�F^���|s��t��5�PW}�<��T�9�c.5B�J���1�&7����.�{f`Ͷ`L��@g���z)_�R���ȁ��C�`S��^�ۦ�t�k�p��Q���PFiS��{1%w)��+�;�VB���3��aH����ʥ��>U��v���m�WEQ�[A�l��ˈ��V��=������;L�Q��<�-?�N�H��]�7��?�Y��1��g���3-�B�1�ɑ��G��r���Hh.�L.v�"1SN[1`Ț�B�9�������O�:)ML�z�R^�?%=�R \!�{���`��P, W�<D0<����M�rt�iM�u�0����&�g,vڏ���v�b�f��-3��%+C��|�H,<8���wy����p-�g�ԣ�"�ͷ@���Dcr$=؃���%�ڏ�A���-��H����J�@d��۾�W��7���49�x�A�:rj����ePt�s
���]����;Kw�U~���D6!�{��d�jlO���Y�_0o�Ğ�))�,i�5���˵	�6�E�V"�XB��v��f�a�2fu�Իi�8Px(^Id<��@̝9�J�2kټ���:@��J��`���?:Ւ�.q��Q�j�
{z���^g	q΋$�d5�P\�����o������X��6��'T�O�S���+�rJ�-ES\J�A��,YZ� �ƴS���Y`�cv�4*��kn�kh�p{����e��n� �f�n�B�A���7�#���R����O����R��y	�o���o �����c9!3�0��[�����U�o����Y��}�����3�B�l��"�ʊ�ꀌ��[E52���"�����Ũ	����y�5r�$�ݭ3��=��+��B�Z1�K��ye�$���U(? AM;&�8��|b"؈��w"���C_k7s��@lK�$�6�`�?u*��8Vp�����)��o�/Sv䐃�(����~��x�ə�hk�MHW�/�t1�
.�M�/-�^�u2�Aų%j�5�5j��±�;K��`l��h�х`������+8�0�w]��05l�~�N2i�P\�������+j6~��N��	#|�3�FiS��ٕ	ĘSV��z��L�s�z%Ķ3)( ��d�X��x��;1�7�!]�����e��mG�)��m-��Mv�ے�Hq�ے��'���$�[g�&V�LA,��;m�#&͝���b>��_�+�\�|�Ɍ����� ��W��so��s�NQ�pa��a��?$_P��/��4��W��if��j!�)s���J���iҡ"�`��	��O Vxi��HW���D�$�N��I8���Q���s�@&�a���b�/q��`�,v���=ͯkjnB[�e��u=�W$���AAl�������z?���jCVc<�f�(�������b;i
����E"e	�M� ^�y���bΏ�/a����*(!�߸mʟ%�3�>�9_��uN7�=��T/����!*�Y�Е<`cb����������x��}9P}�N�H.��r���qP��J�[��`��D�L�W����Z+'�"z*��v�4~�
D����
��]�E�ER�W�V�V@�.��7+�<�~j��\���W��E��=2-l�^Z��~�u53h�8�6�`\�0���˝s��7QaK���#�GՅy7T����Ӭ��X�K���ss) 6��� �czR3$?��/�"cw�D���Hq"���D�X+	Bt�c$(O��!��7� z80L�OҬ����fy�~!D�L�p��ײf�;us֜Q��l�C#Z���0ZT�=��<~0ܫ�;0#��ʇ���,W��3���.q���j�2ͲWOpQ�h!��FG+�Ŝ��.`6�p�W},s̀�U�xD��@�wl���HEȕ���c�eu+��]�:�A�����`T��$1g�=�p�~N�1I]w��O�.�aӥʟ��pxԤ/IԤ�tz�9D��=���D��shu����~�$iʛT��~v+\�i9xo�$Ca�.�FK3w�G�)���1�0�P�è]oa�9�ڹ��:8#�t���[���=�!R��k.��3��v8�,�G���RoOj�<Az^P�cҘ�b�3�@/�C(K2/,�H3���NJ���eƽ�Ɩ�������[��0[�A�~4��0�B�2�x��\�w#W:� ��}~���ڞ�b��o��e)f����[W�e���y���o�+���7!Dr�H;!+��=f��	䀼�������J�W��"��柉�ܬt�n�G�����ip�`,�lo,���� mG��4��p��S+FҘ|
+��8��:ǯtG�Ӡ<� oO���\���xd�0��ܾ�cQOչ��A"ļp�_���!�.|��Z��H����=t��Szܗ
���P�y��c�b�y¢C��I��b^�Q&`�]�P>��$t���X�)�����VH8�w΁��׭g��y
�[4*�hr0ꌧ9݄`Gzi@j{Z�k���P�äb���0+���{+oiEj����I���(G�tӸӰ�B\\-�cU"�A�V=�W���"�+s�jM%t빨,��I"P�Y0-7���E��Bm������c�1���V�\���`I�BN����/,O%�G)$x�S�7�_O6�A��^���:]�^1�V�kg7�rݧ,Işc"���ǘ�
J���-�\P�Zsg6�M��aznͺ�����t�kGz�Ǔ�
Ą}�S�c�r��#"��9��C�\�X�愍}'�~�%)���X0s�:ؿ��X
U�r ~�Qv|���*��H���W�#~r��A'z�|z��w�,Ƞ4w�|ym�0�x�~��U�y5����������F�t�/�&�v��_�-am͐��:p���g�t9��U*�x���η3I�`��wó��RS>3���L����!6&�?Jl������:�/����h�c2��oI��n�=P�q^�����?Ӡ�
���DO.:F�4��B�}����TRPO��	�MDw�\.t�g� ��w�2�l������c��Ӯ2S�muNESO�ad�V�:��d�o�d^-u@�5+}��l�N��V]�Fir��ܪZzNϋn��%1��:k�G�C���vei�=p7C�[3p�,�D��b�� �J�}	�q�̱�U�R����ܰӰ�(���}�������T����^�.��-Q�?>�m�(@�I��K����D&Ԓ���7�����I󾸦	#RO���p���w��J�~'�����)��h�Z����!�۴ߖ	�����^��NT��鵅MaQ�p���QG��	�ݴOK��܈m�cl_Is<nph�K�	p�3���w���(���Ĉ����9�H�{.l�&��l�Io`[��}�L�_��
�[�J�h����b� �l���^��]�T·j����|�_�VǮu�
6��G�[�]&e��j�CY�Y�W�`1/X��{�"�0V�� 1~�QX�:�b�3<*̺�>'��j��<-�t8�[�h���HO�2wn�6���%������%�Vx��
=��yg���6�}��P⠴Qč�;03T����e���nor�cP`9�>k�c����PY����7�d�eE���j��LZ���U�od���	>���9�ًi�j�$d�����20m�i1L�y��
�ql\r��Պ�k��s	�5j, �R�k�=�g����I�6uOC�]r���m��"8T)����WB���E�:ț0~!#�CS���u�.�G�U����{6���O��cS"8�|��y5�H��NҢ�F��?M���Z9��m�ȩ��)]�� VD��]6���w����)�p}��7�n���j/2E��s�
r��������pN6x���i|�o�B��2ŶzB�u�ۢ����BgAb�Lx�,��h�{��d������R?*���*�T��2��M��#t�n#���G���xNE��V"�,�	0�^^�����p��
�{��]��#HC�Nf���V�l��� �=_��u�R<y�-At�;��b���[d��R�K����j�8�1K.zQ��`��J��htr���Wds!�Ց&��K���h=�D�Y�hݣ��
un�Ai�u8԰�7$�t� L���G2qS..J�\�������-)�`�a�
�LJ'��Z�u�=��$��<#{z�#,x���i�R��#���n3��'P����� k���_�\tf�P\%����ڨx��%i/�B��֏��:EA}E�c�,[V-����e�/ �e�m��Y��k�)"�5��[Vr����{$���=u@�H��$�:0��x�3�� 1� �y�����`��ғ���l�[��.āc��QL�����8W�E����.�B�F��!M�ļ����|S���9E�6���8�n�+�W�W@Bm�"�^e�Xb�3�el���¬nV�ŸgIJa�ED1P�a��_J%�|��B��V�FTL�<��Z�d=����,c�O����#z������o>I��(݄�û� ��J4{���$K�c�N@dw�c2	��Xaïb�ɝ��q����;�H�4l	����5EOnR�̐�J��GZ��}�����D(g���}T-�T���Xdp�'�p��8h\|�>s������R���[�ܕF�yd� ��\*���d:�C�����$Щ��m�7�����9��s��󿽋!5Ӷ���^�$�3�����'4%pnVbհ�*ٱPr�C^���"�tA�Wo1l��<{�Ա4��D����M�2�i*9�����!�r���,���i��F�u�>�R3t4��3%L�|��:�zR���O�ǖ��tCC�"�l`�X�z���<t���o��'�����;_�_~(n���A�'�p8��c���^���l�7�'��R���,�}���X�<�5O?eĸK���.�z<s��"�J���*�b\*�>Pl��/�v0����8�W��U����5p�S�PVr�Ej�~���Z����M��\2� {S��ʨb@%!)R������c�5��kn<2����o���Z͉���[ӿ'�Q
Ƙ���	�[�94�x���E�D�L���cq����R�]�k+���P���2l-���e�����ӝQ����AVw�`֕"	"5￵ZE!m����7��v��9�Pց/�}��4.�<�9�T"ߦL1�7_�Ma��!��z$�;W�}/����;Re��8��V��º�/C���U�_�wh�� �8cWf`�|��E��\0�h�T�#>��z�{��� ��4�8�KE��[�O��������Dă�P&�$���"k 2�K���e�����n���H�1]^FO�Z�ɀb���MOn��Q�+tc��W�%R�y5��z��Ȥ�&5��M�����8�2���ԡd�)�d��B�j�lҹ#��?%7h7��?D|�F��$��Čͳt"�k�o�"C5�U+[u�+� �1_����F?w��U˩]�d�����OU��iR�i�������_�a<�u�7�p�P���=�F�΄������ȷ�	�Ԇj�	�χ�g��UL���\7�1/���ü���\�h��/�gߐ��!�Q���N5S�Rd�����2-ȋ�%=�1��u��g�b�@zC|����m��nY�\�W1����;�+,0ף�Bi��tM!��zϸ�-�~.0�ր�s�6�G	O���4(8���	ڃ�+���ɂ�5޶{��=K��o��	P8vH��#�O�oO��+���s2��Э[�N�j��燛��cn���q�A&�I
깕��y��ʂ.UUNg6&�pE���˗-BJ��Q��/��[�&hGCwJ����dE����sκ��E{ʌ�u���ҥ�`8�>���U�0�'q�Z\{:T��[��MX�,-L�,j����g_�HMii�tTK��k�}�?�/�{�B 3��RҲ��FkM��7�!ۜ\��f�:kV�6����8ĸZ8���_x�׳"ឋ� )x�@��7�$��q���nY����.�L����wo`�x�,�r�:����i7`D�&�L�#�pp@�'Vɗ���9��*�^��Rp����>j�G[��)Yƍ��dI���j�Z�h�\b�/�[{�9�P��������%�����6��p
5��lZ���FѦ?-p ۱�rh/$�cvߘ8�	k���W7 ,��F�9�i�z}�xb�p(�l��C|C�힛����2!	� ]��D�_ב��w��?��p�G>��W��;)F=����+2$��'%���A���O'��
ꏞc	�mO���s��l6��-ߙk�c��P"�q&8��TAJY�(UI�%��������a�*�|۴���ݚK�hώh�*�|q�Vur�okp��I��k�݄|���ĖO0B��au?�v_lZ1��x�d&�>�.���zkC��lڛH8u艧��"�\���Ã���*�e�Z�� J�(���E,&��N�\e��d�<�iՕ)f�bĎ�.�ͪi"ݢ6)Y?����#-A7�]�`L]��a�s3]�.
\(�]a^�hd�VZW#��Hf1$=����T���-�'�E~aup�7�j��W�;xS�����%;o��x�
�I��>��x�hf�{��@P�8���7.��=�J�+ܹ��kL�Cyo��Q׃l�57��vX���Ѳ�߁%t�ld41�@��׃�-B��6��
���T���Vȶt\�Q�����4P$�Z.�����F��>(g|��4�I��g�$���JS��L�
��%���c\lo6��&<PV\5H�����J��+��C�!S�7�d�lԖ�2=�PW��k��C5v-�xm��%LY/Ǭg�ÿ��*Jד��Uo9����%����u5Jޓ�,�c��}��/���Y��}��~��E"��d��u���إh]�}Ԍ��#��j��L�c�e��Ϩ�h�{G��M�^�����6�IT+ɋ�V�a�ɮN�����O_W��k�i4��M�z���%��J;��DDt��������[�#v���ʽv��ze(r� �)~��[�1�m_�]���:cG�vI�fa�<�'�,�( 6k;��ȣ��=�J�7|��ߢ+�[�����J��}ï�x�]KJ�x�nIsk~~W/��޶!�]��P�60$ځ`{���}w���"�zr}��f��>���~
xlM4�֓�F��������W��Q�x	����-%=�\o??���>��4(�*�+�d^�j~@�*���;�O��H6�%6�%�}.�$B���\��#�t˪�07��Nc����G�:�>H��>�R�W�2�+�ɶY�o�^~�`"
�iLU����!�`S^a�W+9���Z��4�<=��\sy��{������]�کX��v�\~@@'�e�̀�� �j���`LYJ-o����
��2���c>Dr�L��Z�!b�����i�υ�n6�N��"L�����Z&-#RuR��{1�Y[=�!z�Jk��D���u( �\2�2Y����H��|s㈼"Wӂhvw�����o��Ǩ��~��΅ iBy3��a��qiRF�i&AJ)Z6UqT��ks�v��6�t�R���f��l��r_=�L��5���ԓ���ÕL�b�;�T<p�ӯ«7��oAC�6���pM\a�Y�\�Nj��m�P��<�z{T��4�+��ӵ��>M�\}�?;�~�
����?/ڲ (c���CK"WDO��ݵZ��g�����N������Q�dl��I"����Ox�L$�ũyل��'�-��jI���1�f8�:0�/���75�j侉D���������W��Y�Ù"/M%��f���)��W`3H�X��N$�ϣ��V��P_}z%���Π��G,ر���&�N2���+v"$�W��@Ow�!��a�7�j����������`���y>��aj`�<�1.��{X�r
�9$�*�`A=ebm�1�ef��BWZcy�4��<�1�[��_>��N���I���D�e����L����b6��)�̵E�&Uo��������'�7BY5*��R)tw�H�PԘz�ȸV�MP	b�ma�"&2֧�"�l1� ��++��-B#@<	��d�!�$&I�C�?�g���
�3Hu�8�>sZ.�t��#������ʲ� B^V�D��WN���
8�������/����:�0��$yx�a��H۾�{��u]
��1T?�*�0Y]�Љ�9�$�4�M�\��7#�t�MI��(cf����,�'�[h�rs�j'����%�}�*��lJ��k2b&��hyQ�'e�jD��(v�]+[Ľ8��SS�������
�7��(���1�9J3RE.���tc׏OX��G��< �$������ϟ����T*�Yn8�n�*4#;|��2��`���I+z�yD�x���Y*3h�X0�}�0�9E�>-��(NN�T�П����L�x������|��XM��;���Z�N�=��0�Rc��ZE�λx��4�uݯ�=)����!�v�z�N��������A��:�����Gd�B�I����'﫡�1�nS,���V���P=�Y��[F��2���}��|äozV6N��4�7�41�t�
�����EV~G��ѡDX����6o����YYJ�F�1��_�Q��_B�J�}�	��lBh�'$���&'*w��|#]ǌM*侵Q�� _f��j�T����1�b Fw�8�1<��bVŨ��}�r�Ҩ�{<�������iGGԻ'��dq�D�#����r�p*�)7޹N3�]Zi%/�\4� e���fR�}ݬ��˧X��5�Ʌ�f�4z�a�	?�פ�7���P(C�
���M�׺k�ޫk���� ЏGDF��%�/�� �^��"T<|8(U�c�Ir'���D�;�D1_�����7���)bi���i|�r�v�j"�b��U֖�iGcMa�`q���7�����"�@���+����r�+Fn��g�M���'�x'�p`�!���;���{������,�;u�GLD�����L�?fѹ�\�%Q�FƟ��<���H�E���Al\@�=ݪ3>G�x��;�9wq�l?�C~�%/�6�UK���/��q��^{�t�?�)F����&/���>9�8�A|ld��]����e�D���xN�#��ę%�����T��������H3g�D��f�w��%-��1a�"x�JhA]S��%�o��2�q�KL��Q�i��I���*�=�)��鋇a�ťN�� �++�����0OIL��T��Ypo`4���L&�ذ�޴�@~�(���I�q�j�<SlH�e��P}�?��ZBt"$Ȣ�T�Sxf�޹��Z�]k���[t��SG���<~�G���ܰb�(�6z�(��Tn\�{3�~��E��'����r�	U�R?�{�'#c{� ,�u0Rǎ��s� �B�G�����*����ˤ�ȥ���	d)
����Ѵ�o+M"�h4m�%�-Lpu�O�uI�a�^�sԪ���]y	�v��4יc@�친�-[)�v�Л/��U.X��'�^���ݚ���~>꺃��jzЄ�Һ��9�8�䕚h$|���sP�����i|%FM�w��?&�ɳQ���!W�;���/��B7j#B�jl{P_zW��@Ê��&V��ꏴ;a�!z����n�
U���/�9�i�l��ɵ9���<R9W���W�J>P������wr��E���:P��5j�^8b���[C�
���I�wJ0v|�����bahP�X�G�v:�Ӱ?/Z#��3��ezDJ�m!!��N�[]�Y��Y5��*�(�h@r� ��S5[�Y0��OP�@��"���\]���D@��o@fd3�U*���42F)=�G3��s��f�)NqR�M�ݖ����E��H������<�Q
����j2V�nɱ�g8�`��d��pdL���e��v�����*��ь�3�p�E���J�5Z�A�-B���H�Y��`��7��v�_Bی��a?�Y�9^��=���A��\]� �]w�Q�|�UL͋X�z8d�(�JWb>��@C�@'�{�Z�����8.��G����{�zRr|&!����(S��¥?ۡZn�J�<4��-���M ��}�c�*������(\'̬(0L�P��J5�m5P�W��7װ.v;ۏ����%�����07���:(���;�mRrG�i���	� �v�> 7f��̦�oJ�eH��D~��/��"�_%l��!��� �L�A���p%aT�]�|=U��?l��zL����Ф���tk�(:ы+��o/:Oh�'�"�:r`��lB3�f=�/	��A�D��J��֐�<k�2{�)��	�d���~�����Q!�1�S.x$�i"Ǩ������w {e��%1��ha�g�l\�k�``Y��G�?�kݡ��.fo��Ӵl*5X#%9�2_y�	�{�5 ͊��:���$�QM�h3�[=�M~�u��^�ؕ��[��r����>݁ܫ������v�&��9K��_�r�Ao���}���_����'<�J^��.O|��LG�Du�f�S�r@��c���yߵ���*���#n������.?+��=�o���E3y3<�-6���hj�ր�M�y���!����v|�5�'��t�ƗhA,��N���xԕ�+"*Q�	&�Uǐ���B�8D�\��P��ZK��Jɰ�z����S���0؅�38�sd�6�:7J����-������x�9v�\���G|���s`[���c�HrL'�����^�K�,�y�������[
��!�|;���+���HJ���.W�z�b�*h](�2q�q�\9-��Ts�6��[w��=��C�kY�t�B����x�8�[)�CH0��,�q,`U&��\����'�Gǒ@��Y��ɩ����-jCUT¸l���}�q� nPˑ��3)R����C�R:5������D7���И�&t�xF�oP8��g����jA��*�|i��I�K�t�b��?��ٌ� ��v�}g����=)��b�����u^���}7o�w�_���vMWlʕ!�/�6ȯ�	�(�MJ���
������ǵQ�7?"��������@�2<����l�O9��ӿ�{ܮ �W���%/�C��o駿eS4`6 ��t���qPL`��ZE�"��,�]�k�j���Od��>i^h�C����`,�^z�K>`IC���4����\2/Oom�ѽ�B!��5�l��k8��t|��l�sf�J��_g� �D$+���3����}�W�s��Rǧh/��j��Eޒ,��<���·oƞ
�g(x��?�Y�$�V@��m�xQB{�m.�����~�yb]4=K'�J�}>���׋�:��HF��k��	�%�r�+xm7Ȭ-<��`w«m��ta�=O���YQ\��]��B;�����'ĵ}S0ٌd�Q�1v@n�V/���O����.�,�oz&_J�;�]f�w~d�ƞSZx�T.�&��k[w����U�m�$�
�q��,�v��-+p�S�QV�v�#���VRR� y�
ǎi��|��L�9�@���u�_�H��6�1��8�{�� ����6zd�Rn�]-9�ޤ<���#)����T�+W��E�Jj� TY�A�V�'W&�o{���lA�����L��3/�/�q0"@������eӒC0-匌�ɼ�_7��Y�2�M�#���p���X}�p�M�TAd.�=�f'9��lg۷G����0�i������ޚ��v�ׂK�Ǣ��:��{�ǹ [B��)5t����i�6%t�5����52� �vQp2��q<0{�M�A�S�Z3������7�ț`+r���"��&$�P��|~*vSiy�o��|	�Vj�s;Y���Y��*%$��=�]�ĸ�VDO�~ �W-R?��фe�����h�V�P�FAŰgV2y����n��U��w���ڒa�ڰ�(�]*u�J#�z|0mاˠX�yE���e`�k䆬Mw5.�d׻�q4���Z��bA��_U��@ ���:p�d��<��'C�rD��!��Α=_Nw�+�U����	Go��E�����߯+*@��� ���vubh��?_�;�^� �=��A[b<�j}&E;	LWJ���rh#�|�w\���Po�<I7��s6��`�"�C��ǯm��Jg��y��1{V��P��+P\�����#��� N��тU�����)nn$
/'D�A{�g�o�(e]�(u5�����W1�����DJ�.�yg�=�yxc�'���U����7�����X>8�L�����=Y��r�'���>�ߐ�]?A����]#�#�Yᢌ��� �S��6�B��tD��TQ�OxaI�-Io:�-B�h+��h���t����d��򾣕<y(	�~��˻�-�,1o�!��K!�D��$,����%�=KQ�|#��"��f^,�i{{��f�!X�,����q P����	9�u6�_�Z	]U���mS4��������:�|yٯ��Eq��s�s1����Iܾ5r��t�����z�Xtes*8}�_Y�����(y��Bn�3��� �͹��Nl~�~�M2�UE0����OH�{��6J�MA�Sa:���U�gEC6F|?��_F����I�?!�@ao�I�_*�R	�ΖD�O!�xw�K�⭒�儙�a�����q�'����؇�v|�|n�+HAoXڻ|O��aRq�� w�8�����vDP��(�I�/\�؂�Մ�nJ'�922ׄ��/�e��w{~�^��I����le������vե�ra_+�!P�g������
g?S�Z�8���g1�)jrb[���fJ	��$x_k��6���V9�u�Z3BtM��M� ̵�G�qT�JA�D��址#����E�(|��~�Qtob�0�	�	�����^ujz;��Bq]-�J�Ze���6ZY�]�Z>YT��u�e���1�ʙ���Y���DUϑt=�^�8V
��\�w^T�
jZ��.9}�x;o�0[y3��*�a2[2@=	k��G$v�liH�h@'Bp��vZ�?�.����)��a��}� �Ph��n"U;���@b�H`�)�E)�31`�&3���3�.N(dw�FA�͞'�������쾏��sI�7�(��W�:��̔��65�3�Q`�>I]���.�:I07r��[�d�/��$����z�2�C��#Y���;��
�2���}c�õh��V��Zaѱ�����w,�Q֭��=�zN����&tp��PS�*ʞy���42>�x�ѵݾқ����k:��0`��A���'~�j�����zg,9�=URc�
��7c,/�Sj��|���
���ű)F�\v���E�	��E�,+T/ȷ/��Qb�Y�9�d��+�=_�c�Z��ۨ�Y���y�d�uj0��	-m�N�fq;�ҭ��8 �]D��� I�-1���7#ˡ�*>Z��ta$L#�x�_ʡ�j�g��j�!��s 9������K�Ԟ��Xv�vB��౞'Z}a�N�*����
������*�
���}���L�O���IB�x�u?>��Go�h(�5U���`��t��=�hAx;�1,x���MpC�?��QBtM���#0C%C��&��#P��{��"�]�3���C�P���3���EP!�D�b��̖��i���ͧY�U
k
J���]�59��gZ-���K3��t:7nkSPa����E�,���0DH-d�.�E82' �)�(;u�fJ�
p����X�a{�ʒ�@+�ě��WZ��@���!=�+־��ȍ~��X,���:����ؚkTH� j��.Y�U�C�ö��)�N�v a���ʿ�l�ڔI7�,+�n���b�vš���<���9;��@6<�|}.ۮJ3�a��au?u�a��:��:�t�6�Ka�'ԽW�n$m��[��a�� )����l,�����AW5'3���y<$4%�;aDS��Ȧ%>\{��ʥ����k��陊�Ҭ!T��I]�y�U����ʀ2�MA�{�~2�{�y �ы,�������"�(� �y���eDW8�xഃ�����p@�B�@eK���E�ZWSC���̼x�F��8h�����Xt">���v�)s��W�ͩ���s�Z�D]�f��{��� �2�N�����4��V�����$%�JDsn/�H?�#}.\(�g�:�IK�G�/d�(X3���Z����U%:��u�[��`r�`�4��PFs��ܐ˗b��.���̽%x���9�Ş.ï��(��K&x�u���{8������_�� l,��Gr �:��[�g�6�Ե�&��ةX��D���b�ӨKdO\���r��k���J+�kp��]�-�ZU���:���9��B�R�@dZӆ�m�\O��K��4���ldf�̜�Պ��p�|���vA��iDD0d.�w��H�Bƶ]��������	/2��fD���,K��w���3�M=�:s��mx�%^b�üO�k'a��t���Z^� xy���.�l��)��ʍ�*���:��O��N�[�P��SRvbw]@�>x���RT�����˕4Ю<U��	M�?���?e�R��T#_e�c,��50���wLaWoTn�Nj�;C��7!Z&!�;@�SX����4$�(L ���MF���;��
w���^M,���*��4�}Z�����M�V�n�y�2����\sU��V��-4\<_f�nM�p��4���T7��Es���h�d�BUN�KWI��L������.� ��5��^+s�%�$b��Ӕ�z<;;�+��9��p���� �1��4�� ��U%�3�T��jn�y����݆��MZꜭ�hI�`�/� =R݁���*�8���n,������"*�FȤ��;�Y�߸s�4��bs�R	��~e^�e�5�M����:b���Y02v��C�`K(�7�%������ W�3��_%����z2z��b�
n9��� �2 ��6-��l�f�;Lz ���/�1�8uwIӅdg'��_Y�B1Q�6�m�c��+q֢�m��_ Q/��5�f�6
��<���!Pפ���)	�Ĥ��G�-��el�?��7v2yE����]��Q�^�p����[���4<�K�E�ݥ	�-wj����:
�@\��X�%Y��if�^(m^�:(��4��#���ݽ�
��?�|~�j'>�a�$�we�Ⅽw(�d���M�E��u1h�UB4�D��5�X�0�}0,�"������� -,Z��y���\�C���<��L�|�d7��i�R�Vn�6-�,�T�>�*����9x$P�X�S(��e�~.�;+@�,A@/���	d�8�f�'��9bث�Dʙ�c$vK�d�Afh+�v��z�2��Y�If)�.lQ�8�[��qR"�R�.�
m���m��rᭃ�cc�*U���1o#v�5�꺾�;S��&��r�0�#O��DM����ڙ1�d8�
t���Yz�����십K-(��#"�5��в0d?j,P�8�E��}���^�E z��$��O���}-OQ4yw�:��\e#T�ޒ/2"z_aZ�Lsk�J��F��I60��sdi&I�����������AY>Lɲa4�d"\z���îS���1�gZ�'��7����ƣ)ΜsJH"xR'Ǡ����1�����{��r��E�a�a.?�Mݽ��e��W�7@�^h#�=q�cr�BF	�:���Bu@Xmv�Ù*fؓ����L].�;XU.6e��1��j�r~( %z�XAAg%�1�q���h<�:�t7rIFX�2�=��\�j�BBG������0o$h�����2o��k@�2�z�D}�U�*f��5q����XM�~ېCb�\Ks��8��t޷T��� D^�E���I#�Y��L�a�13�y�����;o�dI(����`���TQo0�������p1������X�\O�@vD-k2^�*���,�����ٔ����9Q�BFZ�b
J0���sc;qm��B��wSOO��w��oldټ_Q~�F�ab�kc��9�s�R2����}Φea,�#���I}�|`!��U�0�w��^ ��Q�Kٽ��OEIf.�o#�.@-~?����q���T�4�a�(Z欮��In��D2����l�s�C|:����^���C��]�'b�YV��rx?(w��>/���Q���+Rrߐ�X�r�1�~O��\k[�*a\�T�p�M#*��wh�=�c�D�&)�L����k3����-�L?��n�c�9�"`#.�Z���W��*���]|+>��;X�:�'܈V���+�m��b3e��\2��9v���_����TB���t��(�x\�]�A�Pl2߼6����Wy8��G?�r-c����r��)�t��^#�jD��Z�c���^G���zC��I�Rxbd�������so�FZ�2��J3Sӄ��<�I��Yv�9�̫� �����jG�s�;�3�����~��Ws�*��"�ْ "h�_�M��0|{����g��v�/ހ�t����.V{�SɅ奶�{gxl��^���q̉S�w:�2�#pN�wU��p�zM	,"u�\n�|�"��e1��f��A|�_�@���C��5Yx,�h�"fc#�A�xL:J{D�0�aNg�����_Z�E0U���kTV`]�+���wI�0a�}����,�`�N�rɳ��W��j���N�]W�ؖ�ۖ��|��|��,�B�Hr�<�����v�|�<|�hpф�7�N(�����I�⃛�,T({gS��aJ_Ft,Cm�Z®E�mD�W�v��r�( @�Ы�JTm�
y����=����+��j:�@gW8u��n���ү��J��T�� ��i)W[R�߱���$,Tu9��>|�V�zR��=�
p� ����	�[�R���l��d�g��N'T�.��d�a���>٢&�#߶4�G}x��#�����'X����n�M(��p��,�qf�7���N�h�v�� �8�|/"�"���ez�w-��<��[�4�,��O#���g.i6�j�|�B��	���n)�yd;�biEJ�F�{7���_`�B3��w0n��&�X�s��,���T�^I),�U+*ӂ�_Z�R+������v�������c��s*��r���%BrJg��v[<6M �m�fg��X�����ۭ��N�-��B���|ve+�
Ž%�J���.{N0'}��2�T�a=����b��S�~�]����z�R���=�hT}���qc��|�]��X�F���л��'?���7���d�΁�p�/����;�t�^4���5��
���s3/z^��2��qC��'����5�u^X��E2�Z���T�"D24.�,����r,}�0 :ŕ��^��ӟɸq���췹����m�:���'�3��=��C^z�Zw�%oh���:�գ�0G,��]�e�)�5���HQ=��/�����8$�-�lzA�p�7��rp�x�LH4F��?�	YΠԀ��&Mr-���������>q�����n`c��)]"yk�@D���95��a'H]J��@��V�O�\<OїL-��7�:R:��Lz$��Y��k�Y�P�T��o��.j#�.�ן �����UM���r�3$����tr��R��r�ܘ�u��ཷ7�lO~��?�P\�m�(�]��e$�������PެsO�~��!�(H���Q	�M,/[P+ެ�[:-�R�X�`�|�`ҋ��Bg�'j�B\�����k`v�7bخ��;��Y�e[3E�l��i�EѾ��5���t۾�%�h.cr�xPW�E��;�eT5�C\�d�t�	�Х蹗�� ��'e'�[d���!Ο7�1Q郢����IT��_�q(��d�J�M$�H5h]2����(���QA����Ѳb�"�c��{�J��R+����Agg"`2�v|�fG����_�W0��j��9��.n�˜2�2*z�GF��d�E�)m�I<���.�U�� [~���+xz;IN���fHH*4���c���[vӥ0?���g��'���Cpk����"s�y�!ݯu"=���+���p)�LyO�u0D	���*B[vR%b�*Y/�jR3�ʽ�'�v���ZC9��
r��]͔l0�z*A��n��sГ(S��εx�1��q�}.��J�-k���.�PW���>��"m��S�I'}��uzo�w�w������K�D�fa�/��8���n����[��������īg>0�̑�ńc�Y�r
e���jl�A��1��[JH͎�`�
�Mv6C�(~�U��S��������� i��K�c~U��.h��r�� ��q��*l=p���Mb	���I�� �/b��j)��}�
��g@� �71��)�X����n�'�{Ń��hzgp��T��^���X{����-��N1��@R�l	;�������*��,G�g�(ϧ�X�kQ�&��2���u��,l���Y���,������k	�cQ
���Nc�G�2�bQ��m���@x��w�C
�}ۖЍ�3��I�P4�~w��IZ�]{�3kro��q7P�Zxh�#Y%�\V[�0��f��g�
i������ȉǪ21��=�ylw��Z���X����y�n��NՅ`�O��>���0tm����b!o�C��
M[��7�>�K�=���>xJ���U2%���T�0��Ԇ���n��*L�ӓ�x�.D`��74>^���Z}�@.�@��F��y��+�D{
4	�Y3r`�}N�E2���qe���(`�ə�Hb�X_k@T%Vp���4�G �Q-"lr<j:�tŌ;Pz
 �b����X�t�ę�w��"&"�ʙl¹ޕȱx�m�Rx�؃JK���&��cI��v%��yɯ7( �mW�M*�Gn�R���N0� �s>�ELQ���j�FTH�ҕ�Ƥ"G�I��i�C���gq��7D���Qz\�����й��LS!��>�#'����'��\;���w�k�n1,���
iLM��m��Tq��e.��s�/0��ѝ�ZR�˖s�3̣KQq������2���|�Fw�zd-�
˶w�L���W�X#�t�yo��4�-���
�G0I��Bޗ#��^4(�7�uQ����]����+
@/���ڸ}����к��С�a�[�5"�t
y�����A����sr�m�<�6v��~�4蹳��ER��� �Y�mm���R<FO������^w���>8��\�}��GZ�Td%cΝ(��l����7�u���:��c���	��au2�`�b)( �n��� ��;X��sT�m,CΙ3m��6��*��}F�#����₴Fق���Dd��T�[�'�����a�I�3��7l/$(�j��Z3�&�N�9����z�V���"��.ʼ�O7��/� ��ښ�\�|N�2�P+��*�����o�*���X�"���fn��sTa��ۤ.�(p8�?���@!F�\~������ǻ+��_ʴ�����UW�I���(Ѝ+W���F`'-�c�1��m��:��$���+��[ݑp Z��od'kd?#�ly^�_�[�
U���Ђ?c����j�s{�}�	}Ko~�C<Wh���������Co�M�"�0Y2�C��0W���H��.#�����em��5d���$
N���tL��Ds�S�ΐ|Wz	Ar�p`=�����̉/�O�5�nt�����X��f]k��H,3ń���6�"ŘH���9_� �E��J�v�Wj2�}���ev�Z�T�șM:4~GA�����zY��1�`����h�׆+�"�w����$o&��jL'�F9�(��|O��_E�s����,��F��	S'[c��ڗ�5+�|���hKF�V^��Xd���<�Y����P�F�����Q��9v��1�4MÃz��ʽ�1�#C&�1n083ѹ�1�'N ������1���hŖ{�5t����o
{P\���^�Z	
��Ҙ����&�:�����ÀC��q������k�c��(������鞻�a���:�������8��u���:�N>��>�-���9d�3<��Z��q����6��x%S�,O>�dW_��=�_��7�i��ʛ� /Vi%���ȿ]�⠀F�a2�2���`�B8�>0���>Y�/�O	�=�������W��z�Ѽj�DD�36p#~F���XV᩠�����O�"X5<m�Ff���F^�*�|}iSV��6��|�������~����T��Y 	�G�����tXku��p�X���A7,�Їa5���q$�:8�[����aH�SF�]���o�k<>@��ʝ�/54Y�O�ym��ZG���)n��O!uu0�%C��|;�û��fi�b�J�g��9��8�	�C�߂��t�6�=@��Է�z��"5+#q�ς�MaA_bx�*��J������c����5 5pǷ���jm�7�W����Y��R�ckm�9�י��z��Q��O�#��(�?��W�����ЫE�i��Hȟ��6��B�+����ga��O����^�h鵚ZUY%�TU����*+�|��B�!R��Y#K*�o��k�l<۲��'�4�G���%�6뗐����Le ���P�r�q ��)7��Y ���Sa�n�z�	4�̍��6$�=4�j�pɛ�@R=v)��g�c�D��샳�u�>$��w��T�𹏐Ҝ�h�u���e�w������1�v|D�����S�#���H7�K�mP@���se,���
��Aӭ�W!���
��E���0��d�]��1��S��ʳv.Q7��4��5�Z��� /�(ܖ?=��������!s���oCo��1�U�]�lLq��`���P�9�+sX����0,�rM`C�$O��:7�*6a������3"��k�����,�D�%��EAt;�+�C�tv�Q)x7��� �YO��z* <:�+���.���?+ɵ;�KË��� #�\�|�FfV�X`M7��,�^�M~�Lo���5G�9�r�R(���RXd�MD��zi3H k?�l���ۗ�Y�{���y|�W�-C#�����B"ĖH[�Z����h��=<�� �H����t�/X�KǄ&���X�1��"�^#��:��Z�t���b��G} y�N	����7s+�$���8��}�e�n��Ehr�,�(su'g�s�TX$�'���3��Sx�L��s�'�f\<�8�MU0�s>XҊd��p����z���KK� ��_jR.���މ����=�L�g��_�!��D����1���8�%��J�+[4E�LU��[.�s� ������q�rMH�|��"�Δ�ϦB����St�n�_�KL|׫��=uj+V&����y�q���J��75���F�߈B��
F������������W�#pk"��O,��m���1��>���1�l�H!����O�U������qko�V�g�2 �a�oCb��D�bMi�X�E�++gW8V�{ы_��s�:J�oH��BZ+n� �8��ԩ�����R��m�[ȩ������/�該/d�Vjq?|����-�|}m���d�"ZA�U�?���>�����x�|�΃rM���M�*�ǌ�?MFMu��(]C?�NxP���j����̈́��}��p�{���V�\Z��u����H��ڡ�f�������it�~�8���ᗦ����Q�ZA�"{��1qk ���˄�iI=��3M�)(�~�N
�/q4LM��D��:����� ]\pnW���~��9�!~��x޲��T�'d���n���xo��G6x�	����
qJ<а\U䨁�v�ʉ�ZD��T����i�O#f��R'�P��������w�h�����%0T�{��G=�ߐ�낅s�ZS�!���k�3�Ur?�v��=�D�9��-�n����~���NSZ��RqKy?�ɮ���#��5�<��?�������k9�u���Ҝٳ��g^�F�|����,`����׃�g�z|�{�,痄;�`��!�u��Inh�X!�c������56O�׭!���}���=m��<
RR��Ä����;h����rF�΁=����:��!9lrȰ�V�v���O<k1ct!h����}�T�y�Pb
6ʂ�7�����Ȼڡ�W�輴��v� S]��a޶`q߿�<s��1VџOj�C�x.]�z ��/���EAȮ}��K������Tz��"��)�#0&��^��1���L���k"� �*:7^���K�_�ݔ�?�"���5c����5�Ɍ_0T;��槯&븨�dh�6��[\�~Ѱ��)1�)}�4�3-[�Ͱ�}c=�ڱ0�pHo��I� �m��[]�����#S��iˤӿ��z�ާ��y����*�rY1=�{����?�e5�N���S`S<�>k����,�&�0�ʙt��	�3��s��[���},��	H�n<Q�+�l�$d3��f�aa��]�A�vK��r4�1�X1E1[��7����}��$*�0(�Fx���}�θ\�\4�\Y�Sг�o�?l�'r���n����;���TU��c�2K��#u?o |e������J�v���,���v �&M�X�ƞ~5U g���:�чd�[�����	���b�| �b5*�s���@�����r�:���\D�g>$Xq
PhN�>(}�P��<P��^1t�d�G��KEF̈��T��s���3^O��&��{"���k�����?8��7����ѵ��Z|�j��"��xN�_H�U[AC����~�p�uE�~���5Ge��T3K�"�J���h��X��&I��<�Q{�uD}O0$�u^���o����2>�ZZ^�t4n�΁��4��V��PT��Nϱ���ǁ� ��:��¶A�v��6��Fΰ%��h�l�6��P�"C��f�wU�V�ݮHe�
�$j�����Ȏ[�q��kY��,��i��_L(,�]Iḡ�u��#���a(��I�p��逆/O6����u�\�E��Ko�M�!�Sn�!		͡w�ؾ]Ј�>���p�g��?xYN�©���H��#W�*�5[���k>i�������BB�+ZHn����5)8Y:�E-�E�kc������3՜��>�S(���s���W��=!~r٨�k���UOV��Z�f�=8����sB��Fl�!dE9��.��`f15���"�[
!k��GZc���KCWXr�$����TA����v]�
A�A� �
�q)��3D���# ���7M���KY�;���s];�\H;V»4	�����y�3�_^�����;6o�. Y]����:��Y��Ϫ��B�/�*f`A/N/_H��ٰa����,.���.s������}ܯ<�y��m!�e�?:���i��6��o�ߙa�o���sn���X啷(���>�H-%o��$���k�5#�{~��������V�v}w�@�j��vQP�F�J�a�MiS��記� -��}����������)��F;�c�X�i�`���5H��Vl�5���0uq���id�[�������fr���=C�Rv
�ir\�b����:�Fyۡ���g����m̢�i��9�WJ�8�M��ݢ��8�m(f�8�/g_fo�z�������Tey�W��(�
̂`d���X�QƱ�eN�.��I{����3��6$�1f0�v�=�z����nVێ� i���(a���m���Tǆ���n����$��l�_A���2����-/Q��3�y{��;D�~�&e�.h���
1��� 6I �Uym�T��"$���	��N2��bf�z�r:�}V��R�E��z@���o���kO�2�~DNx�A�.��wL_�p���9cj�:�ȊQx�J��I��oI'�}��n�Tdڈs��)���М�n�����w�O+/�����P�<װ]�xm��$暴��Y���n�_/�6ᕕ�Q��0�Y�u��1Ҳ�
��p�a����ڎ~�N�++�B˅�~��gk�D]u�߿�Χ!d~��ŷ|et�&�ȑ����i���|_�;
XK�XlEm#�A�ߩ����iԩ�!_��a��??��T)�%��hr^�D�1���������kbL��y��K�|�y�lTw\��B����՛4�q �G+x��ѳ��5�:�ި;T�Nc�͑'f9��U�)bsZ;e������ �>t�T�N�Y��.@29#��eeQ���e��"���tR���L�/��{Er��5���b{����?�,uEy��
�A0�pd�y���YC"����G�o;�(���(��t'�ޤEVGr��&
U�VU�e1������G��<�<�i���,�MG}�[3$�x�'ǆk_�0������\z������K�
G���H�����:�VK'�0�?�KoTµA�Q�<��X*|�\"81X�<��	0�>v2<���(v��wQ���)h���O�UG=9�RH�����\�:��_Nr�m2�qZ0�17J�bAt ��4��ZAA]���g�~���+Y-7#r�7ÖT���s�W�ץ�O����z�.by�nj�M��6�(3�]�H�M�v�`{����>��5�����*+�W������t�J��U�1�4��D8~_0�W��>�8ឪ�֯�,�;e�Fu�ᘺ��3�c<�oH)6�2�YGȓaogw��m٦�\Fڜ ��0�N>����c�EN6�f�#л���g8���*��VXJ2��p��Y�Ʒt�81.�ks�8�N^��m��e�ܓ}�����.���F����� �a���U����=k{k���8J!����gX&h)9g �U'���c���R �jMjWE������{4C��7pv,�8�ic4c�|�K#��` Q[��fz�PWvlk��Ci*��I���a#�T��Vi	���VjKx��WW�y�;���.[��$J�G�*��[x6)^�*{���X������'ѯr�����!9�fz�r��-�+ԫ�O���|�_��J��V7{;����E���f ��L�ץ�l֗rF^��<59b�,qU$����5�6GAWƘU.�g��Y1��l6f+��V�Q37�������1�vGS��!v��h\#��_s��/b+$.��|�Y�����3���fR�v��ǿM�%�KS_���9��~���S�;�4�k�m4y�d�	sx�Yl�"���ޓ��y/7�W���g��L�è�YH}���ޡSD�#6p§�aC>�ȭ%5��SїE���	:���;7�g�W�6�:��j���~[��=��p-'g�F�d.@�u��q�L� �.ߗK�!f!��ď�P�50�:�P������n�J�!<�ꕯF�+xQ�N�)�1�Q�A-d���,[4�����"EX�R�Gn>�,�μ�>���U_t�pAۥk��F�����iP�=\+��%EJxxP1��c�̏"�F�;:��h7i.�NEL�h#����)v��+���K��s�j�p|o�X}�e\��u��f*@�. $�HI�>���@��,���I�!,��0@���ajju�s�(��qel�����z)Qƈ����� &�2���}'0���	~�J]�շdl��P�����ؾ�U9�?��s��ǳ���ߎz�7O��Z�c�����*����Zۓ�KD����`��#�\y�D�0��;��\K�H�P�R4Zg��}�h��C�1���;.��	bu�Nyrbdi�����{haƓ��k"��hڜ�3]�����g��!���[Lx�/��%�����R��E�`Q���U��'��cЀ	��-ǂj��b`43ɴ����1*�(r
�&e��y�h��c����}��HxC.���hjJ�/�U�w\���^�Af��(o4�{�M?+�gf�g�\A|V�xl�\mnҌ�AʭҶ���M��})��^�iG���y��:���<%�=�z@����.c�i���'�v��@���T4F{vغ��C����9O�V��>+��k#�/�j-���a�eF��rC�����B�p٪ԯ�(�&ޙ����&�:Pf���o�^�F]snHi`
s>&�AWj�IW:yeB��%=;�ԫ������y�UJz~I�L�#�m��4*	�3�&>M�h�eI������I'D���%mA��S-���F������v��*�,-Dj��4��t�,H��~.��p�������jY���j��b|Ȉ=}c�t䪉�\�j�f��d��tN�����P$��vNʡ��x̟��j�akݫ����/�N��U�W	����	��Ri�Z6G�1����&����Tf�7�0��P27�%��V��H�d��E��w[�E[Y[c,���|֋Y;��qx́�o��L�P��y�ٛ� ���ⳈH����G���l��-8C#d_j��z����&�C�B�vW�݉X���m���3\#Z��9D���#��~A�6��]��ԯT�H֨d����aW����Rɪ��n�2�+�2���9��}��%�}Q�Zf����5i��ʒ��"��ӈ�M֜�uvy�jo��$)zRE�s���+�X6�!!�'�(���ᣥ���k1I��Hp������>�w�g��{�U��#������>�MoZ"�z$�>%�
��1�[��Ll�@U�yd��շ s�-�C��.�tC@:W�D�
���iȁ��[a�׍���,��#k�[�.��]�޾eV#Tc�'f�˔?���RY�d�����|�Zt�3�NSG�2�6�L֊ʮ�6�Q26JCǣU����!.�dZI�	Z�,t$;���p`���a^�!��H&#�Lk��p��F:e0v�&V� |��LI�TG<zj�24^Ǭ\�CUF��BJ��X%�B����{83�H`#���'es2{��[IOi��u�ʲ�G�V7�y��b�:ˉh��Jֲ����u������9�
�C���C�y '��N�(�r���8��t<���}�"|k��T��$�sg?����v(��*B>���(ΚZ�R�!�)4BthF��|+�����g��Y���b�'<���
(��=vC�[�ڷt1��?��L�=�v��E&%�z�O�C9��cCQ��7rfE���i�)���M����ewTmم@^Q2�i��H��H�c�W�	���q&9����:�R�]]_��o�~f ѭO�3,=޺�&��^��.^�⋆VZ��˳���*��qeh��?���k~ �b����~��c�h��C�B	�m��s��z���?u��O�q�����!��<�Ԯ����j��D˟m�IH�^�s�M�(���?�C��tl�_�wR�ݙ1O6����"kݕ�:�I��Dz�#��!�U3.�����h���`��1����)��X�sB���ZpE��2�P��-��t�����>W�E6�{��&�U��`��~;��b>��,0�]=fm�:�u}�PvR�f׻�#�q©���4��R�m���s
�!혌I�c�P��z�˓a�� m`�*;��]�v+�E�B<��$bw����<E���������1�
bF�rǴ���߽�ȩ��3�.}�z�����`��r�r�|��i��ܬ���'�b'k�]�!���YϢ蹽yjg���C��f�5a���������}�t��n�΋�D$|��u���fU�c'r^}b��G6a�
q����{�Ԟ0�T	Jn��p.t�O���CrT����>�5tEke�L+��Q3���.��z�ҡmY)�l�I3�-���EEs��m�l1M̻N�?<s���t���On���28z��&�ߴ�1_5�j��D��	��|e��A%�_4=��j�ǫ{���ݰ02�����q���s"O�~����_y"5Bݬ#�����gԥ�@���Tsx�A���6�Q=bSZ��W�P�Á����?�������(� SO��k�2݃G� �Ս��TG�� 7�V�;n�P?U�I��ʕ0�J����ě,�X]�G/%�/-C�%K��M��zu=�f)W���vL�VAY����v,��4U�T�@��T" et�����3S�~���Y-M�?h55_b��DS������3�}��}ӂV�o���q�<
�M̶�{�w9�Î!���d~�n�:	�eD�պmH Ş4�����ϫ�]2�`#39�V��v��LY��]_�dU�)j�+q���$�Dj*�H�d���G���[x�-����Ό{I�'7��n)O[�p�� ����,�uUU׷���I�1�	5��~d�q�R��Y���6Uor�+o�jڝ�#.�$�Ү���ǀ���8�H��<����JZ����O�a���7I�`��|��s���ܷ'��2�+��&f�*��oJ�O)�7�%�c�����ؒMQ�ՐM�V���&��o4�<�u�d�XjD�*>o��8��!�Ku@Z����m��9�ytMQ8��|�l��薘mQi�6hyՌ��g킁	h|c��;0��\c���c���eK�c0��3cR�|�z?��Hf~rHm�������Ed͗�`� G� �n�m�$6�3 `_T��9�s�Ւ%����M�s�̽�,F%$���e:�zPF�sw���m���oM�-�Z�x�X8^_+p@��3����q�[�gP1��!1�ְ��oK��9߾g����eK�IXa�J��h�?7�\]q��vp�ظ�4�C�,��m#�sM��ft�����\������?�p鰂`u�~n��]���.j�j(`R���UxT��!b0�Qt������|�PJqY�k3m�D���޾�zDw��/���T�jv^;�P�������A�IfDTqd!2h����"=�iH�/Q;�Ž�9hV�ץbM��L�q���Y�\�e� 
do���j7=/�q���N����D�"6�̎�$g<��yG�H��9���#�C���) aٲ�/�v���ŕ�-�d�<�4l�ö�1x��{-�`V���N�F�~E�Ř�'(������Qx�R����fT��3Ť;��k��#�b)l��
��]�]P�V~�'1Z+BZ��K=����qq�0����dX}�//�	�p��������sT�(�)fy��r���1i�^{0�\n�SmzE�P��)��Ք'G�! +��[n ��Hok!j�³C{�Kb]�zG$�AjR偟�����mT��=�r*�'�vŪWT1Í���͒u���a��$���.�M	�9Pl�<$2����*F�x�3ASw63w���K/���X�ĩ�Z����v�8#�
�<@k2dX�$�CO�����q-��TV�z��7�](�8/�Iy<޿p��A��X#�>L������<���5�TC�C �4�mnX|>m�6ۍǗ~��1��~�)-1�g&�h;�z�z�5_q?��(����:�����Z��i���D��	p�!�ݒ	�M����$���Kkie�@.��	��b!\I�0����v��W]�1�����!/���Ї��۷#�2�I����_��]˝/n�d,H�6ԡ�ɺ�A��r�D?k�k���д1>��� 7���Y-^ �7�[D1��h|Z�@��Q�J�'����'���Rޝ����׉7�Aܗ��//rI2ȽR� ��SEe������|%=�҆N��H��N<<�L���ŲB���C�A��B���1���,��ւ��!A��Rt�ċ$$w2�=�1W�2�% ����&|�]�������?Q�����L@��Aί�(��F}�� ���9%P+�}�9�K��<+	&�B�5��9�G[������QK��-�-�t@L�A�'�5(�u� �`Z3A ��X�WU+2��,��R�NF�D_��O4��������4h��G�W?��&�E�*M�5j~�ߟ����w�]E���/9W��2���5�==�ի�]��8&�4LA	X�KL�7t	�z�;�R��L C$�6�Rst7�B$�}�oY-/3��3�z�o(3{AN��u�W�5���}�?��\����ak�"�9�7���U"B!sЕ�e�}�?��ל��be*��9q��I��e��Lf54�-9����0!���3�� 	~��O��8�3�I�M�6���,�)ű�w\����ݥ��+���CrQ���t� T��rH>(�4�!h�Mt��pk�j�l�0�������#Ӱ��3>�9a���֨ޠx�(���|���}P޷���:�VF$ߴhR�ɩ��oSUj�D��fJzP%
���'o���/��mm����o�Ӱ�I;g�[���M��_�|]�lbR�O��T�vD��p:t�ܑ�YM�
Z݋��}��ت���cM�xA���"����~^�*n㭖 ��Kk��]Vk є%)!��x��bZ���%�]ߣ��x��lv�D�@�=3C�KD�O���TԓɁ�V�+��:X��(��JaI�ݟ&LS&�zZ�Z�1uFl(6�{>�<�┿��Rj�_�;����:��X'���0p��@��7}2}��VSn'�K�j6�e�b�nVG�o��W�}/$��ws�Ԝl�jrL��A�~8�3P]}�5���ֽ:�~��R��w���g���y	�� ��(1m3��+���*���nF+H���.���%��S�?k����M ʕ��(�C�&��nPt�Z�M�s4z���I����]��V�,��n��)��������x�Í<<���6�0i�����¬th X	Q�Z�Y��5���*�*�O����`�}���
�tR9%\M�R#�QX��@H%�d��T7���n#��b�֋��+dH�r�3֍�%�]G>�A�K����0�/ m�A��X�� V�k��S{o�t�ꛒF����QD,s�� /	o�������&?-�o�fXV
��׈K�X�ܘB	�_7�{���$S*�X�n��; ���x���'
H�xj��{Q�=mr��f��9������O�ge3�\e3.���w�?�I���d�N ��_���'1(g���M�7b��sx�Q�N��oa�$����MK�<�{/0�Z��l|�;.N?O�	ŔF�8��k��ԽrAH9*�1�&�t�2�g�lo:��P�a�=�Z�r����\z/����( P�	�.�D���g�Ab�MgK��'c���;�T!��r{t+���Afu}qo�j��D(F� ����R��z����9��2�?�SG?\�"|�;���Q��0���������o|E���9��+$�f��5[�t�Ԑe���_���s|���^I/�䃵�m;��s�Q������ezJ�,�D�C�'oќ���n��lѹG��S� �Le^i�i��acg����b�dN�݀k�_���M#Zb�_��	S�E�@����c�
t
���"���S��@Hq��p���5�<U�!ы?$��6t�B<����Y^PD�\���Y��ʟ+X��{�T�;>�G����B8���T[�3��cjԁ���m������0����ȸ7r�
vyB�\R���@~�>�NdH@w*�_ �ٱx�P�!�쾜Kޢ��kf���s�XWd&�G^���Ct��k��{���!�x,��	Bb�m�n¶^��������c��v�W�׆�DB0��12' ����q�WV��S�3��>�-�)�����(�Mp�==1�K� ]��� H�X��ǰ��=�g���B[I�Sf���V.K���R�l���nm&i����rN�T	��Hr�}�oV,'�8��~oܻ�����ɚ�����y�%2<����	\�p$J�A5s ��ղS���/ó;gPyQNeI�GZ�O�S�.gi@�wB��:��29fS����Y"�)��gȷ���o�	���!Bz��ܤ�̧K����
]^_}ꩇ���������/�t�$/��[����1�pTNsd����-�*dv�˔m�ޟ�;�<��Uㇿ��1�Q
7����]�Z�� ��ݑZ\�#D��Y��븵��Wm�����j)ʡ�p�Nܑ��ډ+�X�E����(].c"n ��>�# b�Y���`Y�0��h&F+��	@ �}�@�b�]v�Iٓ��(�D���WDf1T-fr��'��?`��d������B�zp�����~ߥE�8�)Y��4� .��6S�=kvzGY7RgW�'���`_^�,���<#(~0�1_��P:J�Z\F>�.n�ڇT�O\�.�hgv�Z���M���-S�,���A 5-a	��Z���w�}0B��=�T��z�,����PBu�/-��M�����H衖:�{^b�x�D�	}F�	��XJ��T��Ɇ�6?��A�~��@��&4ٞ�Ϥ}bڜ��F����;?�8�:�Ait�񞞙;�76�0�L���8��:����?��t�ֱ������,����T?G��Ÿ�9=ģ��Z?k<.�� |ռ+�G����2���E��֭��pl9�`�j�>�����f�h�8�)��k�Ua�t|}Tm���Kֿ<a/M�0�����Y��z�yk�ǛH`_7�����ÁU)�ΰ�/_0�Bl9݃��W.�r�!�)@@��X�I�<zp4!�ѷ�����H� �bH�W�b}B�<_�LJ�EM*����o���K�6Z�g�p�!h�˭��Y	� �����4
����12!�q�ߠ1-�=�������T�%����H��e�mx��D<��q���ھјY�DCQR�Σ�����{��/'O����8�c����#PZ-Dd鬽�fb}KִX�£Ȅ²�񬕲����Y64O�7�	h��8���oR��؅G�Աʊ�AyO�J�3å��^�
]qUv��[�Nj)�'BW�H,�S~oa���"���Á�
'�����߄��7��:^��'w�J�f�ٰ�h ���#8����(
6�'��b�6'@��(6�+����ȹ�`n�T+�� ��U�x�8����?K���呹� R���������5���P9�h>䨍�ۄwn4Y��/BVԙ����|�>�ͭ�^����la!���\��+��ɡ�6�P����f��ș�2�@��¦ciBA��W<3��L���7�pk�inK?�W���`�����a�-����s.*����#��I�q��C���.�SS������@MO��lj��ڡ�_g���=��xB����pu�����8�;|��Tw�C�����:��R|�q����\�M��;��]�a[D6mΫR�B�8��]U�N`@����V�+ǋ,=0�����#G�
X+ʭ��:��2�'�@�	aa�B�d�����!$#wU��"�'E����+t����)o��o��U�27�ӗ)���J��C�0դ~� &f � מ�S��/�L�\�zh҉�,*�Y�F�H�Z����Y*71˯]8�·�a�Lk;�����_���� ����v�-ЃT�^��_i}^fyy9����䭯v�U�Ph���g�'��8	z���{�q��,%�+�@K�7�Q�t�Ô�j�n�0��Vm��f"�Qu��s�d�YN �]y�q@�
.a�嚘�!$a��~r�!Ђ�(��&��WA>sG�噌4 =�)�dV-C�����5o �1H0/^��Cj�&�ږ���'G���Ĺ����ldņ�^O��0�����hC�v�����m2y�~t"�����pO�"����P�5��6�1��<f��)�#��I���E��(�,�ɔox��ͽ���Wp�S���(��rܰM��)p�X����7ݖ�R�NXcnO��{�o�/,��c>��k���n���S��-I<��{l�����R��!�i����7� �"����lFSi^�Y�@����r+��i�D�WÞ�\N�t�?ڠa�@�ч��2���#P:r�/��X0x褕����ٖ�JFZF҆3��#�AL	R������(뜬1Zͪr�����-��*�W#g ,3��:@8��S�}wv��e�^���c��E���-c�z�+��Z���!��*⨏��!�ܑ͋��z�1�X~�k_1�7�Ɯ��{�ְ·u�W8CǶC36�"p�7^�*GjADQ�	�Qf�P���|z�0n̵K����`�?QWUE�
zlS����ro��a�Q�ȥ�A�� T����"���(}kDs�����9DQ֨$�C:R_K��:��s�l�j{v	KT��x"��ˎ9��j�!�#��k~���9�?�˽C�����c��U'�3��l|
3e���d*ǈ��Q����6�*�,Ҧ���oM[�xm�4����tT+�j�Vq�{D?>fC�.}�F=M�Pa;�x�$��̗w/.�b��i�j�N�~8��:�أA��w�W^��7L��Jki�`���I)��5���!k��{�%HB �$G����mwx$��P �!g��G�|@�zJ������혔���M��m�Tف*Ld�=uE�����_24�v��\R�mA�:�K�U���X�pm�C��G��Nc�\ڃ��c��C��9���4Ԍ�p<�����8{3��m�!5+����Z'?b8���|X���eCR-LS�`��z��}v����]uD�LgD�3a�A�v���g�Ov�G˵�~�����)MKky2��Ε�^��A-#�S�6$LT��Ϳ'�d��K��)�5a*�b�J�
���G��Sr��S��^���}����J�,�Eh[f-��97�0K�Ն	ٟv��}�g�pb���O��K�<BL�v�m�X�d#XX�������U��\�\�9+XN��G��9��#-B��~$�-XQ�$D�r)Z֎�dQ�e7��	�n�F*P�P%�B�P/w�8�
��tK��q`�K�Y��K��c�^S�L���V�CS�!�*��]av96���k�ln�f�(+֠A��Qq���������y�D��7]G�{e�c�{�c�/aE�=]��˺g	1������a��r�dFl)�W�"�w�\��HÍ!q��$����	ҧT `'�"?���D�UȷhC��<�
d���]���fՓ<(K�G,~{L���̫�F��}�t3ѥeVJ���:Ȅ�fS"����p��;���=��%�j��A΍x ��{�Sn�P*�d<�y��u7fR�d�$xS��5߉9��5�[�y7�BD^���:$d�tw�����b������;�0���2/Cf,����V��pcAﴱH�
�4��"Ѓ��2�y\�����&K7��������
�&qe��b��<d17�v%=�m�Hn�IזS-���t��4ځ�>�����[X��%�a~Q[M
��eة�y���%�Z܊�� ��tE|��HO�'J���7�Q���,(��G�I3I�=d�%ǋz�u�?kG
��K6#��ǔ��-ȇ�d�|�(?�}���6�]��A�b���"� -��E�l��7t����ܻ����q�i���\r�Oqbdvz��L��[��i�A!����^�X (�s�����6z�Gj�j>h�m�,!ǯq�ٜ�pÁ����;:0�X�c�<3������!�꭪r�_�{��[9oz��j���:A�7I"t���T��z���OO�����5<`O���Ky0%���S¾�=�7�J�ᮨ��ǅ3�EC��T���<ӌ�h��g�0����S4�3+^ggCy��47z���;����uQBr���W����0*��O��zV�4i�9��}��߲:
M��� �F���2ګg��Ώ��ӿa�E���:*�1 ���rZ�{��n$���5U�E8�ɏ��OBª����0��,� h�N>�:���o���K������]�L@�x?�yy�#h)
8�Ń��MoI~��b9�ŧ��h-�%�eE�Cnځ��}�Ŀ�=� �O���I'OnS��<�>2F�n��ǘm�4�������M�눒��x��Y6Lp*�C���t,�u�	�\�[1���Q"<��%��ܻ���QG��xۧ��'�F�0%B��E�yMeB�|ƕ!�H���%��D���!�GA��09	���5�V�ٖI*8�=�b$̑&�s�^��z�7���:��80�+0" @�r��v2�P\U*b�mY�z�||�!�G*�|�9}�!���!?���!���b��_����)z��5�� U&>��қ�ݡ�Ѭ�+��%��ڨ����y���3�)��V���>�W�26�mѺ��]M�IS�Q�X��L��k�]��t� 8��!ft3= B 0��5�?�Kݬ}3�.w0��9�7x�L�h?�9j�^-N@Mi"��zq^�xJQ]枕�3��^��;ۚ�-k����>=��1�"Ӈݨ453�G���uN(���]@���> �N�BT�D��UAc���f�ړ��xMc���	�5!��SA$�t�|�:]083;��BlpGߡG�# Ƭ�P-5(�O�2�1���.4�zI�{x���u�||����Z�9T��Z�g�1�}���G1z�~|�X�=�4�%o�$�i�΂��v�2�Ӽ��q�Qy�vq��Pl!~~٪���?�B_����g��^��3ɠ|�OnF_u7Z���])Kq=�x�?%�`5��2;g�@�k"����bb���Ǵ�Ǧc(e<j$������j��Bf��������,�i��Wj8!���b¬����>yi��ؠ$�d����X,t�')�h]�eh�vбZ��a��gx:餗��m[�k�h�^�t 8���"c�s�z�^].|�!���r#ec}G	���|~a�����y�w[Rb̧���H��!_Y$��f$$�^���3�|d?O }l�����9��íB���O�6\e��1���I�8��PI|�!l��҆�u�]O+��?�jr��py&�&�	�����t�vE�ҫ�+�}.i��bgG��u���&�׸����%^;�74]6�*��d,��,�����[B���Fg���ŭ̡�j��`�N�t{b���]�Tar�⧄�0Q9kF_9xU�蟖�xLm`�:ن���>|����f���\��ꚣS�� 	
���9ll�Au���4�8ƪX����+�����-��k�! �⟖�q����l������6��ZAQ��~dM�w2W�x����Oj�X�~NK��N"Ek���⑜��.@�;C#Y:�(�y ��:���a�2��Ĳ��A��=B$q��l�K��E^�>���KRv܀pS76ߢ�Oչo�ɳ�_Aq���㪨����H	fp�1�?e�k1h�8�)�����9ꆁ;^��~;��f�\/��0����O��QT�X�����'����ы�vЬ��F��c�9�h�O�� �I^��[3#�<%�b����\A:��:)�Aj�!xr�j�N�_C^$��#œX����C��y����g��9Y�5��FeE+�u|�\)�� o��5�zF�Q	�>�
��:�~۱+�('�pM�j��t��q�X���~���tf��.ຂ�Gُ����n�X�۾�
 01�Y,b�E�G��YK(�^�c�A�A/j�:��M�o�����6�L�%�nΉA��˫�\ߦ��4��Ha\�2�jV"z�Ù�'yY���J+x��1��譒ANE<��$ [?z���xG�����Zh��p_U=}P�۰^��W�D8�� ��*���Uzҏz�[3��=8�i��_ѳ{6�0��[��9������~?,�V�}k�H,8�^�]R	 q�JRd�����Fա�B�=���T���3��dli��^I�M��po\y��9	�E�ut�LS� $ ���"0=�_x�?�3�lDa��x*�<e���"T��ǉ���{7�1��JzǑ���ᅳ6p����0A�m�I*�toV��=l3��C�1��ʯo�hub	e�|�
y��}E!O:��X�ڶ�'��IZ�)�pL���a�0�\�t�@�Y�A�[�Ff����T�F��ʠ֝����ݔ�s�&�d؎	'���VN�*g2>�3�6�m���=�)��k&��1�o�#he�"�Q�\��-HYD�F�n��=��'>sp�I��kYRl�q���֢=���zF���ˢbr��X��a�M�}�^����@���o���M�?� �����Jc*S��̥2� ~]���Km<˧�{t�w�#�̳7�w[ ���'��8Sׁ���ݬ;����ك�#�Z3蝷��Q�h������1NS*�+2��F�;�5,<3�%���^��G5;�D.U{*��q�.��e�oN<�[���A<dHgu�jM	$;p$I�ً�M�}h-8J(6$�У��2�v��O��ˋe��&������.X����&zv��Sޢ����'��*m�r��b>� �ջ�?Hܹ�L�����!@�DnC-)�r��krh��L馚-��e�~z�,�V�/(�G�Oޥ�s5�rk� uHf�[6Vr��o.���\Y�;�x��F���
ޙ�qȢj���p
K	��Vǖ9<�K6�LfCn-�e���Ǜ�o[�� �:��۹��>-qQ���0=�2'!�α�_��0 [��}ۥtX�㶁J��E�#z�Ȝ��Nv%� j���C���W�J��mk���Ԍ�\�?�		��t`i}�Ey�4q��Du�0�Z�~��Z��) =L7u�d�d� i�c�
7�/�f�����3����@ŭ���)�����|I�"t<�³�8(��7�n'Hy�
\:-��6�۱A�Y
Y�~r�x�r������fh ����м	�/�V?��oMu��ͬ���A��עn�3��}H	,�?���Z�D���W��e>mb20o���/���@�L{ջ��W�4水iK�(Ws�B���ᜯW��Q\:�� �q�d�?�&9y�`�i5����7$h`/ߍ�tă�|���\lUԼ�6�M�HpV�v2s�Y9�ԕ�Ⰿ3Xd�p%���Ⱦ��	UR�m\?�j�Us�\c�UE��I��%i��׊D�H��F��L]%�kx?+i������~9�%�T�Ѫ�*|Ȳ�.�&C�LC�{4M�i�?��������ѫ�ĩL��r��׀���VO�Y�kuE��䂖�ba�q��^�-%xW�����A�];:��&j���۟N���� ��V̩j�~��'\�V�H�b�襈�E�m������v	�`�wP�֡F0+�Yb/f���E�d��0q�}��M�
D�a���Ty���x������f�Ӡy��SG>U#Y�-$��xV���xZ���U��yq�&��/fs���>��r��}I҈�ݟ�e/�l�R����'c�\���䁭�����H^/��t���1���.�~�J���w��{�V4����FM����>�Q���
I��^��z6�3�S&K��]�1�^�is�kv�����I�zbXN�wB�Z����v�D}��+��B�s�w�x ��_�\1�x����g$0��}qq_4N&�H�_exw�����q�7��uE��g�׸�-������m2AӘ��u곌�ĉY�H͵�)��m���ą��=Ӭ'o&օV޸bO�9E�p_�8)�}"ɮ�թ�T7��K�6�4�T��S��X�
TxT̷I�}L�,�+��}n`���qրߵ���^k;�i�"y2ҧ�<cr��
����~���^4OD�mz�'�XΦ�Q~&��{��Z jدT���-��'�u�1`��U�>��ް	���U4�Ay��jB}]xA~~�X��cXF-d���=�QY6�5��޴ǍP�a�1���pTr�ٜ�c%_K�z����,981˛,ʲ\���g�+�1�x<���9��L���j�}3�g����������Q�R���<W�3�؁.�	��).\P�`�7Sn���ʆ+�/��:�׎*ӽܵ���Ρ��C��j�*JO$�śt�O��r뷔b��](�EY�̵���)av;���*�vd��T�.�-0�*E��%y�F&1�������Jn���#q񗡂Lx���T�A��ğ��SDf����D�JjѭR^��L=�a�o�>����S��/X�I�J?U��#d��"��J0u�2pp�{��x���V�H�H!�^�rW��q�j����~̞���h�Y�	M���'��jZܥ�#51��w���1�k�L}p�W2T0y�6+�	}�: kv�����$���]�ek΁Rh)	S}$�V%��ߎ�t�*�H���򭙺���e�}��3�߸��{D��y`��..t[�w�/�	�6``�Bq+�X�����;0��'����0Π�p93���l�g�(���q��/I�ZDQ�	1�B=/�u���P$�+K��?n�V�(8oQ� ���J7sT�̞�]���d�af�?��G�t�Y���lL���R�t�`_��]��Xrǀ-e���6�4,��!E8�sȌ�H�Ռ��`%�pl\>f��4|2���mf�~�(���B����%��Sv�e4���+�]��k�a�YO�f�c�����)��,�3��6q�L��y�u�O�����e�f*B��S���.KA���|���8�܉��g�OF7��%v�/|T��	C�%��ק��w��9xg ;&D��Վ?�����_s�<G,.�@���T��Id�~�U�ѡ�$ǡ���ٽ?���I�Fr����7q*��0�U\o J�t�*�<{za��	�����Uu<�!�s���/���u*��w�>d�+�I�w�W���:�.��k�5��2�}E;|{�J�/���;(D�0��cɃ�u�3��(��mˣ��Ch�T�]��#^�G���.õ*R�(��lH�Y?Q����_�}7Exn���@����f��q���I�ibw����Wy�{tUG�p>�	��2��*����G��Y��	n^����t�`J3�>��S���I	p�R�$�mP���2uny{�^����f�erC�:~�w���c��_Z=ީ�I�
p�w�x��"⃜c����}Nޠurj�낣�H.���֢b�Q����.ɶ�G�����qh�#��t([O�$)7Mz}��p3�� B-3z�k.
\�EI�����Ad������lo�%���� fOzS*l]�;u�\��B�0�T�oߘ�����u�2���0S����珠wm�2��'�ɚ����3΂D����9� �o���O��7�	�T�2h��J�P������2��6>�8c��B`����	��}1���R}|';`���7���A ���~o6�J����pF�C��������eo���4�g�r)b��]ǯ���� n\`�"������J�66�����d�ק�EY�7�0:y
��"fW��L7�恌�po�t��u;�!D�ؐ��^�N '��St�g�z=v�YC��,?�jB��?�D���Q~�/��(�℈�;�0�f�q�/J������o�6F����4[ �$1�`������_5O��#GpX�g��k=�Kޞ���0����q�|B��^�l�j_}��0u���f�D����+�����U��͢��_�t�/V�Έ�������1�@��X�3�[�޿��j�C$�G��t�ы4BIO2"��,��F-.��k� �t�|���6ƥ��r�^��_~�
g�.���i77OC#"?@�ߒ�j\˹Z�O��gZz�87a�R!w�@F	2��H���4��&4�N:�}�V�� 5����Qn��M�r2Y��No���+t�ǹf�/��;�jt�y�,�ԱٞJ��;�� �������o)v��Dn(II&��&D/-A��[A��'o��V���[w?��VÈ�6�ח����sՎ[[�#�UCJ5|���u�ͤ����5��dٛ=<@���k�ԓl����lhGюw���S}���V�*��˄�L-.����h+�i���I��wؚ�A�D֗�}��n�.onH��z���5�GaH�_��� �9���@�d�˝qȚ�� 9Y�:����/͆"��/�����j(��U�ϰ������	�QQ����l'�<�d �kͿ�{[�U���J�т�$��&��KB���!p�J��}j�gjq��f����.���^ֆWӞ��1R[��!/�xR7�zn��_��C�ut+T�[�*m��
očXމ����O�Q��\��wR,)g���fxf�$�|)�������nh�T����/��
��?�CI'(&>�<_5�~��pt��a�����+�\<��w��J����u����^}�.x���7`J?���<8��.0 ��k&7.���D.�-�y����l_�[߭$1D2x��n�����y� ��9���- ��mHi6&���/ua�O�>���ßan�]D%�h����i�]�����I�02E���Z霰�x1�Wig�<CWy׀�K�!�cO���]FI�0��5��V�BhW�QW��N
�����0�ý�^��":1��a{O$&Z�/g��)�wyh�w��̲�����ݷ�{���Ouej?�#˓onN�r�C̙<6NiO�%K�gP�߻�8��$_2��d�9#q�׭��kn}�A��l��@0o��ǭ�X'��p����2J���]�j�1��gV�����/���P�E��S*!�� ���4�հ¤��|�W��ٚ	�m��;�4�w�d��D(˨{W~���i-�4�I�u΢ɚ�Ʈ}��g�,d��f�5Yl�. �c��XG�ղT$-i�E���"ytW���fp�����ǌ	�Z<�"��x���w� �n$LN�Wu:���O$�zv�q`�
���J��>f�AW`�9)��SH�`kWE�x�����1K�Fƈɽ&W(��B@E���Qu���� j�Y�^��J�p���`6�P�E��ǜ�D���q�h�G�C�eymC������a�΀?�����3p)��	���Atk���������(`޶/e��� <�D����+D��X�в��ن�&S|��l5�D�KM�%�ny����'�zW2�6�D��,�w�u�o1$�x�$�G��*�:�^"@�!�;���*��Z�R(����aAF�H'���t�6����KG=��$H��Y�_���j16�������	,����KǿAs�\C�űj��fZ����rW�^�,̒�z��L�˥� �u��&���xc6��GK�N��r媊�{B��9h�5�rj�v�@�sh�����{��=p ���N�atm�?.ǼZ0N��	�Ѻ����D^%1������f�JK�Mj�w���T�+�����$�V,�T�^ؘ�ceo/<fV'���JP�tfM1^�-c�������X��H�Y8=���P�ۇ0�$G������e�υ;���o��IJ4R�{:e��@S+N��RK��'j�/���8�)��cԿ���l�D��>��I��:P�&_ki��|��x'���D����C��	�����L����3B1tO���lՓG�)h�q��$E�kG��zW��СZCk{8G�(�!��G����%�H�zp�����fB7��W5ID$^�\$�5Lci�����w�kTZL��ݛ�����|ޜU����C�,��;��x �0�L�Q|a o�����B=�m�{0�f��o��Mf���8se�
�3)�fBɅ1����廲kl{FZK	Ta���	������d����jRmM�9T�IW�# B+k	D�u�/�~"�4��r�(���8�5��{���_��bT��&�YlG趈t��OR����t��Ҕ�]n 2�Z&@2Jo�hx�Og���� ��ˮ�,�8	\s�'>�D�v-��9�}ⲖL:������_=Ce4��W�Z�&j'�6��i��i��IMc\��1�t�oOX�OOQ��~�i�n��߈��J�<R�&[˜]{�B��S�Y���=��"(�����g��u���i ����l+4����(���H8Ѽ��"�/I8
��c�����M$&�a�r��a�΄���Sj��e�9���N1�s�|bz�"�C��"����u�!j��|��u�l�4��J�>ۨ�"�ǲZ�A���F[w<"�фX��2k܎�x�.�id�m�����tQ��ɡ���1��O��-�A|i��	��.G�ibG�G
���p�vΔ:ե�.+��J�������`+_�K���?�A2Ԡ2�;;��x]:��u�	K�p���-Ujby�v3�m�R�w8_��-t��u�l��{��/O*�%E�����Ec+Ff�p��/�J$���� Z��,��N������+l��4?�6*Ιf�!8J������kv���/Dl� a��Hf������fƯ��pg��?�Z�%�k *�KYy�	ޑ	r����S�Zw�Qs��'W�#XM8�@k�f﹚����۽ھ���f]�4���ۥ�
Lm�a�J��ߎ�xc�Mܫ�*Ѥd??@��E0F�t ��%=!�����FC���P#����7����_���A>��M-^�V�rj����r!h�s��{��5�y9��3k�D^]�p��t�5��M>��Ċr0�Ǖ�N�&��R��CvE����		7�Wת\��M0d�T5zw�y�-�bo2�a:#U�w2��~�'Jt}[�20D0*r�L����۴2�]�Ցxa���-V�ռ��&� ���=4�������_A(�0׈�e���&�U'�&�#�4xD�r踢�z�Ym���{�"vQvaަYм�ȸ7:Y�'��3SeP:�񃡯�sq�&�d�͔L�ZxZ����4���6�A��lqV4��MGi��71j,�����KK�6���-Iµ�E�V��1�7�<V%eI��������I�*Y���we��}')Cdr�,�F��[�QH��|�''��>�����+�:VL���R���ɿ�AԢD���V
�9�����(g�3u�ٳ�a<�̭��tG-xVmҒ��2�M0����a��7��e8s�%YCA��Y�-��ե�V ���4R�E�3�\����a����\��J�դC|���0�
���o+S9�b�������}�T�?ns����N�d�Φ�P�Ҙ�e�����C���:dX�WI=	��/����YXQi'u�{ҎZ�{&��F�fȪ���֌���|ْT\	�����f�"5,�7ോ����禠��@����	'UVd5�J����aH�P�
a�����]�Жm,a� ��w"FRK������~|���W%/���;��� "(S$V�fXO��O	�N~��
��D�����"N���/`�P������heu�]�� �y��R�߮1|�j�(kI}��>�@�YxS���mBG5u�ѭ
`��o"�Sz�,E��7a����v�XH�[�;`����$�À���V�n��`3�R�G�Xɔ�M҂��t�̠W�*>����Ӆ[0�0H��֦�B�X�-�(��V�[�U�_a�{�cU�Օ��6�Be�z������ �J��PF��Ԛ$�C�5�l9���U�*d��I�*�������m<i�V�L�]��f�RB���
T��:׬t���ŻO�,��ح�E���}���)Q*Ē���A��hQ�g`��j֡�xr+�R����E������H��L�h��ex�e}��T�����Aw1-��:���G��q���
��z	�];NF�2'�����`���=�|_��Pw�Z��s���^5|(�����J���ʯX�x�',I{��	�;�.Q�⹌�ɮ�����l�^'�?A�#�_C�!
t�(E�е�	0��%�~KԮ\����5�L`��Bj��p�s�XRq�T�M��Q#�k�	�dG�ݩ
%���k�b���Tէ�Ksq����F6mT�_��.�ˠ �ɑ�]�4�p�1����UB�X�G\dg���GC�Р%>1!�6�f���k�j$�%�ut�j��2�,ՏNE��������>�����»o�Vq�͘_��e+@;i��'u^�R	�|뤐�t�>��h����Jl9mG)�N��>���V�w9�f�7C����ϛĖP���IfL'��F�����
��8�$�JY�r�����b�wjs�_�abA��ԛG�*���Rr T�"H7���A������a�T�
E鸓̀}�K��?�~�g�4��we!�����&��M0�Cv�V�ܬ��Xہ����m�����B����7��s4��/�mZ���Uܸ�mҶ7��F�;l���H�e��-�A��,T/�#���Bp��f~X)_�m��mF_�Y%��W��a�H�kO�l��4'2�Ny"�[�U}٩�PX��Y��pK�H�����c�7򆐬�j�2[�i�r���p����Yph�\�&�IJ���M���ʴeGc�~�`]���q\��A����=�c;���|�� �����:��<�K����.�>������uє<��	$��)�uJ7��i���ϪfW��y~OS���d\_ i��ʏG+���lU�H)ŃgS䐭Q�Re*�x����ȃN��Wl^A�������b���S��eW=E�Zg����3��*6V^},���7iuĥ��?��΋����;s�f���t=��Zr!+�a��Ӻ�V�0����&Ę^���Di�<��y{j��X�D���C�+����
�����H��sd�l��"v�.�W�7�9!j,_�S�FQ������[ng�'J���¡�����������f�k�VcE���9qr��U<��Ek��/�˥�87����W�i�'��3���1����"��p �id; ���/X�_�	��2���cı0��|���:v�U��7�|�76�*w�p�\��·����*�+^\r�����/9��'��@3)������M��O���kШ���PufO�FHx�9v}��)9�X� \:�U��rMC��O[�z�vi�ָ����EL:.-~!2��s;���:�x�0�s9H�o�*�"�ʉ@�`�	�۝�]*ތ�tK~4*��70������a�t-yЀ׎�>FO�Z��y:T�.W�a<zb$dQ� E��^DWql���UɈ���LW�mK���/���1ͥR2�U�#����5�s���k�<پ*X����|$u}�r:gA�ɷtר~P�Nk�|�@M�����h�
N5�q�>۰�my5�5��z����(���U��O�Q����ڜ�ӟՈ�]�n�V�g���혦{d68�篪(H�R'� �3�Կhy3W»�N��6C0@F��*�oa�ô�,��|�\���?k��v��	��U��CH ;��XK�T���lf�)-�jF=}��xa��tS� ,w;�3#
�J��J�{��ځٺ39)U�Gp;��:Q�T���XNO4N�4 �%b��,��\�KS� s~�eq��FÒ4�xv����'=�=T��T�p��aEt(�����q�������)�������f��[BBp�f~MW��	1�xB��\�p�?P*��4�W�,oc�yY�l#����[���w�h�D`  �
�n�Uq����־z~])13��n�*|>	G_�iCKz�
٩��ݡ9��b��8��[��Z��GQKk��)���F���n����-��5:����ֲ����E�Q�}ޔa�Vu���HOwI��_R�C�6��h]�1�R�7sQ!���A�b�A��Zv���|�hva�)�-� js�:�eX�{��e�����Β��A�q]:Ϯh �`^�
R���Z��[�0�[��K��B|���t�e��c��*5��'!d5��L���%�G��ƹ<�N��h<l�η$y���`���t���C�1S�g�M��U��Ft���w\os�Om @y���?��v�E�ǻT��L��o��S"Mp�t5͊',�xY�+9��n3���ɖ&�z�?px�2��}�y	�N�f]�h�!�9���y�|;�]D���)�2a&8�U�ƷFB�8���O֔��+9'����}���k�Z�8Y���qÂ����!�.��Y6y%fM�5��đ9M�pε�f}���	��X��"�x�4�2��NH�;�� m)�@�:ū�<��5���11��d�U��&&=0�B�����{��AdT↉ek�!���%��\Pf1�g��<��	�oI�Z�H#Ag�}��+`����4���7�Q�;mU��,�7�.�KC�,9���mO�yG�긄�RB��t3:��c��.C�g�y@�nߠ�$�f�	ӵRN~��1�<s���I�2F�G�Es��O��(�Z��{Q�~k����u�`s�m�	hvn�]=9�"��/�Rŏ�P�ӎ�����Ts�ER\�,ex���ŀ�y�/�Q��n\,��~b�\�-� �|��=�7���`�'�%��X�L�^����]�����Kl@!l�]����c�:�wOi�e�t���-��%'�Y�V��~6=��-©�s�q�}ŉ�ԫ��H�y<�^b:.��ﯮ�cL�k��M0k((�d#Fm������Ì��&�e0��� �g=��XL�Ў�����>~2�p�ZGE��X+K޸��rd �`�N�۬W<6.g���K�e�Km�).rf_����v	�5�mFSn�
D�����G�٥W��� H'��#�6e� �o���τ=���w�\B��&���_�(�t���w����r���<ŭ�57�Ф�^�f��t�?�������כ)o�6m�Q��#����Z��Z�K��;������rk1_�W��l�,<ۑ;��5c(�Γߡ��D�1��\�������uHgi�1?���	Nq��A��;k��=n��xnۨ��_x: ��y�G�D�|cc�*In��ފ��ߜ�������J���&@k����n5���SBCf�+a�p��.�zp=�/�qn�J�+=B����>���sx���En����.������??����z�ٝ�ݕ�5n�͢^������^�{��AS*��R��������#���ɣ�6Ү#����Ld8n��,��k#:�d�,|J��1iV�y`����5�}��8p.��Vml�񑮸�kx�yx�Ju �n��F�\˼��hB�[Oo��z��M	������T?wLOG��c�|�Ƒ�(��C�.Sӎڵ�l}4C��<	�ᏴAm�#?`�)��xO|��|e��S�:�<J�)��'�ڙ\ 7uT�n�N�I�?5��vHnfe����j��4cU�g���b&�A$N��uMF#Ku��	��iB׻R�> ��Y�	]u@3�0�S�#��XS�U��mn�]��qj��%���+i:��+:ބ,� d����5/\2&�!rub�i���N:�u,tq:?�g 2G�%е�iA��u���vD�H"
�L(�-t��ZM�` �*�6ܵ @��"�����6�dy{[�޸`��4qHm�(}������Ө��
4�$]>!����3~�wミ���$�`��i`i>f��k�5A�'��^Q[��<��Z���a����3�����#�9��P�ǹs	,�ٹ�4��_дU�<.�r����Ŀ`�����������r�ٰ!��#�!oM�sU�U�z_ҿ��+�[�D�N_�K:`>��|���H�h�l�`rT+��U	��h�A� �Yg��ǧs������?w ѯ�,�����ᒣ(�_����^�<���R-��5nus2��_�����N}�����?�JV#�����(��͊/D��������9h����7��d!��W��4��D���V��q� �%�,`s���Rf^<�n����w?�{B{x�w����y�%)tum
�iF{�� j���vdU6��V���o�_?Ĕ� �����
��B\U�'.�������Vխ�WT� �ɖr�X�O4ЩX�)��W[����-�o�&[qi��{(	�,��S�E�9�7�8��l��y�F?7��R`^
��0[�Pm{��"�֭#�ڎ�H��7��^]0.A�9����FQ]q�ZOU�=����}K�uڂ1����]z��/oK���C��W�R�(]�<im��*h��+����-�w�R���9G����I1��L��ot^�VV��*�
m�g�џO+�].|@H�ն,�.�n$�3��}C�; ���*�&su=����r)�O��H�S��w��IZx!\��o�J����Jk�c^�e�MG/~�z!}v��t�fho�z,Yn�w0Nu`@�(t%���N� �`ө��C��%�Vm��#O75�I쥵���k���iʟ���y�|�Ũ(�츺�j7��6�%��
5�
�k>�ک�7�[s)DV��H#�P�����#[���N,�=��UC�p�����qe�a��&�O=�g��KC�wn�SN���K޼ѵ����=�����2�1E�3W2S�YU��e�i�)���<c��wNo(�D)��~��1uW�\�ϣ�12<4�Q7k��'��l�dHD�z}g\����,�j�2�Q�wá�	��
�CO�i]�]m� Χ_�fe�-}ldJ.�}"�N&�VJ�,��G���b�,~b�=�lH�3�m=B��Vv����4Q���:Xm�bn�2�'��F��������3@�ַ��/:v����c���M�T���I���SL�������I��M��[����cb��'�}���Y-}��>�(\s��o8g2-�9��\�2\za�$U�x��N8t^x��%m��+�Gu�z$-�s[� ��VQ��«������Hd������y��a͋�����E`d�.&t�� �|{"��,M�B~qI�a_9�>�7g�oB�as#
C��~�>���3y�Ƽ����;<*�3H7�,\pYz�{�Lq]}�]䈡���k�ؐc��G&91^��1jC��g��R�u?*�w	-)bS/���t�/d� {Ju4���9|�h���C� �m��H��y�d��<+x�t����t+/��}F�ޮWy٪& ��^�����c�7��#�w崤As�"v6�* h����t�2�� �+71�j������
��|���@L�u)C�d�qD�r�����&jŤ&}ڕ̢�*�8����=z����Y��l_�������.nn=��jQO��q�zy9�R]�h�H���D�ED�U$}=|V�(�a��x�;;u�H�"���Ɖ�K%|�1�!,�-4���+ֺR7������/(���QL�p�E=oo=ލ�dBi[s@�:��Q_İFJ���\�M�i]��K��鷕Rwp�K�(��E�����lA�-�Eɧ5�I����	�H�,h���{�;ݮ;��}����մ��˛��g�����m���=�^~$��O�㽠V.�n��!k6/���0PxN�n#OBr�\�践̤r�����H�:��)���������+%m�'�T��-��0�f/������|~�ZX��y o�@��O��m$�A����k�"rz��{��."�����ա Ud�l0'򪦾�x� < �e)�Ќ��m��ޚ���@ �6fjvu&jw�_��a4cS�,=#�lt���M2s�C��*2,�x���w�s�W)>���㏋�����|��<gx���P)wCwB�D*cgA�W�]��}�JC��&l1�D'Lq����ߦ�����5XzZRFiž�L�y_���~�3c��	��	��sW�+���P^��i��M'e�X��s��J����	�%ߋ�g2V5%$Qu"^'k��[��}�XaF��'O�W4y��X�K|�ygw���|���e�&���r��6����nf`�ǑD�Z(�f`��J?�~3`�-B�b�nכ��oq�Xu���un���3��I�T�@K��$�J�M��c$�=����9� ��;Ha/� �Y�n�Xҝ�Y�/Ķ����p��;8Ʒ�������?~=��K��|Ҧ�o�ڴ8v�:��h11���O��$��\��9l6p*v{Pw+�6dA1{�@9|���G2�'P�=pPX�=]
���
��J�jA�8ْ�+dU�d�|��&Gyt!�w��jf��h_�\���� <(���xAf���{)T�))T��uȍh��È&p�g���RkCV�l�����B4��7�3gv٬R�Y������G����Bp��D��v9��2� ��z�--�`ń�n��I�(��u��Ȣ�2,�yy��g�LR��Ȼ���LE٤W�r��GP�V�0�t��uZ��?�E�R���z:�h����L��&�3���1�Y⿖���������J\��u!t9���[;Q�l�A�d��]�����8��*jt�#�2Bz��􄥙��E�Y��W��qHg "a�2F�<n��>��z��������V߅q�k[6�|d����-����[�b���dFj<��Pc:,$R��n9q����?5N���Vq��6��e7AiC�LqbB����9	�D'�f5;�O�Y6�:{�%F�V��2�x�$���z3>��n��5�8��p�A��lK���7L�Y�1������|��^i@���Ť����WBַ�$=�UI��߷������}���4�@x�>I�.Μ62a�4�='7\�� �А�,�I�&�Pƪz	����q6��6p�:8��kj����|�D�d�!1�����{�JN�Gp�� �ԑ7��7�Y��)��e��~�3��4�Ȩ��**hƐ �]g�g�g�����l����7)�2�\����%��Vgq>�����#��w+��<�:Fq}Ɠ��k��)�6)JŜ�+�X캶 8����
J�"�~��&�����e\$U��C�(D�o��RЋ,;<�p��كP�xM�f�w  1�W�z���!t��%G�:�5q�X�j��r�1"iE��"�QV=FB9F�W���~��ުS(g\�}�+:�,s&���}�d8\ ]�(\��\�"K���t;ԓ�i���)�\�>�z������(��!��IPU�'�1�������l(K�p�#6��������'f�<�U��������� �1���B�=�x���(��J����[�*���js�	���v��ڲ=χ�E�\�����q����*I�B�V�>Xpf����	|��n�Lx���`.U�����PA[�pm�eK��R|ίU {K��,��PEe�a����C��3�P���wHA��\������w;�}��(�9�`��q�m�Ǝ}������˞\��b+}�{�	��Mpc�k���M���:��P��W�(	��=H��5UT��V8+Ba���K@t�u��i$�V�g���nk�y���>�#��Ǐk`v�H�� �S|���;��������ǎ���d�V�v\�5�1Q�����t(h�{O�Z1~�y}[逾)J��z�9��4��������n���Kq�c�|/2:Hk����I���Sc�^�t��lU�+薌�-��4�#�O��2��C���8k��n�7_rx�sZH�Ci*�'/�-/4��Eѽ9�����n�F���R�@Z��39Ը`����%��H9�������U�b�O?y3����%6xJ��__k�3�3�e����:�?�eM��u�sh��C�GWcQo�ca����J��ΒE+����S4p��m�γ/�t���|;XE��Qk���.���l�$�����Ub�`Zc��?� �����$u@!�L�n�P�`�����c��b����Yl��C���wڗV��Z:�������GU(H,�]�.����"���.��g��K'=�YL%��g��=̱;��3���Q�w�}����.�����q8�TQ&��sVc ��@���N{ϑ4�����K��YP�4�����]��J7� -�s�TV	�.k,�VL��!w+1.�;-*�:�S����n���:r�y�
B
]P�0V�H��C������Rqgc����v���?j֖m���(���7z!ˋo٩Kq����wV����yC�Bzٶ�a�U�6�2��e��/zO�v)W�7��
�{�~���ԧ.ST��s�)�����nԂv�u�/)˸H/��B�~���;|/��3�I�2qߩӆJ34Ͼ��AR�Aq���C)��X��4�%�k�xS�v�����'~ܘ���p>���^�^��dQ�i�<��,x�z���3a����l���Ԯ:[WBXI�P� ���\�C�^ǭcy�̭c��C)X,z5y���|?��j��n��S�2U��B�!6�T6�;�2`�`M��̄���!�L�g�_�m�[�p=`q��FKj��-6��q9SC�g.8�>�7S���ۢ&v��ެh��zlW=�y�3�^E��`��;� �F�����:5�L���Ġh��}۷4�ʢ�f�o� ^OP�
*��A"��m�����tNC1��֥�����tK�I�2N�BEg�Ap�w)��w�"U�襙��^�D��ު�9�\��3B�F1)�S���v�̓�\pU*��C���mv�˝$�,���ux'�?�G�=�-�-Ke��XJHzX���@����I4�8�Ѝ�l�C����E.�����n}к�jy_��)�Ұ�r?TuA��Ƒۚ'���?�siD��oF!���,�����3��o�,�����!3<�X\%['!�=��53��1pJ�of%H<���'3�&�ҭ�o�H!�3s�ʭ�{ժ�6i��u�E�����+\X���A���CXf�*	���\�k2>j2 �5@��3ƙ  n�-�8��q��bE!{]ÂS�ۼj}A���%EBCQ��,B�V���.@��F$�K�G4���j`�c\����Y'^�'�T��V�ȥ��{oI�
�3%�/��[��l��"������/�<�^�d����������l!i%nUG7��O�CT�]8���*����;W��K7�aE�����|��*-�z�@{\����P��K�'�����$GJr�T�%���?�mb���Jv?i��1>y�O752����6 ������`~���dB���o�\�<}_�Z���(��9�����m�py� {r��͘?�.u��F��0n��u}��xXF��#�_�T��́z����"҂iq��u�S�_�v�*�R'���KR�d�ʽ���j�!��F�{��O9ٕ��G|�o�|�*���\���@��~����l�ag��D{	�`�~���8�0Z�䝪�QX@]����.�x�6�"����_�e#��څ�)����2��u¥��\���X���62҂����S���Vx�z��I^<�x�cV���v����SΚb;^rȭ���e���g;&�&^� ��>�`}���c���Ib@'>�0[k~�zê��MR�ߗ����wΚwS�E�<$!臓�=ڌ��0�e�5q�P6�`�b�j�-�zbVu�Ä��l=�F�u��'ו�83	=�@_�@l�����-B5W9H��0��h��߹�ϫv�xw���Mf�gW�y����f�W��R%��^��:U�%����#(){t6jG��:	���z�;�#߮H���1*�K���վ���yR�_���U��iɶ�`x�}����2��u��f�%%�L�m�=�D:	����-�B��XP�M�� �Se��*��"��fkbz�įJ3u���tS �ָB���{��K��Z���0�G�\��x��et�#�k���$���;�$��ao��&�k�b�� =��&�w���MSS1�o�P���qߣw����K���&����:*^���
��߂�1�X�����)a��h����vh�Lc��b�a�B?~�-� fi�*�|���)�x�K�%>��l�k��oov�l�k�v�#>�.�RC:�ij��uC�ڼgDɕ�L��	������ nm*�H�A:�9�SQx���Q��:_�ѿ5�L�Y�2�!��xiU����l"xk���l�YZv�ua��u���8�TͲΪ��S�E���<��iViy�Z��>J��)��e�}j��^� �cĉ�`���P��0ق�b�P��C�GX0���{'���	�M�ӤK���K_p�E4&�;��C���;]*3�('�T�s4��!�'�KT��`�ڇ�<�����֊����Y�������������-����f��ñѤW�5KP�
��:�R����̧��)�~�����zeP���9*����]���ݕ"�eh�8�$�Gq�~ ����"��K�a��kg�A�`�S����[10P&j�P9�=|���p:8�©� g�:(lS�����@��х��@�@2��),��C���	J���=�O&)(��`��緃ԝ�k���L7>�j�U_0���9R�R�셰�G#?�ئI�VY�p:2Rh�Y�� ��ڍA͓@ʜ8%�:3�ɡ��6JV4;�ʧr�sAפl�V��	�D���NNmv��1m�`6�18X 
7���+��v*0���*\�qf��< �8`u���m	�!���#9�x�C�#_�~?�CU�������̜�P���TM�C��4�"��y;e@��Z���zh����_�I�|CC:?�,�wZ�KG�n��%����p�	�i�b��5~'N�D帬	�>��[73v5,���4%�N�T��L<#�D,�������';\.����f7fMFo�UA4�nH�{���X��"�Бşu^=�����z
g����|�����"�KE��i3�s2�\�!q�{׏�JD��?J�޴$��Q�8�<���k�n}�����!����`�j�b���
�s!�6@�44���/��R�w��I^_r*�~��Hl�#�Rl�[���"�1�����nO�Ak�x�ຊ1�W��<g]2����9[��+U;�'�,��%��}+�`&�S�%��z�<�T(����K1v���练�f����=�8I�۷��?R�{2��Y��uȠ+����9��/S.>wO\�i��Rn��Z9�M�c��=2�3e�G�p|2�G`�ŘM����;�<S
2TB�uDv'1GA��w�Ksmw��m�z�X����f.e�Vsd_��䍦�(�P���y/#�rA���'���t�[�ﴅ4=����3������6�����	Gr
�|�ʊ3�+�:�����.$ r��:z��f�)C�0���2��D��F�@k�m]�G=�i�h�	aEt��P_?�����>e�zb�����e������
��i��#m��0������|�
C�+���a�7�	��_%�I��Xg?܁t��P\M2��?q0���)vÂ���!t��q\h��w�+���0S5�
nN8�,r�Tġlyʭޯs�]l4��p(.8�סҎ(m�m�yCU��t�U��
��G}Z�Q17������'�V9 �D�j�[N��(	o�W�3�@��b�.Je�L��ͱ��,MQ�RQO�oQ�1��o�x@:�|�.��pv�^��dki�HƑ�oYD��-��81��mlƹ�\���2- �F<���q�BL�Ip���	/�hO�{�/*���.v��ՙ�T�����[_���x�7ZuB7��qo#{61��
nd��	� Z�F���+^�-FR����� ������^�� �T�&1,8�5e,9���R^��[I�Ta@����fbn���5S���&W�ln0%�5��ɐW��;�>�$�W?FZ+7��xYKK��?�k��.fl��Wd�!s$�|��F���	r���S:	��n�G`6���	����i̝�[L
�YP%]uЏ�U�DNO*���%��WL���&�O=�A1�"�� �U�M��"1G�9�ْ���D�l�6\����@ޜ�#���sKsƗof"�$q��m�3��j������y�R�ф���Q5UN���WV�]�����8TΡ����mT���c��˱�\ڬ��>�� W{O��VpK��}ؕd/fI�,S�&{m�ۢ�������<NA<ۭW؍�At��1Q�\@(F�;��T8o���+��_g�5��޽8�&��u��P�}h/�?>��ܑ�1��" ���fG�k+k��A���D���z���z��g]<+��X4�T��E�o�dZ�-hP�H��i��uV��?���G2HXo<�(f ?F������>4$�>����o�ࠥ��y���$��<T��2�l��>u���Q
^^��b��Zy��>J|��F�l]?A8�D|�98;Jw�z� 3Ϙ��$�0G�t�խ���S.Tn��^L"'¸���|c�2����(T;J��M�~x�K,�D[i���r �W��f� ުGbx��U}!3g�������_��s�mQk�#�!�p�@�����AB;^Զl:'`}*����'`�e��z��Қ}�%|ee�y���;��	��D)ih�AY����$Br;w�� � �t1�Ut!c��8��Oa�:_V�rh���E��
1>00�]��4W�T�2���t�nlG�L1%�vC�IH���N��U��bD�I���4_\����v��Q��Y��;���T���p)Fn����blkcz�E`���D�>�/��W��ds1�7��E0T�>�e��������'�h�7�i��vڧ8i�ćm:D�%��\���=C[k�R4v�>�9*qx0�c��c���ޟ��No���)��}K��κ�Dl΃a��Ԕ��,qtP�V
c_R��p�za��>�Bx�a\����}���j!b�`��i,UĆ��[ԾT�_l�������\�����s��v��� �pل8��hH kJ��Zь�\�]�%n�/�tgqJ};t�2���.X������lo��=�!�lr2G�l��$M��wI��
��e��'s�y����)��DL��o`��;&��8������&!�2�z�2ܪ�}K?�)��BI����/is֏$M�q���0�[� s��he��h�W����čMX�dC�2�u���D�V�o9�}�Nݎv�t2_t����/A�<6��R�i�M�ܧ���AݡJ �KĲ�+������_�����V`��D+�j����+d���Y��7ۨ�C���@>v�"�U��7�i��UO`�9�������;��%ƃ%S� k��c����(;H��y�\Ԋ0���܁o��!§P�x��8����8�\��z}x閞5�fw%���Xar�Tz��i�ɬ�Qf90u��
���U�;�O1>�q�`���,����#ަC��2R昵��O��CM�j~��ӓ�y�ޗ��?FX���cUʷա���T@�Y��F�v/;{��'�H�|ɯBD[�CKn� �I5�v]�����\M9Z���/1�Ԛ�4�b�Ti"&S(K��@�uk��/�a!J���$Z�Ӓ��P<_��ZW�c�� �Z((YU��N& ���������҅)|�о>�T:M?�*�պ��>%��$�2k��ۖ���7Q����&�-�w��$�r��al�qY*����>�b�<�B���EG�˸��l)�q]Hj����!���n�M�zM���K�#�W�D�#T{��d#�#i�nf o~��Δ*�y4)�Ph�+L��#�42�~ؘ����5���=�QkU����X��=�!
ϛ�|�����%*cv��#�VT آ~�Fl���V�Z����? �m�m��V��@�u�����{�Pb�"�ĝ7��r@�zʐ�u��f�u������liE�4���w�à��ح��X�ޒ�VO4$ @xo1�4��!�)�'c=�{+��G��.\����W3&�t��1?�y�����n)����2��؄_�\� OLrAsK/o�ֱF���CX���w�R��S�����I�pw��0»�
U�Gt���*��3]��G�,�s~�]߄	�^�G�:Z�B�����!��Z�����LL9xC��	8-_N*D�$d�s8i2��gwF�"��G�i՞��br킻맻>x耴�=��ٟ* �MwԉmM�s/$�j���#��b�|� +�~.r?t=��do�Ŏ�*�X�NS?��-�B�<���wA�Y���j��`PU�w|oC}�'`��s��b�S����Y�(�d(�r��z�����q`1�e33'S=_����<�	 q�d$C�~��F��l}�,9����I�i2<v����y��b�F3���M?����,�%�`7�����/�h�	?�iZ��0���D~�B�p����@�X�l��9�q-�\M�:B�r�w�Q����f=�|����;�x��������W�䜃.d���\��P�t���lgSn��:uf���:P��P��Tv;�	�olm�4��7��2!T����_�9�����%�[ؚ!V�	0G����ݲWA���r�4Bk�=މ�.�� ��	�Rc�Nr���X����O�NA0���,��rS��Qa=��T�O��x}cB�>qk��9��'n�Y�nO�<o8�X��r�s_-�,���/;:����Zp;yh���\��58, �><��(Q>�T��5
��4&�W�+[�ﶊ_ȣ���ٔ�7�gA�V�E^-�D�^���y��Uuek���ɍxmpK1�}��pI�oe(���D�q'���`@�0���{��`m��b�_s_	���^\?�<��cX¹:f��R����@e������*�&����|z��$���Ȯ
��
���OA����Qb���p�]��mi`�i�2��B��v^E�G(��={?D̥r���u���v3�N�;��o�0�ӃR��O���i88L��bz���G�?X^��C%�̝0E�B=?����T���p@�aӇ��P��UN��V�A"�&,�Y�ѵG�	��3�c�p4h�$��� '���N_�@X��Ŕ��|�vdrUje�����+L�mJdu��{�se/>u��c#v����Fϡ�7tm*�n(?v��K1$�!aX׼=-�^�{.[�;s�`��*"r�F`���{E�Khj����Ё~#v���v�M�}�.�C��U��y�#}�H�p{�t��"��W^�����5i$�jV��Ã���ً��&�_�b^!.�ILჭ2tq肛��Ԙ�I>����{n��!��M7���T�'	�+p0�@B2�EjQB!�j�=�9n�Z��4V{�y��[h߶�x�����m�9��$�:�s�}���޵=��DI:^e�;9��
�߰�;7)���T�T,�_��^7�[������V�����Ġ)ӂWc:V�r2Y�hYQ���l�=sl#3����r�=i�`y�-%MY㘞*Cn�6���iN�XAU�RJ5Ea����V�8��!KJ@��04ӽ�&�E�<Ks�kn(`E��=�V�)��������y0{�zp�%Y������6^2���h��ْ�~�Zw� �Qհ�h�ܟ��oʹ�,�h�%+�C��l�;�~	F\ �b�?�}�q=���G�P�-��1�GU4��jƓPd*)�A���������DGW���	���4����AS�g�0�]�U�ӛ��a��"���8J��?�{�K3n՝3�>I����yFĺ�^b��*�5F�w�4�K�^�֬e�� ����#�fh�J�CKR~ֆu��퉻*����*�Q�k����C`�e�[��w�d�����n�
�T�Y�,�'�'��l�3L�|@�|��?� I⃈BS7�.Jryf���������/u5�,0M�/)A���R��!s����C��Fnu��#1����!�&P4&��FJ'���6���{4o6�ּ7Ȋ�mi툺A�������偈��˭�C����$&F��<tD!D��n�::�u�y�5��5��g_r��N�y�r��e<ۤ0�I/����A�TU
n�(Y��炣�2�X+r��ze/�@^a,��wgA�N�ǔ���f(3�}	��$U�8b6�E���^� -Q$q@|��.C�;��ca�L,Iz�у�_`I��Z��%I{p�l�{��}���VS�6� ;�D���6��h�z�&w�[�����8�z�Wjm-2מѹ�8V�m�g؝�8��a�Wj�@ش���.��;��>:z ���XnH����Uf�열�pv؈��T�-\��Ss��b��
��yٗ{-����c���&1�vz���zŞA��/'`���.�иNOQ�S�ij����LQ���Ĺ�XӼ�V����C4Mx�[���Cl^�MBzf�`��q�8�ώ��,�/ �-�S�Ju��'��s1\B� E���	Xl�d�{E/��������덮>[)v�q�����뛴��������7B.�,�n�K���"}I���X�x:!W�:�X0A&��b{c'�{���G?/�����t�G��X��������i�=�o+K�1)j��Ԓ��-��%X�<�:M7��)�&\�(��c��N����ۍ3�F���E��|tt��J��3��&��X��4D�S��b%Cӫ���8��MWRg��8��8���0����K�Øoٜ�ˀ��گ���X�s��B_��u����t��S����<i=ǁ)� %�Ö�X��3�JA�/o~���͓\���G1��I�a(yio@�
bkX��v�����V���#4�zE1/��QESt��S��Rnw
Ն��|��g\6����釋���#t� >JƉ���r���u�r��,�����4������P��V ��d�Sv�Va�u>��Q��+ƃL�X����묐IZ�2�;co�W����s mp�D����+a����Zw#�>}�O�[���Vet�D6X�\��H`���G
	�����I�-{����������H���ۿ��ײ9��a)��o�=���P��=&�+�[m�a¾%�(|[���~��RY+u���Up=�����o؜����ޓ7�0~�!4����R�4z�den���H�9]���}'k����8/��o�Н�1�'Ve\b��-����Y;�@G�5UJW@`i"?D.	���3ߩ�D��.��
�۾3���lJӇ5��/B�>�OQ���͓\�y51���9�SL{.���ia}��bH�	v�hѨ/�ʘ[F�V�x��5_��Z J�v�����8���d��[S�j��r5��f�"�uqt�X*�{��b9ކ�h�!݁L.��V�M�-��<>s=�U�F�2�����������B�VE��-C�O�rmI��S��o�=�%��eJ���cAPPB[:w�)�����7���`5"��2H#���K��z��엢I���vC&�VMP%4Ƽ�*�-ȧ��Zo���+uV��M���DMY�4�]ܳ��G&��2����_x���_�Ӽ�+q���G�s�� A��
��l���q�b��@v�c �����P�����lB�����*J��(.>��j���)0�b��S;7͑
D��A@@N�D�e�Vx��0��20w��
UK���6K�����+�	���ΐ��JF��0	��k�:a��"����P7��x5j:X{{��X.P<�'R5�2y/�j�Q�1��'��GݟI䞁��w��A�w���^�o/�{��"eVb��~��;՗z�r7]�R����;����_���ւ6����T(���Bg�������}�Z$4���+[~x�O��p�'X�.*�g�g��
 R�p�B1ܞCc%�]��#Ɏ	������hB#�κ���ۤ>[ʨE�$�Y���'�H��4	4��$Ƣ���u=v4�e���*��齴٣��X�6�G$��T�UM�W�z�\y��Vs�]@]�Ϸ�Z���_����%��a_<���^��S��0��lZe�����A 6a�h��A��3�'rd����ťn��X)����%Ge�Cϳ�;s)фS[�:���GxD)��uW�$�s����f��b's�3��O"X���U_P�o�g���N�'�Y�6A�U��X��r�h3��Κ��F:�<�`7?�e���?+9� fD�����uk���og����6��'p|��?D��8$��h��ď�^�J��x�,�\�����7/N�-�g�:��Lp�X9{���d
3w$3��Q1e�F�!�*Ai�9��������KXh���7: *�3<�*
�vil��Yoh�c���
�VD>_��>���&�!�TR��-���"YS�E�8���x.��?N�JeNHf�O��-�l�	�v�`/�1E�$�q9Mǔ��bo��t�K]ʢ!w�.���J�-ۧ�X�1q�¿�Eͧ�&��cVGGn�ֶ|	�8y�7�Q>{p''<�Nf�L=�¬�Q15�U����J
���wD^C:.[U�,�ܞu4�M6���R�Y֛r�uP�������^(�Fr9���3�"�`
��5Ϋ� O�-2ֳ�0s	�Y�r����e�_�+J��v0���A%q��Te���9�~� ���))�L���L��q]�C��r����������u����w�Yށ��o�0N�%��Zˠ�W	�U43��_�ȅ?cVqֵփ�"嫰hZ�1���	K}TB��q
'F�6 �r�R<��}C��U�,cd�:W���C��N�+B͞�9b'���Y�K�|�����mX�J;)<���[Q�$�z)��iؽ��@|�����ϟ�E��jܖjD�������i8��Ao�T�V�9ƺ$_�`"��yW�*8c�>�ɺt�T;]�9�2:^<�"H�$
 xhWQ'i1&E�q3�{e�f���P2���!ć�9�c���E}�[{���G��2���͘��ۅK�@��G*�)4S������es�JA��~i¼t����&�Һx:tB@o���ײ� L�}k�T3sŁ���a8�BT����S��#�����X
��$�xI���!��s�!��mi5S�� �ٺH����q'�]��F�z�M�xZ�8TĠ�{�HS��g�u�x �Ukʾ��Y���3M7��@�K	HMX%f�F9��uh��P" s�JW�9�6:��Ua-k�d��#��Xy��<���g�0ֺ��*h��&�1����h�����o�95�3�o��n�����}'iy#�X�z�u�1�7������(�	i	5k�37`2�q��5�}I��>�5�uCM�v��v$�t|6#��c���@��ssҌ)��xeZ����ZHH9��=lHn,�U=��K��չ�����w���Q�Z����ޟ������ �,�U�WO���j�Q8�f��в$���Hh��mNuu���t.��c*m�oqh�Z�r���!$��x����2n�Ȓ�癱���Q��6���<��*�a����8÷�N�jL�\]���D8�	�I��L��:�*]Cl���}�U�.�A���/�~��O������kǜBKl�GbϥFR�-F��*�|M��r[HD4R�9R}�iz	y����.PG��mz>��p�)t�@������<Q��ݓ6�����i>a�v�P$�/0���Kn������X���lK&��m�Yc��Vn�;�P�~�7c
��.0�#�@�[V�\��"Y��5X�~08�+��~}�7�C�^��cDf���֬���ɺʪ��υ_wLQ2a��7`�dا��z[�������@��cxT�Ş9��}(����q��� &�P���z�t�o�u�d�f��K�A �1Ŷ����udbX�65����|�%��xk�;�u�8#�%_�G̠�%9q���i�����*A��e���Ye�O1�Aw�f��J��f�>�jR	��%[7�x����c��]�2_;�'�e���*7���W���3.Þ����b��RBg�E�<�I!�ݩE�H�Z�9�#�uu��+�����$�:�5 iyiK��uM�lЗb,n�ϝ�>u�K6}��ɸ;��-F:�����d��������t�2h^)��0.�`#�0Ϳ0i��21��!��h_ة~��L�6�X���{d�I���Od�׵t2n� up�t@�s�DR��0�/�'huA��P�T�`�|��)��7�
��P���.?P���Ѕ�Kd�(�1d]	7~�ż��=�@��ϖfo@B�0��2/?��Ӧ��D�g,��k'�@��qj@=hQ|~MN�c��Ⱦά�4��r�F}��}sO�
6̄�h�0[� J(�<^r���%�HU/�f���G��*���4ܑ^k�� 3`��c,2����{
{1 �,W`����~_!�/�>����>4i-��}�����>ͼO��2Dᶳ�����/�t*��=��O��I�	�j.�A�Y��~ѶK�c��d�C�V�	�ܦ�p�Zg�8J�r�Y|��$r|N���陇0�nBw�[�5(fV��1���Ú�*Be"�0͂�J��fSl��ψ��Ĳ�p�}gx��+2U��n�-r4��G|�YƝ�H�6���1[C�ݶ���s��-z����j�A�\��0�FA�ۉux��]ތjռJv��i��40���ҥBg'���1!ణaiX��r��P�'U������å��X�:\�F3��f �6���΢#XP��?�@�B�Kz%���eE���!���/%�d��/�՟�?'�pY) VG`[e�2c���r^
�P�o	���0r� =�[
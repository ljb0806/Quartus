-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S5ZSIZwTX4ceo8Awp5vZF0JVPKlHB2gEuXGUVUXxhGyVsUDYy4T88Yr5zDxhoPS3S9KDHecNA3Rn
5PmXyW2qtdniYqrkPsnzIeKhtex1z15RQcYOLGGGxMEirQPMzwUs7Hi7exp/lYuxAwPFOzBsVVi7
eiz2D19DCdCvZ3xqgYM723u0B00aZ5++MgWu25tp+laSgZTUdGtnKLZ2K8PJzc8SII3ae9o8pSn5
Fg1a0tNEwJqNv7jgXVnErMa7Qg0/ITTQm5m0DCjeR72bCUHacDsJDgEgLg5mSpuIPe+UjxI5ZhSa
jpArBtP1I8jh33FnL6uv5nFwSyh+rIe8bHu2FA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30096)
`protect data_block
Ew1zNKnw0qn0aNxO9Ep9U/KF4B2YqenxIL0B34paZ4woLMFbOv6I8Pu8vnVJXHdkBSB6C4OubQoa
QbnfTou/ogYDOXk7OW79Q3UkSpa9E1cI1v3pNqA0Exa6naVxLWe32DUrU7g1KGEXUKQZ2qlnhlrm
VaWnjmLY1yEa7WOYGxov+TzbYkhPp1gmo2Ptr1luBcjv0LMcg5yb91RSmZnWzgr52mQKF9dsaA9H
dVmuajmN47RYhShNpHDnRqs30FDfhHkx/HrqzpfLOcq6/r6RO9JoW2P4K6jqNWDPv0xYai+6aGV/
y9O9FDENowpchh8cY0lAuy8Ktd7eUMvPSU1sCr8UhOK6WJyLDYjp2otSFGLks+9BvcBTCrAuOKcD
Gv7hjxFM+unvV/t6goKLq+iN+ch12geqTJQQbUzHILwLpsMIvRgkO0CNcQTSZmnek7+LPyEpavu3
t4rKjjUHLWtlCIK2epEXlC1yuAOfnPTZHKdKo1TTYO9z7XijWL4sHevQ7NZHA9xiwEhEUQEp3+/j
Y0NMyOqZKTs8hmRlTPLMrNGg+dX3r4GjenIawYszTDXlys7XIzfqH2WdD7bquWOm8HBF5VZWfHaS
Op2Gv4LoqQtkro7ifVhjZVDzY6toJaMULB0NIthhew/YgRBgUqBnoVAGK6enjKuWMAkVkUNVlPzL
2i9McykA6FxvZrPbCjJqVqx5ZtT5T2LS+oIaJT2cK+TnaxPQToAIPzGxKdeKXOIp40M/oFyCO6da
rYL88ch5tOzDUPdwshvJeorzz7cmIdkIaVl57Ie6zL1l7VZ9sd+ZHXyVPa5xxQtmtO8HzPOjGDWZ
NfOdlUP97Hi0eDMl1JXH+I5mPqA//H4Od/OI0+Y7Ue+FUCVBOlRXwMegc56aHJyU9ne90gwFPVyK
4508Sz3cOXgdz1emoFpbrL5jFWDAKZ/CGPyHLxnrTP6sk7mdprAAIil//U5Ee+nkmYJFcULcC+Ih
9UuZ085EUBswKDrY1NxCzkplSzhG1FeuCQO0jEQxPWZ5sjJBfe6W054JYupIv8W3v8yuH4rx06pr
D+2z54LmS/3tbN/DjhfXJ0rdgxS4PAPZEwt6+RoFR0pBvZqWuf41YvQBh3DJ4CXTOz4L00KeeeEo
ouIeO0RqlMDoXMvdJejMm8/x3Dv/trhWeIa/keGnK/YN11JjzGDR8e3xFC1fTZbuExPrQKE0a2lx
6s0t519EOSJX9KJOt4aUyReJIm8ZtQWOe+gtkZVnWTCY37j/6w3YRIcE3ssnKsuRuJW2epifwGSM
PUphY6tTNAR9JD/GsjlyQiswUkv/3m5PDaAv8/tiT4tbIOfmJwp+V16Yy5FJk4memI/iFw58ESeB
xH+aQcWdHeuhMUGv/iIAbj3bKXu3xWSiAzYuWhU1W5X9bM2sq3zlslLgtLdD//2RXuavpn3/uri6
tZJFC5hRQTTymud1zWAjNF+Bx7lfoUAm2nkEFZzkmlXBz+RAeHcDGfdVr23usQ5efcQxkhlyEPKg
xLQiAnla5vF3oLoSByceZDOzyHajuPEniVcOPVwRyfvB+YhxvXtXD1yW3T0FOiZmoAmPYrzRyl/b
2pZEir/PiZoku05HInb4r6SqRJWpSFwgYnRC0vn3Q4992CpvejvEuW9naSwl7noWHcQQWiKfMFyc
KGx2Dn64T5wrKE0ButcJJCjH2RG4ABw4OGwDAtWBW5bxsijCKEsyC0BbuQdh+0nNeWwImyKS6vpU
vO7pIK9iOCHBVHvTePJeYh7pf0/+lXRFBaA3cEALuep2PDhx8Is5qWSR3RN+SlsgTBtu4Fn0BVzW
BKFuIYueZ7o8k0VCnQAX/1mQKdnGt7nDsVD+extfE/pLvDz7x02CW9szfjhzONEKuh2747zrjF1G
DUIqf3CeNORTwJPcouWIXRDs3s9YvCDShdNtPU/VgM+o/kNy8yZJs4ZsPxyhKuEk/eeptu8YoldX
ANZJTRiK9xHo+v53yg0NsdwUdHEAMVVf32YnfLHfpyhTwXYVB97shR2+fBKDnZ+xhOhVBdq2SsHe
NwwUUXmhcN9JHaMBKAKjZNQfkDk2mCroDLjw2XtgqLrPdzkO7ow0n5xwmuvoDST8PfpDJdzbejig
CwxzBVmGgAHZY7Ccb/SDzvjqom9whyi/H4qDnw1rGJCqh4cPlf6E5CDYwByS1w0UwMbdL3EUiiCy
h37YwKC+ZHW4929IYF4J79yerHup/YH01f6rXef7ikXs3FbiWedOfCzQG05/KXy+ZIfmNo4IKTLU
aKeVB6zqcEwSP1IkdsDK3m8/KnVco9eVvlgYFzo8M5l6qdci+zvFC+5pxtCOjEJ6zGrlteOZ7Bqm
IjavGXN16sbPHsL3jLgROWgcHeBxow+EEjVdp6X0LExX5084TWhnhbPZOzD41iBMc3GQpuHEV1DW
vGr3RoPMbvi8WMKtvy8FpB8NDUzZPhMIXhcxhc7AD+IvHklG538EGHPT8sYSvq+G239IM/w+ag8l
xM6gMJHHpvwbE+rA/IaLJCcYON/0JP9e1JifbIAaSUAaEYpNJkdE4/wHH2Qqy1qWhm0aen81bmDR
TyB9SXVfN2xWadhm8cguo8zu0PewevRhnNxLkJheIn7XKprFceILvmSHV6dfheErL4sr7XeAV8D0
9tXbxXr9uF+P21Qr/iDhkdOPV6W5B+FWHsXbBysFszHkQhfSrBGojB/4N2/Sz3xGCL8rbvf4pVAW
x7Pef+u1OZukWJ6ISvn5pdQg1fmXXkkOH0tXkkKq5nJTrf9uDlDSVLOJsUEOGbqMfYgtOxPIUoxm
3NMUK86IJWrFFsrUcCdeDw04dttRuYlSC9CP2wUS96BbZCKIRnPSi5u7cV3SYMwVkal6Gm960ut3
JOvPYsyk+nj8EahAZo6o7NBlhGmvbsKnmsF8PICRuxp41gHyIULxQuwVLFWCNFDrNVsbLuG0O1ly
Uw0i4ukg0KiqhNhMSmnYngSYdcjPAo0vYyTkWz1naJX0qkut4rfE5aCSkd3oXnpLvQfYeGpgM+lc
Pg6F9svymOEqDFVN3Uekosm9KB8GurdzZiPFvXVCQP2QjIWf9IT1DMpqxqfoaQ9xnfPx7McXeXmU
/l+AGAt+QMouUaYO7lP4GeWl14mjngsmZY2C92J9QIGgjWaAa6VYXLhK+K4EdkJ6WaIlA+tNvikC
oDeFkn9P1xWFMJRVmHcwiOkJ4JQJXt0/L4OctGI+lZgI20eHho/fEnNqfbUdO0/neNWunO1v7wbs
bQtAEhS9GI42obRxFVBP987T7CxSCki5CS5D8frGBI6JPJgCkb8TP82S0tMvJwgjHqgH+RbgRXBp
xcRZhsCTtNjfF2y6+3qxo6aO24Bn4TPmyED4Yd17bmEdvNII1LMN6YvAXKum9ny2/Mgxs+XVDr+L
V61qM5hq8r41+uIYxZhHLdFD5JCq+MLZCw/ciUPOIzHEX7G3TbCq0XIwWQfAp2xyyCjLbqGhO73e
6ERZhzLK/ItTgZMTdXSE3k/6VCcTjHiiN9BXp0COqkl7Xwb4DFa5yKRa/TE5x/hkf8PTUdojCo2k
GymQT8SeB9Ez+EAF5pcwHcuADf3Mp5dknT6R/tvO0zq2e13tN1zNKKz0GMmmFxnRBueso8feqmaT
u8ugfp5r0DtYERAZ4Ih2iTAG495kb7BxEjlHKdTxCMN2tpFOe/DJUwShT+OR74nWcZO4H01r7/NG
rRfhMKHohVSkzkNCmkjlAZtU5vRgXQXTg8NUTYSWtR8GpcHpkNBqD7FXUMKVERbYSdkGfjpNurPk
JdysmKz4OI5DP67/HGowmDHdbfpDQoOdcRk21Vh8OQ97Eqfo5L3lBhG/JhJtLpAxfrx0JfgW4p0z
fywfGDkr5XUmMtqmrtTWouiyTLzY3ioG0pVwKaGobSBVqUKRZ1ULwezLX8M5T2Xa8nMafb2OtOTX
pyTc3ZO6ealwlDO4iauxcZfnT5eqFckh2fA2PuyfWCTjpTydtAU4XFAPRRrirxI9IR+dZE1eTC61
oDykKA3sIk7jV/AGk9QqHrA3jrO0NVoJ94X5fcYZGwhLm2OA5wHWbWF/wQm3gr9ZY8YGEfLl5FHE
sZlbGaBdimlj8n+0+g7nur5Ha3hKgpkpn9q6Q/oj/sIJHFQDwWaaEbQjht2bLq2cT5gsbqswRe4p
/mXB+XQGd2tr6NxLLqX3hyS/Aw9IBvOEF6eqH38HWIgZHeKDFyn2QKEIhfzP8NXkTE0nUV36TSoC
d6K7FyShmldhKEf5ExmVyXBiFquvHA2oUjXxuybvJD3uTUwEZHI0I1AM8Oi9Kip+/6oSxvxAN3qP
8wQ5I+Vix5KN6th3AJFN4og9F+N7tYM/LwBSvkkQD1fJ+7522aRIH5zXrXBGfKnNS/KZW971pImo
5Eqo4oETXtOH5dtCADemWyVA520pk90WAxUABC3ZvB7IvAdIXr7UV8QyRHgsXT/KKPI/5cswtDBq
Sz7S9G/D4kmcID12Yi0kiCi35S0/V1HhdSxX+w36hqGmwboM325gyHqWorwcxUklWUp3oOgW4dFy
gpIqwwa3QN2oYv7GlvKnPuChlrUicyp0TlWe+YIztSwlAvma4qZ9M/d8XWA+Qstp1arxPCgRPmyv
Te9FyFTMfaSJI/EJj0EaLiCQ4bQtth3R/tQfhzEzfNSliQHDefFmkoRMl1rvpodhDrBJDsbJQYxp
dzVxrkR0rFWe/QjatoP5iTdpqpgg/dMyEjk5sKOyNM4fDGRu7xvXD7eTSKQvDkPFxj+lgLrPyzst
fX0aha0evaI3v2U+E78f8trC2RxwdRinIZa4DPQRLkOQHZD+kLBxICW+JcX0gmk7qnSphJUzsAvI
LFFgLGo8YZGA6NHZ0/qOHoEmr+hDZOWvKJ4jaAChaimfWS0DfC/O9YcwPUmpBzi8awjr2wNgsFTS
c4P09H8yTdL1ig+ttU5OUS8WE487M2oUehc8DFHExrRLp9bXHW13B5JQGuA9NiMm/HpJWjVgmDQd
+vHBIT//gVu3GqFKWmfRmSf0ufsYJgLwiwMGCSV30WUSKWXjfGtQF6D9Iikr0iOBs5RuyF5CubsT
wyuLVTCPbLfHqV9+xdaZy7nJBCNoNd9Hp41wJMKfeCuvUfxfSoFrL6Pptw9hMALgbL4fbDkv/AdT
/RRn6Te6jZq3ywR3CsMuWkikn6wKGhXGKcHF9VhUv9RgXnI6mu3djhHNCeXNp1jpOvnuYto3ili/
3sAPG+6feMMbcQr2qdDW1yk+K4gRI6X+lYlRsIfV667ZTa/SuALnXd9Bkz/x8VYxbBK5Ums7tgek
Tr29g6GjZNdF64HqlhEsvx40mA3tMreObtHUAxCO0iBQPqrrMXxHSET808L/06SZHN9b15XyErfa
rigoyhe3FEYfy1bZZcz/xcVFnzakHRffE1+wnhcX30OLxwDsgPFrGLVYeyzIPcF4fXsuuBF8WNk4
VOdsDetSNL3vLw84vTe09n51zxbqTl3PO6Y4mlYK1CKX4zkRihLK0U1qh7rshph062ZujQOxdg5b
OMAqpI8Zc64ZqIfHaUUktUPYEmUKWZ1ujKq1zLORBOwmmRLSdUUorOmU5ruADVYQcS8TNy+62goL
OxU5KtWKdxVfHVetgQ++VmDOKx92wmqUM7O/3tQ3h+FG8m50s8BRT+CcSa0TNG0/4jisudpS2Xvy
+S+wW5nt4jMa8eiUlsZmgfIYQ8cVyM3edYe5y5jgRTIbM8YBMQ4vLLhyQ7eYUUC4vMalkFVlHV/M
bvy7263urOVgBx0Yr1DXqP//LRExl81J9gnFu/lkdJZTTNvj2RLyYZRoEtTAcu1ui4Aw6neclVI8
D2prqe9iJvWg/FhLx3HnwoClsbf/3507oK+/Z8ASPfjaeWYS5TKinmoiUkjWNTLb7Auv4b0tGBA3
xKUnfvSFoM4HEd0LSewL3HEWGgx0sZhzj4KJXdccVTU/k1eyUaI6V5IfWfWdfNe6OPcKC8uU+7My
SnNHcSBx4UuN5pEKalGTwCspQZvH/Tb8HJtQXCivEeL6sT4KW9JTnIT8WGc0rT7x6ikYptEnkcZo
Ef5MLVgCNjPxy2Qu2Msed6ZIBpIzmVN3TctnQWi2SzxwZcBZjI5CdcTVUReag2aGyIJkSYcp77DE
0TscbogK6vqBOlKf3Rms6CRtG0A1pMmgp0s/oRIqIp/YrAbfKjjoNgJQk5sB2/MLmlc+52ONStSU
rbwncvB5GkSZ876NMj/jj5Kf6lI/LykuCu+DAl1rJ7FCgEcLkHuTUjs38lI2XJVh4ln2RVt0qSKU
Y8iNX9tBgoM7BaGjqdcpV+mZIwMpSywPOdWRN8QMLrYO1Dn3vTP+p+MqxmNY6Y8rBmI20aB3MYpK
cRnjSCyxoghX9mf+tL7wsZsqSQQEYmBCucpNUewzOcy8MolNK9gURhWkfqmAZYdscFcjglNRx3hn
DP2vSo+yPFrobuxG21oLmkMOoWiZ4g1wbvVijbhoNpR0dc486o1ihIll65Oz3VM8T0bpO40/hbKu
RYDy3jvy9W25mi+Q9U2Pk3/3cPPZPHLZNjU/TMaBPpdeUezzVuLOHx41G2FZSUAjgwo8Y7KJJ+oB
AOPawJnAVhd2aHjAh/5EgYxY+22HaoNi2hceSzSuBw6H5FvJJeNtpM2HltZVERNd3Y66ndMFNyJ0
XV4rrD4lvDRRHhjpthsZROuXTkKfJK1Hd9GBO4hwyeNC9H7SdgBxy6fzDEBrH0+5Td5UKO7w+bi+
QChWf76f2VW9oPozBd2ARHnsxF8/AbTr4BJLEjJopW90zEZXoppKlaEzVHL/itzYzpAu0E9NhRuQ
AM2rFwXqqo36v86fVHNC2F81O6PBw9jtQWLzjdCGrDRxbCwQoq/Lbq3PWfyVdTSr4SCJ67U69SrI
p3OnpE2FpAmMobQ9XmLbo3ea7f9XsTlt58YbO7szA8dGyx61HMMc/zzKhMMEgTwzwqrVW7LnhW2y
BSZ1ybD7PO5t5WglZDy78RNwPCj3YwqiQoBRbeqoIYIOU/iAb8HQjBC/jlIm/UIGovRKXNQ6NX/+
RseCwZuZRE3N3GR2YHDHyHlIZPhtknXUtJUXMJxDkO2WVRC25LLeYi7EovrK5+N9AsNxs5HSJo4d
U18isa/7lSlTMDz2K2ZYYi6Yv01PyzMj8GdHRs0Z2fdUHTC7cUZV/DjE8IlComeHnNsJ7vyxFE0s
GAzXC5q9KliYn8PPbMHIzNkMVFgqQhg1MYUShFW6dQx0ifJzZs74vtiXeDG65NJx5XHmXwQUUlzB
HcJjeM/rBJWNlgcP/3Tt3UYEPb54FRI1/RQpuEDXtcyFttj7KzJDoTgbxjQhsW8cTG14MKDLmt8y
/fPabSTTIzmM27Vkn6+F/23gcAVzsMxu97lEb5iMfNGunVSg2XuvQZKbkKgiEbo4V00eJGNxlLrN
a8xlNT5BmvLjzwhzZvoMWX4zJ2QhgUTSk1TaxVzwLGoQ+uLfHTnyKVz759YxsUqmhy6zLlOw7HiX
tPP/FuHYM8Kv8yZ91EAnrwL6TKqafHqYr7t1rON7TP0cTxKE+CmXGgCgR5JjfUHnjC6vf/5SFlqo
UzqylWX1F0oTQROHFuAbC06bGDxk3Knm6k49bm0xP+ltG0mL2+K2Avu1EgU2eS3I02NxNQfQ8ojR
gVrYtQzX/8jaXo72xt/jPHgHS1la6cjuI41uUHLjezXedZc6VJPXF1NkJWSj3x3oaSBr8t2uOQ6c
2f2gzyon7FFnh+7tN+MD0qAjStan6sdN9vGgjRi2TJOXFNnWq1BaF/I0wdJ3VJa3yZKr0DkbNobN
fCZ4u34j+Z7qE0Qxc8/sE1e9Vawj5zSg3r74Cue3UVSyjyUPfLmRp5OkHMmaoxD0UfXed5eaFMeQ
ga9j1ZHVOA0JogEakGiB9OjR6O4vLeOMIWLgL6yie+4RgrEL1IIHELLWBPlyR60ozpJm3hBMGI0L
qXPFD8layuuq9C6uEbu6q9+sEZmXA6IDTyHGDdAOSV+PKaG9GBi1rw+T/wPsGejQ/2/FMgvRoKsg
oLdUgBExlah6CwBCvmhhKDh4gfyml24R/fdh9O/dqaWvFb4DU9bT72Fr1CMDTQANHKr9qkv+ct+2
ozjAurbu6wmwitcBRfd8h+Gi0+NoA/OD5D1Oi0FCBAxtaNmNMG+0psVp4/9ELYy+PuatsFtdUQyR
QhCWHN5UXC+JchYNLBH4xr37RcaG36A3YEZm5pFfBRcOGvX7cHfvc0nq3ZgcJltW9jxOkHatKR+R
H77fM4FxNEXgc0bT1ul9QAB005lgDtwRy853t9ccok3V5hvsZgxPO2XE7wyVP6kLZSrBtFrBZABi
L92nTM7vCnrgE4A2XVjwamaGV8p4qysRzAfLtSE7VFLoTaU/AHFBjm8UL/aYZ52lpQj78kUeK0ie
0WSW+0ulacNj8yo5AGrikvprkbN3u8wT5Pve7+OHijseFPRHqnLYOcGf/wznfkqeNLF6S50TE75N
OTO+CYDABf8WIP1K2jf6GQuJNxUnxr0FdvEG4oAyqSvaFcGcf9o9XcN4XBP8CE4FkBL+uCP2KpE1
a7jz93YBRUIQzxk6hL7RTvDh3Wprqu3AytbuWu5W+cCUcThGMBMXs1ZRrH/pnF5WV1uxFYVU5UK9
rBIrCRCzdXcYvZe8QwzoPBOR+iHC/EkMrjZDoEtzAiqXLNd2GNtFxD8k4CYyzRhcdoMEvLmhTwuM
ykrs/yS0S5/uZxuSsypwDi+7+7jNxAfdpfPpK0WLoHLtSaMSthG7A6/fEK9ibbp22NaZIlmvWZ3y
/fOVtU7JQ0AUgQ0/ybx6Fm45Dqeo1XsQ8DBpA/MoxrF7WcwPc/U4S7HCkFKbRY/KyeaY3aKCPJB4
VVCUexIf6y3V25w8erAv9iPxNh3mbUNZmArwa8vRyVvIWCG1Dp9KDm2Iz6lL4P2yK7154/bGGHf1
O2lf3EBV/XRR+o8/34PvPHs55DRyz3ZPPqeU3NSTfAKR7lncMQ6laI7PQEmX/4hcerpOVix6aHRX
DZ0fyLmuDTTuv/8ybkNribotI3Hfwr8jGmrlIdgmLVFPSOhPovW1lAQyGK0bO5JI25WMKBy7qoMQ
0mgkmGOjUSkYpqNzdSYm4WBuNEoksqMvdvIZRyiuSfR9/CvvxX1EM+Ttj7ZU2vFk9mqqGdzAKPKn
R7IgxratANgs7uPsrfIlIH5a0WKgtG1zxMY2RLFqfJkt4aw02PJ3FYgMIt/qo6CtsHpSxZGrbQbC
Oic9pHwTkCVnRgEP3R0vZ1qDL/9MpdovxmC8Kp6OdyRUmG2IHmxm48hj/j5FuUfIK09B39WPqws6
6H48EyXmwE93kkgX4zFPgKKt7E5fW+ilpM71TxD1QvxzhXMyUhBt+71TWsPJUq/FrRBVmhfC9Yp4
l0OS69Pgps67IqKtw88S70Vl7dhQ1Ws9MJ51zmipZFmEKi2ZApDWjwqrQ+T4tpF+ZShbRVRxV0Zb
cr4YAedjUWDc42ifim1FeJyAXmMFycwj72hrirqcWo2ojKhKLBbZTMDY4vb3hbBNU7P7jt/IilxK
y3g+5/ryMEEZMUFyNUgUkzKDgwRKllKnlzs7BqP+imzdQLr8L3qcNWKGF4m2chPaYCMIwX4UFt0w
9O+AJtjSpI2tOTifeJVAZF7UyvuZ/LGauQKvZ8M9ZbAQQlVXCOE8Q3deAy/Kuva6ZmaDhaUVSCgy
J5UGRvehJLkzxooDyXA0s534Um8jKnNwDOWWzuPEsaXv6Rk6ncSrrvuOmqXHFlNh+OxbHOWOkO+V
qcIz0kImaydix8WUDk5FDnkWvi5rXpEWHSuky1eN6N1U+Hxb887dbRr/rMgE+IFHUHjxJk5SjisJ
HUOqjCfdUt4VXhWnwbV8ju2C6SerZPpa3HUHGIGHKEBr3Nr6pD5+1sKUAM3uQi1khUBIlwhyYQNj
gj1nrmqzQ9mbSB1VP5WM3jhAls+Whg9+5BeOudA3Nz8ARLPwCo8Fn8SUgLCOC9E0UzYStTo1oYyJ
ZoU/SNp/6V/D/Q9xZfRrtGNypDbdCZtzp4fcHmgb2IiDDK0Nk5p4KQ8uUpZOE2CtOSdosyZU2qCj
VrOiVUOYIuCyvbCf5Nyxz0/rIRK7UtuMO6MlG5powOXb+yClQqweVogk3usfyHK4ILPF0lX0wLBm
yvWfdn8Z+LSqanh1Yp4ATTCqsAreui8lImfxw/0TOUzoRthocexSUQMXXnsZz0SDrnSuWDaSIW83
zFthihSz08HaIPclxNRPxUadjuOzM3v4VVXLtGrn/KEkaoRaqtwHWSy6rtMkK7Kc121tp/lEVO85
mdIL04iIDH7vNodjGe0gdbRLInYJKp83JzOYTdy/4EzPMlPeQlgKzoPVTyN9ILPlL/aMJ3CgVvkf
OZY+Gk9lhWz1HRwWEBO1EH2AlIrVGRoHbqYdChwWkaByv2ca9sl37KVYjMNR8y2eASk6ZgJHmAc2
+59Yeg8+7wlo4gTQkkt420UCuQOLNOrOjjBVcOPATnBCsLFxr66K9H7Ek2fszuMSlQmBtSAntamZ
HNPTgcZ3k0wpM0o927Pc4YJ3KO+qDjFuzIsPu+eAaTjcROjIyfDECmawtJ2JmTO+nTCSLeHsMOcp
R6JH97VFmvvp6HmATZCFkc18ppSfEsmZQIf8dtNzUxjzEWJUHQ3jQ2Q5xjEExXgUWBAxvHpB+yMB
zaj4obv72zsMDd2ifkzkSELIRNBKC9e+QHoNGzyEX1JvAECn4LGyl8VtUG+S9QXLiNQiOhtp5r7X
QUhJyVAQ/G5muOBiWXxoEvZQWOiZfYOvsfARcDvrhxajrp04mEMN7wphL+p2Fd8EvIrSBBdfVUr9
y6cEE6Bnuv6jSdUv7JjfBIvocA43uZVWf4wmKyYB3A90k3ZwNO1LA/QC/JkZVm0l/5zcV4RDFNGc
ECpfohZUQ/VqG7Klro4j+aTF8rTzvnpFIgzZTTwOzjcZCejE4xZd0Btk/SHSThuqEzEro6lEiu+5
lA7duHJRev8ql2R5IhQcK3o1yHInuxu3R7wWtNKFQzAoKUsCSWL1G59h+L8M+d5WLEqvwDqX+cZ+
hsfxzoJGRFULtHt8Tsd5Sy/D2HXU39uxRCKDzrZE4SVf291rya+gUnefVLbHh+pUX7DTChfEv0Jt
MoOlM2wB3cAYEy47FZamrnzTp3JrKk8zEoAm/3qTZXvgFmCDnWn2eEIF6n1ycoSs8jWoAz9ZkVU6
OUumbVnuHxraPLsiqid1nMFX78ZRPl5Le/YrikVrgANqU4ADKVisHEw2knzSUumfeaZO3LwI7kT2
7K2XUUtlxScJP7n9aRRcLSTy4PTURgmTXWRetEYdslr/m+0PTz2a7NaEYci2eJOipT+Cy0aECZwR
unSJbzFWjWez19WvTra+g4lUywH8ZORqetyzluJtNEgify9yY+yrBPMnTGYnk/QYmDC1/bHFb1+1
6f25EHlEk4wTjdAfChmNaNQPZEbpp/lmU2v4LvJp6eDcz2F5RA4iFRXVjH52rDIG5cdFwd3MyRx8
Q0fqXkl4bF5P3vB4usmFj6nomhKK+biTKXCbqI5mX92AVFSdBe5wExnjTLUP9Uy/BQQPAnmT/ZSB
dg4z2Ko4GxQboLu1qlTWW7hmkgjmqti8/WaW145bt011tmYfOQaacJNe3RQdYXuDrDq9yE2DK+KH
tpmuO62u6CFhRrKZ2Wi/eILPdrLSixYqd4ol8RpBfov0IkHhz+5QdkErMJVP0G4RkwmoS+SYJA6Z
wRmaYWSRVN7L+8OPiRae5jzihuPq9pjueI6UY2oMuRR2o1X4rIIGE19nGOLR310ts+8pv82JTfuU
cWM6+2tv6A3wWS6BCgtugMKwE2KB8FshWyQgxEHzxy1qOiIBi9uz6YMuUhkyi66lkVH361JRJPUq
v+D5eEnt4oWdatLYFJUl3FsPW3VwH7dNyikXJKr4X8zRxA+Ry4JjA+t2oxtRNMhm086NTvkxBJrb
n0+UggC3PIWd0DGtAL+lFIFaFaaCmguTvnfWhmOOhcbVvjWa5o+dO4RzrdqMewX2SorEGnE8ZPXT
JsYmkm9j/CwYU95gogl6Ntsb3ebjatdHzrjyqLOpoEVkxvmadSBo6zOAXi7pG7iioKsd537ub1df
SneqM2xo1KvzQW9eQbr1GTZuKOxrEqx6697T0H9AR5XRn9gpoQ/dbFeaexp3bwJye9/9rycEpl1v
57GjdiBMI/NAZuigauBHRWh+/6PuefVUX54wT45yIft5X0h+gbSz8rAERl23xpCNHtGzobkw4aHl
2iYR6Y77pRX/nfZMOhdqinpTEK+a/sI8dLNgW9j/jWAN1PxrMyNtndp/omnE+npG3pdjdXtcce06
r38wzk2zpvz4CxsmVFtTiO3f3vfGt9ehOAiHyiCG0C4JvuIfPTYqi0+pnhylwfz9PvpUHjeKtB9n
XVxkMkm1LKXTGpsItUzlOquTX8juevaUK3Az+s+cb3wlurwxHBXL4uKmUmim/dOTsqvadlzIcKt3
oENiAfLP5uh1uO0BS6IK0tZIljd+glEwHFAYjVU2NNl3w8QQENIyOCU331ukj7DZKD7X+T4OEroT
LElIJyRgNQtjV4e9R0b6AA0J/gO++5Me9cqvgGZO+hd8JuiLBipljYljdqqseHp8VCrpObILLzOP
F/tlLNxQ5pEetGLkn+PRdHIo09+Vk+C2dKQGYvu9dXO4aOj/9p1jGCFfZUD3voN2AOZzRXuzROYL
rA7zRoM9IxWU/ozOeKCiFaI+sCsTVtfvNr5gxNWS5temWt1hQOshWEYirtFJ+mHGKWKL5HcMqcth
YIz84X47192fSvTvSdTEjNOtnT1sVvSfJ8z09QqLWyNOBDT0OPKrdqFD4n+H2FVm2cNZEU0Telb/
M9ryprgar2Omy3EEz50P5pMqBI80G/v577Gc39W8jED5GY+u0/n+nWpba9KGwdqDphpEdDFsCohw
fYx6Le60Vg9FhgdNBdlzdszoe6lU2kQCjP/q46UKlJe6lgGaZljlOP2AWZjFH5L7CKOXygYKbyUd
HXw2n7YU16tm3O/82gkLk8e4tv+8azbvWDPHSxcszCKt/Z2iEY+uQyTTjWyxs/n8FjeWYv9mnd0e
YNU4qCIwaVay61fhijZBG15QIgp9yM1tK7f/lVJYsYRDWHoV5qv/9QgI7WCZWBKVEqMaPRxE2H5v
9ibBYj3nS19DrC9LjrJFlaeespkzmlA+zF12ZeoDF73AIn8vLd1Xv+z4UCvwlKWHVSu7rCp5Qe91
Qmfe+jENYyMC5MT5YRQZbSgOWBAesmVVZITFCBYgLVKFcZLDPDX4i6hcIwyjI4/Ze++emLAPbtQ1
0ZFq5GUgSXpwRGVHp4tct3APo+XYhrGKJXZqBkZVon/JcNIJw7hOYyLBHWnSEtz7uxDykUYGP4w0
+cOGjw5JBpKqdmJrqsDWInEHaBGjSkGGgR9M6MP/ox9sOWXJWs4XgIWRxA3YbO12EoXs4eJZdiVK
hPogkRWoOOTPvVnmEC9Yq+/cYO4VYw4GyNfpiy50MRXLiAf/iBN1xdfkTLseZ3+ENkCAWE/KxigS
+G8stwFYahjyVkoz3ngpfVepsohOr+eni64G53qhb2E3eZVFGYcj+Hc+KMs8dfbY6V7ljTxUOTAT
+1xP8m9BK3+6MYho1xbSSm1GA9+EgjDTBbfs0KqDq3wuCFs/UOgA8N+tDtehjUaLgGa7RFLiuLr+
1d5M3bzyJ4m+aWX/nax0dPzVxWUk3WiSpGBOfdNC0aB8vUx9dVYfMRoCp9myeMTK8Lu0rM092wwe
zg3JFMvXIxPh3I4UgOWFH/SeUs6kk5Oul4BYvnBgkkbdZAg3gHfwMR6E+Gi8ryYKOHKy4pE6PP1Q
3QdC+sqnxMwXT9qIx7GTE0JhmkeoIGmIhB1fLt1gi/D6FOhOB7Aaoatrg2s54SvE6XC8AAoDSKmf
N/PKZkgajNNMJWwZwWul+VSntKSus8fH2qLTBKl6iyvbam5yWlLUuEzSpBh4pLbVFS7+1HSvsc2b
fRRbf2M7k52zC9/Huvd/4xPOMr+3E6+1V/n3Wxysc9Vn5RUq5fHcm/FR4e1S9J9hrBLORGMJcGKu
TJQXrf9wPHTD4Z3kdNrLAE4GulYIMcDLoG1Le1x9GFsTlfJ2CfRyEGx2Sa/krViNMMYAORiLpwFv
ADrmvX6jdsbQJEwSqcLHgLEPqcwiQa5Zr0I6Sa1MwXND9HgZm0ON3OV86SZksGdtVOw1iuZ4EY8s
vbpSwjdNd82MfrLCDQmI0l5c/QrOiq1Sy1qql91U4MyON4mTJratZ9UtzQeJLsgb6bB8ggvdqsUp
P3o6zw0jZrvG/XxaDrzNra8fNZz2o5Usv/CB2yOGx+/kUaTfdCcLgYPZZ4GiKJXotV7aeAbb1d0p
TF+0nXKAwRZorJmqGG5w5tZIlvfHtgJrdznXBmYmDut/PlG2NuJc9X2uYMK47jN+QNNOOuiH/A/n
W73QnPNgWdIKmDSZaJ0IrL8Wgp9IdV7CToGqRNSTkdahdhHEtT4fsHx4Rlx3r9i+oXsEcaR9AZPi
jqHpf8ZWwjWdYASeOPBVnukrAfwdkd+SayqFVidgYfCcJfbtWB8CKtankizeFUmdbAc+FsvwzfwR
4BzTL9Vz6/DG3FqYHSxxsqjm3R52LXhFfJniZPQgJfT3hjVU30WV+Hb26G71FwU/yQ7SEG6XMJxQ
xFS83FuwE9kUkTiF26OjJDqlBPenMJSCvckboEV3gnnZFFcW4AobCBsGGppT2LH3CYZf+K2+hy28
f4uR4B4pv7ttLKJ1x9riOjftEJzUDgZi+oUMJEdJna3kQILVgd4l7T37OTbnQjsd9XHKFeRt7hRt
L1aLssxTsAatF8x2BbK/sZy3bwrWjjwawVXi09KB4dGeFhZB0vGRqJu858T5OyAsCEoOhv/QFRYT
PwYSk4/tJ1pE+Xig0BKBQtmCwTcshIKc1QPI0c7pOvTfpgKd63VBX6mx/w4xvfNXpbFeRQPVIIlA
0wGZxRtMODCrlMPD1PbtI+kfUzrNXx9QDlzinXJAAUHJPHgKaxegEF/GnesJnMRA9M1JpJLtmiXw
GjnErp54kHhwuRLhp5esDe98bBNxOdZVAKNWyqnYRQVJbbCcc+CWBioinyEt+mBG0Eab/z+degje
s6ZWkKipz+f27UEExDxzHQROunXJ6niWuMHy2Thnlrsfmk68n9VCGKYRf3DE1lFVIm4KtXWnTGEO
we8LjzLK9HP7EBVE2mJvpek8nYMVZkJYTJom896RsLtmhCoqpeNI1nnIXEoIinSoA4G4Ol3Du8EV
sF0lQDSOpdepMaR5NRRfqh6Nr243/esOYk9a11fqLerTtLEIkthh4tO0Soep77/TZnEQ0oxrtxgH
n6MLowbPsC9jQExhojn7qdTUcG/7hffmjzAS0tGSV2RnBeX2RdJtDXoByfBgVMAp87KmU/WcQ+QE
N5vdUHxQY6+RUv7BGRF091ftSy0OhDtg6u8mzYxZDCGfEXHO+7Ifl79VJUw3NBsNVD+xiQg5sc7q
/eFip6vPhzghh7gq7jsSEB4ZRgZGLCTcilBqceSta+mMG++DdBUHUYE59Y4Tqaf3z7/NjDx10m/F
BwSuChDvHnWPl1LqHdGeWx3GhitgRxrNo+Wx75QNKF2nb6mdNokzOe2RJY0eGRnXgOKdSYy+/kt/
H8Kh4h6w9d4rzQtbclYuwsEz+ICAWQl2tcZLZ0QfJMq2Cq2AoyTCL0ApP3WU6igHGJMMUN6UYu0N
TnJo8zroMc5KPD2QKI7U5WKLHCdzlaVNDcODXLE+TS8ZRehUupwOABVGJLvDu+Gj+8+s5+t3GeQ4
2qxD0WVYHNZPcWMOS8JqkBOtQuWSPYDNfGRnH3mcZ15waP5F8KXVcW1mBWB50QyiWpLK7BPpVYrJ
sdw1+7TCVt8iBU+pct/3icVLQpI4cAfRn1I/5cmLGjiZBto8CEcyOm11l1nltcHRlIdc4wk8xbzD
xXEkAiIw/yMJW4zMzvyoi2uCMaPjyhd+1jp2+sR2H1HsCTT3D/3Z9eUvyijAVwWKzXe3IAVhvOWD
cYgnvjN/GPgHqKfLIUopPox9nmlYwJqKrUKbMjtU0yyaBb9ePhCto7mSgqw7Al41+U8oBC0mDrP/
PUrhHoDngpazX+JjuiaJsp4ZlOKtBHOUdPiX8BzboCwQsdcTargQO+hpG3b2gfUVH2m+0zVdiI2o
l1hy/IzKu9xpqohK6SBQtjNIz9r/nU6vCEo+O5lwNEzHeQ9Pnnb9QGEMGLV6J3NPxWd5XMPtDbTd
fHeJ2GyltwGQp7nwb1XPRp1+JQpM3sWE64Yph8wuvaX1MJY6QYVY5Jfo0RX33Go+6PG3KFJV7xZV
EkSkJ5f4QGzUuINuuB7B9fawAblmhz6yQAbY4hUzQoCGr826+Wai3G1/PmxLPV0kb/wrT+Kylc4a
8cmF8ObNB3HMG4ce1r8SHt4B4JwpdHzYOEvFA0ETSGuDwBnJMXhjtYmtHilicNm6aa5rmrKEOBEU
WpWsqZgkzHF9CNczkRRw8N+yPkdVFinOrLZWLBA2WsSLtIblLfB+ycXk1o/yiV+Qq9OXEDu+5BRX
dlVcczOdK2CcpwoD/oH810Fdsm0TZuhCVjr0dQsOiQYPJv1Pabr/LnwXEBC9df+4SeyjIUi7DtTS
kl12Slm/jLRMFieXP0bmpJavd06+G7CGXvSgRTNTxgguEhLGe4ew1GXVF/PUYMc7VbsvbaYD311g
jKeBxake2liGDvOC4+JuLkVsIytOhOgGqlY59yv4sC3euTvFYUdhsP+mMpPsFXVTFWAAOGXdGyAK
G9HJzeD7/f72lQCIIzz0Aa9vlWN79RbIvZS6iWQWX4vsguP7iITx/Am680o7q0bJMxrvynWeRxSM
otZK/VoNkDFffLhfdiJKAcQ5RJMWV+LzxyK85+zEAQ83Gd05V9mrpBvFx/+bLlEWQKuAkTzaj76O
74FmorB9MJ7NI48EKu7nugkBYLfLShRxu/zbdphtTikOlV5U9AKGzM8j71rc5z9hd9hXzDzK1QHk
TaFsU6lsh6qLJD4nnwjvH5sfjuri3O2xkNAW12EEncCmFW/yNnuJLlvEmmlxT2U6q1b10c5Qalrk
mNO+AMEiOCXyY4FBx79Wr60iyIRyIqBmVGsIC/AX3Dddd/kbD38IVEM+7A2zQQWh4CP73w6g3eqH
TI6fAl8GygJVkTjsgmpo0tQ9OUonSsquGz6MHU5Oo0ADpviCH5r05vmHIGY1XfmMmGabRKDi54v7
uar8+54de06+EBjacTYkVUIsx6Sjcwx83pImSGhoGhm6D+eJkRygfO5sSqTh5ApmlFTF9dKscluN
Pz+FAqH+2U1GJURDZX/XHlICnqxtRzfCG7AsxTAPIjwt2WPgj4bK/NsSj2yfA8LpnDrADhRzbM27
0ACCmbFzRwIIl7fRRlhC48LNqDU5J6nLl7wSlRTFWyZERBCwpSlXBEeKOYl9H1C/kbgpm/tPbp6h
flSS++x9oij6CA09EPwcUcQw/mA4s7mMF9Pf9baXP6yisN2C8lCi5JV4dfLHJmlplXSYTV8hgwow
v68d7iY1xNmEEGLkZELmSPRJRca3IPubngqMIzaE5nsPweeOXXn6IXQZEyzh6dHA7g3f8Qbssj62
xg4QKaZDxNhjFKQ10SLsRYIJWXr0UZaElGY+zTfQ4mM4JSd0hTyQicbU4FV11NW95X9hW9NIzvaP
TMaAUIUGXVVaDg2smUNSsEoKbmM2AWq/RQpEGNLTY2ECesPt6oOh3UoWyPEsWajqR9F+okzTlGDw
YXFt8+6ifCgXGqeuC2l0mqxQ6XoHQxqANOZXJf/bzC5xFxkafT+Y0gw3uuhWgZYi9M+gcRc49q9I
u5+Gde94QUxHN55vln+xvT3J8hbEYgVSE+QBXqap16Pc5E/QratT3XPbiLGghc6SrMpTT+1f939L
XYcikP9sYw9RmldIJX8gHEUFXrkAmES+LbqB/Fv9ujC53EusSkDIiY0kkr5He5Erw9bRtRgEQAOx
hwGvX9mkgxfYFxf32ogxqVeZM844gWZq4AmDr1vhh+jRwbMdea0BZsnf3Wtf4jT7B3yFSt1gvHK0
G1rTBLd/r9QQbmm2eI6DBqR98ZdlpEErwnDz6skpgCkxBVyVmNUaOOtEL2HeS8VWT4xaaYlFivGk
brfw6ivnyIQYfpleTHAoJk9uPMnM+f1nVLjI/K7s9TtA6nzqfY8W3X6Nu+zcxXyHnNrpwoClaGD5
SLPqB7kZXMtR6twS4JOOYNC6jB/M/7kGyx/A/KniE2hEtDGO8UMfZ41zMHVdSGV7ZtFL0L1tjX9Z
JV2HsnvHUbJpuY7DNgN2/jNk6+HIV0XuyOurSXfD+aRxnSCjjZ2O5+FGNvJGpd4hcdGCFlIUPbJ8
s1c/PPk5Nzcr0m+3C/Ek+QJfB+ckJ+M+Zk5GYJ42pWl9JGovAPeM0BMBDOG/+TNZukC2ZSm9VyMl
t1GU/c/O5CuYadRyia+Am5XkUqJOOcDYZ9Pd7ZVm/ByIuZtuqoc3N1GuqEbJbsfKTcC198Q1QivB
R0jeCWd8TBaY53446flb+PdikifFcqit21DIvo6X6uEhjBCyz4mIs1gYS27eF6qNvw01ufvPNXIE
2D4W/8l8KhmbUvzdVem22vsA5/kYy9ESENhA7nkT4p9EpP32VrX00Dq53YMVm2f+OMOEHLTjrK/c
pHH/qDAgLU1IiVNtSr21xnXtn2udckFFfmYxLX7yiy4touULmiiOaEIIaTLRzvjKOIZTGKsjcCS9
d0PopeWb2MsIKVpsiJterxhvNzxxDlCgWVjH9yNtI3Mgmwup5/v2XWybZbpD0kJqZ9zm90rx8HZN
c5jQ4BGAcHClwNslNZx237Z5h8mPSftb3osqXangWo6MJ8C4sK5kB2kPdQzla8yfs1wMlhN3UG5I
bW+sQjmcAfJB9bPZJRbHchoQUIReyj8GqQ9l2KHF5MdJq/wvUz5KXekdHL7YpVjh30AMfI6vEsCe
KXwkC7/Rva2rgLhLW9MJKzIJMpVVCK1IvLHpUNQEesqkHPV8JXjRQDKESgM52JAadYIabZ2Oi6DI
/gXhFOUXAVAfEmblthWfvdn0ARGgF80AWPINNA9mrfNOm8txR3nUcwjxktMV/dyG1q4ri/S5yEzY
DLryNjBKoEChSKJ4492qfh6SlCNLhVoPyLFnFN4U3c+GF1Ql4XSDwK+bQKzKsaNRrGlimao088rf
aosjyHcLqR5icO3Ie0NXtGHlj7Nz5dacs/Np7jJN+QyHlSgyY9t1VjyZvuHOzE53z+ZB9f9QQJVS
luvjRNMwk3x7fg/5odCiQj5In21bFSAvhhOdcFpEfmL96sS9f0aKNCIq1ABywcvtSXcSWVNmgzRc
BkjHG987RauIWBANn+lqKvf3rXGluBeT8uVz8o2yFidd/yfxBm1GtMjywhdi6PvzkVHsoklSHrk0
lMazz6q7xO/OzuhnJb5hZk27wlIdyGgfEB/VxBTpwBD2Bmz7+gc6HPzJ88UjKu5QWLmJBioMVfan
JcjBOda0gtFTKgw7V6Pxild//lT+CME4+0SjqwJ49KKGHtwxKR4+2IeNirsEVL6RxBkonAX6JH7k
Le8atjkpLnugwi/Fgp1RXoC75IA+1LeD914+Ht7a2ZaJPPGGYrci8dBTcU3AfSBHqDGnj8xVNZUi
jT7qYKC6brsVO3LTBJp7osd4s4jVthaWTRGYvwvDtR85o5tFhYWF5cy+nJlblvvN9t39yqpRFJ1+
7sQatpiadPQXp3xRISHaOz3moZVdkvT1AGEuoC3tWYjq+7OzDyRZ7oVBq2/bmzjAtUuMM20PNg3U
k10l4BjKUUU3DEt4AiySpdArjX8LvblOBTE2/uGRrXn8T8ELhNVTfZDidqY6fsu7VhDIOnqrw6lu
dTUAiXJ/6+fnot4v8rAQr2/8idc2E7KiB6ljBqOhkCCfdC5KQDOp+smqr01CXj8qD3i4LPgrzMpy
Eojn28MY3nhHTGofY5NdmWpZadkBXqNWvz6c0kgkTNyO31pmxDOsbY2PduBWzNahi9i0MbRsvEui
B8LSfy1bbdajD/CRshx81cwrftjZZkXMhPWXifgewfUe0HnYIQzqTgRB1B6fs2uhQS6dyE3wUiek
bmVGsVWCEzzGbFWTyj2IW8oNxVxzmTOM7HX/IJLmhbOO/ZUhLqiePCZYFYtBRQfAFv3MkjU86KuY
v1Y0zCMEkxboUvd5TM+0NwVTxOl0VyyOLd5c3mCC1aMPWaiGJcS3sI0Z4MCvzSMycIUrnS2xmmJ5
7zJSPej8HmBZXFsQYhGN3bnWjpfp8Pfe4rGaWkPkJhpDOsbvIsnrk9Y3dVv31sxxBu7iC5Z3B+r6
d3aabz9BHHoMH6+RpaPYLY5JXEhbLGR9uX1sKTPzxPso4jXEI5KfwxVtI47bzQuMMzE65hcemEa8
Xe0MQCmyBdyTgrlZ+Fx8gqCm5B7KtH1HQWLseEytgUrwkXDMVSVRmpFnEtT4B2lnTV4GkteJGHoi
FrH2HaB8LXDTd4DE9xL+cX4HJRFfjz5Q6n6OMaKYiAUY2B5LJYWYn0KsTZ/dyV6PyMSqeR3AmsGf
5+YtFDhEypY6mV5LFrTuXw2BWbgIKfCgEOClW971CzMdu0OPQqS7L1y/WKVguDjbMoCSwfDBDYVW
6AK5oix6zw2F5oDfG5JZBcQGqQrYoGwdmT1pS01JGoGvqsjAuzdPAGt5gpqpK5MubZyBlT6q8/n2
CyC9VkTtp6tpBC7uu9369MUwcEo7/X6z7WltyPKSffNWjOTb7JE0QFPtqXX/1Cjbwd52dTr5NP5p
E9bpV4RAIXQmj5yZDDuhf/zque/Nbe3dZ2+a0d9Etqto+zeM8IhDtIfcsekB57cEMnimZnZUXON5
ESIk94bq2foOO2hptX4R+8ljInK6zNyAAlIuQoTJfL3DkJJU5UrmNBsqdCuGs61UevsAvHZGgGLi
DVohkybkkH7l+9TI29BFiF+4A0F+PsnA2E/9JZ84N7JRQLWJ1x4srr8B0B/7bJo30ipSAXLxeha/
LB/XP7vYbGr9FJ5zixT1qb6Chth1yCxbOM+FNcGyGM1ZYO8AUEKdkWtpwdpH33cyWI8d1d+bs0Pe
8200Ki6vNOe+XbSxh/1TYyD3qwKe1tLipjzR+fEW0IwR/SBtVxWCuHwelLk65/9m3qL+sbWrW9zs
4HAUkG7CaJZXki0+oHE03aHfA9Zo7eJKEzTP3ZhPyKIp+Hu28s0vFU7Cldmd/Cms1VmEbR03vr9O
u5jWcraecOwwHKk9isBq0auU8uDTFLaK/mc8ju7XwXKmfGuUmtIH8O0gxqpAAX7pI7daNwLRDTIt
LblOLq0f2TY0ev320AYuFlzfUk0Du4k0VqGl9CF3/YGRwCqpo2U9H+3mY9F5nsZPn84UBfsyQV+r
bCfUNqKL0ZkhVf84XtGa+VEkXvTrbS8g1Ru2OVmjq8Y51soCKVNbJaRbX6CKAO8YOtyQQP2Gi0yi
PpCVkW8mwF6DHhxZRVRm99fJqwR6HUiEh2Q8xgYGsEihhjBqV3Ps+qZI0UtP1QgofL9hYBglTrvs
4E9fXrvj+ONgH5xn1dvtSl2pj7ezdwJyHyoK0TYjqVbMTlxR+TtRl/Df08N2gSF8p80Oq8y8+Rvi
GR1QFSYJE1lnCzYqNaJALi92hpwPO5XJ8ObNK8m3kHAKqEIAHKXDhA/pdr7ya0HhABN8DSKaP3xo
e/YleS36Wr8Q7n2pBz+v9bdrzKlCgWoX2EdwpcEQJinnyuqOunAO4uvVEaAHK+PXNvlnWRXAU3aY
ILyY0XHY5wyKOStXF9Z2flT1aFke/gxMxYPoi/eJxJedpKOBUZVPgnMv6eMr8hpNZggkweIJBIu5
H8145gXy8L4J7pXlkFHOPxKTQpoxmpNgSJz6kjLiSY199T3H8kFzpNPLpQZb43VUC7arleJ2xait
ncIFA9dqNUF6wFLk1FKnCzpqB4OpuVi9loBFC6Xw4q5kqd1BarQ+hhICvmiuw+E+f7j3/127FDmN
IyYREkX+hEJiAi2TzH4vQOdROB4lbqaugBdptlLASrBYItG4dCvrgy+lRf9FAJ1veVAkNfkkS22B
LgO2dJTij1yP7IkWpS5aPubl64VI+wqnUVG0jpxCFoa2840irjBR1BVXeLzcba5Ja+TBS4HXCQKF
YphXtTJqIZrBmOffOjHNp4phVlxNtruL36FLnrlJIfNGIb8Uc250T6QLsAjfMfEoXO2q3aWIPoii
bMajw/C/kjgiE6eM+MpUlLoABnIkv5fUID+PvI6+nZedMA/8E93SiosLhN1sWLeBtHYyx/4MOaCi
Tqxa6yXNgWTOOcy3U+7XOXJO8gUbtb0/sCAEdFjlHcLszTRL6l1wJQczSwVO6OovFAkerU+P1FL1
16D6W4FUNZjeEAPdP8e/SzH5bd+Ytc211aLvdZIbJYNP4INVeBMTQZHzAKrs9tBsqceFvNhJc6eO
Su2BMt1j8hVmb54+zgeqS+H3fChR4uYebMkR8NHI5GtU06+QW8HeEhZCCLr+OwEhELC7sK0nNXzi
Byxm9Rc7zRacCwiURZ/BE23oHzSFdUKvTZezwcGNbvvrYtkYQpt72DGwduwrtP655eT1MxRgqz2D
4kyW2Q7+bOL0lJV8uDD9J6Tsehsb8q1R5bsYhmo8BXTTCHPCjyMSaF3ILV2VXIfPHGNbsrjisHq7
UmsUYow+rUZpl305YJU0BA7/y3A1UX156kn47dggjPKwIUeaPGt9lSUJvnlzHo1GIt0+NA7z85b6
s+14xtY7MK4vN2y6HCUnh7kjQW0R6D6EMlgp+SSaOWH4shXAPDArTyrS+yzOBO8h2Thdk27YZjst
PN1Q28WKgycinKubgqkf6kPknMvYT2vc31tlQ6z3WXQQA02k9fdKDKfEI2g1VgGAK9n8911dgrsm
Nv86fC9qC7HhTcPpl5l248IfM+NscQSeMZ+9P7/UVH/A8M6VX0KGJJoAv6F0tbKduOoChoyfrIgo
25DV2/9rkCqK+jOFxRltV2U1QPNvRxAJlT/UAzkHlHHishI5mQpipDW4hheIuY0EVb+PcULPGClS
JrwRcs2LWENEFU5X3uJQEYCFr2ET/NdMSSidXZBXidUAEgwdziM7w6QhGeSpaA2DiQcu9rdiBnlg
lZ32JMvMQ9QtyEgyS9Fyz5Qbtfvicw95HTP2Rtp3REysiAK/7L+PKeqltxzldeGkgJLKeBRZ6pvG
c4RvwzPCSNRJEmRbqfhSE/rpH+C2DESedEJrfcxwGXDxyd05dqt1dkS/fo6vz3yvhdvezaQMAEIn
icRLStyywr5YMw4ZbAzRSAJ8KX3K42WWsGn0mTJgVAgHp1fjjw8dj3AG1+OTf+118C8kKI2tygcq
R9peFPTv9XCa+lxwFEpYb2/xjPYvHgnpJSfL5SlShHPxpuF2Tms4D9ZCcDAC5Zk16rqQ3IXdwSzP
jnYtDdvWN6PyL+A6PFgC8Jbz5cWOyHoHgwQzId6ng7gCb0as+BOFvQpDYAJnhNIPhvtcYhl3hqDh
SRE8YUF7Es+xR64EWFlmca3+spxX9FUflTqOltKWKUmDugd/lyUrS9zdWNQLx8CGEJ8rXE8J8b8a
95riZbh3iiRV20H+ZKxlmF4EoPGxoIksgNi/YkLvZ1LOY6KlhSh4W2P0ZdROeQBdk3DBj8Z0WZgE
H2Po/VOzg13ZPIy8ljKlQlXSKlGP6OEcDCLmQgQ0pvI40PSRJd1SsRlREQBL1gox1qZIs+C1rX5x
ef4DIc1GttpJ6z+41lBgTvgEELyWVuxU6q/AJyQpfdCAFPOs702ctMklV4X2rZmuZiU4A3znwxqI
wvUjpt+QRefQTuH7+s39A1ypqL0cEhg1JJwFn8G2Lais6OoCR/Z29jMwrRAF/YZ1RlwxGJn3+E6V
bNv6mqTAxbpUeOnu7dt+wb4LCncGRmNFCIcHkttGL6q740CG4p4uQOfA6Yl0v8XcWyHlk1yrCaMr
WPf8nYj/MdklQD2tdY2Hpyhej6tdhO/KqvKI4v96cysMteqU/sKmqhP4kTtz4bvDdajxzJHpOv23
ovKks0r29WXGoGs6VNSVmeI4VgufIdN5TtK3iBVjPoYiWaGkwDsww86/xndV5X3iG7AkFN++Gk6k
Ek2erYj4gWS8jxjOuL5DoEdxe7DchvIqJIBoDDYkaZPGjAQOr0BiMPzbwdq9Xqi0HXhQ/E7X9oS4
2/uCjFwJ4CdYakgGgMeqZa+/8hCTluSED6fwmgL22VE0wP8bk6K7UnP/eYc+pVMUn7j+TJ62il24
kVosl2sA3b/X3FZbGyP1ZzNbCGtgAhpy9d3I/mKy4B5OUgGKeYMKqnqjS89eeofjqWNFK/xvvzck
KJs4dmMxL5jpU1BhyBSj/mlIxnCgS0AFF321yucrLY2loD5Jv57RgxtML8/iQEJFJmJOl3GNWOaL
P5V61bR3wkehgOfXYbCllHzNEXBMNTGG0R02J9SmpN43Q44+38yQ1mICQUfNNzQIOu05ofQC4AVS
F46XuKZRbv4yYfSVhs/hwMjrtxh6ISueeSOGilpk8nXhZvR/hJNmo1pq8M76Nu8qSzCw7ER7R2Zi
JjF1jhWvrEAs1/Uz3z2fYMDF1lOcxv4unAc22rwCG5s9zqi56hfKRMDLRdHnOy+5JRBdhU32NsEE
oYJho6Q0uOlYtbWFIoj/xPSsTkxf4tQzPolYmUeYSFjknxUhfhQwloC4xnmGhVSLmOJSkHclr+Zs
PqkfKMD76ipTjspBaAM0DvfdaoVcqrXQZ1m9iMVUfEOAy9/aM886lpK+pbVfDWTRCM1+Aytd1ilK
8L5xEj77vCeHn1xqBW3xn/B6EpIyA+cuhCypPELjCfb+CFg7ErMing3JMsrqqL6AihPlq3QDpiIO
BsL+TPT3Lw8CuVzweHWLOjSRsM3vGOyjvZXVPr1MKx7GBYTzp9rAFxNs7Itl/c3JsBsNVE03cxUC
edLlaeznRJDdTg8I3X3DliI61Rg1gT6XO6tCwb1e9efPEHVu7IsFsUmVoO3d8MWgwb9V/b1U5ZnY
+updFTA6INbqj2Ty7mVVXWUBn3Yu92kzHeT0yUINb81dVxw5FQV6yTs/OVNfcLMy6xt7qdi0WMV/
YhHoWhMO8EQ6Rr824MkqdLkT3XBGOXlXw3MlEVPU9YE26d26GJCnE1xZUweX7T9/hnXvxUQ0yRbS
CSK3zi6qyQfozaZKR1ean3RBug5iqXAqnIrd5cWqAQc6BN1KI9Iy5uIWyGBjriW3+eIGfROoXcYe
R+chRxcvtMwcKaZorvOr6WFB4oiqugU6377v8hGZz7SOxbW0Pb3RyaZr136X3yFgHZ+Ttm01ukV6
XYElu7s5R1hqMG5jOVXtSOHMNRN6lugfpjWGQhmYdc1j9/NHd6ucOpnRmv6zGkr4kkWvMShT8OgV
mDCSj/ouAfDT+ImkW1oPWlCauU/UpXRA3QDp1LIoh+0vO6tt6dZL8khR7+SlDIN5SsgM4aKisLRO
TWIylPue/9Oq4tJk72wG4EIX8uCwXmM1j0yC1lgTXIx+woyPWx3j9DYpPOokUpiMvXAaU/jzRfic
vCWQ+Sz4nV2g/GfWBp8cXYEM6VSDCpL+vNooswpyAOBKkgPxt9dFQ9/NnZNgKmlGRKWz/D/gxX3Y
Ac+Vv3efxRrxpeADIkWxhd9c8DngxcD5Yy5WcIcBpCCGzBiE5qsN6k1YNft5BFudeOsFHnwvi60Y
HG+e1x/09t8BzbnARXGlMIA2sm1QG3/fKLOXtI8Yxenfinm8o37CVQaOXaVqTWsyq5f91W6Cuf+/
fhuCnTPx9wXUwlrWrhnLaAket8Fw3W8NMMVBm9EYqwjPkxxkdmp9sF4EsNuymoAVY86tAnkY9Mnj
lqGjc/Fl2GohJCZm4a7zSXbJ3uHlf4s5ZM8jXqQaaK5G5e+tEGqOwKGZgfXE89R+Hk8xT5+ANukN
lfhm/6WSErWz1hh92LsmgcxcI5JO3hJAJpWrTuTXSCnooVhPWewgG5ru76dMOU1ctXkoSW7QH42/
qou98J25B/XIcrh1P3Q9uIpEp8j4l1xjRROvggWDAPcuK6QErMJPwxJEsZo+Nr02Q0urZ+7+1gwu
/QuDcvAwG3fP7lGNx9AQvZgUiMDwgnP6M+lElMYnZc9D3LMh8yMHlgTqZSzekXpi4LIMi99gH1Wo
JMoepC/SHdgwDabFvb22nUOEgFhSl6PzfQTQ3b7kV8PxB0oMLcnPYN9zObk/g9FXcAZjirbEU5uW
L47C7rt6QsHXz0NPDxMUoQV9zCMH4aP0auMhHOqTyD0pq8/7Imhgn45IWcb9heqy/GMln85QQcUv
4RObzx0aqAvpOlaH7NpFTptQ5NAG7cWQUgLyS28rMytmbkc6iIalrfaXm2n5JRhF6E5P2vd+EiJw
mgMb8AbzdlbYyUFpM8Hosean5J0mhIThJrDR5PK47Ut39SnBu8rEkEKwlxy9K0RyYFCWiOj1jWwB
Z1HrzQnc+awfaqT+yT0fTqnC6S99h4r6uK0i35ZfSqXVCQS//OaUJRx2uXQjYZVcUw6p95SRjaWo
3y0Sol4brvfrO85zgI6cACRd7FBPMjKW/xUcYjaPrWMukB+WIK5uEba2DY/1Fz3b4IuOO8Z9W320
BEqK8/lUBVWPZae4+Sh5uVS16jLZtFnzD2MdIk3nOnUWYoqbG6Ul/HGyinqaVUbfAJYfrP6q3Pxh
zm5CoThaG8SAMqRwU9GfDsYAzhz0y0NyZDLnb58dtqooINLSVyGVYOEri62+xeYg/BBZsiwpjMQh
3nKV+fVmb4jlOq3pYaH/ouNtWh5jJnbvoeBT0n6MHSBajStxZ8KCUrUKvBwILqi8scXyoExWcE+t
4gO9bJv+v34fAZ0SllAAxwnFP4G0NDn36PU3FYQ0sNRmBmEihCkoTNDYwgotNeZaeQiXfppYHEm4
SXc1H1xs4ici4q12AkWyyrvnV3CZNWw+C3DLvviQSaGEY4hP3+NrhfA/GwRHEysVRw25uqo0RI3X
Z4Toqn9ijs1/6Fn1L2fMe73taGlccP4RIVM7rie+buaMrLHiYtNo8nzdqCNXsYW+sgXJUp73xmxA
VtSIxN+YcFYL4qdYCJU2+LE5W/UNcpG2rcFQV8BZIC2exnc9pFWTIAIqTz1APx3aQVt3mz5KdrQu
MZVmAtIiL3OaUZ8A3lN3SBDl7UIRUVXoiKFQP9rge7gwH0VwzVqqouv1cYW3qmOZB24eeZQRqfnB
GA7gzyVd5ZsVQwILoTpEny5wxiloO3pNxw+ke9TWqf7ASgk4klr97x1zOsW51Y0xJgf1YzFzeu+H
Lz3hPgFcnFcb5sr6/r7B67iYukIMbJusdHVfzjdnzoUKeryg3ptOF66vHbiWj/XErSXE4gfJ5NIl
COIdZihhMFQIec+0qP8hGWXZDNJ1ZLhx0nplM0wv3Bou/I9818rtoPBeeCeIYrGR3a/GhN7vOviq
8XUOJjuLWjuhFJ7k1vyL1XV2+FCtnAMktCACFjwrhbnh1eTGMa1drSUBmx/r0pItTgbf7xt+ThfX
xd7MKJ12zBps6+FTn45P60oiSltshtHXcRv9RG+2dnebhMTjpw55ig250DFplYlX0w5EhM7FpJUo
se34gOxHZvyTqAmcHE7lSj0dYU8GU5Ip/cQ7NarWXt/oam/YwDJPNdwf1oPeVu92qMDYOzQSnlG3
HbVhU1vNdkau9p2Py/rOES1/eIYQ09EP+El2bn1b1kfJnltCm/R95Qr06UTW1AH8O06f9XCU+udP
EvwU8dfoGystKkmT3Py+2ng1pASDOSsOwA4mGDwywyFQuUZ1UPvrWsGA04c51LhyVcfFHVor3i0P
kFp4vYUW9B8tvuvUsbZp6PYUfxBSleoYNN+dSDIWMduhHw9uALwcUNlYoGKbcs/Bvn0/TTvQXZtf
giSWwBoNJrZtS+P9FpWHUo8vBb9YRWhgGUnxyc7DgDhQNJKCg52bKQ/AwtEcrcIkWmVPLl/tK3wA
C53X4Wtco7lPkCbhJO1RZclHvck2auatT5cgqTguojXyIaVllxO4tiRjzWlrr05+HOGsHuWKzqK8
BsBB3n4PP0eLx9rbvt1CjrOAqK0sgIiwE2r2qQwKx0ejB9Eek2sNxWoCIh5CEHzZYudeZG2DLabt
FSHk03re7CVHBfvbFP0b+TneZMMZO3DDDuiYzbPVJCZYcu+qpI1CBFYel03xqMqTedD08RDtWZut
kPC9yr4aVxywfgoOmCBxR5Kha6f9ujQ/wp2Lqt6ddxGjkFi5libMdRwvMYywWdNteYH4nnGmg5RO
UkiOTdrKWIuSO6A5rCElt8pZKL98rGqOBkjPSEwbeoOvSOgWAY63/MCNfATcGs1vmdm2O3SjTJ00
uiuSxeD9LKztM812hsM4sphBIDGbrsRMvOKEMeJ9fIKRvH7FCJs41lE4OH7Cjlszp+jfkfQmzFsq
8p3kCA9NJOhhzhLKXdIcC73+/A5Q2tXOamTakb8PpqikeqHXU6gPRg0mMS9Je/4d7AHWqJ/K9AHs
BinYU+vn+fIPwswsf6unVP21aJeQwUR+Js7gi81D/Y760WBUiElBI03a1l1RWKzOlYFQ+TY36w1K
b/t4Bvqwi7Yt/4mRqBsgbjl6SdBMXZMiThpNBK6mwhqpQRSNrSxssxuNhiLzaAnIzjf8nZcExF/4
aufS0FpcBcq0y/7PtgSuvdpjWziTdD51elesS0WG2pWncbn2n+STKuBkzoRBh1Ak/mLuybumfC5Y
jKesAOVM//s/uRmWoWRN6AUNrIVdODLtbGOr4qfBV8UbhbzXFimtUg5A4WY1I8yOtYKnkG6aiWo5
H/Ii/akFPnL+thlGiuoi56BlOS2OCB2ZvBtjRfsmkXIDNhK0ZVBl3Mz0jZXgo6aOO/ba3JdT5Rou
fncJZb2K9b8LhPBARZUtQCnxIJs32LaWUtIRQDIAwaGNMe4jT55hBio5X7VfE9YmAp/Q67YQy5fW
Tmvc24W8XJG6VLiyMHXJknl1MDiJmRJO7I8NfvWZwZxYtkWBDHQkIF4TXQbXGprC5I5paBhX77eS
l2tnsJRDx2nd1tq14wmf+Dw/yw/stx4CEvZycP2iyCCWlLqZGxDStWAcrH/tAcIxge4R3z4xmDan
ES9eAAQMcTAAtMDOkKPvDa9LDbjB4rJoGdFqwow5K+c9b9qJADFvQFmfXDJnxRFsWtF0Qiws+/G5
cpWk1XkbkHo0EsHy7ycHeHrxclyROZHi9PGuKMKUuaQ6oaq4G0JVbmGdAmEP9t1usZ6IS6PdxKfd
1O17chQ66EDpWEKlUJSuy+Cl00QdDkCRnu5F0FGpWP4+6JKoPnnJNqdeJGTlnmytCaU7c+zEHAZV
XvLdKdUPQVQ1qMutFG2VhvzKM+p0ZmFlOIr6IDDacgBDrfa33bbmegwAhttvJu1PY+n1GnpMLak7
tZIT33ZIA9i6tjh6NxDgAmyDEL/ZekjJvzaEwapu/tIxC1BHUJHgCFye6KOvBXQlg4H7fTvOiYr5
JLXqWtA1s4Zp+2ckZFiP4Me0wE8lwiySJQmnK+6NmjQBpAWW4o1iJoYmvrE2Q+8cO5Bs2OJ04t8P
VenklzKle5GLHdNxjH4nAqvVAm9rhcnxeuJY/GC6GudxtMc7SjUvvYeXwsnPeP5bzonbGCWmIKEj
/PUNRkin7ner17/p4h5mk+KxeCBzlsABUOroDx3cqUdkUsNz0gIhwC2Qf511iSraO6+EmalH9eaE
6GWVY0ytcCILAxMNWhcp1lKQaFxMNZ43vfruoZS0phYjcKFemkoXDSvc5IUwfUE3x66jIpSKcq7C
iLvxFa4nDcAP4RqOo+2WzU/nSrF21D5t3CK8Lw7JZa9Vw6a+ygSPZvmixTWmHroanvNWYvpEbDrN
tV3HvdEJltZX7ptyXSKxZ6/moJUymxkuRNwPoHH0AvZeSnh+/z/eoQ5k1rWBshwsohaUlkj4mAA8
WAU7GCDGWuqdGcPc6olHgDr2lfT77RwfLHgus6UIucZh4CscDei8SzVfL7ft9cp4wKFwt9PMQBi8
ObaGZcYF0HZqPB++M2xZ+bF038mbMJT+BpWIjC6KzlZhDaSOWp9WQZuh4aAlnBTbvpjNFmxMklMO
5VjIV2imp+YYWD60npC+5XrOmq7fzHXinkKK6x+ay5MjDPDB8XnvvNPrCXZJr+DMQwqv+QUQELnq
gK5PV30WWghHcK+E6G0pc/P9h8n+hciyqpGV1DAdub/mmGUXnH5uLMMX66jFCi3iGmwAgpS79g3B
jYCr9yhwfUsr7n6BAk1ipTwuCRWU6uaCkBMUw5QpVECoGY+h0A4giCBo5CVzBzFMNDxL4ltMg/wO
7skQ2c4lbyD9dZHwq4bdwk07ohLwYLI3Qdzm4m+GpSPrmB/FMdWiqI1UN2M8nOjatrRd3miIBfKG
qjNbxTMbPuay5Zv0AxVA1Vp/+b24MOEUM1WmvMvePFtBGN36GuiYM+AqHeXTO6l71GEMj5LuYkc5
D6D3RUNtf3whb0Hv79cm7Oq+yDHCJLovDgxfXv96pd8XVryJQZ2tiKFYjLyvdMAmCtO0K3F7FBCD
MJHvz05deGbCIFe0Sxpn+N2RHy7GIONO3FllaVKYyzQcMUivOYIeVPFlSJTexF9n6SIKkQQmjNZq
tRYPmhuiNaIs5/jUAGIM25Gl+MYcdyZF9OrfVepnnzFBewH7EhhVJmHRQdCkT70494ncXN2fsu6J
rdwBnyZA9TCsFJ3lKVQoANgnIw6ogx2zgwWCQToqDlS2h8sUB4W0gipxzi4rYS1CZvOieXJS0sCM
ZjuFy0Nv8+wFC0GB0ZicKoUNs9uyMzOIcrlMOUY1DiM3BMBIl/vMFxmAuD/0GyX81az5CzuTk83h
eS4pgEM+YjSHUEYCpf8TONIpn28liqM2Zs0fpnQoKhRpUCJ7QpHRZH6EyYxbpPMglV23A3DoLht2
+DnE03DjVy1/UTqusRW4M76Tfe/E+HvyFKrU8YdjT7S4wKbwNXtyBhhq7Os8KdnL8lHPaTNHAVUJ
zNf48U+MOhfBKNCzHwtjPVzhEICzruU4K7wvsYU4pGx9vX3Gz6syN0fRFIo/pE6Sz7ge7WJWDNkL
sTdg6VXZ6w0PfQHsvrbyjsczcNHUqez7iM/KcpuB5hbF9nKnRwjZywDaYvlOWgroRclWChr6RXkC
U5isVQW5kOYxb1t4OGmBGziw9d46shRgh+V0kLlJ7a05O16rHKarQ/TzDLlwnqlN+LBLy1KRj9Kg
V3guQRX8RwIOsTFCeXxe0xve4xyYH8w2h1wteZy5iK3ul6lboJDbGM0RT+8hA2PpvU+hQPIiR2ED
bqkA0qWDv+F3xbBVW58UQJtf9nDWGeO/mRG0GWMOfrOIjdtAwuY7+sFRWiqiyDyMA4uf7Ij3PpDd
c72Jcu6TmsD9N7p0W7MpTMzezlaa0ahdS+O2UnOSC9/gGVMCFYoOwE1T6Dz35yDOZSeWrTsmqUhs
XaV74MUbt3pkZFrHTnB9oNZtGKOEvJsGvTaJGR16tl6vfWktFxQ8wmnaLvT2gvdNgsBT6bCSGjpK
4HdlhTd0PyRPM4JjMKQWBFq6gvn7aYaM4MQ+qq/+aXn/8yrqEmkdMD/LzpS5Qryz6WfnZduHBHc7
DGPv3JNH9m/m9KsQRNB05p6K0rVe4Ulucx39CFgUEm+UhgrBvblLxnkZYQYQO2TsFY7MF/xQkbgr
vOTE1L/5dkwg/9T5EqATXgK3TZLnqmro6fNmWGfkbZ0xyL91CfBQDrAGA7aEaVrULf+en8K5tkOq
T4/Fd9dv5fu6RpJW9uCeRlZ/91icAA1yX6f8Hnjlqb5xWwO/DQFVgMLeesuAcvvNeqTg2qzAIR7a
MzWT8qMbj/bZDfKwaBmFEp7tvDJlW5HbX4Q5O/b9SMkk4/f4fQdDrj9ecYOIgbjIfbIDaeXEFqIA
pfaceiUCyam+jkwlhx9677P3of62opsAP6THFA3UMhnFhKDEUOPLyueuK39Z95jcjyNMZrQ8imOk
HoGI32kdFKKt0meDahhZsa4Qe8/rFyXXqaOu03sEs+N5X1WY7Dmq2jEWgIKa3ICx4SIB0fZjvNO/
7GTyvIDBj/urumLTS7wIDMU+bXO3DbWsS40kuypjKDsS1D5wDkYrWPP30j3O3V/EmVLlNIZOIRCb
UZCVka7Ax1nL3wUoDj99OraO+7190Q9jbknk/2+Wzg9WtIng+qE2+ExQHsOJz1z+sOhfhbIxkdFh
zp1nM/y6rLndZ2hwoZZNmXGZnd0LAcBs708YP8s9Sr6Db46IISvGUDncTJrC2osoBJxUa9bgho0S
C6gWVDXtN7DdVR50fRBgB6xd9u2fWVR0udGI13e1XQotWkCEDBX+xhdKbFB+QqBkECRMEaXYDIFj
O2KLO8gVaS5XKRLSVKTeD3bGVf1Cpk9WgR5f2gELwO1IztTLr7zjeYLlW/wQZM/NfoUcZXICPSPd
8pznN+SJa+4W2niYB79qae5xv9mnLOIwoUwcECCu0B2NDARu3gauyQEMIes3IirFy6SUAXMSC+e3
b8Puyv3xD8ha6rnKq/lxTnENspJ4HOorZAXzw6BY6F5G4f2Ks/CVee0Lx/p8D1IZpogIXk2cIreS
I/zZuWrziEGBobRnD/+BLnF4p+zTG8T1VLo0wPI8JcLCLwXArCj2svg1zQqR436TLV9DuTcMXTiF
28tHDVSbmffgO16J5y08DCo1SI8ZGM9uApzjdKw7NE/24XgbtkbjHFE7BwcvNc/Cz5tlmivr+wr1
jkEqwRp5xpAqCHQzKJAGBJoihR7bCEefa0MRssKGFsDQ7CXc3SrDLHLiyyhns0/JjtRTMlVMoHwO
+MigI1aWRLm9NqGCW6JVv9ohxCv1a3TanQnvWs/SRpmTRt15BrzKl8akZXckFcEffV+DsFFMk8F7
odc3rCCIcYaCjnbtl9OIeJV39LStRT6rOPC/EUQsEtFHzOV0egO94Nww+hFfpGgeqYRmPhqTIpve
lMLZSIlLjs0MjVWQT82bFVbg6moz/dDwzN35rYlhABLqXDhGqxyDXKFRwJQgI1TCu3DWJTyVUrz9
tbsswVJJTDBf64KQUv6dtMlJSlK7Jl6CgURCh6ZcXh9kYYxNlu9+WWVV3rr2gjTjwd09HjKCpwWA
5WBEHZhP7ikMSkdtXXnBNyMcBClIvGM+ScaiX+uSYQvv0Uqep5eDYD9DJfDOJ7naNiY9wcWtxrwV
M5asc0OBPpkO2N3ZHSm5om34kJmjW6IRUwm/6BASFZBovAA8vI7+Xbz5solxfTGOd9SDYhseT9gJ
QCudWRcSZiaYWXDDe4t7nMeb1qrEoZugZm9nW6PNDFbDBIslBDm8KBkIe0KunVE5DUw0xDIAKRpP
Kj6JA4/YDOZEV59m4x+Um70EZxkztvmfV1GXU032xGPTxD/mowLRC2o6YH9iHFdbBnZd2OJtA58u
AS54AvkJ/ulei2c88N4Bfl8DHSsXNGU94hxSUuisFwncwW57ENKLorf5Q24443uomp1NhFtW7oeM
tiVllRYr4KbUpRR1RLJg+5AQISqugZcTMPstb4N7CEdD0Rgm97p7QWEPt2dRrSA5xuPOODE1CEMK
03bHFCtIFz2vYe8GY/tS3mLxKkVs/DwUaVQlINm3Or81fKb++YAJ1XHH9RLDA7iFFv3cARaAjRFL
SL0B5d3TxBEipWt/f2wgaWNXLWmJMWpMLbNeC3bkQiFeTRCsjJvYrHUKiL5CYtx5GuegQJmIJQnE
etMSN/ptM05aK/1etAhpB1eD4LQ1mSnW30l/53LBS0TWfMnXoetrBN4RBcGg+qly1vrFBonvSRIC
1gbze3cmyep1OvKzOcIzepz5JC4Z63EyeuPXszIuA8FVDVvxY8nQJ2l9NcHZtSMIPjrt1n/BBy5e
fcx3YgoPAzzl4YO/0kVMnGbOqUV2zGP+heh6RE3/tqFlMEzE+6qymN88Tn75ItCV6VBcAFtyVkHZ
vS19masNB56FsVh162Hsil1nefo+cfx+XUp7xPhu7zmXtyZd6TcRnhLcOrAg4P1+/EBkbktn5ZFK
V42mi5OuIY2tTY+UdUTGmfR0jt4MdZbDGIcI8Fl8LqIdowOSYIz7XDUgE2agRT2awxrEHHtnT/e3
6ZfiDSLqVPn4BnKaYrBIYvphwMf5QPthL/bYt6xUl0OwsuZK/S8Y9DARfIQHBwlBh8swz+IZIOUZ
GtQLLMLxxVxXiqVXsFTIJlGcMZkRjTHYWTj4JBS7V7QpXarXfEA3t59/kAzEuXZId7UlspOPuZJS
EYNm9w8wNRw0xz2oFfZjf9spoXfoc5rm/Gj1Vubac8UAGCNauFwU1QrlqaIMjY4DTr2rUjYxSdAj
Jh+McTKAaRtuHgSUrvBO6p6zVpwJwXdO18k56WRFF9o0zWcPSkSMobZCLhuF3Apcri0Madart6fm
ffpy+PhEqf7cUCa8QVdO4Fj0UFRLPclIQJ/Wg9gZY+s3MdMW0P73+OnoeRclWo7itm4mbeimnaPp
utrfUlxOLjnsIpAtBOxA9j7vGzfwu5e1CITtbx0IGvfZyu9Sw+LdBCpf0s4qV+qJL4vieEwx081w
YyjO1+6M4Gwr7DRRZvMvkYryUurSua+xO4KRJtukaVLcDJq84pW3jvo30/AAGgWr9VqvGICoNXv6
a8Dtg9m8slm4FbQK4vpe2YSECqomLZBNnrU7H6Y3fcqA5TRVR2TQFx43rIzuURE9wkVz0hkY286g
xoWLOe5yvxmob/w6E7928USBDHPWkpfirsWCii/3fgaSDuk31JvCsmCZdhap+p+1p9CD9zpM1/SK
0dYESEtjU4RvSyCn8UDNA8yfmmwCo1gOdA2L1MiD2Bpl/gRpLFB2OP6XPcBCxnVT3ihYxAIjuX5Z
yieMS5C62JjEMdIsRKgkphvlr527p9xCM4NYDmeFX73u6Jz57fLraBqqHuLnpiQGcW5/orRRYAsQ
eFC2Z6tg3aXCAl1y2C/BUbKvyBru1ojISAFUcnYaXrkv2g+cSORU1q/nbjcbTMfOcbOj1gNLI929
D06oWjfJEa+oERguDDpyN9Q7CjxqwC1GhzzNbtWkQ3fcgpfc1FFtTziIW2Nro6eZGQXP57JBSZh/
IKTEaHawcBmRYPIT2Ec6ppGmfCrKPxtP3vrgZnIO29xWITzGEy7KBRwunWza0dtEB+YcwcGz3Sdl
bdPZyCojrYzp90zXCASHvUYd9cpOc8wrzkIoV3G28IgpYRG9zG3Upf/6d18g8rv0AakuO8cRzxtA
lAETpjhe5Z89DdFIoD2+/JcLrh+Z0A++seJAXz2Zjk1n24rgyHiKyq7irsT6njNep5LsSgtFa4Bg
qeZQ6tjCS6PdfWdjNCnfxbbxtKsjfmCrka65X3bl/B8srUfB68LU/QYhB/olJCae2DBUwEKmxRsc
poHAhgXZA5xljI8ZJ2qvUOSzLX6rbNpTkMbQRMU6aNPQBB/Q9yeBWuh8Ws6SMyGZuFmBu2RyxbYl
A4ap8HSK+Vtb1lJnbefsonsZvPQokpyRJcKczUB+X8BFUxSraz+4ORDbP0aShqwKvaHaA0UbbkvP
SwbzVM+vrC+PzMJbyUc4uYAQReGJfaQWhxdCo0CzMbdWNCKplUWkNGS8hIChX90j2xYlJ2HNEPpa
kXgdxUxgY+QgK8GvVXiZOCjwsJWJn96+O9ntkoff1BeTZVgRlDL6rIMQAWtegzTcSXKtwNnnF6dU
UV3ECMGj8uuZkjZatfwsO+6+5yAccBmkmj6CZ7j239cqhecMJW4YwZcvXSe+X4F1yI0iX120jijb
grptVyyIIEzMBPD4ZXPG7dZQyZ96nM8RHcJtJUFJwXr1GwMzhGtv9aIkNqnIwq9n/QiLIb6+FHRa
wyivyD/47YkbXphl9MNPiI4VAICcfhBxmZ6b0J0AishlUsvP42PCUCUeUEmchJ4RvSZ3mzFPjXs1
7428byTe8yt7YiDbG9jqXikjWaAX5oLU4eSW05UPzVSX+BszfPouC33kmK668fk8uII6oKYbSvGU
f3uYTpg5AgzTM6UDE2mr1IzhKXBREok2LyJ+bzA8Ees/UZqx+5Ypa0a/u+fc6BOrkDkP69pFLJ1Q
+O2U3TZST2y89h/ynSBemyqXPnHwVXsaEP63Ho12oEH5v6wDnKf5go1F99xvVKVVDOL25MAjxiZ0
mAR70ElCnf791oG/YV3UaCNKdJ+OihDvUKwA4OKDGgONG4xraYD0WHyF91kCqbyErq0N/qRyMjib
WDmxcQ8lbN6tblcI8t2Qf5CB5tX+oCYMXPX8KDHYT5yYFRrnWTA46nhkLAiv8+nwLfvNg2390Ud/
bPd7WxPMLuicVP+ts3DWVP22ly3coB/xCkrJvYfbwTXDuc3KyoCiUESOZsKiCwa7xndkz3H00XtK
0TPuDkAPUjVyGBPX1tb/3+F8GnOlm0WBwhg3WHTyR26z8gkprXofjRIwgHTQkx9WuvWn3R3LoTAe
yMzpvKJr+tBkxLb0oQhqRfQrm+ySDyzbmlXvHBaUA0ezl1YDLYjxc2LcWlBjaa8qovml6o7GpiK2
R2eA8PBHG1Z3n1ycBJ5TZ/eJHoW6Le8YsirnUh6ijy8bs+LtkRTRxaFdoXsbdOYTHSl+ng8uRCb5
6ARcanxjBiCZMJXACpknu/+Kty1jz6yk9pcVOS29ri4r/QCXmhF9NLQploIyBKBv6lD3W7ndRMj+
4931Iy9h1KMTj/mx6VjjSNIv6LN+VE3hASARrh5I2ItJrK16YiVYQux4qJK6izf2VTPx4IG/GJc1
NsU/0ca8t1qdg7rNPKD4LXlJnCt6I/DlwYzi8+7cuV8SrF74hRRSTfU4UpCsrUesynxU+LWzcdyW
IO7B3YmO2V6yMabDCBqjQMmSkPWlyQT/zUtKwnKqP5VQy3kVXVsnnMs7mHCnUHKYKDvxQpqZJoI1
oQi98DZfhz88YDtTVaZ2sTMKu9NfMpODdZbQ/Z6Vv4ftgp/3G26fnZx2wAkmu/D5Ln9o9sVQxPEL
yUTDpSRs9Mt6KGRnEa7HjVsyW11WhZFlG9UGmdYEjXb2iOcTsFZRPtA69BPu2hlqtSm1Oo5weUl8
gUk+LY2BD1VxJEpq32odIg0WNZH77I9GiGdDKdx8AszxF2DRJoznO+yKiZTnWtKEIFT5NHJSGaQT
MNRgbTuNJv/lUR6gM8L3BwqHX+9SLDVNFswnSD87qd7vJWpRdt8izJfjMWobiZTzOTjQd+Cc7D3Q
NqmYlQoyCbR/vovomghrhdewpRolbfB5d6+5R5+CLhxgE1TeOB4XQqbSWrAMdTMEXNI0jUum/hZV
dseZdR9IumVoF9M1X4urvYfpFjSprdV0XSNLDVadu1Bj4f8ehCWgX2WHGSTa4UOiBvi7FpSgalcl
kaBtg4G6IlEvQZBdwcnzaSuDe5dpEbxdV+YGBbBkkfF/61oAixrFXQiBDzCIHXbir0WnSOsJjKmE
n5ylAgB8aJxk37A9DSGeiN9QWXJm4d+pi6Nf8J3kNJPSRjtSTo8Py79LE205BG8UQtPyIU9Vdbvf
FHVJn/vfTGFuPk6yzO1NdpxB697Wnguynb6hNL/aD45vm5CEey1Qq6PL2Uh++KQuDlkHqm49I8k3
zseh29mvFoUMssU59XyvK3s9K4EQZ4GocDUMgEZKiz478spe6jgY18epQ2PYj5CSc4oj2ljSD0n2
c5VsNeFo6G6wg2N6u3ClDINTzuyb9PgRnk3RfKisUk2lZHxlCMNUoTkgZgdik+R2aaKZzyYHWmJt
+bvWo1LBym0YCABIHcPetA0cu/ilOTeHnk380sgW6vEMmavZRrVGjLA6mEpuQ8jLL6efhi41MiLH
PkmB346A//aTw28uYurl1EgWYMS7ibYlYMt2I3i9VpJ/OnK3wpZfP4yAjXJn6JT3QVeJ1NOpFZ2G
kO5Yko1bH0MYUnKZ+vmit0JJQUfRaBVUoHkzRZHknjajEa+g1Ays52twbtInxOxos2DRxCSKWlzn
Yfqk9FQAo3No74c0B5uD5S73oKDfePUy4O16gx8UnWsMP/O16jCg50LvU6cyVz6wKcpjj8hzX7n9
HCF6a9SKS/6VqiUwyxsPXa9TaxJohKuptzoGg0LGG5Mr2ZYXLHtTqPYCrZA6FxmnGyLSCE/0nWqI
QSGB1kI5D6WHCw59hPkoAyFWbHduzNCAJW8rLTfNS7hLMTc+9oMKtVAkwU3koLFE1eM2b7OWKVIe
ZHc1aU9vf8zpYwCo50Hejc2rUCvZbGdtTe9xtlfpestgnE8kTLlx9DHQEOj17l/Rgfgc/qkI8axg
wGiesvJxplmigUNyk5UdaCLZPXCC0dWuwQgnN44EnHlkNolMafm1pFYdYgTxcxx9h6mSjb8DgAdQ
e3v0Cc/CtMWTZ+GKMPpWgiO+J4xxgl6v9mSmJwOgUhcRDxNMfmkpvNgKBmDooDVRk0rTQfF6IJL9
D8+lPwGnxXNZk8OWICBNzV6JnPckGRP4om77SVrgKCovgZlDgUpt6FQhKSJB92yNqJkkQYsoxMDg
WqT5oAtF4uPB0pKB06mZx0sa0Y6wcEi4NHAJP8qD/5mLDMwMSYahP+DvwKztGQCZRhTRPOAvMXNM
ioHhQ6yURX/jAp7Cr3h1Fe8ppbjrBb6ou7WIZIDnWjHeQhY25oSyrjUGM84VnNmSgie3258wK7h1
4JVD9HpAxo97RPz0bf8v8KMU2eGCVFHRdn9Vw2BxJ06EE6DI4b6GhK0mKibDTPOKMtZbFhC/x9P+
KSbuSstSrfuF1FOxGfU3okeigWfUvfZ2gzn/TVy10Yu6c4h0vp+vZrnl/QoWpQbK1QIq8YfZGAf0
qEmMIXPP/ab+AGzsNh6KdhL92RFVk0cNxmI1lSYc5yGLwR+BOQdRW+l6gkJG7m1XaFciQ15N5Hv1
kgShlmjUSs7BZObVEu6sttzB5ra/L2HTXs0N47juflbqDBguvLLm2qgFVy5J+W91Aayondz+Cgjo
Gl4Gx4QL+l57cLBSmcEWN+1I2m1A8v9r0pf9TTinxIE9lyqEe6G61wjqVsCCc7Ja7U4a1bGRNJ6C
D4aSqI5WwK/Qo3STFTHsnu1Wos9jb4pawx5nQXY1/7Cr+lOULj5S+D2cWw1vBj3QoChQZeXixD6w
f80tHwmFJHGfwxRiuA4FVNAqjYclB//RHu2lDxfHlDksxFzaEk2WysnteH39rCea09+TyN06QG5i
gdtLaUDX8TDlmyBSYuK+Nr7wyfTXatIKdOYF6yRxnxNn0JluRZjkEgnzVlSoDZjC+uNFqaFL3Wx/
Rns7fpwP8L+ykK0BTcoen3zY7GudUdmkvClEkATMigIdrqWqViIKGXQHVghfsoaCpOKu5ytVz9NP
ktTo0GJ6xxS0vwTvYEXizuBmc7GN0xqSlNt0GM91ft6ll/mfnmazR/V5kl7u/Re8DzQVBfrp5HXk
tUSkdHKzczwUUGFm9LI4k0Ahh0VMwyt+I++EbQ+Jgwm8rC9gyEY1n6rl/abD1uZJG1LnM2p2c6w7
Emld6ENUg4ijsdsG0rxvI/8Q3zNwwOhWhtugMM6DtpUe0+xL+f4ULex9LQSCtThkd/Ybb3elhtD0
7V2eOw/yHD7tDLE2Tf7Ysac2nQ4GUn5ndP0pzDcrsDSC+cYRHwLiQ2cZjucVW01zxBvxiXmI9A3z
6K7RFXWxc1FWumBhNFu1UkiWcXmnzPTgZrVxyhnywQexopSlesomGs0aWiFtGkIzE392PFCEFkV6
7OaHEdj8ZkIHNYQpYlEXJS8pDU6eCCUAR4bBgSzZ+cMGZFfB6PYTahGRdkGIKqKEOyogC3SFdkpv
gfRB8KjAPEUyfuTt1cUNCREPyXMWO14zK78tleKsmXWlvtN3WmRlqg3zBTqajwW8vqyrmX9uUo4i
CrJvJA143l2gpD+kWV28Xp4Y/74R7FwGWVyCRUJxPOeeKkBxvJtIguYO8s6wd5iVo2qQNao6z1Hp
`protect end_protected
